magic
tech sky130A
timestamp 1749382696
<< nwell >>
rect 2545 1880 5285 2950
<< pwell >>
rect 11240 8880 11460 8943
rect 11570 8880 11970 8960
rect 12080 8875 12600 8935
rect 10955 8550 11100 8580
rect 10490 8230 10710 8293
rect 10820 8230 11100 8550
rect 11220 8175 12580 8575
rect 18455 8550 18600 8580
rect 12895 7940 14145 8240
rect 17990 8230 18210 8293
rect 18320 8230 18600 8550
rect 18720 8175 20080 8575
rect 20390 7940 21640 8240
rect 9680 7520 10930 7620
rect 11220 7495 12580 7895
rect 12895 7520 14145 7620
rect 17180 7520 18430 7620
rect 18720 7495 20080 7895
rect 20390 7520 21640 7620
rect 9680 7020 10930 7170
rect 11275 6980 12525 7130
rect 12895 7020 14145 7170
rect 17180 7020 18430 7170
rect 18775 6980 20025 7130
rect 20390 7020 21640 7170
rect 20490 6705 20860 6855
rect 11030 6515 11730 6665
rect 11770 6515 12030 6665
rect 12070 6515 12770 6665
rect 18530 6515 19230 6665
rect 19270 6515 19530 6665
rect 19570 6515 20270 6665
rect 20395 6370 20655 6520
rect 20695 6370 20955 6520
rect 9665 6005 10905 6285
rect 11205 5935 12620 6185
rect 12895 6005 14135 6285
rect 18705 5975 20120 6225
rect 20545 6030 20805 6180
rect 11240 4340 11460 4403
rect 11570 4340 11970 4420
rect 12080 4335 12600 4395
rect 11250 4105 12500 4155
rect 11195 3800 11895 3850
rect 11935 3800 12635 3850
rect 10155 2985 10855 3585
rect 11220 3175 12580 3575
rect 12945 2985 13645 3585
rect 25955 3550 26100 3580
rect 25490 3230 25710 3293
rect 25820 3230 26100 3550
rect 26220 3175 27580 3575
rect 27890 2940 29140 3240
rect 10155 2455 10855 2655
rect 11220 2495 12580 2895
rect 12945 2455 13645 2655
rect 24680 2520 25930 2620
rect 26220 2495 27580 2895
rect 27890 2520 29140 2620
rect 10155 1965 10855 2265
rect 11275 1980 12525 2130
rect 12945 1965 13645 2265
rect 24680 2020 25930 2170
rect 26275 1980 27525 2130
rect 27890 2020 29140 2170
rect -45 1685 130 1725
rect 27990 1705 28360 1855
rect 3165 1615 3805 1665
rect 4205 1615 4845 1665
rect 2835 1205 3955 1455
rect 4055 1205 5175 1455
rect 2945 975 5065 1075
rect 10155 955 10795 1655
rect 11030 1515 11730 1665
rect 11770 1515 12030 1665
rect 12070 1515 12770 1665
rect 11205 935 12620 1185
rect 13005 955 13645 1655
rect 26030 1515 26730 1665
rect 26770 1515 27030 1665
rect 27070 1515 27770 1665
rect 27895 1370 28155 1520
rect 28195 1370 28455 1520
rect 26205 975 27620 1225
rect 28045 1030 28305 1180
rect 2995 780 5015 880
rect 11260 645 11530 745
rect 11880 700 12580 750
rect 10955 -1450 11100 -1420
rect 10490 -1770 10710 -1707
rect 10820 -1770 11100 -1450
rect 11220 -1825 12580 -1425
rect 11220 -2505 12580 -2105
rect 12895 -2315 14145 -2015
rect 12895 -2545 14145 -2445
rect 11275 -3020 12525 -2870
rect 12895 -2885 14145 -2735
rect 12895 -3295 14135 -3015
rect 11030 -3485 11730 -3335
rect 11770 -3485 12030 -3335
rect 12070 -3485 12770 -3335
rect 11205 -4065 12620 -3815
<< nmos >>
rect 11280 8880 11300 8943
rect 11340 8880 11360 8943
rect 11400 8880 11420 8943
rect 11610 8880 11630 8960
rect 11670 8880 11690 8960
rect 11730 8880 11750 8960
rect 11790 8880 11810 8960
rect 11850 8880 11870 8960
rect 11910 8880 11930 8960
rect 12120 8875 12140 8935
rect 12180 8875 12200 8935
rect 12240 8875 12260 8935
rect 12300 8875 12320 8935
rect 12360 8875 12380 8935
rect 12420 8875 12440 8935
rect 12480 8875 12500 8935
rect 12540 8875 12560 8935
rect 10530 8230 10550 8293
rect 10590 8230 10610 8293
rect 10650 8230 10670 8293
rect 10860 8230 10880 8550
rect 10920 8230 10940 8550
rect 10980 8230 11000 8580
rect 11040 8230 11060 8580
rect 11260 8175 11280 8575
rect 11320 8175 11340 8575
rect 11380 8175 11400 8575
rect 11440 8175 11460 8575
rect 11500 8175 11520 8575
rect 11560 8175 11580 8575
rect 11620 8175 11640 8575
rect 11680 8175 11700 8575
rect 11740 8175 11760 8575
rect 11800 8175 11820 8575
rect 11860 8175 11880 8575
rect 11920 8175 11940 8575
rect 11980 8175 12000 8575
rect 12040 8175 12060 8575
rect 12100 8175 12120 8575
rect 12160 8175 12180 8575
rect 12220 8175 12240 8575
rect 12280 8175 12300 8575
rect 12340 8175 12360 8575
rect 12400 8175 12420 8575
rect 12460 8175 12480 8575
rect 12520 8175 12540 8575
rect 12935 7940 12950 8240
rect 12990 7940 13005 8240
rect 13045 7940 13060 8240
rect 13100 7940 13115 8240
rect 13155 7940 13170 8240
rect 13210 7940 13225 8240
rect 13265 7940 13280 8240
rect 13320 7940 13335 8240
rect 13375 7940 13390 8240
rect 13430 7940 13445 8240
rect 13485 7940 13500 8240
rect 13540 7940 13555 8240
rect 13595 7940 13610 8240
rect 13650 7940 13665 8240
rect 13705 7940 13720 8240
rect 13760 7940 13775 8240
rect 13815 7940 13830 8240
rect 13870 7940 13885 8240
rect 13925 7940 13940 8240
rect 13980 7940 13995 8240
rect 14035 7940 14050 8240
rect 14090 7940 14105 8240
rect 18030 8230 18050 8293
rect 18090 8230 18110 8293
rect 18150 8230 18170 8293
rect 18360 8230 18380 8550
rect 18420 8230 18440 8550
rect 18480 8230 18500 8580
rect 18540 8230 18560 8580
rect 18760 8175 18780 8575
rect 18820 8175 18840 8575
rect 18880 8175 18900 8575
rect 18940 8175 18960 8575
rect 19000 8175 19020 8575
rect 19060 8175 19080 8575
rect 19120 8175 19140 8575
rect 19180 8175 19200 8575
rect 19240 8175 19260 8575
rect 19300 8175 19320 8575
rect 19360 8175 19380 8575
rect 19420 8175 19440 8575
rect 19480 8175 19500 8575
rect 19540 8175 19560 8575
rect 19600 8175 19620 8575
rect 19660 8175 19680 8575
rect 19720 8175 19740 8575
rect 19780 8175 19800 8575
rect 19840 8175 19860 8575
rect 19900 8175 19920 8575
rect 19960 8175 19980 8575
rect 20020 8175 20040 8575
rect 9720 7520 9735 7620
rect 9775 7520 9790 7620
rect 9830 7520 9845 7620
rect 9885 7520 9900 7620
rect 9940 7520 9955 7620
rect 9995 7520 10010 7620
rect 10050 7520 10065 7620
rect 10105 7520 10120 7620
rect 10160 7520 10175 7620
rect 10215 7520 10230 7620
rect 10270 7520 10285 7620
rect 10325 7520 10340 7620
rect 10380 7520 10395 7620
rect 10435 7520 10450 7620
rect 10490 7520 10505 7620
rect 10545 7520 10560 7620
rect 10600 7520 10615 7620
rect 10655 7520 10670 7620
rect 10710 7520 10725 7620
rect 10765 7520 10780 7620
rect 10820 7520 10835 7620
rect 10875 7520 10890 7620
rect 11260 7495 11280 7895
rect 11320 7495 11340 7895
rect 11380 7495 11400 7895
rect 11440 7495 11460 7895
rect 11500 7495 11520 7895
rect 11560 7495 11580 7895
rect 11620 7495 11640 7895
rect 11680 7495 11700 7895
rect 11740 7495 11760 7895
rect 11800 7495 11820 7895
rect 11860 7495 11880 7895
rect 11920 7495 11940 7895
rect 11980 7495 12000 7895
rect 12040 7495 12060 7895
rect 12100 7495 12120 7895
rect 12160 7495 12180 7895
rect 12220 7495 12240 7895
rect 12280 7495 12300 7895
rect 12340 7495 12360 7895
rect 12400 7495 12420 7895
rect 12460 7495 12480 7895
rect 12520 7495 12540 7895
rect 20430 7940 20445 8240
rect 20485 7940 20500 8240
rect 20540 7940 20555 8240
rect 20595 7940 20610 8240
rect 20650 7940 20665 8240
rect 20705 7940 20720 8240
rect 20760 7940 20775 8240
rect 20815 7940 20830 8240
rect 20870 7940 20885 8240
rect 20925 7940 20940 8240
rect 20980 7940 20995 8240
rect 21035 7940 21050 8240
rect 21090 7940 21105 8240
rect 21145 7940 21160 8240
rect 21200 7940 21215 8240
rect 21255 7940 21270 8240
rect 21310 7940 21325 8240
rect 21365 7940 21380 8240
rect 21420 7940 21435 8240
rect 21475 7940 21490 8240
rect 21530 7940 21545 8240
rect 21585 7940 21600 8240
rect 12935 7520 12950 7620
rect 12990 7520 13005 7620
rect 13045 7520 13060 7620
rect 13100 7520 13115 7620
rect 13155 7520 13170 7620
rect 13210 7520 13225 7620
rect 13265 7520 13280 7620
rect 13320 7520 13335 7620
rect 13375 7520 13390 7620
rect 13430 7520 13445 7620
rect 13485 7520 13500 7620
rect 13540 7520 13555 7620
rect 13595 7520 13610 7620
rect 13650 7520 13665 7620
rect 13705 7520 13720 7620
rect 13760 7520 13775 7620
rect 13815 7520 13830 7620
rect 13870 7520 13885 7620
rect 13925 7520 13940 7620
rect 13980 7520 13995 7620
rect 14035 7520 14050 7620
rect 14090 7520 14105 7620
rect 17220 7520 17235 7620
rect 17275 7520 17290 7620
rect 17330 7520 17345 7620
rect 17385 7520 17400 7620
rect 17440 7520 17455 7620
rect 17495 7520 17510 7620
rect 17550 7520 17565 7620
rect 17605 7520 17620 7620
rect 17660 7520 17675 7620
rect 17715 7520 17730 7620
rect 17770 7520 17785 7620
rect 17825 7520 17840 7620
rect 17880 7520 17895 7620
rect 17935 7520 17950 7620
rect 17990 7520 18005 7620
rect 18045 7520 18060 7620
rect 18100 7520 18115 7620
rect 18155 7520 18170 7620
rect 18210 7520 18225 7620
rect 18265 7520 18280 7620
rect 18320 7520 18335 7620
rect 18375 7520 18390 7620
rect 18760 7495 18780 7895
rect 18820 7495 18840 7895
rect 18880 7495 18900 7895
rect 18940 7495 18960 7895
rect 19000 7495 19020 7895
rect 19060 7495 19080 7895
rect 19120 7495 19140 7895
rect 19180 7495 19200 7895
rect 19240 7495 19260 7895
rect 19300 7495 19320 7895
rect 19360 7495 19380 7895
rect 19420 7495 19440 7895
rect 19480 7495 19500 7895
rect 19540 7495 19560 7895
rect 19600 7495 19620 7895
rect 19660 7495 19680 7895
rect 19720 7495 19740 7895
rect 19780 7495 19800 7895
rect 19840 7495 19860 7895
rect 19900 7495 19920 7895
rect 19960 7495 19980 7895
rect 20020 7495 20040 7895
rect 20430 7520 20445 7620
rect 20485 7520 20500 7620
rect 20540 7520 20555 7620
rect 20595 7520 20610 7620
rect 20650 7520 20665 7620
rect 20705 7520 20720 7620
rect 20760 7520 20775 7620
rect 20815 7520 20830 7620
rect 20870 7520 20885 7620
rect 20925 7520 20940 7620
rect 20980 7520 20995 7620
rect 21035 7520 21050 7620
rect 21090 7520 21105 7620
rect 21145 7520 21160 7620
rect 21200 7520 21215 7620
rect 21255 7520 21270 7620
rect 21310 7520 21325 7620
rect 21365 7520 21380 7620
rect 21420 7520 21435 7620
rect 21475 7520 21490 7620
rect 21530 7520 21545 7620
rect 21585 7520 21600 7620
rect 9720 7020 9735 7170
rect 9775 7020 9790 7170
rect 9830 7020 9845 7170
rect 9885 7020 9900 7170
rect 9940 7020 9955 7170
rect 9995 7020 10010 7170
rect 10050 7020 10065 7170
rect 10105 7020 10120 7170
rect 10160 7020 10175 7170
rect 10215 7020 10230 7170
rect 10270 7020 10285 7170
rect 10325 7020 10340 7170
rect 10380 7020 10395 7170
rect 10435 7020 10450 7170
rect 10490 7020 10505 7170
rect 10545 7020 10560 7170
rect 10600 7020 10615 7170
rect 10655 7020 10670 7170
rect 10710 7020 10725 7170
rect 10765 7020 10780 7170
rect 10820 7020 10835 7170
rect 10875 7020 10890 7170
rect 11315 6980 11330 7130
rect 11370 6980 11385 7130
rect 11425 6980 11440 7130
rect 11480 6980 11495 7130
rect 11535 6980 11550 7130
rect 11590 6980 11605 7130
rect 11645 6980 11660 7130
rect 11700 6980 11715 7130
rect 11755 6980 11770 7130
rect 11810 6980 11825 7130
rect 11865 6980 11880 7130
rect 11920 6980 11935 7130
rect 11975 6980 11990 7130
rect 12030 6980 12045 7130
rect 12085 6980 12100 7130
rect 12140 6980 12155 7130
rect 12195 6980 12210 7130
rect 12250 6980 12265 7130
rect 12305 6980 12320 7130
rect 12360 6980 12375 7130
rect 12415 6980 12430 7130
rect 12470 6980 12485 7130
rect 12935 7020 12950 7170
rect 12990 7020 13005 7170
rect 13045 7020 13060 7170
rect 13100 7020 13115 7170
rect 13155 7020 13170 7170
rect 13210 7020 13225 7170
rect 13265 7020 13280 7170
rect 13320 7020 13335 7170
rect 13375 7020 13390 7170
rect 13430 7020 13445 7170
rect 13485 7020 13500 7170
rect 13540 7020 13555 7170
rect 13595 7020 13610 7170
rect 13650 7020 13665 7170
rect 13705 7020 13720 7170
rect 13760 7020 13775 7170
rect 13815 7020 13830 7170
rect 13870 7020 13885 7170
rect 13925 7020 13940 7170
rect 13980 7020 13995 7170
rect 14035 7020 14050 7170
rect 14090 7020 14105 7170
rect 17220 7020 17235 7170
rect 17275 7020 17290 7170
rect 17330 7020 17345 7170
rect 17385 7020 17400 7170
rect 17440 7020 17455 7170
rect 17495 7020 17510 7170
rect 17550 7020 17565 7170
rect 17605 7020 17620 7170
rect 17660 7020 17675 7170
rect 17715 7020 17730 7170
rect 17770 7020 17785 7170
rect 17825 7020 17840 7170
rect 17880 7020 17895 7170
rect 17935 7020 17950 7170
rect 17990 7020 18005 7170
rect 18045 7020 18060 7170
rect 18100 7020 18115 7170
rect 18155 7020 18170 7170
rect 18210 7020 18225 7170
rect 18265 7020 18280 7170
rect 18320 7020 18335 7170
rect 18375 7020 18390 7170
rect 18815 6980 18830 7130
rect 18870 6980 18885 7130
rect 18925 6980 18940 7130
rect 18980 6980 18995 7130
rect 19035 6980 19050 7130
rect 19090 6980 19105 7130
rect 19145 6980 19160 7130
rect 19200 6980 19215 7130
rect 19255 6980 19270 7130
rect 19310 6980 19325 7130
rect 19365 6980 19380 7130
rect 19420 6980 19435 7130
rect 19475 6980 19490 7130
rect 19530 6980 19545 7130
rect 19585 6980 19600 7130
rect 19640 6980 19655 7130
rect 19695 6980 19710 7130
rect 19750 6980 19765 7130
rect 19805 6980 19820 7130
rect 19860 6980 19875 7130
rect 19915 6980 19930 7130
rect 19970 6980 19985 7130
rect 20430 7020 20445 7170
rect 20485 7020 20500 7170
rect 20540 7020 20555 7170
rect 20595 7020 20610 7170
rect 20650 7020 20665 7170
rect 20705 7020 20720 7170
rect 20760 7020 20775 7170
rect 20815 7020 20830 7170
rect 20870 7020 20885 7170
rect 20925 7020 20940 7170
rect 20980 7020 20995 7170
rect 21035 7020 21050 7170
rect 21090 7020 21105 7170
rect 21145 7020 21160 7170
rect 21200 7020 21215 7170
rect 21255 7020 21270 7170
rect 21310 7020 21325 7170
rect 21365 7020 21380 7170
rect 21420 7020 21435 7170
rect 21475 7020 21490 7170
rect 21530 7020 21545 7170
rect 21585 7020 21600 7170
rect 20530 6705 20545 6855
rect 20585 6705 20600 6855
rect 20640 6705 20655 6855
rect 20695 6705 20710 6855
rect 20750 6705 20765 6855
rect 20805 6705 20820 6855
rect 11070 6515 11085 6665
rect 11125 6515 11140 6665
rect 11180 6515 11195 6665
rect 11235 6515 11250 6665
rect 11290 6515 11305 6665
rect 11345 6515 11360 6665
rect 11400 6515 11415 6665
rect 11455 6515 11470 6665
rect 11510 6515 11525 6665
rect 11565 6515 11580 6665
rect 11620 6515 11635 6665
rect 11675 6515 11690 6665
rect 11810 6515 11825 6665
rect 11865 6515 11880 6665
rect 11920 6515 11935 6665
rect 11975 6515 11990 6665
rect 12110 6515 12125 6665
rect 12165 6515 12180 6665
rect 12220 6515 12235 6665
rect 12275 6515 12290 6665
rect 12330 6515 12345 6665
rect 12385 6515 12400 6665
rect 12440 6515 12455 6665
rect 12495 6515 12510 6665
rect 12550 6515 12565 6665
rect 12605 6515 12620 6665
rect 12660 6515 12675 6665
rect 12715 6515 12730 6665
rect 18570 6515 18585 6665
rect 18625 6515 18640 6665
rect 18680 6515 18695 6665
rect 18735 6515 18750 6665
rect 18790 6515 18805 6665
rect 18845 6515 18860 6665
rect 18900 6515 18915 6665
rect 18955 6515 18970 6665
rect 19010 6515 19025 6665
rect 19065 6515 19080 6665
rect 19120 6515 19135 6665
rect 19175 6515 19190 6665
rect 19310 6515 19325 6665
rect 19365 6515 19380 6665
rect 19420 6515 19435 6665
rect 19475 6515 19490 6665
rect 19610 6515 19625 6665
rect 19665 6515 19680 6665
rect 19720 6515 19735 6665
rect 19775 6515 19790 6665
rect 19830 6515 19845 6665
rect 19885 6515 19900 6665
rect 19940 6515 19955 6665
rect 19995 6515 20010 6665
rect 20050 6515 20065 6665
rect 20105 6515 20120 6665
rect 20160 6515 20175 6665
rect 20215 6515 20230 6665
rect 20435 6370 20450 6520
rect 20490 6370 20505 6520
rect 20545 6370 20560 6520
rect 20600 6370 20615 6520
rect 20735 6370 20750 6520
rect 20790 6370 20805 6520
rect 20845 6370 20860 6520
rect 20900 6370 20915 6520
rect 9705 6005 9765 6285
rect 9805 6005 9865 6285
rect 9905 6005 9965 6285
rect 10005 6005 10065 6285
rect 10105 6005 10165 6285
rect 10205 6005 10265 6285
rect 10305 6005 10365 6285
rect 10405 6005 10465 6285
rect 10505 6005 10565 6285
rect 10605 6005 10665 6285
rect 10705 6005 10765 6285
rect 10805 6005 10865 6285
rect 11245 5935 11260 6185
rect 11300 5935 11315 6185
rect 11355 5935 11370 6185
rect 11410 5935 11425 6185
rect 11465 5935 11480 6185
rect 11520 5935 11535 6185
rect 11575 5935 11590 6185
rect 11630 5935 11645 6185
rect 11685 5935 11700 6185
rect 11740 5935 11755 6185
rect 11795 5935 11810 6185
rect 11850 5935 11865 6185
rect 11905 5935 11920 6185
rect 11960 5935 11975 6185
rect 12015 5935 12030 6185
rect 12070 5935 12085 6185
rect 12125 5935 12140 6185
rect 12180 5935 12195 6185
rect 12235 5935 12250 6185
rect 12290 5935 12305 6185
rect 12345 5935 12360 6185
rect 12400 5935 12415 6185
rect 12455 5935 12470 6185
rect 12510 5935 12525 6185
rect 12565 5935 12580 6185
rect 12935 6005 12995 6285
rect 13035 6005 13095 6285
rect 13135 6005 13195 6285
rect 13235 6005 13295 6285
rect 13335 6005 13395 6285
rect 13435 6005 13495 6285
rect 13535 6005 13595 6285
rect 13635 6005 13695 6285
rect 13735 6005 13795 6285
rect 13835 6005 13895 6285
rect 13935 6005 13995 6285
rect 14035 6005 14095 6285
rect 18745 5975 18760 6225
rect 18800 5975 18815 6225
rect 18855 5975 18870 6225
rect 18910 5975 18925 6225
rect 18965 5975 18980 6225
rect 19020 5975 19035 6225
rect 19075 5975 19090 6225
rect 19130 5975 19145 6225
rect 19185 5975 19200 6225
rect 19240 5975 19255 6225
rect 19295 5975 19310 6225
rect 19350 5975 19365 6225
rect 19405 5975 19420 6225
rect 19460 5975 19475 6225
rect 19515 5975 19530 6225
rect 19570 5975 19585 6225
rect 19625 5975 19640 6225
rect 19680 5975 19695 6225
rect 19735 5975 19750 6225
rect 19790 5975 19805 6225
rect 19845 5975 19860 6225
rect 19900 5975 19915 6225
rect 19955 5975 19970 6225
rect 20010 5975 20025 6225
rect 20065 5975 20080 6225
rect 20585 6030 20600 6180
rect 20640 6030 20655 6180
rect 20695 6030 20710 6180
rect 20750 6030 20765 6180
rect 11280 4340 11300 4403
rect 11340 4340 11360 4403
rect 11400 4340 11420 4403
rect 11610 4340 11630 4420
rect 11670 4340 11690 4420
rect 11730 4340 11750 4420
rect 11790 4340 11810 4420
rect 11850 4340 11870 4420
rect 11910 4340 11930 4420
rect 12120 4335 12140 4395
rect 12180 4335 12200 4395
rect 12240 4335 12260 4395
rect 12300 4335 12320 4395
rect 12360 4335 12380 4395
rect 12420 4335 12440 4395
rect 12480 4335 12500 4395
rect 12540 4335 12560 4395
rect 11290 4105 11305 4155
rect 11345 4105 11360 4155
rect 11400 4105 11415 4155
rect 11455 4105 11470 4155
rect 11510 4105 11525 4155
rect 11565 4105 11580 4155
rect 11620 4105 11635 4155
rect 11675 4105 11690 4155
rect 11730 4105 11745 4155
rect 11785 4105 11800 4155
rect 11840 4105 11855 4155
rect 11895 4105 11910 4155
rect 11950 4105 11965 4155
rect 12005 4105 12020 4155
rect 12060 4105 12075 4155
rect 12115 4105 12130 4155
rect 12170 4105 12185 4155
rect 12225 4105 12240 4155
rect 12280 4105 12295 4155
rect 12335 4105 12350 4155
rect 12390 4105 12405 4155
rect 12445 4105 12460 4155
rect 11235 3800 11250 3850
rect 11290 3800 11305 3850
rect 11345 3800 11360 3850
rect 11400 3800 11415 3850
rect 11455 3800 11470 3850
rect 11510 3800 11525 3850
rect 11565 3800 11580 3850
rect 11620 3800 11635 3850
rect 11675 3800 11690 3850
rect 11730 3800 11745 3850
rect 11785 3800 11800 3850
rect 11840 3800 11855 3850
rect 11975 3800 11990 3850
rect 12030 3800 12045 3850
rect 12085 3800 12100 3850
rect 12140 3800 12155 3850
rect 12195 3800 12210 3850
rect 12250 3800 12265 3850
rect 12305 3800 12320 3850
rect 12360 3800 12375 3850
rect 12415 3800 12430 3850
rect 12470 3800 12485 3850
rect 12525 3800 12540 3850
rect 12580 3800 12595 3850
rect 10195 2985 10210 3585
rect 10250 2985 10265 3585
rect 10305 2985 10320 3585
rect 10360 2985 10375 3585
rect 10415 2985 10430 3585
rect 10470 2985 10485 3585
rect 10525 2985 10540 3585
rect 10580 2985 10595 3585
rect 10635 2985 10650 3585
rect 10690 2985 10705 3585
rect 10745 2985 10760 3585
rect 10800 2985 10815 3585
rect 11260 3175 11280 3575
rect 11320 3175 11340 3575
rect 11380 3175 11400 3575
rect 11440 3175 11460 3575
rect 11500 3175 11520 3575
rect 11560 3175 11580 3575
rect 11620 3175 11640 3575
rect 11680 3175 11700 3575
rect 11740 3175 11760 3575
rect 11800 3175 11820 3575
rect 11860 3175 11880 3575
rect 11920 3175 11940 3575
rect 11980 3175 12000 3575
rect 12040 3175 12060 3575
rect 12100 3175 12120 3575
rect 12160 3175 12180 3575
rect 12220 3175 12240 3575
rect 12280 3175 12300 3575
rect 12340 3175 12360 3575
rect 12400 3175 12420 3575
rect 12460 3175 12480 3575
rect 12520 3175 12540 3575
rect 12985 2985 13000 3585
rect 13040 2985 13055 3585
rect 13095 2985 13110 3585
rect 13150 2985 13165 3585
rect 13205 2985 13220 3585
rect 13260 2985 13275 3585
rect 13315 2985 13330 3585
rect 13370 2985 13385 3585
rect 13425 2985 13440 3585
rect 13480 2985 13495 3585
rect 13535 2985 13550 3585
rect 13590 2985 13605 3585
rect 25530 3230 25550 3293
rect 25590 3230 25610 3293
rect 25650 3230 25670 3293
rect 25860 3230 25880 3550
rect 25920 3230 25940 3550
rect 25980 3230 26000 3580
rect 26040 3230 26060 3580
rect 26260 3175 26280 3575
rect 26320 3175 26340 3575
rect 26380 3175 26400 3575
rect 26440 3175 26460 3575
rect 26500 3175 26520 3575
rect 26560 3175 26580 3575
rect 26620 3175 26640 3575
rect 26680 3175 26700 3575
rect 26740 3175 26760 3575
rect 26800 3175 26820 3575
rect 26860 3175 26880 3575
rect 26920 3175 26940 3575
rect 26980 3175 27000 3575
rect 27040 3175 27060 3575
rect 27100 3175 27120 3575
rect 27160 3175 27180 3575
rect 27220 3175 27240 3575
rect 27280 3175 27300 3575
rect 27340 3175 27360 3575
rect 27400 3175 27420 3575
rect 27460 3175 27480 3575
rect 27520 3175 27540 3575
rect 27930 2940 27945 3240
rect 27985 2940 28000 3240
rect 28040 2940 28055 3240
rect 28095 2940 28110 3240
rect 28150 2940 28165 3240
rect 28205 2940 28220 3240
rect 28260 2940 28275 3240
rect 28315 2940 28330 3240
rect 28370 2940 28385 3240
rect 28425 2940 28440 3240
rect 28480 2940 28495 3240
rect 28535 2940 28550 3240
rect 28590 2940 28605 3240
rect 28645 2940 28660 3240
rect 28700 2940 28715 3240
rect 28755 2940 28770 3240
rect 28810 2940 28825 3240
rect 28865 2940 28880 3240
rect 28920 2940 28935 3240
rect 28975 2940 28990 3240
rect 29030 2940 29045 3240
rect 29085 2940 29100 3240
rect 10195 2455 10210 2655
rect 10250 2455 10265 2655
rect 10305 2455 10320 2655
rect 10360 2455 10375 2655
rect 10415 2455 10430 2655
rect 10470 2455 10485 2655
rect 10525 2455 10540 2655
rect 10580 2455 10595 2655
rect 10635 2455 10650 2655
rect 10690 2455 10705 2655
rect 10745 2455 10760 2655
rect 10800 2455 10815 2655
rect 11260 2495 11280 2895
rect 11320 2495 11340 2895
rect 11380 2495 11400 2895
rect 11440 2495 11460 2895
rect 11500 2495 11520 2895
rect 11560 2495 11580 2895
rect 11620 2495 11640 2895
rect 11680 2495 11700 2895
rect 11740 2495 11760 2895
rect 11800 2495 11820 2895
rect 11860 2495 11880 2895
rect 11920 2495 11940 2895
rect 11980 2495 12000 2895
rect 12040 2495 12060 2895
rect 12100 2495 12120 2895
rect 12160 2495 12180 2895
rect 12220 2495 12240 2895
rect 12280 2495 12300 2895
rect 12340 2495 12360 2895
rect 12400 2495 12420 2895
rect 12460 2495 12480 2895
rect 12520 2495 12540 2895
rect 12985 2455 13000 2655
rect 13040 2455 13055 2655
rect 13095 2455 13110 2655
rect 13150 2455 13165 2655
rect 13205 2455 13220 2655
rect 13260 2455 13275 2655
rect 13315 2455 13330 2655
rect 13370 2455 13385 2655
rect 13425 2455 13440 2655
rect 13480 2455 13495 2655
rect 13535 2455 13550 2655
rect 13590 2455 13605 2655
rect 10195 1965 10210 2265
rect 10250 1965 10265 2265
rect 10305 1965 10320 2265
rect 10360 1965 10375 2265
rect 10415 1965 10430 2265
rect 10470 1965 10485 2265
rect 10525 1965 10540 2265
rect 10580 1965 10595 2265
rect 10635 1965 10650 2265
rect 10690 1965 10705 2265
rect 10745 1965 10760 2265
rect 10800 1965 10815 2265
rect 11315 1980 11330 2130
rect 11370 1980 11385 2130
rect 11425 1980 11440 2130
rect 11480 1980 11495 2130
rect 11535 1980 11550 2130
rect 11590 1980 11605 2130
rect 11645 1980 11660 2130
rect 11700 1980 11715 2130
rect 11755 1980 11770 2130
rect 11810 1980 11825 2130
rect 11865 1980 11880 2130
rect 11920 1980 11935 2130
rect 11975 1980 11990 2130
rect 12030 1980 12045 2130
rect 12085 1980 12100 2130
rect 12140 1980 12155 2130
rect 12195 1980 12210 2130
rect 12250 1980 12265 2130
rect 12305 1980 12320 2130
rect 12360 1980 12375 2130
rect 12415 1980 12430 2130
rect 12470 1980 12485 2130
rect 12985 1965 13000 2265
rect 13040 1965 13055 2265
rect 13095 1965 13110 2265
rect 13150 1965 13165 2265
rect 13205 1965 13220 2265
rect 13260 1965 13275 2265
rect 13315 1965 13330 2265
rect 13370 1965 13385 2265
rect 13425 1965 13440 2265
rect 13480 1965 13495 2265
rect 13535 1965 13550 2265
rect 13590 1965 13605 2265
rect 24720 2520 24735 2620
rect 24775 2520 24790 2620
rect 24830 2520 24845 2620
rect 24885 2520 24900 2620
rect 24940 2520 24955 2620
rect 24995 2520 25010 2620
rect 25050 2520 25065 2620
rect 25105 2520 25120 2620
rect 25160 2520 25175 2620
rect 25215 2520 25230 2620
rect 25270 2520 25285 2620
rect 25325 2520 25340 2620
rect 25380 2520 25395 2620
rect 25435 2520 25450 2620
rect 25490 2520 25505 2620
rect 25545 2520 25560 2620
rect 25600 2520 25615 2620
rect 25655 2520 25670 2620
rect 25710 2520 25725 2620
rect 25765 2520 25780 2620
rect 25820 2520 25835 2620
rect 25875 2520 25890 2620
rect 26260 2495 26280 2895
rect 26320 2495 26340 2895
rect 26380 2495 26400 2895
rect 26440 2495 26460 2895
rect 26500 2495 26520 2895
rect 26560 2495 26580 2895
rect 26620 2495 26640 2895
rect 26680 2495 26700 2895
rect 26740 2495 26760 2895
rect 26800 2495 26820 2895
rect 26860 2495 26880 2895
rect 26920 2495 26940 2895
rect 26980 2495 27000 2895
rect 27040 2495 27060 2895
rect 27100 2495 27120 2895
rect 27160 2495 27180 2895
rect 27220 2495 27240 2895
rect 27280 2495 27300 2895
rect 27340 2495 27360 2895
rect 27400 2495 27420 2895
rect 27460 2495 27480 2895
rect 27520 2495 27540 2895
rect 27930 2520 27945 2620
rect 27985 2520 28000 2620
rect 28040 2520 28055 2620
rect 28095 2520 28110 2620
rect 28150 2520 28165 2620
rect 28205 2520 28220 2620
rect 28260 2520 28275 2620
rect 28315 2520 28330 2620
rect 28370 2520 28385 2620
rect 28425 2520 28440 2620
rect 28480 2520 28495 2620
rect 28535 2520 28550 2620
rect 28590 2520 28605 2620
rect 28645 2520 28660 2620
rect 28700 2520 28715 2620
rect 28755 2520 28770 2620
rect 28810 2520 28825 2620
rect 28865 2520 28880 2620
rect 28920 2520 28935 2620
rect 28975 2520 28990 2620
rect 29030 2520 29045 2620
rect 29085 2520 29100 2620
rect 24720 2020 24735 2170
rect 24775 2020 24790 2170
rect 24830 2020 24845 2170
rect 24885 2020 24900 2170
rect 24940 2020 24955 2170
rect 24995 2020 25010 2170
rect 25050 2020 25065 2170
rect 25105 2020 25120 2170
rect 25160 2020 25175 2170
rect 25215 2020 25230 2170
rect 25270 2020 25285 2170
rect 25325 2020 25340 2170
rect 25380 2020 25395 2170
rect 25435 2020 25450 2170
rect 25490 2020 25505 2170
rect 25545 2020 25560 2170
rect 25600 2020 25615 2170
rect 25655 2020 25670 2170
rect 25710 2020 25725 2170
rect 25765 2020 25780 2170
rect 25820 2020 25835 2170
rect 25875 2020 25890 2170
rect 26315 1980 26330 2130
rect 26370 1980 26385 2130
rect 26425 1980 26440 2130
rect 26480 1980 26495 2130
rect 26535 1980 26550 2130
rect 26590 1980 26605 2130
rect 26645 1980 26660 2130
rect 26700 1980 26715 2130
rect 26755 1980 26770 2130
rect 26810 1980 26825 2130
rect 26865 1980 26880 2130
rect 26920 1980 26935 2130
rect 26975 1980 26990 2130
rect 27030 1980 27045 2130
rect 27085 1980 27100 2130
rect 27140 1980 27155 2130
rect 27195 1980 27210 2130
rect 27250 1980 27265 2130
rect 27305 1980 27320 2130
rect 27360 1980 27375 2130
rect 27415 1980 27430 2130
rect 27470 1980 27485 2130
rect 27930 2020 27945 2170
rect 27985 2020 28000 2170
rect 28040 2020 28055 2170
rect 28095 2020 28110 2170
rect 28150 2020 28165 2170
rect 28205 2020 28220 2170
rect 28260 2020 28275 2170
rect 28315 2020 28330 2170
rect 28370 2020 28385 2170
rect 28425 2020 28440 2170
rect 28480 2020 28495 2170
rect 28535 2020 28550 2170
rect 28590 2020 28605 2170
rect 28645 2020 28660 2170
rect 28700 2020 28715 2170
rect 28755 2020 28770 2170
rect 28810 2020 28825 2170
rect 28865 2020 28880 2170
rect 28920 2020 28935 2170
rect 28975 2020 28990 2170
rect 29030 2020 29045 2170
rect 29085 2020 29100 2170
rect 28030 1705 28045 1855
rect 28085 1705 28100 1855
rect 28140 1705 28155 1855
rect 28195 1705 28210 1855
rect 28250 1705 28265 1855
rect 28305 1705 28320 1855
rect 3205 1615 3225 1665
rect 3265 1615 3285 1665
rect 3325 1615 3345 1665
rect 3385 1615 3405 1665
rect 3445 1615 3465 1665
rect 3505 1615 3525 1665
rect 3565 1615 3585 1665
rect 3625 1615 3645 1665
rect 3685 1615 3705 1665
rect 3745 1615 3765 1665
rect 4245 1615 4265 1665
rect 4305 1615 4325 1665
rect 4365 1615 4385 1665
rect 4425 1615 4445 1665
rect 4485 1615 4505 1665
rect 4545 1615 4565 1665
rect 4605 1615 4625 1665
rect 4665 1615 4685 1665
rect 4725 1615 4745 1665
rect 4785 1615 4805 1665
rect 2875 1205 3375 1455
rect 3415 1205 3915 1455
rect 4095 1205 4595 1455
rect 4635 1205 5135 1455
rect 2985 975 3985 1075
rect 4025 975 5025 1075
rect 10195 955 10255 1655
rect 10295 955 10355 1655
rect 10395 955 10455 1655
rect 10495 955 10555 1655
rect 10595 955 10655 1655
rect 10695 955 10755 1655
rect 11070 1515 11085 1665
rect 11125 1515 11140 1665
rect 11180 1515 11195 1665
rect 11235 1515 11250 1665
rect 11290 1515 11305 1665
rect 11345 1515 11360 1665
rect 11400 1515 11415 1665
rect 11455 1515 11470 1665
rect 11510 1515 11525 1665
rect 11565 1515 11580 1665
rect 11620 1515 11635 1665
rect 11675 1515 11690 1665
rect 11810 1515 11825 1665
rect 11865 1515 11880 1665
rect 11920 1515 11935 1665
rect 11975 1515 11990 1665
rect 12110 1515 12125 1665
rect 12165 1515 12180 1665
rect 12220 1515 12235 1665
rect 12275 1515 12290 1665
rect 12330 1515 12345 1665
rect 12385 1515 12400 1665
rect 12440 1515 12455 1665
rect 12495 1515 12510 1665
rect 12550 1515 12565 1665
rect 12605 1515 12620 1665
rect 12660 1515 12675 1665
rect 12715 1515 12730 1665
rect 11245 935 11260 1185
rect 11300 935 11315 1185
rect 11355 935 11370 1185
rect 11410 935 11425 1185
rect 11465 935 11480 1185
rect 11520 935 11535 1185
rect 11575 935 11590 1185
rect 11630 935 11645 1185
rect 11685 935 11700 1185
rect 11740 935 11755 1185
rect 11795 935 11810 1185
rect 11850 935 11865 1185
rect 11905 935 11920 1185
rect 11960 935 11975 1185
rect 12015 935 12030 1185
rect 12070 935 12085 1185
rect 12125 935 12140 1185
rect 12180 935 12195 1185
rect 12235 935 12250 1185
rect 12290 935 12305 1185
rect 12345 935 12360 1185
rect 12400 935 12415 1185
rect 12455 935 12470 1185
rect 12510 935 12525 1185
rect 12565 935 12580 1185
rect 13045 955 13105 1655
rect 13145 955 13205 1655
rect 13245 955 13305 1655
rect 13345 955 13405 1655
rect 13445 955 13505 1655
rect 13545 955 13605 1655
rect 26070 1515 26085 1665
rect 26125 1515 26140 1665
rect 26180 1515 26195 1665
rect 26235 1515 26250 1665
rect 26290 1515 26305 1665
rect 26345 1515 26360 1665
rect 26400 1515 26415 1665
rect 26455 1515 26470 1665
rect 26510 1515 26525 1665
rect 26565 1515 26580 1665
rect 26620 1515 26635 1665
rect 26675 1515 26690 1665
rect 26810 1515 26825 1665
rect 26865 1515 26880 1665
rect 26920 1515 26935 1665
rect 26975 1515 26990 1665
rect 27110 1515 27125 1665
rect 27165 1515 27180 1665
rect 27220 1515 27235 1665
rect 27275 1515 27290 1665
rect 27330 1515 27345 1665
rect 27385 1515 27400 1665
rect 27440 1515 27455 1665
rect 27495 1515 27510 1665
rect 27550 1515 27565 1665
rect 27605 1515 27620 1665
rect 27660 1515 27675 1665
rect 27715 1515 27730 1665
rect 27935 1370 27950 1520
rect 27990 1370 28005 1520
rect 28045 1370 28060 1520
rect 28100 1370 28115 1520
rect 28235 1370 28250 1520
rect 28290 1370 28305 1520
rect 28345 1370 28360 1520
rect 28400 1370 28415 1520
rect 26245 975 26260 1225
rect 26300 975 26315 1225
rect 26355 975 26370 1225
rect 26410 975 26425 1225
rect 26465 975 26480 1225
rect 26520 975 26535 1225
rect 26575 975 26590 1225
rect 26630 975 26645 1225
rect 26685 975 26700 1225
rect 26740 975 26755 1225
rect 26795 975 26810 1225
rect 26850 975 26865 1225
rect 26905 975 26920 1225
rect 26960 975 26975 1225
rect 27015 975 27030 1225
rect 27070 975 27085 1225
rect 27125 975 27140 1225
rect 27180 975 27195 1225
rect 27235 975 27250 1225
rect 27290 975 27305 1225
rect 27345 975 27360 1225
rect 27400 975 27415 1225
rect 27455 975 27470 1225
rect 27510 975 27525 1225
rect 27565 975 27580 1225
rect 28085 1030 28100 1180
rect 28140 1030 28155 1180
rect 28195 1030 28210 1180
rect 28250 1030 28265 1180
rect 3035 780 3085 880
rect 3125 780 3175 880
rect 3215 780 3265 880
rect 3305 780 3355 880
rect 3395 780 3445 880
rect 3485 780 3535 880
rect 3575 780 3625 880
rect 3665 780 3715 880
rect 3755 780 3805 880
rect 3845 780 3895 880
rect 3935 780 3985 880
rect 4025 780 4075 880
rect 4115 780 4165 880
rect 4205 780 4255 880
rect 4295 780 4345 880
rect 4385 780 4435 880
rect 4475 780 4525 880
rect 4565 780 4615 880
rect 4655 780 4705 880
rect 4745 780 4795 880
rect 4835 780 4885 880
rect 4925 780 4975 880
rect 11300 645 11490 745
rect 11920 700 11935 750
rect 11975 700 11990 750
rect 12030 700 12045 750
rect 12085 700 12100 750
rect 12140 700 12155 750
rect 12195 700 12210 750
rect 12250 700 12265 750
rect 12305 700 12320 750
rect 12360 700 12375 750
rect 12415 700 12430 750
rect 12470 700 12485 750
rect 12525 700 12540 750
rect 10530 -1770 10550 -1707
rect 10590 -1770 10610 -1707
rect 10650 -1770 10670 -1707
rect 10860 -1770 10880 -1450
rect 10920 -1770 10940 -1450
rect 10980 -1770 11000 -1420
rect 11040 -1770 11060 -1420
rect 11260 -1825 11280 -1425
rect 11320 -1825 11340 -1425
rect 11380 -1825 11400 -1425
rect 11440 -1825 11460 -1425
rect 11500 -1825 11520 -1425
rect 11560 -1825 11580 -1425
rect 11620 -1825 11640 -1425
rect 11680 -1825 11700 -1425
rect 11740 -1825 11760 -1425
rect 11800 -1825 11820 -1425
rect 11860 -1825 11880 -1425
rect 11920 -1825 11940 -1425
rect 11980 -1825 12000 -1425
rect 12040 -1825 12060 -1425
rect 12100 -1825 12120 -1425
rect 12160 -1825 12180 -1425
rect 12220 -1825 12240 -1425
rect 12280 -1825 12300 -1425
rect 12340 -1825 12360 -1425
rect 12400 -1825 12420 -1425
rect 12460 -1825 12480 -1425
rect 12520 -1825 12540 -1425
rect 11260 -2505 11280 -2105
rect 11320 -2505 11340 -2105
rect 11380 -2505 11400 -2105
rect 11440 -2505 11460 -2105
rect 11500 -2505 11520 -2105
rect 11560 -2505 11580 -2105
rect 11620 -2505 11640 -2105
rect 11680 -2505 11700 -2105
rect 11740 -2505 11760 -2105
rect 11800 -2505 11820 -2105
rect 11860 -2505 11880 -2105
rect 11920 -2505 11940 -2105
rect 11980 -2505 12000 -2105
rect 12040 -2505 12060 -2105
rect 12100 -2505 12120 -2105
rect 12160 -2505 12180 -2105
rect 12220 -2505 12240 -2105
rect 12280 -2505 12300 -2105
rect 12340 -2505 12360 -2105
rect 12400 -2505 12420 -2105
rect 12460 -2505 12480 -2105
rect 12520 -2505 12540 -2105
rect 12935 -2315 12950 -2015
rect 12990 -2315 13005 -2015
rect 13045 -2315 13060 -2015
rect 13100 -2315 13115 -2015
rect 13155 -2315 13170 -2015
rect 13210 -2315 13225 -2015
rect 13265 -2315 13280 -2015
rect 13320 -2315 13335 -2015
rect 13375 -2315 13390 -2015
rect 13430 -2315 13445 -2015
rect 13485 -2315 13500 -2015
rect 13540 -2315 13555 -2015
rect 13595 -2315 13610 -2015
rect 13650 -2315 13665 -2015
rect 13705 -2315 13720 -2015
rect 13760 -2315 13775 -2015
rect 13815 -2315 13830 -2015
rect 13870 -2315 13885 -2015
rect 13925 -2315 13940 -2015
rect 13980 -2315 13995 -2015
rect 14035 -2315 14050 -2015
rect 14090 -2315 14105 -2015
rect 12935 -2545 12950 -2445
rect 12990 -2545 13005 -2445
rect 13045 -2545 13060 -2445
rect 13100 -2545 13115 -2445
rect 13155 -2545 13170 -2445
rect 13210 -2545 13225 -2445
rect 13265 -2545 13280 -2445
rect 13320 -2545 13335 -2445
rect 13375 -2545 13390 -2445
rect 13430 -2545 13445 -2445
rect 13485 -2545 13500 -2445
rect 13540 -2545 13555 -2445
rect 13595 -2545 13610 -2445
rect 13650 -2545 13665 -2445
rect 13705 -2545 13720 -2445
rect 13760 -2545 13775 -2445
rect 13815 -2545 13830 -2445
rect 13870 -2545 13885 -2445
rect 13925 -2545 13940 -2445
rect 13980 -2545 13995 -2445
rect 14035 -2545 14050 -2445
rect 14090 -2545 14105 -2445
rect 11315 -3020 11330 -2870
rect 11370 -3020 11385 -2870
rect 11425 -3020 11440 -2870
rect 11480 -3020 11495 -2870
rect 11535 -3020 11550 -2870
rect 11590 -3020 11605 -2870
rect 11645 -3020 11660 -2870
rect 11700 -3020 11715 -2870
rect 11755 -3020 11770 -2870
rect 11810 -3020 11825 -2870
rect 11865 -3020 11880 -2870
rect 11920 -3020 11935 -2870
rect 11975 -3020 11990 -2870
rect 12030 -3020 12045 -2870
rect 12085 -3020 12100 -2870
rect 12140 -3020 12155 -2870
rect 12195 -3020 12210 -2870
rect 12250 -3020 12265 -2870
rect 12305 -3020 12320 -2870
rect 12360 -3020 12375 -2870
rect 12415 -3020 12430 -2870
rect 12470 -3020 12485 -2870
rect 12935 -2885 12950 -2735
rect 12990 -2885 13005 -2735
rect 13045 -2885 13060 -2735
rect 13100 -2885 13115 -2735
rect 13155 -2885 13170 -2735
rect 13210 -2885 13225 -2735
rect 13265 -2885 13280 -2735
rect 13320 -2885 13335 -2735
rect 13375 -2885 13390 -2735
rect 13430 -2885 13445 -2735
rect 13485 -2885 13500 -2735
rect 13540 -2885 13555 -2735
rect 13595 -2885 13610 -2735
rect 13650 -2885 13665 -2735
rect 13705 -2885 13720 -2735
rect 13760 -2885 13775 -2735
rect 13815 -2885 13830 -2735
rect 13870 -2885 13885 -2735
rect 13925 -2885 13940 -2735
rect 13980 -2885 13995 -2735
rect 14035 -2885 14050 -2735
rect 14090 -2885 14105 -2735
rect 12935 -3295 12995 -3015
rect 13035 -3295 13095 -3015
rect 13135 -3295 13195 -3015
rect 13235 -3295 13295 -3015
rect 13335 -3295 13395 -3015
rect 13435 -3295 13495 -3015
rect 13535 -3295 13595 -3015
rect 13635 -3295 13695 -3015
rect 13735 -3295 13795 -3015
rect 13835 -3295 13895 -3015
rect 13935 -3295 13995 -3015
rect 14035 -3295 14095 -3015
rect 11070 -3485 11085 -3335
rect 11125 -3485 11140 -3335
rect 11180 -3485 11195 -3335
rect 11235 -3485 11250 -3335
rect 11290 -3485 11305 -3335
rect 11345 -3485 11360 -3335
rect 11400 -3485 11415 -3335
rect 11455 -3485 11470 -3335
rect 11510 -3485 11525 -3335
rect 11565 -3485 11580 -3335
rect 11620 -3485 11635 -3335
rect 11675 -3485 11690 -3335
rect 11810 -3485 11825 -3335
rect 11865 -3485 11880 -3335
rect 11920 -3485 11935 -3335
rect 11975 -3485 11990 -3335
rect 12110 -3485 12125 -3335
rect 12165 -3485 12180 -3335
rect 12220 -3485 12235 -3335
rect 12275 -3485 12290 -3335
rect 12330 -3485 12345 -3335
rect 12385 -3485 12400 -3335
rect 12440 -3485 12455 -3335
rect 12495 -3485 12510 -3335
rect 12550 -3485 12565 -3335
rect 12605 -3485 12620 -3335
rect 12660 -3485 12675 -3335
rect 12715 -3485 12730 -3335
rect 11245 -4065 11260 -3815
rect 11300 -4065 11315 -3815
rect 11355 -4065 11370 -3815
rect 11410 -4065 11425 -3815
rect 11465 -4065 11480 -3815
rect 11520 -4065 11535 -3815
rect 11575 -4065 11590 -3815
rect 11630 -4065 11645 -3815
rect 11685 -4065 11700 -3815
rect 11740 -4065 11755 -3815
rect 11795 -4065 11810 -3815
rect 11850 -4065 11865 -3815
rect 11905 -4065 11920 -3815
rect 11960 -4065 11975 -3815
rect 12015 -4065 12030 -3815
rect 12070 -4065 12085 -3815
rect 12125 -4065 12140 -3815
rect 12180 -4065 12195 -3815
rect 12235 -4065 12250 -3815
rect 12290 -4065 12305 -3815
rect 12345 -4065 12360 -3815
rect 12400 -4065 12415 -3815
rect 12455 -4065 12470 -3815
rect 12510 -4065 12525 -3815
rect 12565 -4065 12580 -3815
<< pmos >>
rect 3035 2830 3085 2930
rect 3125 2830 3175 2930
rect 3215 2830 3265 2930
rect 3305 2830 3355 2930
rect 3395 2830 3445 2930
rect 3485 2830 3535 2930
rect 3575 2830 3625 2930
rect 3665 2830 3715 2930
rect 3755 2830 3805 2930
rect 3845 2830 3895 2930
rect 3935 2830 3985 2930
rect 4025 2830 4075 2930
rect 4115 2830 4165 2930
rect 4205 2830 4255 2930
rect 4295 2830 4345 2930
rect 4385 2830 4435 2930
rect 4475 2830 4525 2930
rect 4565 2830 4615 2930
rect 4655 2830 4705 2930
rect 4745 2830 4795 2930
rect 4835 2830 4885 2930
rect 4925 2830 4975 2930
rect 3215 2400 3265 2700
rect 3305 2400 3355 2700
rect 3395 2400 3445 2700
rect 3485 2400 3535 2700
rect 3575 2400 3625 2700
rect 3665 2400 3715 2700
rect 3755 2400 3805 2700
rect 3845 2400 3895 2700
rect 3935 2400 3985 2700
rect 4025 2400 4075 2700
rect 4115 2400 4165 2700
rect 4205 2400 4255 2700
rect 4295 2400 4345 2700
rect 4385 2400 4435 2700
rect 4475 2400 4525 2700
rect 4565 2400 4615 2700
rect 4655 2400 4705 2700
rect 4745 2400 4795 2700
rect 2605 1900 2620 2000
rect 2660 1900 2675 2000
rect 2785 1900 2805 2000
rect 2845 1900 2865 2000
rect 2905 1900 2925 2000
rect 2965 1900 2985 2000
rect 3025 1900 3045 2000
rect 3085 1900 3105 2000
rect 3145 1900 3165 2000
rect 3205 1900 3225 2000
rect 3265 1900 3285 2000
rect 3325 1900 3345 2000
rect 3385 1900 3405 2000
rect 3445 1900 3465 2000
rect 3505 1900 3525 2000
rect 3565 1900 3585 2000
rect 3625 1900 3645 2000
rect 3685 1900 3705 2000
rect 3745 1900 3765 2000
rect 3805 1900 3825 2000
rect 3865 1900 3885 2000
rect 3925 1900 3945 2000
rect 4065 1900 4085 2000
rect 4125 1900 4145 2000
rect 4185 1900 4205 2000
rect 4245 1900 4265 2000
rect 4305 1900 4325 2000
rect 4365 1900 4385 2000
rect 4425 1900 4445 2000
rect 4485 1900 4505 2000
rect 4545 1900 4565 2000
rect 4605 1900 4625 2000
rect 4665 1900 4685 2000
rect 4725 1900 4745 2000
rect 4785 1900 4805 2000
rect 4845 1900 4865 2000
rect 4905 1900 4925 2000
rect 4965 1900 4985 2000
rect 5025 1900 5045 2000
rect 5085 1900 5105 2000
rect 5145 1900 5165 2000
rect 5205 1900 5225 2000
<< ndiff >>
rect 11240 8915 11280 8943
rect 11240 8895 11250 8915
rect 11270 8895 11280 8915
rect 11240 8880 11280 8895
rect 11300 8920 11340 8943
rect 11300 8900 11310 8920
rect 11330 8900 11340 8920
rect 11300 8880 11340 8900
rect 11360 8920 11400 8943
rect 11360 8900 11370 8920
rect 11390 8900 11400 8920
rect 11360 8880 11400 8900
rect 11420 8915 11460 8943
rect 11420 8895 11430 8915
rect 11450 8895 11460 8915
rect 11420 8880 11460 8895
rect 11570 8930 11610 8960
rect 11570 8910 11580 8930
rect 11600 8910 11610 8930
rect 11570 8880 11610 8910
rect 11630 8930 11670 8960
rect 11630 8910 11640 8930
rect 11660 8910 11670 8930
rect 11630 8880 11670 8910
rect 11690 8930 11730 8960
rect 11690 8910 11700 8930
rect 11720 8910 11730 8930
rect 11690 8880 11730 8910
rect 11750 8930 11790 8960
rect 11750 8910 11760 8930
rect 11780 8910 11790 8930
rect 11750 8880 11790 8910
rect 11810 8930 11850 8960
rect 11810 8910 11820 8930
rect 11840 8910 11850 8930
rect 11810 8880 11850 8910
rect 11870 8930 11910 8960
rect 11870 8910 11880 8930
rect 11900 8910 11910 8930
rect 11870 8880 11910 8910
rect 11930 8930 11970 8960
rect 11930 8910 11940 8930
rect 11960 8910 11970 8930
rect 11930 8880 11970 8910
rect 12080 8915 12120 8935
rect 12080 8895 12090 8915
rect 12110 8895 12120 8915
rect 12080 8875 12120 8895
rect 12140 8915 12180 8935
rect 12140 8895 12150 8915
rect 12170 8895 12180 8915
rect 12140 8875 12180 8895
rect 12200 8915 12240 8935
rect 12200 8895 12210 8915
rect 12230 8895 12240 8915
rect 12200 8875 12240 8895
rect 12260 8915 12300 8935
rect 12260 8895 12270 8915
rect 12290 8895 12300 8915
rect 12260 8875 12300 8895
rect 12320 8915 12360 8935
rect 12320 8895 12330 8915
rect 12350 8895 12360 8915
rect 12320 8875 12360 8895
rect 12380 8915 12420 8935
rect 12380 8895 12390 8915
rect 12410 8895 12420 8915
rect 12380 8875 12420 8895
rect 12440 8915 12480 8935
rect 12440 8895 12450 8915
rect 12470 8895 12480 8915
rect 12440 8875 12480 8895
rect 12500 8915 12540 8935
rect 12500 8895 12510 8915
rect 12530 8895 12540 8915
rect 12500 8875 12540 8895
rect 12560 8915 12600 8935
rect 12560 8895 12570 8915
rect 12590 8895 12600 8915
rect 12560 8875 12600 8895
rect 10955 8550 10980 8580
rect 10820 8515 10860 8550
rect 10820 8495 10830 8515
rect 10850 8495 10860 8515
rect 10820 8465 10860 8495
rect 10820 8445 10830 8465
rect 10850 8445 10860 8465
rect 10820 8415 10860 8445
rect 10820 8395 10830 8415
rect 10850 8395 10860 8415
rect 10820 8365 10860 8395
rect 10820 8345 10830 8365
rect 10850 8345 10860 8365
rect 10820 8315 10860 8345
rect 10820 8295 10830 8315
rect 10850 8295 10860 8315
rect 10490 8265 10530 8293
rect 10490 8245 10500 8265
rect 10520 8245 10530 8265
rect 10490 8230 10530 8245
rect 10550 8270 10590 8293
rect 10550 8250 10560 8270
rect 10580 8250 10590 8270
rect 10550 8230 10590 8250
rect 10610 8270 10650 8293
rect 10610 8250 10620 8270
rect 10640 8250 10650 8270
rect 10610 8230 10650 8250
rect 10670 8265 10710 8293
rect 10670 8245 10680 8265
rect 10700 8245 10710 8265
rect 10670 8230 10710 8245
rect 10820 8265 10860 8295
rect 10820 8245 10830 8265
rect 10850 8245 10860 8265
rect 10820 8230 10860 8245
rect 10880 8515 10920 8550
rect 10880 8495 10890 8515
rect 10910 8495 10920 8515
rect 10880 8465 10920 8495
rect 10880 8445 10890 8465
rect 10910 8445 10920 8465
rect 10880 8415 10920 8445
rect 10880 8395 10890 8415
rect 10910 8395 10920 8415
rect 10880 8365 10920 8395
rect 10880 8345 10890 8365
rect 10910 8345 10920 8365
rect 10880 8315 10920 8345
rect 10880 8295 10890 8315
rect 10910 8295 10920 8315
rect 10880 8265 10920 8295
rect 10880 8245 10890 8265
rect 10910 8245 10920 8265
rect 10880 8230 10920 8245
rect 10940 8515 10980 8550
rect 10940 8495 10950 8515
rect 10970 8495 10980 8515
rect 10940 8465 10980 8495
rect 10940 8445 10950 8465
rect 10970 8445 10980 8465
rect 10940 8415 10980 8445
rect 10940 8395 10950 8415
rect 10970 8395 10980 8415
rect 10940 8365 10980 8395
rect 10940 8345 10950 8365
rect 10970 8345 10980 8365
rect 10940 8315 10980 8345
rect 10940 8295 10950 8315
rect 10970 8295 10980 8315
rect 10940 8265 10980 8295
rect 10940 8245 10950 8265
rect 10970 8245 10980 8265
rect 10940 8230 10980 8245
rect 11000 8565 11040 8580
rect 11000 8545 11010 8565
rect 11030 8545 11040 8565
rect 11000 8515 11040 8545
rect 11000 8495 11010 8515
rect 11030 8495 11040 8515
rect 11000 8465 11040 8495
rect 11000 8445 11010 8465
rect 11030 8445 11040 8465
rect 11000 8415 11040 8445
rect 11000 8395 11010 8415
rect 11030 8395 11040 8415
rect 11000 8365 11040 8395
rect 11000 8345 11010 8365
rect 11030 8345 11040 8365
rect 11000 8315 11040 8345
rect 11000 8295 11010 8315
rect 11030 8295 11040 8315
rect 11000 8265 11040 8295
rect 11000 8245 11010 8265
rect 11030 8245 11040 8265
rect 11000 8230 11040 8245
rect 11060 8565 11100 8580
rect 11060 8545 11070 8565
rect 11090 8545 11100 8565
rect 11060 8515 11100 8545
rect 11060 8495 11070 8515
rect 11090 8495 11100 8515
rect 11060 8465 11100 8495
rect 11060 8445 11070 8465
rect 11090 8445 11100 8465
rect 11060 8415 11100 8445
rect 11060 8395 11070 8415
rect 11090 8395 11100 8415
rect 11060 8365 11100 8395
rect 11060 8345 11070 8365
rect 11090 8345 11100 8365
rect 11060 8315 11100 8345
rect 11060 8295 11070 8315
rect 11090 8295 11100 8315
rect 11060 8265 11100 8295
rect 11060 8245 11070 8265
rect 11090 8245 11100 8265
rect 11060 8230 11100 8245
rect 11220 8560 11260 8575
rect 11220 8540 11230 8560
rect 11250 8540 11260 8560
rect 11220 8510 11260 8540
rect 11220 8490 11230 8510
rect 11250 8490 11260 8510
rect 11220 8460 11260 8490
rect 11220 8440 11230 8460
rect 11250 8440 11260 8460
rect 11220 8410 11260 8440
rect 11220 8390 11230 8410
rect 11250 8390 11260 8410
rect 11220 8360 11260 8390
rect 11220 8340 11230 8360
rect 11250 8340 11260 8360
rect 11220 8310 11260 8340
rect 11220 8290 11230 8310
rect 11250 8290 11260 8310
rect 11220 8260 11260 8290
rect 11220 8240 11230 8260
rect 11250 8240 11260 8260
rect 11220 8210 11260 8240
rect 11220 8190 11230 8210
rect 11250 8190 11260 8210
rect 11220 8175 11260 8190
rect 11280 8560 11320 8575
rect 11280 8540 11290 8560
rect 11310 8540 11320 8560
rect 11280 8510 11320 8540
rect 11280 8490 11290 8510
rect 11310 8490 11320 8510
rect 11280 8460 11320 8490
rect 11280 8440 11290 8460
rect 11310 8440 11320 8460
rect 11280 8410 11320 8440
rect 11280 8390 11290 8410
rect 11310 8390 11320 8410
rect 11280 8360 11320 8390
rect 11280 8340 11290 8360
rect 11310 8340 11320 8360
rect 11280 8310 11320 8340
rect 11280 8290 11290 8310
rect 11310 8290 11320 8310
rect 11280 8260 11320 8290
rect 11280 8240 11290 8260
rect 11310 8240 11320 8260
rect 11280 8210 11320 8240
rect 11280 8190 11290 8210
rect 11310 8190 11320 8210
rect 11280 8175 11320 8190
rect 11340 8560 11380 8575
rect 11340 8540 11350 8560
rect 11370 8540 11380 8560
rect 11340 8510 11380 8540
rect 11340 8490 11350 8510
rect 11370 8490 11380 8510
rect 11340 8460 11380 8490
rect 11340 8440 11350 8460
rect 11370 8440 11380 8460
rect 11340 8410 11380 8440
rect 11340 8390 11350 8410
rect 11370 8390 11380 8410
rect 11340 8360 11380 8390
rect 11340 8340 11350 8360
rect 11370 8340 11380 8360
rect 11340 8310 11380 8340
rect 11340 8290 11350 8310
rect 11370 8290 11380 8310
rect 11340 8260 11380 8290
rect 11340 8240 11350 8260
rect 11370 8240 11380 8260
rect 11340 8210 11380 8240
rect 11340 8190 11350 8210
rect 11370 8190 11380 8210
rect 11340 8175 11380 8190
rect 11400 8560 11440 8575
rect 11400 8540 11410 8560
rect 11430 8540 11440 8560
rect 11400 8510 11440 8540
rect 11400 8490 11410 8510
rect 11430 8490 11440 8510
rect 11400 8460 11440 8490
rect 11400 8440 11410 8460
rect 11430 8440 11440 8460
rect 11400 8410 11440 8440
rect 11400 8390 11410 8410
rect 11430 8390 11440 8410
rect 11400 8360 11440 8390
rect 11400 8340 11410 8360
rect 11430 8340 11440 8360
rect 11400 8310 11440 8340
rect 11400 8290 11410 8310
rect 11430 8290 11440 8310
rect 11400 8260 11440 8290
rect 11400 8240 11410 8260
rect 11430 8240 11440 8260
rect 11400 8210 11440 8240
rect 11400 8190 11410 8210
rect 11430 8190 11440 8210
rect 11400 8175 11440 8190
rect 11460 8560 11500 8575
rect 11460 8540 11470 8560
rect 11490 8540 11500 8560
rect 11460 8510 11500 8540
rect 11460 8490 11470 8510
rect 11490 8490 11500 8510
rect 11460 8460 11500 8490
rect 11460 8440 11470 8460
rect 11490 8440 11500 8460
rect 11460 8410 11500 8440
rect 11460 8390 11470 8410
rect 11490 8390 11500 8410
rect 11460 8360 11500 8390
rect 11460 8340 11470 8360
rect 11490 8340 11500 8360
rect 11460 8310 11500 8340
rect 11460 8290 11470 8310
rect 11490 8290 11500 8310
rect 11460 8260 11500 8290
rect 11460 8240 11470 8260
rect 11490 8240 11500 8260
rect 11460 8210 11500 8240
rect 11460 8190 11470 8210
rect 11490 8190 11500 8210
rect 11460 8175 11500 8190
rect 11520 8560 11560 8575
rect 11520 8540 11530 8560
rect 11550 8540 11560 8560
rect 11520 8510 11560 8540
rect 11520 8490 11530 8510
rect 11550 8490 11560 8510
rect 11520 8460 11560 8490
rect 11520 8440 11530 8460
rect 11550 8440 11560 8460
rect 11520 8410 11560 8440
rect 11520 8390 11530 8410
rect 11550 8390 11560 8410
rect 11520 8360 11560 8390
rect 11520 8340 11530 8360
rect 11550 8340 11560 8360
rect 11520 8310 11560 8340
rect 11520 8290 11530 8310
rect 11550 8290 11560 8310
rect 11520 8260 11560 8290
rect 11520 8240 11530 8260
rect 11550 8240 11560 8260
rect 11520 8210 11560 8240
rect 11520 8190 11530 8210
rect 11550 8190 11560 8210
rect 11520 8175 11560 8190
rect 11580 8560 11620 8575
rect 11580 8540 11590 8560
rect 11610 8540 11620 8560
rect 11580 8510 11620 8540
rect 11580 8490 11590 8510
rect 11610 8490 11620 8510
rect 11580 8460 11620 8490
rect 11580 8440 11590 8460
rect 11610 8440 11620 8460
rect 11580 8410 11620 8440
rect 11580 8390 11590 8410
rect 11610 8390 11620 8410
rect 11580 8360 11620 8390
rect 11580 8340 11590 8360
rect 11610 8340 11620 8360
rect 11580 8310 11620 8340
rect 11580 8290 11590 8310
rect 11610 8290 11620 8310
rect 11580 8260 11620 8290
rect 11580 8240 11590 8260
rect 11610 8240 11620 8260
rect 11580 8210 11620 8240
rect 11580 8190 11590 8210
rect 11610 8190 11620 8210
rect 11580 8175 11620 8190
rect 11640 8560 11680 8575
rect 11640 8540 11650 8560
rect 11670 8540 11680 8560
rect 11640 8510 11680 8540
rect 11640 8490 11650 8510
rect 11670 8490 11680 8510
rect 11640 8460 11680 8490
rect 11640 8440 11650 8460
rect 11670 8440 11680 8460
rect 11640 8410 11680 8440
rect 11640 8390 11650 8410
rect 11670 8390 11680 8410
rect 11640 8360 11680 8390
rect 11640 8340 11650 8360
rect 11670 8340 11680 8360
rect 11640 8310 11680 8340
rect 11640 8290 11650 8310
rect 11670 8290 11680 8310
rect 11640 8260 11680 8290
rect 11640 8240 11650 8260
rect 11670 8240 11680 8260
rect 11640 8210 11680 8240
rect 11640 8190 11650 8210
rect 11670 8190 11680 8210
rect 11640 8175 11680 8190
rect 11700 8560 11740 8575
rect 11700 8540 11710 8560
rect 11730 8540 11740 8560
rect 11700 8510 11740 8540
rect 11700 8490 11710 8510
rect 11730 8490 11740 8510
rect 11700 8460 11740 8490
rect 11700 8440 11710 8460
rect 11730 8440 11740 8460
rect 11700 8410 11740 8440
rect 11700 8390 11710 8410
rect 11730 8390 11740 8410
rect 11700 8360 11740 8390
rect 11700 8340 11710 8360
rect 11730 8340 11740 8360
rect 11700 8310 11740 8340
rect 11700 8290 11710 8310
rect 11730 8290 11740 8310
rect 11700 8260 11740 8290
rect 11700 8240 11710 8260
rect 11730 8240 11740 8260
rect 11700 8210 11740 8240
rect 11700 8190 11710 8210
rect 11730 8190 11740 8210
rect 11700 8175 11740 8190
rect 11760 8560 11800 8575
rect 11760 8540 11770 8560
rect 11790 8540 11800 8560
rect 11760 8510 11800 8540
rect 11760 8490 11770 8510
rect 11790 8490 11800 8510
rect 11760 8460 11800 8490
rect 11760 8440 11770 8460
rect 11790 8440 11800 8460
rect 11760 8410 11800 8440
rect 11760 8390 11770 8410
rect 11790 8390 11800 8410
rect 11760 8360 11800 8390
rect 11760 8340 11770 8360
rect 11790 8340 11800 8360
rect 11760 8310 11800 8340
rect 11760 8290 11770 8310
rect 11790 8290 11800 8310
rect 11760 8260 11800 8290
rect 11760 8240 11770 8260
rect 11790 8240 11800 8260
rect 11760 8210 11800 8240
rect 11760 8190 11770 8210
rect 11790 8190 11800 8210
rect 11760 8175 11800 8190
rect 11820 8560 11860 8575
rect 11820 8540 11830 8560
rect 11850 8540 11860 8560
rect 11820 8510 11860 8540
rect 11820 8490 11830 8510
rect 11850 8490 11860 8510
rect 11820 8460 11860 8490
rect 11820 8440 11830 8460
rect 11850 8440 11860 8460
rect 11820 8410 11860 8440
rect 11820 8390 11830 8410
rect 11850 8390 11860 8410
rect 11820 8360 11860 8390
rect 11820 8340 11830 8360
rect 11850 8340 11860 8360
rect 11820 8310 11860 8340
rect 11820 8290 11830 8310
rect 11850 8290 11860 8310
rect 11820 8260 11860 8290
rect 11820 8240 11830 8260
rect 11850 8240 11860 8260
rect 11820 8210 11860 8240
rect 11820 8190 11830 8210
rect 11850 8190 11860 8210
rect 11820 8175 11860 8190
rect 11880 8560 11920 8575
rect 11880 8540 11890 8560
rect 11910 8540 11920 8560
rect 11880 8510 11920 8540
rect 11880 8490 11890 8510
rect 11910 8490 11920 8510
rect 11880 8460 11920 8490
rect 11880 8440 11890 8460
rect 11910 8440 11920 8460
rect 11880 8410 11920 8440
rect 11880 8390 11890 8410
rect 11910 8390 11920 8410
rect 11880 8360 11920 8390
rect 11880 8340 11890 8360
rect 11910 8340 11920 8360
rect 11880 8310 11920 8340
rect 11880 8290 11890 8310
rect 11910 8290 11920 8310
rect 11880 8260 11920 8290
rect 11880 8240 11890 8260
rect 11910 8240 11920 8260
rect 11880 8210 11920 8240
rect 11880 8190 11890 8210
rect 11910 8190 11920 8210
rect 11880 8175 11920 8190
rect 11940 8560 11980 8575
rect 11940 8540 11950 8560
rect 11970 8540 11980 8560
rect 11940 8510 11980 8540
rect 11940 8490 11950 8510
rect 11970 8490 11980 8510
rect 11940 8460 11980 8490
rect 11940 8440 11950 8460
rect 11970 8440 11980 8460
rect 11940 8410 11980 8440
rect 11940 8390 11950 8410
rect 11970 8390 11980 8410
rect 11940 8360 11980 8390
rect 11940 8340 11950 8360
rect 11970 8340 11980 8360
rect 11940 8310 11980 8340
rect 11940 8290 11950 8310
rect 11970 8290 11980 8310
rect 11940 8260 11980 8290
rect 11940 8240 11950 8260
rect 11970 8240 11980 8260
rect 11940 8210 11980 8240
rect 11940 8190 11950 8210
rect 11970 8190 11980 8210
rect 11940 8175 11980 8190
rect 12000 8560 12040 8575
rect 12000 8540 12010 8560
rect 12030 8540 12040 8560
rect 12000 8510 12040 8540
rect 12000 8490 12010 8510
rect 12030 8490 12040 8510
rect 12000 8460 12040 8490
rect 12000 8440 12010 8460
rect 12030 8440 12040 8460
rect 12000 8410 12040 8440
rect 12000 8390 12010 8410
rect 12030 8390 12040 8410
rect 12000 8360 12040 8390
rect 12000 8340 12010 8360
rect 12030 8340 12040 8360
rect 12000 8310 12040 8340
rect 12000 8290 12010 8310
rect 12030 8290 12040 8310
rect 12000 8260 12040 8290
rect 12000 8240 12010 8260
rect 12030 8240 12040 8260
rect 12000 8210 12040 8240
rect 12000 8190 12010 8210
rect 12030 8190 12040 8210
rect 12000 8175 12040 8190
rect 12060 8560 12100 8575
rect 12060 8540 12070 8560
rect 12090 8540 12100 8560
rect 12060 8510 12100 8540
rect 12060 8490 12070 8510
rect 12090 8490 12100 8510
rect 12060 8460 12100 8490
rect 12060 8440 12070 8460
rect 12090 8440 12100 8460
rect 12060 8410 12100 8440
rect 12060 8390 12070 8410
rect 12090 8390 12100 8410
rect 12060 8360 12100 8390
rect 12060 8340 12070 8360
rect 12090 8340 12100 8360
rect 12060 8310 12100 8340
rect 12060 8290 12070 8310
rect 12090 8290 12100 8310
rect 12060 8260 12100 8290
rect 12060 8240 12070 8260
rect 12090 8240 12100 8260
rect 12060 8210 12100 8240
rect 12060 8190 12070 8210
rect 12090 8190 12100 8210
rect 12060 8175 12100 8190
rect 12120 8560 12160 8575
rect 12120 8540 12130 8560
rect 12150 8540 12160 8560
rect 12120 8510 12160 8540
rect 12120 8490 12130 8510
rect 12150 8490 12160 8510
rect 12120 8460 12160 8490
rect 12120 8440 12130 8460
rect 12150 8440 12160 8460
rect 12120 8410 12160 8440
rect 12120 8390 12130 8410
rect 12150 8390 12160 8410
rect 12120 8360 12160 8390
rect 12120 8340 12130 8360
rect 12150 8340 12160 8360
rect 12120 8310 12160 8340
rect 12120 8290 12130 8310
rect 12150 8290 12160 8310
rect 12120 8260 12160 8290
rect 12120 8240 12130 8260
rect 12150 8240 12160 8260
rect 12120 8210 12160 8240
rect 12120 8190 12130 8210
rect 12150 8190 12160 8210
rect 12120 8175 12160 8190
rect 12180 8560 12220 8575
rect 12180 8540 12190 8560
rect 12210 8540 12220 8560
rect 12180 8510 12220 8540
rect 12180 8490 12190 8510
rect 12210 8490 12220 8510
rect 12180 8460 12220 8490
rect 12180 8440 12190 8460
rect 12210 8440 12220 8460
rect 12180 8410 12220 8440
rect 12180 8390 12190 8410
rect 12210 8390 12220 8410
rect 12180 8360 12220 8390
rect 12180 8340 12190 8360
rect 12210 8340 12220 8360
rect 12180 8310 12220 8340
rect 12180 8290 12190 8310
rect 12210 8290 12220 8310
rect 12180 8260 12220 8290
rect 12180 8240 12190 8260
rect 12210 8240 12220 8260
rect 12180 8210 12220 8240
rect 12180 8190 12190 8210
rect 12210 8190 12220 8210
rect 12180 8175 12220 8190
rect 12240 8560 12280 8575
rect 12240 8540 12250 8560
rect 12270 8540 12280 8560
rect 12240 8510 12280 8540
rect 12240 8490 12250 8510
rect 12270 8490 12280 8510
rect 12240 8460 12280 8490
rect 12240 8440 12250 8460
rect 12270 8440 12280 8460
rect 12240 8410 12280 8440
rect 12240 8390 12250 8410
rect 12270 8390 12280 8410
rect 12240 8360 12280 8390
rect 12240 8340 12250 8360
rect 12270 8340 12280 8360
rect 12240 8310 12280 8340
rect 12240 8290 12250 8310
rect 12270 8290 12280 8310
rect 12240 8260 12280 8290
rect 12240 8240 12250 8260
rect 12270 8240 12280 8260
rect 12240 8210 12280 8240
rect 12240 8190 12250 8210
rect 12270 8190 12280 8210
rect 12240 8175 12280 8190
rect 12300 8560 12340 8575
rect 12300 8540 12310 8560
rect 12330 8540 12340 8560
rect 12300 8510 12340 8540
rect 12300 8490 12310 8510
rect 12330 8490 12340 8510
rect 12300 8460 12340 8490
rect 12300 8440 12310 8460
rect 12330 8440 12340 8460
rect 12300 8410 12340 8440
rect 12300 8390 12310 8410
rect 12330 8390 12340 8410
rect 12300 8360 12340 8390
rect 12300 8340 12310 8360
rect 12330 8340 12340 8360
rect 12300 8310 12340 8340
rect 12300 8290 12310 8310
rect 12330 8290 12340 8310
rect 12300 8260 12340 8290
rect 12300 8240 12310 8260
rect 12330 8240 12340 8260
rect 12300 8210 12340 8240
rect 12300 8190 12310 8210
rect 12330 8190 12340 8210
rect 12300 8175 12340 8190
rect 12360 8560 12400 8575
rect 12360 8540 12370 8560
rect 12390 8540 12400 8560
rect 12360 8510 12400 8540
rect 12360 8490 12370 8510
rect 12390 8490 12400 8510
rect 12360 8460 12400 8490
rect 12360 8440 12370 8460
rect 12390 8440 12400 8460
rect 12360 8410 12400 8440
rect 12360 8390 12370 8410
rect 12390 8390 12400 8410
rect 12360 8360 12400 8390
rect 12360 8340 12370 8360
rect 12390 8340 12400 8360
rect 12360 8310 12400 8340
rect 12360 8290 12370 8310
rect 12390 8290 12400 8310
rect 12360 8260 12400 8290
rect 12360 8240 12370 8260
rect 12390 8240 12400 8260
rect 12360 8210 12400 8240
rect 12360 8190 12370 8210
rect 12390 8190 12400 8210
rect 12360 8175 12400 8190
rect 12420 8560 12460 8575
rect 12420 8540 12430 8560
rect 12450 8540 12460 8560
rect 12420 8510 12460 8540
rect 12420 8490 12430 8510
rect 12450 8490 12460 8510
rect 12420 8460 12460 8490
rect 12420 8440 12430 8460
rect 12450 8440 12460 8460
rect 12420 8410 12460 8440
rect 12420 8390 12430 8410
rect 12450 8390 12460 8410
rect 12420 8360 12460 8390
rect 12420 8340 12430 8360
rect 12450 8340 12460 8360
rect 12420 8310 12460 8340
rect 12420 8290 12430 8310
rect 12450 8290 12460 8310
rect 12420 8260 12460 8290
rect 12420 8240 12430 8260
rect 12450 8240 12460 8260
rect 12420 8210 12460 8240
rect 12420 8190 12430 8210
rect 12450 8190 12460 8210
rect 12420 8175 12460 8190
rect 12480 8560 12520 8575
rect 12480 8540 12490 8560
rect 12510 8540 12520 8560
rect 12480 8510 12520 8540
rect 12480 8490 12490 8510
rect 12510 8490 12520 8510
rect 12480 8460 12520 8490
rect 12480 8440 12490 8460
rect 12510 8440 12520 8460
rect 12480 8410 12520 8440
rect 12480 8390 12490 8410
rect 12510 8390 12520 8410
rect 12480 8360 12520 8390
rect 12480 8340 12490 8360
rect 12510 8340 12520 8360
rect 12480 8310 12520 8340
rect 12480 8290 12490 8310
rect 12510 8290 12520 8310
rect 12480 8260 12520 8290
rect 12480 8240 12490 8260
rect 12510 8240 12520 8260
rect 12480 8210 12520 8240
rect 12480 8190 12490 8210
rect 12510 8190 12520 8210
rect 12480 8175 12520 8190
rect 12540 8560 12580 8575
rect 12540 8540 12550 8560
rect 12570 8540 12580 8560
rect 18455 8550 18480 8580
rect 12540 8510 12580 8540
rect 12540 8490 12550 8510
rect 12570 8490 12580 8510
rect 12540 8460 12580 8490
rect 12540 8440 12550 8460
rect 12570 8440 12580 8460
rect 12540 8410 12580 8440
rect 12540 8390 12550 8410
rect 12570 8390 12580 8410
rect 12540 8360 12580 8390
rect 12540 8340 12550 8360
rect 12570 8340 12580 8360
rect 18320 8515 18360 8550
rect 18320 8495 18330 8515
rect 18350 8495 18360 8515
rect 18320 8465 18360 8495
rect 18320 8445 18330 8465
rect 18350 8445 18360 8465
rect 18320 8415 18360 8445
rect 18320 8395 18330 8415
rect 18350 8395 18360 8415
rect 18320 8365 18360 8395
rect 12540 8310 12580 8340
rect 12540 8290 12550 8310
rect 12570 8290 12580 8310
rect 18320 8345 18330 8365
rect 18350 8345 18360 8365
rect 18320 8315 18360 8345
rect 18320 8295 18330 8315
rect 18350 8295 18360 8315
rect 12540 8260 12580 8290
rect 12540 8240 12550 8260
rect 12570 8240 12580 8260
rect 17990 8265 18030 8293
rect 17990 8245 18000 8265
rect 18020 8245 18030 8265
rect 12540 8210 12580 8240
rect 12540 8190 12550 8210
rect 12570 8190 12580 8210
rect 12540 8175 12580 8190
rect 12895 8225 12935 8240
rect 12895 8205 12905 8225
rect 12925 8205 12935 8225
rect 12895 8175 12935 8205
rect 12895 8155 12905 8175
rect 12925 8155 12935 8175
rect 12895 8125 12935 8155
rect 12895 8105 12905 8125
rect 12925 8105 12935 8125
rect 12895 8075 12935 8105
rect 12895 8055 12905 8075
rect 12925 8055 12935 8075
rect 12895 8025 12935 8055
rect 12895 8005 12905 8025
rect 12925 8005 12935 8025
rect 12895 7975 12935 8005
rect 12895 7955 12905 7975
rect 12925 7955 12935 7975
rect 12895 7940 12935 7955
rect 12950 8225 12990 8240
rect 12950 8205 12960 8225
rect 12980 8205 12990 8225
rect 12950 8175 12990 8205
rect 12950 8155 12960 8175
rect 12980 8155 12990 8175
rect 12950 8125 12990 8155
rect 12950 8105 12960 8125
rect 12980 8105 12990 8125
rect 12950 8075 12990 8105
rect 12950 8055 12960 8075
rect 12980 8055 12990 8075
rect 12950 8025 12990 8055
rect 12950 8005 12960 8025
rect 12980 8005 12990 8025
rect 12950 7975 12990 8005
rect 12950 7955 12960 7975
rect 12980 7955 12990 7975
rect 12950 7940 12990 7955
rect 13005 8225 13045 8240
rect 13005 8205 13015 8225
rect 13035 8205 13045 8225
rect 13005 8175 13045 8205
rect 13005 8155 13015 8175
rect 13035 8155 13045 8175
rect 13005 8125 13045 8155
rect 13005 8105 13015 8125
rect 13035 8105 13045 8125
rect 13005 8075 13045 8105
rect 13005 8055 13015 8075
rect 13035 8055 13045 8075
rect 13005 8025 13045 8055
rect 13005 8005 13015 8025
rect 13035 8005 13045 8025
rect 13005 7975 13045 8005
rect 13005 7955 13015 7975
rect 13035 7955 13045 7975
rect 13005 7940 13045 7955
rect 13060 8225 13100 8240
rect 13060 8205 13070 8225
rect 13090 8205 13100 8225
rect 13060 8175 13100 8205
rect 13060 8155 13070 8175
rect 13090 8155 13100 8175
rect 13060 8125 13100 8155
rect 13060 8105 13070 8125
rect 13090 8105 13100 8125
rect 13060 8075 13100 8105
rect 13060 8055 13070 8075
rect 13090 8055 13100 8075
rect 13060 8025 13100 8055
rect 13060 8005 13070 8025
rect 13090 8005 13100 8025
rect 13060 7975 13100 8005
rect 13060 7955 13070 7975
rect 13090 7955 13100 7975
rect 13060 7940 13100 7955
rect 13115 8225 13155 8240
rect 13115 8205 13125 8225
rect 13145 8205 13155 8225
rect 13115 8175 13155 8205
rect 13115 8155 13125 8175
rect 13145 8155 13155 8175
rect 13115 8125 13155 8155
rect 13115 8105 13125 8125
rect 13145 8105 13155 8125
rect 13115 8075 13155 8105
rect 13115 8055 13125 8075
rect 13145 8055 13155 8075
rect 13115 8025 13155 8055
rect 13115 8005 13125 8025
rect 13145 8005 13155 8025
rect 13115 7975 13155 8005
rect 13115 7955 13125 7975
rect 13145 7955 13155 7975
rect 13115 7940 13155 7955
rect 13170 8225 13210 8240
rect 13170 8205 13180 8225
rect 13200 8205 13210 8225
rect 13170 8175 13210 8205
rect 13170 8155 13180 8175
rect 13200 8155 13210 8175
rect 13170 8125 13210 8155
rect 13170 8105 13180 8125
rect 13200 8105 13210 8125
rect 13170 8075 13210 8105
rect 13170 8055 13180 8075
rect 13200 8055 13210 8075
rect 13170 8025 13210 8055
rect 13170 8005 13180 8025
rect 13200 8005 13210 8025
rect 13170 7975 13210 8005
rect 13170 7955 13180 7975
rect 13200 7955 13210 7975
rect 13170 7940 13210 7955
rect 13225 8225 13265 8240
rect 13225 8205 13235 8225
rect 13255 8205 13265 8225
rect 13225 8175 13265 8205
rect 13225 8155 13235 8175
rect 13255 8155 13265 8175
rect 13225 8125 13265 8155
rect 13225 8105 13235 8125
rect 13255 8105 13265 8125
rect 13225 8075 13265 8105
rect 13225 8055 13235 8075
rect 13255 8055 13265 8075
rect 13225 8025 13265 8055
rect 13225 8005 13235 8025
rect 13255 8005 13265 8025
rect 13225 7975 13265 8005
rect 13225 7955 13235 7975
rect 13255 7955 13265 7975
rect 13225 7940 13265 7955
rect 13280 8225 13320 8240
rect 13280 8205 13290 8225
rect 13310 8205 13320 8225
rect 13280 8175 13320 8205
rect 13280 8155 13290 8175
rect 13310 8155 13320 8175
rect 13280 8125 13320 8155
rect 13280 8105 13290 8125
rect 13310 8105 13320 8125
rect 13280 8075 13320 8105
rect 13280 8055 13290 8075
rect 13310 8055 13320 8075
rect 13280 8025 13320 8055
rect 13280 8005 13290 8025
rect 13310 8005 13320 8025
rect 13280 7975 13320 8005
rect 13280 7955 13290 7975
rect 13310 7955 13320 7975
rect 13280 7940 13320 7955
rect 13335 8225 13375 8240
rect 13335 8205 13345 8225
rect 13365 8205 13375 8225
rect 13335 8175 13375 8205
rect 13335 8155 13345 8175
rect 13365 8155 13375 8175
rect 13335 8125 13375 8155
rect 13335 8105 13345 8125
rect 13365 8105 13375 8125
rect 13335 8075 13375 8105
rect 13335 8055 13345 8075
rect 13365 8055 13375 8075
rect 13335 8025 13375 8055
rect 13335 8005 13345 8025
rect 13365 8005 13375 8025
rect 13335 7975 13375 8005
rect 13335 7955 13345 7975
rect 13365 7955 13375 7975
rect 13335 7940 13375 7955
rect 13390 8225 13430 8240
rect 13390 8205 13400 8225
rect 13420 8205 13430 8225
rect 13390 8175 13430 8205
rect 13390 8155 13400 8175
rect 13420 8155 13430 8175
rect 13390 8125 13430 8155
rect 13390 8105 13400 8125
rect 13420 8105 13430 8125
rect 13390 8075 13430 8105
rect 13390 8055 13400 8075
rect 13420 8055 13430 8075
rect 13390 8025 13430 8055
rect 13390 8005 13400 8025
rect 13420 8005 13430 8025
rect 13390 7975 13430 8005
rect 13390 7955 13400 7975
rect 13420 7955 13430 7975
rect 13390 7940 13430 7955
rect 13445 8225 13485 8240
rect 13445 8205 13455 8225
rect 13475 8205 13485 8225
rect 13445 8175 13485 8205
rect 13445 8155 13455 8175
rect 13475 8155 13485 8175
rect 13445 8125 13485 8155
rect 13445 8105 13455 8125
rect 13475 8105 13485 8125
rect 13445 8075 13485 8105
rect 13445 8055 13455 8075
rect 13475 8055 13485 8075
rect 13445 8025 13485 8055
rect 13445 8005 13455 8025
rect 13475 8005 13485 8025
rect 13445 7975 13485 8005
rect 13445 7955 13455 7975
rect 13475 7955 13485 7975
rect 13445 7940 13485 7955
rect 13500 8225 13540 8240
rect 13500 8205 13510 8225
rect 13530 8205 13540 8225
rect 13500 8175 13540 8205
rect 13500 8155 13510 8175
rect 13530 8155 13540 8175
rect 13500 8125 13540 8155
rect 13500 8105 13510 8125
rect 13530 8105 13540 8125
rect 13500 8075 13540 8105
rect 13500 8055 13510 8075
rect 13530 8055 13540 8075
rect 13500 8025 13540 8055
rect 13500 8005 13510 8025
rect 13530 8005 13540 8025
rect 13500 7975 13540 8005
rect 13500 7955 13510 7975
rect 13530 7955 13540 7975
rect 13500 7940 13540 7955
rect 13555 8225 13595 8240
rect 13555 8205 13565 8225
rect 13585 8205 13595 8225
rect 13555 8175 13595 8205
rect 13555 8155 13565 8175
rect 13585 8155 13595 8175
rect 13555 8125 13595 8155
rect 13555 8105 13565 8125
rect 13585 8105 13595 8125
rect 13555 8075 13595 8105
rect 13555 8055 13565 8075
rect 13585 8055 13595 8075
rect 13555 8025 13595 8055
rect 13555 8005 13565 8025
rect 13585 8005 13595 8025
rect 13555 7975 13595 8005
rect 13555 7955 13565 7975
rect 13585 7955 13595 7975
rect 13555 7940 13595 7955
rect 13610 8225 13650 8240
rect 13610 8205 13620 8225
rect 13640 8205 13650 8225
rect 13610 8175 13650 8205
rect 13610 8155 13620 8175
rect 13640 8155 13650 8175
rect 13610 8125 13650 8155
rect 13610 8105 13620 8125
rect 13640 8105 13650 8125
rect 13610 8075 13650 8105
rect 13610 8055 13620 8075
rect 13640 8055 13650 8075
rect 13610 8025 13650 8055
rect 13610 8005 13620 8025
rect 13640 8005 13650 8025
rect 13610 7975 13650 8005
rect 13610 7955 13620 7975
rect 13640 7955 13650 7975
rect 13610 7940 13650 7955
rect 13665 8225 13705 8240
rect 13665 8205 13675 8225
rect 13695 8205 13705 8225
rect 13665 8175 13705 8205
rect 13665 8155 13675 8175
rect 13695 8155 13705 8175
rect 13665 8125 13705 8155
rect 13665 8105 13675 8125
rect 13695 8105 13705 8125
rect 13665 8075 13705 8105
rect 13665 8055 13675 8075
rect 13695 8055 13705 8075
rect 13665 8025 13705 8055
rect 13665 8005 13675 8025
rect 13695 8005 13705 8025
rect 13665 7975 13705 8005
rect 13665 7955 13675 7975
rect 13695 7955 13705 7975
rect 13665 7940 13705 7955
rect 13720 8225 13760 8240
rect 13720 8205 13730 8225
rect 13750 8205 13760 8225
rect 13720 8175 13760 8205
rect 13720 8155 13730 8175
rect 13750 8155 13760 8175
rect 13720 8125 13760 8155
rect 13720 8105 13730 8125
rect 13750 8105 13760 8125
rect 13720 8075 13760 8105
rect 13720 8055 13730 8075
rect 13750 8055 13760 8075
rect 13720 8025 13760 8055
rect 13720 8005 13730 8025
rect 13750 8005 13760 8025
rect 13720 7975 13760 8005
rect 13720 7955 13730 7975
rect 13750 7955 13760 7975
rect 13720 7940 13760 7955
rect 13775 8225 13815 8240
rect 13775 8205 13785 8225
rect 13805 8205 13815 8225
rect 13775 8175 13815 8205
rect 13775 8155 13785 8175
rect 13805 8155 13815 8175
rect 13775 8125 13815 8155
rect 13775 8105 13785 8125
rect 13805 8105 13815 8125
rect 13775 8075 13815 8105
rect 13775 8055 13785 8075
rect 13805 8055 13815 8075
rect 13775 8025 13815 8055
rect 13775 8005 13785 8025
rect 13805 8005 13815 8025
rect 13775 7975 13815 8005
rect 13775 7955 13785 7975
rect 13805 7955 13815 7975
rect 13775 7940 13815 7955
rect 13830 8225 13870 8240
rect 13830 8205 13840 8225
rect 13860 8205 13870 8225
rect 13830 8175 13870 8205
rect 13830 8155 13840 8175
rect 13860 8155 13870 8175
rect 13830 8125 13870 8155
rect 13830 8105 13840 8125
rect 13860 8105 13870 8125
rect 13830 8075 13870 8105
rect 13830 8055 13840 8075
rect 13860 8055 13870 8075
rect 13830 8025 13870 8055
rect 13830 8005 13840 8025
rect 13860 8005 13870 8025
rect 13830 7975 13870 8005
rect 13830 7955 13840 7975
rect 13860 7955 13870 7975
rect 13830 7940 13870 7955
rect 13885 8225 13925 8240
rect 13885 8205 13895 8225
rect 13915 8205 13925 8225
rect 13885 8175 13925 8205
rect 13885 8155 13895 8175
rect 13915 8155 13925 8175
rect 13885 8125 13925 8155
rect 13885 8105 13895 8125
rect 13915 8105 13925 8125
rect 13885 8075 13925 8105
rect 13885 8055 13895 8075
rect 13915 8055 13925 8075
rect 13885 8025 13925 8055
rect 13885 8005 13895 8025
rect 13915 8005 13925 8025
rect 13885 7975 13925 8005
rect 13885 7955 13895 7975
rect 13915 7955 13925 7975
rect 13885 7940 13925 7955
rect 13940 8225 13980 8240
rect 13940 8205 13950 8225
rect 13970 8205 13980 8225
rect 13940 8175 13980 8205
rect 13940 8155 13950 8175
rect 13970 8155 13980 8175
rect 13940 8125 13980 8155
rect 13940 8105 13950 8125
rect 13970 8105 13980 8125
rect 13940 8075 13980 8105
rect 13940 8055 13950 8075
rect 13970 8055 13980 8075
rect 13940 8025 13980 8055
rect 13940 8005 13950 8025
rect 13970 8005 13980 8025
rect 13940 7975 13980 8005
rect 13940 7955 13950 7975
rect 13970 7955 13980 7975
rect 13940 7940 13980 7955
rect 13995 8225 14035 8240
rect 13995 8205 14005 8225
rect 14025 8205 14035 8225
rect 13995 8175 14035 8205
rect 13995 8155 14005 8175
rect 14025 8155 14035 8175
rect 13995 8125 14035 8155
rect 13995 8105 14005 8125
rect 14025 8105 14035 8125
rect 13995 8075 14035 8105
rect 13995 8055 14005 8075
rect 14025 8055 14035 8075
rect 13995 8025 14035 8055
rect 13995 8005 14005 8025
rect 14025 8005 14035 8025
rect 13995 7975 14035 8005
rect 13995 7955 14005 7975
rect 14025 7955 14035 7975
rect 13995 7940 14035 7955
rect 14050 8225 14090 8240
rect 14050 8205 14060 8225
rect 14080 8205 14090 8225
rect 14050 8175 14090 8205
rect 14050 8155 14060 8175
rect 14080 8155 14090 8175
rect 14050 8125 14090 8155
rect 14050 8105 14060 8125
rect 14080 8105 14090 8125
rect 14050 8075 14090 8105
rect 14050 8055 14060 8075
rect 14080 8055 14090 8075
rect 14050 8025 14090 8055
rect 14050 8005 14060 8025
rect 14080 8005 14090 8025
rect 14050 7975 14090 8005
rect 14050 7955 14060 7975
rect 14080 7955 14090 7975
rect 14050 7940 14090 7955
rect 14105 8225 14145 8240
rect 17990 8230 18030 8245
rect 18050 8270 18090 8293
rect 18050 8250 18060 8270
rect 18080 8250 18090 8270
rect 18050 8230 18090 8250
rect 18110 8270 18150 8293
rect 18110 8250 18120 8270
rect 18140 8250 18150 8270
rect 18110 8230 18150 8250
rect 18170 8265 18210 8293
rect 18170 8245 18180 8265
rect 18200 8245 18210 8265
rect 18170 8230 18210 8245
rect 18320 8265 18360 8295
rect 18320 8245 18330 8265
rect 18350 8245 18360 8265
rect 18320 8230 18360 8245
rect 18380 8515 18420 8550
rect 18380 8495 18390 8515
rect 18410 8495 18420 8515
rect 18380 8465 18420 8495
rect 18380 8445 18390 8465
rect 18410 8445 18420 8465
rect 18380 8415 18420 8445
rect 18380 8395 18390 8415
rect 18410 8395 18420 8415
rect 18380 8365 18420 8395
rect 18380 8345 18390 8365
rect 18410 8345 18420 8365
rect 18380 8315 18420 8345
rect 18380 8295 18390 8315
rect 18410 8295 18420 8315
rect 18380 8265 18420 8295
rect 18380 8245 18390 8265
rect 18410 8245 18420 8265
rect 18380 8230 18420 8245
rect 18440 8515 18480 8550
rect 18440 8495 18450 8515
rect 18470 8495 18480 8515
rect 18440 8465 18480 8495
rect 18440 8445 18450 8465
rect 18470 8445 18480 8465
rect 18440 8415 18480 8445
rect 18440 8395 18450 8415
rect 18470 8395 18480 8415
rect 18440 8365 18480 8395
rect 18440 8345 18450 8365
rect 18470 8345 18480 8365
rect 18440 8315 18480 8345
rect 18440 8295 18450 8315
rect 18470 8295 18480 8315
rect 18440 8265 18480 8295
rect 18440 8245 18450 8265
rect 18470 8245 18480 8265
rect 18440 8230 18480 8245
rect 18500 8565 18540 8580
rect 18500 8545 18510 8565
rect 18530 8545 18540 8565
rect 18500 8515 18540 8545
rect 18500 8495 18510 8515
rect 18530 8495 18540 8515
rect 18500 8465 18540 8495
rect 18500 8445 18510 8465
rect 18530 8445 18540 8465
rect 18500 8415 18540 8445
rect 18500 8395 18510 8415
rect 18530 8395 18540 8415
rect 18500 8365 18540 8395
rect 18500 8345 18510 8365
rect 18530 8345 18540 8365
rect 18500 8315 18540 8345
rect 18500 8295 18510 8315
rect 18530 8295 18540 8315
rect 18500 8265 18540 8295
rect 18500 8245 18510 8265
rect 18530 8245 18540 8265
rect 18500 8230 18540 8245
rect 18560 8565 18600 8580
rect 18560 8545 18570 8565
rect 18590 8545 18600 8565
rect 18560 8515 18600 8545
rect 18560 8495 18570 8515
rect 18590 8495 18600 8515
rect 18560 8465 18600 8495
rect 18560 8445 18570 8465
rect 18590 8445 18600 8465
rect 18560 8415 18600 8445
rect 18560 8395 18570 8415
rect 18590 8395 18600 8415
rect 18560 8365 18600 8395
rect 18560 8345 18570 8365
rect 18590 8345 18600 8365
rect 18560 8315 18600 8345
rect 18560 8295 18570 8315
rect 18590 8295 18600 8315
rect 18560 8265 18600 8295
rect 18560 8245 18570 8265
rect 18590 8245 18600 8265
rect 18560 8230 18600 8245
rect 18720 8560 18760 8575
rect 18720 8540 18730 8560
rect 18750 8540 18760 8560
rect 18720 8510 18760 8540
rect 18720 8490 18730 8510
rect 18750 8490 18760 8510
rect 18720 8460 18760 8490
rect 18720 8440 18730 8460
rect 18750 8440 18760 8460
rect 18720 8410 18760 8440
rect 18720 8390 18730 8410
rect 18750 8390 18760 8410
rect 18720 8360 18760 8390
rect 18720 8340 18730 8360
rect 18750 8340 18760 8360
rect 18720 8310 18760 8340
rect 18720 8290 18730 8310
rect 18750 8290 18760 8310
rect 18720 8260 18760 8290
rect 18720 8240 18730 8260
rect 18750 8240 18760 8260
rect 14105 8205 14115 8225
rect 14135 8205 14145 8225
rect 14105 8175 14145 8205
rect 18720 8210 18760 8240
rect 18720 8190 18730 8210
rect 18750 8190 18760 8210
rect 18720 8175 18760 8190
rect 18780 8560 18820 8575
rect 18780 8540 18790 8560
rect 18810 8540 18820 8560
rect 18780 8510 18820 8540
rect 18780 8490 18790 8510
rect 18810 8490 18820 8510
rect 18780 8460 18820 8490
rect 18780 8440 18790 8460
rect 18810 8440 18820 8460
rect 18780 8410 18820 8440
rect 18780 8390 18790 8410
rect 18810 8390 18820 8410
rect 18780 8360 18820 8390
rect 18780 8340 18790 8360
rect 18810 8340 18820 8360
rect 18780 8310 18820 8340
rect 18780 8290 18790 8310
rect 18810 8290 18820 8310
rect 18780 8260 18820 8290
rect 18780 8240 18790 8260
rect 18810 8240 18820 8260
rect 18780 8210 18820 8240
rect 18780 8190 18790 8210
rect 18810 8190 18820 8210
rect 18780 8175 18820 8190
rect 18840 8560 18880 8575
rect 18840 8540 18850 8560
rect 18870 8540 18880 8560
rect 18840 8510 18880 8540
rect 18840 8490 18850 8510
rect 18870 8490 18880 8510
rect 18840 8460 18880 8490
rect 18840 8440 18850 8460
rect 18870 8440 18880 8460
rect 18840 8410 18880 8440
rect 18840 8390 18850 8410
rect 18870 8390 18880 8410
rect 18840 8360 18880 8390
rect 18840 8340 18850 8360
rect 18870 8340 18880 8360
rect 18840 8310 18880 8340
rect 18840 8290 18850 8310
rect 18870 8290 18880 8310
rect 18840 8260 18880 8290
rect 18840 8240 18850 8260
rect 18870 8240 18880 8260
rect 18840 8210 18880 8240
rect 18840 8190 18850 8210
rect 18870 8190 18880 8210
rect 18840 8175 18880 8190
rect 18900 8560 18940 8575
rect 18900 8540 18910 8560
rect 18930 8540 18940 8560
rect 18900 8510 18940 8540
rect 18900 8490 18910 8510
rect 18930 8490 18940 8510
rect 18900 8460 18940 8490
rect 18900 8440 18910 8460
rect 18930 8440 18940 8460
rect 18900 8410 18940 8440
rect 18900 8390 18910 8410
rect 18930 8390 18940 8410
rect 18900 8360 18940 8390
rect 18900 8340 18910 8360
rect 18930 8340 18940 8360
rect 18900 8310 18940 8340
rect 18900 8290 18910 8310
rect 18930 8290 18940 8310
rect 18900 8260 18940 8290
rect 18900 8240 18910 8260
rect 18930 8240 18940 8260
rect 18900 8210 18940 8240
rect 18900 8190 18910 8210
rect 18930 8190 18940 8210
rect 18900 8175 18940 8190
rect 18960 8560 19000 8575
rect 18960 8540 18970 8560
rect 18990 8540 19000 8560
rect 18960 8510 19000 8540
rect 18960 8490 18970 8510
rect 18990 8490 19000 8510
rect 18960 8460 19000 8490
rect 18960 8440 18970 8460
rect 18990 8440 19000 8460
rect 18960 8410 19000 8440
rect 18960 8390 18970 8410
rect 18990 8390 19000 8410
rect 18960 8360 19000 8390
rect 18960 8340 18970 8360
rect 18990 8340 19000 8360
rect 18960 8310 19000 8340
rect 18960 8290 18970 8310
rect 18990 8290 19000 8310
rect 18960 8260 19000 8290
rect 18960 8240 18970 8260
rect 18990 8240 19000 8260
rect 18960 8210 19000 8240
rect 18960 8190 18970 8210
rect 18990 8190 19000 8210
rect 18960 8175 19000 8190
rect 19020 8560 19060 8575
rect 19020 8540 19030 8560
rect 19050 8540 19060 8560
rect 19020 8510 19060 8540
rect 19020 8490 19030 8510
rect 19050 8490 19060 8510
rect 19020 8460 19060 8490
rect 19020 8440 19030 8460
rect 19050 8440 19060 8460
rect 19020 8410 19060 8440
rect 19020 8390 19030 8410
rect 19050 8390 19060 8410
rect 19020 8360 19060 8390
rect 19020 8340 19030 8360
rect 19050 8340 19060 8360
rect 19020 8310 19060 8340
rect 19020 8290 19030 8310
rect 19050 8290 19060 8310
rect 19020 8260 19060 8290
rect 19020 8240 19030 8260
rect 19050 8240 19060 8260
rect 19020 8210 19060 8240
rect 19020 8190 19030 8210
rect 19050 8190 19060 8210
rect 19020 8175 19060 8190
rect 19080 8560 19120 8575
rect 19080 8540 19090 8560
rect 19110 8540 19120 8560
rect 19080 8510 19120 8540
rect 19080 8490 19090 8510
rect 19110 8490 19120 8510
rect 19080 8460 19120 8490
rect 19080 8440 19090 8460
rect 19110 8440 19120 8460
rect 19080 8410 19120 8440
rect 19080 8390 19090 8410
rect 19110 8390 19120 8410
rect 19080 8360 19120 8390
rect 19080 8340 19090 8360
rect 19110 8340 19120 8360
rect 19080 8310 19120 8340
rect 19080 8290 19090 8310
rect 19110 8290 19120 8310
rect 19080 8260 19120 8290
rect 19080 8240 19090 8260
rect 19110 8240 19120 8260
rect 19080 8210 19120 8240
rect 19080 8190 19090 8210
rect 19110 8190 19120 8210
rect 19080 8175 19120 8190
rect 19140 8560 19180 8575
rect 19140 8540 19150 8560
rect 19170 8540 19180 8560
rect 19140 8510 19180 8540
rect 19140 8490 19150 8510
rect 19170 8490 19180 8510
rect 19140 8460 19180 8490
rect 19140 8440 19150 8460
rect 19170 8440 19180 8460
rect 19140 8410 19180 8440
rect 19140 8390 19150 8410
rect 19170 8390 19180 8410
rect 19140 8360 19180 8390
rect 19140 8340 19150 8360
rect 19170 8340 19180 8360
rect 19140 8310 19180 8340
rect 19140 8290 19150 8310
rect 19170 8290 19180 8310
rect 19140 8260 19180 8290
rect 19140 8240 19150 8260
rect 19170 8240 19180 8260
rect 19140 8210 19180 8240
rect 19140 8190 19150 8210
rect 19170 8190 19180 8210
rect 19140 8175 19180 8190
rect 19200 8560 19240 8575
rect 19200 8540 19210 8560
rect 19230 8540 19240 8560
rect 19200 8510 19240 8540
rect 19200 8490 19210 8510
rect 19230 8490 19240 8510
rect 19200 8460 19240 8490
rect 19200 8440 19210 8460
rect 19230 8440 19240 8460
rect 19200 8410 19240 8440
rect 19200 8390 19210 8410
rect 19230 8390 19240 8410
rect 19200 8360 19240 8390
rect 19200 8340 19210 8360
rect 19230 8340 19240 8360
rect 19200 8310 19240 8340
rect 19200 8290 19210 8310
rect 19230 8290 19240 8310
rect 19200 8260 19240 8290
rect 19200 8240 19210 8260
rect 19230 8240 19240 8260
rect 19200 8210 19240 8240
rect 19200 8190 19210 8210
rect 19230 8190 19240 8210
rect 19200 8175 19240 8190
rect 19260 8560 19300 8575
rect 19260 8540 19270 8560
rect 19290 8540 19300 8560
rect 19260 8510 19300 8540
rect 19260 8490 19270 8510
rect 19290 8490 19300 8510
rect 19260 8460 19300 8490
rect 19260 8440 19270 8460
rect 19290 8440 19300 8460
rect 19260 8410 19300 8440
rect 19260 8390 19270 8410
rect 19290 8390 19300 8410
rect 19260 8360 19300 8390
rect 19260 8340 19270 8360
rect 19290 8340 19300 8360
rect 19260 8310 19300 8340
rect 19260 8290 19270 8310
rect 19290 8290 19300 8310
rect 19260 8260 19300 8290
rect 19260 8240 19270 8260
rect 19290 8240 19300 8260
rect 19260 8210 19300 8240
rect 19260 8190 19270 8210
rect 19290 8190 19300 8210
rect 19260 8175 19300 8190
rect 19320 8560 19360 8575
rect 19320 8540 19330 8560
rect 19350 8540 19360 8560
rect 19320 8510 19360 8540
rect 19320 8490 19330 8510
rect 19350 8490 19360 8510
rect 19320 8460 19360 8490
rect 19320 8440 19330 8460
rect 19350 8440 19360 8460
rect 19320 8410 19360 8440
rect 19320 8390 19330 8410
rect 19350 8390 19360 8410
rect 19320 8360 19360 8390
rect 19320 8340 19330 8360
rect 19350 8340 19360 8360
rect 19320 8310 19360 8340
rect 19320 8290 19330 8310
rect 19350 8290 19360 8310
rect 19320 8260 19360 8290
rect 19320 8240 19330 8260
rect 19350 8240 19360 8260
rect 19320 8210 19360 8240
rect 19320 8190 19330 8210
rect 19350 8190 19360 8210
rect 19320 8175 19360 8190
rect 19380 8560 19420 8575
rect 19380 8540 19390 8560
rect 19410 8540 19420 8560
rect 19380 8510 19420 8540
rect 19380 8490 19390 8510
rect 19410 8490 19420 8510
rect 19380 8460 19420 8490
rect 19380 8440 19390 8460
rect 19410 8440 19420 8460
rect 19380 8410 19420 8440
rect 19380 8390 19390 8410
rect 19410 8390 19420 8410
rect 19380 8360 19420 8390
rect 19380 8340 19390 8360
rect 19410 8340 19420 8360
rect 19380 8310 19420 8340
rect 19380 8290 19390 8310
rect 19410 8290 19420 8310
rect 19380 8260 19420 8290
rect 19380 8240 19390 8260
rect 19410 8240 19420 8260
rect 19380 8210 19420 8240
rect 19380 8190 19390 8210
rect 19410 8190 19420 8210
rect 19380 8175 19420 8190
rect 19440 8560 19480 8575
rect 19440 8540 19450 8560
rect 19470 8540 19480 8560
rect 19440 8510 19480 8540
rect 19440 8490 19450 8510
rect 19470 8490 19480 8510
rect 19440 8460 19480 8490
rect 19440 8440 19450 8460
rect 19470 8440 19480 8460
rect 19440 8410 19480 8440
rect 19440 8390 19450 8410
rect 19470 8390 19480 8410
rect 19440 8360 19480 8390
rect 19440 8340 19450 8360
rect 19470 8340 19480 8360
rect 19440 8310 19480 8340
rect 19440 8290 19450 8310
rect 19470 8290 19480 8310
rect 19440 8260 19480 8290
rect 19440 8240 19450 8260
rect 19470 8240 19480 8260
rect 19440 8210 19480 8240
rect 19440 8190 19450 8210
rect 19470 8190 19480 8210
rect 19440 8175 19480 8190
rect 19500 8560 19540 8575
rect 19500 8540 19510 8560
rect 19530 8540 19540 8560
rect 19500 8510 19540 8540
rect 19500 8490 19510 8510
rect 19530 8490 19540 8510
rect 19500 8460 19540 8490
rect 19500 8440 19510 8460
rect 19530 8440 19540 8460
rect 19500 8410 19540 8440
rect 19500 8390 19510 8410
rect 19530 8390 19540 8410
rect 19500 8360 19540 8390
rect 19500 8340 19510 8360
rect 19530 8340 19540 8360
rect 19500 8310 19540 8340
rect 19500 8290 19510 8310
rect 19530 8290 19540 8310
rect 19500 8260 19540 8290
rect 19500 8240 19510 8260
rect 19530 8240 19540 8260
rect 19500 8210 19540 8240
rect 19500 8190 19510 8210
rect 19530 8190 19540 8210
rect 19500 8175 19540 8190
rect 19560 8560 19600 8575
rect 19560 8540 19570 8560
rect 19590 8540 19600 8560
rect 19560 8510 19600 8540
rect 19560 8490 19570 8510
rect 19590 8490 19600 8510
rect 19560 8460 19600 8490
rect 19560 8440 19570 8460
rect 19590 8440 19600 8460
rect 19560 8410 19600 8440
rect 19560 8390 19570 8410
rect 19590 8390 19600 8410
rect 19560 8360 19600 8390
rect 19560 8340 19570 8360
rect 19590 8340 19600 8360
rect 19560 8310 19600 8340
rect 19560 8290 19570 8310
rect 19590 8290 19600 8310
rect 19560 8260 19600 8290
rect 19560 8240 19570 8260
rect 19590 8240 19600 8260
rect 19560 8210 19600 8240
rect 19560 8190 19570 8210
rect 19590 8190 19600 8210
rect 19560 8175 19600 8190
rect 19620 8560 19660 8575
rect 19620 8540 19630 8560
rect 19650 8540 19660 8560
rect 19620 8510 19660 8540
rect 19620 8490 19630 8510
rect 19650 8490 19660 8510
rect 19620 8460 19660 8490
rect 19620 8440 19630 8460
rect 19650 8440 19660 8460
rect 19620 8410 19660 8440
rect 19620 8390 19630 8410
rect 19650 8390 19660 8410
rect 19620 8360 19660 8390
rect 19620 8340 19630 8360
rect 19650 8340 19660 8360
rect 19620 8310 19660 8340
rect 19620 8290 19630 8310
rect 19650 8290 19660 8310
rect 19620 8260 19660 8290
rect 19620 8240 19630 8260
rect 19650 8240 19660 8260
rect 19620 8210 19660 8240
rect 19620 8190 19630 8210
rect 19650 8190 19660 8210
rect 19620 8175 19660 8190
rect 19680 8560 19720 8575
rect 19680 8540 19690 8560
rect 19710 8540 19720 8560
rect 19680 8510 19720 8540
rect 19680 8490 19690 8510
rect 19710 8490 19720 8510
rect 19680 8460 19720 8490
rect 19680 8440 19690 8460
rect 19710 8440 19720 8460
rect 19680 8410 19720 8440
rect 19680 8390 19690 8410
rect 19710 8390 19720 8410
rect 19680 8360 19720 8390
rect 19680 8340 19690 8360
rect 19710 8340 19720 8360
rect 19680 8310 19720 8340
rect 19680 8290 19690 8310
rect 19710 8290 19720 8310
rect 19680 8260 19720 8290
rect 19680 8240 19690 8260
rect 19710 8240 19720 8260
rect 19680 8210 19720 8240
rect 19680 8190 19690 8210
rect 19710 8190 19720 8210
rect 19680 8175 19720 8190
rect 19740 8560 19780 8575
rect 19740 8540 19750 8560
rect 19770 8540 19780 8560
rect 19740 8510 19780 8540
rect 19740 8490 19750 8510
rect 19770 8490 19780 8510
rect 19740 8460 19780 8490
rect 19740 8440 19750 8460
rect 19770 8440 19780 8460
rect 19740 8410 19780 8440
rect 19740 8390 19750 8410
rect 19770 8390 19780 8410
rect 19740 8360 19780 8390
rect 19740 8340 19750 8360
rect 19770 8340 19780 8360
rect 19740 8310 19780 8340
rect 19740 8290 19750 8310
rect 19770 8290 19780 8310
rect 19740 8260 19780 8290
rect 19740 8240 19750 8260
rect 19770 8240 19780 8260
rect 19740 8210 19780 8240
rect 19740 8190 19750 8210
rect 19770 8190 19780 8210
rect 19740 8175 19780 8190
rect 19800 8560 19840 8575
rect 19800 8540 19810 8560
rect 19830 8540 19840 8560
rect 19800 8510 19840 8540
rect 19800 8490 19810 8510
rect 19830 8490 19840 8510
rect 19800 8460 19840 8490
rect 19800 8440 19810 8460
rect 19830 8440 19840 8460
rect 19800 8410 19840 8440
rect 19800 8390 19810 8410
rect 19830 8390 19840 8410
rect 19800 8360 19840 8390
rect 19800 8340 19810 8360
rect 19830 8340 19840 8360
rect 19800 8310 19840 8340
rect 19800 8290 19810 8310
rect 19830 8290 19840 8310
rect 19800 8260 19840 8290
rect 19800 8240 19810 8260
rect 19830 8240 19840 8260
rect 19800 8210 19840 8240
rect 19800 8190 19810 8210
rect 19830 8190 19840 8210
rect 19800 8175 19840 8190
rect 19860 8560 19900 8575
rect 19860 8540 19870 8560
rect 19890 8540 19900 8560
rect 19860 8510 19900 8540
rect 19860 8490 19870 8510
rect 19890 8490 19900 8510
rect 19860 8460 19900 8490
rect 19860 8440 19870 8460
rect 19890 8440 19900 8460
rect 19860 8410 19900 8440
rect 19860 8390 19870 8410
rect 19890 8390 19900 8410
rect 19860 8360 19900 8390
rect 19860 8340 19870 8360
rect 19890 8340 19900 8360
rect 19860 8310 19900 8340
rect 19860 8290 19870 8310
rect 19890 8290 19900 8310
rect 19860 8260 19900 8290
rect 19860 8240 19870 8260
rect 19890 8240 19900 8260
rect 19860 8210 19900 8240
rect 19860 8190 19870 8210
rect 19890 8190 19900 8210
rect 19860 8175 19900 8190
rect 19920 8560 19960 8575
rect 19920 8540 19930 8560
rect 19950 8540 19960 8560
rect 19920 8510 19960 8540
rect 19920 8490 19930 8510
rect 19950 8490 19960 8510
rect 19920 8460 19960 8490
rect 19920 8440 19930 8460
rect 19950 8440 19960 8460
rect 19920 8410 19960 8440
rect 19920 8390 19930 8410
rect 19950 8390 19960 8410
rect 19920 8360 19960 8390
rect 19920 8340 19930 8360
rect 19950 8340 19960 8360
rect 19920 8310 19960 8340
rect 19920 8290 19930 8310
rect 19950 8290 19960 8310
rect 19920 8260 19960 8290
rect 19920 8240 19930 8260
rect 19950 8240 19960 8260
rect 19920 8210 19960 8240
rect 19920 8190 19930 8210
rect 19950 8190 19960 8210
rect 19920 8175 19960 8190
rect 19980 8560 20020 8575
rect 19980 8540 19990 8560
rect 20010 8540 20020 8560
rect 19980 8510 20020 8540
rect 19980 8490 19990 8510
rect 20010 8490 20020 8510
rect 19980 8460 20020 8490
rect 19980 8440 19990 8460
rect 20010 8440 20020 8460
rect 19980 8410 20020 8440
rect 19980 8390 19990 8410
rect 20010 8390 20020 8410
rect 19980 8360 20020 8390
rect 19980 8340 19990 8360
rect 20010 8340 20020 8360
rect 19980 8310 20020 8340
rect 19980 8290 19990 8310
rect 20010 8290 20020 8310
rect 19980 8260 20020 8290
rect 19980 8240 19990 8260
rect 20010 8240 20020 8260
rect 19980 8210 20020 8240
rect 19980 8190 19990 8210
rect 20010 8190 20020 8210
rect 19980 8175 20020 8190
rect 20040 8560 20080 8575
rect 20040 8540 20050 8560
rect 20070 8540 20080 8560
rect 20040 8510 20080 8540
rect 20040 8490 20050 8510
rect 20070 8490 20080 8510
rect 20040 8460 20080 8490
rect 20040 8440 20050 8460
rect 20070 8440 20080 8460
rect 20040 8410 20080 8440
rect 20040 8390 20050 8410
rect 20070 8390 20080 8410
rect 20040 8360 20080 8390
rect 20040 8340 20050 8360
rect 20070 8340 20080 8360
rect 20040 8310 20080 8340
rect 20040 8290 20050 8310
rect 20070 8290 20080 8310
rect 20040 8260 20080 8290
rect 20040 8240 20050 8260
rect 20070 8240 20080 8260
rect 20040 8210 20080 8240
rect 20040 8190 20050 8210
rect 20070 8190 20080 8210
rect 20040 8175 20080 8190
rect 20390 8225 20430 8240
rect 20390 8205 20400 8225
rect 20420 8205 20430 8225
rect 20390 8175 20430 8205
rect 14105 8155 14115 8175
rect 14135 8155 14145 8175
rect 14105 8125 14145 8155
rect 20390 8155 20400 8175
rect 20420 8155 20430 8175
rect 14105 8105 14115 8125
rect 14135 8105 14145 8125
rect 20390 8125 20430 8155
rect 14105 8075 14145 8105
rect 14105 8055 14115 8075
rect 14135 8055 14145 8075
rect 14105 8025 14145 8055
rect 14105 8005 14115 8025
rect 14135 8005 14145 8025
rect 14105 7975 14145 8005
rect 14105 7955 14115 7975
rect 14135 7955 14145 7975
rect 14105 7940 14145 7955
rect 20390 8105 20400 8125
rect 20420 8105 20430 8125
rect 20390 8075 20430 8105
rect 20390 8055 20400 8075
rect 20420 8055 20430 8075
rect 20390 8025 20430 8055
rect 20390 8005 20400 8025
rect 20420 8005 20430 8025
rect 20390 7975 20430 8005
rect 20390 7955 20400 7975
rect 20420 7955 20430 7975
rect 11220 7880 11260 7895
rect 11220 7860 11230 7880
rect 11250 7860 11260 7880
rect 11220 7830 11260 7860
rect 11220 7810 11230 7830
rect 11250 7810 11260 7830
rect 11220 7780 11260 7810
rect 11220 7760 11230 7780
rect 11250 7760 11260 7780
rect 11220 7730 11260 7760
rect 11220 7710 11230 7730
rect 11250 7710 11260 7730
rect 11220 7680 11260 7710
rect 11220 7660 11230 7680
rect 11250 7660 11260 7680
rect 11220 7630 11260 7660
rect 9680 7605 9720 7620
rect 9680 7585 9690 7605
rect 9710 7585 9720 7605
rect 9680 7555 9720 7585
rect 9680 7535 9690 7555
rect 9710 7535 9720 7555
rect 9680 7520 9720 7535
rect 9735 7605 9775 7620
rect 9735 7585 9745 7605
rect 9765 7585 9775 7605
rect 9735 7555 9775 7585
rect 9735 7535 9745 7555
rect 9765 7535 9775 7555
rect 9735 7520 9775 7535
rect 9790 7605 9830 7620
rect 9790 7585 9800 7605
rect 9820 7585 9830 7605
rect 9790 7555 9830 7585
rect 9790 7535 9800 7555
rect 9820 7535 9830 7555
rect 9790 7520 9830 7535
rect 9845 7605 9885 7620
rect 9845 7585 9855 7605
rect 9875 7585 9885 7605
rect 9845 7555 9885 7585
rect 9845 7535 9855 7555
rect 9875 7535 9885 7555
rect 9845 7520 9885 7535
rect 9900 7605 9940 7620
rect 9900 7585 9910 7605
rect 9930 7585 9940 7605
rect 9900 7555 9940 7585
rect 9900 7535 9910 7555
rect 9930 7535 9940 7555
rect 9900 7520 9940 7535
rect 9955 7605 9995 7620
rect 9955 7585 9965 7605
rect 9985 7585 9995 7605
rect 9955 7555 9995 7585
rect 9955 7535 9965 7555
rect 9985 7535 9995 7555
rect 9955 7520 9995 7535
rect 10010 7605 10050 7620
rect 10010 7585 10020 7605
rect 10040 7585 10050 7605
rect 10010 7555 10050 7585
rect 10010 7535 10020 7555
rect 10040 7535 10050 7555
rect 10010 7520 10050 7535
rect 10065 7605 10105 7620
rect 10065 7585 10075 7605
rect 10095 7585 10105 7605
rect 10065 7555 10105 7585
rect 10065 7535 10075 7555
rect 10095 7535 10105 7555
rect 10065 7520 10105 7535
rect 10120 7605 10160 7620
rect 10120 7585 10130 7605
rect 10150 7585 10160 7605
rect 10120 7555 10160 7585
rect 10120 7535 10130 7555
rect 10150 7535 10160 7555
rect 10120 7520 10160 7535
rect 10175 7605 10215 7620
rect 10175 7585 10185 7605
rect 10205 7585 10215 7605
rect 10175 7555 10215 7585
rect 10175 7535 10185 7555
rect 10205 7535 10215 7555
rect 10175 7520 10215 7535
rect 10230 7605 10270 7620
rect 10230 7585 10240 7605
rect 10260 7585 10270 7605
rect 10230 7555 10270 7585
rect 10230 7535 10240 7555
rect 10260 7535 10270 7555
rect 10230 7520 10270 7535
rect 10285 7605 10325 7620
rect 10285 7585 10295 7605
rect 10315 7585 10325 7605
rect 10285 7555 10325 7585
rect 10285 7535 10295 7555
rect 10315 7535 10325 7555
rect 10285 7520 10325 7535
rect 10340 7605 10380 7620
rect 10340 7585 10350 7605
rect 10370 7585 10380 7605
rect 10340 7555 10380 7585
rect 10340 7535 10350 7555
rect 10370 7535 10380 7555
rect 10340 7520 10380 7535
rect 10395 7605 10435 7620
rect 10395 7585 10405 7605
rect 10425 7585 10435 7605
rect 10395 7555 10435 7585
rect 10395 7535 10405 7555
rect 10425 7535 10435 7555
rect 10395 7520 10435 7535
rect 10450 7605 10490 7620
rect 10450 7585 10460 7605
rect 10480 7585 10490 7605
rect 10450 7555 10490 7585
rect 10450 7535 10460 7555
rect 10480 7535 10490 7555
rect 10450 7520 10490 7535
rect 10505 7605 10545 7620
rect 10505 7585 10515 7605
rect 10535 7585 10545 7605
rect 10505 7555 10545 7585
rect 10505 7535 10515 7555
rect 10535 7535 10545 7555
rect 10505 7520 10545 7535
rect 10560 7605 10600 7620
rect 10560 7585 10570 7605
rect 10590 7585 10600 7605
rect 10560 7555 10600 7585
rect 10560 7535 10570 7555
rect 10590 7535 10600 7555
rect 10560 7520 10600 7535
rect 10615 7605 10655 7620
rect 10615 7585 10625 7605
rect 10645 7585 10655 7605
rect 10615 7555 10655 7585
rect 10615 7535 10625 7555
rect 10645 7535 10655 7555
rect 10615 7520 10655 7535
rect 10670 7605 10710 7620
rect 10670 7585 10680 7605
rect 10700 7585 10710 7605
rect 10670 7555 10710 7585
rect 10670 7535 10680 7555
rect 10700 7535 10710 7555
rect 10670 7520 10710 7535
rect 10725 7605 10765 7620
rect 10725 7585 10735 7605
rect 10755 7585 10765 7605
rect 10725 7555 10765 7585
rect 10725 7535 10735 7555
rect 10755 7535 10765 7555
rect 10725 7520 10765 7535
rect 10780 7605 10820 7620
rect 10780 7585 10790 7605
rect 10810 7585 10820 7605
rect 10780 7555 10820 7585
rect 10780 7535 10790 7555
rect 10810 7535 10820 7555
rect 10780 7520 10820 7535
rect 10835 7605 10875 7620
rect 10835 7585 10845 7605
rect 10865 7585 10875 7605
rect 10835 7555 10875 7585
rect 10835 7535 10845 7555
rect 10865 7535 10875 7555
rect 10835 7520 10875 7535
rect 10890 7605 10930 7620
rect 10890 7585 10900 7605
rect 10920 7585 10930 7605
rect 10890 7555 10930 7585
rect 10890 7535 10900 7555
rect 10920 7535 10930 7555
rect 10890 7520 10930 7535
rect 11220 7610 11230 7630
rect 11250 7610 11260 7630
rect 11220 7580 11260 7610
rect 11220 7560 11230 7580
rect 11250 7560 11260 7580
rect 11220 7530 11260 7560
rect 11220 7510 11230 7530
rect 11250 7510 11260 7530
rect 11220 7495 11260 7510
rect 11280 7880 11320 7895
rect 11280 7860 11290 7880
rect 11310 7860 11320 7880
rect 11280 7830 11320 7860
rect 11280 7810 11290 7830
rect 11310 7810 11320 7830
rect 11280 7780 11320 7810
rect 11280 7760 11290 7780
rect 11310 7760 11320 7780
rect 11280 7730 11320 7760
rect 11280 7710 11290 7730
rect 11310 7710 11320 7730
rect 11280 7680 11320 7710
rect 11280 7660 11290 7680
rect 11310 7660 11320 7680
rect 11280 7630 11320 7660
rect 11280 7610 11290 7630
rect 11310 7610 11320 7630
rect 11280 7580 11320 7610
rect 11280 7560 11290 7580
rect 11310 7560 11320 7580
rect 11280 7530 11320 7560
rect 11280 7510 11290 7530
rect 11310 7510 11320 7530
rect 11280 7495 11320 7510
rect 11340 7880 11380 7895
rect 11340 7860 11350 7880
rect 11370 7860 11380 7880
rect 11340 7830 11380 7860
rect 11340 7810 11350 7830
rect 11370 7810 11380 7830
rect 11340 7780 11380 7810
rect 11340 7760 11350 7780
rect 11370 7760 11380 7780
rect 11340 7730 11380 7760
rect 11340 7710 11350 7730
rect 11370 7710 11380 7730
rect 11340 7680 11380 7710
rect 11340 7660 11350 7680
rect 11370 7660 11380 7680
rect 11340 7630 11380 7660
rect 11340 7610 11350 7630
rect 11370 7610 11380 7630
rect 11340 7580 11380 7610
rect 11340 7560 11350 7580
rect 11370 7560 11380 7580
rect 11340 7530 11380 7560
rect 11340 7510 11350 7530
rect 11370 7510 11380 7530
rect 11340 7495 11380 7510
rect 11400 7880 11440 7895
rect 11400 7860 11410 7880
rect 11430 7860 11440 7880
rect 11400 7830 11440 7860
rect 11400 7810 11410 7830
rect 11430 7810 11440 7830
rect 11400 7780 11440 7810
rect 11400 7760 11410 7780
rect 11430 7760 11440 7780
rect 11400 7730 11440 7760
rect 11400 7710 11410 7730
rect 11430 7710 11440 7730
rect 11400 7680 11440 7710
rect 11400 7660 11410 7680
rect 11430 7660 11440 7680
rect 11400 7630 11440 7660
rect 11400 7610 11410 7630
rect 11430 7610 11440 7630
rect 11400 7580 11440 7610
rect 11400 7560 11410 7580
rect 11430 7560 11440 7580
rect 11400 7530 11440 7560
rect 11400 7510 11410 7530
rect 11430 7510 11440 7530
rect 11400 7495 11440 7510
rect 11460 7880 11500 7895
rect 11460 7860 11470 7880
rect 11490 7860 11500 7880
rect 11460 7830 11500 7860
rect 11460 7810 11470 7830
rect 11490 7810 11500 7830
rect 11460 7780 11500 7810
rect 11460 7760 11470 7780
rect 11490 7760 11500 7780
rect 11460 7730 11500 7760
rect 11460 7710 11470 7730
rect 11490 7710 11500 7730
rect 11460 7680 11500 7710
rect 11460 7660 11470 7680
rect 11490 7660 11500 7680
rect 11460 7630 11500 7660
rect 11460 7610 11470 7630
rect 11490 7610 11500 7630
rect 11460 7580 11500 7610
rect 11460 7560 11470 7580
rect 11490 7560 11500 7580
rect 11460 7530 11500 7560
rect 11460 7510 11470 7530
rect 11490 7510 11500 7530
rect 11460 7495 11500 7510
rect 11520 7880 11560 7895
rect 11520 7860 11530 7880
rect 11550 7860 11560 7880
rect 11520 7830 11560 7860
rect 11520 7810 11530 7830
rect 11550 7810 11560 7830
rect 11520 7780 11560 7810
rect 11520 7760 11530 7780
rect 11550 7760 11560 7780
rect 11520 7730 11560 7760
rect 11520 7710 11530 7730
rect 11550 7710 11560 7730
rect 11520 7680 11560 7710
rect 11520 7660 11530 7680
rect 11550 7660 11560 7680
rect 11520 7630 11560 7660
rect 11520 7610 11530 7630
rect 11550 7610 11560 7630
rect 11520 7580 11560 7610
rect 11520 7560 11530 7580
rect 11550 7560 11560 7580
rect 11520 7530 11560 7560
rect 11520 7510 11530 7530
rect 11550 7510 11560 7530
rect 11520 7495 11560 7510
rect 11580 7880 11620 7895
rect 11580 7860 11590 7880
rect 11610 7860 11620 7880
rect 11580 7830 11620 7860
rect 11580 7810 11590 7830
rect 11610 7810 11620 7830
rect 11580 7780 11620 7810
rect 11580 7760 11590 7780
rect 11610 7760 11620 7780
rect 11580 7730 11620 7760
rect 11580 7710 11590 7730
rect 11610 7710 11620 7730
rect 11580 7680 11620 7710
rect 11580 7660 11590 7680
rect 11610 7660 11620 7680
rect 11580 7630 11620 7660
rect 11580 7610 11590 7630
rect 11610 7610 11620 7630
rect 11580 7580 11620 7610
rect 11580 7560 11590 7580
rect 11610 7560 11620 7580
rect 11580 7530 11620 7560
rect 11580 7510 11590 7530
rect 11610 7510 11620 7530
rect 11580 7495 11620 7510
rect 11640 7880 11680 7895
rect 11640 7860 11650 7880
rect 11670 7860 11680 7880
rect 11640 7830 11680 7860
rect 11640 7810 11650 7830
rect 11670 7810 11680 7830
rect 11640 7780 11680 7810
rect 11640 7760 11650 7780
rect 11670 7760 11680 7780
rect 11640 7730 11680 7760
rect 11640 7710 11650 7730
rect 11670 7710 11680 7730
rect 11640 7680 11680 7710
rect 11640 7660 11650 7680
rect 11670 7660 11680 7680
rect 11640 7630 11680 7660
rect 11640 7610 11650 7630
rect 11670 7610 11680 7630
rect 11640 7580 11680 7610
rect 11640 7560 11650 7580
rect 11670 7560 11680 7580
rect 11640 7530 11680 7560
rect 11640 7510 11650 7530
rect 11670 7510 11680 7530
rect 11640 7495 11680 7510
rect 11700 7880 11740 7895
rect 11700 7860 11710 7880
rect 11730 7860 11740 7880
rect 11700 7830 11740 7860
rect 11700 7810 11710 7830
rect 11730 7810 11740 7830
rect 11700 7780 11740 7810
rect 11700 7760 11710 7780
rect 11730 7760 11740 7780
rect 11700 7730 11740 7760
rect 11700 7710 11710 7730
rect 11730 7710 11740 7730
rect 11700 7680 11740 7710
rect 11700 7660 11710 7680
rect 11730 7660 11740 7680
rect 11700 7630 11740 7660
rect 11700 7610 11710 7630
rect 11730 7610 11740 7630
rect 11700 7580 11740 7610
rect 11700 7560 11710 7580
rect 11730 7560 11740 7580
rect 11700 7530 11740 7560
rect 11700 7510 11710 7530
rect 11730 7510 11740 7530
rect 11700 7495 11740 7510
rect 11760 7880 11800 7895
rect 11760 7860 11770 7880
rect 11790 7860 11800 7880
rect 11760 7830 11800 7860
rect 11760 7810 11770 7830
rect 11790 7810 11800 7830
rect 11760 7780 11800 7810
rect 11760 7760 11770 7780
rect 11790 7760 11800 7780
rect 11760 7730 11800 7760
rect 11760 7710 11770 7730
rect 11790 7710 11800 7730
rect 11760 7680 11800 7710
rect 11760 7660 11770 7680
rect 11790 7660 11800 7680
rect 11760 7630 11800 7660
rect 11760 7610 11770 7630
rect 11790 7610 11800 7630
rect 11760 7580 11800 7610
rect 11760 7560 11770 7580
rect 11790 7560 11800 7580
rect 11760 7530 11800 7560
rect 11760 7510 11770 7530
rect 11790 7510 11800 7530
rect 11760 7495 11800 7510
rect 11820 7880 11860 7895
rect 11820 7860 11830 7880
rect 11850 7860 11860 7880
rect 11820 7830 11860 7860
rect 11820 7810 11830 7830
rect 11850 7810 11860 7830
rect 11820 7780 11860 7810
rect 11820 7760 11830 7780
rect 11850 7760 11860 7780
rect 11820 7730 11860 7760
rect 11820 7710 11830 7730
rect 11850 7710 11860 7730
rect 11820 7680 11860 7710
rect 11820 7660 11830 7680
rect 11850 7660 11860 7680
rect 11820 7630 11860 7660
rect 11820 7610 11830 7630
rect 11850 7610 11860 7630
rect 11820 7580 11860 7610
rect 11820 7560 11830 7580
rect 11850 7560 11860 7580
rect 11820 7530 11860 7560
rect 11820 7510 11830 7530
rect 11850 7510 11860 7530
rect 11820 7495 11860 7510
rect 11880 7880 11920 7895
rect 11880 7860 11890 7880
rect 11910 7860 11920 7880
rect 11880 7830 11920 7860
rect 11880 7810 11890 7830
rect 11910 7810 11920 7830
rect 11880 7780 11920 7810
rect 11880 7760 11890 7780
rect 11910 7760 11920 7780
rect 11880 7730 11920 7760
rect 11880 7710 11890 7730
rect 11910 7710 11920 7730
rect 11880 7680 11920 7710
rect 11880 7660 11890 7680
rect 11910 7660 11920 7680
rect 11880 7630 11920 7660
rect 11880 7610 11890 7630
rect 11910 7610 11920 7630
rect 11880 7580 11920 7610
rect 11880 7560 11890 7580
rect 11910 7560 11920 7580
rect 11880 7530 11920 7560
rect 11880 7510 11890 7530
rect 11910 7510 11920 7530
rect 11880 7495 11920 7510
rect 11940 7880 11980 7895
rect 11940 7860 11950 7880
rect 11970 7860 11980 7880
rect 11940 7830 11980 7860
rect 11940 7810 11950 7830
rect 11970 7810 11980 7830
rect 11940 7780 11980 7810
rect 11940 7760 11950 7780
rect 11970 7760 11980 7780
rect 11940 7730 11980 7760
rect 11940 7710 11950 7730
rect 11970 7710 11980 7730
rect 11940 7680 11980 7710
rect 11940 7660 11950 7680
rect 11970 7660 11980 7680
rect 11940 7630 11980 7660
rect 11940 7610 11950 7630
rect 11970 7610 11980 7630
rect 11940 7580 11980 7610
rect 11940 7560 11950 7580
rect 11970 7560 11980 7580
rect 11940 7530 11980 7560
rect 11940 7510 11950 7530
rect 11970 7510 11980 7530
rect 11940 7495 11980 7510
rect 12000 7880 12040 7895
rect 12000 7860 12010 7880
rect 12030 7860 12040 7880
rect 12000 7830 12040 7860
rect 12000 7810 12010 7830
rect 12030 7810 12040 7830
rect 12000 7780 12040 7810
rect 12000 7760 12010 7780
rect 12030 7760 12040 7780
rect 12000 7730 12040 7760
rect 12000 7710 12010 7730
rect 12030 7710 12040 7730
rect 12000 7680 12040 7710
rect 12000 7660 12010 7680
rect 12030 7660 12040 7680
rect 12000 7630 12040 7660
rect 12000 7610 12010 7630
rect 12030 7610 12040 7630
rect 12000 7580 12040 7610
rect 12000 7560 12010 7580
rect 12030 7560 12040 7580
rect 12000 7530 12040 7560
rect 12000 7510 12010 7530
rect 12030 7510 12040 7530
rect 12000 7495 12040 7510
rect 12060 7880 12100 7895
rect 12060 7860 12070 7880
rect 12090 7860 12100 7880
rect 12060 7830 12100 7860
rect 12060 7810 12070 7830
rect 12090 7810 12100 7830
rect 12060 7780 12100 7810
rect 12060 7760 12070 7780
rect 12090 7760 12100 7780
rect 12060 7730 12100 7760
rect 12060 7710 12070 7730
rect 12090 7710 12100 7730
rect 12060 7680 12100 7710
rect 12060 7660 12070 7680
rect 12090 7660 12100 7680
rect 12060 7630 12100 7660
rect 12060 7610 12070 7630
rect 12090 7610 12100 7630
rect 12060 7580 12100 7610
rect 12060 7560 12070 7580
rect 12090 7560 12100 7580
rect 12060 7530 12100 7560
rect 12060 7510 12070 7530
rect 12090 7510 12100 7530
rect 12060 7495 12100 7510
rect 12120 7880 12160 7895
rect 12120 7860 12130 7880
rect 12150 7860 12160 7880
rect 12120 7830 12160 7860
rect 12120 7810 12130 7830
rect 12150 7810 12160 7830
rect 12120 7780 12160 7810
rect 12120 7760 12130 7780
rect 12150 7760 12160 7780
rect 12120 7730 12160 7760
rect 12120 7710 12130 7730
rect 12150 7710 12160 7730
rect 12120 7680 12160 7710
rect 12120 7660 12130 7680
rect 12150 7660 12160 7680
rect 12120 7630 12160 7660
rect 12120 7610 12130 7630
rect 12150 7610 12160 7630
rect 12120 7580 12160 7610
rect 12120 7560 12130 7580
rect 12150 7560 12160 7580
rect 12120 7530 12160 7560
rect 12120 7510 12130 7530
rect 12150 7510 12160 7530
rect 12120 7495 12160 7510
rect 12180 7880 12220 7895
rect 12180 7860 12190 7880
rect 12210 7860 12220 7880
rect 12180 7830 12220 7860
rect 12180 7810 12190 7830
rect 12210 7810 12220 7830
rect 12180 7780 12220 7810
rect 12180 7760 12190 7780
rect 12210 7760 12220 7780
rect 12180 7730 12220 7760
rect 12180 7710 12190 7730
rect 12210 7710 12220 7730
rect 12180 7680 12220 7710
rect 12180 7660 12190 7680
rect 12210 7660 12220 7680
rect 12180 7630 12220 7660
rect 12180 7610 12190 7630
rect 12210 7610 12220 7630
rect 12180 7580 12220 7610
rect 12180 7560 12190 7580
rect 12210 7560 12220 7580
rect 12180 7530 12220 7560
rect 12180 7510 12190 7530
rect 12210 7510 12220 7530
rect 12180 7495 12220 7510
rect 12240 7880 12280 7895
rect 12240 7860 12250 7880
rect 12270 7860 12280 7880
rect 12240 7830 12280 7860
rect 12240 7810 12250 7830
rect 12270 7810 12280 7830
rect 12240 7780 12280 7810
rect 12240 7760 12250 7780
rect 12270 7760 12280 7780
rect 12240 7730 12280 7760
rect 12240 7710 12250 7730
rect 12270 7710 12280 7730
rect 12240 7680 12280 7710
rect 12240 7660 12250 7680
rect 12270 7660 12280 7680
rect 12240 7630 12280 7660
rect 12240 7610 12250 7630
rect 12270 7610 12280 7630
rect 12240 7580 12280 7610
rect 12240 7560 12250 7580
rect 12270 7560 12280 7580
rect 12240 7530 12280 7560
rect 12240 7510 12250 7530
rect 12270 7510 12280 7530
rect 12240 7495 12280 7510
rect 12300 7880 12340 7895
rect 12300 7860 12310 7880
rect 12330 7860 12340 7880
rect 12300 7830 12340 7860
rect 12300 7810 12310 7830
rect 12330 7810 12340 7830
rect 12300 7780 12340 7810
rect 12300 7760 12310 7780
rect 12330 7760 12340 7780
rect 12300 7730 12340 7760
rect 12300 7710 12310 7730
rect 12330 7710 12340 7730
rect 12300 7680 12340 7710
rect 12300 7660 12310 7680
rect 12330 7660 12340 7680
rect 12300 7630 12340 7660
rect 12300 7610 12310 7630
rect 12330 7610 12340 7630
rect 12300 7580 12340 7610
rect 12300 7560 12310 7580
rect 12330 7560 12340 7580
rect 12300 7530 12340 7560
rect 12300 7510 12310 7530
rect 12330 7510 12340 7530
rect 12300 7495 12340 7510
rect 12360 7880 12400 7895
rect 12360 7860 12370 7880
rect 12390 7860 12400 7880
rect 12360 7830 12400 7860
rect 12360 7810 12370 7830
rect 12390 7810 12400 7830
rect 12360 7780 12400 7810
rect 12360 7760 12370 7780
rect 12390 7760 12400 7780
rect 12360 7730 12400 7760
rect 12360 7710 12370 7730
rect 12390 7710 12400 7730
rect 12360 7680 12400 7710
rect 12360 7660 12370 7680
rect 12390 7660 12400 7680
rect 12360 7630 12400 7660
rect 12360 7610 12370 7630
rect 12390 7610 12400 7630
rect 12360 7580 12400 7610
rect 12360 7560 12370 7580
rect 12390 7560 12400 7580
rect 12360 7530 12400 7560
rect 12360 7510 12370 7530
rect 12390 7510 12400 7530
rect 12360 7495 12400 7510
rect 12420 7880 12460 7895
rect 12420 7860 12430 7880
rect 12450 7860 12460 7880
rect 12420 7830 12460 7860
rect 12420 7810 12430 7830
rect 12450 7810 12460 7830
rect 12420 7780 12460 7810
rect 12420 7760 12430 7780
rect 12450 7760 12460 7780
rect 12420 7730 12460 7760
rect 12420 7710 12430 7730
rect 12450 7710 12460 7730
rect 12420 7680 12460 7710
rect 12420 7660 12430 7680
rect 12450 7660 12460 7680
rect 12420 7630 12460 7660
rect 12420 7610 12430 7630
rect 12450 7610 12460 7630
rect 12420 7580 12460 7610
rect 12420 7560 12430 7580
rect 12450 7560 12460 7580
rect 12420 7530 12460 7560
rect 12420 7510 12430 7530
rect 12450 7510 12460 7530
rect 12420 7495 12460 7510
rect 12480 7880 12520 7895
rect 12480 7860 12490 7880
rect 12510 7860 12520 7880
rect 12480 7830 12520 7860
rect 12480 7810 12490 7830
rect 12510 7810 12520 7830
rect 12480 7780 12520 7810
rect 12480 7760 12490 7780
rect 12510 7760 12520 7780
rect 12480 7730 12520 7760
rect 12480 7710 12490 7730
rect 12510 7710 12520 7730
rect 12480 7680 12520 7710
rect 12480 7660 12490 7680
rect 12510 7660 12520 7680
rect 12480 7630 12520 7660
rect 12480 7610 12490 7630
rect 12510 7610 12520 7630
rect 12480 7580 12520 7610
rect 12480 7560 12490 7580
rect 12510 7560 12520 7580
rect 12480 7530 12520 7560
rect 12480 7510 12490 7530
rect 12510 7510 12520 7530
rect 12480 7495 12520 7510
rect 12540 7880 12580 7895
rect 20390 7940 20430 7955
rect 20445 8225 20485 8240
rect 20445 8205 20455 8225
rect 20475 8205 20485 8225
rect 20445 8175 20485 8205
rect 20445 8155 20455 8175
rect 20475 8155 20485 8175
rect 20445 8125 20485 8155
rect 20445 8105 20455 8125
rect 20475 8105 20485 8125
rect 20445 8075 20485 8105
rect 20445 8055 20455 8075
rect 20475 8055 20485 8075
rect 20445 8025 20485 8055
rect 20445 8005 20455 8025
rect 20475 8005 20485 8025
rect 20445 7975 20485 8005
rect 20445 7955 20455 7975
rect 20475 7955 20485 7975
rect 20445 7940 20485 7955
rect 20500 8225 20540 8240
rect 20500 8205 20510 8225
rect 20530 8205 20540 8225
rect 20500 8175 20540 8205
rect 20500 8155 20510 8175
rect 20530 8155 20540 8175
rect 20500 8125 20540 8155
rect 20500 8105 20510 8125
rect 20530 8105 20540 8125
rect 20500 8075 20540 8105
rect 20500 8055 20510 8075
rect 20530 8055 20540 8075
rect 20500 8025 20540 8055
rect 20500 8005 20510 8025
rect 20530 8005 20540 8025
rect 20500 7975 20540 8005
rect 20500 7955 20510 7975
rect 20530 7955 20540 7975
rect 20500 7940 20540 7955
rect 20555 8225 20595 8240
rect 20555 8205 20565 8225
rect 20585 8205 20595 8225
rect 20555 8175 20595 8205
rect 20555 8155 20565 8175
rect 20585 8155 20595 8175
rect 20555 8125 20595 8155
rect 20555 8105 20565 8125
rect 20585 8105 20595 8125
rect 20555 8075 20595 8105
rect 20555 8055 20565 8075
rect 20585 8055 20595 8075
rect 20555 8025 20595 8055
rect 20555 8005 20565 8025
rect 20585 8005 20595 8025
rect 20555 7975 20595 8005
rect 20555 7955 20565 7975
rect 20585 7955 20595 7975
rect 20555 7940 20595 7955
rect 20610 8225 20650 8240
rect 20610 8205 20620 8225
rect 20640 8205 20650 8225
rect 20610 8175 20650 8205
rect 20610 8155 20620 8175
rect 20640 8155 20650 8175
rect 20610 8125 20650 8155
rect 20610 8105 20620 8125
rect 20640 8105 20650 8125
rect 20610 8075 20650 8105
rect 20610 8055 20620 8075
rect 20640 8055 20650 8075
rect 20610 8025 20650 8055
rect 20610 8005 20620 8025
rect 20640 8005 20650 8025
rect 20610 7975 20650 8005
rect 20610 7955 20620 7975
rect 20640 7955 20650 7975
rect 20610 7940 20650 7955
rect 20665 8225 20705 8240
rect 20665 8205 20675 8225
rect 20695 8205 20705 8225
rect 20665 8175 20705 8205
rect 20665 8155 20675 8175
rect 20695 8155 20705 8175
rect 20665 8125 20705 8155
rect 20665 8105 20675 8125
rect 20695 8105 20705 8125
rect 20665 8075 20705 8105
rect 20665 8055 20675 8075
rect 20695 8055 20705 8075
rect 20665 8025 20705 8055
rect 20665 8005 20675 8025
rect 20695 8005 20705 8025
rect 20665 7975 20705 8005
rect 20665 7955 20675 7975
rect 20695 7955 20705 7975
rect 20665 7940 20705 7955
rect 20720 8225 20760 8240
rect 20720 8205 20730 8225
rect 20750 8205 20760 8225
rect 20720 8175 20760 8205
rect 20720 8155 20730 8175
rect 20750 8155 20760 8175
rect 20720 8125 20760 8155
rect 20720 8105 20730 8125
rect 20750 8105 20760 8125
rect 20720 8075 20760 8105
rect 20720 8055 20730 8075
rect 20750 8055 20760 8075
rect 20720 8025 20760 8055
rect 20720 8005 20730 8025
rect 20750 8005 20760 8025
rect 20720 7975 20760 8005
rect 20720 7955 20730 7975
rect 20750 7955 20760 7975
rect 20720 7940 20760 7955
rect 20775 8225 20815 8240
rect 20775 8205 20785 8225
rect 20805 8205 20815 8225
rect 20775 8175 20815 8205
rect 20775 8155 20785 8175
rect 20805 8155 20815 8175
rect 20775 8125 20815 8155
rect 20775 8105 20785 8125
rect 20805 8105 20815 8125
rect 20775 8075 20815 8105
rect 20775 8055 20785 8075
rect 20805 8055 20815 8075
rect 20775 8025 20815 8055
rect 20775 8005 20785 8025
rect 20805 8005 20815 8025
rect 20775 7975 20815 8005
rect 20775 7955 20785 7975
rect 20805 7955 20815 7975
rect 20775 7940 20815 7955
rect 20830 8225 20870 8240
rect 20830 8205 20840 8225
rect 20860 8205 20870 8225
rect 20830 8175 20870 8205
rect 20830 8155 20840 8175
rect 20860 8155 20870 8175
rect 20830 8125 20870 8155
rect 20830 8105 20840 8125
rect 20860 8105 20870 8125
rect 20830 8075 20870 8105
rect 20830 8055 20840 8075
rect 20860 8055 20870 8075
rect 20830 8025 20870 8055
rect 20830 8005 20840 8025
rect 20860 8005 20870 8025
rect 20830 7975 20870 8005
rect 20830 7955 20840 7975
rect 20860 7955 20870 7975
rect 20830 7940 20870 7955
rect 20885 8225 20925 8240
rect 20885 8205 20895 8225
rect 20915 8205 20925 8225
rect 20885 8175 20925 8205
rect 20885 8155 20895 8175
rect 20915 8155 20925 8175
rect 20885 8125 20925 8155
rect 20885 8105 20895 8125
rect 20915 8105 20925 8125
rect 20885 8075 20925 8105
rect 20885 8055 20895 8075
rect 20915 8055 20925 8075
rect 20885 8025 20925 8055
rect 20885 8005 20895 8025
rect 20915 8005 20925 8025
rect 20885 7975 20925 8005
rect 20885 7955 20895 7975
rect 20915 7955 20925 7975
rect 20885 7940 20925 7955
rect 20940 8225 20980 8240
rect 20940 8205 20950 8225
rect 20970 8205 20980 8225
rect 20940 8175 20980 8205
rect 20940 8155 20950 8175
rect 20970 8155 20980 8175
rect 20940 8125 20980 8155
rect 20940 8105 20950 8125
rect 20970 8105 20980 8125
rect 20940 8075 20980 8105
rect 20940 8055 20950 8075
rect 20970 8055 20980 8075
rect 20940 8025 20980 8055
rect 20940 8005 20950 8025
rect 20970 8005 20980 8025
rect 20940 7975 20980 8005
rect 20940 7955 20950 7975
rect 20970 7955 20980 7975
rect 20940 7940 20980 7955
rect 20995 8225 21035 8240
rect 20995 8205 21005 8225
rect 21025 8205 21035 8225
rect 20995 8175 21035 8205
rect 20995 8155 21005 8175
rect 21025 8155 21035 8175
rect 20995 8125 21035 8155
rect 20995 8105 21005 8125
rect 21025 8105 21035 8125
rect 20995 8075 21035 8105
rect 20995 8055 21005 8075
rect 21025 8055 21035 8075
rect 20995 8025 21035 8055
rect 20995 8005 21005 8025
rect 21025 8005 21035 8025
rect 20995 7975 21035 8005
rect 20995 7955 21005 7975
rect 21025 7955 21035 7975
rect 20995 7940 21035 7955
rect 21050 8225 21090 8240
rect 21050 8205 21060 8225
rect 21080 8205 21090 8225
rect 21050 8175 21090 8205
rect 21050 8155 21060 8175
rect 21080 8155 21090 8175
rect 21050 8125 21090 8155
rect 21050 8105 21060 8125
rect 21080 8105 21090 8125
rect 21050 8075 21090 8105
rect 21050 8055 21060 8075
rect 21080 8055 21090 8075
rect 21050 8025 21090 8055
rect 21050 8005 21060 8025
rect 21080 8005 21090 8025
rect 21050 7975 21090 8005
rect 21050 7955 21060 7975
rect 21080 7955 21090 7975
rect 21050 7940 21090 7955
rect 21105 8225 21145 8240
rect 21105 8205 21115 8225
rect 21135 8205 21145 8225
rect 21105 8175 21145 8205
rect 21105 8155 21115 8175
rect 21135 8155 21145 8175
rect 21105 8125 21145 8155
rect 21105 8105 21115 8125
rect 21135 8105 21145 8125
rect 21105 8075 21145 8105
rect 21105 8055 21115 8075
rect 21135 8055 21145 8075
rect 21105 8025 21145 8055
rect 21105 8005 21115 8025
rect 21135 8005 21145 8025
rect 21105 7975 21145 8005
rect 21105 7955 21115 7975
rect 21135 7955 21145 7975
rect 21105 7940 21145 7955
rect 21160 8225 21200 8240
rect 21160 8205 21170 8225
rect 21190 8205 21200 8225
rect 21160 8175 21200 8205
rect 21160 8155 21170 8175
rect 21190 8155 21200 8175
rect 21160 8125 21200 8155
rect 21160 8105 21170 8125
rect 21190 8105 21200 8125
rect 21160 8075 21200 8105
rect 21160 8055 21170 8075
rect 21190 8055 21200 8075
rect 21160 8025 21200 8055
rect 21160 8005 21170 8025
rect 21190 8005 21200 8025
rect 21160 7975 21200 8005
rect 21160 7955 21170 7975
rect 21190 7955 21200 7975
rect 21160 7940 21200 7955
rect 21215 8225 21255 8240
rect 21215 8205 21225 8225
rect 21245 8205 21255 8225
rect 21215 8175 21255 8205
rect 21215 8155 21225 8175
rect 21245 8155 21255 8175
rect 21215 8125 21255 8155
rect 21215 8105 21225 8125
rect 21245 8105 21255 8125
rect 21215 8075 21255 8105
rect 21215 8055 21225 8075
rect 21245 8055 21255 8075
rect 21215 8025 21255 8055
rect 21215 8005 21225 8025
rect 21245 8005 21255 8025
rect 21215 7975 21255 8005
rect 21215 7955 21225 7975
rect 21245 7955 21255 7975
rect 21215 7940 21255 7955
rect 21270 8225 21310 8240
rect 21270 8205 21280 8225
rect 21300 8205 21310 8225
rect 21270 8175 21310 8205
rect 21270 8155 21280 8175
rect 21300 8155 21310 8175
rect 21270 8125 21310 8155
rect 21270 8105 21280 8125
rect 21300 8105 21310 8125
rect 21270 8075 21310 8105
rect 21270 8055 21280 8075
rect 21300 8055 21310 8075
rect 21270 8025 21310 8055
rect 21270 8005 21280 8025
rect 21300 8005 21310 8025
rect 21270 7975 21310 8005
rect 21270 7955 21280 7975
rect 21300 7955 21310 7975
rect 21270 7940 21310 7955
rect 21325 8225 21365 8240
rect 21325 8205 21335 8225
rect 21355 8205 21365 8225
rect 21325 8175 21365 8205
rect 21325 8155 21335 8175
rect 21355 8155 21365 8175
rect 21325 8125 21365 8155
rect 21325 8105 21335 8125
rect 21355 8105 21365 8125
rect 21325 8075 21365 8105
rect 21325 8055 21335 8075
rect 21355 8055 21365 8075
rect 21325 8025 21365 8055
rect 21325 8005 21335 8025
rect 21355 8005 21365 8025
rect 21325 7975 21365 8005
rect 21325 7955 21335 7975
rect 21355 7955 21365 7975
rect 21325 7940 21365 7955
rect 21380 8225 21420 8240
rect 21380 8205 21390 8225
rect 21410 8205 21420 8225
rect 21380 8175 21420 8205
rect 21380 8155 21390 8175
rect 21410 8155 21420 8175
rect 21380 8125 21420 8155
rect 21380 8105 21390 8125
rect 21410 8105 21420 8125
rect 21380 8075 21420 8105
rect 21380 8055 21390 8075
rect 21410 8055 21420 8075
rect 21380 8025 21420 8055
rect 21380 8005 21390 8025
rect 21410 8005 21420 8025
rect 21380 7975 21420 8005
rect 21380 7955 21390 7975
rect 21410 7955 21420 7975
rect 21380 7940 21420 7955
rect 21435 8225 21475 8240
rect 21435 8205 21445 8225
rect 21465 8205 21475 8225
rect 21435 8175 21475 8205
rect 21435 8155 21445 8175
rect 21465 8155 21475 8175
rect 21435 8125 21475 8155
rect 21435 8105 21445 8125
rect 21465 8105 21475 8125
rect 21435 8075 21475 8105
rect 21435 8055 21445 8075
rect 21465 8055 21475 8075
rect 21435 8025 21475 8055
rect 21435 8005 21445 8025
rect 21465 8005 21475 8025
rect 21435 7975 21475 8005
rect 21435 7955 21445 7975
rect 21465 7955 21475 7975
rect 21435 7940 21475 7955
rect 21490 8225 21530 8240
rect 21490 8205 21500 8225
rect 21520 8205 21530 8225
rect 21490 8175 21530 8205
rect 21490 8155 21500 8175
rect 21520 8155 21530 8175
rect 21490 8125 21530 8155
rect 21490 8105 21500 8125
rect 21520 8105 21530 8125
rect 21490 8075 21530 8105
rect 21490 8055 21500 8075
rect 21520 8055 21530 8075
rect 21490 8025 21530 8055
rect 21490 8005 21500 8025
rect 21520 8005 21530 8025
rect 21490 7975 21530 8005
rect 21490 7955 21500 7975
rect 21520 7955 21530 7975
rect 21490 7940 21530 7955
rect 21545 8225 21585 8240
rect 21545 8205 21555 8225
rect 21575 8205 21585 8225
rect 21545 8175 21585 8205
rect 21545 8155 21555 8175
rect 21575 8155 21585 8175
rect 21545 8125 21585 8155
rect 21545 8105 21555 8125
rect 21575 8105 21585 8125
rect 21545 8075 21585 8105
rect 21545 8055 21555 8075
rect 21575 8055 21585 8075
rect 21545 8025 21585 8055
rect 21545 8005 21555 8025
rect 21575 8005 21585 8025
rect 21545 7975 21585 8005
rect 21545 7955 21555 7975
rect 21575 7955 21585 7975
rect 21545 7940 21585 7955
rect 21600 8225 21640 8240
rect 21600 8205 21610 8225
rect 21630 8205 21640 8225
rect 21600 8175 21640 8205
rect 21600 8155 21610 8175
rect 21630 8155 21640 8175
rect 21600 8125 21640 8155
rect 21600 8105 21610 8125
rect 21630 8105 21640 8125
rect 21600 8075 21640 8105
rect 21600 8055 21610 8075
rect 21630 8055 21640 8075
rect 21600 8025 21640 8055
rect 21600 8005 21610 8025
rect 21630 8005 21640 8025
rect 21600 7975 21640 8005
rect 21600 7955 21610 7975
rect 21630 7955 21640 7975
rect 21600 7940 21640 7955
rect 12540 7860 12550 7880
rect 12570 7860 12580 7880
rect 12540 7830 12580 7860
rect 18720 7880 18760 7895
rect 18720 7860 18730 7880
rect 18750 7860 18760 7880
rect 12540 7810 12550 7830
rect 12570 7810 12580 7830
rect 12540 7780 12580 7810
rect 12540 7760 12550 7780
rect 12570 7760 12580 7780
rect 12540 7730 12580 7760
rect 12540 7710 12550 7730
rect 12570 7710 12580 7730
rect 12540 7680 12580 7710
rect 18720 7830 18760 7860
rect 18720 7810 18730 7830
rect 18750 7810 18760 7830
rect 18720 7780 18760 7810
rect 18720 7760 18730 7780
rect 18750 7760 18760 7780
rect 18720 7730 18760 7760
rect 18720 7710 18730 7730
rect 18750 7710 18760 7730
rect 12540 7660 12550 7680
rect 12570 7660 12580 7680
rect 12540 7630 12580 7660
rect 18720 7680 18760 7710
rect 18720 7660 18730 7680
rect 18750 7660 18760 7680
rect 12540 7610 12550 7630
rect 12570 7610 12580 7630
rect 18720 7630 18760 7660
rect 12540 7580 12580 7610
rect 12540 7560 12550 7580
rect 12570 7560 12580 7580
rect 12540 7530 12580 7560
rect 12540 7510 12550 7530
rect 12570 7510 12580 7530
rect 12895 7605 12935 7620
rect 12895 7585 12905 7605
rect 12925 7585 12935 7605
rect 12895 7555 12935 7585
rect 12895 7535 12905 7555
rect 12925 7535 12935 7555
rect 12895 7520 12935 7535
rect 12950 7605 12990 7620
rect 12950 7585 12960 7605
rect 12980 7585 12990 7605
rect 12950 7555 12990 7585
rect 12950 7535 12960 7555
rect 12980 7535 12990 7555
rect 12950 7520 12990 7535
rect 13005 7605 13045 7620
rect 13005 7585 13015 7605
rect 13035 7585 13045 7605
rect 13005 7555 13045 7585
rect 13005 7535 13015 7555
rect 13035 7535 13045 7555
rect 13005 7520 13045 7535
rect 13060 7605 13100 7620
rect 13060 7585 13070 7605
rect 13090 7585 13100 7605
rect 13060 7555 13100 7585
rect 13060 7535 13070 7555
rect 13090 7535 13100 7555
rect 13060 7520 13100 7535
rect 13115 7605 13155 7620
rect 13115 7585 13125 7605
rect 13145 7585 13155 7605
rect 13115 7555 13155 7585
rect 13115 7535 13125 7555
rect 13145 7535 13155 7555
rect 13115 7520 13155 7535
rect 13170 7605 13210 7620
rect 13170 7585 13180 7605
rect 13200 7585 13210 7605
rect 13170 7555 13210 7585
rect 13170 7535 13180 7555
rect 13200 7535 13210 7555
rect 13170 7520 13210 7535
rect 13225 7605 13265 7620
rect 13225 7585 13235 7605
rect 13255 7585 13265 7605
rect 13225 7555 13265 7585
rect 13225 7535 13235 7555
rect 13255 7535 13265 7555
rect 13225 7520 13265 7535
rect 13280 7605 13320 7620
rect 13280 7585 13290 7605
rect 13310 7585 13320 7605
rect 13280 7555 13320 7585
rect 13280 7535 13290 7555
rect 13310 7535 13320 7555
rect 13280 7520 13320 7535
rect 13335 7605 13375 7620
rect 13335 7585 13345 7605
rect 13365 7585 13375 7605
rect 13335 7555 13375 7585
rect 13335 7535 13345 7555
rect 13365 7535 13375 7555
rect 13335 7520 13375 7535
rect 13390 7605 13430 7620
rect 13390 7585 13400 7605
rect 13420 7585 13430 7605
rect 13390 7555 13430 7585
rect 13390 7535 13400 7555
rect 13420 7535 13430 7555
rect 13390 7520 13430 7535
rect 13445 7605 13485 7620
rect 13445 7585 13455 7605
rect 13475 7585 13485 7605
rect 13445 7555 13485 7585
rect 13445 7535 13455 7555
rect 13475 7535 13485 7555
rect 13445 7520 13485 7535
rect 13500 7605 13540 7620
rect 13500 7585 13510 7605
rect 13530 7585 13540 7605
rect 13500 7555 13540 7585
rect 13500 7535 13510 7555
rect 13530 7535 13540 7555
rect 13500 7520 13540 7535
rect 13555 7605 13595 7620
rect 13555 7585 13565 7605
rect 13585 7585 13595 7605
rect 13555 7555 13595 7585
rect 13555 7535 13565 7555
rect 13585 7535 13595 7555
rect 13555 7520 13595 7535
rect 13610 7605 13650 7620
rect 13610 7585 13620 7605
rect 13640 7585 13650 7605
rect 13610 7555 13650 7585
rect 13610 7535 13620 7555
rect 13640 7535 13650 7555
rect 13610 7520 13650 7535
rect 13665 7605 13705 7620
rect 13665 7585 13675 7605
rect 13695 7585 13705 7605
rect 13665 7555 13705 7585
rect 13665 7535 13675 7555
rect 13695 7535 13705 7555
rect 13665 7520 13705 7535
rect 13720 7605 13760 7620
rect 13720 7585 13730 7605
rect 13750 7585 13760 7605
rect 13720 7555 13760 7585
rect 13720 7535 13730 7555
rect 13750 7535 13760 7555
rect 13720 7520 13760 7535
rect 13775 7605 13815 7620
rect 13775 7585 13785 7605
rect 13805 7585 13815 7605
rect 13775 7555 13815 7585
rect 13775 7535 13785 7555
rect 13805 7535 13815 7555
rect 13775 7520 13815 7535
rect 13830 7605 13870 7620
rect 13830 7585 13840 7605
rect 13860 7585 13870 7605
rect 13830 7555 13870 7585
rect 13830 7535 13840 7555
rect 13860 7535 13870 7555
rect 13830 7520 13870 7535
rect 13885 7605 13925 7620
rect 13885 7585 13895 7605
rect 13915 7585 13925 7605
rect 13885 7555 13925 7585
rect 13885 7535 13895 7555
rect 13915 7535 13925 7555
rect 13885 7520 13925 7535
rect 13940 7605 13980 7620
rect 13940 7585 13950 7605
rect 13970 7585 13980 7605
rect 13940 7555 13980 7585
rect 13940 7535 13950 7555
rect 13970 7535 13980 7555
rect 13940 7520 13980 7535
rect 13995 7605 14035 7620
rect 13995 7585 14005 7605
rect 14025 7585 14035 7605
rect 13995 7555 14035 7585
rect 13995 7535 14005 7555
rect 14025 7535 14035 7555
rect 13995 7520 14035 7535
rect 14050 7605 14090 7620
rect 14050 7585 14060 7605
rect 14080 7585 14090 7605
rect 14050 7555 14090 7585
rect 14050 7535 14060 7555
rect 14080 7535 14090 7555
rect 14050 7520 14090 7535
rect 14105 7605 14145 7620
rect 14105 7585 14115 7605
rect 14135 7585 14145 7605
rect 14105 7555 14145 7585
rect 14105 7535 14115 7555
rect 14135 7535 14145 7555
rect 14105 7520 14145 7535
rect 17180 7605 17220 7620
rect 17180 7585 17190 7605
rect 17210 7585 17220 7605
rect 17180 7555 17220 7585
rect 17180 7535 17190 7555
rect 17210 7535 17220 7555
rect 17180 7520 17220 7535
rect 17235 7605 17275 7620
rect 17235 7585 17245 7605
rect 17265 7585 17275 7605
rect 17235 7555 17275 7585
rect 17235 7535 17245 7555
rect 17265 7535 17275 7555
rect 17235 7520 17275 7535
rect 17290 7605 17330 7620
rect 17290 7585 17300 7605
rect 17320 7585 17330 7605
rect 17290 7555 17330 7585
rect 17290 7535 17300 7555
rect 17320 7535 17330 7555
rect 17290 7520 17330 7535
rect 17345 7605 17385 7620
rect 17345 7585 17355 7605
rect 17375 7585 17385 7605
rect 17345 7555 17385 7585
rect 17345 7535 17355 7555
rect 17375 7535 17385 7555
rect 17345 7520 17385 7535
rect 17400 7605 17440 7620
rect 17400 7585 17410 7605
rect 17430 7585 17440 7605
rect 17400 7555 17440 7585
rect 17400 7535 17410 7555
rect 17430 7535 17440 7555
rect 17400 7520 17440 7535
rect 17455 7605 17495 7620
rect 17455 7585 17465 7605
rect 17485 7585 17495 7605
rect 17455 7555 17495 7585
rect 17455 7535 17465 7555
rect 17485 7535 17495 7555
rect 17455 7520 17495 7535
rect 17510 7605 17550 7620
rect 17510 7585 17520 7605
rect 17540 7585 17550 7605
rect 17510 7555 17550 7585
rect 17510 7535 17520 7555
rect 17540 7535 17550 7555
rect 17510 7520 17550 7535
rect 17565 7605 17605 7620
rect 17565 7585 17575 7605
rect 17595 7585 17605 7605
rect 17565 7555 17605 7585
rect 17565 7535 17575 7555
rect 17595 7535 17605 7555
rect 17565 7520 17605 7535
rect 17620 7605 17660 7620
rect 17620 7585 17630 7605
rect 17650 7585 17660 7605
rect 17620 7555 17660 7585
rect 17620 7535 17630 7555
rect 17650 7535 17660 7555
rect 17620 7520 17660 7535
rect 17675 7605 17715 7620
rect 17675 7585 17685 7605
rect 17705 7585 17715 7605
rect 17675 7555 17715 7585
rect 17675 7535 17685 7555
rect 17705 7535 17715 7555
rect 17675 7520 17715 7535
rect 17730 7605 17770 7620
rect 17730 7585 17740 7605
rect 17760 7585 17770 7605
rect 17730 7555 17770 7585
rect 17730 7535 17740 7555
rect 17760 7535 17770 7555
rect 17730 7520 17770 7535
rect 17785 7605 17825 7620
rect 17785 7585 17795 7605
rect 17815 7585 17825 7605
rect 17785 7555 17825 7585
rect 17785 7535 17795 7555
rect 17815 7535 17825 7555
rect 17785 7520 17825 7535
rect 17840 7605 17880 7620
rect 17840 7585 17850 7605
rect 17870 7585 17880 7605
rect 17840 7555 17880 7585
rect 17840 7535 17850 7555
rect 17870 7535 17880 7555
rect 17840 7520 17880 7535
rect 17895 7605 17935 7620
rect 17895 7585 17905 7605
rect 17925 7585 17935 7605
rect 17895 7555 17935 7585
rect 17895 7535 17905 7555
rect 17925 7535 17935 7555
rect 17895 7520 17935 7535
rect 17950 7605 17990 7620
rect 17950 7585 17960 7605
rect 17980 7585 17990 7605
rect 17950 7555 17990 7585
rect 17950 7535 17960 7555
rect 17980 7535 17990 7555
rect 17950 7520 17990 7535
rect 18005 7605 18045 7620
rect 18005 7585 18015 7605
rect 18035 7585 18045 7605
rect 18005 7555 18045 7585
rect 18005 7535 18015 7555
rect 18035 7535 18045 7555
rect 18005 7520 18045 7535
rect 18060 7605 18100 7620
rect 18060 7585 18070 7605
rect 18090 7585 18100 7605
rect 18060 7555 18100 7585
rect 18060 7535 18070 7555
rect 18090 7535 18100 7555
rect 18060 7520 18100 7535
rect 18115 7605 18155 7620
rect 18115 7585 18125 7605
rect 18145 7585 18155 7605
rect 18115 7555 18155 7585
rect 18115 7535 18125 7555
rect 18145 7535 18155 7555
rect 18115 7520 18155 7535
rect 18170 7605 18210 7620
rect 18170 7585 18180 7605
rect 18200 7585 18210 7605
rect 18170 7555 18210 7585
rect 18170 7535 18180 7555
rect 18200 7535 18210 7555
rect 18170 7520 18210 7535
rect 18225 7605 18265 7620
rect 18225 7585 18235 7605
rect 18255 7585 18265 7605
rect 18225 7555 18265 7585
rect 18225 7535 18235 7555
rect 18255 7535 18265 7555
rect 18225 7520 18265 7535
rect 18280 7605 18320 7620
rect 18280 7585 18290 7605
rect 18310 7585 18320 7605
rect 18280 7555 18320 7585
rect 18280 7535 18290 7555
rect 18310 7535 18320 7555
rect 18280 7520 18320 7535
rect 18335 7605 18375 7620
rect 18335 7585 18345 7605
rect 18365 7585 18375 7605
rect 18335 7555 18375 7585
rect 18335 7535 18345 7555
rect 18365 7535 18375 7555
rect 18335 7520 18375 7535
rect 18390 7605 18430 7620
rect 18390 7585 18400 7605
rect 18420 7585 18430 7605
rect 18390 7555 18430 7585
rect 18390 7535 18400 7555
rect 18420 7535 18430 7555
rect 18390 7520 18430 7535
rect 18720 7610 18730 7630
rect 18750 7610 18760 7630
rect 18720 7580 18760 7610
rect 18720 7560 18730 7580
rect 18750 7560 18760 7580
rect 18720 7530 18760 7560
rect 12540 7495 12580 7510
rect 18720 7510 18730 7530
rect 18750 7510 18760 7530
rect 18720 7495 18760 7510
rect 18780 7880 18820 7895
rect 18780 7860 18790 7880
rect 18810 7860 18820 7880
rect 18780 7830 18820 7860
rect 18780 7810 18790 7830
rect 18810 7810 18820 7830
rect 18780 7780 18820 7810
rect 18780 7760 18790 7780
rect 18810 7760 18820 7780
rect 18780 7730 18820 7760
rect 18780 7710 18790 7730
rect 18810 7710 18820 7730
rect 18780 7680 18820 7710
rect 18780 7660 18790 7680
rect 18810 7660 18820 7680
rect 18780 7630 18820 7660
rect 18780 7610 18790 7630
rect 18810 7610 18820 7630
rect 18780 7580 18820 7610
rect 18780 7560 18790 7580
rect 18810 7560 18820 7580
rect 18780 7530 18820 7560
rect 18780 7510 18790 7530
rect 18810 7510 18820 7530
rect 18780 7495 18820 7510
rect 18840 7880 18880 7895
rect 18840 7860 18850 7880
rect 18870 7860 18880 7880
rect 18840 7830 18880 7860
rect 18840 7810 18850 7830
rect 18870 7810 18880 7830
rect 18840 7780 18880 7810
rect 18840 7760 18850 7780
rect 18870 7760 18880 7780
rect 18840 7730 18880 7760
rect 18840 7710 18850 7730
rect 18870 7710 18880 7730
rect 18840 7680 18880 7710
rect 18840 7660 18850 7680
rect 18870 7660 18880 7680
rect 18840 7630 18880 7660
rect 18840 7610 18850 7630
rect 18870 7610 18880 7630
rect 18840 7580 18880 7610
rect 18840 7560 18850 7580
rect 18870 7560 18880 7580
rect 18840 7530 18880 7560
rect 18840 7510 18850 7530
rect 18870 7510 18880 7530
rect 18840 7495 18880 7510
rect 18900 7880 18940 7895
rect 18900 7860 18910 7880
rect 18930 7860 18940 7880
rect 18900 7830 18940 7860
rect 18900 7810 18910 7830
rect 18930 7810 18940 7830
rect 18900 7780 18940 7810
rect 18900 7760 18910 7780
rect 18930 7760 18940 7780
rect 18900 7730 18940 7760
rect 18900 7710 18910 7730
rect 18930 7710 18940 7730
rect 18900 7680 18940 7710
rect 18900 7660 18910 7680
rect 18930 7660 18940 7680
rect 18900 7630 18940 7660
rect 18900 7610 18910 7630
rect 18930 7610 18940 7630
rect 18900 7580 18940 7610
rect 18900 7560 18910 7580
rect 18930 7560 18940 7580
rect 18900 7530 18940 7560
rect 18900 7510 18910 7530
rect 18930 7510 18940 7530
rect 18900 7495 18940 7510
rect 18960 7880 19000 7895
rect 18960 7860 18970 7880
rect 18990 7860 19000 7880
rect 18960 7830 19000 7860
rect 18960 7810 18970 7830
rect 18990 7810 19000 7830
rect 18960 7780 19000 7810
rect 18960 7760 18970 7780
rect 18990 7760 19000 7780
rect 18960 7730 19000 7760
rect 18960 7710 18970 7730
rect 18990 7710 19000 7730
rect 18960 7680 19000 7710
rect 18960 7660 18970 7680
rect 18990 7660 19000 7680
rect 18960 7630 19000 7660
rect 18960 7610 18970 7630
rect 18990 7610 19000 7630
rect 18960 7580 19000 7610
rect 18960 7560 18970 7580
rect 18990 7560 19000 7580
rect 18960 7530 19000 7560
rect 18960 7510 18970 7530
rect 18990 7510 19000 7530
rect 18960 7495 19000 7510
rect 19020 7880 19060 7895
rect 19020 7860 19030 7880
rect 19050 7860 19060 7880
rect 19020 7830 19060 7860
rect 19020 7810 19030 7830
rect 19050 7810 19060 7830
rect 19020 7780 19060 7810
rect 19020 7760 19030 7780
rect 19050 7760 19060 7780
rect 19020 7730 19060 7760
rect 19020 7710 19030 7730
rect 19050 7710 19060 7730
rect 19020 7680 19060 7710
rect 19020 7660 19030 7680
rect 19050 7660 19060 7680
rect 19020 7630 19060 7660
rect 19020 7610 19030 7630
rect 19050 7610 19060 7630
rect 19020 7580 19060 7610
rect 19020 7560 19030 7580
rect 19050 7560 19060 7580
rect 19020 7530 19060 7560
rect 19020 7510 19030 7530
rect 19050 7510 19060 7530
rect 19020 7495 19060 7510
rect 19080 7880 19120 7895
rect 19080 7860 19090 7880
rect 19110 7860 19120 7880
rect 19080 7830 19120 7860
rect 19080 7810 19090 7830
rect 19110 7810 19120 7830
rect 19080 7780 19120 7810
rect 19080 7760 19090 7780
rect 19110 7760 19120 7780
rect 19080 7730 19120 7760
rect 19080 7710 19090 7730
rect 19110 7710 19120 7730
rect 19080 7680 19120 7710
rect 19080 7660 19090 7680
rect 19110 7660 19120 7680
rect 19080 7630 19120 7660
rect 19080 7610 19090 7630
rect 19110 7610 19120 7630
rect 19080 7580 19120 7610
rect 19080 7560 19090 7580
rect 19110 7560 19120 7580
rect 19080 7530 19120 7560
rect 19080 7510 19090 7530
rect 19110 7510 19120 7530
rect 19080 7495 19120 7510
rect 19140 7880 19180 7895
rect 19140 7860 19150 7880
rect 19170 7860 19180 7880
rect 19140 7830 19180 7860
rect 19140 7810 19150 7830
rect 19170 7810 19180 7830
rect 19140 7780 19180 7810
rect 19140 7760 19150 7780
rect 19170 7760 19180 7780
rect 19140 7730 19180 7760
rect 19140 7710 19150 7730
rect 19170 7710 19180 7730
rect 19140 7680 19180 7710
rect 19140 7660 19150 7680
rect 19170 7660 19180 7680
rect 19140 7630 19180 7660
rect 19140 7610 19150 7630
rect 19170 7610 19180 7630
rect 19140 7580 19180 7610
rect 19140 7560 19150 7580
rect 19170 7560 19180 7580
rect 19140 7530 19180 7560
rect 19140 7510 19150 7530
rect 19170 7510 19180 7530
rect 19140 7495 19180 7510
rect 19200 7880 19240 7895
rect 19200 7860 19210 7880
rect 19230 7860 19240 7880
rect 19200 7830 19240 7860
rect 19200 7810 19210 7830
rect 19230 7810 19240 7830
rect 19200 7780 19240 7810
rect 19200 7760 19210 7780
rect 19230 7760 19240 7780
rect 19200 7730 19240 7760
rect 19200 7710 19210 7730
rect 19230 7710 19240 7730
rect 19200 7680 19240 7710
rect 19200 7660 19210 7680
rect 19230 7660 19240 7680
rect 19200 7630 19240 7660
rect 19200 7610 19210 7630
rect 19230 7610 19240 7630
rect 19200 7580 19240 7610
rect 19200 7560 19210 7580
rect 19230 7560 19240 7580
rect 19200 7530 19240 7560
rect 19200 7510 19210 7530
rect 19230 7510 19240 7530
rect 19200 7495 19240 7510
rect 19260 7880 19300 7895
rect 19260 7860 19270 7880
rect 19290 7860 19300 7880
rect 19260 7830 19300 7860
rect 19260 7810 19270 7830
rect 19290 7810 19300 7830
rect 19260 7780 19300 7810
rect 19260 7760 19270 7780
rect 19290 7760 19300 7780
rect 19260 7730 19300 7760
rect 19260 7710 19270 7730
rect 19290 7710 19300 7730
rect 19260 7680 19300 7710
rect 19260 7660 19270 7680
rect 19290 7660 19300 7680
rect 19260 7630 19300 7660
rect 19260 7610 19270 7630
rect 19290 7610 19300 7630
rect 19260 7580 19300 7610
rect 19260 7560 19270 7580
rect 19290 7560 19300 7580
rect 19260 7530 19300 7560
rect 19260 7510 19270 7530
rect 19290 7510 19300 7530
rect 19260 7495 19300 7510
rect 19320 7880 19360 7895
rect 19320 7860 19330 7880
rect 19350 7860 19360 7880
rect 19320 7830 19360 7860
rect 19320 7810 19330 7830
rect 19350 7810 19360 7830
rect 19320 7780 19360 7810
rect 19320 7760 19330 7780
rect 19350 7760 19360 7780
rect 19320 7730 19360 7760
rect 19320 7710 19330 7730
rect 19350 7710 19360 7730
rect 19320 7680 19360 7710
rect 19320 7660 19330 7680
rect 19350 7660 19360 7680
rect 19320 7630 19360 7660
rect 19320 7610 19330 7630
rect 19350 7610 19360 7630
rect 19320 7580 19360 7610
rect 19320 7560 19330 7580
rect 19350 7560 19360 7580
rect 19320 7530 19360 7560
rect 19320 7510 19330 7530
rect 19350 7510 19360 7530
rect 19320 7495 19360 7510
rect 19380 7880 19420 7895
rect 19380 7860 19390 7880
rect 19410 7860 19420 7880
rect 19380 7830 19420 7860
rect 19380 7810 19390 7830
rect 19410 7810 19420 7830
rect 19380 7780 19420 7810
rect 19380 7760 19390 7780
rect 19410 7760 19420 7780
rect 19380 7730 19420 7760
rect 19380 7710 19390 7730
rect 19410 7710 19420 7730
rect 19380 7680 19420 7710
rect 19380 7660 19390 7680
rect 19410 7660 19420 7680
rect 19380 7630 19420 7660
rect 19380 7610 19390 7630
rect 19410 7610 19420 7630
rect 19380 7580 19420 7610
rect 19380 7560 19390 7580
rect 19410 7560 19420 7580
rect 19380 7530 19420 7560
rect 19380 7510 19390 7530
rect 19410 7510 19420 7530
rect 19380 7495 19420 7510
rect 19440 7880 19480 7895
rect 19440 7860 19450 7880
rect 19470 7860 19480 7880
rect 19440 7830 19480 7860
rect 19440 7810 19450 7830
rect 19470 7810 19480 7830
rect 19440 7780 19480 7810
rect 19440 7760 19450 7780
rect 19470 7760 19480 7780
rect 19440 7730 19480 7760
rect 19440 7710 19450 7730
rect 19470 7710 19480 7730
rect 19440 7680 19480 7710
rect 19440 7660 19450 7680
rect 19470 7660 19480 7680
rect 19440 7630 19480 7660
rect 19440 7610 19450 7630
rect 19470 7610 19480 7630
rect 19440 7580 19480 7610
rect 19440 7560 19450 7580
rect 19470 7560 19480 7580
rect 19440 7530 19480 7560
rect 19440 7510 19450 7530
rect 19470 7510 19480 7530
rect 19440 7495 19480 7510
rect 19500 7880 19540 7895
rect 19500 7860 19510 7880
rect 19530 7860 19540 7880
rect 19500 7830 19540 7860
rect 19500 7810 19510 7830
rect 19530 7810 19540 7830
rect 19500 7780 19540 7810
rect 19500 7760 19510 7780
rect 19530 7760 19540 7780
rect 19500 7730 19540 7760
rect 19500 7710 19510 7730
rect 19530 7710 19540 7730
rect 19500 7680 19540 7710
rect 19500 7660 19510 7680
rect 19530 7660 19540 7680
rect 19500 7630 19540 7660
rect 19500 7610 19510 7630
rect 19530 7610 19540 7630
rect 19500 7580 19540 7610
rect 19500 7560 19510 7580
rect 19530 7560 19540 7580
rect 19500 7530 19540 7560
rect 19500 7510 19510 7530
rect 19530 7510 19540 7530
rect 19500 7495 19540 7510
rect 19560 7880 19600 7895
rect 19560 7860 19570 7880
rect 19590 7860 19600 7880
rect 19560 7830 19600 7860
rect 19560 7810 19570 7830
rect 19590 7810 19600 7830
rect 19560 7780 19600 7810
rect 19560 7760 19570 7780
rect 19590 7760 19600 7780
rect 19560 7730 19600 7760
rect 19560 7710 19570 7730
rect 19590 7710 19600 7730
rect 19560 7680 19600 7710
rect 19560 7660 19570 7680
rect 19590 7660 19600 7680
rect 19560 7630 19600 7660
rect 19560 7610 19570 7630
rect 19590 7610 19600 7630
rect 19560 7580 19600 7610
rect 19560 7560 19570 7580
rect 19590 7560 19600 7580
rect 19560 7530 19600 7560
rect 19560 7510 19570 7530
rect 19590 7510 19600 7530
rect 19560 7495 19600 7510
rect 19620 7880 19660 7895
rect 19620 7860 19630 7880
rect 19650 7860 19660 7880
rect 19620 7830 19660 7860
rect 19620 7810 19630 7830
rect 19650 7810 19660 7830
rect 19620 7780 19660 7810
rect 19620 7760 19630 7780
rect 19650 7760 19660 7780
rect 19620 7730 19660 7760
rect 19620 7710 19630 7730
rect 19650 7710 19660 7730
rect 19620 7680 19660 7710
rect 19620 7660 19630 7680
rect 19650 7660 19660 7680
rect 19620 7630 19660 7660
rect 19620 7610 19630 7630
rect 19650 7610 19660 7630
rect 19620 7580 19660 7610
rect 19620 7560 19630 7580
rect 19650 7560 19660 7580
rect 19620 7530 19660 7560
rect 19620 7510 19630 7530
rect 19650 7510 19660 7530
rect 19620 7495 19660 7510
rect 19680 7880 19720 7895
rect 19680 7860 19690 7880
rect 19710 7860 19720 7880
rect 19680 7830 19720 7860
rect 19680 7810 19690 7830
rect 19710 7810 19720 7830
rect 19680 7780 19720 7810
rect 19680 7760 19690 7780
rect 19710 7760 19720 7780
rect 19680 7730 19720 7760
rect 19680 7710 19690 7730
rect 19710 7710 19720 7730
rect 19680 7680 19720 7710
rect 19680 7660 19690 7680
rect 19710 7660 19720 7680
rect 19680 7630 19720 7660
rect 19680 7610 19690 7630
rect 19710 7610 19720 7630
rect 19680 7580 19720 7610
rect 19680 7560 19690 7580
rect 19710 7560 19720 7580
rect 19680 7530 19720 7560
rect 19680 7510 19690 7530
rect 19710 7510 19720 7530
rect 19680 7495 19720 7510
rect 19740 7880 19780 7895
rect 19740 7860 19750 7880
rect 19770 7860 19780 7880
rect 19740 7830 19780 7860
rect 19740 7810 19750 7830
rect 19770 7810 19780 7830
rect 19740 7780 19780 7810
rect 19740 7760 19750 7780
rect 19770 7760 19780 7780
rect 19740 7730 19780 7760
rect 19740 7710 19750 7730
rect 19770 7710 19780 7730
rect 19740 7680 19780 7710
rect 19740 7660 19750 7680
rect 19770 7660 19780 7680
rect 19740 7630 19780 7660
rect 19740 7610 19750 7630
rect 19770 7610 19780 7630
rect 19740 7580 19780 7610
rect 19740 7560 19750 7580
rect 19770 7560 19780 7580
rect 19740 7530 19780 7560
rect 19740 7510 19750 7530
rect 19770 7510 19780 7530
rect 19740 7495 19780 7510
rect 19800 7880 19840 7895
rect 19800 7860 19810 7880
rect 19830 7860 19840 7880
rect 19800 7830 19840 7860
rect 19800 7810 19810 7830
rect 19830 7810 19840 7830
rect 19800 7780 19840 7810
rect 19800 7760 19810 7780
rect 19830 7760 19840 7780
rect 19800 7730 19840 7760
rect 19800 7710 19810 7730
rect 19830 7710 19840 7730
rect 19800 7680 19840 7710
rect 19800 7660 19810 7680
rect 19830 7660 19840 7680
rect 19800 7630 19840 7660
rect 19800 7610 19810 7630
rect 19830 7610 19840 7630
rect 19800 7580 19840 7610
rect 19800 7560 19810 7580
rect 19830 7560 19840 7580
rect 19800 7530 19840 7560
rect 19800 7510 19810 7530
rect 19830 7510 19840 7530
rect 19800 7495 19840 7510
rect 19860 7880 19900 7895
rect 19860 7860 19870 7880
rect 19890 7860 19900 7880
rect 19860 7830 19900 7860
rect 19860 7810 19870 7830
rect 19890 7810 19900 7830
rect 19860 7780 19900 7810
rect 19860 7760 19870 7780
rect 19890 7760 19900 7780
rect 19860 7730 19900 7760
rect 19860 7710 19870 7730
rect 19890 7710 19900 7730
rect 19860 7680 19900 7710
rect 19860 7660 19870 7680
rect 19890 7660 19900 7680
rect 19860 7630 19900 7660
rect 19860 7610 19870 7630
rect 19890 7610 19900 7630
rect 19860 7580 19900 7610
rect 19860 7560 19870 7580
rect 19890 7560 19900 7580
rect 19860 7530 19900 7560
rect 19860 7510 19870 7530
rect 19890 7510 19900 7530
rect 19860 7495 19900 7510
rect 19920 7880 19960 7895
rect 19920 7860 19930 7880
rect 19950 7860 19960 7880
rect 19920 7830 19960 7860
rect 19920 7810 19930 7830
rect 19950 7810 19960 7830
rect 19920 7780 19960 7810
rect 19920 7760 19930 7780
rect 19950 7760 19960 7780
rect 19920 7730 19960 7760
rect 19920 7710 19930 7730
rect 19950 7710 19960 7730
rect 19920 7680 19960 7710
rect 19920 7660 19930 7680
rect 19950 7660 19960 7680
rect 19920 7630 19960 7660
rect 19920 7610 19930 7630
rect 19950 7610 19960 7630
rect 19920 7580 19960 7610
rect 19920 7560 19930 7580
rect 19950 7560 19960 7580
rect 19920 7530 19960 7560
rect 19920 7510 19930 7530
rect 19950 7510 19960 7530
rect 19920 7495 19960 7510
rect 19980 7880 20020 7895
rect 19980 7860 19990 7880
rect 20010 7860 20020 7880
rect 19980 7830 20020 7860
rect 19980 7810 19990 7830
rect 20010 7810 20020 7830
rect 19980 7780 20020 7810
rect 19980 7760 19990 7780
rect 20010 7760 20020 7780
rect 19980 7730 20020 7760
rect 19980 7710 19990 7730
rect 20010 7710 20020 7730
rect 19980 7680 20020 7710
rect 19980 7660 19990 7680
rect 20010 7660 20020 7680
rect 19980 7630 20020 7660
rect 19980 7610 19990 7630
rect 20010 7610 20020 7630
rect 19980 7580 20020 7610
rect 19980 7560 19990 7580
rect 20010 7560 20020 7580
rect 19980 7530 20020 7560
rect 19980 7510 19990 7530
rect 20010 7510 20020 7530
rect 19980 7495 20020 7510
rect 20040 7880 20080 7895
rect 20040 7860 20050 7880
rect 20070 7860 20080 7880
rect 20040 7830 20080 7860
rect 20040 7810 20050 7830
rect 20070 7810 20080 7830
rect 20040 7780 20080 7810
rect 20040 7760 20050 7780
rect 20070 7760 20080 7780
rect 20040 7730 20080 7760
rect 20040 7710 20050 7730
rect 20070 7710 20080 7730
rect 20040 7680 20080 7710
rect 20040 7660 20050 7680
rect 20070 7660 20080 7680
rect 20040 7630 20080 7660
rect 20040 7610 20050 7630
rect 20070 7610 20080 7630
rect 20040 7580 20080 7610
rect 20040 7560 20050 7580
rect 20070 7560 20080 7580
rect 20040 7530 20080 7560
rect 20040 7510 20050 7530
rect 20070 7510 20080 7530
rect 20390 7605 20430 7620
rect 20390 7585 20400 7605
rect 20420 7585 20430 7605
rect 20390 7555 20430 7585
rect 20390 7535 20400 7555
rect 20420 7535 20430 7555
rect 20390 7520 20430 7535
rect 20445 7605 20485 7620
rect 20445 7585 20455 7605
rect 20475 7585 20485 7605
rect 20445 7555 20485 7585
rect 20445 7535 20455 7555
rect 20475 7535 20485 7555
rect 20445 7520 20485 7535
rect 20500 7605 20540 7620
rect 20500 7585 20510 7605
rect 20530 7585 20540 7605
rect 20500 7555 20540 7585
rect 20500 7535 20510 7555
rect 20530 7535 20540 7555
rect 20500 7520 20540 7535
rect 20555 7605 20595 7620
rect 20555 7585 20565 7605
rect 20585 7585 20595 7605
rect 20555 7555 20595 7585
rect 20555 7535 20565 7555
rect 20585 7535 20595 7555
rect 20555 7520 20595 7535
rect 20610 7605 20650 7620
rect 20610 7585 20620 7605
rect 20640 7585 20650 7605
rect 20610 7555 20650 7585
rect 20610 7535 20620 7555
rect 20640 7535 20650 7555
rect 20610 7520 20650 7535
rect 20665 7605 20705 7620
rect 20665 7585 20675 7605
rect 20695 7585 20705 7605
rect 20665 7555 20705 7585
rect 20665 7535 20675 7555
rect 20695 7535 20705 7555
rect 20665 7520 20705 7535
rect 20720 7605 20760 7620
rect 20720 7585 20730 7605
rect 20750 7585 20760 7605
rect 20720 7555 20760 7585
rect 20720 7535 20730 7555
rect 20750 7535 20760 7555
rect 20720 7520 20760 7535
rect 20775 7605 20815 7620
rect 20775 7585 20785 7605
rect 20805 7585 20815 7605
rect 20775 7555 20815 7585
rect 20775 7535 20785 7555
rect 20805 7535 20815 7555
rect 20775 7520 20815 7535
rect 20830 7605 20870 7620
rect 20830 7585 20840 7605
rect 20860 7585 20870 7605
rect 20830 7555 20870 7585
rect 20830 7535 20840 7555
rect 20860 7535 20870 7555
rect 20830 7520 20870 7535
rect 20885 7605 20925 7620
rect 20885 7585 20895 7605
rect 20915 7585 20925 7605
rect 20885 7555 20925 7585
rect 20885 7535 20895 7555
rect 20915 7535 20925 7555
rect 20885 7520 20925 7535
rect 20940 7605 20980 7620
rect 20940 7585 20950 7605
rect 20970 7585 20980 7605
rect 20940 7555 20980 7585
rect 20940 7535 20950 7555
rect 20970 7535 20980 7555
rect 20940 7520 20980 7535
rect 20995 7605 21035 7620
rect 20995 7585 21005 7605
rect 21025 7585 21035 7605
rect 20995 7555 21035 7585
rect 20995 7535 21005 7555
rect 21025 7535 21035 7555
rect 20995 7520 21035 7535
rect 21050 7605 21090 7620
rect 21050 7585 21060 7605
rect 21080 7585 21090 7605
rect 21050 7555 21090 7585
rect 21050 7535 21060 7555
rect 21080 7535 21090 7555
rect 21050 7520 21090 7535
rect 21105 7605 21145 7620
rect 21105 7585 21115 7605
rect 21135 7585 21145 7605
rect 21105 7555 21145 7585
rect 21105 7535 21115 7555
rect 21135 7535 21145 7555
rect 21105 7520 21145 7535
rect 21160 7605 21200 7620
rect 21160 7585 21170 7605
rect 21190 7585 21200 7605
rect 21160 7555 21200 7585
rect 21160 7535 21170 7555
rect 21190 7535 21200 7555
rect 21160 7520 21200 7535
rect 21215 7605 21255 7620
rect 21215 7585 21225 7605
rect 21245 7585 21255 7605
rect 21215 7555 21255 7585
rect 21215 7535 21225 7555
rect 21245 7535 21255 7555
rect 21215 7520 21255 7535
rect 21270 7605 21310 7620
rect 21270 7585 21280 7605
rect 21300 7585 21310 7605
rect 21270 7555 21310 7585
rect 21270 7535 21280 7555
rect 21300 7535 21310 7555
rect 21270 7520 21310 7535
rect 21325 7605 21365 7620
rect 21325 7585 21335 7605
rect 21355 7585 21365 7605
rect 21325 7555 21365 7585
rect 21325 7535 21335 7555
rect 21355 7535 21365 7555
rect 21325 7520 21365 7535
rect 21380 7605 21420 7620
rect 21380 7585 21390 7605
rect 21410 7585 21420 7605
rect 21380 7555 21420 7585
rect 21380 7535 21390 7555
rect 21410 7535 21420 7555
rect 21380 7520 21420 7535
rect 21435 7605 21475 7620
rect 21435 7585 21445 7605
rect 21465 7585 21475 7605
rect 21435 7555 21475 7585
rect 21435 7535 21445 7555
rect 21465 7535 21475 7555
rect 21435 7520 21475 7535
rect 21490 7605 21530 7620
rect 21490 7585 21500 7605
rect 21520 7585 21530 7605
rect 21490 7555 21530 7585
rect 21490 7535 21500 7555
rect 21520 7535 21530 7555
rect 21490 7520 21530 7535
rect 21545 7605 21585 7620
rect 21545 7585 21555 7605
rect 21575 7585 21585 7605
rect 21545 7555 21585 7585
rect 21545 7535 21555 7555
rect 21575 7535 21585 7555
rect 21545 7520 21585 7535
rect 21600 7605 21640 7620
rect 21600 7585 21610 7605
rect 21630 7585 21640 7605
rect 21600 7555 21640 7585
rect 21600 7535 21610 7555
rect 21630 7535 21640 7555
rect 21600 7520 21640 7535
rect 20040 7495 20080 7510
rect 9680 7155 9720 7170
rect 9680 7135 9690 7155
rect 9710 7135 9720 7155
rect 9680 7105 9720 7135
rect 9680 7085 9690 7105
rect 9710 7085 9720 7105
rect 9680 7055 9720 7085
rect 9680 7035 9690 7055
rect 9710 7035 9720 7055
rect 9680 7020 9720 7035
rect 9735 7155 9775 7170
rect 9735 7135 9745 7155
rect 9765 7135 9775 7155
rect 9735 7105 9775 7135
rect 9735 7085 9745 7105
rect 9765 7085 9775 7105
rect 9735 7055 9775 7085
rect 9735 7035 9745 7055
rect 9765 7035 9775 7055
rect 9735 7020 9775 7035
rect 9790 7155 9830 7170
rect 9790 7135 9800 7155
rect 9820 7135 9830 7155
rect 9790 7105 9830 7135
rect 9790 7085 9800 7105
rect 9820 7085 9830 7105
rect 9790 7055 9830 7085
rect 9790 7035 9800 7055
rect 9820 7035 9830 7055
rect 9790 7020 9830 7035
rect 9845 7155 9885 7170
rect 9845 7135 9855 7155
rect 9875 7135 9885 7155
rect 9845 7105 9885 7135
rect 9845 7085 9855 7105
rect 9875 7085 9885 7105
rect 9845 7055 9885 7085
rect 9845 7035 9855 7055
rect 9875 7035 9885 7055
rect 9845 7020 9885 7035
rect 9900 7155 9940 7170
rect 9900 7135 9910 7155
rect 9930 7135 9940 7155
rect 9900 7105 9940 7135
rect 9900 7085 9910 7105
rect 9930 7085 9940 7105
rect 9900 7055 9940 7085
rect 9900 7035 9910 7055
rect 9930 7035 9940 7055
rect 9900 7020 9940 7035
rect 9955 7155 9995 7170
rect 9955 7135 9965 7155
rect 9985 7135 9995 7155
rect 9955 7105 9995 7135
rect 9955 7085 9965 7105
rect 9985 7085 9995 7105
rect 9955 7055 9995 7085
rect 9955 7035 9965 7055
rect 9985 7035 9995 7055
rect 9955 7020 9995 7035
rect 10010 7155 10050 7170
rect 10010 7135 10020 7155
rect 10040 7135 10050 7155
rect 10010 7105 10050 7135
rect 10010 7085 10020 7105
rect 10040 7085 10050 7105
rect 10010 7055 10050 7085
rect 10010 7035 10020 7055
rect 10040 7035 10050 7055
rect 10010 7020 10050 7035
rect 10065 7155 10105 7170
rect 10065 7135 10075 7155
rect 10095 7135 10105 7155
rect 10065 7105 10105 7135
rect 10065 7085 10075 7105
rect 10095 7085 10105 7105
rect 10065 7055 10105 7085
rect 10065 7035 10075 7055
rect 10095 7035 10105 7055
rect 10065 7020 10105 7035
rect 10120 7155 10160 7170
rect 10120 7135 10130 7155
rect 10150 7135 10160 7155
rect 10120 7105 10160 7135
rect 10120 7085 10130 7105
rect 10150 7085 10160 7105
rect 10120 7055 10160 7085
rect 10120 7035 10130 7055
rect 10150 7035 10160 7055
rect 10120 7020 10160 7035
rect 10175 7155 10215 7170
rect 10175 7135 10185 7155
rect 10205 7135 10215 7155
rect 10175 7105 10215 7135
rect 10175 7085 10185 7105
rect 10205 7085 10215 7105
rect 10175 7055 10215 7085
rect 10175 7035 10185 7055
rect 10205 7035 10215 7055
rect 10175 7020 10215 7035
rect 10230 7155 10270 7170
rect 10230 7135 10240 7155
rect 10260 7135 10270 7155
rect 10230 7105 10270 7135
rect 10230 7085 10240 7105
rect 10260 7085 10270 7105
rect 10230 7055 10270 7085
rect 10230 7035 10240 7055
rect 10260 7035 10270 7055
rect 10230 7020 10270 7035
rect 10285 7155 10325 7170
rect 10285 7135 10295 7155
rect 10315 7135 10325 7155
rect 10285 7105 10325 7135
rect 10285 7085 10295 7105
rect 10315 7085 10325 7105
rect 10285 7055 10325 7085
rect 10285 7035 10295 7055
rect 10315 7035 10325 7055
rect 10285 7020 10325 7035
rect 10340 7155 10380 7170
rect 10340 7135 10350 7155
rect 10370 7135 10380 7155
rect 10340 7105 10380 7135
rect 10340 7085 10350 7105
rect 10370 7085 10380 7105
rect 10340 7055 10380 7085
rect 10340 7035 10350 7055
rect 10370 7035 10380 7055
rect 10340 7020 10380 7035
rect 10395 7155 10435 7170
rect 10395 7135 10405 7155
rect 10425 7135 10435 7155
rect 10395 7105 10435 7135
rect 10395 7085 10405 7105
rect 10425 7085 10435 7105
rect 10395 7055 10435 7085
rect 10395 7035 10405 7055
rect 10425 7035 10435 7055
rect 10395 7020 10435 7035
rect 10450 7155 10490 7170
rect 10450 7135 10460 7155
rect 10480 7135 10490 7155
rect 10450 7105 10490 7135
rect 10450 7085 10460 7105
rect 10480 7085 10490 7105
rect 10450 7055 10490 7085
rect 10450 7035 10460 7055
rect 10480 7035 10490 7055
rect 10450 7020 10490 7035
rect 10505 7155 10545 7170
rect 10505 7135 10515 7155
rect 10535 7135 10545 7155
rect 10505 7105 10545 7135
rect 10505 7085 10515 7105
rect 10535 7085 10545 7105
rect 10505 7055 10545 7085
rect 10505 7035 10515 7055
rect 10535 7035 10545 7055
rect 10505 7020 10545 7035
rect 10560 7155 10600 7170
rect 10560 7135 10570 7155
rect 10590 7135 10600 7155
rect 10560 7105 10600 7135
rect 10560 7085 10570 7105
rect 10590 7085 10600 7105
rect 10560 7055 10600 7085
rect 10560 7035 10570 7055
rect 10590 7035 10600 7055
rect 10560 7020 10600 7035
rect 10615 7155 10655 7170
rect 10615 7135 10625 7155
rect 10645 7135 10655 7155
rect 10615 7105 10655 7135
rect 10615 7085 10625 7105
rect 10645 7085 10655 7105
rect 10615 7055 10655 7085
rect 10615 7035 10625 7055
rect 10645 7035 10655 7055
rect 10615 7020 10655 7035
rect 10670 7155 10710 7170
rect 10670 7135 10680 7155
rect 10700 7135 10710 7155
rect 10670 7105 10710 7135
rect 10670 7085 10680 7105
rect 10700 7085 10710 7105
rect 10670 7055 10710 7085
rect 10670 7035 10680 7055
rect 10700 7035 10710 7055
rect 10670 7020 10710 7035
rect 10725 7155 10765 7170
rect 10725 7135 10735 7155
rect 10755 7135 10765 7155
rect 10725 7105 10765 7135
rect 10725 7085 10735 7105
rect 10755 7085 10765 7105
rect 10725 7055 10765 7085
rect 10725 7035 10735 7055
rect 10755 7035 10765 7055
rect 10725 7020 10765 7035
rect 10780 7155 10820 7170
rect 10780 7135 10790 7155
rect 10810 7135 10820 7155
rect 10780 7105 10820 7135
rect 10780 7085 10790 7105
rect 10810 7085 10820 7105
rect 10780 7055 10820 7085
rect 10780 7035 10790 7055
rect 10810 7035 10820 7055
rect 10780 7020 10820 7035
rect 10835 7155 10875 7170
rect 10835 7135 10845 7155
rect 10865 7135 10875 7155
rect 10835 7105 10875 7135
rect 10835 7085 10845 7105
rect 10865 7085 10875 7105
rect 10835 7055 10875 7085
rect 10835 7035 10845 7055
rect 10865 7035 10875 7055
rect 10835 7020 10875 7035
rect 10890 7155 10930 7170
rect 12895 7155 12935 7170
rect 10890 7135 10900 7155
rect 10920 7135 10930 7155
rect 10890 7105 10930 7135
rect 12895 7135 12905 7155
rect 12925 7135 12935 7155
rect 10890 7085 10900 7105
rect 10920 7085 10930 7105
rect 10890 7055 10930 7085
rect 10890 7035 10900 7055
rect 10920 7035 10930 7055
rect 10890 7020 10930 7035
rect 11275 7115 11315 7130
rect 11275 7095 11285 7115
rect 11305 7095 11315 7115
rect 11275 7065 11315 7095
rect 11275 7045 11285 7065
rect 11305 7045 11315 7065
rect 11275 7015 11315 7045
rect 11275 6995 11285 7015
rect 11305 6995 11315 7015
rect 11275 6980 11315 6995
rect 11330 7115 11370 7130
rect 11330 7095 11340 7115
rect 11360 7095 11370 7115
rect 11330 7065 11370 7095
rect 11330 7045 11340 7065
rect 11360 7045 11370 7065
rect 11330 7015 11370 7045
rect 11330 6995 11340 7015
rect 11360 6995 11370 7015
rect 11330 6980 11370 6995
rect 11385 7115 11425 7130
rect 11385 7095 11395 7115
rect 11415 7095 11425 7115
rect 11385 7065 11425 7095
rect 11385 7045 11395 7065
rect 11415 7045 11425 7065
rect 11385 7015 11425 7045
rect 11385 6995 11395 7015
rect 11415 6995 11425 7015
rect 11385 6980 11425 6995
rect 11440 7115 11480 7130
rect 11440 7095 11450 7115
rect 11470 7095 11480 7115
rect 11440 7065 11480 7095
rect 11440 7045 11450 7065
rect 11470 7045 11480 7065
rect 11440 7015 11480 7045
rect 11440 6995 11450 7015
rect 11470 6995 11480 7015
rect 11440 6980 11480 6995
rect 11495 7115 11535 7130
rect 11495 7095 11505 7115
rect 11525 7095 11535 7115
rect 11495 7065 11535 7095
rect 11495 7045 11505 7065
rect 11525 7045 11535 7065
rect 11495 7015 11535 7045
rect 11495 6995 11505 7015
rect 11525 6995 11535 7015
rect 11495 6980 11535 6995
rect 11550 7115 11590 7130
rect 11550 7095 11560 7115
rect 11580 7095 11590 7115
rect 11550 7065 11590 7095
rect 11550 7045 11560 7065
rect 11580 7045 11590 7065
rect 11550 7015 11590 7045
rect 11550 6995 11560 7015
rect 11580 6995 11590 7015
rect 11550 6980 11590 6995
rect 11605 7115 11645 7130
rect 11605 7095 11615 7115
rect 11635 7095 11645 7115
rect 11605 7065 11645 7095
rect 11605 7045 11615 7065
rect 11635 7045 11645 7065
rect 11605 7015 11645 7045
rect 11605 6995 11615 7015
rect 11635 6995 11645 7015
rect 11605 6980 11645 6995
rect 11660 7115 11700 7130
rect 11660 7095 11670 7115
rect 11690 7095 11700 7115
rect 11660 7065 11700 7095
rect 11660 7045 11670 7065
rect 11690 7045 11700 7065
rect 11660 7015 11700 7045
rect 11660 6995 11670 7015
rect 11690 6995 11700 7015
rect 11660 6980 11700 6995
rect 11715 7115 11755 7130
rect 11715 7095 11725 7115
rect 11745 7095 11755 7115
rect 11715 7065 11755 7095
rect 11715 7045 11725 7065
rect 11745 7045 11755 7065
rect 11715 7015 11755 7045
rect 11715 6995 11725 7015
rect 11745 6995 11755 7015
rect 11715 6980 11755 6995
rect 11770 7115 11810 7130
rect 11770 7095 11780 7115
rect 11800 7095 11810 7115
rect 11770 7065 11810 7095
rect 11770 7045 11780 7065
rect 11800 7045 11810 7065
rect 11770 7015 11810 7045
rect 11770 6995 11780 7015
rect 11800 6995 11810 7015
rect 11770 6980 11810 6995
rect 11825 7115 11865 7130
rect 11825 7095 11835 7115
rect 11855 7095 11865 7115
rect 11825 7065 11865 7095
rect 11825 7045 11835 7065
rect 11855 7045 11865 7065
rect 11825 7015 11865 7045
rect 11825 6995 11835 7015
rect 11855 6995 11865 7015
rect 11825 6980 11865 6995
rect 11880 7115 11920 7130
rect 11880 7095 11890 7115
rect 11910 7095 11920 7115
rect 11880 7065 11920 7095
rect 11880 7045 11890 7065
rect 11910 7045 11920 7065
rect 11880 7015 11920 7045
rect 11880 6995 11890 7015
rect 11910 6995 11920 7015
rect 11880 6980 11920 6995
rect 11935 7115 11975 7130
rect 11935 7095 11945 7115
rect 11965 7095 11975 7115
rect 11935 7065 11975 7095
rect 11935 7045 11945 7065
rect 11965 7045 11975 7065
rect 11935 7015 11975 7045
rect 11935 6995 11945 7015
rect 11965 6995 11975 7015
rect 11935 6980 11975 6995
rect 11990 7115 12030 7130
rect 11990 7095 12000 7115
rect 12020 7095 12030 7115
rect 11990 7065 12030 7095
rect 11990 7045 12000 7065
rect 12020 7045 12030 7065
rect 11990 7015 12030 7045
rect 11990 6995 12000 7015
rect 12020 6995 12030 7015
rect 11990 6980 12030 6995
rect 12045 7115 12085 7130
rect 12045 7095 12055 7115
rect 12075 7095 12085 7115
rect 12045 7065 12085 7095
rect 12045 7045 12055 7065
rect 12075 7045 12085 7065
rect 12045 7015 12085 7045
rect 12045 6995 12055 7015
rect 12075 6995 12085 7015
rect 12045 6980 12085 6995
rect 12100 7115 12140 7130
rect 12100 7095 12110 7115
rect 12130 7095 12140 7115
rect 12100 7065 12140 7095
rect 12100 7045 12110 7065
rect 12130 7045 12140 7065
rect 12100 7015 12140 7045
rect 12100 6995 12110 7015
rect 12130 6995 12140 7015
rect 12100 6980 12140 6995
rect 12155 7115 12195 7130
rect 12155 7095 12165 7115
rect 12185 7095 12195 7115
rect 12155 7065 12195 7095
rect 12155 7045 12165 7065
rect 12185 7045 12195 7065
rect 12155 7015 12195 7045
rect 12155 6995 12165 7015
rect 12185 6995 12195 7015
rect 12155 6980 12195 6995
rect 12210 7115 12250 7130
rect 12210 7095 12220 7115
rect 12240 7095 12250 7115
rect 12210 7065 12250 7095
rect 12210 7045 12220 7065
rect 12240 7045 12250 7065
rect 12210 7015 12250 7045
rect 12210 6995 12220 7015
rect 12240 6995 12250 7015
rect 12210 6980 12250 6995
rect 12265 7115 12305 7130
rect 12265 7095 12275 7115
rect 12295 7095 12305 7115
rect 12265 7065 12305 7095
rect 12265 7045 12275 7065
rect 12295 7045 12305 7065
rect 12265 7015 12305 7045
rect 12265 6995 12275 7015
rect 12295 6995 12305 7015
rect 12265 6980 12305 6995
rect 12320 7115 12360 7130
rect 12320 7095 12330 7115
rect 12350 7095 12360 7115
rect 12320 7065 12360 7095
rect 12320 7045 12330 7065
rect 12350 7045 12360 7065
rect 12320 7015 12360 7045
rect 12320 6995 12330 7015
rect 12350 6995 12360 7015
rect 12320 6980 12360 6995
rect 12375 7115 12415 7130
rect 12375 7095 12385 7115
rect 12405 7095 12415 7115
rect 12375 7065 12415 7095
rect 12375 7045 12385 7065
rect 12405 7045 12415 7065
rect 12375 7015 12415 7045
rect 12375 6995 12385 7015
rect 12405 6995 12415 7015
rect 12375 6980 12415 6995
rect 12430 7115 12470 7130
rect 12430 7095 12440 7115
rect 12460 7095 12470 7115
rect 12430 7065 12470 7095
rect 12430 7045 12440 7065
rect 12460 7045 12470 7065
rect 12430 7015 12470 7045
rect 12430 6995 12440 7015
rect 12460 6995 12470 7015
rect 12430 6980 12470 6995
rect 12485 7115 12525 7130
rect 12485 7095 12495 7115
rect 12515 7095 12525 7115
rect 12485 7065 12525 7095
rect 12485 7045 12495 7065
rect 12515 7045 12525 7065
rect 12485 7015 12525 7045
rect 12895 7105 12935 7135
rect 12895 7085 12905 7105
rect 12925 7085 12935 7105
rect 12895 7055 12935 7085
rect 12895 7035 12905 7055
rect 12925 7035 12935 7055
rect 12895 7020 12935 7035
rect 12950 7155 12990 7170
rect 12950 7135 12960 7155
rect 12980 7135 12990 7155
rect 12950 7105 12990 7135
rect 12950 7085 12960 7105
rect 12980 7085 12990 7105
rect 12950 7055 12990 7085
rect 12950 7035 12960 7055
rect 12980 7035 12990 7055
rect 12950 7020 12990 7035
rect 13005 7155 13045 7170
rect 13005 7135 13015 7155
rect 13035 7135 13045 7155
rect 13005 7105 13045 7135
rect 13005 7085 13015 7105
rect 13035 7085 13045 7105
rect 13005 7055 13045 7085
rect 13005 7035 13015 7055
rect 13035 7035 13045 7055
rect 13005 7020 13045 7035
rect 13060 7155 13100 7170
rect 13060 7135 13070 7155
rect 13090 7135 13100 7155
rect 13060 7105 13100 7135
rect 13060 7085 13070 7105
rect 13090 7085 13100 7105
rect 13060 7055 13100 7085
rect 13060 7035 13070 7055
rect 13090 7035 13100 7055
rect 13060 7020 13100 7035
rect 13115 7155 13155 7170
rect 13115 7135 13125 7155
rect 13145 7135 13155 7155
rect 13115 7105 13155 7135
rect 13115 7085 13125 7105
rect 13145 7085 13155 7105
rect 13115 7055 13155 7085
rect 13115 7035 13125 7055
rect 13145 7035 13155 7055
rect 13115 7020 13155 7035
rect 13170 7155 13210 7170
rect 13170 7135 13180 7155
rect 13200 7135 13210 7155
rect 13170 7105 13210 7135
rect 13170 7085 13180 7105
rect 13200 7085 13210 7105
rect 13170 7055 13210 7085
rect 13170 7035 13180 7055
rect 13200 7035 13210 7055
rect 13170 7020 13210 7035
rect 13225 7155 13265 7170
rect 13225 7135 13235 7155
rect 13255 7135 13265 7155
rect 13225 7105 13265 7135
rect 13225 7085 13235 7105
rect 13255 7085 13265 7105
rect 13225 7055 13265 7085
rect 13225 7035 13235 7055
rect 13255 7035 13265 7055
rect 13225 7020 13265 7035
rect 13280 7155 13320 7170
rect 13280 7135 13290 7155
rect 13310 7135 13320 7155
rect 13280 7105 13320 7135
rect 13280 7085 13290 7105
rect 13310 7085 13320 7105
rect 13280 7055 13320 7085
rect 13280 7035 13290 7055
rect 13310 7035 13320 7055
rect 13280 7020 13320 7035
rect 13335 7155 13375 7170
rect 13335 7135 13345 7155
rect 13365 7135 13375 7155
rect 13335 7105 13375 7135
rect 13335 7085 13345 7105
rect 13365 7085 13375 7105
rect 13335 7055 13375 7085
rect 13335 7035 13345 7055
rect 13365 7035 13375 7055
rect 13335 7020 13375 7035
rect 13390 7155 13430 7170
rect 13390 7135 13400 7155
rect 13420 7135 13430 7155
rect 13390 7105 13430 7135
rect 13390 7085 13400 7105
rect 13420 7085 13430 7105
rect 13390 7055 13430 7085
rect 13390 7035 13400 7055
rect 13420 7035 13430 7055
rect 13390 7020 13430 7035
rect 13445 7155 13485 7170
rect 13445 7135 13455 7155
rect 13475 7135 13485 7155
rect 13445 7105 13485 7135
rect 13445 7085 13455 7105
rect 13475 7085 13485 7105
rect 13445 7055 13485 7085
rect 13445 7035 13455 7055
rect 13475 7035 13485 7055
rect 13445 7020 13485 7035
rect 13500 7155 13540 7170
rect 13500 7135 13510 7155
rect 13530 7135 13540 7155
rect 13500 7105 13540 7135
rect 13500 7085 13510 7105
rect 13530 7085 13540 7105
rect 13500 7055 13540 7085
rect 13500 7035 13510 7055
rect 13530 7035 13540 7055
rect 13500 7020 13540 7035
rect 13555 7155 13595 7170
rect 13555 7135 13565 7155
rect 13585 7135 13595 7155
rect 13555 7105 13595 7135
rect 13555 7085 13565 7105
rect 13585 7085 13595 7105
rect 13555 7055 13595 7085
rect 13555 7035 13565 7055
rect 13585 7035 13595 7055
rect 13555 7020 13595 7035
rect 13610 7155 13650 7170
rect 13610 7135 13620 7155
rect 13640 7135 13650 7155
rect 13610 7105 13650 7135
rect 13610 7085 13620 7105
rect 13640 7085 13650 7105
rect 13610 7055 13650 7085
rect 13610 7035 13620 7055
rect 13640 7035 13650 7055
rect 13610 7020 13650 7035
rect 13665 7155 13705 7170
rect 13665 7135 13675 7155
rect 13695 7135 13705 7155
rect 13665 7105 13705 7135
rect 13665 7085 13675 7105
rect 13695 7085 13705 7105
rect 13665 7055 13705 7085
rect 13665 7035 13675 7055
rect 13695 7035 13705 7055
rect 13665 7020 13705 7035
rect 13720 7155 13760 7170
rect 13720 7135 13730 7155
rect 13750 7135 13760 7155
rect 13720 7105 13760 7135
rect 13720 7085 13730 7105
rect 13750 7085 13760 7105
rect 13720 7055 13760 7085
rect 13720 7035 13730 7055
rect 13750 7035 13760 7055
rect 13720 7020 13760 7035
rect 13775 7155 13815 7170
rect 13775 7135 13785 7155
rect 13805 7135 13815 7155
rect 13775 7105 13815 7135
rect 13775 7085 13785 7105
rect 13805 7085 13815 7105
rect 13775 7055 13815 7085
rect 13775 7035 13785 7055
rect 13805 7035 13815 7055
rect 13775 7020 13815 7035
rect 13830 7155 13870 7170
rect 13830 7135 13840 7155
rect 13860 7135 13870 7155
rect 13830 7105 13870 7135
rect 13830 7085 13840 7105
rect 13860 7085 13870 7105
rect 13830 7055 13870 7085
rect 13830 7035 13840 7055
rect 13860 7035 13870 7055
rect 13830 7020 13870 7035
rect 13885 7155 13925 7170
rect 13885 7135 13895 7155
rect 13915 7135 13925 7155
rect 13885 7105 13925 7135
rect 13885 7085 13895 7105
rect 13915 7085 13925 7105
rect 13885 7055 13925 7085
rect 13885 7035 13895 7055
rect 13915 7035 13925 7055
rect 13885 7020 13925 7035
rect 13940 7155 13980 7170
rect 13940 7135 13950 7155
rect 13970 7135 13980 7155
rect 13940 7105 13980 7135
rect 13940 7085 13950 7105
rect 13970 7085 13980 7105
rect 13940 7055 13980 7085
rect 13940 7035 13950 7055
rect 13970 7035 13980 7055
rect 13940 7020 13980 7035
rect 13995 7155 14035 7170
rect 13995 7135 14005 7155
rect 14025 7135 14035 7155
rect 13995 7105 14035 7135
rect 13995 7085 14005 7105
rect 14025 7085 14035 7105
rect 13995 7055 14035 7085
rect 13995 7035 14005 7055
rect 14025 7035 14035 7055
rect 13995 7020 14035 7035
rect 14050 7155 14090 7170
rect 14050 7135 14060 7155
rect 14080 7135 14090 7155
rect 14050 7105 14090 7135
rect 14050 7085 14060 7105
rect 14080 7085 14090 7105
rect 14050 7055 14090 7085
rect 14050 7035 14060 7055
rect 14080 7035 14090 7055
rect 14050 7020 14090 7035
rect 14105 7155 14145 7170
rect 14105 7135 14115 7155
rect 14135 7135 14145 7155
rect 14105 7105 14145 7135
rect 14105 7085 14115 7105
rect 14135 7085 14145 7105
rect 14105 7055 14145 7085
rect 14105 7035 14115 7055
rect 14135 7035 14145 7055
rect 14105 7020 14145 7035
rect 17180 7155 17220 7170
rect 17180 7135 17190 7155
rect 17210 7135 17220 7155
rect 17180 7105 17220 7135
rect 17180 7085 17190 7105
rect 17210 7085 17220 7105
rect 17180 7055 17220 7085
rect 17180 7035 17190 7055
rect 17210 7035 17220 7055
rect 17180 7020 17220 7035
rect 17235 7155 17275 7170
rect 17235 7135 17245 7155
rect 17265 7135 17275 7155
rect 17235 7105 17275 7135
rect 17235 7085 17245 7105
rect 17265 7085 17275 7105
rect 17235 7055 17275 7085
rect 17235 7035 17245 7055
rect 17265 7035 17275 7055
rect 17235 7020 17275 7035
rect 17290 7155 17330 7170
rect 17290 7135 17300 7155
rect 17320 7135 17330 7155
rect 17290 7105 17330 7135
rect 17290 7085 17300 7105
rect 17320 7085 17330 7105
rect 17290 7055 17330 7085
rect 17290 7035 17300 7055
rect 17320 7035 17330 7055
rect 17290 7020 17330 7035
rect 17345 7155 17385 7170
rect 17345 7135 17355 7155
rect 17375 7135 17385 7155
rect 17345 7105 17385 7135
rect 17345 7085 17355 7105
rect 17375 7085 17385 7105
rect 17345 7055 17385 7085
rect 17345 7035 17355 7055
rect 17375 7035 17385 7055
rect 17345 7020 17385 7035
rect 17400 7155 17440 7170
rect 17400 7135 17410 7155
rect 17430 7135 17440 7155
rect 17400 7105 17440 7135
rect 17400 7085 17410 7105
rect 17430 7085 17440 7105
rect 17400 7055 17440 7085
rect 17400 7035 17410 7055
rect 17430 7035 17440 7055
rect 17400 7020 17440 7035
rect 17455 7155 17495 7170
rect 17455 7135 17465 7155
rect 17485 7135 17495 7155
rect 17455 7105 17495 7135
rect 17455 7085 17465 7105
rect 17485 7085 17495 7105
rect 17455 7055 17495 7085
rect 17455 7035 17465 7055
rect 17485 7035 17495 7055
rect 17455 7020 17495 7035
rect 17510 7155 17550 7170
rect 17510 7135 17520 7155
rect 17540 7135 17550 7155
rect 17510 7105 17550 7135
rect 17510 7085 17520 7105
rect 17540 7085 17550 7105
rect 17510 7055 17550 7085
rect 17510 7035 17520 7055
rect 17540 7035 17550 7055
rect 17510 7020 17550 7035
rect 17565 7155 17605 7170
rect 17565 7135 17575 7155
rect 17595 7135 17605 7155
rect 17565 7105 17605 7135
rect 17565 7085 17575 7105
rect 17595 7085 17605 7105
rect 17565 7055 17605 7085
rect 17565 7035 17575 7055
rect 17595 7035 17605 7055
rect 17565 7020 17605 7035
rect 17620 7155 17660 7170
rect 17620 7135 17630 7155
rect 17650 7135 17660 7155
rect 17620 7105 17660 7135
rect 17620 7085 17630 7105
rect 17650 7085 17660 7105
rect 17620 7055 17660 7085
rect 17620 7035 17630 7055
rect 17650 7035 17660 7055
rect 17620 7020 17660 7035
rect 17675 7155 17715 7170
rect 17675 7135 17685 7155
rect 17705 7135 17715 7155
rect 17675 7105 17715 7135
rect 17675 7085 17685 7105
rect 17705 7085 17715 7105
rect 17675 7055 17715 7085
rect 17675 7035 17685 7055
rect 17705 7035 17715 7055
rect 17675 7020 17715 7035
rect 17730 7155 17770 7170
rect 17730 7135 17740 7155
rect 17760 7135 17770 7155
rect 17730 7105 17770 7135
rect 17730 7085 17740 7105
rect 17760 7085 17770 7105
rect 17730 7055 17770 7085
rect 17730 7035 17740 7055
rect 17760 7035 17770 7055
rect 17730 7020 17770 7035
rect 17785 7155 17825 7170
rect 17785 7135 17795 7155
rect 17815 7135 17825 7155
rect 17785 7105 17825 7135
rect 17785 7085 17795 7105
rect 17815 7085 17825 7105
rect 17785 7055 17825 7085
rect 17785 7035 17795 7055
rect 17815 7035 17825 7055
rect 17785 7020 17825 7035
rect 17840 7155 17880 7170
rect 17840 7135 17850 7155
rect 17870 7135 17880 7155
rect 17840 7105 17880 7135
rect 17840 7085 17850 7105
rect 17870 7085 17880 7105
rect 17840 7055 17880 7085
rect 17840 7035 17850 7055
rect 17870 7035 17880 7055
rect 17840 7020 17880 7035
rect 17895 7155 17935 7170
rect 17895 7135 17905 7155
rect 17925 7135 17935 7155
rect 17895 7105 17935 7135
rect 17895 7085 17905 7105
rect 17925 7085 17935 7105
rect 17895 7055 17935 7085
rect 17895 7035 17905 7055
rect 17925 7035 17935 7055
rect 17895 7020 17935 7035
rect 17950 7155 17990 7170
rect 17950 7135 17960 7155
rect 17980 7135 17990 7155
rect 17950 7105 17990 7135
rect 17950 7085 17960 7105
rect 17980 7085 17990 7105
rect 17950 7055 17990 7085
rect 17950 7035 17960 7055
rect 17980 7035 17990 7055
rect 17950 7020 17990 7035
rect 18005 7155 18045 7170
rect 18005 7135 18015 7155
rect 18035 7135 18045 7155
rect 18005 7105 18045 7135
rect 18005 7085 18015 7105
rect 18035 7085 18045 7105
rect 18005 7055 18045 7085
rect 18005 7035 18015 7055
rect 18035 7035 18045 7055
rect 18005 7020 18045 7035
rect 18060 7155 18100 7170
rect 18060 7135 18070 7155
rect 18090 7135 18100 7155
rect 18060 7105 18100 7135
rect 18060 7085 18070 7105
rect 18090 7085 18100 7105
rect 18060 7055 18100 7085
rect 18060 7035 18070 7055
rect 18090 7035 18100 7055
rect 18060 7020 18100 7035
rect 18115 7155 18155 7170
rect 18115 7135 18125 7155
rect 18145 7135 18155 7155
rect 18115 7105 18155 7135
rect 18115 7085 18125 7105
rect 18145 7085 18155 7105
rect 18115 7055 18155 7085
rect 18115 7035 18125 7055
rect 18145 7035 18155 7055
rect 18115 7020 18155 7035
rect 18170 7155 18210 7170
rect 18170 7135 18180 7155
rect 18200 7135 18210 7155
rect 18170 7105 18210 7135
rect 18170 7085 18180 7105
rect 18200 7085 18210 7105
rect 18170 7055 18210 7085
rect 18170 7035 18180 7055
rect 18200 7035 18210 7055
rect 18170 7020 18210 7035
rect 18225 7155 18265 7170
rect 18225 7135 18235 7155
rect 18255 7135 18265 7155
rect 18225 7105 18265 7135
rect 18225 7085 18235 7105
rect 18255 7085 18265 7105
rect 18225 7055 18265 7085
rect 18225 7035 18235 7055
rect 18255 7035 18265 7055
rect 18225 7020 18265 7035
rect 18280 7155 18320 7170
rect 18280 7135 18290 7155
rect 18310 7135 18320 7155
rect 18280 7105 18320 7135
rect 18280 7085 18290 7105
rect 18310 7085 18320 7105
rect 18280 7055 18320 7085
rect 18280 7035 18290 7055
rect 18310 7035 18320 7055
rect 18280 7020 18320 7035
rect 18335 7155 18375 7170
rect 18335 7135 18345 7155
rect 18365 7135 18375 7155
rect 18335 7105 18375 7135
rect 18335 7085 18345 7105
rect 18365 7085 18375 7105
rect 18335 7055 18375 7085
rect 18335 7035 18345 7055
rect 18365 7035 18375 7055
rect 18335 7020 18375 7035
rect 18390 7155 18430 7170
rect 20390 7155 20430 7170
rect 18390 7135 18400 7155
rect 18420 7135 18430 7155
rect 18390 7105 18430 7135
rect 20390 7135 20400 7155
rect 20420 7135 20430 7155
rect 18390 7085 18400 7105
rect 18420 7085 18430 7105
rect 18390 7055 18430 7085
rect 18390 7035 18400 7055
rect 18420 7035 18430 7055
rect 18390 7020 18430 7035
rect 18775 7115 18815 7130
rect 18775 7095 18785 7115
rect 18805 7095 18815 7115
rect 18775 7065 18815 7095
rect 18775 7045 18785 7065
rect 18805 7045 18815 7065
rect 12485 6995 12495 7015
rect 12515 6995 12525 7015
rect 18775 7015 18815 7045
rect 12485 6980 12525 6995
rect 18775 6995 18785 7015
rect 18805 6995 18815 7015
rect 18775 6980 18815 6995
rect 18830 7115 18870 7130
rect 18830 7095 18840 7115
rect 18860 7095 18870 7115
rect 18830 7065 18870 7095
rect 18830 7045 18840 7065
rect 18860 7045 18870 7065
rect 18830 7015 18870 7045
rect 18830 6995 18840 7015
rect 18860 6995 18870 7015
rect 18830 6980 18870 6995
rect 18885 7115 18925 7130
rect 18885 7095 18895 7115
rect 18915 7095 18925 7115
rect 18885 7065 18925 7095
rect 18885 7045 18895 7065
rect 18915 7045 18925 7065
rect 18885 7015 18925 7045
rect 18885 6995 18895 7015
rect 18915 6995 18925 7015
rect 18885 6980 18925 6995
rect 18940 7115 18980 7130
rect 18940 7095 18950 7115
rect 18970 7095 18980 7115
rect 18940 7065 18980 7095
rect 18940 7045 18950 7065
rect 18970 7045 18980 7065
rect 18940 7015 18980 7045
rect 18940 6995 18950 7015
rect 18970 6995 18980 7015
rect 18940 6980 18980 6995
rect 18995 7115 19035 7130
rect 18995 7095 19005 7115
rect 19025 7095 19035 7115
rect 18995 7065 19035 7095
rect 18995 7045 19005 7065
rect 19025 7045 19035 7065
rect 18995 7015 19035 7045
rect 18995 6995 19005 7015
rect 19025 6995 19035 7015
rect 18995 6980 19035 6995
rect 19050 7115 19090 7130
rect 19050 7095 19060 7115
rect 19080 7095 19090 7115
rect 19050 7065 19090 7095
rect 19050 7045 19060 7065
rect 19080 7045 19090 7065
rect 19050 7015 19090 7045
rect 19050 6995 19060 7015
rect 19080 6995 19090 7015
rect 19050 6980 19090 6995
rect 19105 7115 19145 7130
rect 19105 7095 19115 7115
rect 19135 7095 19145 7115
rect 19105 7065 19145 7095
rect 19105 7045 19115 7065
rect 19135 7045 19145 7065
rect 19105 7015 19145 7045
rect 19105 6995 19115 7015
rect 19135 6995 19145 7015
rect 19105 6980 19145 6995
rect 19160 7115 19200 7130
rect 19160 7095 19170 7115
rect 19190 7095 19200 7115
rect 19160 7065 19200 7095
rect 19160 7045 19170 7065
rect 19190 7045 19200 7065
rect 19160 7015 19200 7045
rect 19160 6995 19170 7015
rect 19190 6995 19200 7015
rect 19160 6980 19200 6995
rect 19215 7115 19255 7130
rect 19215 7095 19225 7115
rect 19245 7095 19255 7115
rect 19215 7065 19255 7095
rect 19215 7045 19225 7065
rect 19245 7045 19255 7065
rect 19215 7015 19255 7045
rect 19215 6995 19225 7015
rect 19245 6995 19255 7015
rect 19215 6980 19255 6995
rect 19270 7115 19310 7130
rect 19270 7095 19280 7115
rect 19300 7095 19310 7115
rect 19270 7065 19310 7095
rect 19270 7045 19280 7065
rect 19300 7045 19310 7065
rect 19270 7015 19310 7045
rect 19270 6995 19280 7015
rect 19300 6995 19310 7015
rect 19270 6980 19310 6995
rect 19325 7115 19365 7130
rect 19325 7095 19335 7115
rect 19355 7095 19365 7115
rect 19325 7065 19365 7095
rect 19325 7045 19335 7065
rect 19355 7045 19365 7065
rect 19325 7015 19365 7045
rect 19325 6995 19335 7015
rect 19355 6995 19365 7015
rect 19325 6980 19365 6995
rect 19380 7115 19420 7130
rect 19380 7095 19390 7115
rect 19410 7095 19420 7115
rect 19380 7065 19420 7095
rect 19380 7045 19390 7065
rect 19410 7045 19420 7065
rect 19380 7015 19420 7045
rect 19380 6995 19390 7015
rect 19410 6995 19420 7015
rect 19380 6980 19420 6995
rect 19435 7115 19475 7130
rect 19435 7095 19445 7115
rect 19465 7095 19475 7115
rect 19435 7065 19475 7095
rect 19435 7045 19445 7065
rect 19465 7045 19475 7065
rect 19435 7015 19475 7045
rect 19435 6995 19445 7015
rect 19465 6995 19475 7015
rect 19435 6980 19475 6995
rect 19490 7115 19530 7130
rect 19490 7095 19500 7115
rect 19520 7095 19530 7115
rect 19490 7065 19530 7095
rect 19490 7045 19500 7065
rect 19520 7045 19530 7065
rect 19490 7015 19530 7045
rect 19490 6995 19500 7015
rect 19520 6995 19530 7015
rect 19490 6980 19530 6995
rect 19545 7115 19585 7130
rect 19545 7095 19555 7115
rect 19575 7095 19585 7115
rect 19545 7065 19585 7095
rect 19545 7045 19555 7065
rect 19575 7045 19585 7065
rect 19545 7015 19585 7045
rect 19545 6995 19555 7015
rect 19575 6995 19585 7015
rect 19545 6980 19585 6995
rect 19600 7115 19640 7130
rect 19600 7095 19610 7115
rect 19630 7095 19640 7115
rect 19600 7065 19640 7095
rect 19600 7045 19610 7065
rect 19630 7045 19640 7065
rect 19600 7015 19640 7045
rect 19600 6995 19610 7015
rect 19630 6995 19640 7015
rect 19600 6980 19640 6995
rect 19655 7115 19695 7130
rect 19655 7095 19665 7115
rect 19685 7095 19695 7115
rect 19655 7065 19695 7095
rect 19655 7045 19665 7065
rect 19685 7045 19695 7065
rect 19655 7015 19695 7045
rect 19655 6995 19665 7015
rect 19685 6995 19695 7015
rect 19655 6980 19695 6995
rect 19710 7115 19750 7130
rect 19710 7095 19720 7115
rect 19740 7095 19750 7115
rect 19710 7065 19750 7095
rect 19710 7045 19720 7065
rect 19740 7045 19750 7065
rect 19710 7015 19750 7045
rect 19710 6995 19720 7015
rect 19740 6995 19750 7015
rect 19710 6980 19750 6995
rect 19765 7115 19805 7130
rect 19765 7095 19775 7115
rect 19795 7095 19805 7115
rect 19765 7065 19805 7095
rect 19765 7045 19775 7065
rect 19795 7045 19805 7065
rect 19765 7015 19805 7045
rect 19765 6995 19775 7015
rect 19795 6995 19805 7015
rect 19765 6980 19805 6995
rect 19820 7115 19860 7130
rect 19820 7095 19830 7115
rect 19850 7095 19860 7115
rect 19820 7065 19860 7095
rect 19820 7045 19830 7065
rect 19850 7045 19860 7065
rect 19820 7015 19860 7045
rect 19820 6995 19830 7015
rect 19850 6995 19860 7015
rect 19820 6980 19860 6995
rect 19875 7115 19915 7130
rect 19875 7095 19885 7115
rect 19905 7095 19915 7115
rect 19875 7065 19915 7095
rect 19875 7045 19885 7065
rect 19905 7045 19915 7065
rect 19875 7015 19915 7045
rect 19875 6995 19885 7015
rect 19905 6995 19915 7015
rect 19875 6980 19915 6995
rect 19930 7115 19970 7130
rect 19930 7095 19940 7115
rect 19960 7095 19970 7115
rect 19930 7065 19970 7095
rect 19930 7045 19940 7065
rect 19960 7045 19970 7065
rect 19930 7015 19970 7045
rect 19930 6995 19940 7015
rect 19960 6995 19970 7015
rect 19930 6980 19970 6995
rect 19985 7115 20025 7130
rect 19985 7095 19995 7115
rect 20015 7095 20025 7115
rect 19985 7065 20025 7095
rect 19985 7045 19995 7065
rect 20015 7045 20025 7065
rect 19985 7015 20025 7045
rect 20390 7105 20430 7135
rect 20390 7085 20400 7105
rect 20420 7085 20430 7105
rect 20390 7055 20430 7085
rect 20390 7035 20400 7055
rect 20420 7035 20430 7055
rect 20390 7020 20430 7035
rect 20445 7155 20485 7170
rect 20445 7135 20455 7155
rect 20475 7135 20485 7155
rect 20445 7105 20485 7135
rect 20445 7085 20455 7105
rect 20475 7085 20485 7105
rect 20445 7055 20485 7085
rect 20445 7035 20455 7055
rect 20475 7035 20485 7055
rect 20445 7020 20485 7035
rect 20500 7155 20540 7170
rect 20500 7135 20510 7155
rect 20530 7135 20540 7155
rect 20500 7105 20540 7135
rect 20500 7085 20510 7105
rect 20530 7085 20540 7105
rect 20500 7055 20540 7085
rect 20500 7035 20510 7055
rect 20530 7035 20540 7055
rect 20500 7020 20540 7035
rect 20555 7155 20595 7170
rect 20555 7135 20565 7155
rect 20585 7135 20595 7155
rect 20555 7105 20595 7135
rect 20555 7085 20565 7105
rect 20585 7085 20595 7105
rect 20555 7055 20595 7085
rect 20555 7035 20565 7055
rect 20585 7035 20595 7055
rect 20555 7020 20595 7035
rect 20610 7155 20650 7170
rect 20610 7135 20620 7155
rect 20640 7135 20650 7155
rect 20610 7105 20650 7135
rect 20610 7085 20620 7105
rect 20640 7085 20650 7105
rect 20610 7055 20650 7085
rect 20610 7035 20620 7055
rect 20640 7035 20650 7055
rect 20610 7020 20650 7035
rect 20665 7155 20705 7170
rect 20665 7135 20675 7155
rect 20695 7135 20705 7155
rect 20665 7105 20705 7135
rect 20665 7085 20675 7105
rect 20695 7085 20705 7105
rect 20665 7055 20705 7085
rect 20665 7035 20675 7055
rect 20695 7035 20705 7055
rect 20665 7020 20705 7035
rect 20720 7155 20760 7170
rect 20720 7135 20730 7155
rect 20750 7135 20760 7155
rect 20720 7105 20760 7135
rect 20720 7085 20730 7105
rect 20750 7085 20760 7105
rect 20720 7055 20760 7085
rect 20720 7035 20730 7055
rect 20750 7035 20760 7055
rect 20720 7020 20760 7035
rect 20775 7155 20815 7170
rect 20775 7135 20785 7155
rect 20805 7135 20815 7155
rect 20775 7105 20815 7135
rect 20775 7085 20785 7105
rect 20805 7085 20815 7105
rect 20775 7055 20815 7085
rect 20775 7035 20785 7055
rect 20805 7035 20815 7055
rect 20775 7020 20815 7035
rect 20830 7155 20870 7170
rect 20830 7135 20840 7155
rect 20860 7135 20870 7155
rect 20830 7105 20870 7135
rect 20830 7085 20840 7105
rect 20860 7085 20870 7105
rect 20830 7055 20870 7085
rect 20830 7035 20840 7055
rect 20860 7035 20870 7055
rect 20830 7020 20870 7035
rect 20885 7155 20925 7170
rect 20885 7135 20895 7155
rect 20915 7135 20925 7155
rect 20885 7105 20925 7135
rect 20885 7085 20895 7105
rect 20915 7085 20925 7105
rect 20885 7055 20925 7085
rect 20885 7035 20895 7055
rect 20915 7035 20925 7055
rect 20885 7020 20925 7035
rect 20940 7155 20980 7170
rect 20940 7135 20950 7155
rect 20970 7135 20980 7155
rect 20940 7105 20980 7135
rect 20940 7085 20950 7105
rect 20970 7085 20980 7105
rect 20940 7055 20980 7085
rect 20940 7035 20950 7055
rect 20970 7035 20980 7055
rect 20940 7020 20980 7035
rect 20995 7155 21035 7170
rect 20995 7135 21005 7155
rect 21025 7135 21035 7155
rect 20995 7105 21035 7135
rect 20995 7085 21005 7105
rect 21025 7085 21035 7105
rect 20995 7055 21035 7085
rect 20995 7035 21005 7055
rect 21025 7035 21035 7055
rect 20995 7020 21035 7035
rect 21050 7155 21090 7170
rect 21050 7135 21060 7155
rect 21080 7135 21090 7155
rect 21050 7105 21090 7135
rect 21050 7085 21060 7105
rect 21080 7085 21090 7105
rect 21050 7055 21090 7085
rect 21050 7035 21060 7055
rect 21080 7035 21090 7055
rect 21050 7020 21090 7035
rect 21105 7155 21145 7170
rect 21105 7135 21115 7155
rect 21135 7135 21145 7155
rect 21105 7105 21145 7135
rect 21105 7085 21115 7105
rect 21135 7085 21145 7105
rect 21105 7055 21145 7085
rect 21105 7035 21115 7055
rect 21135 7035 21145 7055
rect 21105 7020 21145 7035
rect 21160 7155 21200 7170
rect 21160 7135 21170 7155
rect 21190 7135 21200 7155
rect 21160 7105 21200 7135
rect 21160 7085 21170 7105
rect 21190 7085 21200 7105
rect 21160 7055 21200 7085
rect 21160 7035 21170 7055
rect 21190 7035 21200 7055
rect 21160 7020 21200 7035
rect 21215 7155 21255 7170
rect 21215 7135 21225 7155
rect 21245 7135 21255 7155
rect 21215 7105 21255 7135
rect 21215 7085 21225 7105
rect 21245 7085 21255 7105
rect 21215 7055 21255 7085
rect 21215 7035 21225 7055
rect 21245 7035 21255 7055
rect 21215 7020 21255 7035
rect 21270 7155 21310 7170
rect 21270 7135 21280 7155
rect 21300 7135 21310 7155
rect 21270 7105 21310 7135
rect 21270 7085 21280 7105
rect 21300 7085 21310 7105
rect 21270 7055 21310 7085
rect 21270 7035 21280 7055
rect 21300 7035 21310 7055
rect 21270 7020 21310 7035
rect 21325 7155 21365 7170
rect 21325 7135 21335 7155
rect 21355 7135 21365 7155
rect 21325 7105 21365 7135
rect 21325 7085 21335 7105
rect 21355 7085 21365 7105
rect 21325 7055 21365 7085
rect 21325 7035 21335 7055
rect 21355 7035 21365 7055
rect 21325 7020 21365 7035
rect 21380 7155 21420 7170
rect 21380 7135 21390 7155
rect 21410 7135 21420 7155
rect 21380 7105 21420 7135
rect 21380 7085 21390 7105
rect 21410 7085 21420 7105
rect 21380 7055 21420 7085
rect 21380 7035 21390 7055
rect 21410 7035 21420 7055
rect 21380 7020 21420 7035
rect 21435 7155 21475 7170
rect 21435 7135 21445 7155
rect 21465 7135 21475 7155
rect 21435 7105 21475 7135
rect 21435 7085 21445 7105
rect 21465 7085 21475 7105
rect 21435 7055 21475 7085
rect 21435 7035 21445 7055
rect 21465 7035 21475 7055
rect 21435 7020 21475 7035
rect 21490 7155 21530 7170
rect 21490 7135 21500 7155
rect 21520 7135 21530 7155
rect 21490 7105 21530 7135
rect 21490 7085 21500 7105
rect 21520 7085 21530 7105
rect 21490 7055 21530 7085
rect 21490 7035 21500 7055
rect 21520 7035 21530 7055
rect 21490 7020 21530 7035
rect 21545 7155 21585 7170
rect 21545 7135 21555 7155
rect 21575 7135 21585 7155
rect 21545 7105 21585 7135
rect 21545 7085 21555 7105
rect 21575 7085 21585 7105
rect 21545 7055 21585 7085
rect 21545 7035 21555 7055
rect 21575 7035 21585 7055
rect 21545 7020 21585 7035
rect 21600 7155 21640 7170
rect 21600 7135 21610 7155
rect 21630 7135 21640 7155
rect 21600 7105 21640 7135
rect 21600 7085 21610 7105
rect 21630 7085 21640 7105
rect 21600 7055 21640 7085
rect 21600 7035 21610 7055
rect 21630 7035 21640 7055
rect 21600 7020 21640 7035
rect 19985 6995 19995 7015
rect 20015 6995 20025 7015
rect 19985 6980 20025 6995
rect 20490 6840 20530 6855
rect 20490 6820 20500 6840
rect 20520 6820 20530 6840
rect 20490 6790 20530 6820
rect 20490 6770 20500 6790
rect 20520 6770 20530 6790
rect 20490 6740 20530 6770
rect 20490 6720 20500 6740
rect 20520 6720 20530 6740
rect 20490 6705 20530 6720
rect 20545 6840 20585 6855
rect 20545 6820 20555 6840
rect 20575 6820 20585 6840
rect 20545 6790 20585 6820
rect 20545 6770 20555 6790
rect 20575 6770 20585 6790
rect 20545 6740 20585 6770
rect 20545 6720 20555 6740
rect 20575 6720 20585 6740
rect 20545 6705 20585 6720
rect 20600 6840 20640 6855
rect 20600 6820 20610 6840
rect 20630 6820 20640 6840
rect 20600 6790 20640 6820
rect 20600 6770 20610 6790
rect 20630 6770 20640 6790
rect 20600 6740 20640 6770
rect 20600 6720 20610 6740
rect 20630 6720 20640 6740
rect 20600 6705 20640 6720
rect 20655 6840 20695 6855
rect 20655 6820 20665 6840
rect 20685 6820 20695 6840
rect 20655 6790 20695 6820
rect 20655 6770 20665 6790
rect 20685 6770 20695 6790
rect 20655 6740 20695 6770
rect 20655 6720 20665 6740
rect 20685 6720 20695 6740
rect 20655 6705 20695 6720
rect 20710 6840 20750 6855
rect 20710 6820 20720 6840
rect 20740 6820 20750 6840
rect 20710 6790 20750 6820
rect 20710 6770 20720 6790
rect 20740 6770 20750 6790
rect 20710 6740 20750 6770
rect 20710 6720 20720 6740
rect 20740 6720 20750 6740
rect 20710 6705 20750 6720
rect 20765 6840 20805 6855
rect 20765 6820 20775 6840
rect 20795 6820 20805 6840
rect 20765 6790 20805 6820
rect 20765 6770 20775 6790
rect 20795 6770 20805 6790
rect 20765 6740 20805 6770
rect 20765 6720 20775 6740
rect 20795 6720 20805 6740
rect 20765 6705 20805 6720
rect 20820 6840 20860 6855
rect 20820 6820 20830 6840
rect 20850 6820 20860 6840
rect 20820 6790 20860 6820
rect 20820 6770 20830 6790
rect 20850 6770 20860 6790
rect 20820 6740 20860 6770
rect 20820 6720 20830 6740
rect 20850 6720 20860 6740
rect 20820 6705 20860 6720
rect 11030 6650 11070 6665
rect 11030 6630 11040 6650
rect 11060 6630 11070 6650
rect 11030 6600 11070 6630
rect 11030 6580 11040 6600
rect 11060 6580 11070 6600
rect 11030 6550 11070 6580
rect 11030 6530 11040 6550
rect 11060 6530 11070 6550
rect 11030 6515 11070 6530
rect 11085 6650 11125 6665
rect 11085 6630 11095 6650
rect 11115 6630 11125 6650
rect 11085 6600 11125 6630
rect 11085 6580 11095 6600
rect 11115 6580 11125 6600
rect 11085 6550 11125 6580
rect 11085 6530 11095 6550
rect 11115 6530 11125 6550
rect 11085 6515 11125 6530
rect 11140 6650 11180 6665
rect 11140 6630 11150 6650
rect 11170 6630 11180 6650
rect 11140 6600 11180 6630
rect 11140 6580 11150 6600
rect 11170 6580 11180 6600
rect 11140 6550 11180 6580
rect 11140 6530 11150 6550
rect 11170 6530 11180 6550
rect 11140 6515 11180 6530
rect 11195 6650 11235 6665
rect 11195 6630 11205 6650
rect 11225 6630 11235 6650
rect 11195 6600 11235 6630
rect 11195 6580 11205 6600
rect 11225 6580 11235 6600
rect 11195 6550 11235 6580
rect 11195 6530 11205 6550
rect 11225 6530 11235 6550
rect 11195 6515 11235 6530
rect 11250 6650 11290 6665
rect 11250 6630 11260 6650
rect 11280 6630 11290 6650
rect 11250 6600 11290 6630
rect 11250 6580 11260 6600
rect 11280 6580 11290 6600
rect 11250 6550 11290 6580
rect 11250 6530 11260 6550
rect 11280 6530 11290 6550
rect 11250 6515 11290 6530
rect 11305 6650 11345 6665
rect 11305 6630 11315 6650
rect 11335 6630 11345 6650
rect 11305 6600 11345 6630
rect 11305 6580 11315 6600
rect 11335 6580 11345 6600
rect 11305 6550 11345 6580
rect 11305 6530 11315 6550
rect 11335 6530 11345 6550
rect 11305 6515 11345 6530
rect 11360 6650 11400 6665
rect 11360 6630 11370 6650
rect 11390 6630 11400 6650
rect 11360 6600 11400 6630
rect 11360 6580 11370 6600
rect 11390 6580 11400 6600
rect 11360 6550 11400 6580
rect 11360 6530 11370 6550
rect 11390 6530 11400 6550
rect 11360 6515 11400 6530
rect 11415 6650 11455 6665
rect 11415 6630 11425 6650
rect 11445 6630 11455 6650
rect 11415 6600 11455 6630
rect 11415 6580 11425 6600
rect 11445 6580 11455 6600
rect 11415 6550 11455 6580
rect 11415 6530 11425 6550
rect 11445 6530 11455 6550
rect 11415 6515 11455 6530
rect 11470 6650 11510 6665
rect 11470 6630 11480 6650
rect 11500 6630 11510 6650
rect 11470 6600 11510 6630
rect 11470 6580 11480 6600
rect 11500 6580 11510 6600
rect 11470 6550 11510 6580
rect 11470 6530 11480 6550
rect 11500 6530 11510 6550
rect 11470 6515 11510 6530
rect 11525 6650 11565 6665
rect 11525 6630 11535 6650
rect 11555 6630 11565 6650
rect 11525 6600 11565 6630
rect 11525 6580 11535 6600
rect 11555 6580 11565 6600
rect 11525 6550 11565 6580
rect 11525 6530 11535 6550
rect 11555 6530 11565 6550
rect 11525 6515 11565 6530
rect 11580 6650 11620 6665
rect 11580 6630 11590 6650
rect 11610 6630 11620 6650
rect 11580 6600 11620 6630
rect 11580 6580 11590 6600
rect 11610 6580 11620 6600
rect 11580 6550 11620 6580
rect 11580 6530 11590 6550
rect 11610 6530 11620 6550
rect 11580 6515 11620 6530
rect 11635 6650 11675 6665
rect 11635 6630 11645 6650
rect 11665 6630 11675 6650
rect 11635 6600 11675 6630
rect 11635 6580 11645 6600
rect 11665 6580 11675 6600
rect 11635 6550 11675 6580
rect 11635 6530 11645 6550
rect 11665 6530 11675 6550
rect 11635 6515 11675 6530
rect 11690 6650 11730 6665
rect 11770 6650 11810 6665
rect 11690 6630 11700 6650
rect 11720 6630 11730 6650
rect 11770 6630 11780 6650
rect 11800 6630 11810 6650
rect 11690 6600 11730 6630
rect 11770 6600 11810 6630
rect 11690 6580 11700 6600
rect 11720 6580 11730 6600
rect 11770 6580 11780 6600
rect 11800 6580 11810 6600
rect 11690 6550 11730 6580
rect 11770 6550 11810 6580
rect 11690 6530 11700 6550
rect 11720 6530 11730 6550
rect 11770 6530 11780 6550
rect 11800 6530 11810 6550
rect 11690 6515 11730 6530
rect 11770 6515 11810 6530
rect 11825 6650 11865 6665
rect 11825 6630 11835 6650
rect 11855 6630 11865 6650
rect 11825 6600 11865 6630
rect 11825 6580 11835 6600
rect 11855 6580 11865 6600
rect 11825 6550 11865 6580
rect 11825 6530 11835 6550
rect 11855 6530 11865 6550
rect 11825 6515 11865 6530
rect 11880 6650 11920 6665
rect 11880 6630 11890 6650
rect 11910 6630 11920 6650
rect 11880 6600 11920 6630
rect 11880 6580 11890 6600
rect 11910 6580 11920 6600
rect 11880 6550 11920 6580
rect 11880 6530 11890 6550
rect 11910 6530 11920 6550
rect 11880 6515 11920 6530
rect 11935 6650 11975 6665
rect 11935 6630 11945 6650
rect 11965 6630 11975 6650
rect 11935 6600 11975 6630
rect 11935 6580 11945 6600
rect 11965 6580 11975 6600
rect 11935 6550 11975 6580
rect 11935 6530 11945 6550
rect 11965 6530 11975 6550
rect 11935 6515 11975 6530
rect 11990 6650 12030 6665
rect 12070 6650 12110 6665
rect 11990 6630 12000 6650
rect 12020 6630 12030 6650
rect 12070 6630 12080 6650
rect 12100 6630 12110 6650
rect 11990 6600 12030 6630
rect 12070 6600 12110 6630
rect 11990 6580 12000 6600
rect 12020 6580 12030 6600
rect 12070 6580 12080 6600
rect 12100 6580 12110 6600
rect 11990 6550 12030 6580
rect 12070 6550 12110 6580
rect 11990 6530 12000 6550
rect 12020 6530 12030 6550
rect 12070 6530 12080 6550
rect 12100 6530 12110 6550
rect 11990 6515 12030 6530
rect 12070 6515 12110 6530
rect 12125 6650 12165 6665
rect 12125 6630 12135 6650
rect 12155 6630 12165 6650
rect 12125 6600 12165 6630
rect 12125 6580 12135 6600
rect 12155 6580 12165 6600
rect 12125 6550 12165 6580
rect 12125 6530 12135 6550
rect 12155 6530 12165 6550
rect 12125 6515 12165 6530
rect 12180 6650 12220 6665
rect 12180 6630 12190 6650
rect 12210 6630 12220 6650
rect 12180 6600 12220 6630
rect 12180 6580 12190 6600
rect 12210 6580 12220 6600
rect 12180 6550 12220 6580
rect 12180 6530 12190 6550
rect 12210 6530 12220 6550
rect 12180 6515 12220 6530
rect 12235 6650 12275 6665
rect 12235 6630 12245 6650
rect 12265 6630 12275 6650
rect 12235 6600 12275 6630
rect 12235 6580 12245 6600
rect 12265 6580 12275 6600
rect 12235 6550 12275 6580
rect 12235 6530 12245 6550
rect 12265 6530 12275 6550
rect 12235 6515 12275 6530
rect 12290 6650 12330 6665
rect 12290 6630 12300 6650
rect 12320 6630 12330 6650
rect 12290 6600 12330 6630
rect 12290 6580 12300 6600
rect 12320 6580 12330 6600
rect 12290 6550 12330 6580
rect 12290 6530 12300 6550
rect 12320 6530 12330 6550
rect 12290 6515 12330 6530
rect 12345 6650 12385 6665
rect 12345 6630 12355 6650
rect 12375 6630 12385 6650
rect 12345 6600 12385 6630
rect 12345 6580 12355 6600
rect 12375 6580 12385 6600
rect 12345 6550 12385 6580
rect 12345 6530 12355 6550
rect 12375 6530 12385 6550
rect 12345 6515 12385 6530
rect 12400 6650 12440 6665
rect 12400 6630 12410 6650
rect 12430 6630 12440 6650
rect 12400 6600 12440 6630
rect 12400 6580 12410 6600
rect 12430 6580 12440 6600
rect 12400 6550 12440 6580
rect 12400 6530 12410 6550
rect 12430 6530 12440 6550
rect 12400 6515 12440 6530
rect 12455 6650 12495 6665
rect 12455 6630 12465 6650
rect 12485 6630 12495 6650
rect 12455 6600 12495 6630
rect 12455 6580 12465 6600
rect 12485 6580 12495 6600
rect 12455 6550 12495 6580
rect 12455 6530 12465 6550
rect 12485 6530 12495 6550
rect 12455 6515 12495 6530
rect 12510 6650 12550 6665
rect 12510 6630 12520 6650
rect 12540 6630 12550 6650
rect 12510 6600 12550 6630
rect 12510 6580 12520 6600
rect 12540 6580 12550 6600
rect 12510 6550 12550 6580
rect 12510 6530 12520 6550
rect 12540 6530 12550 6550
rect 12510 6515 12550 6530
rect 12565 6650 12605 6665
rect 12565 6630 12575 6650
rect 12595 6630 12605 6650
rect 12565 6600 12605 6630
rect 12565 6580 12575 6600
rect 12595 6580 12605 6600
rect 12565 6550 12605 6580
rect 12565 6530 12575 6550
rect 12595 6530 12605 6550
rect 12565 6515 12605 6530
rect 12620 6650 12660 6665
rect 12620 6630 12630 6650
rect 12650 6630 12660 6650
rect 12620 6600 12660 6630
rect 12620 6580 12630 6600
rect 12650 6580 12660 6600
rect 12620 6550 12660 6580
rect 12620 6530 12630 6550
rect 12650 6530 12660 6550
rect 12620 6515 12660 6530
rect 12675 6650 12715 6665
rect 12675 6630 12685 6650
rect 12705 6630 12715 6650
rect 12675 6600 12715 6630
rect 12675 6580 12685 6600
rect 12705 6580 12715 6600
rect 12675 6550 12715 6580
rect 12675 6530 12685 6550
rect 12705 6530 12715 6550
rect 12675 6515 12715 6530
rect 12730 6650 12770 6665
rect 12730 6630 12740 6650
rect 12760 6630 12770 6650
rect 12730 6600 12770 6630
rect 12730 6580 12740 6600
rect 12760 6580 12770 6600
rect 12730 6550 12770 6580
rect 12730 6530 12740 6550
rect 12760 6530 12770 6550
rect 12730 6515 12770 6530
rect 18530 6650 18570 6665
rect 18530 6630 18540 6650
rect 18560 6630 18570 6650
rect 18530 6600 18570 6630
rect 18530 6580 18540 6600
rect 18560 6580 18570 6600
rect 18530 6550 18570 6580
rect 18530 6530 18540 6550
rect 18560 6530 18570 6550
rect 18530 6515 18570 6530
rect 18585 6650 18625 6665
rect 18585 6630 18595 6650
rect 18615 6630 18625 6650
rect 18585 6600 18625 6630
rect 18585 6580 18595 6600
rect 18615 6580 18625 6600
rect 18585 6550 18625 6580
rect 18585 6530 18595 6550
rect 18615 6530 18625 6550
rect 18585 6515 18625 6530
rect 18640 6650 18680 6665
rect 18640 6630 18650 6650
rect 18670 6630 18680 6650
rect 18640 6600 18680 6630
rect 18640 6580 18650 6600
rect 18670 6580 18680 6600
rect 18640 6550 18680 6580
rect 18640 6530 18650 6550
rect 18670 6530 18680 6550
rect 18640 6515 18680 6530
rect 18695 6650 18735 6665
rect 18695 6630 18705 6650
rect 18725 6630 18735 6650
rect 18695 6600 18735 6630
rect 18695 6580 18705 6600
rect 18725 6580 18735 6600
rect 18695 6550 18735 6580
rect 18695 6530 18705 6550
rect 18725 6530 18735 6550
rect 18695 6515 18735 6530
rect 18750 6650 18790 6665
rect 18750 6630 18760 6650
rect 18780 6630 18790 6650
rect 18750 6600 18790 6630
rect 18750 6580 18760 6600
rect 18780 6580 18790 6600
rect 18750 6550 18790 6580
rect 18750 6530 18760 6550
rect 18780 6530 18790 6550
rect 18750 6515 18790 6530
rect 18805 6650 18845 6665
rect 18805 6630 18815 6650
rect 18835 6630 18845 6650
rect 18805 6600 18845 6630
rect 18805 6580 18815 6600
rect 18835 6580 18845 6600
rect 18805 6550 18845 6580
rect 18805 6530 18815 6550
rect 18835 6530 18845 6550
rect 18805 6515 18845 6530
rect 18860 6650 18900 6665
rect 18860 6630 18870 6650
rect 18890 6630 18900 6650
rect 18860 6600 18900 6630
rect 18860 6580 18870 6600
rect 18890 6580 18900 6600
rect 18860 6550 18900 6580
rect 18860 6530 18870 6550
rect 18890 6530 18900 6550
rect 18860 6515 18900 6530
rect 18915 6650 18955 6665
rect 18915 6630 18925 6650
rect 18945 6630 18955 6650
rect 18915 6600 18955 6630
rect 18915 6580 18925 6600
rect 18945 6580 18955 6600
rect 18915 6550 18955 6580
rect 18915 6530 18925 6550
rect 18945 6530 18955 6550
rect 18915 6515 18955 6530
rect 18970 6650 19010 6665
rect 18970 6630 18980 6650
rect 19000 6630 19010 6650
rect 18970 6600 19010 6630
rect 18970 6580 18980 6600
rect 19000 6580 19010 6600
rect 18970 6550 19010 6580
rect 18970 6530 18980 6550
rect 19000 6530 19010 6550
rect 18970 6515 19010 6530
rect 19025 6650 19065 6665
rect 19025 6630 19035 6650
rect 19055 6630 19065 6650
rect 19025 6600 19065 6630
rect 19025 6580 19035 6600
rect 19055 6580 19065 6600
rect 19025 6550 19065 6580
rect 19025 6530 19035 6550
rect 19055 6530 19065 6550
rect 19025 6515 19065 6530
rect 19080 6650 19120 6665
rect 19080 6630 19090 6650
rect 19110 6630 19120 6650
rect 19080 6600 19120 6630
rect 19080 6580 19090 6600
rect 19110 6580 19120 6600
rect 19080 6550 19120 6580
rect 19080 6530 19090 6550
rect 19110 6530 19120 6550
rect 19080 6515 19120 6530
rect 19135 6650 19175 6665
rect 19135 6630 19145 6650
rect 19165 6630 19175 6650
rect 19135 6600 19175 6630
rect 19135 6580 19145 6600
rect 19165 6580 19175 6600
rect 19135 6550 19175 6580
rect 19135 6530 19145 6550
rect 19165 6530 19175 6550
rect 19135 6515 19175 6530
rect 19190 6650 19230 6665
rect 19270 6650 19310 6665
rect 19190 6630 19200 6650
rect 19220 6630 19230 6650
rect 19270 6630 19280 6650
rect 19300 6630 19310 6650
rect 19190 6600 19230 6630
rect 19270 6600 19310 6630
rect 19190 6580 19200 6600
rect 19220 6580 19230 6600
rect 19270 6580 19280 6600
rect 19300 6580 19310 6600
rect 19190 6550 19230 6580
rect 19270 6550 19310 6580
rect 19190 6530 19200 6550
rect 19220 6530 19230 6550
rect 19270 6530 19280 6550
rect 19300 6530 19310 6550
rect 19190 6515 19230 6530
rect 19270 6515 19310 6530
rect 19325 6650 19365 6665
rect 19325 6630 19335 6650
rect 19355 6630 19365 6650
rect 19325 6600 19365 6630
rect 19325 6580 19335 6600
rect 19355 6580 19365 6600
rect 19325 6550 19365 6580
rect 19325 6530 19335 6550
rect 19355 6530 19365 6550
rect 19325 6515 19365 6530
rect 19380 6650 19420 6665
rect 19380 6630 19390 6650
rect 19410 6630 19420 6650
rect 19380 6600 19420 6630
rect 19380 6580 19390 6600
rect 19410 6580 19420 6600
rect 19380 6550 19420 6580
rect 19380 6530 19390 6550
rect 19410 6530 19420 6550
rect 19380 6515 19420 6530
rect 19435 6650 19475 6665
rect 19435 6630 19445 6650
rect 19465 6630 19475 6650
rect 19435 6600 19475 6630
rect 19435 6580 19445 6600
rect 19465 6580 19475 6600
rect 19435 6550 19475 6580
rect 19435 6530 19445 6550
rect 19465 6530 19475 6550
rect 19435 6515 19475 6530
rect 19490 6650 19530 6665
rect 19570 6650 19610 6665
rect 19490 6630 19500 6650
rect 19520 6630 19530 6650
rect 19570 6630 19580 6650
rect 19600 6630 19610 6650
rect 19490 6600 19530 6630
rect 19570 6600 19610 6630
rect 19490 6580 19500 6600
rect 19520 6580 19530 6600
rect 19570 6580 19580 6600
rect 19600 6580 19610 6600
rect 19490 6550 19530 6580
rect 19570 6550 19610 6580
rect 19490 6530 19500 6550
rect 19520 6530 19530 6550
rect 19570 6530 19580 6550
rect 19600 6530 19610 6550
rect 19490 6515 19530 6530
rect 19570 6515 19610 6530
rect 19625 6650 19665 6665
rect 19625 6630 19635 6650
rect 19655 6630 19665 6650
rect 19625 6600 19665 6630
rect 19625 6580 19635 6600
rect 19655 6580 19665 6600
rect 19625 6550 19665 6580
rect 19625 6530 19635 6550
rect 19655 6530 19665 6550
rect 19625 6515 19665 6530
rect 19680 6650 19720 6665
rect 19680 6630 19690 6650
rect 19710 6630 19720 6650
rect 19680 6600 19720 6630
rect 19680 6580 19690 6600
rect 19710 6580 19720 6600
rect 19680 6550 19720 6580
rect 19680 6530 19690 6550
rect 19710 6530 19720 6550
rect 19680 6515 19720 6530
rect 19735 6650 19775 6665
rect 19735 6630 19745 6650
rect 19765 6630 19775 6650
rect 19735 6600 19775 6630
rect 19735 6580 19745 6600
rect 19765 6580 19775 6600
rect 19735 6550 19775 6580
rect 19735 6530 19745 6550
rect 19765 6530 19775 6550
rect 19735 6515 19775 6530
rect 19790 6650 19830 6665
rect 19790 6630 19800 6650
rect 19820 6630 19830 6650
rect 19790 6600 19830 6630
rect 19790 6580 19800 6600
rect 19820 6580 19830 6600
rect 19790 6550 19830 6580
rect 19790 6530 19800 6550
rect 19820 6530 19830 6550
rect 19790 6515 19830 6530
rect 19845 6650 19885 6665
rect 19845 6630 19855 6650
rect 19875 6630 19885 6650
rect 19845 6600 19885 6630
rect 19845 6580 19855 6600
rect 19875 6580 19885 6600
rect 19845 6550 19885 6580
rect 19845 6530 19855 6550
rect 19875 6530 19885 6550
rect 19845 6515 19885 6530
rect 19900 6650 19940 6665
rect 19900 6630 19910 6650
rect 19930 6630 19940 6650
rect 19900 6600 19940 6630
rect 19900 6580 19910 6600
rect 19930 6580 19940 6600
rect 19900 6550 19940 6580
rect 19900 6530 19910 6550
rect 19930 6530 19940 6550
rect 19900 6515 19940 6530
rect 19955 6650 19995 6665
rect 19955 6630 19965 6650
rect 19985 6630 19995 6650
rect 19955 6600 19995 6630
rect 19955 6580 19965 6600
rect 19985 6580 19995 6600
rect 19955 6550 19995 6580
rect 19955 6530 19965 6550
rect 19985 6530 19995 6550
rect 19955 6515 19995 6530
rect 20010 6650 20050 6665
rect 20010 6630 20020 6650
rect 20040 6630 20050 6650
rect 20010 6600 20050 6630
rect 20010 6580 20020 6600
rect 20040 6580 20050 6600
rect 20010 6550 20050 6580
rect 20010 6530 20020 6550
rect 20040 6530 20050 6550
rect 20010 6515 20050 6530
rect 20065 6650 20105 6665
rect 20065 6630 20075 6650
rect 20095 6630 20105 6650
rect 20065 6600 20105 6630
rect 20065 6580 20075 6600
rect 20095 6580 20105 6600
rect 20065 6550 20105 6580
rect 20065 6530 20075 6550
rect 20095 6530 20105 6550
rect 20065 6515 20105 6530
rect 20120 6650 20160 6665
rect 20120 6630 20130 6650
rect 20150 6630 20160 6650
rect 20120 6600 20160 6630
rect 20120 6580 20130 6600
rect 20150 6580 20160 6600
rect 20120 6550 20160 6580
rect 20120 6530 20130 6550
rect 20150 6530 20160 6550
rect 20120 6515 20160 6530
rect 20175 6650 20215 6665
rect 20175 6630 20185 6650
rect 20205 6630 20215 6650
rect 20175 6600 20215 6630
rect 20175 6580 20185 6600
rect 20205 6580 20215 6600
rect 20175 6550 20215 6580
rect 20175 6530 20185 6550
rect 20205 6530 20215 6550
rect 20175 6515 20215 6530
rect 20230 6650 20270 6665
rect 20230 6630 20240 6650
rect 20260 6630 20270 6650
rect 20230 6600 20270 6630
rect 20230 6580 20240 6600
rect 20260 6580 20270 6600
rect 20230 6550 20270 6580
rect 20230 6530 20240 6550
rect 20260 6530 20270 6550
rect 20230 6515 20270 6530
rect 20395 6505 20435 6520
rect 20395 6485 20405 6505
rect 20425 6485 20435 6505
rect 20395 6455 20435 6485
rect 20395 6435 20405 6455
rect 20425 6435 20435 6455
rect 20395 6405 20435 6435
rect 20395 6385 20405 6405
rect 20425 6385 20435 6405
rect 20395 6370 20435 6385
rect 20450 6505 20490 6520
rect 20450 6485 20460 6505
rect 20480 6485 20490 6505
rect 20450 6455 20490 6485
rect 20450 6435 20460 6455
rect 20480 6435 20490 6455
rect 20450 6405 20490 6435
rect 20450 6385 20460 6405
rect 20480 6385 20490 6405
rect 20450 6370 20490 6385
rect 20505 6505 20545 6520
rect 20505 6485 20515 6505
rect 20535 6485 20545 6505
rect 20505 6455 20545 6485
rect 20505 6435 20515 6455
rect 20535 6435 20545 6455
rect 20505 6405 20545 6435
rect 20505 6385 20515 6405
rect 20535 6385 20545 6405
rect 20505 6370 20545 6385
rect 20560 6505 20600 6520
rect 20560 6485 20570 6505
rect 20590 6485 20600 6505
rect 20560 6455 20600 6485
rect 20560 6435 20570 6455
rect 20590 6435 20600 6455
rect 20560 6405 20600 6435
rect 20560 6385 20570 6405
rect 20590 6385 20600 6405
rect 20560 6370 20600 6385
rect 20615 6505 20655 6520
rect 20695 6505 20735 6520
rect 20615 6485 20625 6505
rect 20645 6485 20655 6505
rect 20695 6485 20705 6505
rect 20725 6485 20735 6505
rect 20615 6455 20655 6485
rect 20695 6455 20735 6485
rect 20615 6435 20625 6455
rect 20645 6435 20655 6455
rect 20695 6435 20705 6455
rect 20725 6435 20735 6455
rect 20615 6405 20655 6435
rect 20695 6405 20735 6435
rect 20615 6385 20625 6405
rect 20645 6385 20655 6405
rect 20695 6385 20705 6405
rect 20725 6385 20735 6405
rect 20615 6370 20655 6385
rect 20695 6370 20735 6385
rect 20750 6505 20790 6520
rect 20750 6485 20760 6505
rect 20780 6485 20790 6505
rect 20750 6455 20790 6485
rect 20750 6435 20760 6455
rect 20780 6435 20790 6455
rect 20750 6405 20790 6435
rect 20750 6385 20760 6405
rect 20780 6385 20790 6405
rect 20750 6370 20790 6385
rect 20805 6505 20845 6520
rect 20805 6485 20815 6505
rect 20835 6485 20845 6505
rect 20805 6455 20845 6485
rect 20805 6435 20815 6455
rect 20835 6435 20845 6455
rect 20805 6405 20845 6435
rect 20805 6385 20815 6405
rect 20835 6385 20845 6405
rect 20805 6370 20845 6385
rect 20860 6505 20900 6520
rect 20860 6485 20870 6505
rect 20890 6485 20900 6505
rect 20860 6455 20900 6485
rect 20860 6435 20870 6455
rect 20890 6435 20900 6455
rect 20860 6405 20900 6435
rect 20860 6385 20870 6405
rect 20890 6385 20900 6405
rect 20860 6370 20900 6385
rect 20915 6505 20955 6520
rect 20915 6485 20925 6505
rect 20945 6485 20955 6505
rect 20915 6455 20955 6485
rect 20915 6435 20925 6455
rect 20945 6435 20955 6455
rect 20915 6405 20955 6435
rect 20915 6385 20925 6405
rect 20945 6385 20955 6405
rect 20915 6370 20955 6385
rect 9665 6270 9705 6285
rect 9665 6250 9675 6270
rect 9695 6250 9705 6270
rect 9665 6225 9705 6250
rect 9665 6205 9675 6225
rect 9695 6205 9705 6225
rect 9665 6180 9705 6205
rect 9665 6160 9675 6180
rect 9695 6160 9705 6180
rect 9665 6130 9705 6160
rect 9665 6110 9675 6130
rect 9695 6110 9705 6130
rect 9665 6085 9705 6110
rect 9665 6065 9675 6085
rect 9695 6065 9705 6085
rect 9665 6040 9705 6065
rect 9665 6020 9675 6040
rect 9695 6020 9705 6040
rect 9665 6005 9705 6020
rect 9765 6270 9805 6285
rect 9765 6250 9775 6270
rect 9795 6250 9805 6270
rect 9765 6225 9805 6250
rect 9765 6205 9775 6225
rect 9795 6205 9805 6225
rect 9765 6180 9805 6205
rect 9765 6160 9775 6180
rect 9795 6160 9805 6180
rect 9765 6130 9805 6160
rect 9765 6110 9775 6130
rect 9795 6110 9805 6130
rect 9765 6085 9805 6110
rect 9765 6065 9775 6085
rect 9795 6065 9805 6085
rect 9765 6040 9805 6065
rect 9765 6020 9775 6040
rect 9795 6020 9805 6040
rect 9765 6005 9805 6020
rect 9865 6270 9905 6285
rect 9865 6250 9875 6270
rect 9895 6250 9905 6270
rect 9865 6225 9905 6250
rect 9865 6205 9875 6225
rect 9895 6205 9905 6225
rect 9865 6180 9905 6205
rect 9865 6160 9875 6180
rect 9895 6160 9905 6180
rect 9865 6130 9905 6160
rect 9865 6110 9875 6130
rect 9895 6110 9905 6130
rect 9865 6085 9905 6110
rect 9865 6065 9875 6085
rect 9895 6065 9905 6085
rect 9865 6040 9905 6065
rect 9865 6020 9875 6040
rect 9895 6020 9905 6040
rect 9865 6005 9905 6020
rect 9965 6270 10005 6285
rect 9965 6250 9975 6270
rect 9995 6250 10005 6270
rect 9965 6225 10005 6250
rect 9965 6205 9975 6225
rect 9995 6205 10005 6225
rect 9965 6180 10005 6205
rect 9965 6160 9975 6180
rect 9995 6160 10005 6180
rect 9965 6130 10005 6160
rect 9965 6110 9975 6130
rect 9995 6110 10005 6130
rect 9965 6085 10005 6110
rect 9965 6065 9975 6085
rect 9995 6065 10005 6085
rect 9965 6040 10005 6065
rect 9965 6020 9975 6040
rect 9995 6020 10005 6040
rect 9965 6005 10005 6020
rect 10065 6270 10105 6285
rect 10065 6250 10075 6270
rect 10095 6250 10105 6270
rect 10065 6225 10105 6250
rect 10065 6205 10075 6225
rect 10095 6205 10105 6225
rect 10065 6180 10105 6205
rect 10065 6160 10075 6180
rect 10095 6160 10105 6180
rect 10065 6130 10105 6160
rect 10065 6110 10075 6130
rect 10095 6110 10105 6130
rect 10065 6085 10105 6110
rect 10065 6065 10075 6085
rect 10095 6065 10105 6085
rect 10065 6040 10105 6065
rect 10065 6020 10075 6040
rect 10095 6020 10105 6040
rect 10065 6005 10105 6020
rect 10165 6270 10205 6285
rect 10165 6250 10175 6270
rect 10195 6250 10205 6270
rect 10165 6225 10205 6250
rect 10165 6205 10175 6225
rect 10195 6205 10205 6225
rect 10165 6180 10205 6205
rect 10165 6160 10175 6180
rect 10195 6160 10205 6180
rect 10165 6130 10205 6160
rect 10165 6110 10175 6130
rect 10195 6110 10205 6130
rect 10165 6085 10205 6110
rect 10165 6065 10175 6085
rect 10195 6065 10205 6085
rect 10165 6040 10205 6065
rect 10165 6020 10175 6040
rect 10195 6020 10205 6040
rect 10165 6005 10205 6020
rect 10265 6270 10305 6285
rect 10265 6250 10275 6270
rect 10295 6250 10305 6270
rect 10265 6225 10305 6250
rect 10265 6205 10275 6225
rect 10295 6205 10305 6225
rect 10265 6180 10305 6205
rect 10265 6160 10275 6180
rect 10295 6160 10305 6180
rect 10265 6130 10305 6160
rect 10265 6110 10275 6130
rect 10295 6110 10305 6130
rect 10265 6085 10305 6110
rect 10265 6065 10275 6085
rect 10295 6065 10305 6085
rect 10265 6040 10305 6065
rect 10265 6020 10275 6040
rect 10295 6020 10305 6040
rect 10265 6005 10305 6020
rect 10365 6270 10405 6285
rect 10365 6250 10375 6270
rect 10395 6250 10405 6270
rect 10365 6225 10405 6250
rect 10365 6205 10375 6225
rect 10395 6205 10405 6225
rect 10365 6180 10405 6205
rect 10365 6160 10375 6180
rect 10395 6160 10405 6180
rect 10365 6130 10405 6160
rect 10365 6110 10375 6130
rect 10395 6110 10405 6130
rect 10365 6085 10405 6110
rect 10365 6065 10375 6085
rect 10395 6065 10405 6085
rect 10365 6040 10405 6065
rect 10365 6020 10375 6040
rect 10395 6020 10405 6040
rect 10365 6005 10405 6020
rect 10465 6270 10505 6285
rect 10465 6250 10475 6270
rect 10495 6250 10505 6270
rect 10465 6225 10505 6250
rect 10465 6205 10475 6225
rect 10495 6205 10505 6225
rect 10465 6180 10505 6205
rect 10465 6160 10475 6180
rect 10495 6160 10505 6180
rect 10465 6130 10505 6160
rect 10465 6110 10475 6130
rect 10495 6110 10505 6130
rect 10465 6085 10505 6110
rect 10465 6065 10475 6085
rect 10495 6065 10505 6085
rect 10465 6040 10505 6065
rect 10465 6020 10475 6040
rect 10495 6020 10505 6040
rect 10465 6005 10505 6020
rect 10565 6270 10605 6285
rect 10565 6250 10575 6270
rect 10595 6250 10605 6270
rect 10565 6225 10605 6250
rect 10565 6205 10575 6225
rect 10595 6205 10605 6225
rect 10565 6180 10605 6205
rect 10565 6160 10575 6180
rect 10595 6160 10605 6180
rect 10565 6130 10605 6160
rect 10565 6110 10575 6130
rect 10595 6110 10605 6130
rect 10565 6085 10605 6110
rect 10565 6065 10575 6085
rect 10595 6065 10605 6085
rect 10565 6040 10605 6065
rect 10565 6020 10575 6040
rect 10595 6020 10605 6040
rect 10565 6005 10605 6020
rect 10665 6270 10705 6285
rect 10665 6250 10675 6270
rect 10695 6250 10705 6270
rect 10665 6225 10705 6250
rect 10665 6205 10675 6225
rect 10695 6205 10705 6225
rect 10665 6180 10705 6205
rect 10665 6160 10675 6180
rect 10695 6160 10705 6180
rect 10665 6130 10705 6160
rect 10665 6110 10675 6130
rect 10695 6110 10705 6130
rect 10665 6085 10705 6110
rect 10665 6065 10675 6085
rect 10695 6065 10705 6085
rect 10665 6040 10705 6065
rect 10665 6020 10675 6040
rect 10695 6020 10705 6040
rect 10665 6005 10705 6020
rect 10765 6270 10805 6285
rect 10765 6250 10775 6270
rect 10795 6250 10805 6270
rect 10765 6225 10805 6250
rect 10765 6205 10775 6225
rect 10795 6205 10805 6225
rect 10765 6180 10805 6205
rect 10765 6160 10775 6180
rect 10795 6160 10805 6180
rect 10765 6130 10805 6160
rect 10765 6110 10775 6130
rect 10795 6110 10805 6130
rect 10765 6085 10805 6110
rect 10765 6065 10775 6085
rect 10795 6065 10805 6085
rect 10765 6040 10805 6065
rect 10765 6020 10775 6040
rect 10795 6020 10805 6040
rect 10765 6005 10805 6020
rect 10865 6270 10905 6285
rect 10865 6250 10875 6270
rect 10895 6250 10905 6270
rect 12895 6270 12935 6285
rect 10865 6225 10905 6250
rect 10865 6205 10875 6225
rect 10895 6205 10905 6225
rect 10865 6180 10905 6205
rect 12895 6250 12905 6270
rect 12925 6250 12935 6270
rect 12895 6225 12935 6250
rect 12895 6205 12905 6225
rect 12925 6205 12935 6225
rect 10865 6160 10875 6180
rect 10895 6160 10905 6180
rect 10865 6130 10905 6160
rect 10865 6110 10875 6130
rect 10895 6110 10905 6130
rect 10865 6085 10905 6110
rect 10865 6065 10875 6085
rect 10895 6065 10905 6085
rect 10865 6040 10905 6065
rect 10865 6020 10875 6040
rect 10895 6020 10905 6040
rect 10865 6005 10905 6020
rect 11205 6170 11245 6185
rect 11205 6150 11215 6170
rect 11235 6150 11245 6170
rect 11205 6120 11245 6150
rect 11205 6100 11215 6120
rect 11235 6100 11245 6120
rect 11205 6070 11245 6100
rect 11205 6050 11215 6070
rect 11235 6050 11245 6070
rect 11205 6020 11245 6050
rect 11205 6000 11215 6020
rect 11235 6000 11245 6020
rect 11205 5970 11245 6000
rect 11205 5950 11215 5970
rect 11235 5950 11245 5970
rect 11205 5935 11245 5950
rect 11260 6170 11300 6185
rect 11260 6150 11270 6170
rect 11290 6150 11300 6170
rect 11260 6120 11300 6150
rect 11260 6100 11270 6120
rect 11290 6100 11300 6120
rect 11260 6070 11300 6100
rect 11260 6050 11270 6070
rect 11290 6050 11300 6070
rect 11260 6020 11300 6050
rect 11260 6000 11270 6020
rect 11290 6000 11300 6020
rect 11260 5970 11300 6000
rect 11260 5950 11270 5970
rect 11290 5950 11300 5970
rect 11260 5935 11300 5950
rect 11315 6170 11355 6185
rect 11315 6150 11325 6170
rect 11345 6150 11355 6170
rect 11315 6120 11355 6150
rect 11315 6100 11325 6120
rect 11345 6100 11355 6120
rect 11315 6070 11355 6100
rect 11315 6050 11325 6070
rect 11345 6050 11355 6070
rect 11315 6020 11355 6050
rect 11315 6000 11325 6020
rect 11345 6000 11355 6020
rect 11315 5970 11355 6000
rect 11315 5950 11325 5970
rect 11345 5950 11355 5970
rect 11315 5935 11355 5950
rect 11370 6170 11410 6185
rect 11370 6150 11380 6170
rect 11400 6150 11410 6170
rect 11370 6120 11410 6150
rect 11370 6100 11380 6120
rect 11400 6100 11410 6120
rect 11370 6070 11410 6100
rect 11370 6050 11380 6070
rect 11400 6050 11410 6070
rect 11370 6020 11410 6050
rect 11370 6000 11380 6020
rect 11400 6000 11410 6020
rect 11370 5970 11410 6000
rect 11370 5950 11380 5970
rect 11400 5950 11410 5970
rect 11370 5935 11410 5950
rect 11425 6170 11465 6185
rect 11425 6150 11435 6170
rect 11455 6150 11465 6170
rect 11425 6120 11465 6150
rect 11425 6100 11435 6120
rect 11455 6100 11465 6120
rect 11425 6070 11465 6100
rect 11425 6050 11435 6070
rect 11455 6050 11465 6070
rect 11425 6020 11465 6050
rect 11425 6000 11435 6020
rect 11455 6000 11465 6020
rect 11425 5970 11465 6000
rect 11425 5950 11435 5970
rect 11455 5950 11465 5970
rect 11425 5935 11465 5950
rect 11480 6170 11520 6185
rect 11480 6150 11490 6170
rect 11510 6150 11520 6170
rect 11480 6120 11520 6150
rect 11480 6100 11490 6120
rect 11510 6100 11520 6120
rect 11480 6070 11520 6100
rect 11480 6050 11490 6070
rect 11510 6050 11520 6070
rect 11480 6020 11520 6050
rect 11480 6000 11490 6020
rect 11510 6000 11520 6020
rect 11480 5970 11520 6000
rect 11480 5950 11490 5970
rect 11510 5950 11520 5970
rect 11480 5935 11520 5950
rect 11535 6170 11575 6185
rect 11535 6150 11545 6170
rect 11565 6150 11575 6170
rect 11535 6120 11575 6150
rect 11535 6100 11545 6120
rect 11565 6100 11575 6120
rect 11535 6070 11575 6100
rect 11535 6050 11545 6070
rect 11565 6050 11575 6070
rect 11535 6020 11575 6050
rect 11535 6000 11545 6020
rect 11565 6000 11575 6020
rect 11535 5970 11575 6000
rect 11535 5950 11545 5970
rect 11565 5950 11575 5970
rect 11535 5935 11575 5950
rect 11590 6170 11630 6185
rect 11590 6150 11600 6170
rect 11620 6150 11630 6170
rect 11590 6120 11630 6150
rect 11590 6100 11600 6120
rect 11620 6100 11630 6120
rect 11590 6070 11630 6100
rect 11590 6050 11600 6070
rect 11620 6050 11630 6070
rect 11590 6020 11630 6050
rect 11590 6000 11600 6020
rect 11620 6000 11630 6020
rect 11590 5970 11630 6000
rect 11590 5950 11600 5970
rect 11620 5950 11630 5970
rect 11590 5935 11630 5950
rect 11645 6170 11685 6185
rect 11645 6150 11655 6170
rect 11675 6150 11685 6170
rect 11645 6120 11685 6150
rect 11645 6100 11655 6120
rect 11675 6100 11685 6120
rect 11645 6070 11685 6100
rect 11645 6050 11655 6070
rect 11675 6050 11685 6070
rect 11645 6020 11685 6050
rect 11645 6000 11655 6020
rect 11675 6000 11685 6020
rect 11645 5970 11685 6000
rect 11645 5950 11655 5970
rect 11675 5950 11685 5970
rect 11645 5935 11685 5950
rect 11700 6170 11740 6185
rect 11700 6150 11710 6170
rect 11730 6150 11740 6170
rect 11700 6120 11740 6150
rect 11700 6100 11710 6120
rect 11730 6100 11740 6120
rect 11700 6070 11740 6100
rect 11700 6050 11710 6070
rect 11730 6050 11740 6070
rect 11700 6020 11740 6050
rect 11700 6000 11710 6020
rect 11730 6000 11740 6020
rect 11700 5970 11740 6000
rect 11700 5950 11710 5970
rect 11730 5950 11740 5970
rect 11700 5935 11740 5950
rect 11755 6170 11795 6185
rect 11755 6150 11765 6170
rect 11785 6150 11795 6170
rect 11755 6120 11795 6150
rect 11755 6100 11765 6120
rect 11785 6100 11795 6120
rect 11755 6070 11795 6100
rect 11755 6050 11765 6070
rect 11785 6050 11795 6070
rect 11755 6020 11795 6050
rect 11755 6000 11765 6020
rect 11785 6000 11795 6020
rect 11755 5970 11795 6000
rect 11755 5950 11765 5970
rect 11785 5950 11795 5970
rect 11755 5935 11795 5950
rect 11810 6170 11850 6185
rect 11810 6150 11820 6170
rect 11840 6150 11850 6170
rect 11810 6120 11850 6150
rect 11810 6100 11820 6120
rect 11840 6100 11850 6120
rect 11810 6070 11850 6100
rect 11810 6050 11820 6070
rect 11840 6050 11850 6070
rect 11810 6020 11850 6050
rect 11810 6000 11820 6020
rect 11840 6000 11850 6020
rect 11810 5970 11850 6000
rect 11810 5950 11820 5970
rect 11840 5950 11850 5970
rect 11810 5935 11850 5950
rect 11865 6170 11905 6185
rect 11865 6150 11875 6170
rect 11895 6150 11905 6170
rect 11865 6120 11905 6150
rect 11865 6100 11875 6120
rect 11895 6100 11905 6120
rect 11865 6070 11905 6100
rect 11865 6050 11875 6070
rect 11895 6050 11905 6070
rect 11865 6020 11905 6050
rect 11865 6000 11875 6020
rect 11895 6000 11905 6020
rect 11865 5970 11905 6000
rect 11865 5950 11875 5970
rect 11895 5950 11905 5970
rect 11865 5935 11905 5950
rect 11920 6170 11960 6185
rect 11920 6150 11930 6170
rect 11950 6150 11960 6170
rect 11920 6120 11960 6150
rect 11920 6100 11930 6120
rect 11950 6100 11960 6120
rect 11920 6070 11960 6100
rect 11920 6050 11930 6070
rect 11950 6050 11960 6070
rect 11920 6020 11960 6050
rect 11920 6000 11930 6020
rect 11950 6000 11960 6020
rect 11920 5970 11960 6000
rect 11920 5950 11930 5970
rect 11950 5950 11960 5970
rect 11920 5935 11960 5950
rect 11975 6170 12015 6185
rect 11975 6150 11985 6170
rect 12005 6150 12015 6170
rect 11975 6120 12015 6150
rect 11975 6100 11985 6120
rect 12005 6100 12015 6120
rect 11975 6070 12015 6100
rect 11975 6050 11985 6070
rect 12005 6050 12015 6070
rect 11975 6020 12015 6050
rect 11975 6000 11985 6020
rect 12005 6000 12015 6020
rect 11975 5970 12015 6000
rect 11975 5950 11985 5970
rect 12005 5950 12015 5970
rect 11975 5935 12015 5950
rect 12030 6170 12070 6185
rect 12030 6150 12040 6170
rect 12060 6150 12070 6170
rect 12030 6120 12070 6150
rect 12030 6100 12040 6120
rect 12060 6100 12070 6120
rect 12030 6070 12070 6100
rect 12030 6050 12040 6070
rect 12060 6050 12070 6070
rect 12030 6020 12070 6050
rect 12030 6000 12040 6020
rect 12060 6000 12070 6020
rect 12030 5970 12070 6000
rect 12030 5950 12040 5970
rect 12060 5950 12070 5970
rect 12030 5935 12070 5950
rect 12085 6170 12125 6185
rect 12085 6150 12095 6170
rect 12115 6150 12125 6170
rect 12085 6120 12125 6150
rect 12085 6100 12095 6120
rect 12115 6100 12125 6120
rect 12085 6070 12125 6100
rect 12085 6050 12095 6070
rect 12115 6050 12125 6070
rect 12085 6020 12125 6050
rect 12085 6000 12095 6020
rect 12115 6000 12125 6020
rect 12085 5970 12125 6000
rect 12085 5950 12095 5970
rect 12115 5950 12125 5970
rect 12085 5935 12125 5950
rect 12140 6170 12180 6185
rect 12140 6150 12150 6170
rect 12170 6150 12180 6170
rect 12140 6120 12180 6150
rect 12140 6100 12150 6120
rect 12170 6100 12180 6120
rect 12140 6070 12180 6100
rect 12140 6050 12150 6070
rect 12170 6050 12180 6070
rect 12140 6020 12180 6050
rect 12140 6000 12150 6020
rect 12170 6000 12180 6020
rect 12140 5970 12180 6000
rect 12140 5950 12150 5970
rect 12170 5950 12180 5970
rect 12140 5935 12180 5950
rect 12195 6170 12235 6185
rect 12195 6150 12205 6170
rect 12225 6150 12235 6170
rect 12195 6120 12235 6150
rect 12195 6100 12205 6120
rect 12225 6100 12235 6120
rect 12195 6070 12235 6100
rect 12195 6050 12205 6070
rect 12225 6050 12235 6070
rect 12195 6020 12235 6050
rect 12195 6000 12205 6020
rect 12225 6000 12235 6020
rect 12195 5970 12235 6000
rect 12195 5950 12205 5970
rect 12225 5950 12235 5970
rect 12195 5935 12235 5950
rect 12250 6170 12290 6185
rect 12250 6150 12260 6170
rect 12280 6150 12290 6170
rect 12250 6120 12290 6150
rect 12250 6100 12260 6120
rect 12280 6100 12290 6120
rect 12250 6070 12290 6100
rect 12250 6050 12260 6070
rect 12280 6050 12290 6070
rect 12250 6020 12290 6050
rect 12250 6000 12260 6020
rect 12280 6000 12290 6020
rect 12250 5970 12290 6000
rect 12250 5950 12260 5970
rect 12280 5950 12290 5970
rect 12250 5935 12290 5950
rect 12305 6170 12345 6185
rect 12305 6150 12315 6170
rect 12335 6150 12345 6170
rect 12305 6120 12345 6150
rect 12305 6100 12315 6120
rect 12335 6100 12345 6120
rect 12305 6070 12345 6100
rect 12305 6050 12315 6070
rect 12335 6050 12345 6070
rect 12305 6020 12345 6050
rect 12305 6000 12315 6020
rect 12335 6000 12345 6020
rect 12305 5970 12345 6000
rect 12305 5950 12315 5970
rect 12335 5950 12345 5970
rect 12305 5935 12345 5950
rect 12360 6170 12400 6185
rect 12360 6150 12370 6170
rect 12390 6150 12400 6170
rect 12360 6120 12400 6150
rect 12360 6100 12370 6120
rect 12390 6100 12400 6120
rect 12360 6070 12400 6100
rect 12360 6050 12370 6070
rect 12390 6050 12400 6070
rect 12360 6020 12400 6050
rect 12360 6000 12370 6020
rect 12390 6000 12400 6020
rect 12360 5970 12400 6000
rect 12360 5950 12370 5970
rect 12390 5950 12400 5970
rect 12360 5935 12400 5950
rect 12415 6170 12455 6185
rect 12415 6150 12425 6170
rect 12445 6150 12455 6170
rect 12415 6120 12455 6150
rect 12415 6100 12425 6120
rect 12445 6100 12455 6120
rect 12415 6070 12455 6100
rect 12415 6050 12425 6070
rect 12445 6050 12455 6070
rect 12415 6020 12455 6050
rect 12415 6000 12425 6020
rect 12445 6000 12455 6020
rect 12415 5970 12455 6000
rect 12415 5950 12425 5970
rect 12445 5950 12455 5970
rect 12415 5935 12455 5950
rect 12470 6170 12510 6185
rect 12470 6150 12480 6170
rect 12500 6150 12510 6170
rect 12470 6120 12510 6150
rect 12470 6100 12480 6120
rect 12500 6100 12510 6120
rect 12470 6070 12510 6100
rect 12470 6050 12480 6070
rect 12500 6050 12510 6070
rect 12470 6020 12510 6050
rect 12470 6000 12480 6020
rect 12500 6000 12510 6020
rect 12470 5970 12510 6000
rect 12470 5950 12480 5970
rect 12500 5950 12510 5970
rect 12470 5935 12510 5950
rect 12525 6170 12565 6185
rect 12525 6150 12535 6170
rect 12555 6150 12565 6170
rect 12525 6120 12565 6150
rect 12525 6100 12535 6120
rect 12555 6100 12565 6120
rect 12525 6070 12565 6100
rect 12525 6050 12535 6070
rect 12555 6050 12565 6070
rect 12525 6020 12565 6050
rect 12525 6000 12535 6020
rect 12555 6000 12565 6020
rect 12525 5970 12565 6000
rect 12525 5950 12535 5970
rect 12555 5950 12565 5970
rect 12525 5935 12565 5950
rect 12580 6170 12620 6185
rect 12580 6150 12590 6170
rect 12610 6150 12620 6170
rect 12580 6120 12620 6150
rect 12580 6100 12590 6120
rect 12610 6100 12620 6120
rect 12580 6070 12620 6100
rect 12580 6050 12590 6070
rect 12610 6050 12620 6070
rect 12580 6020 12620 6050
rect 12580 6000 12590 6020
rect 12610 6000 12620 6020
rect 12895 6180 12935 6205
rect 12895 6160 12905 6180
rect 12925 6160 12935 6180
rect 12895 6130 12935 6160
rect 12895 6110 12905 6130
rect 12925 6110 12935 6130
rect 12895 6085 12935 6110
rect 12895 6065 12905 6085
rect 12925 6065 12935 6085
rect 12895 6040 12935 6065
rect 12895 6020 12905 6040
rect 12925 6020 12935 6040
rect 12895 6005 12935 6020
rect 12995 6270 13035 6285
rect 12995 6250 13005 6270
rect 13025 6250 13035 6270
rect 12995 6225 13035 6250
rect 12995 6205 13005 6225
rect 13025 6205 13035 6225
rect 12995 6180 13035 6205
rect 12995 6160 13005 6180
rect 13025 6160 13035 6180
rect 12995 6130 13035 6160
rect 12995 6110 13005 6130
rect 13025 6110 13035 6130
rect 12995 6085 13035 6110
rect 12995 6065 13005 6085
rect 13025 6065 13035 6085
rect 12995 6040 13035 6065
rect 12995 6020 13005 6040
rect 13025 6020 13035 6040
rect 12995 6005 13035 6020
rect 13095 6270 13135 6285
rect 13095 6250 13105 6270
rect 13125 6250 13135 6270
rect 13095 6225 13135 6250
rect 13095 6205 13105 6225
rect 13125 6205 13135 6225
rect 13095 6180 13135 6205
rect 13095 6160 13105 6180
rect 13125 6160 13135 6180
rect 13095 6130 13135 6160
rect 13095 6110 13105 6130
rect 13125 6110 13135 6130
rect 13095 6085 13135 6110
rect 13095 6065 13105 6085
rect 13125 6065 13135 6085
rect 13095 6040 13135 6065
rect 13095 6020 13105 6040
rect 13125 6020 13135 6040
rect 13095 6005 13135 6020
rect 13195 6270 13235 6285
rect 13195 6250 13205 6270
rect 13225 6250 13235 6270
rect 13195 6225 13235 6250
rect 13195 6205 13205 6225
rect 13225 6205 13235 6225
rect 13195 6180 13235 6205
rect 13195 6160 13205 6180
rect 13225 6160 13235 6180
rect 13195 6130 13235 6160
rect 13195 6110 13205 6130
rect 13225 6110 13235 6130
rect 13195 6085 13235 6110
rect 13195 6065 13205 6085
rect 13225 6065 13235 6085
rect 13195 6040 13235 6065
rect 13195 6020 13205 6040
rect 13225 6020 13235 6040
rect 13195 6005 13235 6020
rect 13295 6270 13335 6285
rect 13295 6250 13305 6270
rect 13325 6250 13335 6270
rect 13295 6225 13335 6250
rect 13295 6205 13305 6225
rect 13325 6205 13335 6225
rect 13295 6180 13335 6205
rect 13295 6160 13305 6180
rect 13325 6160 13335 6180
rect 13295 6130 13335 6160
rect 13295 6110 13305 6130
rect 13325 6110 13335 6130
rect 13295 6085 13335 6110
rect 13295 6065 13305 6085
rect 13325 6065 13335 6085
rect 13295 6040 13335 6065
rect 13295 6020 13305 6040
rect 13325 6020 13335 6040
rect 13295 6005 13335 6020
rect 13395 6270 13435 6285
rect 13395 6250 13405 6270
rect 13425 6250 13435 6270
rect 13395 6225 13435 6250
rect 13395 6205 13405 6225
rect 13425 6205 13435 6225
rect 13395 6180 13435 6205
rect 13395 6160 13405 6180
rect 13425 6160 13435 6180
rect 13395 6130 13435 6160
rect 13395 6110 13405 6130
rect 13425 6110 13435 6130
rect 13395 6085 13435 6110
rect 13395 6065 13405 6085
rect 13425 6065 13435 6085
rect 13395 6040 13435 6065
rect 13395 6020 13405 6040
rect 13425 6020 13435 6040
rect 13395 6005 13435 6020
rect 13495 6270 13535 6285
rect 13495 6250 13505 6270
rect 13525 6250 13535 6270
rect 13495 6225 13535 6250
rect 13495 6205 13505 6225
rect 13525 6205 13535 6225
rect 13495 6180 13535 6205
rect 13495 6160 13505 6180
rect 13525 6160 13535 6180
rect 13495 6130 13535 6160
rect 13495 6110 13505 6130
rect 13525 6110 13535 6130
rect 13495 6085 13535 6110
rect 13495 6065 13505 6085
rect 13525 6065 13535 6085
rect 13495 6040 13535 6065
rect 13495 6020 13505 6040
rect 13525 6020 13535 6040
rect 13495 6005 13535 6020
rect 13595 6270 13635 6285
rect 13595 6250 13605 6270
rect 13625 6250 13635 6270
rect 13595 6225 13635 6250
rect 13595 6205 13605 6225
rect 13625 6205 13635 6225
rect 13595 6180 13635 6205
rect 13595 6160 13605 6180
rect 13625 6160 13635 6180
rect 13595 6130 13635 6160
rect 13595 6110 13605 6130
rect 13625 6110 13635 6130
rect 13595 6085 13635 6110
rect 13595 6065 13605 6085
rect 13625 6065 13635 6085
rect 13595 6040 13635 6065
rect 13595 6020 13605 6040
rect 13625 6020 13635 6040
rect 13595 6005 13635 6020
rect 13695 6270 13735 6285
rect 13695 6250 13705 6270
rect 13725 6250 13735 6270
rect 13695 6225 13735 6250
rect 13695 6205 13705 6225
rect 13725 6205 13735 6225
rect 13695 6180 13735 6205
rect 13695 6160 13705 6180
rect 13725 6160 13735 6180
rect 13695 6130 13735 6160
rect 13695 6110 13705 6130
rect 13725 6110 13735 6130
rect 13695 6085 13735 6110
rect 13695 6065 13705 6085
rect 13725 6065 13735 6085
rect 13695 6040 13735 6065
rect 13695 6020 13705 6040
rect 13725 6020 13735 6040
rect 13695 6005 13735 6020
rect 13795 6270 13835 6285
rect 13795 6250 13805 6270
rect 13825 6250 13835 6270
rect 13795 6225 13835 6250
rect 13795 6205 13805 6225
rect 13825 6205 13835 6225
rect 13795 6180 13835 6205
rect 13795 6160 13805 6180
rect 13825 6160 13835 6180
rect 13795 6130 13835 6160
rect 13795 6110 13805 6130
rect 13825 6110 13835 6130
rect 13795 6085 13835 6110
rect 13795 6065 13805 6085
rect 13825 6065 13835 6085
rect 13795 6040 13835 6065
rect 13795 6020 13805 6040
rect 13825 6020 13835 6040
rect 13795 6005 13835 6020
rect 13895 6270 13935 6285
rect 13895 6250 13905 6270
rect 13925 6250 13935 6270
rect 13895 6225 13935 6250
rect 13895 6205 13905 6225
rect 13925 6205 13935 6225
rect 13895 6180 13935 6205
rect 13895 6160 13905 6180
rect 13925 6160 13935 6180
rect 13895 6130 13935 6160
rect 13895 6110 13905 6130
rect 13925 6110 13935 6130
rect 13895 6085 13935 6110
rect 13895 6065 13905 6085
rect 13925 6065 13935 6085
rect 13895 6040 13935 6065
rect 13895 6020 13905 6040
rect 13925 6020 13935 6040
rect 13895 6005 13935 6020
rect 13995 6270 14035 6285
rect 13995 6250 14005 6270
rect 14025 6250 14035 6270
rect 13995 6225 14035 6250
rect 13995 6205 14005 6225
rect 14025 6205 14035 6225
rect 13995 6180 14035 6205
rect 13995 6160 14005 6180
rect 14025 6160 14035 6180
rect 13995 6130 14035 6160
rect 13995 6110 14005 6130
rect 14025 6110 14035 6130
rect 13995 6085 14035 6110
rect 13995 6065 14005 6085
rect 14025 6065 14035 6085
rect 13995 6040 14035 6065
rect 13995 6020 14005 6040
rect 14025 6020 14035 6040
rect 13995 6005 14035 6020
rect 14095 6270 14135 6285
rect 14095 6250 14105 6270
rect 14125 6250 14135 6270
rect 14095 6225 14135 6250
rect 14095 6205 14105 6225
rect 14125 6205 14135 6225
rect 14095 6180 14135 6205
rect 14095 6160 14105 6180
rect 14125 6160 14135 6180
rect 14095 6130 14135 6160
rect 14095 6110 14105 6130
rect 14125 6110 14135 6130
rect 14095 6085 14135 6110
rect 14095 6065 14105 6085
rect 14125 6065 14135 6085
rect 14095 6040 14135 6065
rect 14095 6020 14105 6040
rect 14125 6020 14135 6040
rect 14095 6005 14135 6020
rect 18705 6210 18745 6225
rect 18705 6190 18715 6210
rect 18735 6190 18745 6210
rect 18705 6160 18745 6190
rect 18705 6140 18715 6160
rect 18735 6140 18745 6160
rect 18705 6110 18745 6140
rect 18705 6090 18715 6110
rect 18735 6090 18745 6110
rect 18705 6060 18745 6090
rect 18705 6040 18715 6060
rect 18735 6040 18745 6060
rect 18705 6010 18745 6040
rect 12580 5970 12620 6000
rect 12580 5950 12590 5970
rect 12610 5950 12620 5970
rect 18705 5990 18715 6010
rect 18735 5990 18745 6010
rect 18705 5975 18745 5990
rect 18760 6210 18800 6225
rect 18760 6190 18770 6210
rect 18790 6190 18800 6210
rect 18760 6160 18800 6190
rect 18760 6140 18770 6160
rect 18790 6140 18800 6160
rect 18760 6110 18800 6140
rect 18760 6090 18770 6110
rect 18790 6090 18800 6110
rect 18760 6060 18800 6090
rect 18760 6040 18770 6060
rect 18790 6040 18800 6060
rect 18760 6010 18800 6040
rect 18760 5990 18770 6010
rect 18790 5990 18800 6010
rect 18760 5975 18800 5990
rect 18815 6210 18855 6225
rect 18815 6190 18825 6210
rect 18845 6190 18855 6210
rect 18815 6160 18855 6190
rect 18815 6140 18825 6160
rect 18845 6140 18855 6160
rect 18815 6110 18855 6140
rect 18815 6090 18825 6110
rect 18845 6090 18855 6110
rect 18815 6060 18855 6090
rect 18815 6040 18825 6060
rect 18845 6040 18855 6060
rect 18815 6010 18855 6040
rect 18815 5990 18825 6010
rect 18845 5990 18855 6010
rect 18815 5975 18855 5990
rect 18870 6210 18910 6225
rect 18870 6190 18880 6210
rect 18900 6190 18910 6210
rect 18870 6160 18910 6190
rect 18870 6140 18880 6160
rect 18900 6140 18910 6160
rect 18870 6110 18910 6140
rect 18870 6090 18880 6110
rect 18900 6090 18910 6110
rect 18870 6060 18910 6090
rect 18870 6040 18880 6060
rect 18900 6040 18910 6060
rect 18870 6010 18910 6040
rect 18870 5990 18880 6010
rect 18900 5990 18910 6010
rect 18870 5975 18910 5990
rect 18925 6210 18965 6225
rect 18925 6190 18935 6210
rect 18955 6190 18965 6210
rect 18925 6160 18965 6190
rect 18925 6140 18935 6160
rect 18955 6140 18965 6160
rect 18925 6110 18965 6140
rect 18925 6090 18935 6110
rect 18955 6090 18965 6110
rect 18925 6060 18965 6090
rect 18925 6040 18935 6060
rect 18955 6040 18965 6060
rect 18925 6010 18965 6040
rect 18925 5990 18935 6010
rect 18955 5990 18965 6010
rect 18925 5975 18965 5990
rect 18980 6210 19020 6225
rect 18980 6190 18990 6210
rect 19010 6190 19020 6210
rect 18980 6160 19020 6190
rect 18980 6140 18990 6160
rect 19010 6140 19020 6160
rect 18980 6110 19020 6140
rect 18980 6090 18990 6110
rect 19010 6090 19020 6110
rect 18980 6060 19020 6090
rect 18980 6040 18990 6060
rect 19010 6040 19020 6060
rect 18980 6010 19020 6040
rect 18980 5990 18990 6010
rect 19010 5990 19020 6010
rect 18980 5975 19020 5990
rect 19035 6210 19075 6225
rect 19035 6190 19045 6210
rect 19065 6190 19075 6210
rect 19035 6160 19075 6190
rect 19035 6140 19045 6160
rect 19065 6140 19075 6160
rect 19035 6110 19075 6140
rect 19035 6090 19045 6110
rect 19065 6090 19075 6110
rect 19035 6060 19075 6090
rect 19035 6040 19045 6060
rect 19065 6040 19075 6060
rect 19035 6010 19075 6040
rect 19035 5990 19045 6010
rect 19065 5990 19075 6010
rect 19035 5975 19075 5990
rect 19090 6210 19130 6225
rect 19090 6190 19100 6210
rect 19120 6190 19130 6210
rect 19090 6160 19130 6190
rect 19090 6140 19100 6160
rect 19120 6140 19130 6160
rect 19090 6110 19130 6140
rect 19090 6090 19100 6110
rect 19120 6090 19130 6110
rect 19090 6060 19130 6090
rect 19090 6040 19100 6060
rect 19120 6040 19130 6060
rect 19090 6010 19130 6040
rect 19090 5990 19100 6010
rect 19120 5990 19130 6010
rect 19090 5975 19130 5990
rect 19145 6210 19185 6225
rect 19145 6190 19155 6210
rect 19175 6190 19185 6210
rect 19145 6160 19185 6190
rect 19145 6140 19155 6160
rect 19175 6140 19185 6160
rect 19145 6110 19185 6140
rect 19145 6090 19155 6110
rect 19175 6090 19185 6110
rect 19145 6060 19185 6090
rect 19145 6040 19155 6060
rect 19175 6040 19185 6060
rect 19145 6010 19185 6040
rect 19145 5990 19155 6010
rect 19175 5990 19185 6010
rect 19145 5975 19185 5990
rect 19200 6210 19240 6225
rect 19200 6190 19210 6210
rect 19230 6190 19240 6210
rect 19200 6160 19240 6190
rect 19200 6140 19210 6160
rect 19230 6140 19240 6160
rect 19200 6110 19240 6140
rect 19200 6090 19210 6110
rect 19230 6090 19240 6110
rect 19200 6060 19240 6090
rect 19200 6040 19210 6060
rect 19230 6040 19240 6060
rect 19200 6010 19240 6040
rect 19200 5990 19210 6010
rect 19230 5990 19240 6010
rect 19200 5975 19240 5990
rect 19255 6210 19295 6225
rect 19255 6190 19265 6210
rect 19285 6190 19295 6210
rect 19255 6160 19295 6190
rect 19255 6140 19265 6160
rect 19285 6140 19295 6160
rect 19255 6110 19295 6140
rect 19255 6090 19265 6110
rect 19285 6090 19295 6110
rect 19255 6060 19295 6090
rect 19255 6040 19265 6060
rect 19285 6040 19295 6060
rect 19255 6010 19295 6040
rect 19255 5990 19265 6010
rect 19285 5990 19295 6010
rect 19255 5975 19295 5990
rect 19310 6210 19350 6225
rect 19310 6190 19320 6210
rect 19340 6190 19350 6210
rect 19310 6160 19350 6190
rect 19310 6140 19320 6160
rect 19340 6140 19350 6160
rect 19310 6110 19350 6140
rect 19310 6090 19320 6110
rect 19340 6090 19350 6110
rect 19310 6060 19350 6090
rect 19310 6040 19320 6060
rect 19340 6040 19350 6060
rect 19310 6010 19350 6040
rect 19310 5990 19320 6010
rect 19340 5990 19350 6010
rect 19310 5975 19350 5990
rect 19365 6210 19405 6225
rect 19365 6190 19375 6210
rect 19395 6190 19405 6210
rect 19365 6160 19405 6190
rect 19365 6140 19375 6160
rect 19395 6140 19405 6160
rect 19365 6110 19405 6140
rect 19365 6090 19375 6110
rect 19395 6090 19405 6110
rect 19365 6060 19405 6090
rect 19365 6040 19375 6060
rect 19395 6040 19405 6060
rect 19365 6010 19405 6040
rect 19365 5990 19375 6010
rect 19395 5990 19405 6010
rect 19365 5975 19405 5990
rect 19420 6210 19460 6225
rect 19420 6190 19430 6210
rect 19450 6190 19460 6210
rect 19420 6160 19460 6190
rect 19420 6140 19430 6160
rect 19450 6140 19460 6160
rect 19420 6110 19460 6140
rect 19420 6090 19430 6110
rect 19450 6090 19460 6110
rect 19420 6060 19460 6090
rect 19420 6040 19430 6060
rect 19450 6040 19460 6060
rect 19420 6010 19460 6040
rect 19420 5990 19430 6010
rect 19450 5990 19460 6010
rect 19420 5975 19460 5990
rect 19475 6210 19515 6225
rect 19475 6190 19485 6210
rect 19505 6190 19515 6210
rect 19475 6160 19515 6190
rect 19475 6140 19485 6160
rect 19505 6140 19515 6160
rect 19475 6110 19515 6140
rect 19475 6090 19485 6110
rect 19505 6090 19515 6110
rect 19475 6060 19515 6090
rect 19475 6040 19485 6060
rect 19505 6040 19515 6060
rect 19475 6010 19515 6040
rect 19475 5990 19485 6010
rect 19505 5990 19515 6010
rect 19475 5975 19515 5990
rect 19530 6210 19570 6225
rect 19530 6190 19540 6210
rect 19560 6190 19570 6210
rect 19530 6160 19570 6190
rect 19530 6140 19540 6160
rect 19560 6140 19570 6160
rect 19530 6110 19570 6140
rect 19530 6090 19540 6110
rect 19560 6090 19570 6110
rect 19530 6060 19570 6090
rect 19530 6040 19540 6060
rect 19560 6040 19570 6060
rect 19530 6010 19570 6040
rect 19530 5990 19540 6010
rect 19560 5990 19570 6010
rect 19530 5975 19570 5990
rect 19585 6210 19625 6225
rect 19585 6190 19595 6210
rect 19615 6190 19625 6210
rect 19585 6160 19625 6190
rect 19585 6140 19595 6160
rect 19615 6140 19625 6160
rect 19585 6110 19625 6140
rect 19585 6090 19595 6110
rect 19615 6090 19625 6110
rect 19585 6060 19625 6090
rect 19585 6040 19595 6060
rect 19615 6040 19625 6060
rect 19585 6010 19625 6040
rect 19585 5990 19595 6010
rect 19615 5990 19625 6010
rect 19585 5975 19625 5990
rect 19640 6210 19680 6225
rect 19640 6190 19650 6210
rect 19670 6190 19680 6210
rect 19640 6160 19680 6190
rect 19640 6140 19650 6160
rect 19670 6140 19680 6160
rect 19640 6110 19680 6140
rect 19640 6090 19650 6110
rect 19670 6090 19680 6110
rect 19640 6060 19680 6090
rect 19640 6040 19650 6060
rect 19670 6040 19680 6060
rect 19640 6010 19680 6040
rect 19640 5990 19650 6010
rect 19670 5990 19680 6010
rect 19640 5975 19680 5990
rect 19695 6210 19735 6225
rect 19695 6190 19705 6210
rect 19725 6190 19735 6210
rect 19695 6160 19735 6190
rect 19695 6140 19705 6160
rect 19725 6140 19735 6160
rect 19695 6110 19735 6140
rect 19695 6090 19705 6110
rect 19725 6090 19735 6110
rect 19695 6060 19735 6090
rect 19695 6040 19705 6060
rect 19725 6040 19735 6060
rect 19695 6010 19735 6040
rect 19695 5990 19705 6010
rect 19725 5990 19735 6010
rect 19695 5975 19735 5990
rect 19750 6210 19790 6225
rect 19750 6190 19760 6210
rect 19780 6190 19790 6210
rect 19750 6160 19790 6190
rect 19750 6140 19760 6160
rect 19780 6140 19790 6160
rect 19750 6110 19790 6140
rect 19750 6090 19760 6110
rect 19780 6090 19790 6110
rect 19750 6060 19790 6090
rect 19750 6040 19760 6060
rect 19780 6040 19790 6060
rect 19750 6010 19790 6040
rect 19750 5990 19760 6010
rect 19780 5990 19790 6010
rect 19750 5975 19790 5990
rect 19805 6210 19845 6225
rect 19805 6190 19815 6210
rect 19835 6190 19845 6210
rect 19805 6160 19845 6190
rect 19805 6140 19815 6160
rect 19835 6140 19845 6160
rect 19805 6110 19845 6140
rect 19805 6090 19815 6110
rect 19835 6090 19845 6110
rect 19805 6060 19845 6090
rect 19805 6040 19815 6060
rect 19835 6040 19845 6060
rect 19805 6010 19845 6040
rect 19805 5990 19815 6010
rect 19835 5990 19845 6010
rect 19805 5975 19845 5990
rect 19860 6210 19900 6225
rect 19860 6190 19870 6210
rect 19890 6190 19900 6210
rect 19860 6160 19900 6190
rect 19860 6140 19870 6160
rect 19890 6140 19900 6160
rect 19860 6110 19900 6140
rect 19860 6090 19870 6110
rect 19890 6090 19900 6110
rect 19860 6060 19900 6090
rect 19860 6040 19870 6060
rect 19890 6040 19900 6060
rect 19860 6010 19900 6040
rect 19860 5990 19870 6010
rect 19890 5990 19900 6010
rect 19860 5975 19900 5990
rect 19915 6210 19955 6225
rect 19915 6190 19925 6210
rect 19945 6190 19955 6210
rect 19915 6160 19955 6190
rect 19915 6140 19925 6160
rect 19945 6140 19955 6160
rect 19915 6110 19955 6140
rect 19915 6090 19925 6110
rect 19945 6090 19955 6110
rect 19915 6060 19955 6090
rect 19915 6040 19925 6060
rect 19945 6040 19955 6060
rect 19915 6010 19955 6040
rect 19915 5990 19925 6010
rect 19945 5990 19955 6010
rect 19915 5975 19955 5990
rect 19970 6210 20010 6225
rect 19970 6190 19980 6210
rect 20000 6190 20010 6210
rect 19970 6160 20010 6190
rect 19970 6140 19980 6160
rect 20000 6140 20010 6160
rect 19970 6110 20010 6140
rect 19970 6090 19980 6110
rect 20000 6090 20010 6110
rect 19970 6060 20010 6090
rect 19970 6040 19980 6060
rect 20000 6040 20010 6060
rect 19970 6010 20010 6040
rect 19970 5990 19980 6010
rect 20000 5990 20010 6010
rect 19970 5975 20010 5990
rect 20025 6210 20065 6225
rect 20025 6190 20035 6210
rect 20055 6190 20065 6210
rect 20025 6160 20065 6190
rect 20025 6140 20035 6160
rect 20055 6140 20065 6160
rect 20025 6110 20065 6140
rect 20025 6090 20035 6110
rect 20055 6090 20065 6110
rect 20025 6060 20065 6090
rect 20025 6040 20035 6060
rect 20055 6040 20065 6060
rect 20025 6010 20065 6040
rect 20025 5990 20035 6010
rect 20055 5990 20065 6010
rect 20025 5975 20065 5990
rect 20080 6210 20120 6225
rect 20080 6190 20090 6210
rect 20110 6190 20120 6210
rect 20080 6160 20120 6190
rect 20080 6140 20090 6160
rect 20110 6140 20120 6160
rect 20080 6110 20120 6140
rect 20080 6090 20090 6110
rect 20110 6090 20120 6110
rect 20080 6060 20120 6090
rect 20080 6040 20090 6060
rect 20110 6040 20120 6060
rect 20080 6010 20120 6040
rect 20545 6165 20585 6180
rect 20545 6145 20555 6165
rect 20575 6145 20585 6165
rect 20545 6115 20585 6145
rect 20545 6095 20555 6115
rect 20575 6095 20585 6115
rect 20545 6065 20585 6095
rect 20545 6045 20555 6065
rect 20575 6045 20585 6065
rect 20545 6030 20585 6045
rect 20600 6165 20640 6180
rect 20600 6145 20610 6165
rect 20630 6145 20640 6165
rect 20600 6115 20640 6145
rect 20600 6095 20610 6115
rect 20630 6095 20640 6115
rect 20600 6065 20640 6095
rect 20600 6045 20610 6065
rect 20630 6045 20640 6065
rect 20600 6030 20640 6045
rect 20655 6165 20695 6180
rect 20655 6145 20665 6165
rect 20685 6145 20695 6165
rect 20655 6115 20695 6145
rect 20655 6095 20665 6115
rect 20685 6095 20695 6115
rect 20655 6065 20695 6095
rect 20655 6045 20665 6065
rect 20685 6045 20695 6065
rect 20655 6030 20695 6045
rect 20710 6165 20750 6180
rect 20710 6145 20720 6165
rect 20740 6145 20750 6165
rect 20710 6115 20750 6145
rect 20710 6095 20720 6115
rect 20740 6095 20750 6115
rect 20710 6065 20750 6095
rect 20710 6045 20720 6065
rect 20740 6045 20750 6065
rect 20710 6030 20750 6045
rect 20765 6165 20805 6180
rect 20765 6145 20775 6165
rect 20795 6145 20805 6165
rect 20765 6115 20805 6145
rect 20765 6095 20775 6115
rect 20795 6095 20805 6115
rect 20765 6065 20805 6095
rect 20765 6045 20775 6065
rect 20795 6045 20805 6065
rect 20765 6030 20805 6045
rect 20080 5990 20090 6010
rect 20110 5990 20120 6010
rect 20080 5975 20120 5990
rect 12580 5935 12620 5950
rect 11240 4375 11280 4403
rect 11240 4355 11250 4375
rect 11270 4355 11280 4375
rect 11240 4340 11280 4355
rect 11300 4380 11340 4403
rect 11300 4360 11310 4380
rect 11330 4360 11340 4380
rect 11300 4340 11340 4360
rect 11360 4380 11400 4403
rect 11360 4360 11370 4380
rect 11390 4360 11400 4380
rect 11360 4340 11400 4360
rect 11420 4375 11460 4403
rect 11420 4355 11430 4375
rect 11450 4355 11460 4375
rect 11420 4340 11460 4355
rect 11570 4390 11610 4420
rect 11570 4370 11580 4390
rect 11600 4370 11610 4390
rect 11570 4340 11610 4370
rect 11630 4390 11670 4420
rect 11630 4370 11640 4390
rect 11660 4370 11670 4390
rect 11630 4340 11670 4370
rect 11690 4390 11730 4420
rect 11690 4370 11700 4390
rect 11720 4370 11730 4390
rect 11690 4340 11730 4370
rect 11750 4390 11790 4420
rect 11750 4370 11760 4390
rect 11780 4370 11790 4390
rect 11750 4340 11790 4370
rect 11810 4390 11850 4420
rect 11810 4370 11820 4390
rect 11840 4370 11850 4390
rect 11810 4340 11850 4370
rect 11870 4390 11910 4420
rect 11870 4370 11880 4390
rect 11900 4370 11910 4390
rect 11870 4340 11910 4370
rect 11930 4390 11970 4420
rect 11930 4370 11940 4390
rect 11960 4370 11970 4390
rect 11930 4340 11970 4370
rect 12080 4375 12120 4395
rect 12080 4355 12090 4375
rect 12110 4355 12120 4375
rect 12080 4335 12120 4355
rect 12140 4375 12180 4395
rect 12140 4355 12150 4375
rect 12170 4355 12180 4375
rect 12140 4335 12180 4355
rect 12200 4375 12240 4395
rect 12200 4355 12210 4375
rect 12230 4355 12240 4375
rect 12200 4335 12240 4355
rect 12260 4375 12300 4395
rect 12260 4355 12270 4375
rect 12290 4355 12300 4375
rect 12260 4335 12300 4355
rect 12320 4375 12360 4395
rect 12320 4355 12330 4375
rect 12350 4355 12360 4375
rect 12320 4335 12360 4355
rect 12380 4375 12420 4395
rect 12380 4355 12390 4375
rect 12410 4355 12420 4375
rect 12380 4335 12420 4355
rect 12440 4375 12480 4395
rect 12440 4355 12450 4375
rect 12470 4355 12480 4375
rect 12440 4335 12480 4355
rect 12500 4375 12540 4395
rect 12500 4355 12510 4375
rect 12530 4355 12540 4375
rect 12500 4335 12540 4355
rect 12560 4375 12600 4395
rect 12560 4355 12570 4375
rect 12590 4355 12600 4375
rect 12560 4335 12600 4355
rect 11250 4140 11290 4155
rect 11250 4120 11260 4140
rect 11280 4120 11290 4140
rect 11250 4105 11290 4120
rect 11305 4140 11345 4155
rect 11305 4120 11315 4140
rect 11335 4120 11345 4140
rect 11305 4105 11345 4120
rect 11360 4140 11400 4155
rect 11360 4120 11370 4140
rect 11390 4120 11400 4140
rect 11360 4105 11400 4120
rect 11415 4140 11455 4155
rect 11415 4120 11425 4140
rect 11445 4120 11455 4140
rect 11415 4105 11455 4120
rect 11470 4140 11510 4155
rect 11470 4120 11480 4140
rect 11500 4120 11510 4140
rect 11470 4105 11510 4120
rect 11525 4140 11565 4155
rect 11525 4120 11535 4140
rect 11555 4120 11565 4140
rect 11525 4105 11565 4120
rect 11580 4140 11620 4155
rect 11580 4120 11590 4140
rect 11610 4120 11620 4140
rect 11580 4105 11620 4120
rect 11635 4140 11675 4155
rect 11635 4120 11645 4140
rect 11665 4120 11675 4140
rect 11635 4105 11675 4120
rect 11690 4140 11730 4155
rect 11690 4120 11700 4140
rect 11720 4120 11730 4140
rect 11690 4105 11730 4120
rect 11745 4140 11785 4155
rect 11745 4120 11755 4140
rect 11775 4120 11785 4140
rect 11745 4105 11785 4120
rect 11800 4140 11840 4155
rect 11800 4120 11810 4140
rect 11830 4120 11840 4140
rect 11800 4105 11840 4120
rect 11855 4140 11895 4155
rect 11855 4120 11865 4140
rect 11885 4120 11895 4140
rect 11855 4105 11895 4120
rect 11910 4140 11950 4155
rect 11910 4120 11920 4140
rect 11940 4120 11950 4140
rect 11910 4105 11950 4120
rect 11965 4140 12005 4155
rect 11965 4120 11975 4140
rect 11995 4120 12005 4140
rect 11965 4105 12005 4120
rect 12020 4140 12060 4155
rect 12020 4120 12030 4140
rect 12050 4120 12060 4140
rect 12020 4105 12060 4120
rect 12075 4140 12115 4155
rect 12075 4120 12085 4140
rect 12105 4120 12115 4140
rect 12075 4105 12115 4120
rect 12130 4140 12170 4155
rect 12130 4120 12140 4140
rect 12160 4120 12170 4140
rect 12130 4105 12170 4120
rect 12185 4140 12225 4155
rect 12185 4120 12195 4140
rect 12215 4120 12225 4140
rect 12185 4105 12225 4120
rect 12240 4140 12280 4155
rect 12240 4120 12250 4140
rect 12270 4120 12280 4140
rect 12240 4105 12280 4120
rect 12295 4140 12335 4155
rect 12295 4120 12305 4140
rect 12325 4120 12335 4140
rect 12295 4105 12335 4120
rect 12350 4140 12390 4155
rect 12350 4120 12360 4140
rect 12380 4120 12390 4140
rect 12350 4105 12390 4120
rect 12405 4140 12445 4155
rect 12405 4120 12415 4140
rect 12435 4120 12445 4140
rect 12405 4105 12445 4120
rect 12460 4140 12500 4155
rect 12460 4120 12470 4140
rect 12490 4120 12500 4140
rect 12460 4105 12500 4120
rect 11195 3835 11235 3850
rect 11195 3815 11205 3835
rect 11225 3815 11235 3835
rect 11195 3800 11235 3815
rect 11250 3835 11290 3850
rect 11250 3815 11260 3835
rect 11280 3815 11290 3835
rect 11250 3800 11290 3815
rect 11305 3835 11345 3850
rect 11305 3815 11315 3835
rect 11335 3815 11345 3835
rect 11305 3800 11345 3815
rect 11360 3835 11400 3850
rect 11360 3815 11370 3835
rect 11390 3815 11400 3835
rect 11360 3800 11400 3815
rect 11415 3835 11455 3850
rect 11415 3815 11425 3835
rect 11445 3815 11455 3835
rect 11415 3800 11455 3815
rect 11470 3835 11510 3850
rect 11470 3815 11480 3835
rect 11500 3815 11510 3835
rect 11470 3800 11510 3815
rect 11525 3835 11565 3850
rect 11525 3815 11535 3835
rect 11555 3815 11565 3835
rect 11525 3800 11565 3815
rect 11580 3835 11620 3850
rect 11580 3815 11590 3835
rect 11610 3815 11620 3835
rect 11580 3800 11620 3815
rect 11635 3835 11675 3850
rect 11635 3815 11645 3835
rect 11665 3815 11675 3835
rect 11635 3800 11675 3815
rect 11690 3835 11730 3850
rect 11690 3815 11700 3835
rect 11720 3815 11730 3835
rect 11690 3800 11730 3815
rect 11745 3835 11785 3850
rect 11745 3815 11755 3835
rect 11775 3815 11785 3835
rect 11745 3800 11785 3815
rect 11800 3835 11840 3850
rect 11800 3815 11810 3835
rect 11830 3815 11840 3835
rect 11800 3800 11840 3815
rect 11855 3835 11895 3850
rect 11935 3835 11975 3850
rect 11855 3815 11865 3835
rect 11885 3815 11895 3835
rect 11935 3815 11945 3835
rect 11965 3815 11975 3835
rect 11855 3800 11895 3815
rect 11935 3800 11975 3815
rect 11990 3835 12030 3850
rect 11990 3815 12000 3835
rect 12020 3815 12030 3835
rect 11990 3800 12030 3815
rect 12045 3835 12085 3850
rect 12045 3815 12055 3835
rect 12075 3815 12085 3835
rect 12045 3800 12085 3815
rect 12100 3835 12140 3850
rect 12100 3815 12110 3835
rect 12130 3815 12140 3835
rect 12100 3800 12140 3815
rect 12155 3835 12195 3850
rect 12155 3815 12165 3835
rect 12185 3815 12195 3835
rect 12155 3800 12195 3815
rect 12210 3835 12250 3850
rect 12210 3815 12220 3835
rect 12240 3815 12250 3835
rect 12210 3800 12250 3815
rect 12265 3835 12305 3850
rect 12265 3815 12275 3835
rect 12295 3815 12305 3835
rect 12265 3800 12305 3815
rect 12320 3835 12360 3850
rect 12320 3815 12330 3835
rect 12350 3815 12360 3835
rect 12320 3800 12360 3815
rect 12375 3835 12415 3850
rect 12375 3815 12385 3835
rect 12405 3815 12415 3835
rect 12375 3800 12415 3815
rect 12430 3835 12470 3850
rect 12430 3815 12440 3835
rect 12460 3815 12470 3835
rect 12430 3800 12470 3815
rect 12485 3835 12525 3850
rect 12485 3815 12495 3835
rect 12515 3815 12525 3835
rect 12485 3800 12525 3815
rect 12540 3835 12580 3850
rect 12540 3815 12550 3835
rect 12570 3815 12580 3835
rect 12540 3800 12580 3815
rect 12595 3835 12635 3850
rect 12595 3815 12605 3835
rect 12625 3815 12635 3835
rect 12595 3800 12635 3815
rect 10155 3570 10195 3585
rect 10155 3550 10165 3570
rect 10185 3550 10195 3570
rect 10155 3520 10195 3550
rect 10155 3500 10165 3520
rect 10185 3500 10195 3520
rect 10155 3470 10195 3500
rect 10155 3450 10165 3470
rect 10185 3450 10195 3470
rect 10155 3420 10195 3450
rect 10155 3400 10165 3420
rect 10185 3400 10195 3420
rect 10155 3370 10195 3400
rect 10155 3350 10165 3370
rect 10185 3350 10195 3370
rect 10155 3320 10195 3350
rect 10155 3300 10165 3320
rect 10185 3300 10195 3320
rect 10155 3270 10195 3300
rect 10155 3250 10165 3270
rect 10185 3250 10195 3270
rect 10155 3220 10195 3250
rect 10155 3200 10165 3220
rect 10185 3200 10195 3220
rect 10155 3170 10195 3200
rect 10155 3150 10165 3170
rect 10185 3150 10195 3170
rect 10155 3120 10195 3150
rect 10155 3100 10165 3120
rect 10185 3100 10195 3120
rect 10155 3070 10195 3100
rect 10155 3050 10165 3070
rect 10185 3050 10195 3070
rect 10155 3020 10195 3050
rect 10155 3000 10165 3020
rect 10185 3000 10195 3020
rect 10155 2985 10195 3000
rect 10210 3570 10250 3585
rect 10210 3550 10220 3570
rect 10240 3550 10250 3570
rect 10210 3520 10250 3550
rect 10210 3500 10220 3520
rect 10240 3500 10250 3520
rect 10210 3470 10250 3500
rect 10210 3450 10220 3470
rect 10240 3450 10250 3470
rect 10210 3420 10250 3450
rect 10210 3400 10220 3420
rect 10240 3400 10250 3420
rect 10210 3370 10250 3400
rect 10210 3350 10220 3370
rect 10240 3350 10250 3370
rect 10210 3320 10250 3350
rect 10210 3300 10220 3320
rect 10240 3300 10250 3320
rect 10210 3270 10250 3300
rect 10210 3250 10220 3270
rect 10240 3250 10250 3270
rect 10210 3220 10250 3250
rect 10210 3200 10220 3220
rect 10240 3200 10250 3220
rect 10210 3170 10250 3200
rect 10210 3150 10220 3170
rect 10240 3150 10250 3170
rect 10210 3120 10250 3150
rect 10210 3100 10220 3120
rect 10240 3100 10250 3120
rect 10210 3070 10250 3100
rect 10210 3050 10220 3070
rect 10240 3050 10250 3070
rect 10210 3020 10250 3050
rect 10210 3000 10220 3020
rect 10240 3000 10250 3020
rect 10210 2985 10250 3000
rect 10265 3570 10305 3585
rect 10265 3550 10275 3570
rect 10295 3550 10305 3570
rect 10265 3520 10305 3550
rect 10265 3500 10275 3520
rect 10295 3500 10305 3520
rect 10265 3470 10305 3500
rect 10265 3450 10275 3470
rect 10295 3450 10305 3470
rect 10265 3420 10305 3450
rect 10265 3400 10275 3420
rect 10295 3400 10305 3420
rect 10265 3370 10305 3400
rect 10265 3350 10275 3370
rect 10295 3350 10305 3370
rect 10265 3320 10305 3350
rect 10265 3300 10275 3320
rect 10295 3300 10305 3320
rect 10265 3270 10305 3300
rect 10265 3250 10275 3270
rect 10295 3250 10305 3270
rect 10265 3220 10305 3250
rect 10265 3200 10275 3220
rect 10295 3200 10305 3220
rect 10265 3170 10305 3200
rect 10265 3150 10275 3170
rect 10295 3150 10305 3170
rect 10265 3120 10305 3150
rect 10265 3100 10275 3120
rect 10295 3100 10305 3120
rect 10265 3070 10305 3100
rect 10265 3050 10275 3070
rect 10295 3050 10305 3070
rect 10265 3020 10305 3050
rect 10265 3000 10275 3020
rect 10295 3000 10305 3020
rect 10265 2985 10305 3000
rect 10320 3570 10360 3585
rect 10320 3550 10330 3570
rect 10350 3550 10360 3570
rect 10320 3520 10360 3550
rect 10320 3500 10330 3520
rect 10350 3500 10360 3520
rect 10320 3470 10360 3500
rect 10320 3450 10330 3470
rect 10350 3450 10360 3470
rect 10320 3420 10360 3450
rect 10320 3400 10330 3420
rect 10350 3400 10360 3420
rect 10320 3370 10360 3400
rect 10320 3350 10330 3370
rect 10350 3350 10360 3370
rect 10320 3320 10360 3350
rect 10320 3300 10330 3320
rect 10350 3300 10360 3320
rect 10320 3270 10360 3300
rect 10320 3250 10330 3270
rect 10350 3250 10360 3270
rect 10320 3220 10360 3250
rect 10320 3200 10330 3220
rect 10350 3200 10360 3220
rect 10320 3170 10360 3200
rect 10320 3150 10330 3170
rect 10350 3150 10360 3170
rect 10320 3120 10360 3150
rect 10320 3100 10330 3120
rect 10350 3100 10360 3120
rect 10320 3070 10360 3100
rect 10320 3050 10330 3070
rect 10350 3050 10360 3070
rect 10320 3020 10360 3050
rect 10320 3000 10330 3020
rect 10350 3000 10360 3020
rect 10320 2985 10360 3000
rect 10375 3570 10415 3585
rect 10375 3550 10385 3570
rect 10405 3550 10415 3570
rect 10375 3520 10415 3550
rect 10375 3500 10385 3520
rect 10405 3500 10415 3520
rect 10375 3470 10415 3500
rect 10375 3450 10385 3470
rect 10405 3450 10415 3470
rect 10375 3420 10415 3450
rect 10375 3400 10385 3420
rect 10405 3400 10415 3420
rect 10375 3370 10415 3400
rect 10375 3350 10385 3370
rect 10405 3350 10415 3370
rect 10375 3320 10415 3350
rect 10375 3300 10385 3320
rect 10405 3300 10415 3320
rect 10375 3270 10415 3300
rect 10375 3250 10385 3270
rect 10405 3250 10415 3270
rect 10375 3220 10415 3250
rect 10375 3200 10385 3220
rect 10405 3200 10415 3220
rect 10375 3170 10415 3200
rect 10375 3150 10385 3170
rect 10405 3150 10415 3170
rect 10375 3120 10415 3150
rect 10375 3100 10385 3120
rect 10405 3100 10415 3120
rect 10375 3070 10415 3100
rect 10375 3050 10385 3070
rect 10405 3050 10415 3070
rect 10375 3020 10415 3050
rect 10375 3000 10385 3020
rect 10405 3000 10415 3020
rect 10375 2985 10415 3000
rect 10430 3570 10470 3585
rect 10430 3550 10440 3570
rect 10460 3550 10470 3570
rect 10430 3520 10470 3550
rect 10430 3500 10440 3520
rect 10460 3500 10470 3520
rect 10430 3470 10470 3500
rect 10430 3450 10440 3470
rect 10460 3450 10470 3470
rect 10430 3420 10470 3450
rect 10430 3400 10440 3420
rect 10460 3400 10470 3420
rect 10430 3370 10470 3400
rect 10430 3350 10440 3370
rect 10460 3350 10470 3370
rect 10430 3320 10470 3350
rect 10430 3300 10440 3320
rect 10460 3300 10470 3320
rect 10430 3270 10470 3300
rect 10430 3250 10440 3270
rect 10460 3250 10470 3270
rect 10430 3220 10470 3250
rect 10430 3200 10440 3220
rect 10460 3200 10470 3220
rect 10430 3170 10470 3200
rect 10430 3150 10440 3170
rect 10460 3150 10470 3170
rect 10430 3120 10470 3150
rect 10430 3100 10440 3120
rect 10460 3100 10470 3120
rect 10430 3070 10470 3100
rect 10430 3050 10440 3070
rect 10460 3050 10470 3070
rect 10430 3020 10470 3050
rect 10430 3000 10440 3020
rect 10460 3000 10470 3020
rect 10430 2985 10470 3000
rect 10485 3570 10525 3585
rect 10485 3550 10495 3570
rect 10515 3550 10525 3570
rect 10485 3520 10525 3550
rect 10485 3500 10495 3520
rect 10515 3500 10525 3520
rect 10485 3470 10525 3500
rect 10485 3450 10495 3470
rect 10515 3450 10525 3470
rect 10485 3420 10525 3450
rect 10485 3400 10495 3420
rect 10515 3400 10525 3420
rect 10485 3370 10525 3400
rect 10485 3350 10495 3370
rect 10515 3350 10525 3370
rect 10485 3320 10525 3350
rect 10485 3300 10495 3320
rect 10515 3300 10525 3320
rect 10485 3270 10525 3300
rect 10485 3250 10495 3270
rect 10515 3250 10525 3270
rect 10485 3220 10525 3250
rect 10485 3200 10495 3220
rect 10515 3200 10525 3220
rect 10485 3170 10525 3200
rect 10485 3150 10495 3170
rect 10515 3150 10525 3170
rect 10485 3120 10525 3150
rect 10485 3100 10495 3120
rect 10515 3100 10525 3120
rect 10485 3070 10525 3100
rect 10485 3050 10495 3070
rect 10515 3050 10525 3070
rect 10485 3020 10525 3050
rect 10485 3000 10495 3020
rect 10515 3000 10525 3020
rect 10485 2985 10525 3000
rect 10540 3570 10580 3585
rect 10540 3550 10550 3570
rect 10570 3550 10580 3570
rect 10540 3520 10580 3550
rect 10540 3500 10550 3520
rect 10570 3500 10580 3520
rect 10540 3470 10580 3500
rect 10540 3450 10550 3470
rect 10570 3450 10580 3470
rect 10540 3420 10580 3450
rect 10540 3400 10550 3420
rect 10570 3400 10580 3420
rect 10540 3370 10580 3400
rect 10540 3350 10550 3370
rect 10570 3350 10580 3370
rect 10540 3320 10580 3350
rect 10540 3300 10550 3320
rect 10570 3300 10580 3320
rect 10540 3270 10580 3300
rect 10540 3250 10550 3270
rect 10570 3250 10580 3270
rect 10540 3220 10580 3250
rect 10540 3200 10550 3220
rect 10570 3200 10580 3220
rect 10540 3170 10580 3200
rect 10540 3150 10550 3170
rect 10570 3150 10580 3170
rect 10540 3120 10580 3150
rect 10540 3100 10550 3120
rect 10570 3100 10580 3120
rect 10540 3070 10580 3100
rect 10540 3050 10550 3070
rect 10570 3050 10580 3070
rect 10540 3020 10580 3050
rect 10540 3000 10550 3020
rect 10570 3000 10580 3020
rect 10540 2985 10580 3000
rect 10595 3570 10635 3585
rect 10595 3550 10605 3570
rect 10625 3550 10635 3570
rect 10595 3520 10635 3550
rect 10595 3500 10605 3520
rect 10625 3500 10635 3520
rect 10595 3470 10635 3500
rect 10595 3450 10605 3470
rect 10625 3450 10635 3470
rect 10595 3420 10635 3450
rect 10595 3400 10605 3420
rect 10625 3400 10635 3420
rect 10595 3370 10635 3400
rect 10595 3350 10605 3370
rect 10625 3350 10635 3370
rect 10595 3320 10635 3350
rect 10595 3300 10605 3320
rect 10625 3300 10635 3320
rect 10595 3270 10635 3300
rect 10595 3250 10605 3270
rect 10625 3250 10635 3270
rect 10595 3220 10635 3250
rect 10595 3200 10605 3220
rect 10625 3200 10635 3220
rect 10595 3170 10635 3200
rect 10595 3150 10605 3170
rect 10625 3150 10635 3170
rect 10595 3120 10635 3150
rect 10595 3100 10605 3120
rect 10625 3100 10635 3120
rect 10595 3070 10635 3100
rect 10595 3050 10605 3070
rect 10625 3050 10635 3070
rect 10595 3020 10635 3050
rect 10595 3000 10605 3020
rect 10625 3000 10635 3020
rect 10595 2985 10635 3000
rect 10650 3570 10690 3585
rect 10650 3550 10660 3570
rect 10680 3550 10690 3570
rect 10650 3520 10690 3550
rect 10650 3500 10660 3520
rect 10680 3500 10690 3520
rect 10650 3470 10690 3500
rect 10650 3450 10660 3470
rect 10680 3450 10690 3470
rect 10650 3420 10690 3450
rect 10650 3400 10660 3420
rect 10680 3400 10690 3420
rect 10650 3370 10690 3400
rect 10650 3350 10660 3370
rect 10680 3350 10690 3370
rect 10650 3320 10690 3350
rect 10650 3300 10660 3320
rect 10680 3300 10690 3320
rect 10650 3270 10690 3300
rect 10650 3250 10660 3270
rect 10680 3250 10690 3270
rect 10650 3220 10690 3250
rect 10650 3200 10660 3220
rect 10680 3200 10690 3220
rect 10650 3170 10690 3200
rect 10650 3150 10660 3170
rect 10680 3150 10690 3170
rect 10650 3120 10690 3150
rect 10650 3100 10660 3120
rect 10680 3100 10690 3120
rect 10650 3070 10690 3100
rect 10650 3050 10660 3070
rect 10680 3050 10690 3070
rect 10650 3020 10690 3050
rect 10650 3000 10660 3020
rect 10680 3000 10690 3020
rect 10650 2985 10690 3000
rect 10705 3570 10745 3585
rect 10705 3550 10715 3570
rect 10735 3550 10745 3570
rect 10705 3520 10745 3550
rect 10705 3500 10715 3520
rect 10735 3500 10745 3520
rect 10705 3470 10745 3500
rect 10705 3450 10715 3470
rect 10735 3450 10745 3470
rect 10705 3420 10745 3450
rect 10705 3400 10715 3420
rect 10735 3400 10745 3420
rect 10705 3370 10745 3400
rect 10705 3350 10715 3370
rect 10735 3350 10745 3370
rect 10705 3320 10745 3350
rect 10705 3300 10715 3320
rect 10735 3300 10745 3320
rect 10705 3270 10745 3300
rect 10705 3250 10715 3270
rect 10735 3250 10745 3270
rect 10705 3220 10745 3250
rect 10705 3200 10715 3220
rect 10735 3200 10745 3220
rect 10705 3170 10745 3200
rect 10705 3150 10715 3170
rect 10735 3150 10745 3170
rect 10705 3120 10745 3150
rect 10705 3100 10715 3120
rect 10735 3100 10745 3120
rect 10705 3070 10745 3100
rect 10705 3050 10715 3070
rect 10735 3050 10745 3070
rect 10705 3020 10745 3050
rect 10705 3000 10715 3020
rect 10735 3000 10745 3020
rect 10705 2985 10745 3000
rect 10760 3570 10800 3585
rect 10760 3550 10770 3570
rect 10790 3550 10800 3570
rect 10760 3520 10800 3550
rect 10760 3500 10770 3520
rect 10790 3500 10800 3520
rect 10760 3470 10800 3500
rect 10760 3450 10770 3470
rect 10790 3450 10800 3470
rect 10760 3420 10800 3450
rect 10760 3400 10770 3420
rect 10790 3400 10800 3420
rect 10760 3370 10800 3400
rect 10760 3350 10770 3370
rect 10790 3350 10800 3370
rect 10760 3320 10800 3350
rect 10760 3300 10770 3320
rect 10790 3300 10800 3320
rect 10760 3270 10800 3300
rect 10760 3250 10770 3270
rect 10790 3250 10800 3270
rect 10760 3220 10800 3250
rect 10760 3200 10770 3220
rect 10790 3200 10800 3220
rect 10760 3170 10800 3200
rect 10760 3150 10770 3170
rect 10790 3150 10800 3170
rect 10760 3120 10800 3150
rect 10760 3100 10770 3120
rect 10790 3100 10800 3120
rect 10760 3070 10800 3100
rect 10760 3050 10770 3070
rect 10790 3050 10800 3070
rect 10760 3020 10800 3050
rect 10760 3000 10770 3020
rect 10790 3000 10800 3020
rect 10760 2985 10800 3000
rect 10815 3570 10855 3585
rect 10815 3550 10825 3570
rect 10845 3550 10855 3570
rect 10815 3520 10855 3550
rect 10815 3500 10825 3520
rect 10845 3500 10855 3520
rect 10815 3470 10855 3500
rect 10815 3450 10825 3470
rect 10845 3450 10855 3470
rect 10815 3420 10855 3450
rect 10815 3400 10825 3420
rect 10845 3400 10855 3420
rect 10815 3370 10855 3400
rect 10815 3350 10825 3370
rect 10845 3350 10855 3370
rect 10815 3320 10855 3350
rect 10815 3300 10825 3320
rect 10845 3300 10855 3320
rect 10815 3270 10855 3300
rect 10815 3250 10825 3270
rect 10845 3250 10855 3270
rect 10815 3220 10855 3250
rect 10815 3200 10825 3220
rect 10845 3200 10855 3220
rect 10815 3170 10855 3200
rect 11220 3560 11260 3575
rect 11220 3540 11230 3560
rect 11250 3540 11260 3560
rect 11220 3510 11260 3540
rect 11220 3490 11230 3510
rect 11250 3490 11260 3510
rect 11220 3460 11260 3490
rect 11220 3440 11230 3460
rect 11250 3440 11260 3460
rect 11220 3410 11260 3440
rect 11220 3390 11230 3410
rect 11250 3390 11260 3410
rect 11220 3360 11260 3390
rect 11220 3340 11230 3360
rect 11250 3340 11260 3360
rect 11220 3310 11260 3340
rect 11220 3290 11230 3310
rect 11250 3290 11260 3310
rect 11220 3260 11260 3290
rect 11220 3240 11230 3260
rect 11250 3240 11260 3260
rect 11220 3210 11260 3240
rect 11220 3190 11230 3210
rect 11250 3190 11260 3210
rect 11220 3175 11260 3190
rect 11280 3560 11320 3575
rect 11280 3540 11290 3560
rect 11310 3540 11320 3560
rect 11280 3510 11320 3540
rect 11280 3490 11290 3510
rect 11310 3490 11320 3510
rect 11280 3460 11320 3490
rect 11280 3440 11290 3460
rect 11310 3440 11320 3460
rect 11280 3410 11320 3440
rect 11280 3390 11290 3410
rect 11310 3390 11320 3410
rect 11280 3360 11320 3390
rect 11280 3340 11290 3360
rect 11310 3340 11320 3360
rect 11280 3310 11320 3340
rect 11280 3290 11290 3310
rect 11310 3290 11320 3310
rect 11280 3260 11320 3290
rect 11280 3240 11290 3260
rect 11310 3240 11320 3260
rect 11280 3210 11320 3240
rect 11280 3190 11290 3210
rect 11310 3190 11320 3210
rect 11280 3175 11320 3190
rect 11340 3560 11380 3575
rect 11340 3540 11350 3560
rect 11370 3540 11380 3560
rect 11340 3510 11380 3540
rect 11340 3490 11350 3510
rect 11370 3490 11380 3510
rect 11340 3460 11380 3490
rect 11340 3440 11350 3460
rect 11370 3440 11380 3460
rect 11340 3410 11380 3440
rect 11340 3390 11350 3410
rect 11370 3390 11380 3410
rect 11340 3360 11380 3390
rect 11340 3340 11350 3360
rect 11370 3340 11380 3360
rect 11340 3310 11380 3340
rect 11340 3290 11350 3310
rect 11370 3290 11380 3310
rect 11340 3260 11380 3290
rect 11340 3240 11350 3260
rect 11370 3240 11380 3260
rect 11340 3210 11380 3240
rect 11340 3190 11350 3210
rect 11370 3190 11380 3210
rect 11340 3175 11380 3190
rect 11400 3560 11440 3575
rect 11400 3540 11410 3560
rect 11430 3540 11440 3560
rect 11400 3510 11440 3540
rect 11400 3490 11410 3510
rect 11430 3490 11440 3510
rect 11400 3460 11440 3490
rect 11400 3440 11410 3460
rect 11430 3440 11440 3460
rect 11400 3410 11440 3440
rect 11400 3390 11410 3410
rect 11430 3390 11440 3410
rect 11400 3360 11440 3390
rect 11400 3340 11410 3360
rect 11430 3340 11440 3360
rect 11400 3310 11440 3340
rect 11400 3290 11410 3310
rect 11430 3290 11440 3310
rect 11400 3260 11440 3290
rect 11400 3240 11410 3260
rect 11430 3240 11440 3260
rect 11400 3210 11440 3240
rect 11400 3190 11410 3210
rect 11430 3190 11440 3210
rect 11400 3175 11440 3190
rect 11460 3560 11500 3575
rect 11460 3540 11470 3560
rect 11490 3540 11500 3560
rect 11460 3510 11500 3540
rect 11460 3490 11470 3510
rect 11490 3490 11500 3510
rect 11460 3460 11500 3490
rect 11460 3440 11470 3460
rect 11490 3440 11500 3460
rect 11460 3410 11500 3440
rect 11460 3390 11470 3410
rect 11490 3390 11500 3410
rect 11460 3360 11500 3390
rect 11460 3340 11470 3360
rect 11490 3340 11500 3360
rect 11460 3310 11500 3340
rect 11460 3290 11470 3310
rect 11490 3290 11500 3310
rect 11460 3260 11500 3290
rect 11460 3240 11470 3260
rect 11490 3240 11500 3260
rect 11460 3210 11500 3240
rect 11460 3190 11470 3210
rect 11490 3190 11500 3210
rect 11460 3175 11500 3190
rect 11520 3560 11560 3575
rect 11520 3540 11530 3560
rect 11550 3540 11560 3560
rect 11520 3510 11560 3540
rect 11520 3490 11530 3510
rect 11550 3490 11560 3510
rect 11520 3460 11560 3490
rect 11520 3440 11530 3460
rect 11550 3440 11560 3460
rect 11520 3410 11560 3440
rect 11520 3390 11530 3410
rect 11550 3390 11560 3410
rect 11520 3360 11560 3390
rect 11520 3340 11530 3360
rect 11550 3340 11560 3360
rect 11520 3310 11560 3340
rect 11520 3290 11530 3310
rect 11550 3290 11560 3310
rect 11520 3260 11560 3290
rect 11520 3240 11530 3260
rect 11550 3240 11560 3260
rect 11520 3210 11560 3240
rect 11520 3190 11530 3210
rect 11550 3190 11560 3210
rect 11520 3175 11560 3190
rect 11580 3560 11620 3575
rect 11580 3540 11590 3560
rect 11610 3540 11620 3560
rect 11580 3510 11620 3540
rect 11580 3490 11590 3510
rect 11610 3490 11620 3510
rect 11580 3460 11620 3490
rect 11580 3440 11590 3460
rect 11610 3440 11620 3460
rect 11580 3410 11620 3440
rect 11580 3390 11590 3410
rect 11610 3390 11620 3410
rect 11580 3360 11620 3390
rect 11580 3340 11590 3360
rect 11610 3340 11620 3360
rect 11580 3310 11620 3340
rect 11580 3290 11590 3310
rect 11610 3290 11620 3310
rect 11580 3260 11620 3290
rect 11580 3240 11590 3260
rect 11610 3240 11620 3260
rect 11580 3210 11620 3240
rect 11580 3190 11590 3210
rect 11610 3190 11620 3210
rect 11580 3175 11620 3190
rect 11640 3560 11680 3575
rect 11640 3540 11650 3560
rect 11670 3540 11680 3560
rect 11640 3510 11680 3540
rect 11640 3490 11650 3510
rect 11670 3490 11680 3510
rect 11640 3460 11680 3490
rect 11640 3440 11650 3460
rect 11670 3440 11680 3460
rect 11640 3410 11680 3440
rect 11640 3390 11650 3410
rect 11670 3390 11680 3410
rect 11640 3360 11680 3390
rect 11640 3340 11650 3360
rect 11670 3340 11680 3360
rect 11640 3310 11680 3340
rect 11640 3290 11650 3310
rect 11670 3290 11680 3310
rect 11640 3260 11680 3290
rect 11640 3240 11650 3260
rect 11670 3240 11680 3260
rect 11640 3210 11680 3240
rect 11640 3190 11650 3210
rect 11670 3190 11680 3210
rect 11640 3175 11680 3190
rect 11700 3560 11740 3575
rect 11700 3540 11710 3560
rect 11730 3540 11740 3560
rect 11700 3510 11740 3540
rect 11700 3490 11710 3510
rect 11730 3490 11740 3510
rect 11700 3460 11740 3490
rect 11700 3440 11710 3460
rect 11730 3440 11740 3460
rect 11700 3410 11740 3440
rect 11700 3390 11710 3410
rect 11730 3390 11740 3410
rect 11700 3360 11740 3390
rect 11700 3340 11710 3360
rect 11730 3340 11740 3360
rect 11700 3310 11740 3340
rect 11700 3290 11710 3310
rect 11730 3290 11740 3310
rect 11700 3260 11740 3290
rect 11700 3240 11710 3260
rect 11730 3240 11740 3260
rect 11700 3210 11740 3240
rect 11700 3190 11710 3210
rect 11730 3190 11740 3210
rect 11700 3175 11740 3190
rect 11760 3560 11800 3575
rect 11760 3540 11770 3560
rect 11790 3540 11800 3560
rect 11760 3510 11800 3540
rect 11760 3490 11770 3510
rect 11790 3490 11800 3510
rect 11760 3460 11800 3490
rect 11760 3440 11770 3460
rect 11790 3440 11800 3460
rect 11760 3410 11800 3440
rect 11760 3390 11770 3410
rect 11790 3390 11800 3410
rect 11760 3360 11800 3390
rect 11760 3340 11770 3360
rect 11790 3340 11800 3360
rect 11760 3310 11800 3340
rect 11760 3290 11770 3310
rect 11790 3290 11800 3310
rect 11760 3260 11800 3290
rect 11760 3240 11770 3260
rect 11790 3240 11800 3260
rect 11760 3210 11800 3240
rect 11760 3190 11770 3210
rect 11790 3190 11800 3210
rect 11760 3175 11800 3190
rect 11820 3560 11860 3575
rect 11820 3540 11830 3560
rect 11850 3540 11860 3560
rect 11820 3510 11860 3540
rect 11820 3490 11830 3510
rect 11850 3490 11860 3510
rect 11820 3460 11860 3490
rect 11820 3440 11830 3460
rect 11850 3440 11860 3460
rect 11820 3410 11860 3440
rect 11820 3390 11830 3410
rect 11850 3390 11860 3410
rect 11820 3360 11860 3390
rect 11820 3340 11830 3360
rect 11850 3340 11860 3360
rect 11820 3310 11860 3340
rect 11820 3290 11830 3310
rect 11850 3290 11860 3310
rect 11820 3260 11860 3290
rect 11820 3240 11830 3260
rect 11850 3240 11860 3260
rect 11820 3210 11860 3240
rect 11820 3190 11830 3210
rect 11850 3190 11860 3210
rect 11820 3175 11860 3190
rect 11880 3560 11920 3575
rect 11880 3540 11890 3560
rect 11910 3540 11920 3560
rect 11880 3510 11920 3540
rect 11880 3490 11890 3510
rect 11910 3490 11920 3510
rect 11880 3460 11920 3490
rect 11880 3440 11890 3460
rect 11910 3440 11920 3460
rect 11880 3410 11920 3440
rect 11880 3390 11890 3410
rect 11910 3390 11920 3410
rect 11880 3360 11920 3390
rect 11880 3340 11890 3360
rect 11910 3340 11920 3360
rect 11880 3310 11920 3340
rect 11880 3290 11890 3310
rect 11910 3290 11920 3310
rect 11880 3260 11920 3290
rect 11880 3240 11890 3260
rect 11910 3240 11920 3260
rect 11880 3210 11920 3240
rect 11880 3190 11890 3210
rect 11910 3190 11920 3210
rect 11880 3175 11920 3190
rect 11940 3560 11980 3575
rect 11940 3540 11950 3560
rect 11970 3540 11980 3560
rect 11940 3510 11980 3540
rect 11940 3490 11950 3510
rect 11970 3490 11980 3510
rect 11940 3460 11980 3490
rect 11940 3440 11950 3460
rect 11970 3440 11980 3460
rect 11940 3410 11980 3440
rect 11940 3390 11950 3410
rect 11970 3390 11980 3410
rect 11940 3360 11980 3390
rect 11940 3340 11950 3360
rect 11970 3340 11980 3360
rect 11940 3310 11980 3340
rect 11940 3290 11950 3310
rect 11970 3290 11980 3310
rect 11940 3260 11980 3290
rect 11940 3240 11950 3260
rect 11970 3240 11980 3260
rect 11940 3210 11980 3240
rect 11940 3190 11950 3210
rect 11970 3190 11980 3210
rect 11940 3175 11980 3190
rect 12000 3560 12040 3575
rect 12000 3540 12010 3560
rect 12030 3540 12040 3560
rect 12000 3510 12040 3540
rect 12000 3490 12010 3510
rect 12030 3490 12040 3510
rect 12000 3460 12040 3490
rect 12000 3440 12010 3460
rect 12030 3440 12040 3460
rect 12000 3410 12040 3440
rect 12000 3390 12010 3410
rect 12030 3390 12040 3410
rect 12000 3360 12040 3390
rect 12000 3340 12010 3360
rect 12030 3340 12040 3360
rect 12000 3310 12040 3340
rect 12000 3290 12010 3310
rect 12030 3290 12040 3310
rect 12000 3260 12040 3290
rect 12000 3240 12010 3260
rect 12030 3240 12040 3260
rect 12000 3210 12040 3240
rect 12000 3190 12010 3210
rect 12030 3190 12040 3210
rect 12000 3175 12040 3190
rect 12060 3560 12100 3575
rect 12060 3540 12070 3560
rect 12090 3540 12100 3560
rect 12060 3510 12100 3540
rect 12060 3490 12070 3510
rect 12090 3490 12100 3510
rect 12060 3460 12100 3490
rect 12060 3440 12070 3460
rect 12090 3440 12100 3460
rect 12060 3410 12100 3440
rect 12060 3390 12070 3410
rect 12090 3390 12100 3410
rect 12060 3360 12100 3390
rect 12060 3340 12070 3360
rect 12090 3340 12100 3360
rect 12060 3310 12100 3340
rect 12060 3290 12070 3310
rect 12090 3290 12100 3310
rect 12060 3260 12100 3290
rect 12060 3240 12070 3260
rect 12090 3240 12100 3260
rect 12060 3210 12100 3240
rect 12060 3190 12070 3210
rect 12090 3190 12100 3210
rect 12060 3175 12100 3190
rect 12120 3560 12160 3575
rect 12120 3540 12130 3560
rect 12150 3540 12160 3560
rect 12120 3510 12160 3540
rect 12120 3490 12130 3510
rect 12150 3490 12160 3510
rect 12120 3460 12160 3490
rect 12120 3440 12130 3460
rect 12150 3440 12160 3460
rect 12120 3410 12160 3440
rect 12120 3390 12130 3410
rect 12150 3390 12160 3410
rect 12120 3360 12160 3390
rect 12120 3340 12130 3360
rect 12150 3340 12160 3360
rect 12120 3310 12160 3340
rect 12120 3290 12130 3310
rect 12150 3290 12160 3310
rect 12120 3260 12160 3290
rect 12120 3240 12130 3260
rect 12150 3240 12160 3260
rect 12120 3210 12160 3240
rect 12120 3190 12130 3210
rect 12150 3190 12160 3210
rect 12120 3175 12160 3190
rect 12180 3560 12220 3575
rect 12180 3540 12190 3560
rect 12210 3540 12220 3560
rect 12180 3510 12220 3540
rect 12180 3490 12190 3510
rect 12210 3490 12220 3510
rect 12180 3460 12220 3490
rect 12180 3440 12190 3460
rect 12210 3440 12220 3460
rect 12180 3410 12220 3440
rect 12180 3390 12190 3410
rect 12210 3390 12220 3410
rect 12180 3360 12220 3390
rect 12180 3340 12190 3360
rect 12210 3340 12220 3360
rect 12180 3310 12220 3340
rect 12180 3290 12190 3310
rect 12210 3290 12220 3310
rect 12180 3260 12220 3290
rect 12180 3240 12190 3260
rect 12210 3240 12220 3260
rect 12180 3210 12220 3240
rect 12180 3190 12190 3210
rect 12210 3190 12220 3210
rect 12180 3175 12220 3190
rect 12240 3560 12280 3575
rect 12240 3540 12250 3560
rect 12270 3540 12280 3560
rect 12240 3510 12280 3540
rect 12240 3490 12250 3510
rect 12270 3490 12280 3510
rect 12240 3460 12280 3490
rect 12240 3440 12250 3460
rect 12270 3440 12280 3460
rect 12240 3410 12280 3440
rect 12240 3390 12250 3410
rect 12270 3390 12280 3410
rect 12240 3360 12280 3390
rect 12240 3340 12250 3360
rect 12270 3340 12280 3360
rect 12240 3310 12280 3340
rect 12240 3290 12250 3310
rect 12270 3290 12280 3310
rect 12240 3260 12280 3290
rect 12240 3240 12250 3260
rect 12270 3240 12280 3260
rect 12240 3210 12280 3240
rect 12240 3190 12250 3210
rect 12270 3190 12280 3210
rect 12240 3175 12280 3190
rect 12300 3560 12340 3575
rect 12300 3540 12310 3560
rect 12330 3540 12340 3560
rect 12300 3510 12340 3540
rect 12300 3490 12310 3510
rect 12330 3490 12340 3510
rect 12300 3460 12340 3490
rect 12300 3440 12310 3460
rect 12330 3440 12340 3460
rect 12300 3410 12340 3440
rect 12300 3390 12310 3410
rect 12330 3390 12340 3410
rect 12300 3360 12340 3390
rect 12300 3340 12310 3360
rect 12330 3340 12340 3360
rect 12300 3310 12340 3340
rect 12300 3290 12310 3310
rect 12330 3290 12340 3310
rect 12300 3260 12340 3290
rect 12300 3240 12310 3260
rect 12330 3240 12340 3260
rect 12300 3210 12340 3240
rect 12300 3190 12310 3210
rect 12330 3190 12340 3210
rect 12300 3175 12340 3190
rect 12360 3560 12400 3575
rect 12360 3540 12370 3560
rect 12390 3540 12400 3560
rect 12360 3510 12400 3540
rect 12360 3490 12370 3510
rect 12390 3490 12400 3510
rect 12360 3460 12400 3490
rect 12360 3440 12370 3460
rect 12390 3440 12400 3460
rect 12360 3410 12400 3440
rect 12360 3390 12370 3410
rect 12390 3390 12400 3410
rect 12360 3360 12400 3390
rect 12360 3340 12370 3360
rect 12390 3340 12400 3360
rect 12360 3310 12400 3340
rect 12360 3290 12370 3310
rect 12390 3290 12400 3310
rect 12360 3260 12400 3290
rect 12360 3240 12370 3260
rect 12390 3240 12400 3260
rect 12360 3210 12400 3240
rect 12360 3190 12370 3210
rect 12390 3190 12400 3210
rect 12360 3175 12400 3190
rect 12420 3560 12460 3575
rect 12420 3540 12430 3560
rect 12450 3540 12460 3560
rect 12420 3510 12460 3540
rect 12420 3490 12430 3510
rect 12450 3490 12460 3510
rect 12420 3460 12460 3490
rect 12420 3440 12430 3460
rect 12450 3440 12460 3460
rect 12420 3410 12460 3440
rect 12420 3390 12430 3410
rect 12450 3390 12460 3410
rect 12420 3360 12460 3390
rect 12420 3340 12430 3360
rect 12450 3340 12460 3360
rect 12420 3310 12460 3340
rect 12420 3290 12430 3310
rect 12450 3290 12460 3310
rect 12420 3260 12460 3290
rect 12420 3240 12430 3260
rect 12450 3240 12460 3260
rect 12420 3210 12460 3240
rect 12420 3190 12430 3210
rect 12450 3190 12460 3210
rect 12420 3175 12460 3190
rect 12480 3560 12520 3575
rect 12480 3540 12490 3560
rect 12510 3540 12520 3560
rect 12480 3510 12520 3540
rect 12480 3490 12490 3510
rect 12510 3490 12520 3510
rect 12480 3460 12520 3490
rect 12480 3440 12490 3460
rect 12510 3440 12520 3460
rect 12480 3410 12520 3440
rect 12480 3390 12490 3410
rect 12510 3390 12520 3410
rect 12480 3360 12520 3390
rect 12480 3340 12490 3360
rect 12510 3340 12520 3360
rect 12480 3310 12520 3340
rect 12480 3290 12490 3310
rect 12510 3290 12520 3310
rect 12480 3260 12520 3290
rect 12480 3240 12490 3260
rect 12510 3240 12520 3260
rect 12480 3210 12520 3240
rect 12480 3190 12490 3210
rect 12510 3190 12520 3210
rect 12480 3175 12520 3190
rect 12540 3560 12580 3575
rect 12540 3540 12550 3560
rect 12570 3540 12580 3560
rect 12540 3510 12580 3540
rect 12540 3490 12550 3510
rect 12570 3490 12580 3510
rect 12540 3460 12580 3490
rect 12540 3440 12550 3460
rect 12570 3440 12580 3460
rect 12540 3410 12580 3440
rect 12540 3390 12550 3410
rect 12570 3390 12580 3410
rect 12540 3360 12580 3390
rect 12540 3340 12550 3360
rect 12570 3340 12580 3360
rect 12540 3310 12580 3340
rect 12540 3290 12550 3310
rect 12570 3290 12580 3310
rect 12540 3260 12580 3290
rect 12540 3240 12550 3260
rect 12570 3240 12580 3260
rect 12540 3210 12580 3240
rect 12540 3190 12550 3210
rect 12570 3190 12580 3210
rect 12540 3175 12580 3190
rect 12945 3570 12985 3585
rect 12945 3550 12955 3570
rect 12975 3550 12985 3570
rect 12945 3520 12985 3550
rect 12945 3500 12955 3520
rect 12975 3500 12985 3520
rect 12945 3470 12985 3500
rect 12945 3450 12955 3470
rect 12975 3450 12985 3470
rect 12945 3420 12985 3450
rect 12945 3400 12955 3420
rect 12975 3400 12985 3420
rect 12945 3370 12985 3400
rect 12945 3350 12955 3370
rect 12975 3350 12985 3370
rect 12945 3320 12985 3350
rect 12945 3300 12955 3320
rect 12975 3300 12985 3320
rect 12945 3270 12985 3300
rect 12945 3250 12955 3270
rect 12975 3250 12985 3270
rect 12945 3220 12985 3250
rect 12945 3200 12955 3220
rect 12975 3200 12985 3220
rect 10815 3150 10825 3170
rect 10845 3150 10855 3170
rect 12945 3170 12985 3200
rect 12945 3150 12955 3170
rect 12975 3150 12985 3170
rect 10815 3120 10855 3150
rect 12945 3120 12985 3150
rect 10815 3100 10825 3120
rect 10845 3100 10855 3120
rect 10815 3070 10855 3100
rect 10815 3050 10825 3070
rect 10845 3050 10855 3070
rect 10815 3020 10855 3050
rect 10815 3000 10825 3020
rect 10845 3000 10855 3020
rect 10815 2985 10855 3000
rect 12945 3100 12955 3120
rect 12975 3100 12985 3120
rect 12945 3070 12985 3100
rect 12945 3050 12955 3070
rect 12975 3050 12985 3070
rect 12945 3020 12985 3050
rect 12945 3000 12955 3020
rect 12975 3000 12985 3020
rect 12945 2985 12985 3000
rect 13000 3570 13040 3585
rect 13000 3550 13010 3570
rect 13030 3550 13040 3570
rect 13000 3520 13040 3550
rect 13000 3500 13010 3520
rect 13030 3500 13040 3520
rect 13000 3470 13040 3500
rect 13000 3450 13010 3470
rect 13030 3450 13040 3470
rect 13000 3420 13040 3450
rect 13000 3400 13010 3420
rect 13030 3400 13040 3420
rect 13000 3370 13040 3400
rect 13000 3350 13010 3370
rect 13030 3350 13040 3370
rect 13000 3320 13040 3350
rect 13000 3300 13010 3320
rect 13030 3300 13040 3320
rect 13000 3270 13040 3300
rect 13000 3250 13010 3270
rect 13030 3250 13040 3270
rect 13000 3220 13040 3250
rect 13000 3200 13010 3220
rect 13030 3200 13040 3220
rect 13000 3170 13040 3200
rect 13000 3150 13010 3170
rect 13030 3150 13040 3170
rect 13000 3120 13040 3150
rect 13000 3100 13010 3120
rect 13030 3100 13040 3120
rect 13000 3070 13040 3100
rect 13000 3050 13010 3070
rect 13030 3050 13040 3070
rect 13000 3020 13040 3050
rect 13000 3000 13010 3020
rect 13030 3000 13040 3020
rect 13000 2985 13040 3000
rect 13055 3570 13095 3585
rect 13055 3550 13065 3570
rect 13085 3550 13095 3570
rect 13055 3520 13095 3550
rect 13055 3500 13065 3520
rect 13085 3500 13095 3520
rect 13055 3470 13095 3500
rect 13055 3450 13065 3470
rect 13085 3450 13095 3470
rect 13055 3420 13095 3450
rect 13055 3400 13065 3420
rect 13085 3400 13095 3420
rect 13055 3370 13095 3400
rect 13055 3350 13065 3370
rect 13085 3350 13095 3370
rect 13055 3320 13095 3350
rect 13055 3300 13065 3320
rect 13085 3300 13095 3320
rect 13055 3270 13095 3300
rect 13055 3250 13065 3270
rect 13085 3250 13095 3270
rect 13055 3220 13095 3250
rect 13055 3200 13065 3220
rect 13085 3200 13095 3220
rect 13055 3170 13095 3200
rect 13055 3150 13065 3170
rect 13085 3150 13095 3170
rect 13055 3120 13095 3150
rect 13055 3100 13065 3120
rect 13085 3100 13095 3120
rect 13055 3070 13095 3100
rect 13055 3050 13065 3070
rect 13085 3050 13095 3070
rect 13055 3020 13095 3050
rect 13055 3000 13065 3020
rect 13085 3000 13095 3020
rect 13055 2985 13095 3000
rect 13110 3570 13150 3585
rect 13110 3550 13120 3570
rect 13140 3550 13150 3570
rect 13110 3520 13150 3550
rect 13110 3500 13120 3520
rect 13140 3500 13150 3520
rect 13110 3470 13150 3500
rect 13110 3450 13120 3470
rect 13140 3450 13150 3470
rect 13110 3420 13150 3450
rect 13110 3400 13120 3420
rect 13140 3400 13150 3420
rect 13110 3370 13150 3400
rect 13110 3350 13120 3370
rect 13140 3350 13150 3370
rect 13110 3320 13150 3350
rect 13110 3300 13120 3320
rect 13140 3300 13150 3320
rect 13110 3270 13150 3300
rect 13110 3250 13120 3270
rect 13140 3250 13150 3270
rect 13110 3220 13150 3250
rect 13110 3200 13120 3220
rect 13140 3200 13150 3220
rect 13110 3170 13150 3200
rect 13110 3150 13120 3170
rect 13140 3150 13150 3170
rect 13110 3120 13150 3150
rect 13110 3100 13120 3120
rect 13140 3100 13150 3120
rect 13110 3070 13150 3100
rect 13110 3050 13120 3070
rect 13140 3050 13150 3070
rect 13110 3020 13150 3050
rect 13110 3000 13120 3020
rect 13140 3000 13150 3020
rect 13110 2985 13150 3000
rect 13165 3570 13205 3585
rect 13165 3550 13175 3570
rect 13195 3550 13205 3570
rect 13165 3520 13205 3550
rect 13165 3500 13175 3520
rect 13195 3500 13205 3520
rect 13165 3470 13205 3500
rect 13165 3450 13175 3470
rect 13195 3450 13205 3470
rect 13165 3420 13205 3450
rect 13165 3400 13175 3420
rect 13195 3400 13205 3420
rect 13165 3370 13205 3400
rect 13165 3350 13175 3370
rect 13195 3350 13205 3370
rect 13165 3320 13205 3350
rect 13165 3300 13175 3320
rect 13195 3300 13205 3320
rect 13165 3270 13205 3300
rect 13165 3250 13175 3270
rect 13195 3250 13205 3270
rect 13165 3220 13205 3250
rect 13165 3200 13175 3220
rect 13195 3200 13205 3220
rect 13165 3170 13205 3200
rect 13165 3150 13175 3170
rect 13195 3150 13205 3170
rect 13165 3120 13205 3150
rect 13165 3100 13175 3120
rect 13195 3100 13205 3120
rect 13165 3070 13205 3100
rect 13165 3050 13175 3070
rect 13195 3050 13205 3070
rect 13165 3020 13205 3050
rect 13165 3000 13175 3020
rect 13195 3000 13205 3020
rect 13165 2985 13205 3000
rect 13220 3570 13260 3585
rect 13220 3550 13230 3570
rect 13250 3550 13260 3570
rect 13220 3520 13260 3550
rect 13220 3500 13230 3520
rect 13250 3500 13260 3520
rect 13220 3470 13260 3500
rect 13220 3450 13230 3470
rect 13250 3450 13260 3470
rect 13220 3420 13260 3450
rect 13220 3400 13230 3420
rect 13250 3400 13260 3420
rect 13220 3370 13260 3400
rect 13220 3350 13230 3370
rect 13250 3350 13260 3370
rect 13220 3320 13260 3350
rect 13220 3300 13230 3320
rect 13250 3300 13260 3320
rect 13220 3270 13260 3300
rect 13220 3250 13230 3270
rect 13250 3250 13260 3270
rect 13220 3220 13260 3250
rect 13220 3200 13230 3220
rect 13250 3200 13260 3220
rect 13220 3170 13260 3200
rect 13220 3150 13230 3170
rect 13250 3150 13260 3170
rect 13220 3120 13260 3150
rect 13220 3100 13230 3120
rect 13250 3100 13260 3120
rect 13220 3070 13260 3100
rect 13220 3050 13230 3070
rect 13250 3050 13260 3070
rect 13220 3020 13260 3050
rect 13220 3000 13230 3020
rect 13250 3000 13260 3020
rect 13220 2985 13260 3000
rect 13275 3570 13315 3585
rect 13275 3550 13285 3570
rect 13305 3550 13315 3570
rect 13275 3520 13315 3550
rect 13275 3500 13285 3520
rect 13305 3500 13315 3520
rect 13275 3470 13315 3500
rect 13275 3450 13285 3470
rect 13305 3450 13315 3470
rect 13275 3420 13315 3450
rect 13275 3400 13285 3420
rect 13305 3400 13315 3420
rect 13275 3370 13315 3400
rect 13275 3350 13285 3370
rect 13305 3350 13315 3370
rect 13275 3320 13315 3350
rect 13275 3300 13285 3320
rect 13305 3300 13315 3320
rect 13275 3270 13315 3300
rect 13275 3250 13285 3270
rect 13305 3250 13315 3270
rect 13275 3220 13315 3250
rect 13275 3200 13285 3220
rect 13305 3200 13315 3220
rect 13275 3170 13315 3200
rect 13275 3150 13285 3170
rect 13305 3150 13315 3170
rect 13275 3120 13315 3150
rect 13275 3100 13285 3120
rect 13305 3100 13315 3120
rect 13275 3070 13315 3100
rect 13275 3050 13285 3070
rect 13305 3050 13315 3070
rect 13275 3020 13315 3050
rect 13275 3000 13285 3020
rect 13305 3000 13315 3020
rect 13275 2985 13315 3000
rect 13330 3570 13370 3585
rect 13330 3550 13340 3570
rect 13360 3550 13370 3570
rect 13330 3520 13370 3550
rect 13330 3500 13340 3520
rect 13360 3500 13370 3520
rect 13330 3470 13370 3500
rect 13330 3450 13340 3470
rect 13360 3450 13370 3470
rect 13330 3420 13370 3450
rect 13330 3400 13340 3420
rect 13360 3400 13370 3420
rect 13330 3370 13370 3400
rect 13330 3350 13340 3370
rect 13360 3350 13370 3370
rect 13330 3320 13370 3350
rect 13330 3300 13340 3320
rect 13360 3300 13370 3320
rect 13330 3270 13370 3300
rect 13330 3250 13340 3270
rect 13360 3250 13370 3270
rect 13330 3220 13370 3250
rect 13330 3200 13340 3220
rect 13360 3200 13370 3220
rect 13330 3170 13370 3200
rect 13330 3150 13340 3170
rect 13360 3150 13370 3170
rect 13330 3120 13370 3150
rect 13330 3100 13340 3120
rect 13360 3100 13370 3120
rect 13330 3070 13370 3100
rect 13330 3050 13340 3070
rect 13360 3050 13370 3070
rect 13330 3020 13370 3050
rect 13330 3000 13340 3020
rect 13360 3000 13370 3020
rect 13330 2985 13370 3000
rect 13385 3570 13425 3585
rect 13385 3550 13395 3570
rect 13415 3550 13425 3570
rect 13385 3520 13425 3550
rect 13385 3500 13395 3520
rect 13415 3500 13425 3520
rect 13385 3470 13425 3500
rect 13385 3450 13395 3470
rect 13415 3450 13425 3470
rect 13385 3420 13425 3450
rect 13385 3400 13395 3420
rect 13415 3400 13425 3420
rect 13385 3370 13425 3400
rect 13385 3350 13395 3370
rect 13415 3350 13425 3370
rect 13385 3320 13425 3350
rect 13385 3300 13395 3320
rect 13415 3300 13425 3320
rect 13385 3270 13425 3300
rect 13385 3250 13395 3270
rect 13415 3250 13425 3270
rect 13385 3220 13425 3250
rect 13385 3200 13395 3220
rect 13415 3200 13425 3220
rect 13385 3170 13425 3200
rect 13385 3150 13395 3170
rect 13415 3150 13425 3170
rect 13385 3120 13425 3150
rect 13385 3100 13395 3120
rect 13415 3100 13425 3120
rect 13385 3070 13425 3100
rect 13385 3050 13395 3070
rect 13415 3050 13425 3070
rect 13385 3020 13425 3050
rect 13385 3000 13395 3020
rect 13415 3000 13425 3020
rect 13385 2985 13425 3000
rect 13440 3570 13480 3585
rect 13440 3550 13450 3570
rect 13470 3550 13480 3570
rect 13440 3520 13480 3550
rect 13440 3500 13450 3520
rect 13470 3500 13480 3520
rect 13440 3470 13480 3500
rect 13440 3450 13450 3470
rect 13470 3450 13480 3470
rect 13440 3420 13480 3450
rect 13440 3400 13450 3420
rect 13470 3400 13480 3420
rect 13440 3370 13480 3400
rect 13440 3350 13450 3370
rect 13470 3350 13480 3370
rect 13440 3320 13480 3350
rect 13440 3300 13450 3320
rect 13470 3300 13480 3320
rect 13440 3270 13480 3300
rect 13440 3250 13450 3270
rect 13470 3250 13480 3270
rect 13440 3220 13480 3250
rect 13440 3200 13450 3220
rect 13470 3200 13480 3220
rect 13440 3170 13480 3200
rect 13440 3150 13450 3170
rect 13470 3150 13480 3170
rect 13440 3120 13480 3150
rect 13440 3100 13450 3120
rect 13470 3100 13480 3120
rect 13440 3070 13480 3100
rect 13440 3050 13450 3070
rect 13470 3050 13480 3070
rect 13440 3020 13480 3050
rect 13440 3000 13450 3020
rect 13470 3000 13480 3020
rect 13440 2985 13480 3000
rect 13495 3570 13535 3585
rect 13495 3550 13505 3570
rect 13525 3550 13535 3570
rect 13495 3520 13535 3550
rect 13495 3500 13505 3520
rect 13525 3500 13535 3520
rect 13495 3470 13535 3500
rect 13495 3450 13505 3470
rect 13525 3450 13535 3470
rect 13495 3420 13535 3450
rect 13495 3400 13505 3420
rect 13525 3400 13535 3420
rect 13495 3370 13535 3400
rect 13495 3350 13505 3370
rect 13525 3350 13535 3370
rect 13495 3320 13535 3350
rect 13495 3300 13505 3320
rect 13525 3300 13535 3320
rect 13495 3270 13535 3300
rect 13495 3250 13505 3270
rect 13525 3250 13535 3270
rect 13495 3220 13535 3250
rect 13495 3200 13505 3220
rect 13525 3200 13535 3220
rect 13495 3170 13535 3200
rect 13495 3150 13505 3170
rect 13525 3150 13535 3170
rect 13495 3120 13535 3150
rect 13495 3100 13505 3120
rect 13525 3100 13535 3120
rect 13495 3070 13535 3100
rect 13495 3050 13505 3070
rect 13525 3050 13535 3070
rect 13495 3020 13535 3050
rect 13495 3000 13505 3020
rect 13525 3000 13535 3020
rect 13495 2985 13535 3000
rect 13550 3570 13590 3585
rect 13550 3550 13560 3570
rect 13580 3550 13590 3570
rect 13550 3520 13590 3550
rect 13550 3500 13560 3520
rect 13580 3500 13590 3520
rect 13550 3470 13590 3500
rect 13550 3450 13560 3470
rect 13580 3450 13590 3470
rect 13550 3420 13590 3450
rect 13550 3400 13560 3420
rect 13580 3400 13590 3420
rect 13550 3370 13590 3400
rect 13550 3350 13560 3370
rect 13580 3350 13590 3370
rect 13550 3320 13590 3350
rect 13550 3300 13560 3320
rect 13580 3300 13590 3320
rect 13550 3270 13590 3300
rect 13550 3250 13560 3270
rect 13580 3250 13590 3270
rect 13550 3220 13590 3250
rect 13550 3200 13560 3220
rect 13580 3200 13590 3220
rect 13550 3170 13590 3200
rect 13550 3150 13560 3170
rect 13580 3150 13590 3170
rect 13550 3120 13590 3150
rect 13550 3100 13560 3120
rect 13580 3100 13590 3120
rect 13550 3070 13590 3100
rect 13550 3050 13560 3070
rect 13580 3050 13590 3070
rect 13550 3020 13590 3050
rect 13550 3000 13560 3020
rect 13580 3000 13590 3020
rect 13550 2985 13590 3000
rect 13605 3570 13645 3585
rect 13605 3550 13615 3570
rect 13635 3550 13645 3570
rect 25955 3550 25980 3580
rect 13605 3520 13645 3550
rect 13605 3500 13615 3520
rect 13635 3500 13645 3520
rect 13605 3470 13645 3500
rect 13605 3450 13615 3470
rect 13635 3450 13645 3470
rect 13605 3420 13645 3450
rect 13605 3400 13615 3420
rect 13635 3400 13645 3420
rect 13605 3370 13645 3400
rect 13605 3350 13615 3370
rect 13635 3350 13645 3370
rect 13605 3320 13645 3350
rect 13605 3300 13615 3320
rect 13635 3300 13645 3320
rect 13605 3270 13645 3300
rect 13605 3250 13615 3270
rect 13635 3250 13645 3270
rect 13605 3220 13645 3250
rect 13605 3200 13615 3220
rect 13635 3200 13645 3220
rect 13605 3170 13645 3200
rect 13605 3150 13615 3170
rect 13635 3150 13645 3170
rect 13605 3120 13645 3150
rect 13605 3100 13615 3120
rect 13635 3100 13645 3120
rect 13605 3070 13645 3100
rect 13605 3050 13615 3070
rect 13635 3050 13645 3070
rect 13605 3020 13645 3050
rect 13605 3000 13615 3020
rect 13635 3000 13645 3020
rect 13605 2985 13645 3000
rect 25820 3515 25860 3550
rect 25820 3495 25830 3515
rect 25850 3495 25860 3515
rect 25820 3465 25860 3495
rect 25820 3445 25830 3465
rect 25850 3445 25860 3465
rect 25820 3415 25860 3445
rect 25820 3395 25830 3415
rect 25850 3395 25860 3415
rect 25820 3365 25860 3395
rect 25820 3345 25830 3365
rect 25850 3345 25860 3365
rect 25820 3315 25860 3345
rect 25820 3295 25830 3315
rect 25850 3295 25860 3315
rect 25490 3265 25530 3293
rect 25490 3245 25500 3265
rect 25520 3245 25530 3265
rect 25490 3230 25530 3245
rect 25550 3270 25590 3293
rect 25550 3250 25560 3270
rect 25580 3250 25590 3270
rect 25550 3230 25590 3250
rect 25610 3270 25650 3293
rect 25610 3250 25620 3270
rect 25640 3250 25650 3270
rect 25610 3230 25650 3250
rect 25670 3265 25710 3293
rect 25670 3245 25680 3265
rect 25700 3245 25710 3265
rect 25670 3230 25710 3245
rect 25820 3265 25860 3295
rect 25820 3245 25830 3265
rect 25850 3245 25860 3265
rect 25820 3230 25860 3245
rect 25880 3515 25920 3550
rect 25880 3495 25890 3515
rect 25910 3495 25920 3515
rect 25880 3465 25920 3495
rect 25880 3445 25890 3465
rect 25910 3445 25920 3465
rect 25880 3415 25920 3445
rect 25880 3395 25890 3415
rect 25910 3395 25920 3415
rect 25880 3365 25920 3395
rect 25880 3345 25890 3365
rect 25910 3345 25920 3365
rect 25880 3315 25920 3345
rect 25880 3295 25890 3315
rect 25910 3295 25920 3315
rect 25880 3265 25920 3295
rect 25880 3245 25890 3265
rect 25910 3245 25920 3265
rect 25880 3230 25920 3245
rect 25940 3515 25980 3550
rect 25940 3495 25950 3515
rect 25970 3495 25980 3515
rect 25940 3465 25980 3495
rect 25940 3445 25950 3465
rect 25970 3445 25980 3465
rect 25940 3415 25980 3445
rect 25940 3395 25950 3415
rect 25970 3395 25980 3415
rect 25940 3365 25980 3395
rect 25940 3345 25950 3365
rect 25970 3345 25980 3365
rect 25940 3315 25980 3345
rect 25940 3295 25950 3315
rect 25970 3295 25980 3315
rect 25940 3265 25980 3295
rect 25940 3245 25950 3265
rect 25970 3245 25980 3265
rect 25940 3230 25980 3245
rect 26000 3565 26040 3580
rect 26000 3545 26010 3565
rect 26030 3545 26040 3565
rect 26000 3515 26040 3545
rect 26000 3495 26010 3515
rect 26030 3495 26040 3515
rect 26000 3465 26040 3495
rect 26000 3445 26010 3465
rect 26030 3445 26040 3465
rect 26000 3415 26040 3445
rect 26000 3395 26010 3415
rect 26030 3395 26040 3415
rect 26000 3365 26040 3395
rect 26000 3345 26010 3365
rect 26030 3345 26040 3365
rect 26000 3315 26040 3345
rect 26000 3295 26010 3315
rect 26030 3295 26040 3315
rect 26000 3265 26040 3295
rect 26000 3245 26010 3265
rect 26030 3245 26040 3265
rect 26000 3230 26040 3245
rect 26060 3565 26100 3580
rect 26060 3545 26070 3565
rect 26090 3545 26100 3565
rect 26060 3515 26100 3545
rect 26060 3495 26070 3515
rect 26090 3495 26100 3515
rect 26060 3465 26100 3495
rect 26060 3445 26070 3465
rect 26090 3445 26100 3465
rect 26060 3415 26100 3445
rect 26060 3395 26070 3415
rect 26090 3395 26100 3415
rect 26060 3365 26100 3395
rect 26060 3345 26070 3365
rect 26090 3345 26100 3365
rect 26060 3315 26100 3345
rect 26060 3295 26070 3315
rect 26090 3295 26100 3315
rect 26060 3265 26100 3295
rect 26060 3245 26070 3265
rect 26090 3245 26100 3265
rect 26060 3230 26100 3245
rect 26220 3560 26260 3575
rect 26220 3540 26230 3560
rect 26250 3540 26260 3560
rect 26220 3510 26260 3540
rect 26220 3490 26230 3510
rect 26250 3490 26260 3510
rect 26220 3460 26260 3490
rect 26220 3440 26230 3460
rect 26250 3440 26260 3460
rect 26220 3410 26260 3440
rect 26220 3390 26230 3410
rect 26250 3390 26260 3410
rect 26220 3360 26260 3390
rect 26220 3340 26230 3360
rect 26250 3340 26260 3360
rect 26220 3310 26260 3340
rect 26220 3290 26230 3310
rect 26250 3290 26260 3310
rect 26220 3260 26260 3290
rect 26220 3240 26230 3260
rect 26250 3240 26260 3260
rect 26220 3210 26260 3240
rect 26220 3190 26230 3210
rect 26250 3190 26260 3210
rect 26220 3175 26260 3190
rect 26280 3560 26320 3575
rect 26280 3540 26290 3560
rect 26310 3540 26320 3560
rect 26280 3510 26320 3540
rect 26280 3490 26290 3510
rect 26310 3490 26320 3510
rect 26280 3460 26320 3490
rect 26280 3440 26290 3460
rect 26310 3440 26320 3460
rect 26280 3410 26320 3440
rect 26280 3390 26290 3410
rect 26310 3390 26320 3410
rect 26280 3360 26320 3390
rect 26280 3340 26290 3360
rect 26310 3340 26320 3360
rect 26280 3310 26320 3340
rect 26280 3290 26290 3310
rect 26310 3290 26320 3310
rect 26280 3260 26320 3290
rect 26280 3240 26290 3260
rect 26310 3240 26320 3260
rect 26280 3210 26320 3240
rect 26280 3190 26290 3210
rect 26310 3190 26320 3210
rect 26280 3175 26320 3190
rect 26340 3560 26380 3575
rect 26340 3540 26350 3560
rect 26370 3540 26380 3560
rect 26340 3510 26380 3540
rect 26340 3490 26350 3510
rect 26370 3490 26380 3510
rect 26340 3460 26380 3490
rect 26340 3440 26350 3460
rect 26370 3440 26380 3460
rect 26340 3410 26380 3440
rect 26340 3390 26350 3410
rect 26370 3390 26380 3410
rect 26340 3360 26380 3390
rect 26340 3340 26350 3360
rect 26370 3340 26380 3360
rect 26340 3310 26380 3340
rect 26340 3290 26350 3310
rect 26370 3290 26380 3310
rect 26340 3260 26380 3290
rect 26340 3240 26350 3260
rect 26370 3240 26380 3260
rect 26340 3210 26380 3240
rect 26340 3190 26350 3210
rect 26370 3190 26380 3210
rect 26340 3175 26380 3190
rect 26400 3560 26440 3575
rect 26400 3540 26410 3560
rect 26430 3540 26440 3560
rect 26400 3510 26440 3540
rect 26400 3490 26410 3510
rect 26430 3490 26440 3510
rect 26400 3460 26440 3490
rect 26400 3440 26410 3460
rect 26430 3440 26440 3460
rect 26400 3410 26440 3440
rect 26400 3390 26410 3410
rect 26430 3390 26440 3410
rect 26400 3360 26440 3390
rect 26400 3340 26410 3360
rect 26430 3340 26440 3360
rect 26400 3310 26440 3340
rect 26400 3290 26410 3310
rect 26430 3290 26440 3310
rect 26400 3260 26440 3290
rect 26400 3240 26410 3260
rect 26430 3240 26440 3260
rect 26400 3210 26440 3240
rect 26400 3190 26410 3210
rect 26430 3190 26440 3210
rect 26400 3175 26440 3190
rect 26460 3560 26500 3575
rect 26460 3540 26470 3560
rect 26490 3540 26500 3560
rect 26460 3510 26500 3540
rect 26460 3490 26470 3510
rect 26490 3490 26500 3510
rect 26460 3460 26500 3490
rect 26460 3440 26470 3460
rect 26490 3440 26500 3460
rect 26460 3410 26500 3440
rect 26460 3390 26470 3410
rect 26490 3390 26500 3410
rect 26460 3360 26500 3390
rect 26460 3340 26470 3360
rect 26490 3340 26500 3360
rect 26460 3310 26500 3340
rect 26460 3290 26470 3310
rect 26490 3290 26500 3310
rect 26460 3260 26500 3290
rect 26460 3240 26470 3260
rect 26490 3240 26500 3260
rect 26460 3210 26500 3240
rect 26460 3190 26470 3210
rect 26490 3190 26500 3210
rect 26460 3175 26500 3190
rect 26520 3560 26560 3575
rect 26520 3540 26530 3560
rect 26550 3540 26560 3560
rect 26520 3510 26560 3540
rect 26520 3490 26530 3510
rect 26550 3490 26560 3510
rect 26520 3460 26560 3490
rect 26520 3440 26530 3460
rect 26550 3440 26560 3460
rect 26520 3410 26560 3440
rect 26520 3390 26530 3410
rect 26550 3390 26560 3410
rect 26520 3360 26560 3390
rect 26520 3340 26530 3360
rect 26550 3340 26560 3360
rect 26520 3310 26560 3340
rect 26520 3290 26530 3310
rect 26550 3290 26560 3310
rect 26520 3260 26560 3290
rect 26520 3240 26530 3260
rect 26550 3240 26560 3260
rect 26520 3210 26560 3240
rect 26520 3190 26530 3210
rect 26550 3190 26560 3210
rect 26520 3175 26560 3190
rect 26580 3560 26620 3575
rect 26580 3540 26590 3560
rect 26610 3540 26620 3560
rect 26580 3510 26620 3540
rect 26580 3490 26590 3510
rect 26610 3490 26620 3510
rect 26580 3460 26620 3490
rect 26580 3440 26590 3460
rect 26610 3440 26620 3460
rect 26580 3410 26620 3440
rect 26580 3390 26590 3410
rect 26610 3390 26620 3410
rect 26580 3360 26620 3390
rect 26580 3340 26590 3360
rect 26610 3340 26620 3360
rect 26580 3310 26620 3340
rect 26580 3290 26590 3310
rect 26610 3290 26620 3310
rect 26580 3260 26620 3290
rect 26580 3240 26590 3260
rect 26610 3240 26620 3260
rect 26580 3210 26620 3240
rect 26580 3190 26590 3210
rect 26610 3190 26620 3210
rect 26580 3175 26620 3190
rect 26640 3560 26680 3575
rect 26640 3540 26650 3560
rect 26670 3540 26680 3560
rect 26640 3510 26680 3540
rect 26640 3490 26650 3510
rect 26670 3490 26680 3510
rect 26640 3460 26680 3490
rect 26640 3440 26650 3460
rect 26670 3440 26680 3460
rect 26640 3410 26680 3440
rect 26640 3390 26650 3410
rect 26670 3390 26680 3410
rect 26640 3360 26680 3390
rect 26640 3340 26650 3360
rect 26670 3340 26680 3360
rect 26640 3310 26680 3340
rect 26640 3290 26650 3310
rect 26670 3290 26680 3310
rect 26640 3260 26680 3290
rect 26640 3240 26650 3260
rect 26670 3240 26680 3260
rect 26640 3210 26680 3240
rect 26640 3190 26650 3210
rect 26670 3190 26680 3210
rect 26640 3175 26680 3190
rect 26700 3560 26740 3575
rect 26700 3540 26710 3560
rect 26730 3540 26740 3560
rect 26700 3510 26740 3540
rect 26700 3490 26710 3510
rect 26730 3490 26740 3510
rect 26700 3460 26740 3490
rect 26700 3440 26710 3460
rect 26730 3440 26740 3460
rect 26700 3410 26740 3440
rect 26700 3390 26710 3410
rect 26730 3390 26740 3410
rect 26700 3360 26740 3390
rect 26700 3340 26710 3360
rect 26730 3340 26740 3360
rect 26700 3310 26740 3340
rect 26700 3290 26710 3310
rect 26730 3290 26740 3310
rect 26700 3260 26740 3290
rect 26700 3240 26710 3260
rect 26730 3240 26740 3260
rect 26700 3210 26740 3240
rect 26700 3190 26710 3210
rect 26730 3190 26740 3210
rect 26700 3175 26740 3190
rect 26760 3560 26800 3575
rect 26760 3540 26770 3560
rect 26790 3540 26800 3560
rect 26760 3510 26800 3540
rect 26760 3490 26770 3510
rect 26790 3490 26800 3510
rect 26760 3460 26800 3490
rect 26760 3440 26770 3460
rect 26790 3440 26800 3460
rect 26760 3410 26800 3440
rect 26760 3390 26770 3410
rect 26790 3390 26800 3410
rect 26760 3360 26800 3390
rect 26760 3340 26770 3360
rect 26790 3340 26800 3360
rect 26760 3310 26800 3340
rect 26760 3290 26770 3310
rect 26790 3290 26800 3310
rect 26760 3260 26800 3290
rect 26760 3240 26770 3260
rect 26790 3240 26800 3260
rect 26760 3210 26800 3240
rect 26760 3190 26770 3210
rect 26790 3190 26800 3210
rect 26760 3175 26800 3190
rect 26820 3560 26860 3575
rect 26820 3540 26830 3560
rect 26850 3540 26860 3560
rect 26820 3510 26860 3540
rect 26820 3490 26830 3510
rect 26850 3490 26860 3510
rect 26820 3460 26860 3490
rect 26820 3440 26830 3460
rect 26850 3440 26860 3460
rect 26820 3410 26860 3440
rect 26820 3390 26830 3410
rect 26850 3390 26860 3410
rect 26820 3360 26860 3390
rect 26820 3340 26830 3360
rect 26850 3340 26860 3360
rect 26820 3310 26860 3340
rect 26820 3290 26830 3310
rect 26850 3290 26860 3310
rect 26820 3260 26860 3290
rect 26820 3240 26830 3260
rect 26850 3240 26860 3260
rect 26820 3210 26860 3240
rect 26820 3190 26830 3210
rect 26850 3190 26860 3210
rect 26820 3175 26860 3190
rect 26880 3560 26920 3575
rect 26880 3540 26890 3560
rect 26910 3540 26920 3560
rect 26880 3510 26920 3540
rect 26880 3490 26890 3510
rect 26910 3490 26920 3510
rect 26880 3460 26920 3490
rect 26880 3440 26890 3460
rect 26910 3440 26920 3460
rect 26880 3410 26920 3440
rect 26880 3390 26890 3410
rect 26910 3390 26920 3410
rect 26880 3360 26920 3390
rect 26880 3340 26890 3360
rect 26910 3340 26920 3360
rect 26880 3310 26920 3340
rect 26880 3290 26890 3310
rect 26910 3290 26920 3310
rect 26880 3260 26920 3290
rect 26880 3240 26890 3260
rect 26910 3240 26920 3260
rect 26880 3210 26920 3240
rect 26880 3190 26890 3210
rect 26910 3190 26920 3210
rect 26880 3175 26920 3190
rect 26940 3560 26980 3575
rect 26940 3540 26950 3560
rect 26970 3540 26980 3560
rect 26940 3510 26980 3540
rect 26940 3490 26950 3510
rect 26970 3490 26980 3510
rect 26940 3460 26980 3490
rect 26940 3440 26950 3460
rect 26970 3440 26980 3460
rect 26940 3410 26980 3440
rect 26940 3390 26950 3410
rect 26970 3390 26980 3410
rect 26940 3360 26980 3390
rect 26940 3340 26950 3360
rect 26970 3340 26980 3360
rect 26940 3310 26980 3340
rect 26940 3290 26950 3310
rect 26970 3290 26980 3310
rect 26940 3260 26980 3290
rect 26940 3240 26950 3260
rect 26970 3240 26980 3260
rect 26940 3210 26980 3240
rect 26940 3190 26950 3210
rect 26970 3190 26980 3210
rect 26940 3175 26980 3190
rect 27000 3560 27040 3575
rect 27000 3540 27010 3560
rect 27030 3540 27040 3560
rect 27000 3510 27040 3540
rect 27000 3490 27010 3510
rect 27030 3490 27040 3510
rect 27000 3460 27040 3490
rect 27000 3440 27010 3460
rect 27030 3440 27040 3460
rect 27000 3410 27040 3440
rect 27000 3390 27010 3410
rect 27030 3390 27040 3410
rect 27000 3360 27040 3390
rect 27000 3340 27010 3360
rect 27030 3340 27040 3360
rect 27000 3310 27040 3340
rect 27000 3290 27010 3310
rect 27030 3290 27040 3310
rect 27000 3260 27040 3290
rect 27000 3240 27010 3260
rect 27030 3240 27040 3260
rect 27000 3210 27040 3240
rect 27000 3190 27010 3210
rect 27030 3190 27040 3210
rect 27000 3175 27040 3190
rect 27060 3560 27100 3575
rect 27060 3540 27070 3560
rect 27090 3540 27100 3560
rect 27060 3510 27100 3540
rect 27060 3490 27070 3510
rect 27090 3490 27100 3510
rect 27060 3460 27100 3490
rect 27060 3440 27070 3460
rect 27090 3440 27100 3460
rect 27060 3410 27100 3440
rect 27060 3390 27070 3410
rect 27090 3390 27100 3410
rect 27060 3360 27100 3390
rect 27060 3340 27070 3360
rect 27090 3340 27100 3360
rect 27060 3310 27100 3340
rect 27060 3290 27070 3310
rect 27090 3290 27100 3310
rect 27060 3260 27100 3290
rect 27060 3240 27070 3260
rect 27090 3240 27100 3260
rect 27060 3210 27100 3240
rect 27060 3190 27070 3210
rect 27090 3190 27100 3210
rect 27060 3175 27100 3190
rect 27120 3560 27160 3575
rect 27120 3540 27130 3560
rect 27150 3540 27160 3560
rect 27120 3510 27160 3540
rect 27120 3490 27130 3510
rect 27150 3490 27160 3510
rect 27120 3460 27160 3490
rect 27120 3440 27130 3460
rect 27150 3440 27160 3460
rect 27120 3410 27160 3440
rect 27120 3390 27130 3410
rect 27150 3390 27160 3410
rect 27120 3360 27160 3390
rect 27120 3340 27130 3360
rect 27150 3340 27160 3360
rect 27120 3310 27160 3340
rect 27120 3290 27130 3310
rect 27150 3290 27160 3310
rect 27120 3260 27160 3290
rect 27120 3240 27130 3260
rect 27150 3240 27160 3260
rect 27120 3210 27160 3240
rect 27120 3190 27130 3210
rect 27150 3190 27160 3210
rect 27120 3175 27160 3190
rect 27180 3560 27220 3575
rect 27180 3540 27190 3560
rect 27210 3540 27220 3560
rect 27180 3510 27220 3540
rect 27180 3490 27190 3510
rect 27210 3490 27220 3510
rect 27180 3460 27220 3490
rect 27180 3440 27190 3460
rect 27210 3440 27220 3460
rect 27180 3410 27220 3440
rect 27180 3390 27190 3410
rect 27210 3390 27220 3410
rect 27180 3360 27220 3390
rect 27180 3340 27190 3360
rect 27210 3340 27220 3360
rect 27180 3310 27220 3340
rect 27180 3290 27190 3310
rect 27210 3290 27220 3310
rect 27180 3260 27220 3290
rect 27180 3240 27190 3260
rect 27210 3240 27220 3260
rect 27180 3210 27220 3240
rect 27180 3190 27190 3210
rect 27210 3190 27220 3210
rect 27180 3175 27220 3190
rect 27240 3560 27280 3575
rect 27240 3540 27250 3560
rect 27270 3540 27280 3560
rect 27240 3510 27280 3540
rect 27240 3490 27250 3510
rect 27270 3490 27280 3510
rect 27240 3460 27280 3490
rect 27240 3440 27250 3460
rect 27270 3440 27280 3460
rect 27240 3410 27280 3440
rect 27240 3390 27250 3410
rect 27270 3390 27280 3410
rect 27240 3360 27280 3390
rect 27240 3340 27250 3360
rect 27270 3340 27280 3360
rect 27240 3310 27280 3340
rect 27240 3290 27250 3310
rect 27270 3290 27280 3310
rect 27240 3260 27280 3290
rect 27240 3240 27250 3260
rect 27270 3240 27280 3260
rect 27240 3210 27280 3240
rect 27240 3190 27250 3210
rect 27270 3190 27280 3210
rect 27240 3175 27280 3190
rect 27300 3560 27340 3575
rect 27300 3540 27310 3560
rect 27330 3540 27340 3560
rect 27300 3510 27340 3540
rect 27300 3490 27310 3510
rect 27330 3490 27340 3510
rect 27300 3460 27340 3490
rect 27300 3440 27310 3460
rect 27330 3440 27340 3460
rect 27300 3410 27340 3440
rect 27300 3390 27310 3410
rect 27330 3390 27340 3410
rect 27300 3360 27340 3390
rect 27300 3340 27310 3360
rect 27330 3340 27340 3360
rect 27300 3310 27340 3340
rect 27300 3290 27310 3310
rect 27330 3290 27340 3310
rect 27300 3260 27340 3290
rect 27300 3240 27310 3260
rect 27330 3240 27340 3260
rect 27300 3210 27340 3240
rect 27300 3190 27310 3210
rect 27330 3190 27340 3210
rect 27300 3175 27340 3190
rect 27360 3560 27400 3575
rect 27360 3540 27370 3560
rect 27390 3540 27400 3560
rect 27360 3510 27400 3540
rect 27360 3490 27370 3510
rect 27390 3490 27400 3510
rect 27360 3460 27400 3490
rect 27360 3440 27370 3460
rect 27390 3440 27400 3460
rect 27360 3410 27400 3440
rect 27360 3390 27370 3410
rect 27390 3390 27400 3410
rect 27360 3360 27400 3390
rect 27360 3340 27370 3360
rect 27390 3340 27400 3360
rect 27360 3310 27400 3340
rect 27360 3290 27370 3310
rect 27390 3290 27400 3310
rect 27360 3260 27400 3290
rect 27360 3240 27370 3260
rect 27390 3240 27400 3260
rect 27360 3210 27400 3240
rect 27360 3190 27370 3210
rect 27390 3190 27400 3210
rect 27360 3175 27400 3190
rect 27420 3560 27460 3575
rect 27420 3540 27430 3560
rect 27450 3540 27460 3560
rect 27420 3510 27460 3540
rect 27420 3490 27430 3510
rect 27450 3490 27460 3510
rect 27420 3460 27460 3490
rect 27420 3440 27430 3460
rect 27450 3440 27460 3460
rect 27420 3410 27460 3440
rect 27420 3390 27430 3410
rect 27450 3390 27460 3410
rect 27420 3360 27460 3390
rect 27420 3340 27430 3360
rect 27450 3340 27460 3360
rect 27420 3310 27460 3340
rect 27420 3290 27430 3310
rect 27450 3290 27460 3310
rect 27420 3260 27460 3290
rect 27420 3240 27430 3260
rect 27450 3240 27460 3260
rect 27420 3210 27460 3240
rect 27420 3190 27430 3210
rect 27450 3190 27460 3210
rect 27420 3175 27460 3190
rect 27480 3560 27520 3575
rect 27480 3540 27490 3560
rect 27510 3540 27520 3560
rect 27480 3510 27520 3540
rect 27480 3490 27490 3510
rect 27510 3490 27520 3510
rect 27480 3460 27520 3490
rect 27480 3440 27490 3460
rect 27510 3440 27520 3460
rect 27480 3410 27520 3440
rect 27480 3390 27490 3410
rect 27510 3390 27520 3410
rect 27480 3360 27520 3390
rect 27480 3340 27490 3360
rect 27510 3340 27520 3360
rect 27480 3310 27520 3340
rect 27480 3290 27490 3310
rect 27510 3290 27520 3310
rect 27480 3260 27520 3290
rect 27480 3240 27490 3260
rect 27510 3240 27520 3260
rect 27480 3210 27520 3240
rect 27480 3190 27490 3210
rect 27510 3190 27520 3210
rect 27480 3175 27520 3190
rect 27540 3560 27580 3575
rect 27540 3540 27550 3560
rect 27570 3540 27580 3560
rect 27540 3510 27580 3540
rect 27540 3490 27550 3510
rect 27570 3490 27580 3510
rect 27540 3460 27580 3490
rect 27540 3440 27550 3460
rect 27570 3440 27580 3460
rect 27540 3410 27580 3440
rect 27540 3390 27550 3410
rect 27570 3390 27580 3410
rect 27540 3360 27580 3390
rect 27540 3340 27550 3360
rect 27570 3340 27580 3360
rect 27540 3310 27580 3340
rect 27540 3290 27550 3310
rect 27570 3290 27580 3310
rect 27540 3260 27580 3290
rect 27540 3240 27550 3260
rect 27570 3240 27580 3260
rect 27540 3210 27580 3240
rect 27540 3190 27550 3210
rect 27570 3190 27580 3210
rect 27540 3175 27580 3190
rect 27890 3225 27930 3240
rect 27890 3205 27900 3225
rect 27920 3205 27930 3225
rect 27890 3175 27930 3205
rect 27890 3155 27900 3175
rect 27920 3155 27930 3175
rect 27890 3125 27930 3155
rect 27890 3105 27900 3125
rect 27920 3105 27930 3125
rect 27890 3075 27930 3105
rect 27890 3055 27900 3075
rect 27920 3055 27930 3075
rect 27890 3025 27930 3055
rect 27890 3005 27900 3025
rect 27920 3005 27930 3025
rect 27890 2975 27930 3005
rect 27890 2955 27900 2975
rect 27920 2955 27930 2975
rect 27890 2940 27930 2955
rect 27945 3225 27985 3240
rect 27945 3205 27955 3225
rect 27975 3205 27985 3225
rect 27945 3175 27985 3205
rect 27945 3155 27955 3175
rect 27975 3155 27985 3175
rect 27945 3125 27985 3155
rect 27945 3105 27955 3125
rect 27975 3105 27985 3125
rect 27945 3075 27985 3105
rect 27945 3055 27955 3075
rect 27975 3055 27985 3075
rect 27945 3025 27985 3055
rect 27945 3005 27955 3025
rect 27975 3005 27985 3025
rect 27945 2975 27985 3005
rect 27945 2955 27955 2975
rect 27975 2955 27985 2975
rect 27945 2940 27985 2955
rect 28000 3225 28040 3240
rect 28000 3205 28010 3225
rect 28030 3205 28040 3225
rect 28000 3175 28040 3205
rect 28000 3155 28010 3175
rect 28030 3155 28040 3175
rect 28000 3125 28040 3155
rect 28000 3105 28010 3125
rect 28030 3105 28040 3125
rect 28000 3075 28040 3105
rect 28000 3055 28010 3075
rect 28030 3055 28040 3075
rect 28000 3025 28040 3055
rect 28000 3005 28010 3025
rect 28030 3005 28040 3025
rect 28000 2975 28040 3005
rect 28000 2955 28010 2975
rect 28030 2955 28040 2975
rect 28000 2940 28040 2955
rect 28055 3225 28095 3240
rect 28055 3205 28065 3225
rect 28085 3205 28095 3225
rect 28055 3175 28095 3205
rect 28055 3155 28065 3175
rect 28085 3155 28095 3175
rect 28055 3125 28095 3155
rect 28055 3105 28065 3125
rect 28085 3105 28095 3125
rect 28055 3075 28095 3105
rect 28055 3055 28065 3075
rect 28085 3055 28095 3075
rect 28055 3025 28095 3055
rect 28055 3005 28065 3025
rect 28085 3005 28095 3025
rect 28055 2975 28095 3005
rect 28055 2955 28065 2975
rect 28085 2955 28095 2975
rect 28055 2940 28095 2955
rect 28110 3225 28150 3240
rect 28110 3205 28120 3225
rect 28140 3205 28150 3225
rect 28110 3175 28150 3205
rect 28110 3155 28120 3175
rect 28140 3155 28150 3175
rect 28110 3125 28150 3155
rect 28110 3105 28120 3125
rect 28140 3105 28150 3125
rect 28110 3075 28150 3105
rect 28110 3055 28120 3075
rect 28140 3055 28150 3075
rect 28110 3025 28150 3055
rect 28110 3005 28120 3025
rect 28140 3005 28150 3025
rect 28110 2975 28150 3005
rect 28110 2955 28120 2975
rect 28140 2955 28150 2975
rect 28110 2940 28150 2955
rect 28165 3225 28205 3240
rect 28165 3205 28175 3225
rect 28195 3205 28205 3225
rect 28165 3175 28205 3205
rect 28165 3155 28175 3175
rect 28195 3155 28205 3175
rect 28165 3125 28205 3155
rect 28165 3105 28175 3125
rect 28195 3105 28205 3125
rect 28165 3075 28205 3105
rect 28165 3055 28175 3075
rect 28195 3055 28205 3075
rect 28165 3025 28205 3055
rect 28165 3005 28175 3025
rect 28195 3005 28205 3025
rect 28165 2975 28205 3005
rect 28165 2955 28175 2975
rect 28195 2955 28205 2975
rect 28165 2940 28205 2955
rect 28220 3225 28260 3240
rect 28220 3205 28230 3225
rect 28250 3205 28260 3225
rect 28220 3175 28260 3205
rect 28220 3155 28230 3175
rect 28250 3155 28260 3175
rect 28220 3125 28260 3155
rect 28220 3105 28230 3125
rect 28250 3105 28260 3125
rect 28220 3075 28260 3105
rect 28220 3055 28230 3075
rect 28250 3055 28260 3075
rect 28220 3025 28260 3055
rect 28220 3005 28230 3025
rect 28250 3005 28260 3025
rect 28220 2975 28260 3005
rect 28220 2955 28230 2975
rect 28250 2955 28260 2975
rect 28220 2940 28260 2955
rect 28275 3225 28315 3240
rect 28275 3205 28285 3225
rect 28305 3205 28315 3225
rect 28275 3175 28315 3205
rect 28275 3155 28285 3175
rect 28305 3155 28315 3175
rect 28275 3125 28315 3155
rect 28275 3105 28285 3125
rect 28305 3105 28315 3125
rect 28275 3075 28315 3105
rect 28275 3055 28285 3075
rect 28305 3055 28315 3075
rect 28275 3025 28315 3055
rect 28275 3005 28285 3025
rect 28305 3005 28315 3025
rect 28275 2975 28315 3005
rect 28275 2955 28285 2975
rect 28305 2955 28315 2975
rect 28275 2940 28315 2955
rect 28330 3225 28370 3240
rect 28330 3205 28340 3225
rect 28360 3205 28370 3225
rect 28330 3175 28370 3205
rect 28330 3155 28340 3175
rect 28360 3155 28370 3175
rect 28330 3125 28370 3155
rect 28330 3105 28340 3125
rect 28360 3105 28370 3125
rect 28330 3075 28370 3105
rect 28330 3055 28340 3075
rect 28360 3055 28370 3075
rect 28330 3025 28370 3055
rect 28330 3005 28340 3025
rect 28360 3005 28370 3025
rect 28330 2975 28370 3005
rect 28330 2955 28340 2975
rect 28360 2955 28370 2975
rect 28330 2940 28370 2955
rect 28385 3225 28425 3240
rect 28385 3205 28395 3225
rect 28415 3205 28425 3225
rect 28385 3175 28425 3205
rect 28385 3155 28395 3175
rect 28415 3155 28425 3175
rect 28385 3125 28425 3155
rect 28385 3105 28395 3125
rect 28415 3105 28425 3125
rect 28385 3075 28425 3105
rect 28385 3055 28395 3075
rect 28415 3055 28425 3075
rect 28385 3025 28425 3055
rect 28385 3005 28395 3025
rect 28415 3005 28425 3025
rect 28385 2975 28425 3005
rect 28385 2955 28395 2975
rect 28415 2955 28425 2975
rect 28385 2940 28425 2955
rect 28440 3225 28480 3240
rect 28440 3205 28450 3225
rect 28470 3205 28480 3225
rect 28440 3175 28480 3205
rect 28440 3155 28450 3175
rect 28470 3155 28480 3175
rect 28440 3125 28480 3155
rect 28440 3105 28450 3125
rect 28470 3105 28480 3125
rect 28440 3075 28480 3105
rect 28440 3055 28450 3075
rect 28470 3055 28480 3075
rect 28440 3025 28480 3055
rect 28440 3005 28450 3025
rect 28470 3005 28480 3025
rect 28440 2975 28480 3005
rect 28440 2955 28450 2975
rect 28470 2955 28480 2975
rect 28440 2940 28480 2955
rect 28495 3225 28535 3240
rect 28495 3205 28505 3225
rect 28525 3205 28535 3225
rect 28495 3175 28535 3205
rect 28495 3155 28505 3175
rect 28525 3155 28535 3175
rect 28495 3125 28535 3155
rect 28495 3105 28505 3125
rect 28525 3105 28535 3125
rect 28495 3075 28535 3105
rect 28495 3055 28505 3075
rect 28525 3055 28535 3075
rect 28495 3025 28535 3055
rect 28495 3005 28505 3025
rect 28525 3005 28535 3025
rect 28495 2975 28535 3005
rect 28495 2955 28505 2975
rect 28525 2955 28535 2975
rect 28495 2940 28535 2955
rect 28550 3225 28590 3240
rect 28550 3205 28560 3225
rect 28580 3205 28590 3225
rect 28550 3175 28590 3205
rect 28550 3155 28560 3175
rect 28580 3155 28590 3175
rect 28550 3125 28590 3155
rect 28550 3105 28560 3125
rect 28580 3105 28590 3125
rect 28550 3075 28590 3105
rect 28550 3055 28560 3075
rect 28580 3055 28590 3075
rect 28550 3025 28590 3055
rect 28550 3005 28560 3025
rect 28580 3005 28590 3025
rect 28550 2975 28590 3005
rect 28550 2955 28560 2975
rect 28580 2955 28590 2975
rect 28550 2940 28590 2955
rect 28605 3225 28645 3240
rect 28605 3205 28615 3225
rect 28635 3205 28645 3225
rect 28605 3175 28645 3205
rect 28605 3155 28615 3175
rect 28635 3155 28645 3175
rect 28605 3125 28645 3155
rect 28605 3105 28615 3125
rect 28635 3105 28645 3125
rect 28605 3075 28645 3105
rect 28605 3055 28615 3075
rect 28635 3055 28645 3075
rect 28605 3025 28645 3055
rect 28605 3005 28615 3025
rect 28635 3005 28645 3025
rect 28605 2975 28645 3005
rect 28605 2955 28615 2975
rect 28635 2955 28645 2975
rect 28605 2940 28645 2955
rect 28660 3225 28700 3240
rect 28660 3205 28670 3225
rect 28690 3205 28700 3225
rect 28660 3175 28700 3205
rect 28660 3155 28670 3175
rect 28690 3155 28700 3175
rect 28660 3125 28700 3155
rect 28660 3105 28670 3125
rect 28690 3105 28700 3125
rect 28660 3075 28700 3105
rect 28660 3055 28670 3075
rect 28690 3055 28700 3075
rect 28660 3025 28700 3055
rect 28660 3005 28670 3025
rect 28690 3005 28700 3025
rect 28660 2975 28700 3005
rect 28660 2955 28670 2975
rect 28690 2955 28700 2975
rect 28660 2940 28700 2955
rect 28715 3225 28755 3240
rect 28715 3205 28725 3225
rect 28745 3205 28755 3225
rect 28715 3175 28755 3205
rect 28715 3155 28725 3175
rect 28745 3155 28755 3175
rect 28715 3125 28755 3155
rect 28715 3105 28725 3125
rect 28745 3105 28755 3125
rect 28715 3075 28755 3105
rect 28715 3055 28725 3075
rect 28745 3055 28755 3075
rect 28715 3025 28755 3055
rect 28715 3005 28725 3025
rect 28745 3005 28755 3025
rect 28715 2975 28755 3005
rect 28715 2955 28725 2975
rect 28745 2955 28755 2975
rect 28715 2940 28755 2955
rect 28770 3225 28810 3240
rect 28770 3205 28780 3225
rect 28800 3205 28810 3225
rect 28770 3175 28810 3205
rect 28770 3155 28780 3175
rect 28800 3155 28810 3175
rect 28770 3125 28810 3155
rect 28770 3105 28780 3125
rect 28800 3105 28810 3125
rect 28770 3075 28810 3105
rect 28770 3055 28780 3075
rect 28800 3055 28810 3075
rect 28770 3025 28810 3055
rect 28770 3005 28780 3025
rect 28800 3005 28810 3025
rect 28770 2975 28810 3005
rect 28770 2955 28780 2975
rect 28800 2955 28810 2975
rect 28770 2940 28810 2955
rect 28825 3225 28865 3240
rect 28825 3205 28835 3225
rect 28855 3205 28865 3225
rect 28825 3175 28865 3205
rect 28825 3155 28835 3175
rect 28855 3155 28865 3175
rect 28825 3125 28865 3155
rect 28825 3105 28835 3125
rect 28855 3105 28865 3125
rect 28825 3075 28865 3105
rect 28825 3055 28835 3075
rect 28855 3055 28865 3075
rect 28825 3025 28865 3055
rect 28825 3005 28835 3025
rect 28855 3005 28865 3025
rect 28825 2975 28865 3005
rect 28825 2955 28835 2975
rect 28855 2955 28865 2975
rect 28825 2940 28865 2955
rect 28880 3225 28920 3240
rect 28880 3205 28890 3225
rect 28910 3205 28920 3225
rect 28880 3175 28920 3205
rect 28880 3155 28890 3175
rect 28910 3155 28920 3175
rect 28880 3125 28920 3155
rect 28880 3105 28890 3125
rect 28910 3105 28920 3125
rect 28880 3075 28920 3105
rect 28880 3055 28890 3075
rect 28910 3055 28920 3075
rect 28880 3025 28920 3055
rect 28880 3005 28890 3025
rect 28910 3005 28920 3025
rect 28880 2975 28920 3005
rect 28880 2955 28890 2975
rect 28910 2955 28920 2975
rect 28880 2940 28920 2955
rect 28935 3225 28975 3240
rect 28935 3205 28945 3225
rect 28965 3205 28975 3225
rect 28935 3175 28975 3205
rect 28935 3155 28945 3175
rect 28965 3155 28975 3175
rect 28935 3125 28975 3155
rect 28935 3105 28945 3125
rect 28965 3105 28975 3125
rect 28935 3075 28975 3105
rect 28935 3055 28945 3075
rect 28965 3055 28975 3075
rect 28935 3025 28975 3055
rect 28935 3005 28945 3025
rect 28965 3005 28975 3025
rect 28935 2975 28975 3005
rect 28935 2955 28945 2975
rect 28965 2955 28975 2975
rect 28935 2940 28975 2955
rect 28990 3225 29030 3240
rect 28990 3205 29000 3225
rect 29020 3205 29030 3225
rect 28990 3175 29030 3205
rect 28990 3155 29000 3175
rect 29020 3155 29030 3175
rect 28990 3125 29030 3155
rect 28990 3105 29000 3125
rect 29020 3105 29030 3125
rect 28990 3075 29030 3105
rect 28990 3055 29000 3075
rect 29020 3055 29030 3075
rect 28990 3025 29030 3055
rect 28990 3005 29000 3025
rect 29020 3005 29030 3025
rect 28990 2975 29030 3005
rect 28990 2955 29000 2975
rect 29020 2955 29030 2975
rect 28990 2940 29030 2955
rect 29045 3225 29085 3240
rect 29045 3205 29055 3225
rect 29075 3205 29085 3225
rect 29045 3175 29085 3205
rect 29045 3155 29055 3175
rect 29075 3155 29085 3175
rect 29045 3125 29085 3155
rect 29045 3105 29055 3125
rect 29075 3105 29085 3125
rect 29045 3075 29085 3105
rect 29045 3055 29055 3075
rect 29075 3055 29085 3075
rect 29045 3025 29085 3055
rect 29045 3005 29055 3025
rect 29075 3005 29085 3025
rect 29045 2975 29085 3005
rect 29045 2955 29055 2975
rect 29075 2955 29085 2975
rect 29045 2940 29085 2955
rect 29100 3225 29140 3240
rect 29100 3205 29110 3225
rect 29130 3205 29140 3225
rect 29100 3175 29140 3205
rect 29100 3155 29110 3175
rect 29130 3155 29140 3175
rect 29100 3125 29140 3155
rect 29100 3105 29110 3125
rect 29130 3105 29140 3125
rect 29100 3075 29140 3105
rect 29100 3055 29110 3075
rect 29130 3055 29140 3075
rect 29100 3025 29140 3055
rect 29100 3005 29110 3025
rect 29130 3005 29140 3025
rect 29100 2975 29140 3005
rect 29100 2955 29110 2975
rect 29130 2955 29140 2975
rect 29100 2940 29140 2955
rect 11220 2880 11260 2895
rect 11220 2860 11230 2880
rect 11250 2860 11260 2880
rect 11220 2830 11260 2860
rect 11220 2810 11230 2830
rect 11250 2810 11260 2830
rect 11220 2780 11260 2810
rect 11220 2760 11230 2780
rect 11250 2760 11260 2780
rect 11220 2730 11260 2760
rect 11220 2710 11230 2730
rect 11250 2710 11260 2730
rect 11220 2680 11260 2710
rect 11220 2660 11230 2680
rect 11250 2660 11260 2680
rect 10155 2640 10195 2655
rect 10155 2620 10165 2640
rect 10185 2620 10195 2640
rect 10155 2590 10195 2620
rect 10155 2570 10165 2590
rect 10185 2570 10195 2590
rect 10155 2540 10195 2570
rect 10155 2520 10165 2540
rect 10185 2520 10195 2540
rect 10155 2490 10195 2520
rect 10155 2470 10165 2490
rect 10185 2470 10195 2490
rect 10155 2455 10195 2470
rect 10210 2640 10250 2655
rect 10210 2620 10220 2640
rect 10240 2620 10250 2640
rect 10210 2590 10250 2620
rect 10210 2570 10220 2590
rect 10240 2570 10250 2590
rect 10210 2540 10250 2570
rect 10210 2520 10220 2540
rect 10240 2520 10250 2540
rect 10210 2490 10250 2520
rect 10210 2470 10220 2490
rect 10240 2470 10250 2490
rect 10210 2455 10250 2470
rect 10265 2640 10305 2655
rect 10265 2620 10275 2640
rect 10295 2620 10305 2640
rect 10265 2590 10305 2620
rect 10265 2570 10275 2590
rect 10295 2570 10305 2590
rect 10265 2540 10305 2570
rect 10265 2520 10275 2540
rect 10295 2520 10305 2540
rect 10265 2490 10305 2520
rect 10265 2470 10275 2490
rect 10295 2470 10305 2490
rect 10265 2455 10305 2470
rect 10320 2640 10360 2655
rect 10320 2620 10330 2640
rect 10350 2620 10360 2640
rect 10320 2590 10360 2620
rect 10320 2570 10330 2590
rect 10350 2570 10360 2590
rect 10320 2540 10360 2570
rect 10320 2520 10330 2540
rect 10350 2520 10360 2540
rect 10320 2490 10360 2520
rect 10320 2470 10330 2490
rect 10350 2470 10360 2490
rect 10320 2455 10360 2470
rect 10375 2640 10415 2655
rect 10375 2620 10385 2640
rect 10405 2620 10415 2640
rect 10375 2590 10415 2620
rect 10375 2570 10385 2590
rect 10405 2570 10415 2590
rect 10375 2540 10415 2570
rect 10375 2520 10385 2540
rect 10405 2520 10415 2540
rect 10375 2490 10415 2520
rect 10375 2470 10385 2490
rect 10405 2470 10415 2490
rect 10375 2455 10415 2470
rect 10430 2640 10470 2655
rect 10430 2620 10440 2640
rect 10460 2620 10470 2640
rect 10430 2590 10470 2620
rect 10430 2570 10440 2590
rect 10460 2570 10470 2590
rect 10430 2540 10470 2570
rect 10430 2520 10440 2540
rect 10460 2520 10470 2540
rect 10430 2490 10470 2520
rect 10430 2470 10440 2490
rect 10460 2470 10470 2490
rect 10430 2455 10470 2470
rect 10485 2640 10525 2655
rect 10485 2620 10495 2640
rect 10515 2620 10525 2640
rect 10485 2590 10525 2620
rect 10485 2570 10495 2590
rect 10515 2570 10525 2590
rect 10485 2540 10525 2570
rect 10485 2520 10495 2540
rect 10515 2520 10525 2540
rect 10485 2490 10525 2520
rect 10485 2470 10495 2490
rect 10515 2470 10525 2490
rect 10485 2455 10525 2470
rect 10540 2640 10580 2655
rect 10540 2620 10550 2640
rect 10570 2620 10580 2640
rect 10540 2590 10580 2620
rect 10540 2570 10550 2590
rect 10570 2570 10580 2590
rect 10540 2540 10580 2570
rect 10540 2520 10550 2540
rect 10570 2520 10580 2540
rect 10540 2490 10580 2520
rect 10540 2470 10550 2490
rect 10570 2470 10580 2490
rect 10540 2455 10580 2470
rect 10595 2640 10635 2655
rect 10595 2620 10605 2640
rect 10625 2620 10635 2640
rect 10595 2590 10635 2620
rect 10595 2570 10605 2590
rect 10625 2570 10635 2590
rect 10595 2540 10635 2570
rect 10595 2520 10605 2540
rect 10625 2520 10635 2540
rect 10595 2490 10635 2520
rect 10595 2470 10605 2490
rect 10625 2470 10635 2490
rect 10595 2455 10635 2470
rect 10650 2640 10690 2655
rect 10650 2620 10660 2640
rect 10680 2620 10690 2640
rect 10650 2590 10690 2620
rect 10650 2570 10660 2590
rect 10680 2570 10690 2590
rect 10650 2540 10690 2570
rect 10650 2520 10660 2540
rect 10680 2520 10690 2540
rect 10650 2490 10690 2520
rect 10650 2470 10660 2490
rect 10680 2470 10690 2490
rect 10650 2455 10690 2470
rect 10705 2640 10745 2655
rect 10705 2620 10715 2640
rect 10735 2620 10745 2640
rect 10705 2590 10745 2620
rect 10705 2570 10715 2590
rect 10735 2570 10745 2590
rect 10705 2540 10745 2570
rect 10705 2520 10715 2540
rect 10735 2520 10745 2540
rect 10705 2490 10745 2520
rect 10705 2470 10715 2490
rect 10735 2470 10745 2490
rect 10705 2455 10745 2470
rect 10760 2640 10800 2655
rect 10760 2620 10770 2640
rect 10790 2620 10800 2640
rect 10760 2590 10800 2620
rect 10760 2570 10770 2590
rect 10790 2570 10800 2590
rect 10760 2540 10800 2570
rect 10760 2520 10770 2540
rect 10790 2520 10800 2540
rect 10760 2490 10800 2520
rect 10760 2470 10770 2490
rect 10790 2470 10800 2490
rect 10760 2455 10800 2470
rect 10815 2640 10855 2655
rect 10815 2620 10825 2640
rect 10845 2620 10855 2640
rect 10815 2590 10855 2620
rect 10815 2570 10825 2590
rect 10845 2570 10855 2590
rect 10815 2540 10855 2570
rect 10815 2520 10825 2540
rect 10845 2520 10855 2540
rect 10815 2490 10855 2520
rect 11220 2630 11260 2660
rect 11220 2610 11230 2630
rect 11250 2610 11260 2630
rect 11220 2580 11260 2610
rect 11220 2560 11230 2580
rect 11250 2560 11260 2580
rect 11220 2530 11260 2560
rect 11220 2510 11230 2530
rect 11250 2510 11260 2530
rect 11220 2495 11260 2510
rect 11280 2880 11320 2895
rect 11280 2860 11290 2880
rect 11310 2860 11320 2880
rect 11280 2830 11320 2860
rect 11280 2810 11290 2830
rect 11310 2810 11320 2830
rect 11280 2780 11320 2810
rect 11280 2760 11290 2780
rect 11310 2760 11320 2780
rect 11280 2730 11320 2760
rect 11280 2710 11290 2730
rect 11310 2710 11320 2730
rect 11280 2680 11320 2710
rect 11280 2660 11290 2680
rect 11310 2660 11320 2680
rect 11280 2630 11320 2660
rect 11280 2610 11290 2630
rect 11310 2610 11320 2630
rect 11280 2580 11320 2610
rect 11280 2560 11290 2580
rect 11310 2560 11320 2580
rect 11280 2530 11320 2560
rect 11280 2510 11290 2530
rect 11310 2510 11320 2530
rect 11280 2495 11320 2510
rect 11340 2880 11380 2895
rect 11340 2860 11350 2880
rect 11370 2860 11380 2880
rect 11340 2830 11380 2860
rect 11340 2810 11350 2830
rect 11370 2810 11380 2830
rect 11340 2780 11380 2810
rect 11340 2760 11350 2780
rect 11370 2760 11380 2780
rect 11340 2730 11380 2760
rect 11340 2710 11350 2730
rect 11370 2710 11380 2730
rect 11340 2680 11380 2710
rect 11340 2660 11350 2680
rect 11370 2660 11380 2680
rect 11340 2630 11380 2660
rect 11340 2610 11350 2630
rect 11370 2610 11380 2630
rect 11340 2580 11380 2610
rect 11340 2560 11350 2580
rect 11370 2560 11380 2580
rect 11340 2530 11380 2560
rect 11340 2510 11350 2530
rect 11370 2510 11380 2530
rect 11340 2495 11380 2510
rect 11400 2880 11440 2895
rect 11400 2860 11410 2880
rect 11430 2860 11440 2880
rect 11400 2830 11440 2860
rect 11400 2810 11410 2830
rect 11430 2810 11440 2830
rect 11400 2780 11440 2810
rect 11400 2760 11410 2780
rect 11430 2760 11440 2780
rect 11400 2730 11440 2760
rect 11400 2710 11410 2730
rect 11430 2710 11440 2730
rect 11400 2680 11440 2710
rect 11400 2660 11410 2680
rect 11430 2660 11440 2680
rect 11400 2630 11440 2660
rect 11400 2610 11410 2630
rect 11430 2610 11440 2630
rect 11400 2580 11440 2610
rect 11400 2560 11410 2580
rect 11430 2560 11440 2580
rect 11400 2530 11440 2560
rect 11400 2510 11410 2530
rect 11430 2510 11440 2530
rect 11400 2495 11440 2510
rect 11460 2880 11500 2895
rect 11460 2860 11470 2880
rect 11490 2860 11500 2880
rect 11460 2830 11500 2860
rect 11460 2810 11470 2830
rect 11490 2810 11500 2830
rect 11460 2780 11500 2810
rect 11460 2760 11470 2780
rect 11490 2760 11500 2780
rect 11460 2730 11500 2760
rect 11460 2710 11470 2730
rect 11490 2710 11500 2730
rect 11460 2680 11500 2710
rect 11460 2660 11470 2680
rect 11490 2660 11500 2680
rect 11460 2630 11500 2660
rect 11460 2610 11470 2630
rect 11490 2610 11500 2630
rect 11460 2580 11500 2610
rect 11460 2560 11470 2580
rect 11490 2560 11500 2580
rect 11460 2530 11500 2560
rect 11460 2510 11470 2530
rect 11490 2510 11500 2530
rect 11460 2495 11500 2510
rect 11520 2880 11560 2895
rect 11520 2860 11530 2880
rect 11550 2860 11560 2880
rect 11520 2830 11560 2860
rect 11520 2810 11530 2830
rect 11550 2810 11560 2830
rect 11520 2780 11560 2810
rect 11520 2760 11530 2780
rect 11550 2760 11560 2780
rect 11520 2730 11560 2760
rect 11520 2710 11530 2730
rect 11550 2710 11560 2730
rect 11520 2680 11560 2710
rect 11520 2660 11530 2680
rect 11550 2660 11560 2680
rect 11520 2630 11560 2660
rect 11520 2610 11530 2630
rect 11550 2610 11560 2630
rect 11520 2580 11560 2610
rect 11520 2560 11530 2580
rect 11550 2560 11560 2580
rect 11520 2530 11560 2560
rect 11520 2510 11530 2530
rect 11550 2510 11560 2530
rect 11520 2495 11560 2510
rect 11580 2880 11620 2895
rect 11580 2860 11590 2880
rect 11610 2860 11620 2880
rect 11580 2830 11620 2860
rect 11580 2810 11590 2830
rect 11610 2810 11620 2830
rect 11580 2780 11620 2810
rect 11580 2760 11590 2780
rect 11610 2760 11620 2780
rect 11580 2730 11620 2760
rect 11580 2710 11590 2730
rect 11610 2710 11620 2730
rect 11580 2680 11620 2710
rect 11580 2660 11590 2680
rect 11610 2660 11620 2680
rect 11580 2630 11620 2660
rect 11580 2610 11590 2630
rect 11610 2610 11620 2630
rect 11580 2580 11620 2610
rect 11580 2560 11590 2580
rect 11610 2560 11620 2580
rect 11580 2530 11620 2560
rect 11580 2510 11590 2530
rect 11610 2510 11620 2530
rect 11580 2495 11620 2510
rect 11640 2880 11680 2895
rect 11640 2860 11650 2880
rect 11670 2860 11680 2880
rect 11640 2830 11680 2860
rect 11640 2810 11650 2830
rect 11670 2810 11680 2830
rect 11640 2780 11680 2810
rect 11640 2760 11650 2780
rect 11670 2760 11680 2780
rect 11640 2730 11680 2760
rect 11640 2710 11650 2730
rect 11670 2710 11680 2730
rect 11640 2680 11680 2710
rect 11640 2660 11650 2680
rect 11670 2660 11680 2680
rect 11640 2630 11680 2660
rect 11640 2610 11650 2630
rect 11670 2610 11680 2630
rect 11640 2580 11680 2610
rect 11640 2560 11650 2580
rect 11670 2560 11680 2580
rect 11640 2530 11680 2560
rect 11640 2510 11650 2530
rect 11670 2510 11680 2530
rect 11640 2495 11680 2510
rect 11700 2880 11740 2895
rect 11700 2860 11710 2880
rect 11730 2860 11740 2880
rect 11700 2830 11740 2860
rect 11700 2810 11710 2830
rect 11730 2810 11740 2830
rect 11700 2780 11740 2810
rect 11700 2760 11710 2780
rect 11730 2760 11740 2780
rect 11700 2730 11740 2760
rect 11700 2710 11710 2730
rect 11730 2710 11740 2730
rect 11700 2680 11740 2710
rect 11700 2660 11710 2680
rect 11730 2660 11740 2680
rect 11700 2630 11740 2660
rect 11700 2610 11710 2630
rect 11730 2610 11740 2630
rect 11700 2580 11740 2610
rect 11700 2560 11710 2580
rect 11730 2560 11740 2580
rect 11700 2530 11740 2560
rect 11700 2510 11710 2530
rect 11730 2510 11740 2530
rect 11700 2495 11740 2510
rect 11760 2880 11800 2895
rect 11760 2860 11770 2880
rect 11790 2860 11800 2880
rect 11760 2830 11800 2860
rect 11760 2810 11770 2830
rect 11790 2810 11800 2830
rect 11760 2780 11800 2810
rect 11760 2760 11770 2780
rect 11790 2760 11800 2780
rect 11760 2730 11800 2760
rect 11760 2710 11770 2730
rect 11790 2710 11800 2730
rect 11760 2680 11800 2710
rect 11760 2660 11770 2680
rect 11790 2660 11800 2680
rect 11760 2630 11800 2660
rect 11760 2610 11770 2630
rect 11790 2610 11800 2630
rect 11760 2580 11800 2610
rect 11760 2560 11770 2580
rect 11790 2560 11800 2580
rect 11760 2530 11800 2560
rect 11760 2510 11770 2530
rect 11790 2510 11800 2530
rect 11760 2495 11800 2510
rect 11820 2880 11860 2895
rect 11820 2860 11830 2880
rect 11850 2860 11860 2880
rect 11820 2830 11860 2860
rect 11820 2810 11830 2830
rect 11850 2810 11860 2830
rect 11820 2780 11860 2810
rect 11820 2760 11830 2780
rect 11850 2760 11860 2780
rect 11820 2730 11860 2760
rect 11820 2710 11830 2730
rect 11850 2710 11860 2730
rect 11820 2680 11860 2710
rect 11820 2660 11830 2680
rect 11850 2660 11860 2680
rect 11820 2630 11860 2660
rect 11820 2610 11830 2630
rect 11850 2610 11860 2630
rect 11820 2580 11860 2610
rect 11820 2560 11830 2580
rect 11850 2560 11860 2580
rect 11820 2530 11860 2560
rect 11820 2510 11830 2530
rect 11850 2510 11860 2530
rect 11820 2495 11860 2510
rect 11880 2880 11920 2895
rect 11880 2860 11890 2880
rect 11910 2860 11920 2880
rect 11880 2830 11920 2860
rect 11880 2810 11890 2830
rect 11910 2810 11920 2830
rect 11880 2780 11920 2810
rect 11880 2760 11890 2780
rect 11910 2760 11920 2780
rect 11880 2730 11920 2760
rect 11880 2710 11890 2730
rect 11910 2710 11920 2730
rect 11880 2680 11920 2710
rect 11880 2660 11890 2680
rect 11910 2660 11920 2680
rect 11880 2630 11920 2660
rect 11880 2610 11890 2630
rect 11910 2610 11920 2630
rect 11880 2580 11920 2610
rect 11880 2560 11890 2580
rect 11910 2560 11920 2580
rect 11880 2530 11920 2560
rect 11880 2510 11890 2530
rect 11910 2510 11920 2530
rect 11880 2495 11920 2510
rect 11940 2880 11980 2895
rect 11940 2860 11950 2880
rect 11970 2860 11980 2880
rect 11940 2830 11980 2860
rect 11940 2810 11950 2830
rect 11970 2810 11980 2830
rect 11940 2780 11980 2810
rect 11940 2760 11950 2780
rect 11970 2760 11980 2780
rect 11940 2730 11980 2760
rect 11940 2710 11950 2730
rect 11970 2710 11980 2730
rect 11940 2680 11980 2710
rect 11940 2660 11950 2680
rect 11970 2660 11980 2680
rect 11940 2630 11980 2660
rect 11940 2610 11950 2630
rect 11970 2610 11980 2630
rect 11940 2580 11980 2610
rect 11940 2560 11950 2580
rect 11970 2560 11980 2580
rect 11940 2530 11980 2560
rect 11940 2510 11950 2530
rect 11970 2510 11980 2530
rect 11940 2495 11980 2510
rect 12000 2880 12040 2895
rect 12000 2860 12010 2880
rect 12030 2860 12040 2880
rect 12000 2830 12040 2860
rect 12000 2810 12010 2830
rect 12030 2810 12040 2830
rect 12000 2780 12040 2810
rect 12000 2760 12010 2780
rect 12030 2760 12040 2780
rect 12000 2730 12040 2760
rect 12000 2710 12010 2730
rect 12030 2710 12040 2730
rect 12000 2680 12040 2710
rect 12000 2660 12010 2680
rect 12030 2660 12040 2680
rect 12000 2630 12040 2660
rect 12000 2610 12010 2630
rect 12030 2610 12040 2630
rect 12000 2580 12040 2610
rect 12000 2560 12010 2580
rect 12030 2560 12040 2580
rect 12000 2530 12040 2560
rect 12000 2510 12010 2530
rect 12030 2510 12040 2530
rect 12000 2495 12040 2510
rect 12060 2880 12100 2895
rect 12060 2860 12070 2880
rect 12090 2860 12100 2880
rect 12060 2830 12100 2860
rect 12060 2810 12070 2830
rect 12090 2810 12100 2830
rect 12060 2780 12100 2810
rect 12060 2760 12070 2780
rect 12090 2760 12100 2780
rect 12060 2730 12100 2760
rect 12060 2710 12070 2730
rect 12090 2710 12100 2730
rect 12060 2680 12100 2710
rect 12060 2660 12070 2680
rect 12090 2660 12100 2680
rect 12060 2630 12100 2660
rect 12060 2610 12070 2630
rect 12090 2610 12100 2630
rect 12060 2580 12100 2610
rect 12060 2560 12070 2580
rect 12090 2560 12100 2580
rect 12060 2530 12100 2560
rect 12060 2510 12070 2530
rect 12090 2510 12100 2530
rect 12060 2495 12100 2510
rect 12120 2880 12160 2895
rect 12120 2860 12130 2880
rect 12150 2860 12160 2880
rect 12120 2830 12160 2860
rect 12120 2810 12130 2830
rect 12150 2810 12160 2830
rect 12120 2780 12160 2810
rect 12120 2760 12130 2780
rect 12150 2760 12160 2780
rect 12120 2730 12160 2760
rect 12120 2710 12130 2730
rect 12150 2710 12160 2730
rect 12120 2680 12160 2710
rect 12120 2660 12130 2680
rect 12150 2660 12160 2680
rect 12120 2630 12160 2660
rect 12120 2610 12130 2630
rect 12150 2610 12160 2630
rect 12120 2580 12160 2610
rect 12120 2560 12130 2580
rect 12150 2560 12160 2580
rect 12120 2530 12160 2560
rect 12120 2510 12130 2530
rect 12150 2510 12160 2530
rect 12120 2495 12160 2510
rect 12180 2880 12220 2895
rect 12180 2860 12190 2880
rect 12210 2860 12220 2880
rect 12180 2830 12220 2860
rect 12180 2810 12190 2830
rect 12210 2810 12220 2830
rect 12180 2780 12220 2810
rect 12180 2760 12190 2780
rect 12210 2760 12220 2780
rect 12180 2730 12220 2760
rect 12180 2710 12190 2730
rect 12210 2710 12220 2730
rect 12180 2680 12220 2710
rect 12180 2660 12190 2680
rect 12210 2660 12220 2680
rect 12180 2630 12220 2660
rect 12180 2610 12190 2630
rect 12210 2610 12220 2630
rect 12180 2580 12220 2610
rect 12180 2560 12190 2580
rect 12210 2560 12220 2580
rect 12180 2530 12220 2560
rect 12180 2510 12190 2530
rect 12210 2510 12220 2530
rect 12180 2495 12220 2510
rect 12240 2880 12280 2895
rect 12240 2860 12250 2880
rect 12270 2860 12280 2880
rect 12240 2830 12280 2860
rect 12240 2810 12250 2830
rect 12270 2810 12280 2830
rect 12240 2780 12280 2810
rect 12240 2760 12250 2780
rect 12270 2760 12280 2780
rect 12240 2730 12280 2760
rect 12240 2710 12250 2730
rect 12270 2710 12280 2730
rect 12240 2680 12280 2710
rect 12240 2660 12250 2680
rect 12270 2660 12280 2680
rect 12240 2630 12280 2660
rect 12240 2610 12250 2630
rect 12270 2610 12280 2630
rect 12240 2580 12280 2610
rect 12240 2560 12250 2580
rect 12270 2560 12280 2580
rect 12240 2530 12280 2560
rect 12240 2510 12250 2530
rect 12270 2510 12280 2530
rect 12240 2495 12280 2510
rect 12300 2880 12340 2895
rect 12300 2860 12310 2880
rect 12330 2860 12340 2880
rect 12300 2830 12340 2860
rect 12300 2810 12310 2830
rect 12330 2810 12340 2830
rect 12300 2780 12340 2810
rect 12300 2760 12310 2780
rect 12330 2760 12340 2780
rect 12300 2730 12340 2760
rect 12300 2710 12310 2730
rect 12330 2710 12340 2730
rect 12300 2680 12340 2710
rect 12300 2660 12310 2680
rect 12330 2660 12340 2680
rect 12300 2630 12340 2660
rect 12300 2610 12310 2630
rect 12330 2610 12340 2630
rect 12300 2580 12340 2610
rect 12300 2560 12310 2580
rect 12330 2560 12340 2580
rect 12300 2530 12340 2560
rect 12300 2510 12310 2530
rect 12330 2510 12340 2530
rect 12300 2495 12340 2510
rect 12360 2880 12400 2895
rect 12360 2860 12370 2880
rect 12390 2860 12400 2880
rect 12360 2830 12400 2860
rect 12360 2810 12370 2830
rect 12390 2810 12400 2830
rect 12360 2780 12400 2810
rect 12360 2760 12370 2780
rect 12390 2760 12400 2780
rect 12360 2730 12400 2760
rect 12360 2710 12370 2730
rect 12390 2710 12400 2730
rect 12360 2680 12400 2710
rect 12360 2660 12370 2680
rect 12390 2660 12400 2680
rect 12360 2630 12400 2660
rect 12360 2610 12370 2630
rect 12390 2610 12400 2630
rect 12360 2580 12400 2610
rect 12360 2560 12370 2580
rect 12390 2560 12400 2580
rect 12360 2530 12400 2560
rect 12360 2510 12370 2530
rect 12390 2510 12400 2530
rect 12360 2495 12400 2510
rect 12420 2880 12460 2895
rect 12420 2860 12430 2880
rect 12450 2860 12460 2880
rect 12420 2830 12460 2860
rect 12420 2810 12430 2830
rect 12450 2810 12460 2830
rect 12420 2780 12460 2810
rect 12420 2760 12430 2780
rect 12450 2760 12460 2780
rect 12420 2730 12460 2760
rect 12420 2710 12430 2730
rect 12450 2710 12460 2730
rect 12420 2680 12460 2710
rect 12420 2660 12430 2680
rect 12450 2660 12460 2680
rect 12420 2630 12460 2660
rect 12420 2610 12430 2630
rect 12450 2610 12460 2630
rect 12420 2580 12460 2610
rect 12420 2560 12430 2580
rect 12450 2560 12460 2580
rect 12420 2530 12460 2560
rect 12420 2510 12430 2530
rect 12450 2510 12460 2530
rect 12420 2495 12460 2510
rect 12480 2880 12520 2895
rect 12480 2860 12490 2880
rect 12510 2860 12520 2880
rect 12480 2830 12520 2860
rect 12480 2810 12490 2830
rect 12510 2810 12520 2830
rect 12480 2780 12520 2810
rect 12480 2760 12490 2780
rect 12510 2760 12520 2780
rect 12480 2730 12520 2760
rect 12480 2710 12490 2730
rect 12510 2710 12520 2730
rect 12480 2680 12520 2710
rect 12480 2660 12490 2680
rect 12510 2660 12520 2680
rect 12480 2630 12520 2660
rect 12480 2610 12490 2630
rect 12510 2610 12520 2630
rect 12480 2580 12520 2610
rect 12480 2560 12490 2580
rect 12510 2560 12520 2580
rect 12480 2530 12520 2560
rect 12480 2510 12490 2530
rect 12510 2510 12520 2530
rect 12480 2495 12520 2510
rect 12540 2880 12580 2895
rect 12540 2860 12550 2880
rect 12570 2860 12580 2880
rect 12540 2830 12580 2860
rect 12540 2810 12550 2830
rect 12570 2810 12580 2830
rect 12540 2780 12580 2810
rect 12540 2760 12550 2780
rect 12570 2760 12580 2780
rect 12540 2730 12580 2760
rect 12540 2710 12550 2730
rect 12570 2710 12580 2730
rect 12540 2680 12580 2710
rect 12540 2660 12550 2680
rect 12570 2660 12580 2680
rect 26220 2880 26260 2895
rect 26220 2860 26230 2880
rect 26250 2860 26260 2880
rect 26220 2830 26260 2860
rect 26220 2810 26230 2830
rect 26250 2810 26260 2830
rect 26220 2780 26260 2810
rect 26220 2760 26230 2780
rect 26250 2760 26260 2780
rect 26220 2730 26260 2760
rect 26220 2710 26230 2730
rect 26250 2710 26260 2730
rect 26220 2680 26260 2710
rect 12540 2630 12580 2660
rect 26220 2660 26230 2680
rect 26250 2660 26260 2680
rect 12540 2610 12550 2630
rect 12570 2610 12580 2630
rect 12540 2580 12580 2610
rect 12540 2560 12550 2580
rect 12570 2560 12580 2580
rect 12540 2530 12580 2560
rect 12540 2510 12550 2530
rect 12570 2510 12580 2530
rect 12540 2495 12580 2510
rect 12945 2640 12985 2655
rect 12945 2620 12955 2640
rect 12975 2620 12985 2640
rect 12945 2590 12985 2620
rect 12945 2570 12955 2590
rect 12975 2570 12985 2590
rect 12945 2540 12985 2570
rect 12945 2520 12955 2540
rect 12975 2520 12985 2540
rect 10815 2470 10825 2490
rect 10845 2470 10855 2490
rect 12945 2490 12985 2520
rect 12945 2470 12955 2490
rect 12975 2470 12985 2490
rect 10815 2455 10855 2470
rect 12945 2455 12985 2470
rect 13000 2640 13040 2655
rect 13000 2620 13010 2640
rect 13030 2620 13040 2640
rect 13000 2590 13040 2620
rect 13000 2570 13010 2590
rect 13030 2570 13040 2590
rect 13000 2540 13040 2570
rect 13000 2520 13010 2540
rect 13030 2520 13040 2540
rect 13000 2490 13040 2520
rect 13000 2470 13010 2490
rect 13030 2470 13040 2490
rect 13000 2455 13040 2470
rect 13055 2640 13095 2655
rect 13055 2620 13065 2640
rect 13085 2620 13095 2640
rect 13055 2590 13095 2620
rect 13055 2570 13065 2590
rect 13085 2570 13095 2590
rect 13055 2540 13095 2570
rect 13055 2520 13065 2540
rect 13085 2520 13095 2540
rect 13055 2490 13095 2520
rect 13055 2470 13065 2490
rect 13085 2470 13095 2490
rect 13055 2455 13095 2470
rect 13110 2640 13150 2655
rect 13110 2620 13120 2640
rect 13140 2620 13150 2640
rect 13110 2590 13150 2620
rect 13110 2570 13120 2590
rect 13140 2570 13150 2590
rect 13110 2540 13150 2570
rect 13110 2520 13120 2540
rect 13140 2520 13150 2540
rect 13110 2490 13150 2520
rect 13110 2470 13120 2490
rect 13140 2470 13150 2490
rect 13110 2455 13150 2470
rect 13165 2640 13205 2655
rect 13165 2620 13175 2640
rect 13195 2620 13205 2640
rect 13165 2590 13205 2620
rect 13165 2570 13175 2590
rect 13195 2570 13205 2590
rect 13165 2540 13205 2570
rect 13165 2520 13175 2540
rect 13195 2520 13205 2540
rect 13165 2490 13205 2520
rect 13165 2470 13175 2490
rect 13195 2470 13205 2490
rect 13165 2455 13205 2470
rect 13220 2640 13260 2655
rect 13220 2620 13230 2640
rect 13250 2620 13260 2640
rect 13220 2590 13260 2620
rect 13220 2570 13230 2590
rect 13250 2570 13260 2590
rect 13220 2540 13260 2570
rect 13220 2520 13230 2540
rect 13250 2520 13260 2540
rect 13220 2490 13260 2520
rect 13220 2470 13230 2490
rect 13250 2470 13260 2490
rect 13220 2455 13260 2470
rect 13275 2640 13315 2655
rect 13275 2620 13285 2640
rect 13305 2620 13315 2640
rect 13275 2590 13315 2620
rect 13275 2570 13285 2590
rect 13305 2570 13315 2590
rect 13275 2540 13315 2570
rect 13275 2520 13285 2540
rect 13305 2520 13315 2540
rect 13275 2490 13315 2520
rect 13275 2470 13285 2490
rect 13305 2470 13315 2490
rect 13275 2455 13315 2470
rect 13330 2640 13370 2655
rect 13330 2620 13340 2640
rect 13360 2620 13370 2640
rect 13330 2590 13370 2620
rect 13330 2570 13340 2590
rect 13360 2570 13370 2590
rect 13330 2540 13370 2570
rect 13330 2520 13340 2540
rect 13360 2520 13370 2540
rect 13330 2490 13370 2520
rect 13330 2470 13340 2490
rect 13360 2470 13370 2490
rect 13330 2455 13370 2470
rect 13385 2640 13425 2655
rect 13385 2620 13395 2640
rect 13415 2620 13425 2640
rect 13385 2590 13425 2620
rect 13385 2570 13395 2590
rect 13415 2570 13425 2590
rect 13385 2540 13425 2570
rect 13385 2520 13395 2540
rect 13415 2520 13425 2540
rect 13385 2490 13425 2520
rect 13385 2470 13395 2490
rect 13415 2470 13425 2490
rect 13385 2455 13425 2470
rect 13440 2640 13480 2655
rect 13440 2620 13450 2640
rect 13470 2620 13480 2640
rect 13440 2590 13480 2620
rect 13440 2570 13450 2590
rect 13470 2570 13480 2590
rect 13440 2540 13480 2570
rect 13440 2520 13450 2540
rect 13470 2520 13480 2540
rect 13440 2490 13480 2520
rect 13440 2470 13450 2490
rect 13470 2470 13480 2490
rect 13440 2455 13480 2470
rect 13495 2640 13535 2655
rect 13495 2620 13505 2640
rect 13525 2620 13535 2640
rect 13495 2590 13535 2620
rect 13495 2570 13505 2590
rect 13525 2570 13535 2590
rect 13495 2540 13535 2570
rect 13495 2520 13505 2540
rect 13525 2520 13535 2540
rect 13495 2490 13535 2520
rect 13495 2470 13505 2490
rect 13525 2470 13535 2490
rect 13495 2455 13535 2470
rect 13550 2640 13590 2655
rect 13550 2620 13560 2640
rect 13580 2620 13590 2640
rect 13550 2590 13590 2620
rect 13550 2570 13560 2590
rect 13580 2570 13590 2590
rect 13550 2540 13590 2570
rect 13550 2520 13560 2540
rect 13580 2520 13590 2540
rect 13550 2490 13590 2520
rect 13550 2470 13560 2490
rect 13580 2470 13590 2490
rect 13550 2455 13590 2470
rect 13605 2640 13645 2655
rect 13605 2620 13615 2640
rect 13635 2620 13645 2640
rect 13605 2590 13645 2620
rect 13605 2570 13615 2590
rect 13635 2570 13645 2590
rect 13605 2540 13645 2570
rect 13605 2520 13615 2540
rect 13635 2520 13645 2540
rect 13605 2490 13645 2520
rect 13605 2470 13615 2490
rect 13635 2470 13645 2490
rect 13605 2455 13645 2470
rect 10155 2250 10195 2265
rect 10155 2230 10165 2250
rect 10185 2230 10195 2250
rect 10155 2200 10195 2230
rect 10155 2180 10165 2200
rect 10185 2180 10195 2200
rect 10155 2150 10195 2180
rect 10155 2130 10165 2150
rect 10185 2130 10195 2150
rect 10155 2100 10195 2130
rect 10155 2080 10165 2100
rect 10185 2080 10195 2100
rect 10155 2050 10195 2080
rect 10155 2030 10165 2050
rect 10185 2030 10195 2050
rect 10155 2000 10195 2030
rect 10155 1980 10165 2000
rect 10185 1980 10195 2000
rect 10155 1965 10195 1980
rect 10210 2250 10250 2265
rect 10210 2230 10220 2250
rect 10240 2230 10250 2250
rect 10210 2200 10250 2230
rect 10210 2180 10220 2200
rect 10240 2180 10250 2200
rect 10210 2150 10250 2180
rect 10210 2130 10220 2150
rect 10240 2130 10250 2150
rect 10210 2100 10250 2130
rect 10210 2080 10220 2100
rect 10240 2080 10250 2100
rect 10210 2050 10250 2080
rect 10210 2030 10220 2050
rect 10240 2030 10250 2050
rect 10210 2000 10250 2030
rect 10210 1980 10220 2000
rect 10240 1980 10250 2000
rect 10210 1965 10250 1980
rect 10265 2250 10305 2265
rect 10265 2230 10275 2250
rect 10295 2230 10305 2250
rect 10265 2200 10305 2230
rect 10265 2180 10275 2200
rect 10295 2180 10305 2200
rect 10265 2150 10305 2180
rect 10265 2130 10275 2150
rect 10295 2130 10305 2150
rect 10265 2100 10305 2130
rect 10265 2080 10275 2100
rect 10295 2080 10305 2100
rect 10265 2050 10305 2080
rect 10265 2030 10275 2050
rect 10295 2030 10305 2050
rect 10265 2000 10305 2030
rect 10265 1980 10275 2000
rect 10295 1980 10305 2000
rect 10265 1965 10305 1980
rect 10320 2250 10360 2265
rect 10320 2230 10330 2250
rect 10350 2230 10360 2250
rect 10320 2200 10360 2230
rect 10320 2180 10330 2200
rect 10350 2180 10360 2200
rect 10320 2150 10360 2180
rect 10320 2130 10330 2150
rect 10350 2130 10360 2150
rect 10320 2100 10360 2130
rect 10320 2080 10330 2100
rect 10350 2080 10360 2100
rect 10320 2050 10360 2080
rect 10320 2030 10330 2050
rect 10350 2030 10360 2050
rect 10320 2000 10360 2030
rect 10320 1980 10330 2000
rect 10350 1980 10360 2000
rect 10320 1965 10360 1980
rect 10375 2250 10415 2265
rect 10375 2230 10385 2250
rect 10405 2230 10415 2250
rect 10375 2200 10415 2230
rect 10375 2180 10385 2200
rect 10405 2180 10415 2200
rect 10375 2150 10415 2180
rect 10375 2130 10385 2150
rect 10405 2130 10415 2150
rect 10375 2100 10415 2130
rect 10375 2080 10385 2100
rect 10405 2080 10415 2100
rect 10375 2050 10415 2080
rect 10375 2030 10385 2050
rect 10405 2030 10415 2050
rect 10375 2000 10415 2030
rect 10375 1980 10385 2000
rect 10405 1980 10415 2000
rect 10375 1965 10415 1980
rect 10430 2250 10470 2265
rect 10430 2230 10440 2250
rect 10460 2230 10470 2250
rect 10430 2200 10470 2230
rect 10430 2180 10440 2200
rect 10460 2180 10470 2200
rect 10430 2150 10470 2180
rect 10430 2130 10440 2150
rect 10460 2130 10470 2150
rect 10430 2100 10470 2130
rect 10430 2080 10440 2100
rect 10460 2080 10470 2100
rect 10430 2050 10470 2080
rect 10430 2030 10440 2050
rect 10460 2030 10470 2050
rect 10430 2000 10470 2030
rect 10430 1980 10440 2000
rect 10460 1980 10470 2000
rect 10430 1965 10470 1980
rect 10485 2250 10525 2265
rect 10485 2230 10495 2250
rect 10515 2230 10525 2250
rect 10485 2200 10525 2230
rect 10485 2180 10495 2200
rect 10515 2180 10525 2200
rect 10485 2150 10525 2180
rect 10485 2130 10495 2150
rect 10515 2130 10525 2150
rect 10485 2100 10525 2130
rect 10485 2080 10495 2100
rect 10515 2080 10525 2100
rect 10485 2050 10525 2080
rect 10485 2030 10495 2050
rect 10515 2030 10525 2050
rect 10485 2000 10525 2030
rect 10485 1980 10495 2000
rect 10515 1980 10525 2000
rect 10485 1965 10525 1980
rect 10540 2250 10580 2265
rect 10540 2230 10550 2250
rect 10570 2230 10580 2250
rect 10540 2200 10580 2230
rect 10540 2180 10550 2200
rect 10570 2180 10580 2200
rect 10540 2150 10580 2180
rect 10540 2130 10550 2150
rect 10570 2130 10580 2150
rect 10540 2100 10580 2130
rect 10540 2080 10550 2100
rect 10570 2080 10580 2100
rect 10540 2050 10580 2080
rect 10540 2030 10550 2050
rect 10570 2030 10580 2050
rect 10540 2000 10580 2030
rect 10540 1980 10550 2000
rect 10570 1980 10580 2000
rect 10540 1965 10580 1980
rect 10595 2250 10635 2265
rect 10595 2230 10605 2250
rect 10625 2230 10635 2250
rect 10595 2200 10635 2230
rect 10595 2180 10605 2200
rect 10625 2180 10635 2200
rect 10595 2150 10635 2180
rect 10595 2130 10605 2150
rect 10625 2130 10635 2150
rect 10595 2100 10635 2130
rect 10595 2080 10605 2100
rect 10625 2080 10635 2100
rect 10595 2050 10635 2080
rect 10595 2030 10605 2050
rect 10625 2030 10635 2050
rect 10595 2000 10635 2030
rect 10595 1980 10605 2000
rect 10625 1980 10635 2000
rect 10595 1965 10635 1980
rect 10650 2250 10690 2265
rect 10650 2230 10660 2250
rect 10680 2230 10690 2250
rect 10650 2200 10690 2230
rect 10650 2180 10660 2200
rect 10680 2180 10690 2200
rect 10650 2150 10690 2180
rect 10650 2130 10660 2150
rect 10680 2130 10690 2150
rect 10650 2100 10690 2130
rect 10650 2080 10660 2100
rect 10680 2080 10690 2100
rect 10650 2050 10690 2080
rect 10650 2030 10660 2050
rect 10680 2030 10690 2050
rect 10650 2000 10690 2030
rect 10650 1980 10660 2000
rect 10680 1980 10690 2000
rect 10650 1965 10690 1980
rect 10705 2250 10745 2265
rect 10705 2230 10715 2250
rect 10735 2230 10745 2250
rect 10705 2200 10745 2230
rect 10705 2180 10715 2200
rect 10735 2180 10745 2200
rect 10705 2150 10745 2180
rect 10705 2130 10715 2150
rect 10735 2130 10745 2150
rect 10705 2100 10745 2130
rect 10705 2080 10715 2100
rect 10735 2080 10745 2100
rect 10705 2050 10745 2080
rect 10705 2030 10715 2050
rect 10735 2030 10745 2050
rect 10705 2000 10745 2030
rect 10705 1980 10715 2000
rect 10735 1980 10745 2000
rect 10705 1965 10745 1980
rect 10760 2250 10800 2265
rect 10760 2230 10770 2250
rect 10790 2230 10800 2250
rect 10760 2200 10800 2230
rect 10760 2180 10770 2200
rect 10790 2180 10800 2200
rect 10760 2150 10800 2180
rect 10760 2130 10770 2150
rect 10790 2130 10800 2150
rect 10760 2100 10800 2130
rect 10760 2080 10770 2100
rect 10790 2080 10800 2100
rect 10760 2050 10800 2080
rect 10760 2030 10770 2050
rect 10790 2030 10800 2050
rect 10760 2000 10800 2030
rect 10760 1980 10770 2000
rect 10790 1980 10800 2000
rect 10760 1965 10800 1980
rect 10815 2250 10855 2265
rect 10815 2230 10825 2250
rect 10845 2230 10855 2250
rect 10815 2200 10855 2230
rect 10815 2180 10825 2200
rect 10845 2180 10855 2200
rect 12945 2250 12985 2265
rect 12945 2230 12955 2250
rect 12975 2230 12985 2250
rect 12945 2200 12985 2230
rect 10815 2150 10855 2180
rect 12945 2180 12955 2200
rect 12975 2180 12985 2200
rect 10815 2130 10825 2150
rect 10845 2130 10855 2150
rect 12945 2150 12985 2180
rect 12945 2130 12955 2150
rect 12975 2130 12985 2150
rect 10815 2100 10855 2130
rect 10815 2080 10825 2100
rect 10845 2080 10855 2100
rect 10815 2050 10855 2080
rect 10815 2030 10825 2050
rect 10845 2030 10855 2050
rect 10815 2000 10855 2030
rect 10815 1980 10825 2000
rect 10845 1980 10855 2000
rect 11275 2115 11315 2130
rect 11275 2095 11285 2115
rect 11305 2095 11315 2115
rect 11275 2065 11315 2095
rect 11275 2045 11285 2065
rect 11305 2045 11315 2065
rect 11275 2015 11315 2045
rect 11275 1995 11285 2015
rect 11305 1995 11315 2015
rect 11275 1980 11315 1995
rect 11330 2115 11370 2130
rect 11330 2095 11340 2115
rect 11360 2095 11370 2115
rect 11330 2065 11370 2095
rect 11330 2045 11340 2065
rect 11360 2045 11370 2065
rect 11330 2015 11370 2045
rect 11330 1995 11340 2015
rect 11360 1995 11370 2015
rect 11330 1980 11370 1995
rect 11385 2115 11425 2130
rect 11385 2095 11395 2115
rect 11415 2095 11425 2115
rect 11385 2065 11425 2095
rect 11385 2045 11395 2065
rect 11415 2045 11425 2065
rect 11385 2015 11425 2045
rect 11385 1995 11395 2015
rect 11415 1995 11425 2015
rect 11385 1980 11425 1995
rect 11440 2115 11480 2130
rect 11440 2095 11450 2115
rect 11470 2095 11480 2115
rect 11440 2065 11480 2095
rect 11440 2045 11450 2065
rect 11470 2045 11480 2065
rect 11440 2015 11480 2045
rect 11440 1995 11450 2015
rect 11470 1995 11480 2015
rect 11440 1980 11480 1995
rect 11495 2115 11535 2130
rect 11495 2095 11505 2115
rect 11525 2095 11535 2115
rect 11495 2065 11535 2095
rect 11495 2045 11505 2065
rect 11525 2045 11535 2065
rect 11495 2015 11535 2045
rect 11495 1995 11505 2015
rect 11525 1995 11535 2015
rect 11495 1980 11535 1995
rect 11550 2115 11590 2130
rect 11550 2095 11560 2115
rect 11580 2095 11590 2115
rect 11550 2065 11590 2095
rect 11550 2045 11560 2065
rect 11580 2045 11590 2065
rect 11550 2015 11590 2045
rect 11550 1995 11560 2015
rect 11580 1995 11590 2015
rect 11550 1980 11590 1995
rect 11605 2115 11645 2130
rect 11605 2095 11615 2115
rect 11635 2095 11645 2115
rect 11605 2065 11645 2095
rect 11605 2045 11615 2065
rect 11635 2045 11645 2065
rect 11605 2015 11645 2045
rect 11605 1995 11615 2015
rect 11635 1995 11645 2015
rect 11605 1980 11645 1995
rect 11660 2115 11700 2130
rect 11660 2095 11670 2115
rect 11690 2095 11700 2115
rect 11660 2065 11700 2095
rect 11660 2045 11670 2065
rect 11690 2045 11700 2065
rect 11660 2015 11700 2045
rect 11660 1995 11670 2015
rect 11690 1995 11700 2015
rect 11660 1980 11700 1995
rect 11715 2115 11755 2130
rect 11715 2095 11725 2115
rect 11745 2095 11755 2115
rect 11715 2065 11755 2095
rect 11715 2045 11725 2065
rect 11745 2045 11755 2065
rect 11715 2015 11755 2045
rect 11715 1995 11725 2015
rect 11745 1995 11755 2015
rect 11715 1980 11755 1995
rect 11770 2115 11810 2130
rect 11770 2095 11780 2115
rect 11800 2095 11810 2115
rect 11770 2065 11810 2095
rect 11770 2045 11780 2065
rect 11800 2045 11810 2065
rect 11770 2015 11810 2045
rect 11770 1995 11780 2015
rect 11800 1995 11810 2015
rect 11770 1980 11810 1995
rect 11825 2115 11865 2130
rect 11825 2095 11835 2115
rect 11855 2095 11865 2115
rect 11825 2065 11865 2095
rect 11825 2045 11835 2065
rect 11855 2045 11865 2065
rect 11825 2015 11865 2045
rect 11825 1995 11835 2015
rect 11855 1995 11865 2015
rect 11825 1980 11865 1995
rect 11880 2115 11920 2130
rect 11880 2095 11890 2115
rect 11910 2095 11920 2115
rect 11880 2065 11920 2095
rect 11880 2045 11890 2065
rect 11910 2045 11920 2065
rect 11880 2015 11920 2045
rect 11880 1995 11890 2015
rect 11910 1995 11920 2015
rect 11880 1980 11920 1995
rect 11935 2115 11975 2130
rect 11935 2095 11945 2115
rect 11965 2095 11975 2115
rect 11935 2065 11975 2095
rect 11935 2045 11945 2065
rect 11965 2045 11975 2065
rect 11935 2015 11975 2045
rect 11935 1995 11945 2015
rect 11965 1995 11975 2015
rect 11935 1980 11975 1995
rect 11990 2115 12030 2130
rect 11990 2095 12000 2115
rect 12020 2095 12030 2115
rect 11990 2065 12030 2095
rect 11990 2045 12000 2065
rect 12020 2045 12030 2065
rect 11990 2015 12030 2045
rect 11990 1995 12000 2015
rect 12020 1995 12030 2015
rect 11990 1980 12030 1995
rect 12045 2115 12085 2130
rect 12045 2095 12055 2115
rect 12075 2095 12085 2115
rect 12045 2065 12085 2095
rect 12045 2045 12055 2065
rect 12075 2045 12085 2065
rect 12045 2015 12085 2045
rect 12045 1995 12055 2015
rect 12075 1995 12085 2015
rect 12045 1980 12085 1995
rect 12100 2115 12140 2130
rect 12100 2095 12110 2115
rect 12130 2095 12140 2115
rect 12100 2065 12140 2095
rect 12100 2045 12110 2065
rect 12130 2045 12140 2065
rect 12100 2015 12140 2045
rect 12100 1995 12110 2015
rect 12130 1995 12140 2015
rect 12100 1980 12140 1995
rect 12155 2115 12195 2130
rect 12155 2095 12165 2115
rect 12185 2095 12195 2115
rect 12155 2065 12195 2095
rect 12155 2045 12165 2065
rect 12185 2045 12195 2065
rect 12155 2015 12195 2045
rect 12155 1995 12165 2015
rect 12185 1995 12195 2015
rect 12155 1980 12195 1995
rect 12210 2115 12250 2130
rect 12210 2095 12220 2115
rect 12240 2095 12250 2115
rect 12210 2065 12250 2095
rect 12210 2045 12220 2065
rect 12240 2045 12250 2065
rect 12210 2015 12250 2045
rect 12210 1995 12220 2015
rect 12240 1995 12250 2015
rect 12210 1980 12250 1995
rect 12265 2115 12305 2130
rect 12265 2095 12275 2115
rect 12295 2095 12305 2115
rect 12265 2065 12305 2095
rect 12265 2045 12275 2065
rect 12295 2045 12305 2065
rect 12265 2015 12305 2045
rect 12265 1995 12275 2015
rect 12295 1995 12305 2015
rect 12265 1980 12305 1995
rect 12320 2115 12360 2130
rect 12320 2095 12330 2115
rect 12350 2095 12360 2115
rect 12320 2065 12360 2095
rect 12320 2045 12330 2065
rect 12350 2045 12360 2065
rect 12320 2015 12360 2045
rect 12320 1995 12330 2015
rect 12350 1995 12360 2015
rect 12320 1980 12360 1995
rect 12375 2115 12415 2130
rect 12375 2095 12385 2115
rect 12405 2095 12415 2115
rect 12375 2065 12415 2095
rect 12375 2045 12385 2065
rect 12405 2045 12415 2065
rect 12375 2015 12415 2045
rect 12375 1995 12385 2015
rect 12405 1995 12415 2015
rect 12375 1980 12415 1995
rect 12430 2115 12470 2130
rect 12430 2095 12440 2115
rect 12460 2095 12470 2115
rect 12430 2065 12470 2095
rect 12430 2045 12440 2065
rect 12460 2045 12470 2065
rect 12430 2015 12470 2045
rect 12430 1995 12440 2015
rect 12460 1995 12470 2015
rect 12430 1980 12470 1995
rect 12485 2115 12525 2130
rect 12485 2095 12495 2115
rect 12515 2095 12525 2115
rect 12485 2065 12525 2095
rect 12485 2045 12495 2065
rect 12515 2045 12525 2065
rect 12485 2015 12525 2045
rect 12485 1995 12495 2015
rect 12515 1995 12525 2015
rect 12485 1980 12525 1995
rect 12945 2100 12985 2130
rect 12945 2080 12955 2100
rect 12975 2080 12985 2100
rect 12945 2050 12985 2080
rect 12945 2030 12955 2050
rect 12975 2030 12985 2050
rect 12945 2000 12985 2030
rect 12945 1980 12955 2000
rect 12975 1980 12985 2000
rect 10815 1965 10855 1980
rect 12945 1965 12985 1980
rect 13000 2250 13040 2265
rect 13000 2230 13010 2250
rect 13030 2230 13040 2250
rect 13000 2200 13040 2230
rect 13000 2180 13010 2200
rect 13030 2180 13040 2200
rect 13000 2150 13040 2180
rect 13000 2130 13010 2150
rect 13030 2130 13040 2150
rect 13000 2100 13040 2130
rect 13000 2080 13010 2100
rect 13030 2080 13040 2100
rect 13000 2050 13040 2080
rect 13000 2030 13010 2050
rect 13030 2030 13040 2050
rect 13000 2000 13040 2030
rect 13000 1980 13010 2000
rect 13030 1980 13040 2000
rect 13000 1965 13040 1980
rect 13055 2250 13095 2265
rect 13055 2230 13065 2250
rect 13085 2230 13095 2250
rect 13055 2200 13095 2230
rect 13055 2180 13065 2200
rect 13085 2180 13095 2200
rect 13055 2150 13095 2180
rect 13055 2130 13065 2150
rect 13085 2130 13095 2150
rect 13055 2100 13095 2130
rect 13055 2080 13065 2100
rect 13085 2080 13095 2100
rect 13055 2050 13095 2080
rect 13055 2030 13065 2050
rect 13085 2030 13095 2050
rect 13055 2000 13095 2030
rect 13055 1980 13065 2000
rect 13085 1980 13095 2000
rect 13055 1965 13095 1980
rect 13110 2250 13150 2265
rect 13110 2230 13120 2250
rect 13140 2230 13150 2250
rect 13110 2200 13150 2230
rect 13110 2180 13120 2200
rect 13140 2180 13150 2200
rect 13110 2150 13150 2180
rect 13110 2130 13120 2150
rect 13140 2130 13150 2150
rect 13110 2100 13150 2130
rect 13110 2080 13120 2100
rect 13140 2080 13150 2100
rect 13110 2050 13150 2080
rect 13110 2030 13120 2050
rect 13140 2030 13150 2050
rect 13110 2000 13150 2030
rect 13110 1980 13120 2000
rect 13140 1980 13150 2000
rect 13110 1965 13150 1980
rect 13165 2250 13205 2265
rect 13165 2230 13175 2250
rect 13195 2230 13205 2250
rect 13165 2200 13205 2230
rect 13165 2180 13175 2200
rect 13195 2180 13205 2200
rect 13165 2150 13205 2180
rect 13165 2130 13175 2150
rect 13195 2130 13205 2150
rect 13165 2100 13205 2130
rect 13165 2080 13175 2100
rect 13195 2080 13205 2100
rect 13165 2050 13205 2080
rect 13165 2030 13175 2050
rect 13195 2030 13205 2050
rect 13165 2000 13205 2030
rect 13165 1980 13175 2000
rect 13195 1980 13205 2000
rect 13165 1965 13205 1980
rect 13220 2250 13260 2265
rect 13220 2230 13230 2250
rect 13250 2230 13260 2250
rect 13220 2200 13260 2230
rect 13220 2180 13230 2200
rect 13250 2180 13260 2200
rect 13220 2150 13260 2180
rect 13220 2130 13230 2150
rect 13250 2130 13260 2150
rect 13220 2100 13260 2130
rect 13220 2080 13230 2100
rect 13250 2080 13260 2100
rect 13220 2050 13260 2080
rect 13220 2030 13230 2050
rect 13250 2030 13260 2050
rect 13220 2000 13260 2030
rect 13220 1980 13230 2000
rect 13250 1980 13260 2000
rect 13220 1965 13260 1980
rect 13275 2250 13315 2265
rect 13275 2230 13285 2250
rect 13305 2230 13315 2250
rect 13275 2200 13315 2230
rect 13275 2180 13285 2200
rect 13305 2180 13315 2200
rect 13275 2150 13315 2180
rect 13275 2130 13285 2150
rect 13305 2130 13315 2150
rect 13275 2100 13315 2130
rect 13275 2080 13285 2100
rect 13305 2080 13315 2100
rect 13275 2050 13315 2080
rect 13275 2030 13285 2050
rect 13305 2030 13315 2050
rect 13275 2000 13315 2030
rect 13275 1980 13285 2000
rect 13305 1980 13315 2000
rect 13275 1965 13315 1980
rect 13330 2250 13370 2265
rect 13330 2230 13340 2250
rect 13360 2230 13370 2250
rect 13330 2200 13370 2230
rect 13330 2180 13340 2200
rect 13360 2180 13370 2200
rect 13330 2150 13370 2180
rect 13330 2130 13340 2150
rect 13360 2130 13370 2150
rect 13330 2100 13370 2130
rect 13330 2080 13340 2100
rect 13360 2080 13370 2100
rect 13330 2050 13370 2080
rect 13330 2030 13340 2050
rect 13360 2030 13370 2050
rect 13330 2000 13370 2030
rect 13330 1980 13340 2000
rect 13360 1980 13370 2000
rect 13330 1965 13370 1980
rect 13385 2250 13425 2265
rect 13385 2230 13395 2250
rect 13415 2230 13425 2250
rect 13385 2200 13425 2230
rect 13385 2180 13395 2200
rect 13415 2180 13425 2200
rect 13385 2150 13425 2180
rect 13385 2130 13395 2150
rect 13415 2130 13425 2150
rect 13385 2100 13425 2130
rect 13385 2080 13395 2100
rect 13415 2080 13425 2100
rect 13385 2050 13425 2080
rect 13385 2030 13395 2050
rect 13415 2030 13425 2050
rect 13385 2000 13425 2030
rect 13385 1980 13395 2000
rect 13415 1980 13425 2000
rect 13385 1965 13425 1980
rect 13440 2250 13480 2265
rect 13440 2230 13450 2250
rect 13470 2230 13480 2250
rect 13440 2200 13480 2230
rect 13440 2180 13450 2200
rect 13470 2180 13480 2200
rect 13440 2150 13480 2180
rect 13440 2130 13450 2150
rect 13470 2130 13480 2150
rect 13440 2100 13480 2130
rect 13440 2080 13450 2100
rect 13470 2080 13480 2100
rect 13440 2050 13480 2080
rect 13440 2030 13450 2050
rect 13470 2030 13480 2050
rect 13440 2000 13480 2030
rect 13440 1980 13450 2000
rect 13470 1980 13480 2000
rect 13440 1965 13480 1980
rect 13495 2250 13535 2265
rect 13495 2230 13505 2250
rect 13525 2230 13535 2250
rect 13495 2200 13535 2230
rect 13495 2180 13505 2200
rect 13525 2180 13535 2200
rect 13495 2150 13535 2180
rect 13495 2130 13505 2150
rect 13525 2130 13535 2150
rect 13495 2100 13535 2130
rect 13495 2080 13505 2100
rect 13525 2080 13535 2100
rect 13495 2050 13535 2080
rect 13495 2030 13505 2050
rect 13525 2030 13535 2050
rect 13495 2000 13535 2030
rect 13495 1980 13505 2000
rect 13525 1980 13535 2000
rect 13495 1965 13535 1980
rect 13550 2250 13590 2265
rect 13550 2230 13560 2250
rect 13580 2230 13590 2250
rect 13550 2200 13590 2230
rect 13550 2180 13560 2200
rect 13580 2180 13590 2200
rect 13550 2150 13590 2180
rect 13550 2130 13560 2150
rect 13580 2130 13590 2150
rect 13550 2100 13590 2130
rect 13550 2080 13560 2100
rect 13580 2080 13590 2100
rect 13550 2050 13590 2080
rect 13550 2030 13560 2050
rect 13580 2030 13590 2050
rect 13550 2000 13590 2030
rect 13550 1980 13560 2000
rect 13580 1980 13590 2000
rect 13550 1965 13590 1980
rect 13605 2250 13645 2265
rect 13605 2230 13615 2250
rect 13635 2230 13645 2250
rect 13605 2200 13645 2230
rect 13605 2180 13615 2200
rect 13635 2180 13645 2200
rect 13605 2150 13645 2180
rect 13605 2130 13615 2150
rect 13635 2130 13645 2150
rect 13605 2100 13645 2130
rect 13605 2080 13615 2100
rect 13635 2080 13645 2100
rect 13605 2050 13645 2080
rect 13605 2030 13615 2050
rect 13635 2030 13645 2050
rect 13605 2000 13645 2030
rect 26220 2630 26260 2660
rect 24680 2605 24720 2620
rect 24680 2585 24690 2605
rect 24710 2585 24720 2605
rect 24680 2555 24720 2585
rect 24680 2535 24690 2555
rect 24710 2535 24720 2555
rect 24680 2520 24720 2535
rect 24735 2605 24775 2620
rect 24735 2585 24745 2605
rect 24765 2585 24775 2605
rect 24735 2555 24775 2585
rect 24735 2535 24745 2555
rect 24765 2535 24775 2555
rect 24735 2520 24775 2535
rect 24790 2605 24830 2620
rect 24790 2585 24800 2605
rect 24820 2585 24830 2605
rect 24790 2555 24830 2585
rect 24790 2535 24800 2555
rect 24820 2535 24830 2555
rect 24790 2520 24830 2535
rect 24845 2605 24885 2620
rect 24845 2585 24855 2605
rect 24875 2585 24885 2605
rect 24845 2555 24885 2585
rect 24845 2535 24855 2555
rect 24875 2535 24885 2555
rect 24845 2520 24885 2535
rect 24900 2605 24940 2620
rect 24900 2585 24910 2605
rect 24930 2585 24940 2605
rect 24900 2555 24940 2585
rect 24900 2535 24910 2555
rect 24930 2535 24940 2555
rect 24900 2520 24940 2535
rect 24955 2605 24995 2620
rect 24955 2585 24965 2605
rect 24985 2585 24995 2605
rect 24955 2555 24995 2585
rect 24955 2535 24965 2555
rect 24985 2535 24995 2555
rect 24955 2520 24995 2535
rect 25010 2605 25050 2620
rect 25010 2585 25020 2605
rect 25040 2585 25050 2605
rect 25010 2555 25050 2585
rect 25010 2535 25020 2555
rect 25040 2535 25050 2555
rect 25010 2520 25050 2535
rect 25065 2605 25105 2620
rect 25065 2585 25075 2605
rect 25095 2585 25105 2605
rect 25065 2555 25105 2585
rect 25065 2535 25075 2555
rect 25095 2535 25105 2555
rect 25065 2520 25105 2535
rect 25120 2605 25160 2620
rect 25120 2585 25130 2605
rect 25150 2585 25160 2605
rect 25120 2555 25160 2585
rect 25120 2535 25130 2555
rect 25150 2535 25160 2555
rect 25120 2520 25160 2535
rect 25175 2605 25215 2620
rect 25175 2585 25185 2605
rect 25205 2585 25215 2605
rect 25175 2555 25215 2585
rect 25175 2535 25185 2555
rect 25205 2535 25215 2555
rect 25175 2520 25215 2535
rect 25230 2605 25270 2620
rect 25230 2585 25240 2605
rect 25260 2585 25270 2605
rect 25230 2555 25270 2585
rect 25230 2535 25240 2555
rect 25260 2535 25270 2555
rect 25230 2520 25270 2535
rect 25285 2605 25325 2620
rect 25285 2585 25295 2605
rect 25315 2585 25325 2605
rect 25285 2555 25325 2585
rect 25285 2535 25295 2555
rect 25315 2535 25325 2555
rect 25285 2520 25325 2535
rect 25340 2605 25380 2620
rect 25340 2585 25350 2605
rect 25370 2585 25380 2605
rect 25340 2555 25380 2585
rect 25340 2535 25350 2555
rect 25370 2535 25380 2555
rect 25340 2520 25380 2535
rect 25395 2605 25435 2620
rect 25395 2585 25405 2605
rect 25425 2585 25435 2605
rect 25395 2555 25435 2585
rect 25395 2535 25405 2555
rect 25425 2535 25435 2555
rect 25395 2520 25435 2535
rect 25450 2605 25490 2620
rect 25450 2585 25460 2605
rect 25480 2585 25490 2605
rect 25450 2555 25490 2585
rect 25450 2535 25460 2555
rect 25480 2535 25490 2555
rect 25450 2520 25490 2535
rect 25505 2605 25545 2620
rect 25505 2585 25515 2605
rect 25535 2585 25545 2605
rect 25505 2555 25545 2585
rect 25505 2535 25515 2555
rect 25535 2535 25545 2555
rect 25505 2520 25545 2535
rect 25560 2605 25600 2620
rect 25560 2585 25570 2605
rect 25590 2585 25600 2605
rect 25560 2555 25600 2585
rect 25560 2535 25570 2555
rect 25590 2535 25600 2555
rect 25560 2520 25600 2535
rect 25615 2605 25655 2620
rect 25615 2585 25625 2605
rect 25645 2585 25655 2605
rect 25615 2555 25655 2585
rect 25615 2535 25625 2555
rect 25645 2535 25655 2555
rect 25615 2520 25655 2535
rect 25670 2605 25710 2620
rect 25670 2585 25680 2605
rect 25700 2585 25710 2605
rect 25670 2555 25710 2585
rect 25670 2535 25680 2555
rect 25700 2535 25710 2555
rect 25670 2520 25710 2535
rect 25725 2605 25765 2620
rect 25725 2585 25735 2605
rect 25755 2585 25765 2605
rect 25725 2555 25765 2585
rect 25725 2535 25735 2555
rect 25755 2535 25765 2555
rect 25725 2520 25765 2535
rect 25780 2605 25820 2620
rect 25780 2585 25790 2605
rect 25810 2585 25820 2605
rect 25780 2555 25820 2585
rect 25780 2535 25790 2555
rect 25810 2535 25820 2555
rect 25780 2520 25820 2535
rect 25835 2605 25875 2620
rect 25835 2585 25845 2605
rect 25865 2585 25875 2605
rect 25835 2555 25875 2585
rect 25835 2535 25845 2555
rect 25865 2535 25875 2555
rect 25835 2520 25875 2535
rect 25890 2605 25930 2620
rect 25890 2585 25900 2605
rect 25920 2585 25930 2605
rect 25890 2555 25930 2585
rect 25890 2535 25900 2555
rect 25920 2535 25930 2555
rect 25890 2520 25930 2535
rect 26220 2610 26230 2630
rect 26250 2610 26260 2630
rect 26220 2580 26260 2610
rect 26220 2560 26230 2580
rect 26250 2560 26260 2580
rect 26220 2530 26260 2560
rect 26220 2510 26230 2530
rect 26250 2510 26260 2530
rect 26220 2495 26260 2510
rect 26280 2880 26320 2895
rect 26280 2860 26290 2880
rect 26310 2860 26320 2880
rect 26280 2830 26320 2860
rect 26280 2810 26290 2830
rect 26310 2810 26320 2830
rect 26280 2780 26320 2810
rect 26280 2760 26290 2780
rect 26310 2760 26320 2780
rect 26280 2730 26320 2760
rect 26280 2710 26290 2730
rect 26310 2710 26320 2730
rect 26280 2680 26320 2710
rect 26280 2660 26290 2680
rect 26310 2660 26320 2680
rect 26280 2630 26320 2660
rect 26280 2610 26290 2630
rect 26310 2610 26320 2630
rect 26280 2580 26320 2610
rect 26280 2560 26290 2580
rect 26310 2560 26320 2580
rect 26280 2530 26320 2560
rect 26280 2510 26290 2530
rect 26310 2510 26320 2530
rect 26280 2495 26320 2510
rect 26340 2880 26380 2895
rect 26340 2860 26350 2880
rect 26370 2860 26380 2880
rect 26340 2830 26380 2860
rect 26340 2810 26350 2830
rect 26370 2810 26380 2830
rect 26340 2780 26380 2810
rect 26340 2760 26350 2780
rect 26370 2760 26380 2780
rect 26340 2730 26380 2760
rect 26340 2710 26350 2730
rect 26370 2710 26380 2730
rect 26340 2680 26380 2710
rect 26340 2660 26350 2680
rect 26370 2660 26380 2680
rect 26340 2630 26380 2660
rect 26340 2610 26350 2630
rect 26370 2610 26380 2630
rect 26340 2580 26380 2610
rect 26340 2560 26350 2580
rect 26370 2560 26380 2580
rect 26340 2530 26380 2560
rect 26340 2510 26350 2530
rect 26370 2510 26380 2530
rect 26340 2495 26380 2510
rect 26400 2880 26440 2895
rect 26400 2860 26410 2880
rect 26430 2860 26440 2880
rect 26400 2830 26440 2860
rect 26400 2810 26410 2830
rect 26430 2810 26440 2830
rect 26400 2780 26440 2810
rect 26400 2760 26410 2780
rect 26430 2760 26440 2780
rect 26400 2730 26440 2760
rect 26400 2710 26410 2730
rect 26430 2710 26440 2730
rect 26400 2680 26440 2710
rect 26400 2660 26410 2680
rect 26430 2660 26440 2680
rect 26400 2630 26440 2660
rect 26400 2610 26410 2630
rect 26430 2610 26440 2630
rect 26400 2580 26440 2610
rect 26400 2560 26410 2580
rect 26430 2560 26440 2580
rect 26400 2530 26440 2560
rect 26400 2510 26410 2530
rect 26430 2510 26440 2530
rect 26400 2495 26440 2510
rect 26460 2880 26500 2895
rect 26460 2860 26470 2880
rect 26490 2860 26500 2880
rect 26460 2830 26500 2860
rect 26460 2810 26470 2830
rect 26490 2810 26500 2830
rect 26460 2780 26500 2810
rect 26460 2760 26470 2780
rect 26490 2760 26500 2780
rect 26460 2730 26500 2760
rect 26460 2710 26470 2730
rect 26490 2710 26500 2730
rect 26460 2680 26500 2710
rect 26460 2660 26470 2680
rect 26490 2660 26500 2680
rect 26460 2630 26500 2660
rect 26460 2610 26470 2630
rect 26490 2610 26500 2630
rect 26460 2580 26500 2610
rect 26460 2560 26470 2580
rect 26490 2560 26500 2580
rect 26460 2530 26500 2560
rect 26460 2510 26470 2530
rect 26490 2510 26500 2530
rect 26460 2495 26500 2510
rect 26520 2880 26560 2895
rect 26520 2860 26530 2880
rect 26550 2860 26560 2880
rect 26520 2830 26560 2860
rect 26520 2810 26530 2830
rect 26550 2810 26560 2830
rect 26520 2780 26560 2810
rect 26520 2760 26530 2780
rect 26550 2760 26560 2780
rect 26520 2730 26560 2760
rect 26520 2710 26530 2730
rect 26550 2710 26560 2730
rect 26520 2680 26560 2710
rect 26520 2660 26530 2680
rect 26550 2660 26560 2680
rect 26520 2630 26560 2660
rect 26520 2610 26530 2630
rect 26550 2610 26560 2630
rect 26520 2580 26560 2610
rect 26520 2560 26530 2580
rect 26550 2560 26560 2580
rect 26520 2530 26560 2560
rect 26520 2510 26530 2530
rect 26550 2510 26560 2530
rect 26520 2495 26560 2510
rect 26580 2880 26620 2895
rect 26580 2860 26590 2880
rect 26610 2860 26620 2880
rect 26580 2830 26620 2860
rect 26580 2810 26590 2830
rect 26610 2810 26620 2830
rect 26580 2780 26620 2810
rect 26580 2760 26590 2780
rect 26610 2760 26620 2780
rect 26580 2730 26620 2760
rect 26580 2710 26590 2730
rect 26610 2710 26620 2730
rect 26580 2680 26620 2710
rect 26580 2660 26590 2680
rect 26610 2660 26620 2680
rect 26580 2630 26620 2660
rect 26580 2610 26590 2630
rect 26610 2610 26620 2630
rect 26580 2580 26620 2610
rect 26580 2560 26590 2580
rect 26610 2560 26620 2580
rect 26580 2530 26620 2560
rect 26580 2510 26590 2530
rect 26610 2510 26620 2530
rect 26580 2495 26620 2510
rect 26640 2880 26680 2895
rect 26640 2860 26650 2880
rect 26670 2860 26680 2880
rect 26640 2830 26680 2860
rect 26640 2810 26650 2830
rect 26670 2810 26680 2830
rect 26640 2780 26680 2810
rect 26640 2760 26650 2780
rect 26670 2760 26680 2780
rect 26640 2730 26680 2760
rect 26640 2710 26650 2730
rect 26670 2710 26680 2730
rect 26640 2680 26680 2710
rect 26640 2660 26650 2680
rect 26670 2660 26680 2680
rect 26640 2630 26680 2660
rect 26640 2610 26650 2630
rect 26670 2610 26680 2630
rect 26640 2580 26680 2610
rect 26640 2560 26650 2580
rect 26670 2560 26680 2580
rect 26640 2530 26680 2560
rect 26640 2510 26650 2530
rect 26670 2510 26680 2530
rect 26640 2495 26680 2510
rect 26700 2880 26740 2895
rect 26700 2860 26710 2880
rect 26730 2860 26740 2880
rect 26700 2830 26740 2860
rect 26700 2810 26710 2830
rect 26730 2810 26740 2830
rect 26700 2780 26740 2810
rect 26700 2760 26710 2780
rect 26730 2760 26740 2780
rect 26700 2730 26740 2760
rect 26700 2710 26710 2730
rect 26730 2710 26740 2730
rect 26700 2680 26740 2710
rect 26700 2660 26710 2680
rect 26730 2660 26740 2680
rect 26700 2630 26740 2660
rect 26700 2610 26710 2630
rect 26730 2610 26740 2630
rect 26700 2580 26740 2610
rect 26700 2560 26710 2580
rect 26730 2560 26740 2580
rect 26700 2530 26740 2560
rect 26700 2510 26710 2530
rect 26730 2510 26740 2530
rect 26700 2495 26740 2510
rect 26760 2880 26800 2895
rect 26760 2860 26770 2880
rect 26790 2860 26800 2880
rect 26760 2830 26800 2860
rect 26760 2810 26770 2830
rect 26790 2810 26800 2830
rect 26760 2780 26800 2810
rect 26760 2760 26770 2780
rect 26790 2760 26800 2780
rect 26760 2730 26800 2760
rect 26760 2710 26770 2730
rect 26790 2710 26800 2730
rect 26760 2680 26800 2710
rect 26760 2660 26770 2680
rect 26790 2660 26800 2680
rect 26760 2630 26800 2660
rect 26760 2610 26770 2630
rect 26790 2610 26800 2630
rect 26760 2580 26800 2610
rect 26760 2560 26770 2580
rect 26790 2560 26800 2580
rect 26760 2530 26800 2560
rect 26760 2510 26770 2530
rect 26790 2510 26800 2530
rect 26760 2495 26800 2510
rect 26820 2880 26860 2895
rect 26820 2860 26830 2880
rect 26850 2860 26860 2880
rect 26820 2830 26860 2860
rect 26820 2810 26830 2830
rect 26850 2810 26860 2830
rect 26820 2780 26860 2810
rect 26820 2760 26830 2780
rect 26850 2760 26860 2780
rect 26820 2730 26860 2760
rect 26820 2710 26830 2730
rect 26850 2710 26860 2730
rect 26820 2680 26860 2710
rect 26820 2660 26830 2680
rect 26850 2660 26860 2680
rect 26820 2630 26860 2660
rect 26820 2610 26830 2630
rect 26850 2610 26860 2630
rect 26820 2580 26860 2610
rect 26820 2560 26830 2580
rect 26850 2560 26860 2580
rect 26820 2530 26860 2560
rect 26820 2510 26830 2530
rect 26850 2510 26860 2530
rect 26820 2495 26860 2510
rect 26880 2880 26920 2895
rect 26880 2860 26890 2880
rect 26910 2860 26920 2880
rect 26880 2830 26920 2860
rect 26880 2810 26890 2830
rect 26910 2810 26920 2830
rect 26880 2780 26920 2810
rect 26880 2760 26890 2780
rect 26910 2760 26920 2780
rect 26880 2730 26920 2760
rect 26880 2710 26890 2730
rect 26910 2710 26920 2730
rect 26880 2680 26920 2710
rect 26880 2660 26890 2680
rect 26910 2660 26920 2680
rect 26880 2630 26920 2660
rect 26880 2610 26890 2630
rect 26910 2610 26920 2630
rect 26880 2580 26920 2610
rect 26880 2560 26890 2580
rect 26910 2560 26920 2580
rect 26880 2530 26920 2560
rect 26880 2510 26890 2530
rect 26910 2510 26920 2530
rect 26880 2495 26920 2510
rect 26940 2880 26980 2895
rect 26940 2860 26950 2880
rect 26970 2860 26980 2880
rect 26940 2830 26980 2860
rect 26940 2810 26950 2830
rect 26970 2810 26980 2830
rect 26940 2780 26980 2810
rect 26940 2760 26950 2780
rect 26970 2760 26980 2780
rect 26940 2730 26980 2760
rect 26940 2710 26950 2730
rect 26970 2710 26980 2730
rect 26940 2680 26980 2710
rect 26940 2660 26950 2680
rect 26970 2660 26980 2680
rect 26940 2630 26980 2660
rect 26940 2610 26950 2630
rect 26970 2610 26980 2630
rect 26940 2580 26980 2610
rect 26940 2560 26950 2580
rect 26970 2560 26980 2580
rect 26940 2530 26980 2560
rect 26940 2510 26950 2530
rect 26970 2510 26980 2530
rect 26940 2495 26980 2510
rect 27000 2880 27040 2895
rect 27000 2860 27010 2880
rect 27030 2860 27040 2880
rect 27000 2830 27040 2860
rect 27000 2810 27010 2830
rect 27030 2810 27040 2830
rect 27000 2780 27040 2810
rect 27000 2760 27010 2780
rect 27030 2760 27040 2780
rect 27000 2730 27040 2760
rect 27000 2710 27010 2730
rect 27030 2710 27040 2730
rect 27000 2680 27040 2710
rect 27000 2660 27010 2680
rect 27030 2660 27040 2680
rect 27000 2630 27040 2660
rect 27000 2610 27010 2630
rect 27030 2610 27040 2630
rect 27000 2580 27040 2610
rect 27000 2560 27010 2580
rect 27030 2560 27040 2580
rect 27000 2530 27040 2560
rect 27000 2510 27010 2530
rect 27030 2510 27040 2530
rect 27000 2495 27040 2510
rect 27060 2880 27100 2895
rect 27060 2860 27070 2880
rect 27090 2860 27100 2880
rect 27060 2830 27100 2860
rect 27060 2810 27070 2830
rect 27090 2810 27100 2830
rect 27060 2780 27100 2810
rect 27060 2760 27070 2780
rect 27090 2760 27100 2780
rect 27060 2730 27100 2760
rect 27060 2710 27070 2730
rect 27090 2710 27100 2730
rect 27060 2680 27100 2710
rect 27060 2660 27070 2680
rect 27090 2660 27100 2680
rect 27060 2630 27100 2660
rect 27060 2610 27070 2630
rect 27090 2610 27100 2630
rect 27060 2580 27100 2610
rect 27060 2560 27070 2580
rect 27090 2560 27100 2580
rect 27060 2530 27100 2560
rect 27060 2510 27070 2530
rect 27090 2510 27100 2530
rect 27060 2495 27100 2510
rect 27120 2880 27160 2895
rect 27120 2860 27130 2880
rect 27150 2860 27160 2880
rect 27120 2830 27160 2860
rect 27120 2810 27130 2830
rect 27150 2810 27160 2830
rect 27120 2780 27160 2810
rect 27120 2760 27130 2780
rect 27150 2760 27160 2780
rect 27120 2730 27160 2760
rect 27120 2710 27130 2730
rect 27150 2710 27160 2730
rect 27120 2680 27160 2710
rect 27120 2660 27130 2680
rect 27150 2660 27160 2680
rect 27120 2630 27160 2660
rect 27120 2610 27130 2630
rect 27150 2610 27160 2630
rect 27120 2580 27160 2610
rect 27120 2560 27130 2580
rect 27150 2560 27160 2580
rect 27120 2530 27160 2560
rect 27120 2510 27130 2530
rect 27150 2510 27160 2530
rect 27120 2495 27160 2510
rect 27180 2880 27220 2895
rect 27180 2860 27190 2880
rect 27210 2860 27220 2880
rect 27180 2830 27220 2860
rect 27180 2810 27190 2830
rect 27210 2810 27220 2830
rect 27180 2780 27220 2810
rect 27180 2760 27190 2780
rect 27210 2760 27220 2780
rect 27180 2730 27220 2760
rect 27180 2710 27190 2730
rect 27210 2710 27220 2730
rect 27180 2680 27220 2710
rect 27180 2660 27190 2680
rect 27210 2660 27220 2680
rect 27180 2630 27220 2660
rect 27180 2610 27190 2630
rect 27210 2610 27220 2630
rect 27180 2580 27220 2610
rect 27180 2560 27190 2580
rect 27210 2560 27220 2580
rect 27180 2530 27220 2560
rect 27180 2510 27190 2530
rect 27210 2510 27220 2530
rect 27180 2495 27220 2510
rect 27240 2880 27280 2895
rect 27240 2860 27250 2880
rect 27270 2860 27280 2880
rect 27240 2830 27280 2860
rect 27240 2810 27250 2830
rect 27270 2810 27280 2830
rect 27240 2780 27280 2810
rect 27240 2760 27250 2780
rect 27270 2760 27280 2780
rect 27240 2730 27280 2760
rect 27240 2710 27250 2730
rect 27270 2710 27280 2730
rect 27240 2680 27280 2710
rect 27240 2660 27250 2680
rect 27270 2660 27280 2680
rect 27240 2630 27280 2660
rect 27240 2610 27250 2630
rect 27270 2610 27280 2630
rect 27240 2580 27280 2610
rect 27240 2560 27250 2580
rect 27270 2560 27280 2580
rect 27240 2530 27280 2560
rect 27240 2510 27250 2530
rect 27270 2510 27280 2530
rect 27240 2495 27280 2510
rect 27300 2880 27340 2895
rect 27300 2860 27310 2880
rect 27330 2860 27340 2880
rect 27300 2830 27340 2860
rect 27300 2810 27310 2830
rect 27330 2810 27340 2830
rect 27300 2780 27340 2810
rect 27300 2760 27310 2780
rect 27330 2760 27340 2780
rect 27300 2730 27340 2760
rect 27300 2710 27310 2730
rect 27330 2710 27340 2730
rect 27300 2680 27340 2710
rect 27300 2660 27310 2680
rect 27330 2660 27340 2680
rect 27300 2630 27340 2660
rect 27300 2610 27310 2630
rect 27330 2610 27340 2630
rect 27300 2580 27340 2610
rect 27300 2560 27310 2580
rect 27330 2560 27340 2580
rect 27300 2530 27340 2560
rect 27300 2510 27310 2530
rect 27330 2510 27340 2530
rect 27300 2495 27340 2510
rect 27360 2880 27400 2895
rect 27360 2860 27370 2880
rect 27390 2860 27400 2880
rect 27360 2830 27400 2860
rect 27360 2810 27370 2830
rect 27390 2810 27400 2830
rect 27360 2780 27400 2810
rect 27360 2760 27370 2780
rect 27390 2760 27400 2780
rect 27360 2730 27400 2760
rect 27360 2710 27370 2730
rect 27390 2710 27400 2730
rect 27360 2680 27400 2710
rect 27360 2660 27370 2680
rect 27390 2660 27400 2680
rect 27360 2630 27400 2660
rect 27360 2610 27370 2630
rect 27390 2610 27400 2630
rect 27360 2580 27400 2610
rect 27360 2560 27370 2580
rect 27390 2560 27400 2580
rect 27360 2530 27400 2560
rect 27360 2510 27370 2530
rect 27390 2510 27400 2530
rect 27360 2495 27400 2510
rect 27420 2880 27460 2895
rect 27420 2860 27430 2880
rect 27450 2860 27460 2880
rect 27420 2830 27460 2860
rect 27420 2810 27430 2830
rect 27450 2810 27460 2830
rect 27420 2780 27460 2810
rect 27420 2760 27430 2780
rect 27450 2760 27460 2780
rect 27420 2730 27460 2760
rect 27420 2710 27430 2730
rect 27450 2710 27460 2730
rect 27420 2680 27460 2710
rect 27420 2660 27430 2680
rect 27450 2660 27460 2680
rect 27420 2630 27460 2660
rect 27420 2610 27430 2630
rect 27450 2610 27460 2630
rect 27420 2580 27460 2610
rect 27420 2560 27430 2580
rect 27450 2560 27460 2580
rect 27420 2530 27460 2560
rect 27420 2510 27430 2530
rect 27450 2510 27460 2530
rect 27420 2495 27460 2510
rect 27480 2880 27520 2895
rect 27480 2860 27490 2880
rect 27510 2860 27520 2880
rect 27480 2830 27520 2860
rect 27480 2810 27490 2830
rect 27510 2810 27520 2830
rect 27480 2780 27520 2810
rect 27480 2760 27490 2780
rect 27510 2760 27520 2780
rect 27480 2730 27520 2760
rect 27480 2710 27490 2730
rect 27510 2710 27520 2730
rect 27480 2680 27520 2710
rect 27480 2660 27490 2680
rect 27510 2660 27520 2680
rect 27480 2630 27520 2660
rect 27480 2610 27490 2630
rect 27510 2610 27520 2630
rect 27480 2580 27520 2610
rect 27480 2560 27490 2580
rect 27510 2560 27520 2580
rect 27480 2530 27520 2560
rect 27480 2510 27490 2530
rect 27510 2510 27520 2530
rect 27480 2495 27520 2510
rect 27540 2880 27580 2895
rect 27540 2860 27550 2880
rect 27570 2860 27580 2880
rect 27540 2830 27580 2860
rect 27540 2810 27550 2830
rect 27570 2810 27580 2830
rect 27540 2780 27580 2810
rect 27540 2760 27550 2780
rect 27570 2760 27580 2780
rect 27540 2730 27580 2760
rect 27540 2710 27550 2730
rect 27570 2710 27580 2730
rect 27540 2680 27580 2710
rect 27540 2660 27550 2680
rect 27570 2660 27580 2680
rect 27540 2630 27580 2660
rect 27540 2610 27550 2630
rect 27570 2610 27580 2630
rect 27540 2580 27580 2610
rect 27540 2560 27550 2580
rect 27570 2560 27580 2580
rect 27540 2530 27580 2560
rect 27540 2510 27550 2530
rect 27570 2510 27580 2530
rect 27890 2605 27930 2620
rect 27890 2585 27900 2605
rect 27920 2585 27930 2605
rect 27890 2555 27930 2585
rect 27890 2535 27900 2555
rect 27920 2535 27930 2555
rect 27890 2520 27930 2535
rect 27945 2605 27985 2620
rect 27945 2585 27955 2605
rect 27975 2585 27985 2605
rect 27945 2555 27985 2585
rect 27945 2535 27955 2555
rect 27975 2535 27985 2555
rect 27945 2520 27985 2535
rect 28000 2605 28040 2620
rect 28000 2585 28010 2605
rect 28030 2585 28040 2605
rect 28000 2555 28040 2585
rect 28000 2535 28010 2555
rect 28030 2535 28040 2555
rect 28000 2520 28040 2535
rect 28055 2605 28095 2620
rect 28055 2585 28065 2605
rect 28085 2585 28095 2605
rect 28055 2555 28095 2585
rect 28055 2535 28065 2555
rect 28085 2535 28095 2555
rect 28055 2520 28095 2535
rect 28110 2605 28150 2620
rect 28110 2585 28120 2605
rect 28140 2585 28150 2605
rect 28110 2555 28150 2585
rect 28110 2535 28120 2555
rect 28140 2535 28150 2555
rect 28110 2520 28150 2535
rect 28165 2605 28205 2620
rect 28165 2585 28175 2605
rect 28195 2585 28205 2605
rect 28165 2555 28205 2585
rect 28165 2535 28175 2555
rect 28195 2535 28205 2555
rect 28165 2520 28205 2535
rect 28220 2605 28260 2620
rect 28220 2585 28230 2605
rect 28250 2585 28260 2605
rect 28220 2555 28260 2585
rect 28220 2535 28230 2555
rect 28250 2535 28260 2555
rect 28220 2520 28260 2535
rect 28275 2605 28315 2620
rect 28275 2585 28285 2605
rect 28305 2585 28315 2605
rect 28275 2555 28315 2585
rect 28275 2535 28285 2555
rect 28305 2535 28315 2555
rect 28275 2520 28315 2535
rect 28330 2605 28370 2620
rect 28330 2585 28340 2605
rect 28360 2585 28370 2605
rect 28330 2555 28370 2585
rect 28330 2535 28340 2555
rect 28360 2535 28370 2555
rect 28330 2520 28370 2535
rect 28385 2605 28425 2620
rect 28385 2585 28395 2605
rect 28415 2585 28425 2605
rect 28385 2555 28425 2585
rect 28385 2535 28395 2555
rect 28415 2535 28425 2555
rect 28385 2520 28425 2535
rect 28440 2605 28480 2620
rect 28440 2585 28450 2605
rect 28470 2585 28480 2605
rect 28440 2555 28480 2585
rect 28440 2535 28450 2555
rect 28470 2535 28480 2555
rect 28440 2520 28480 2535
rect 28495 2605 28535 2620
rect 28495 2585 28505 2605
rect 28525 2585 28535 2605
rect 28495 2555 28535 2585
rect 28495 2535 28505 2555
rect 28525 2535 28535 2555
rect 28495 2520 28535 2535
rect 28550 2605 28590 2620
rect 28550 2585 28560 2605
rect 28580 2585 28590 2605
rect 28550 2555 28590 2585
rect 28550 2535 28560 2555
rect 28580 2535 28590 2555
rect 28550 2520 28590 2535
rect 28605 2605 28645 2620
rect 28605 2585 28615 2605
rect 28635 2585 28645 2605
rect 28605 2555 28645 2585
rect 28605 2535 28615 2555
rect 28635 2535 28645 2555
rect 28605 2520 28645 2535
rect 28660 2605 28700 2620
rect 28660 2585 28670 2605
rect 28690 2585 28700 2605
rect 28660 2555 28700 2585
rect 28660 2535 28670 2555
rect 28690 2535 28700 2555
rect 28660 2520 28700 2535
rect 28715 2605 28755 2620
rect 28715 2585 28725 2605
rect 28745 2585 28755 2605
rect 28715 2555 28755 2585
rect 28715 2535 28725 2555
rect 28745 2535 28755 2555
rect 28715 2520 28755 2535
rect 28770 2605 28810 2620
rect 28770 2585 28780 2605
rect 28800 2585 28810 2605
rect 28770 2555 28810 2585
rect 28770 2535 28780 2555
rect 28800 2535 28810 2555
rect 28770 2520 28810 2535
rect 28825 2605 28865 2620
rect 28825 2585 28835 2605
rect 28855 2585 28865 2605
rect 28825 2555 28865 2585
rect 28825 2535 28835 2555
rect 28855 2535 28865 2555
rect 28825 2520 28865 2535
rect 28880 2605 28920 2620
rect 28880 2585 28890 2605
rect 28910 2585 28920 2605
rect 28880 2555 28920 2585
rect 28880 2535 28890 2555
rect 28910 2535 28920 2555
rect 28880 2520 28920 2535
rect 28935 2605 28975 2620
rect 28935 2585 28945 2605
rect 28965 2585 28975 2605
rect 28935 2555 28975 2585
rect 28935 2535 28945 2555
rect 28965 2535 28975 2555
rect 28935 2520 28975 2535
rect 28990 2605 29030 2620
rect 28990 2585 29000 2605
rect 29020 2585 29030 2605
rect 28990 2555 29030 2585
rect 28990 2535 29000 2555
rect 29020 2535 29030 2555
rect 28990 2520 29030 2535
rect 29045 2605 29085 2620
rect 29045 2585 29055 2605
rect 29075 2585 29085 2605
rect 29045 2555 29085 2585
rect 29045 2535 29055 2555
rect 29075 2535 29085 2555
rect 29045 2520 29085 2535
rect 29100 2605 29140 2620
rect 29100 2585 29110 2605
rect 29130 2585 29140 2605
rect 29100 2555 29140 2585
rect 29100 2535 29110 2555
rect 29130 2535 29140 2555
rect 29100 2520 29140 2535
rect 27540 2495 27580 2510
rect 24680 2155 24720 2170
rect 24680 2135 24690 2155
rect 24710 2135 24720 2155
rect 24680 2105 24720 2135
rect 24680 2085 24690 2105
rect 24710 2085 24720 2105
rect 24680 2055 24720 2085
rect 24680 2035 24690 2055
rect 24710 2035 24720 2055
rect 24680 2020 24720 2035
rect 24735 2155 24775 2170
rect 24735 2135 24745 2155
rect 24765 2135 24775 2155
rect 24735 2105 24775 2135
rect 24735 2085 24745 2105
rect 24765 2085 24775 2105
rect 24735 2055 24775 2085
rect 24735 2035 24745 2055
rect 24765 2035 24775 2055
rect 24735 2020 24775 2035
rect 24790 2155 24830 2170
rect 24790 2135 24800 2155
rect 24820 2135 24830 2155
rect 24790 2105 24830 2135
rect 24790 2085 24800 2105
rect 24820 2085 24830 2105
rect 24790 2055 24830 2085
rect 24790 2035 24800 2055
rect 24820 2035 24830 2055
rect 24790 2020 24830 2035
rect 24845 2155 24885 2170
rect 24845 2135 24855 2155
rect 24875 2135 24885 2155
rect 24845 2105 24885 2135
rect 24845 2085 24855 2105
rect 24875 2085 24885 2105
rect 24845 2055 24885 2085
rect 24845 2035 24855 2055
rect 24875 2035 24885 2055
rect 24845 2020 24885 2035
rect 24900 2155 24940 2170
rect 24900 2135 24910 2155
rect 24930 2135 24940 2155
rect 24900 2105 24940 2135
rect 24900 2085 24910 2105
rect 24930 2085 24940 2105
rect 24900 2055 24940 2085
rect 24900 2035 24910 2055
rect 24930 2035 24940 2055
rect 24900 2020 24940 2035
rect 24955 2155 24995 2170
rect 24955 2135 24965 2155
rect 24985 2135 24995 2155
rect 24955 2105 24995 2135
rect 24955 2085 24965 2105
rect 24985 2085 24995 2105
rect 24955 2055 24995 2085
rect 24955 2035 24965 2055
rect 24985 2035 24995 2055
rect 24955 2020 24995 2035
rect 25010 2155 25050 2170
rect 25010 2135 25020 2155
rect 25040 2135 25050 2155
rect 25010 2105 25050 2135
rect 25010 2085 25020 2105
rect 25040 2085 25050 2105
rect 25010 2055 25050 2085
rect 25010 2035 25020 2055
rect 25040 2035 25050 2055
rect 25010 2020 25050 2035
rect 25065 2155 25105 2170
rect 25065 2135 25075 2155
rect 25095 2135 25105 2155
rect 25065 2105 25105 2135
rect 25065 2085 25075 2105
rect 25095 2085 25105 2105
rect 25065 2055 25105 2085
rect 25065 2035 25075 2055
rect 25095 2035 25105 2055
rect 25065 2020 25105 2035
rect 25120 2155 25160 2170
rect 25120 2135 25130 2155
rect 25150 2135 25160 2155
rect 25120 2105 25160 2135
rect 25120 2085 25130 2105
rect 25150 2085 25160 2105
rect 25120 2055 25160 2085
rect 25120 2035 25130 2055
rect 25150 2035 25160 2055
rect 25120 2020 25160 2035
rect 25175 2155 25215 2170
rect 25175 2135 25185 2155
rect 25205 2135 25215 2155
rect 25175 2105 25215 2135
rect 25175 2085 25185 2105
rect 25205 2085 25215 2105
rect 25175 2055 25215 2085
rect 25175 2035 25185 2055
rect 25205 2035 25215 2055
rect 25175 2020 25215 2035
rect 25230 2155 25270 2170
rect 25230 2135 25240 2155
rect 25260 2135 25270 2155
rect 25230 2105 25270 2135
rect 25230 2085 25240 2105
rect 25260 2085 25270 2105
rect 25230 2055 25270 2085
rect 25230 2035 25240 2055
rect 25260 2035 25270 2055
rect 25230 2020 25270 2035
rect 25285 2155 25325 2170
rect 25285 2135 25295 2155
rect 25315 2135 25325 2155
rect 25285 2105 25325 2135
rect 25285 2085 25295 2105
rect 25315 2085 25325 2105
rect 25285 2055 25325 2085
rect 25285 2035 25295 2055
rect 25315 2035 25325 2055
rect 25285 2020 25325 2035
rect 25340 2155 25380 2170
rect 25340 2135 25350 2155
rect 25370 2135 25380 2155
rect 25340 2105 25380 2135
rect 25340 2085 25350 2105
rect 25370 2085 25380 2105
rect 25340 2055 25380 2085
rect 25340 2035 25350 2055
rect 25370 2035 25380 2055
rect 25340 2020 25380 2035
rect 25395 2155 25435 2170
rect 25395 2135 25405 2155
rect 25425 2135 25435 2155
rect 25395 2105 25435 2135
rect 25395 2085 25405 2105
rect 25425 2085 25435 2105
rect 25395 2055 25435 2085
rect 25395 2035 25405 2055
rect 25425 2035 25435 2055
rect 25395 2020 25435 2035
rect 25450 2155 25490 2170
rect 25450 2135 25460 2155
rect 25480 2135 25490 2155
rect 25450 2105 25490 2135
rect 25450 2085 25460 2105
rect 25480 2085 25490 2105
rect 25450 2055 25490 2085
rect 25450 2035 25460 2055
rect 25480 2035 25490 2055
rect 25450 2020 25490 2035
rect 25505 2155 25545 2170
rect 25505 2135 25515 2155
rect 25535 2135 25545 2155
rect 25505 2105 25545 2135
rect 25505 2085 25515 2105
rect 25535 2085 25545 2105
rect 25505 2055 25545 2085
rect 25505 2035 25515 2055
rect 25535 2035 25545 2055
rect 25505 2020 25545 2035
rect 25560 2155 25600 2170
rect 25560 2135 25570 2155
rect 25590 2135 25600 2155
rect 25560 2105 25600 2135
rect 25560 2085 25570 2105
rect 25590 2085 25600 2105
rect 25560 2055 25600 2085
rect 25560 2035 25570 2055
rect 25590 2035 25600 2055
rect 25560 2020 25600 2035
rect 25615 2155 25655 2170
rect 25615 2135 25625 2155
rect 25645 2135 25655 2155
rect 25615 2105 25655 2135
rect 25615 2085 25625 2105
rect 25645 2085 25655 2105
rect 25615 2055 25655 2085
rect 25615 2035 25625 2055
rect 25645 2035 25655 2055
rect 25615 2020 25655 2035
rect 25670 2155 25710 2170
rect 25670 2135 25680 2155
rect 25700 2135 25710 2155
rect 25670 2105 25710 2135
rect 25670 2085 25680 2105
rect 25700 2085 25710 2105
rect 25670 2055 25710 2085
rect 25670 2035 25680 2055
rect 25700 2035 25710 2055
rect 25670 2020 25710 2035
rect 25725 2155 25765 2170
rect 25725 2135 25735 2155
rect 25755 2135 25765 2155
rect 25725 2105 25765 2135
rect 25725 2085 25735 2105
rect 25755 2085 25765 2105
rect 25725 2055 25765 2085
rect 25725 2035 25735 2055
rect 25755 2035 25765 2055
rect 25725 2020 25765 2035
rect 25780 2155 25820 2170
rect 25780 2135 25790 2155
rect 25810 2135 25820 2155
rect 25780 2105 25820 2135
rect 25780 2085 25790 2105
rect 25810 2085 25820 2105
rect 25780 2055 25820 2085
rect 25780 2035 25790 2055
rect 25810 2035 25820 2055
rect 25780 2020 25820 2035
rect 25835 2155 25875 2170
rect 25835 2135 25845 2155
rect 25865 2135 25875 2155
rect 25835 2105 25875 2135
rect 25835 2085 25845 2105
rect 25865 2085 25875 2105
rect 25835 2055 25875 2085
rect 25835 2035 25845 2055
rect 25865 2035 25875 2055
rect 25835 2020 25875 2035
rect 25890 2155 25930 2170
rect 27890 2155 27930 2170
rect 25890 2135 25900 2155
rect 25920 2135 25930 2155
rect 25890 2105 25930 2135
rect 27890 2135 27900 2155
rect 27920 2135 27930 2155
rect 25890 2085 25900 2105
rect 25920 2085 25930 2105
rect 25890 2055 25930 2085
rect 25890 2035 25900 2055
rect 25920 2035 25930 2055
rect 25890 2020 25930 2035
rect 26275 2115 26315 2130
rect 26275 2095 26285 2115
rect 26305 2095 26315 2115
rect 26275 2065 26315 2095
rect 26275 2045 26285 2065
rect 26305 2045 26315 2065
rect 26275 2015 26315 2045
rect 13605 1980 13615 2000
rect 13635 1980 13645 2000
rect 26275 1995 26285 2015
rect 26305 1995 26315 2015
rect 26275 1980 26315 1995
rect 26330 2115 26370 2130
rect 26330 2095 26340 2115
rect 26360 2095 26370 2115
rect 26330 2065 26370 2095
rect 26330 2045 26340 2065
rect 26360 2045 26370 2065
rect 26330 2015 26370 2045
rect 26330 1995 26340 2015
rect 26360 1995 26370 2015
rect 26330 1980 26370 1995
rect 26385 2115 26425 2130
rect 26385 2095 26395 2115
rect 26415 2095 26425 2115
rect 26385 2065 26425 2095
rect 26385 2045 26395 2065
rect 26415 2045 26425 2065
rect 26385 2015 26425 2045
rect 26385 1995 26395 2015
rect 26415 1995 26425 2015
rect 26385 1980 26425 1995
rect 26440 2115 26480 2130
rect 26440 2095 26450 2115
rect 26470 2095 26480 2115
rect 26440 2065 26480 2095
rect 26440 2045 26450 2065
rect 26470 2045 26480 2065
rect 26440 2015 26480 2045
rect 26440 1995 26450 2015
rect 26470 1995 26480 2015
rect 26440 1980 26480 1995
rect 26495 2115 26535 2130
rect 26495 2095 26505 2115
rect 26525 2095 26535 2115
rect 26495 2065 26535 2095
rect 26495 2045 26505 2065
rect 26525 2045 26535 2065
rect 26495 2015 26535 2045
rect 26495 1995 26505 2015
rect 26525 1995 26535 2015
rect 26495 1980 26535 1995
rect 26550 2115 26590 2130
rect 26550 2095 26560 2115
rect 26580 2095 26590 2115
rect 26550 2065 26590 2095
rect 26550 2045 26560 2065
rect 26580 2045 26590 2065
rect 26550 2015 26590 2045
rect 26550 1995 26560 2015
rect 26580 1995 26590 2015
rect 26550 1980 26590 1995
rect 26605 2115 26645 2130
rect 26605 2095 26615 2115
rect 26635 2095 26645 2115
rect 26605 2065 26645 2095
rect 26605 2045 26615 2065
rect 26635 2045 26645 2065
rect 26605 2015 26645 2045
rect 26605 1995 26615 2015
rect 26635 1995 26645 2015
rect 26605 1980 26645 1995
rect 26660 2115 26700 2130
rect 26660 2095 26670 2115
rect 26690 2095 26700 2115
rect 26660 2065 26700 2095
rect 26660 2045 26670 2065
rect 26690 2045 26700 2065
rect 26660 2015 26700 2045
rect 26660 1995 26670 2015
rect 26690 1995 26700 2015
rect 26660 1980 26700 1995
rect 26715 2115 26755 2130
rect 26715 2095 26725 2115
rect 26745 2095 26755 2115
rect 26715 2065 26755 2095
rect 26715 2045 26725 2065
rect 26745 2045 26755 2065
rect 26715 2015 26755 2045
rect 26715 1995 26725 2015
rect 26745 1995 26755 2015
rect 26715 1980 26755 1995
rect 26770 2115 26810 2130
rect 26770 2095 26780 2115
rect 26800 2095 26810 2115
rect 26770 2065 26810 2095
rect 26770 2045 26780 2065
rect 26800 2045 26810 2065
rect 26770 2015 26810 2045
rect 26770 1995 26780 2015
rect 26800 1995 26810 2015
rect 26770 1980 26810 1995
rect 26825 2115 26865 2130
rect 26825 2095 26835 2115
rect 26855 2095 26865 2115
rect 26825 2065 26865 2095
rect 26825 2045 26835 2065
rect 26855 2045 26865 2065
rect 26825 2015 26865 2045
rect 26825 1995 26835 2015
rect 26855 1995 26865 2015
rect 26825 1980 26865 1995
rect 26880 2115 26920 2130
rect 26880 2095 26890 2115
rect 26910 2095 26920 2115
rect 26880 2065 26920 2095
rect 26880 2045 26890 2065
rect 26910 2045 26920 2065
rect 26880 2015 26920 2045
rect 26880 1995 26890 2015
rect 26910 1995 26920 2015
rect 26880 1980 26920 1995
rect 26935 2115 26975 2130
rect 26935 2095 26945 2115
rect 26965 2095 26975 2115
rect 26935 2065 26975 2095
rect 26935 2045 26945 2065
rect 26965 2045 26975 2065
rect 26935 2015 26975 2045
rect 26935 1995 26945 2015
rect 26965 1995 26975 2015
rect 26935 1980 26975 1995
rect 26990 2115 27030 2130
rect 26990 2095 27000 2115
rect 27020 2095 27030 2115
rect 26990 2065 27030 2095
rect 26990 2045 27000 2065
rect 27020 2045 27030 2065
rect 26990 2015 27030 2045
rect 26990 1995 27000 2015
rect 27020 1995 27030 2015
rect 26990 1980 27030 1995
rect 27045 2115 27085 2130
rect 27045 2095 27055 2115
rect 27075 2095 27085 2115
rect 27045 2065 27085 2095
rect 27045 2045 27055 2065
rect 27075 2045 27085 2065
rect 27045 2015 27085 2045
rect 27045 1995 27055 2015
rect 27075 1995 27085 2015
rect 27045 1980 27085 1995
rect 27100 2115 27140 2130
rect 27100 2095 27110 2115
rect 27130 2095 27140 2115
rect 27100 2065 27140 2095
rect 27100 2045 27110 2065
rect 27130 2045 27140 2065
rect 27100 2015 27140 2045
rect 27100 1995 27110 2015
rect 27130 1995 27140 2015
rect 27100 1980 27140 1995
rect 27155 2115 27195 2130
rect 27155 2095 27165 2115
rect 27185 2095 27195 2115
rect 27155 2065 27195 2095
rect 27155 2045 27165 2065
rect 27185 2045 27195 2065
rect 27155 2015 27195 2045
rect 27155 1995 27165 2015
rect 27185 1995 27195 2015
rect 27155 1980 27195 1995
rect 27210 2115 27250 2130
rect 27210 2095 27220 2115
rect 27240 2095 27250 2115
rect 27210 2065 27250 2095
rect 27210 2045 27220 2065
rect 27240 2045 27250 2065
rect 27210 2015 27250 2045
rect 27210 1995 27220 2015
rect 27240 1995 27250 2015
rect 27210 1980 27250 1995
rect 27265 2115 27305 2130
rect 27265 2095 27275 2115
rect 27295 2095 27305 2115
rect 27265 2065 27305 2095
rect 27265 2045 27275 2065
rect 27295 2045 27305 2065
rect 27265 2015 27305 2045
rect 27265 1995 27275 2015
rect 27295 1995 27305 2015
rect 27265 1980 27305 1995
rect 27320 2115 27360 2130
rect 27320 2095 27330 2115
rect 27350 2095 27360 2115
rect 27320 2065 27360 2095
rect 27320 2045 27330 2065
rect 27350 2045 27360 2065
rect 27320 2015 27360 2045
rect 27320 1995 27330 2015
rect 27350 1995 27360 2015
rect 27320 1980 27360 1995
rect 27375 2115 27415 2130
rect 27375 2095 27385 2115
rect 27405 2095 27415 2115
rect 27375 2065 27415 2095
rect 27375 2045 27385 2065
rect 27405 2045 27415 2065
rect 27375 2015 27415 2045
rect 27375 1995 27385 2015
rect 27405 1995 27415 2015
rect 27375 1980 27415 1995
rect 27430 2115 27470 2130
rect 27430 2095 27440 2115
rect 27460 2095 27470 2115
rect 27430 2065 27470 2095
rect 27430 2045 27440 2065
rect 27460 2045 27470 2065
rect 27430 2015 27470 2045
rect 27430 1995 27440 2015
rect 27460 1995 27470 2015
rect 27430 1980 27470 1995
rect 27485 2115 27525 2130
rect 27485 2095 27495 2115
rect 27515 2095 27525 2115
rect 27485 2065 27525 2095
rect 27485 2045 27495 2065
rect 27515 2045 27525 2065
rect 27485 2015 27525 2045
rect 27890 2105 27930 2135
rect 27890 2085 27900 2105
rect 27920 2085 27930 2105
rect 27890 2055 27930 2085
rect 27890 2035 27900 2055
rect 27920 2035 27930 2055
rect 27890 2020 27930 2035
rect 27945 2155 27985 2170
rect 27945 2135 27955 2155
rect 27975 2135 27985 2155
rect 27945 2105 27985 2135
rect 27945 2085 27955 2105
rect 27975 2085 27985 2105
rect 27945 2055 27985 2085
rect 27945 2035 27955 2055
rect 27975 2035 27985 2055
rect 27945 2020 27985 2035
rect 28000 2155 28040 2170
rect 28000 2135 28010 2155
rect 28030 2135 28040 2155
rect 28000 2105 28040 2135
rect 28000 2085 28010 2105
rect 28030 2085 28040 2105
rect 28000 2055 28040 2085
rect 28000 2035 28010 2055
rect 28030 2035 28040 2055
rect 28000 2020 28040 2035
rect 28055 2155 28095 2170
rect 28055 2135 28065 2155
rect 28085 2135 28095 2155
rect 28055 2105 28095 2135
rect 28055 2085 28065 2105
rect 28085 2085 28095 2105
rect 28055 2055 28095 2085
rect 28055 2035 28065 2055
rect 28085 2035 28095 2055
rect 28055 2020 28095 2035
rect 28110 2155 28150 2170
rect 28110 2135 28120 2155
rect 28140 2135 28150 2155
rect 28110 2105 28150 2135
rect 28110 2085 28120 2105
rect 28140 2085 28150 2105
rect 28110 2055 28150 2085
rect 28110 2035 28120 2055
rect 28140 2035 28150 2055
rect 28110 2020 28150 2035
rect 28165 2155 28205 2170
rect 28165 2135 28175 2155
rect 28195 2135 28205 2155
rect 28165 2105 28205 2135
rect 28165 2085 28175 2105
rect 28195 2085 28205 2105
rect 28165 2055 28205 2085
rect 28165 2035 28175 2055
rect 28195 2035 28205 2055
rect 28165 2020 28205 2035
rect 28220 2155 28260 2170
rect 28220 2135 28230 2155
rect 28250 2135 28260 2155
rect 28220 2105 28260 2135
rect 28220 2085 28230 2105
rect 28250 2085 28260 2105
rect 28220 2055 28260 2085
rect 28220 2035 28230 2055
rect 28250 2035 28260 2055
rect 28220 2020 28260 2035
rect 28275 2155 28315 2170
rect 28275 2135 28285 2155
rect 28305 2135 28315 2155
rect 28275 2105 28315 2135
rect 28275 2085 28285 2105
rect 28305 2085 28315 2105
rect 28275 2055 28315 2085
rect 28275 2035 28285 2055
rect 28305 2035 28315 2055
rect 28275 2020 28315 2035
rect 28330 2155 28370 2170
rect 28330 2135 28340 2155
rect 28360 2135 28370 2155
rect 28330 2105 28370 2135
rect 28330 2085 28340 2105
rect 28360 2085 28370 2105
rect 28330 2055 28370 2085
rect 28330 2035 28340 2055
rect 28360 2035 28370 2055
rect 28330 2020 28370 2035
rect 28385 2155 28425 2170
rect 28385 2135 28395 2155
rect 28415 2135 28425 2155
rect 28385 2105 28425 2135
rect 28385 2085 28395 2105
rect 28415 2085 28425 2105
rect 28385 2055 28425 2085
rect 28385 2035 28395 2055
rect 28415 2035 28425 2055
rect 28385 2020 28425 2035
rect 28440 2155 28480 2170
rect 28440 2135 28450 2155
rect 28470 2135 28480 2155
rect 28440 2105 28480 2135
rect 28440 2085 28450 2105
rect 28470 2085 28480 2105
rect 28440 2055 28480 2085
rect 28440 2035 28450 2055
rect 28470 2035 28480 2055
rect 28440 2020 28480 2035
rect 28495 2155 28535 2170
rect 28495 2135 28505 2155
rect 28525 2135 28535 2155
rect 28495 2105 28535 2135
rect 28495 2085 28505 2105
rect 28525 2085 28535 2105
rect 28495 2055 28535 2085
rect 28495 2035 28505 2055
rect 28525 2035 28535 2055
rect 28495 2020 28535 2035
rect 28550 2155 28590 2170
rect 28550 2135 28560 2155
rect 28580 2135 28590 2155
rect 28550 2105 28590 2135
rect 28550 2085 28560 2105
rect 28580 2085 28590 2105
rect 28550 2055 28590 2085
rect 28550 2035 28560 2055
rect 28580 2035 28590 2055
rect 28550 2020 28590 2035
rect 28605 2155 28645 2170
rect 28605 2135 28615 2155
rect 28635 2135 28645 2155
rect 28605 2105 28645 2135
rect 28605 2085 28615 2105
rect 28635 2085 28645 2105
rect 28605 2055 28645 2085
rect 28605 2035 28615 2055
rect 28635 2035 28645 2055
rect 28605 2020 28645 2035
rect 28660 2155 28700 2170
rect 28660 2135 28670 2155
rect 28690 2135 28700 2155
rect 28660 2105 28700 2135
rect 28660 2085 28670 2105
rect 28690 2085 28700 2105
rect 28660 2055 28700 2085
rect 28660 2035 28670 2055
rect 28690 2035 28700 2055
rect 28660 2020 28700 2035
rect 28715 2155 28755 2170
rect 28715 2135 28725 2155
rect 28745 2135 28755 2155
rect 28715 2105 28755 2135
rect 28715 2085 28725 2105
rect 28745 2085 28755 2105
rect 28715 2055 28755 2085
rect 28715 2035 28725 2055
rect 28745 2035 28755 2055
rect 28715 2020 28755 2035
rect 28770 2155 28810 2170
rect 28770 2135 28780 2155
rect 28800 2135 28810 2155
rect 28770 2105 28810 2135
rect 28770 2085 28780 2105
rect 28800 2085 28810 2105
rect 28770 2055 28810 2085
rect 28770 2035 28780 2055
rect 28800 2035 28810 2055
rect 28770 2020 28810 2035
rect 28825 2155 28865 2170
rect 28825 2135 28835 2155
rect 28855 2135 28865 2155
rect 28825 2105 28865 2135
rect 28825 2085 28835 2105
rect 28855 2085 28865 2105
rect 28825 2055 28865 2085
rect 28825 2035 28835 2055
rect 28855 2035 28865 2055
rect 28825 2020 28865 2035
rect 28880 2155 28920 2170
rect 28880 2135 28890 2155
rect 28910 2135 28920 2155
rect 28880 2105 28920 2135
rect 28880 2085 28890 2105
rect 28910 2085 28920 2105
rect 28880 2055 28920 2085
rect 28880 2035 28890 2055
rect 28910 2035 28920 2055
rect 28880 2020 28920 2035
rect 28935 2155 28975 2170
rect 28935 2135 28945 2155
rect 28965 2135 28975 2155
rect 28935 2105 28975 2135
rect 28935 2085 28945 2105
rect 28965 2085 28975 2105
rect 28935 2055 28975 2085
rect 28935 2035 28945 2055
rect 28965 2035 28975 2055
rect 28935 2020 28975 2035
rect 28990 2155 29030 2170
rect 28990 2135 29000 2155
rect 29020 2135 29030 2155
rect 28990 2105 29030 2135
rect 28990 2085 29000 2105
rect 29020 2085 29030 2105
rect 28990 2055 29030 2085
rect 28990 2035 29000 2055
rect 29020 2035 29030 2055
rect 28990 2020 29030 2035
rect 29045 2155 29085 2170
rect 29045 2135 29055 2155
rect 29075 2135 29085 2155
rect 29045 2105 29085 2135
rect 29045 2085 29055 2105
rect 29075 2085 29085 2105
rect 29045 2055 29085 2085
rect 29045 2035 29055 2055
rect 29075 2035 29085 2055
rect 29045 2020 29085 2035
rect 29100 2155 29140 2170
rect 29100 2135 29110 2155
rect 29130 2135 29140 2155
rect 29100 2105 29140 2135
rect 29100 2085 29110 2105
rect 29130 2085 29140 2105
rect 29100 2055 29140 2085
rect 29100 2035 29110 2055
rect 29130 2035 29140 2055
rect 29100 2020 29140 2035
rect 27485 1995 27495 2015
rect 27515 1995 27525 2015
rect 27485 1980 27525 1995
rect 13605 1965 13645 1980
rect 27990 1840 28030 1855
rect 27990 1820 28000 1840
rect 28020 1820 28030 1840
rect 27990 1790 28030 1820
rect 27990 1770 28000 1790
rect 28020 1770 28030 1790
rect 27990 1740 28030 1770
rect 27990 1720 28000 1740
rect 28020 1720 28030 1740
rect 27990 1705 28030 1720
rect 28045 1840 28085 1855
rect 28045 1820 28055 1840
rect 28075 1820 28085 1840
rect 28045 1790 28085 1820
rect 28045 1770 28055 1790
rect 28075 1770 28085 1790
rect 28045 1740 28085 1770
rect 28045 1720 28055 1740
rect 28075 1720 28085 1740
rect 28045 1705 28085 1720
rect 28100 1840 28140 1855
rect 28100 1820 28110 1840
rect 28130 1820 28140 1840
rect 28100 1790 28140 1820
rect 28100 1770 28110 1790
rect 28130 1770 28140 1790
rect 28100 1740 28140 1770
rect 28100 1720 28110 1740
rect 28130 1720 28140 1740
rect 28100 1705 28140 1720
rect 28155 1840 28195 1855
rect 28155 1820 28165 1840
rect 28185 1820 28195 1840
rect 28155 1790 28195 1820
rect 28155 1770 28165 1790
rect 28185 1770 28195 1790
rect 28155 1740 28195 1770
rect 28155 1720 28165 1740
rect 28185 1720 28195 1740
rect 28155 1705 28195 1720
rect 28210 1840 28250 1855
rect 28210 1820 28220 1840
rect 28240 1820 28250 1840
rect 28210 1790 28250 1820
rect 28210 1770 28220 1790
rect 28240 1770 28250 1790
rect 28210 1740 28250 1770
rect 28210 1720 28220 1740
rect 28240 1720 28250 1740
rect 28210 1705 28250 1720
rect 28265 1840 28305 1855
rect 28265 1820 28275 1840
rect 28295 1820 28305 1840
rect 28265 1790 28305 1820
rect 28265 1770 28275 1790
rect 28295 1770 28305 1790
rect 28265 1740 28305 1770
rect 28265 1720 28275 1740
rect 28295 1720 28305 1740
rect 28265 1705 28305 1720
rect 28320 1840 28360 1855
rect 28320 1820 28330 1840
rect 28350 1820 28360 1840
rect 28320 1790 28360 1820
rect 28320 1770 28330 1790
rect 28350 1770 28360 1790
rect 28320 1740 28360 1770
rect 28320 1720 28330 1740
rect 28350 1720 28360 1740
rect 28320 1705 28360 1720
rect 3165 1650 3205 1665
rect 3165 1630 3175 1650
rect 3195 1630 3205 1650
rect 3165 1615 3205 1630
rect 3225 1650 3265 1665
rect 3225 1630 3235 1650
rect 3255 1630 3265 1650
rect 3225 1615 3265 1630
rect 3285 1650 3325 1665
rect 3285 1630 3295 1650
rect 3315 1630 3325 1650
rect 3285 1615 3325 1630
rect 3345 1650 3385 1665
rect 3345 1630 3355 1650
rect 3375 1630 3385 1650
rect 3345 1615 3385 1630
rect 3405 1650 3445 1665
rect 3405 1630 3415 1650
rect 3435 1630 3445 1650
rect 3405 1615 3445 1630
rect 3465 1650 3505 1665
rect 3465 1630 3475 1650
rect 3495 1630 3505 1650
rect 3465 1615 3505 1630
rect 3525 1650 3565 1665
rect 3525 1630 3535 1650
rect 3555 1630 3565 1650
rect 3525 1615 3565 1630
rect 3585 1650 3625 1665
rect 3585 1630 3595 1650
rect 3615 1630 3625 1650
rect 3585 1615 3625 1630
rect 3645 1650 3685 1665
rect 3645 1630 3655 1650
rect 3675 1630 3685 1650
rect 3645 1615 3685 1630
rect 3705 1650 3745 1665
rect 3705 1630 3715 1650
rect 3735 1630 3745 1650
rect 3705 1615 3745 1630
rect 3765 1650 3805 1665
rect 3765 1630 3775 1650
rect 3795 1630 3805 1650
rect 3765 1615 3805 1630
rect 4205 1650 4245 1665
rect 4205 1630 4215 1650
rect 4235 1630 4245 1650
rect 4205 1615 4245 1630
rect 4265 1650 4305 1665
rect 4265 1630 4275 1650
rect 4295 1630 4305 1650
rect 4265 1615 4305 1630
rect 4325 1650 4365 1665
rect 4325 1630 4335 1650
rect 4355 1630 4365 1650
rect 4325 1615 4365 1630
rect 4385 1650 4425 1665
rect 4385 1630 4395 1650
rect 4415 1630 4425 1650
rect 4385 1615 4425 1630
rect 4445 1650 4485 1665
rect 4445 1630 4455 1650
rect 4475 1630 4485 1650
rect 4445 1615 4485 1630
rect 4505 1650 4545 1665
rect 4505 1630 4515 1650
rect 4535 1630 4545 1650
rect 4505 1615 4545 1630
rect 4565 1650 4605 1665
rect 4565 1630 4575 1650
rect 4595 1630 4605 1650
rect 4565 1615 4605 1630
rect 4625 1650 4665 1665
rect 4625 1630 4635 1650
rect 4655 1630 4665 1650
rect 4625 1615 4665 1630
rect 4685 1650 4725 1665
rect 4685 1630 4695 1650
rect 4715 1630 4725 1650
rect 4685 1615 4725 1630
rect 4745 1650 4785 1665
rect 4745 1630 4755 1650
rect 4775 1630 4785 1650
rect 4745 1615 4785 1630
rect 4805 1650 4845 1665
rect 4805 1630 4815 1650
rect 4835 1630 4845 1650
rect 4805 1615 4845 1630
rect 10155 1640 10195 1655
rect 10155 1620 10165 1640
rect 10185 1620 10195 1640
rect 2835 1440 2875 1455
rect 2835 1420 2845 1440
rect 2865 1420 2875 1440
rect 2835 1390 2875 1420
rect 2835 1370 2845 1390
rect 2865 1370 2875 1390
rect 2835 1340 2875 1370
rect 2835 1320 2845 1340
rect 2865 1320 2875 1340
rect 2835 1290 2875 1320
rect 2835 1270 2845 1290
rect 2865 1270 2875 1290
rect 2835 1240 2875 1270
rect 2835 1220 2845 1240
rect 2865 1220 2875 1240
rect 2835 1205 2875 1220
rect 3375 1440 3415 1455
rect 3375 1420 3385 1440
rect 3405 1420 3415 1440
rect 3375 1390 3415 1420
rect 3375 1370 3385 1390
rect 3405 1370 3415 1390
rect 3375 1340 3415 1370
rect 3375 1320 3385 1340
rect 3405 1320 3415 1340
rect 3375 1290 3415 1320
rect 3375 1270 3385 1290
rect 3405 1270 3415 1290
rect 3375 1240 3415 1270
rect 3375 1220 3385 1240
rect 3405 1220 3415 1240
rect 3375 1205 3415 1220
rect 3915 1440 3955 1455
rect 3915 1420 3925 1440
rect 3945 1420 3955 1440
rect 3915 1390 3955 1420
rect 3915 1370 3925 1390
rect 3945 1370 3955 1390
rect 3915 1340 3955 1370
rect 3915 1320 3925 1340
rect 3945 1320 3955 1340
rect 3915 1290 3955 1320
rect 3915 1270 3925 1290
rect 3945 1270 3955 1290
rect 3915 1240 3955 1270
rect 3915 1220 3925 1240
rect 3945 1220 3955 1240
rect 3915 1205 3955 1220
rect 4055 1440 4095 1455
rect 4055 1420 4065 1440
rect 4085 1420 4095 1440
rect 4055 1390 4095 1420
rect 4055 1370 4065 1390
rect 4085 1370 4095 1390
rect 4055 1340 4095 1370
rect 4055 1320 4065 1340
rect 4085 1320 4095 1340
rect 4055 1290 4095 1320
rect 4055 1270 4065 1290
rect 4085 1270 4095 1290
rect 4055 1240 4095 1270
rect 4055 1220 4065 1240
rect 4085 1220 4095 1240
rect 4055 1205 4095 1220
rect 4595 1440 4635 1455
rect 4595 1420 4605 1440
rect 4625 1420 4635 1440
rect 4595 1390 4635 1420
rect 4595 1370 4605 1390
rect 4625 1370 4635 1390
rect 4595 1340 4635 1370
rect 4595 1320 4605 1340
rect 4625 1320 4635 1340
rect 4595 1290 4635 1320
rect 4595 1270 4605 1290
rect 4625 1270 4635 1290
rect 4595 1240 4635 1270
rect 4595 1220 4605 1240
rect 4625 1220 4635 1240
rect 4595 1205 4635 1220
rect 5135 1440 5175 1455
rect 5135 1420 5145 1440
rect 5165 1420 5175 1440
rect 5135 1390 5175 1420
rect 5135 1370 5145 1390
rect 5165 1370 5175 1390
rect 5135 1340 5175 1370
rect 5135 1320 5145 1340
rect 5165 1320 5175 1340
rect 5135 1290 5175 1320
rect 5135 1270 5145 1290
rect 5165 1270 5175 1290
rect 5135 1240 5175 1270
rect 5135 1220 5145 1240
rect 5165 1220 5175 1240
rect 5135 1205 5175 1220
rect 2945 1060 2985 1075
rect 2945 1040 2955 1060
rect 2975 1040 2985 1060
rect 2945 1010 2985 1040
rect 2945 990 2955 1010
rect 2975 990 2985 1010
rect 2945 975 2985 990
rect 3985 1060 4025 1075
rect 3985 1040 3995 1060
rect 4015 1040 4025 1060
rect 3985 1010 4025 1040
rect 3985 990 3995 1010
rect 4015 990 4025 1010
rect 3985 975 4025 990
rect 5025 1060 5065 1075
rect 5025 1040 5035 1060
rect 5055 1040 5065 1060
rect 5025 1010 5065 1040
rect 5025 990 5035 1010
rect 5055 990 5065 1010
rect 5025 975 5065 990
rect 10155 1590 10195 1620
rect 10155 1570 10165 1590
rect 10185 1570 10195 1590
rect 10155 1540 10195 1570
rect 10155 1520 10165 1540
rect 10185 1520 10195 1540
rect 10155 1490 10195 1520
rect 10155 1470 10165 1490
rect 10185 1470 10195 1490
rect 10155 1440 10195 1470
rect 10155 1420 10165 1440
rect 10185 1420 10195 1440
rect 10155 1390 10195 1420
rect 10155 1370 10165 1390
rect 10185 1370 10195 1390
rect 10155 1340 10195 1370
rect 10155 1320 10165 1340
rect 10185 1320 10195 1340
rect 10155 1290 10195 1320
rect 10155 1270 10165 1290
rect 10185 1270 10195 1290
rect 10155 1240 10195 1270
rect 10155 1220 10165 1240
rect 10185 1220 10195 1240
rect 10155 1190 10195 1220
rect 10155 1170 10165 1190
rect 10185 1170 10195 1190
rect 10155 1140 10195 1170
rect 10155 1120 10165 1140
rect 10185 1120 10195 1140
rect 10155 1090 10195 1120
rect 10155 1070 10165 1090
rect 10185 1070 10195 1090
rect 10155 1040 10195 1070
rect 10155 1020 10165 1040
rect 10185 1020 10195 1040
rect 10155 990 10195 1020
rect 10155 970 10165 990
rect 10185 970 10195 990
rect 10155 955 10195 970
rect 10255 1640 10295 1655
rect 10255 1620 10265 1640
rect 10285 1620 10295 1640
rect 10255 1590 10295 1620
rect 10255 1570 10265 1590
rect 10285 1570 10295 1590
rect 10255 1540 10295 1570
rect 10255 1520 10265 1540
rect 10285 1520 10295 1540
rect 10255 1490 10295 1520
rect 10255 1470 10265 1490
rect 10285 1470 10295 1490
rect 10255 1440 10295 1470
rect 10255 1420 10265 1440
rect 10285 1420 10295 1440
rect 10255 1390 10295 1420
rect 10255 1370 10265 1390
rect 10285 1370 10295 1390
rect 10255 1340 10295 1370
rect 10255 1320 10265 1340
rect 10285 1320 10295 1340
rect 10255 1290 10295 1320
rect 10255 1270 10265 1290
rect 10285 1270 10295 1290
rect 10255 1240 10295 1270
rect 10255 1220 10265 1240
rect 10285 1220 10295 1240
rect 10255 1190 10295 1220
rect 10255 1170 10265 1190
rect 10285 1170 10295 1190
rect 10255 1140 10295 1170
rect 10255 1120 10265 1140
rect 10285 1120 10295 1140
rect 10255 1090 10295 1120
rect 10255 1070 10265 1090
rect 10285 1070 10295 1090
rect 10255 1040 10295 1070
rect 10255 1020 10265 1040
rect 10285 1020 10295 1040
rect 10255 990 10295 1020
rect 10255 970 10265 990
rect 10285 970 10295 990
rect 10255 955 10295 970
rect 10355 1640 10395 1655
rect 10355 1620 10365 1640
rect 10385 1620 10395 1640
rect 10355 1590 10395 1620
rect 10355 1570 10365 1590
rect 10385 1570 10395 1590
rect 10355 1540 10395 1570
rect 10355 1520 10365 1540
rect 10385 1520 10395 1540
rect 10355 1490 10395 1520
rect 10355 1470 10365 1490
rect 10385 1470 10395 1490
rect 10355 1440 10395 1470
rect 10355 1420 10365 1440
rect 10385 1420 10395 1440
rect 10355 1390 10395 1420
rect 10355 1370 10365 1390
rect 10385 1370 10395 1390
rect 10355 1340 10395 1370
rect 10355 1320 10365 1340
rect 10385 1320 10395 1340
rect 10355 1290 10395 1320
rect 10355 1270 10365 1290
rect 10385 1270 10395 1290
rect 10355 1240 10395 1270
rect 10355 1220 10365 1240
rect 10385 1220 10395 1240
rect 10355 1190 10395 1220
rect 10355 1170 10365 1190
rect 10385 1170 10395 1190
rect 10355 1140 10395 1170
rect 10355 1120 10365 1140
rect 10385 1120 10395 1140
rect 10355 1090 10395 1120
rect 10355 1070 10365 1090
rect 10385 1070 10395 1090
rect 10355 1040 10395 1070
rect 10355 1020 10365 1040
rect 10385 1020 10395 1040
rect 10355 990 10395 1020
rect 10355 970 10365 990
rect 10385 970 10395 990
rect 10355 955 10395 970
rect 10455 1640 10495 1655
rect 10455 1620 10465 1640
rect 10485 1620 10495 1640
rect 10455 1590 10495 1620
rect 10455 1570 10465 1590
rect 10485 1570 10495 1590
rect 10455 1540 10495 1570
rect 10455 1520 10465 1540
rect 10485 1520 10495 1540
rect 10455 1490 10495 1520
rect 10455 1470 10465 1490
rect 10485 1470 10495 1490
rect 10455 1440 10495 1470
rect 10455 1420 10465 1440
rect 10485 1420 10495 1440
rect 10455 1390 10495 1420
rect 10455 1370 10465 1390
rect 10485 1370 10495 1390
rect 10455 1340 10495 1370
rect 10455 1320 10465 1340
rect 10485 1320 10495 1340
rect 10455 1290 10495 1320
rect 10455 1270 10465 1290
rect 10485 1270 10495 1290
rect 10455 1240 10495 1270
rect 10455 1220 10465 1240
rect 10485 1220 10495 1240
rect 10455 1190 10495 1220
rect 10455 1170 10465 1190
rect 10485 1170 10495 1190
rect 10455 1140 10495 1170
rect 10455 1120 10465 1140
rect 10485 1120 10495 1140
rect 10455 1090 10495 1120
rect 10455 1070 10465 1090
rect 10485 1070 10495 1090
rect 10455 1040 10495 1070
rect 10455 1020 10465 1040
rect 10485 1020 10495 1040
rect 10455 990 10495 1020
rect 10455 970 10465 990
rect 10485 970 10495 990
rect 10455 955 10495 970
rect 10555 1640 10595 1655
rect 10555 1620 10565 1640
rect 10585 1620 10595 1640
rect 10555 1590 10595 1620
rect 10555 1570 10565 1590
rect 10585 1570 10595 1590
rect 10555 1540 10595 1570
rect 10555 1520 10565 1540
rect 10585 1520 10595 1540
rect 10555 1490 10595 1520
rect 10555 1470 10565 1490
rect 10585 1470 10595 1490
rect 10555 1440 10595 1470
rect 10555 1420 10565 1440
rect 10585 1420 10595 1440
rect 10555 1390 10595 1420
rect 10555 1370 10565 1390
rect 10585 1370 10595 1390
rect 10555 1340 10595 1370
rect 10555 1320 10565 1340
rect 10585 1320 10595 1340
rect 10555 1290 10595 1320
rect 10555 1270 10565 1290
rect 10585 1270 10595 1290
rect 10555 1240 10595 1270
rect 10555 1220 10565 1240
rect 10585 1220 10595 1240
rect 10555 1190 10595 1220
rect 10555 1170 10565 1190
rect 10585 1170 10595 1190
rect 10555 1140 10595 1170
rect 10555 1120 10565 1140
rect 10585 1120 10595 1140
rect 10555 1090 10595 1120
rect 10555 1070 10565 1090
rect 10585 1070 10595 1090
rect 10555 1040 10595 1070
rect 10555 1020 10565 1040
rect 10585 1020 10595 1040
rect 10555 990 10595 1020
rect 10555 970 10565 990
rect 10585 970 10595 990
rect 10555 955 10595 970
rect 10655 1640 10695 1655
rect 10655 1620 10665 1640
rect 10685 1620 10695 1640
rect 10655 1590 10695 1620
rect 10655 1570 10665 1590
rect 10685 1570 10695 1590
rect 10655 1540 10695 1570
rect 10655 1520 10665 1540
rect 10685 1520 10695 1540
rect 10655 1490 10695 1520
rect 10655 1470 10665 1490
rect 10685 1470 10695 1490
rect 10655 1440 10695 1470
rect 10655 1420 10665 1440
rect 10685 1420 10695 1440
rect 10655 1390 10695 1420
rect 10655 1370 10665 1390
rect 10685 1370 10695 1390
rect 10655 1340 10695 1370
rect 10655 1320 10665 1340
rect 10685 1320 10695 1340
rect 10655 1290 10695 1320
rect 10655 1270 10665 1290
rect 10685 1270 10695 1290
rect 10655 1240 10695 1270
rect 10655 1220 10665 1240
rect 10685 1220 10695 1240
rect 10655 1190 10695 1220
rect 10655 1170 10665 1190
rect 10685 1170 10695 1190
rect 10655 1140 10695 1170
rect 10655 1120 10665 1140
rect 10685 1120 10695 1140
rect 10655 1090 10695 1120
rect 10655 1070 10665 1090
rect 10685 1070 10695 1090
rect 10655 1040 10695 1070
rect 10655 1020 10665 1040
rect 10685 1020 10695 1040
rect 10655 990 10695 1020
rect 10655 970 10665 990
rect 10685 970 10695 990
rect 10655 955 10695 970
rect 10755 1640 10795 1655
rect 10755 1620 10765 1640
rect 10785 1620 10795 1640
rect 10755 1590 10795 1620
rect 10755 1570 10765 1590
rect 10785 1570 10795 1590
rect 10755 1540 10795 1570
rect 10755 1520 10765 1540
rect 10785 1520 10795 1540
rect 10755 1490 10795 1520
rect 11030 1650 11070 1665
rect 11030 1630 11040 1650
rect 11060 1630 11070 1650
rect 11030 1600 11070 1630
rect 11030 1580 11040 1600
rect 11060 1580 11070 1600
rect 11030 1550 11070 1580
rect 11030 1530 11040 1550
rect 11060 1530 11070 1550
rect 11030 1515 11070 1530
rect 11085 1650 11125 1665
rect 11085 1630 11095 1650
rect 11115 1630 11125 1650
rect 11085 1600 11125 1630
rect 11085 1580 11095 1600
rect 11115 1580 11125 1600
rect 11085 1550 11125 1580
rect 11085 1530 11095 1550
rect 11115 1530 11125 1550
rect 11085 1515 11125 1530
rect 11140 1650 11180 1665
rect 11140 1630 11150 1650
rect 11170 1630 11180 1650
rect 11140 1600 11180 1630
rect 11140 1580 11150 1600
rect 11170 1580 11180 1600
rect 11140 1550 11180 1580
rect 11140 1530 11150 1550
rect 11170 1530 11180 1550
rect 11140 1515 11180 1530
rect 11195 1650 11235 1665
rect 11195 1630 11205 1650
rect 11225 1630 11235 1650
rect 11195 1600 11235 1630
rect 11195 1580 11205 1600
rect 11225 1580 11235 1600
rect 11195 1550 11235 1580
rect 11195 1530 11205 1550
rect 11225 1530 11235 1550
rect 11195 1515 11235 1530
rect 11250 1650 11290 1665
rect 11250 1630 11260 1650
rect 11280 1630 11290 1650
rect 11250 1600 11290 1630
rect 11250 1580 11260 1600
rect 11280 1580 11290 1600
rect 11250 1550 11290 1580
rect 11250 1530 11260 1550
rect 11280 1530 11290 1550
rect 11250 1515 11290 1530
rect 11305 1650 11345 1665
rect 11305 1630 11315 1650
rect 11335 1630 11345 1650
rect 11305 1600 11345 1630
rect 11305 1580 11315 1600
rect 11335 1580 11345 1600
rect 11305 1550 11345 1580
rect 11305 1530 11315 1550
rect 11335 1530 11345 1550
rect 11305 1515 11345 1530
rect 11360 1650 11400 1665
rect 11360 1630 11370 1650
rect 11390 1630 11400 1650
rect 11360 1600 11400 1630
rect 11360 1580 11370 1600
rect 11390 1580 11400 1600
rect 11360 1550 11400 1580
rect 11360 1530 11370 1550
rect 11390 1530 11400 1550
rect 11360 1515 11400 1530
rect 11415 1650 11455 1665
rect 11415 1630 11425 1650
rect 11445 1630 11455 1650
rect 11415 1600 11455 1630
rect 11415 1580 11425 1600
rect 11445 1580 11455 1600
rect 11415 1550 11455 1580
rect 11415 1530 11425 1550
rect 11445 1530 11455 1550
rect 11415 1515 11455 1530
rect 11470 1650 11510 1665
rect 11470 1630 11480 1650
rect 11500 1630 11510 1650
rect 11470 1600 11510 1630
rect 11470 1580 11480 1600
rect 11500 1580 11510 1600
rect 11470 1550 11510 1580
rect 11470 1530 11480 1550
rect 11500 1530 11510 1550
rect 11470 1515 11510 1530
rect 11525 1650 11565 1665
rect 11525 1630 11535 1650
rect 11555 1630 11565 1650
rect 11525 1600 11565 1630
rect 11525 1580 11535 1600
rect 11555 1580 11565 1600
rect 11525 1550 11565 1580
rect 11525 1530 11535 1550
rect 11555 1530 11565 1550
rect 11525 1515 11565 1530
rect 11580 1650 11620 1665
rect 11580 1630 11590 1650
rect 11610 1630 11620 1650
rect 11580 1600 11620 1630
rect 11580 1580 11590 1600
rect 11610 1580 11620 1600
rect 11580 1550 11620 1580
rect 11580 1530 11590 1550
rect 11610 1530 11620 1550
rect 11580 1515 11620 1530
rect 11635 1650 11675 1665
rect 11635 1630 11645 1650
rect 11665 1630 11675 1650
rect 11635 1600 11675 1630
rect 11635 1580 11645 1600
rect 11665 1580 11675 1600
rect 11635 1550 11675 1580
rect 11635 1530 11645 1550
rect 11665 1530 11675 1550
rect 11635 1515 11675 1530
rect 11690 1650 11730 1665
rect 11770 1650 11810 1665
rect 11690 1630 11700 1650
rect 11720 1630 11730 1650
rect 11770 1630 11780 1650
rect 11800 1630 11810 1650
rect 11690 1600 11730 1630
rect 11770 1600 11810 1630
rect 11690 1580 11700 1600
rect 11720 1580 11730 1600
rect 11770 1580 11780 1600
rect 11800 1580 11810 1600
rect 11690 1550 11730 1580
rect 11770 1550 11810 1580
rect 11690 1530 11700 1550
rect 11720 1530 11730 1550
rect 11770 1530 11780 1550
rect 11800 1530 11810 1550
rect 11690 1515 11730 1530
rect 11770 1515 11810 1530
rect 11825 1650 11865 1665
rect 11825 1630 11835 1650
rect 11855 1630 11865 1650
rect 11825 1600 11865 1630
rect 11825 1580 11835 1600
rect 11855 1580 11865 1600
rect 11825 1550 11865 1580
rect 11825 1530 11835 1550
rect 11855 1530 11865 1550
rect 11825 1515 11865 1530
rect 11880 1650 11920 1665
rect 11880 1630 11890 1650
rect 11910 1630 11920 1650
rect 11880 1600 11920 1630
rect 11880 1580 11890 1600
rect 11910 1580 11920 1600
rect 11880 1550 11920 1580
rect 11880 1530 11890 1550
rect 11910 1530 11920 1550
rect 11880 1515 11920 1530
rect 11935 1650 11975 1665
rect 11935 1630 11945 1650
rect 11965 1630 11975 1650
rect 11935 1600 11975 1630
rect 11935 1580 11945 1600
rect 11965 1580 11975 1600
rect 11935 1550 11975 1580
rect 11935 1530 11945 1550
rect 11965 1530 11975 1550
rect 11935 1515 11975 1530
rect 11990 1650 12030 1665
rect 12070 1650 12110 1665
rect 11990 1630 12000 1650
rect 12020 1630 12030 1650
rect 12070 1630 12080 1650
rect 12100 1630 12110 1650
rect 11990 1600 12030 1630
rect 12070 1600 12110 1630
rect 11990 1580 12000 1600
rect 12020 1580 12030 1600
rect 12070 1580 12080 1600
rect 12100 1580 12110 1600
rect 11990 1550 12030 1580
rect 12070 1550 12110 1580
rect 11990 1530 12000 1550
rect 12020 1530 12030 1550
rect 12070 1530 12080 1550
rect 12100 1530 12110 1550
rect 11990 1515 12030 1530
rect 12070 1515 12110 1530
rect 12125 1650 12165 1665
rect 12125 1630 12135 1650
rect 12155 1630 12165 1650
rect 12125 1600 12165 1630
rect 12125 1580 12135 1600
rect 12155 1580 12165 1600
rect 12125 1550 12165 1580
rect 12125 1530 12135 1550
rect 12155 1530 12165 1550
rect 12125 1515 12165 1530
rect 12180 1650 12220 1665
rect 12180 1630 12190 1650
rect 12210 1630 12220 1650
rect 12180 1600 12220 1630
rect 12180 1580 12190 1600
rect 12210 1580 12220 1600
rect 12180 1550 12220 1580
rect 12180 1530 12190 1550
rect 12210 1530 12220 1550
rect 12180 1515 12220 1530
rect 12235 1650 12275 1665
rect 12235 1630 12245 1650
rect 12265 1630 12275 1650
rect 12235 1600 12275 1630
rect 12235 1580 12245 1600
rect 12265 1580 12275 1600
rect 12235 1550 12275 1580
rect 12235 1530 12245 1550
rect 12265 1530 12275 1550
rect 12235 1515 12275 1530
rect 12290 1650 12330 1665
rect 12290 1630 12300 1650
rect 12320 1630 12330 1650
rect 12290 1600 12330 1630
rect 12290 1580 12300 1600
rect 12320 1580 12330 1600
rect 12290 1550 12330 1580
rect 12290 1530 12300 1550
rect 12320 1530 12330 1550
rect 12290 1515 12330 1530
rect 12345 1650 12385 1665
rect 12345 1630 12355 1650
rect 12375 1630 12385 1650
rect 12345 1600 12385 1630
rect 12345 1580 12355 1600
rect 12375 1580 12385 1600
rect 12345 1550 12385 1580
rect 12345 1530 12355 1550
rect 12375 1530 12385 1550
rect 12345 1515 12385 1530
rect 12400 1650 12440 1665
rect 12400 1630 12410 1650
rect 12430 1630 12440 1650
rect 12400 1600 12440 1630
rect 12400 1580 12410 1600
rect 12430 1580 12440 1600
rect 12400 1550 12440 1580
rect 12400 1530 12410 1550
rect 12430 1530 12440 1550
rect 12400 1515 12440 1530
rect 12455 1650 12495 1665
rect 12455 1630 12465 1650
rect 12485 1630 12495 1650
rect 12455 1600 12495 1630
rect 12455 1580 12465 1600
rect 12485 1580 12495 1600
rect 12455 1550 12495 1580
rect 12455 1530 12465 1550
rect 12485 1530 12495 1550
rect 12455 1515 12495 1530
rect 12510 1650 12550 1665
rect 12510 1630 12520 1650
rect 12540 1630 12550 1650
rect 12510 1600 12550 1630
rect 12510 1580 12520 1600
rect 12540 1580 12550 1600
rect 12510 1550 12550 1580
rect 12510 1530 12520 1550
rect 12540 1530 12550 1550
rect 12510 1515 12550 1530
rect 12565 1650 12605 1665
rect 12565 1630 12575 1650
rect 12595 1630 12605 1650
rect 12565 1600 12605 1630
rect 12565 1580 12575 1600
rect 12595 1580 12605 1600
rect 12565 1550 12605 1580
rect 12565 1530 12575 1550
rect 12595 1530 12605 1550
rect 12565 1515 12605 1530
rect 12620 1650 12660 1665
rect 12620 1630 12630 1650
rect 12650 1630 12660 1650
rect 12620 1600 12660 1630
rect 12620 1580 12630 1600
rect 12650 1580 12660 1600
rect 12620 1550 12660 1580
rect 12620 1530 12630 1550
rect 12650 1530 12660 1550
rect 12620 1515 12660 1530
rect 12675 1650 12715 1665
rect 12675 1630 12685 1650
rect 12705 1630 12715 1650
rect 12675 1600 12715 1630
rect 12675 1580 12685 1600
rect 12705 1580 12715 1600
rect 12675 1550 12715 1580
rect 12675 1530 12685 1550
rect 12705 1530 12715 1550
rect 12675 1515 12715 1530
rect 12730 1650 12770 1665
rect 12730 1630 12740 1650
rect 12760 1630 12770 1650
rect 12730 1600 12770 1630
rect 12730 1580 12740 1600
rect 12760 1580 12770 1600
rect 12730 1550 12770 1580
rect 12730 1530 12740 1550
rect 12760 1530 12770 1550
rect 12730 1515 12770 1530
rect 13005 1640 13045 1655
rect 13005 1620 13015 1640
rect 13035 1620 13045 1640
rect 13005 1590 13045 1620
rect 13005 1570 13015 1590
rect 13035 1570 13045 1590
rect 13005 1540 13045 1570
rect 13005 1520 13015 1540
rect 13035 1520 13045 1540
rect 10755 1470 10765 1490
rect 10785 1470 10795 1490
rect 10755 1440 10795 1470
rect 13005 1490 13045 1520
rect 13005 1470 13015 1490
rect 13035 1470 13045 1490
rect 10755 1420 10765 1440
rect 10785 1420 10795 1440
rect 10755 1390 10795 1420
rect 10755 1370 10765 1390
rect 10785 1370 10795 1390
rect 10755 1340 10795 1370
rect 10755 1320 10765 1340
rect 10785 1320 10795 1340
rect 10755 1290 10795 1320
rect 10755 1270 10765 1290
rect 10785 1270 10795 1290
rect 10755 1240 10795 1270
rect 13005 1440 13045 1470
rect 13005 1420 13015 1440
rect 13035 1420 13045 1440
rect 13005 1390 13045 1420
rect 13005 1370 13015 1390
rect 13035 1370 13045 1390
rect 13005 1340 13045 1370
rect 13005 1320 13015 1340
rect 13035 1320 13045 1340
rect 13005 1290 13045 1320
rect 13005 1270 13015 1290
rect 13035 1270 13045 1290
rect 10755 1220 10765 1240
rect 10785 1220 10795 1240
rect 10755 1190 10795 1220
rect 10755 1170 10765 1190
rect 10785 1170 10795 1190
rect 13005 1240 13045 1270
rect 13005 1220 13015 1240
rect 13035 1220 13045 1240
rect 13005 1190 13045 1220
rect 10755 1140 10795 1170
rect 10755 1120 10765 1140
rect 10785 1120 10795 1140
rect 10755 1090 10795 1120
rect 10755 1070 10765 1090
rect 10785 1070 10795 1090
rect 10755 1040 10795 1070
rect 10755 1020 10765 1040
rect 10785 1020 10795 1040
rect 10755 990 10795 1020
rect 10755 970 10765 990
rect 10785 970 10795 990
rect 10755 955 10795 970
rect 11205 1170 11245 1185
rect 11205 1150 11215 1170
rect 11235 1150 11245 1170
rect 11205 1120 11245 1150
rect 11205 1100 11215 1120
rect 11235 1100 11245 1120
rect 11205 1070 11245 1100
rect 11205 1050 11215 1070
rect 11235 1050 11245 1070
rect 11205 1020 11245 1050
rect 11205 1000 11215 1020
rect 11235 1000 11245 1020
rect 11205 970 11245 1000
rect 11205 950 11215 970
rect 11235 950 11245 970
rect 11205 935 11245 950
rect 11260 1170 11300 1185
rect 11260 1150 11270 1170
rect 11290 1150 11300 1170
rect 11260 1120 11300 1150
rect 11260 1100 11270 1120
rect 11290 1100 11300 1120
rect 11260 1070 11300 1100
rect 11260 1050 11270 1070
rect 11290 1050 11300 1070
rect 11260 1020 11300 1050
rect 11260 1000 11270 1020
rect 11290 1000 11300 1020
rect 11260 970 11300 1000
rect 11260 950 11270 970
rect 11290 950 11300 970
rect 11260 935 11300 950
rect 11315 1170 11355 1185
rect 11315 1150 11325 1170
rect 11345 1150 11355 1170
rect 11315 1120 11355 1150
rect 11315 1100 11325 1120
rect 11345 1100 11355 1120
rect 11315 1070 11355 1100
rect 11315 1050 11325 1070
rect 11345 1050 11355 1070
rect 11315 1020 11355 1050
rect 11315 1000 11325 1020
rect 11345 1000 11355 1020
rect 11315 970 11355 1000
rect 11315 950 11325 970
rect 11345 950 11355 970
rect 11315 935 11355 950
rect 11370 1170 11410 1185
rect 11370 1150 11380 1170
rect 11400 1150 11410 1170
rect 11370 1120 11410 1150
rect 11370 1100 11380 1120
rect 11400 1100 11410 1120
rect 11370 1070 11410 1100
rect 11370 1050 11380 1070
rect 11400 1050 11410 1070
rect 11370 1020 11410 1050
rect 11370 1000 11380 1020
rect 11400 1000 11410 1020
rect 11370 970 11410 1000
rect 11370 950 11380 970
rect 11400 950 11410 970
rect 11370 935 11410 950
rect 11425 1170 11465 1185
rect 11425 1150 11435 1170
rect 11455 1150 11465 1170
rect 11425 1120 11465 1150
rect 11425 1100 11435 1120
rect 11455 1100 11465 1120
rect 11425 1070 11465 1100
rect 11425 1050 11435 1070
rect 11455 1050 11465 1070
rect 11425 1020 11465 1050
rect 11425 1000 11435 1020
rect 11455 1000 11465 1020
rect 11425 970 11465 1000
rect 11425 950 11435 970
rect 11455 950 11465 970
rect 11425 935 11465 950
rect 11480 1170 11520 1185
rect 11480 1150 11490 1170
rect 11510 1150 11520 1170
rect 11480 1120 11520 1150
rect 11480 1100 11490 1120
rect 11510 1100 11520 1120
rect 11480 1070 11520 1100
rect 11480 1050 11490 1070
rect 11510 1050 11520 1070
rect 11480 1020 11520 1050
rect 11480 1000 11490 1020
rect 11510 1000 11520 1020
rect 11480 970 11520 1000
rect 11480 950 11490 970
rect 11510 950 11520 970
rect 11480 935 11520 950
rect 11535 1170 11575 1185
rect 11535 1150 11545 1170
rect 11565 1150 11575 1170
rect 11535 1120 11575 1150
rect 11535 1100 11545 1120
rect 11565 1100 11575 1120
rect 11535 1070 11575 1100
rect 11535 1050 11545 1070
rect 11565 1050 11575 1070
rect 11535 1020 11575 1050
rect 11535 1000 11545 1020
rect 11565 1000 11575 1020
rect 11535 970 11575 1000
rect 11535 950 11545 970
rect 11565 950 11575 970
rect 11535 935 11575 950
rect 11590 1170 11630 1185
rect 11590 1150 11600 1170
rect 11620 1150 11630 1170
rect 11590 1120 11630 1150
rect 11590 1100 11600 1120
rect 11620 1100 11630 1120
rect 11590 1070 11630 1100
rect 11590 1050 11600 1070
rect 11620 1050 11630 1070
rect 11590 1020 11630 1050
rect 11590 1000 11600 1020
rect 11620 1000 11630 1020
rect 11590 970 11630 1000
rect 11590 950 11600 970
rect 11620 950 11630 970
rect 11590 935 11630 950
rect 11645 1170 11685 1185
rect 11645 1150 11655 1170
rect 11675 1150 11685 1170
rect 11645 1120 11685 1150
rect 11645 1100 11655 1120
rect 11675 1100 11685 1120
rect 11645 1070 11685 1100
rect 11645 1050 11655 1070
rect 11675 1050 11685 1070
rect 11645 1020 11685 1050
rect 11645 1000 11655 1020
rect 11675 1000 11685 1020
rect 11645 970 11685 1000
rect 11645 950 11655 970
rect 11675 950 11685 970
rect 11645 935 11685 950
rect 11700 1170 11740 1185
rect 11700 1150 11710 1170
rect 11730 1150 11740 1170
rect 11700 1120 11740 1150
rect 11700 1100 11710 1120
rect 11730 1100 11740 1120
rect 11700 1070 11740 1100
rect 11700 1050 11710 1070
rect 11730 1050 11740 1070
rect 11700 1020 11740 1050
rect 11700 1000 11710 1020
rect 11730 1000 11740 1020
rect 11700 970 11740 1000
rect 11700 950 11710 970
rect 11730 950 11740 970
rect 11700 935 11740 950
rect 11755 1170 11795 1185
rect 11755 1150 11765 1170
rect 11785 1150 11795 1170
rect 11755 1120 11795 1150
rect 11755 1100 11765 1120
rect 11785 1100 11795 1120
rect 11755 1070 11795 1100
rect 11755 1050 11765 1070
rect 11785 1050 11795 1070
rect 11755 1020 11795 1050
rect 11755 1000 11765 1020
rect 11785 1000 11795 1020
rect 11755 970 11795 1000
rect 11755 950 11765 970
rect 11785 950 11795 970
rect 11755 935 11795 950
rect 11810 1170 11850 1185
rect 11810 1150 11820 1170
rect 11840 1150 11850 1170
rect 11810 1120 11850 1150
rect 11810 1100 11820 1120
rect 11840 1100 11850 1120
rect 11810 1070 11850 1100
rect 11810 1050 11820 1070
rect 11840 1050 11850 1070
rect 11810 1020 11850 1050
rect 11810 1000 11820 1020
rect 11840 1000 11850 1020
rect 11810 970 11850 1000
rect 11810 950 11820 970
rect 11840 950 11850 970
rect 11810 935 11850 950
rect 11865 1170 11905 1185
rect 11865 1150 11875 1170
rect 11895 1150 11905 1170
rect 11865 1120 11905 1150
rect 11865 1100 11875 1120
rect 11895 1100 11905 1120
rect 11865 1070 11905 1100
rect 11865 1050 11875 1070
rect 11895 1050 11905 1070
rect 11865 1020 11905 1050
rect 11865 1000 11875 1020
rect 11895 1000 11905 1020
rect 11865 970 11905 1000
rect 11865 950 11875 970
rect 11895 950 11905 970
rect 11865 935 11905 950
rect 11920 1170 11960 1185
rect 11920 1150 11930 1170
rect 11950 1150 11960 1170
rect 11920 1120 11960 1150
rect 11920 1100 11930 1120
rect 11950 1100 11960 1120
rect 11920 1070 11960 1100
rect 11920 1050 11930 1070
rect 11950 1050 11960 1070
rect 11920 1020 11960 1050
rect 11920 1000 11930 1020
rect 11950 1000 11960 1020
rect 11920 970 11960 1000
rect 11920 950 11930 970
rect 11950 950 11960 970
rect 11920 935 11960 950
rect 11975 1170 12015 1185
rect 11975 1150 11985 1170
rect 12005 1150 12015 1170
rect 11975 1120 12015 1150
rect 11975 1100 11985 1120
rect 12005 1100 12015 1120
rect 11975 1070 12015 1100
rect 11975 1050 11985 1070
rect 12005 1050 12015 1070
rect 11975 1020 12015 1050
rect 11975 1000 11985 1020
rect 12005 1000 12015 1020
rect 11975 970 12015 1000
rect 11975 950 11985 970
rect 12005 950 12015 970
rect 11975 935 12015 950
rect 12030 1170 12070 1185
rect 12030 1150 12040 1170
rect 12060 1150 12070 1170
rect 12030 1120 12070 1150
rect 12030 1100 12040 1120
rect 12060 1100 12070 1120
rect 12030 1070 12070 1100
rect 12030 1050 12040 1070
rect 12060 1050 12070 1070
rect 12030 1020 12070 1050
rect 12030 1000 12040 1020
rect 12060 1000 12070 1020
rect 12030 970 12070 1000
rect 12030 950 12040 970
rect 12060 950 12070 970
rect 12030 935 12070 950
rect 12085 1170 12125 1185
rect 12085 1150 12095 1170
rect 12115 1150 12125 1170
rect 12085 1120 12125 1150
rect 12085 1100 12095 1120
rect 12115 1100 12125 1120
rect 12085 1070 12125 1100
rect 12085 1050 12095 1070
rect 12115 1050 12125 1070
rect 12085 1020 12125 1050
rect 12085 1000 12095 1020
rect 12115 1000 12125 1020
rect 12085 970 12125 1000
rect 12085 950 12095 970
rect 12115 950 12125 970
rect 12085 935 12125 950
rect 12140 1170 12180 1185
rect 12140 1150 12150 1170
rect 12170 1150 12180 1170
rect 12140 1120 12180 1150
rect 12140 1100 12150 1120
rect 12170 1100 12180 1120
rect 12140 1070 12180 1100
rect 12140 1050 12150 1070
rect 12170 1050 12180 1070
rect 12140 1020 12180 1050
rect 12140 1000 12150 1020
rect 12170 1000 12180 1020
rect 12140 970 12180 1000
rect 12140 950 12150 970
rect 12170 950 12180 970
rect 12140 935 12180 950
rect 12195 1170 12235 1185
rect 12195 1150 12205 1170
rect 12225 1150 12235 1170
rect 12195 1120 12235 1150
rect 12195 1100 12205 1120
rect 12225 1100 12235 1120
rect 12195 1070 12235 1100
rect 12195 1050 12205 1070
rect 12225 1050 12235 1070
rect 12195 1020 12235 1050
rect 12195 1000 12205 1020
rect 12225 1000 12235 1020
rect 12195 970 12235 1000
rect 12195 950 12205 970
rect 12225 950 12235 970
rect 12195 935 12235 950
rect 12250 1170 12290 1185
rect 12250 1150 12260 1170
rect 12280 1150 12290 1170
rect 12250 1120 12290 1150
rect 12250 1100 12260 1120
rect 12280 1100 12290 1120
rect 12250 1070 12290 1100
rect 12250 1050 12260 1070
rect 12280 1050 12290 1070
rect 12250 1020 12290 1050
rect 12250 1000 12260 1020
rect 12280 1000 12290 1020
rect 12250 970 12290 1000
rect 12250 950 12260 970
rect 12280 950 12290 970
rect 12250 935 12290 950
rect 12305 1170 12345 1185
rect 12305 1150 12315 1170
rect 12335 1150 12345 1170
rect 12305 1120 12345 1150
rect 12305 1100 12315 1120
rect 12335 1100 12345 1120
rect 12305 1070 12345 1100
rect 12305 1050 12315 1070
rect 12335 1050 12345 1070
rect 12305 1020 12345 1050
rect 12305 1000 12315 1020
rect 12335 1000 12345 1020
rect 12305 970 12345 1000
rect 12305 950 12315 970
rect 12335 950 12345 970
rect 12305 935 12345 950
rect 12360 1170 12400 1185
rect 12360 1150 12370 1170
rect 12390 1150 12400 1170
rect 12360 1120 12400 1150
rect 12360 1100 12370 1120
rect 12390 1100 12400 1120
rect 12360 1070 12400 1100
rect 12360 1050 12370 1070
rect 12390 1050 12400 1070
rect 12360 1020 12400 1050
rect 12360 1000 12370 1020
rect 12390 1000 12400 1020
rect 12360 970 12400 1000
rect 12360 950 12370 970
rect 12390 950 12400 970
rect 12360 935 12400 950
rect 12415 1170 12455 1185
rect 12415 1150 12425 1170
rect 12445 1150 12455 1170
rect 12415 1120 12455 1150
rect 12415 1100 12425 1120
rect 12445 1100 12455 1120
rect 12415 1070 12455 1100
rect 12415 1050 12425 1070
rect 12445 1050 12455 1070
rect 12415 1020 12455 1050
rect 12415 1000 12425 1020
rect 12445 1000 12455 1020
rect 12415 970 12455 1000
rect 12415 950 12425 970
rect 12445 950 12455 970
rect 12415 935 12455 950
rect 12470 1170 12510 1185
rect 12470 1150 12480 1170
rect 12500 1150 12510 1170
rect 12470 1120 12510 1150
rect 12470 1100 12480 1120
rect 12500 1100 12510 1120
rect 12470 1070 12510 1100
rect 12470 1050 12480 1070
rect 12500 1050 12510 1070
rect 12470 1020 12510 1050
rect 12470 1000 12480 1020
rect 12500 1000 12510 1020
rect 12470 970 12510 1000
rect 12470 950 12480 970
rect 12500 950 12510 970
rect 12470 935 12510 950
rect 12525 1170 12565 1185
rect 12525 1150 12535 1170
rect 12555 1150 12565 1170
rect 12525 1120 12565 1150
rect 12525 1100 12535 1120
rect 12555 1100 12565 1120
rect 12525 1070 12565 1100
rect 12525 1050 12535 1070
rect 12555 1050 12565 1070
rect 12525 1020 12565 1050
rect 12525 1000 12535 1020
rect 12555 1000 12565 1020
rect 12525 970 12565 1000
rect 12525 950 12535 970
rect 12555 950 12565 970
rect 12525 935 12565 950
rect 12580 1170 12620 1185
rect 12580 1150 12590 1170
rect 12610 1150 12620 1170
rect 12580 1120 12620 1150
rect 12580 1100 12590 1120
rect 12610 1100 12620 1120
rect 12580 1070 12620 1100
rect 12580 1050 12590 1070
rect 12610 1050 12620 1070
rect 12580 1020 12620 1050
rect 12580 1000 12590 1020
rect 12610 1000 12620 1020
rect 12580 970 12620 1000
rect 12580 950 12590 970
rect 12610 950 12620 970
rect 13005 1170 13015 1190
rect 13035 1170 13045 1190
rect 13005 1140 13045 1170
rect 13005 1120 13015 1140
rect 13035 1120 13045 1140
rect 13005 1090 13045 1120
rect 13005 1070 13015 1090
rect 13035 1070 13045 1090
rect 13005 1040 13045 1070
rect 13005 1020 13015 1040
rect 13035 1020 13045 1040
rect 13005 990 13045 1020
rect 13005 970 13015 990
rect 13035 970 13045 990
rect 13005 955 13045 970
rect 13105 1640 13145 1655
rect 13105 1620 13115 1640
rect 13135 1620 13145 1640
rect 13105 1590 13145 1620
rect 13105 1570 13115 1590
rect 13135 1570 13145 1590
rect 13105 1540 13145 1570
rect 13105 1520 13115 1540
rect 13135 1520 13145 1540
rect 13105 1490 13145 1520
rect 13105 1470 13115 1490
rect 13135 1470 13145 1490
rect 13105 1440 13145 1470
rect 13105 1420 13115 1440
rect 13135 1420 13145 1440
rect 13105 1390 13145 1420
rect 13105 1370 13115 1390
rect 13135 1370 13145 1390
rect 13105 1340 13145 1370
rect 13105 1320 13115 1340
rect 13135 1320 13145 1340
rect 13105 1290 13145 1320
rect 13105 1270 13115 1290
rect 13135 1270 13145 1290
rect 13105 1240 13145 1270
rect 13105 1220 13115 1240
rect 13135 1220 13145 1240
rect 13105 1190 13145 1220
rect 13105 1170 13115 1190
rect 13135 1170 13145 1190
rect 13105 1140 13145 1170
rect 13105 1120 13115 1140
rect 13135 1120 13145 1140
rect 13105 1090 13145 1120
rect 13105 1070 13115 1090
rect 13135 1070 13145 1090
rect 13105 1040 13145 1070
rect 13105 1020 13115 1040
rect 13135 1020 13145 1040
rect 13105 990 13145 1020
rect 13105 970 13115 990
rect 13135 970 13145 990
rect 13105 955 13145 970
rect 13205 1640 13245 1655
rect 13205 1620 13215 1640
rect 13235 1620 13245 1640
rect 13205 1590 13245 1620
rect 13205 1570 13215 1590
rect 13235 1570 13245 1590
rect 13205 1540 13245 1570
rect 13205 1520 13215 1540
rect 13235 1520 13245 1540
rect 13205 1490 13245 1520
rect 13205 1470 13215 1490
rect 13235 1470 13245 1490
rect 13205 1440 13245 1470
rect 13205 1420 13215 1440
rect 13235 1420 13245 1440
rect 13205 1390 13245 1420
rect 13205 1370 13215 1390
rect 13235 1370 13245 1390
rect 13205 1340 13245 1370
rect 13205 1320 13215 1340
rect 13235 1320 13245 1340
rect 13205 1290 13245 1320
rect 13205 1270 13215 1290
rect 13235 1270 13245 1290
rect 13205 1240 13245 1270
rect 13205 1220 13215 1240
rect 13235 1220 13245 1240
rect 13205 1190 13245 1220
rect 13205 1170 13215 1190
rect 13235 1170 13245 1190
rect 13205 1140 13245 1170
rect 13205 1120 13215 1140
rect 13235 1120 13245 1140
rect 13205 1090 13245 1120
rect 13205 1070 13215 1090
rect 13235 1070 13245 1090
rect 13205 1040 13245 1070
rect 13205 1020 13215 1040
rect 13235 1020 13245 1040
rect 13205 990 13245 1020
rect 13205 970 13215 990
rect 13235 970 13245 990
rect 13205 955 13245 970
rect 13305 1640 13345 1655
rect 13305 1620 13315 1640
rect 13335 1620 13345 1640
rect 13305 1590 13345 1620
rect 13305 1570 13315 1590
rect 13335 1570 13345 1590
rect 13305 1540 13345 1570
rect 13305 1520 13315 1540
rect 13335 1520 13345 1540
rect 13305 1490 13345 1520
rect 13305 1470 13315 1490
rect 13335 1470 13345 1490
rect 13305 1440 13345 1470
rect 13305 1420 13315 1440
rect 13335 1420 13345 1440
rect 13305 1390 13345 1420
rect 13305 1370 13315 1390
rect 13335 1370 13345 1390
rect 13305 1340 13345 1370
rect 13305 1320 13315 1340
rect 13335 1320 13345 1340
rect 13305 1290 13345 1320
rect 13305 1270 13315 1290
rect 13335 1270 13345 1290
rect 13305 1240 13345 1270
rect 13305 1220 13315 1240
rect 13335 1220 13345 1240
rect 13305 1190 13345 1220
rect 13305 1170 13315 1190
rect 13335 1170 13345 1190
rect 13305 1140 13345 1170
rect 13305 1120 13315 1140
rect 13335 1120 13345 1140
rect 13305 1090 13345 1120
rect 13305 1070 13315 1090
rect 13335 1070 13345 1090
rect 13305 1040 13345 1070
rect 13305 1020 13315 1040
rect 13335 1020 13345 1040
rect 13305 990 13345 1020
rect 13305 970 13315 990
rect 13335 970 13345 990
rect 13305 955 13345 970
rect 13405 1640 13445 1655
rect 13405 1620 13415 1640
rect 13435 1620 13445 1640
rect 13405 1590 13445 1620
rect 13405 1570 13415 1590
rect 13435 1570 13445 1590
rect 13405 1540 13445 1570
rect 13405 1520 13415 1540
rect 13435 1520 13445 1540
rect 13405 1490 13445 1520
rect 13405 1470 13415 1490
rect 13435 1470 13445 1490
rect 13405 1440 13445 1470
rect 13405 1420 13415 1440
rect 13435 1420 13445 1440
rect 13405 1390 13445 1420
rect 13405 1370 13415 1390
rect 13435 1370 13445 1390
rect 13405 1340 13445 1370
rect 13405 1320 13415 1340
rect 13435 1320 13445 1340
rect 13405 1290 13445 1320
rect 13405 1270 13415 1290
rect 13435 1270 13445 1290
rect 13405 1240 13445 1270
rect 13405 1220 13415 1240
rect 13435 1220 13445 1240
rect 13405 1190 13445 1220
rect 13405 1170 13415 1190
rect 13435 1170 13445 1190
rect 13405 1140 13445 1170
rect 13405 1120 13415 1140
rect 13435 1120 13445 1140
rect 13405 1090 13445 1120
rect 13405 1070 13415 1090
rect 13435 1070 13445 1090
rect 13405 1040 13445 1070
rect 13405 1020 13415 1040
rect 13435 1020 13445 1040
rect 13405 990 13445 1020
rect 13405 970 13415 990
rect 13435 970 13445 990
rect 13405 955 13445 970
rect 13505 1640 13545 1655
rect 13505 1620 13515 1640
rect 13535 1620 13545 1640
rect 13505 1590 13545 1620
rect 13505 1570 13515 1590
rect 13535 1570 13545 1590
rect 13505 1540 13545 1570
rect 13505 1520 13515 1540
rect 13535 1520 13545 1540
rect 13505 1490 13545 1520
rect 13505 1470 13515 1490
rect 13535 1470 13545 1490
rect 13505 1440 13545 1470
rect 13505 1420 13515 1440
rect 13535 1420 13545 1440
rect 13505 1390 13545 1420
rect 13505 1370 13515 1390
rect 13535 1370 13545 1390
rect 13505 1340 13545 1370
rect 13505 1320 13515 1340
rect 13535 1320 13545 1340
rect 13505 1290 13545 1320
rect 13505 1270 13515 1290
rect 13535 1270 13545 1290
rect 13505 1240 13545 1270
rect 13505 1220 13515 1240
rect 13535 1220 13545 1240
rect 13505 1190 13545 1220
rect 13505 1170 13515 1190
rect 13535 1170 13545 1190
rect 13505 1140 13545 1170
rect 13505 1120 13515 1140
rect 13535 1120 13545 1140
rect 13505 1090 13545 1120
rect 13505 1070 13515 1090
rect 13535 1070 13545 1090
rect 13505 1040 13545 1070
rect 13505 1020 13515 1040
rect 13535 1020 13545 1040
rect 13505 990 13545 1020
rect 13505 970 13515 990
rect 13535 970 13545 990
rect 13505 955 13545 970
rect 13605 1640 13645 1655
rect 13605 1620 13615 1640
rect 13635 1620 13645 1640
rect 13605 1590 13645 1620
rect 26030 1650 26070 1665
rect 26030 1630 26040 1650
rect 26060 1630 26070 1650
rect 13605 1570 13615 1590
rect 13635 1570 13645 1590
rect 13605 1540 13645 1570
rect 13605 1520 13615 1540
rect 13635 1520 13645 1540
rect 13605 1490 13645 1520
rect 13605 1470 13615 1490
rect 13635 1470 13645 1490
rect 13605 1440 13645 1470
rect 13605 1420 13615 1440
rect 13635 1420 13645 1440
rect 13605 1390 13645 1420
rect 13605 1370 13615 1390
rect 13635 1370 13645 1390
rect 13605 1340 13645 1370
rect 13605 1320 13615 1340
rect 13635 1320 13645 1340
rect 13605 1290 13645 1320
rect 13605 1270 13615 1290
rect 13635 1270 13645 1290
rect 13605 1240 13645 1270
rect 13605 1220 13615 1240
rect 13635 1220 13645 1240
rect 13605 1190 13645 1220
rect 13605 1170 13615 1190
rect 13635 1170 13645 1190
rect 13605 1140 13645 1170
rect 13605 1120 13615 1140
rect 13635 1120 13645 1140
rect 13605 1090 13645 1120
rect 13605 1070 13615 1090
rect 13635 1070 13645 1090
rect 13605 1040 13645 1070
rect 13605 1020 13615 1040
rect 13635 1020 13645 1040
rect 13605 990 13645 1020
rect 13605 970 13615 990
rect 13635 970 13645 990
rect 13605 955 13645 970
rect 12580 935 12620 950
rect 26030 1600 26070 1630
rect 26030 1580 26040 1600
rect 26060 1580 26070 1600
rect 26030 1550 26070 1580
rect 26030 1530 26040 1550
rect 26060 1530 26070 1550
rect 26030 1515 26070 1530
rect 26085 1650 26125 1665
rect 26085 1630 26095 1650
rect 26115 1630 26125 1650
rect 26085 1600 26125 1630
rect 26085 1580 26095 1600
rect 26115 1580 26125 1600
rect 26085 1550 26125 1580
rect 26085 1530 26095 1550
rect 26115 1530 26125 1550
rect 26085 1515 26125 1530
rect 26140 1650 26180 1665
rect 26140 1630 26150 1650
rect 26170 1630 26180 1650
rect 26140 1600 26180 1630
rect 26140 1580 26150 1600
rect 26170 1580 26180 1600
rect 26140 1550 26180 1580
rect 26140 1530 26150 1550
rect 26170 1530 26180 1550
rect 26140 1515 26180 1530
rect 26195 1650 26235 1665
rect 26195 1630 26205 1650
rect 26225 1630 26235 1650
rect 26195 1600 26235 1630
rect 26195 1580 26205 1600
rect 26225 1580 26235 1600
rect 26195 1550 26235 1580
rect 26195 1530 26205 1550
rect 26225 1530 26235 1550
rect 26195 1515 26235 1530
rect 26250 1650 26290 1665
rect 26250 1630 26260 1650
rect 26280 1630 26290 1650
rect 26250 1600 26290 1630
rect 26250 1580 26260 1600
rect 26280 1580 26290 1600
rect 26250 1550 26290 1580
rect 26250 1530 26260 1550
rect 26280 1530 26290 1550
rect 26250 1515 26290 1530
rect 26305 1650 26345 1665
rect 26305 1630 26315 1650
rect 26335 1630 26345 1650
rect 26305 1600 26345 1630
rect 26305 1580 26315 1600
rect 26335 1580 26345 1600
rect 26305 1550 26345 1580
rect 26305 1530 26315 1550
rect 26335 1530 26345 1550
rect 26305 1515 26345 1530
rect 26360 1650 26400 1665
rect 26360 1630 26370 1650
rect 26390 1630 26400 1650
rect 26360 1600 26400 1630
rect 26360 1580 26370 1600
rect 26390 1580 26400 1600
rect 26360 1550 26400 1580
rect 26360 1530 26370 1550
rect 26390 1530 26400 1550
rect 26360 1515 26400 1530
rect 26415 1650 26455 1665
rect 26415 1630 26425 1650
rect 26445 1630 26455 1650
rect 26415 1600 26455 1630
rect 26415 1580 26425 1600
rect 26445 1580 26455 1600
rect 26415 1550 26455 1580
rect 26415 1530 26425 1550
rect 26445 1530 26455 1550
rect 26415 1515 26455 1530
rect 26470 1650 26510 1665
rect 26470 1630 26480 1650
rect 26500 1630 26510 1650
rect 26470 1600 26510 1630
rect 26470 1580 26480 1600
rect 26500 1580 26510 1600
rect 26470 1550 26510 1580
rect 26470 1530 26480 1550
rect 26500 1530 26510 1550
rect 26470 1515 26510 1530
rect 26525 1650 26565 1665
rect 26525 1630 26535 1650
rect 26555 1630 26565 1650
rect 26525 1600 26565 1630
rect 26525 1580 26535 1600
rect 26555 1580 26565 1600
rect 26525 1550 26565 1580
rect 26525 1530 26535 1550
rect 26555 1530 26565 1550
rect 26525 1515 26565 1530
rect 26580 1650 26620 1665
rect 26580 1630 26590 1650
rect 26610 1630 26620 1650
rect 26580 1600 26620 1630
rect 26580 1580 26590 1600
rect 26610 1580 26620 1600
rect 26580 1550 26620 1580
rect 26580 1530 26590 1550
rect 26610 1530 26620 1550
rect 26580 1515 26620 1530
rect 26635 1650 26675 1665
rect 26635 1630 26645 1650
rect 26665 1630 26675 1650
rect 26635 1600 26675 1630
rect 26635 1580 26645 1600
rect 26665 1580 26675 1600
rect 26635 1550 26675 1580
rect 26635 1530 26645 1550
rect 26665 1530 26675 1550
rect 26635 1515 26675 1530
rect 26690 1650 26730 1665
rect 26770 1650 26810 1665
rect 26690 1630 26700 1650
rect 26720 1630 26730 1650
rect 26770 1630 26780 1650
rect 26800 1630 26810 1650
rect 26690 1600 26730 1630
rect 26770 1600 26810 1630
rect 26690 1580 26700 1600
rect 26720 1580 26730 1600
rect 26770 1580 26780 1600
rect 26800 1580 26810 1600
rect 26690 1550 26730 1580
rect 26770 1550 26810 1580
rect 26690 1530 26700 1550
rect 26720 1530 26730 1550
rect 26770 1530 26780 1550
rect 26800 1530 26810 1550
rect 26690 1515 26730 1530
rect 26770 1515 26810 1530
rect 26825 1650 26865 1665
rect 26825 1630 26835 1650
rect 26855 1630 26865 1650
rect 26825 1600 26865 1630
rect 26825 1580 26835 1600
rect 26855 1580 26865 1600
rect 26825 1550 26865 1580
rect 26825 1530 26835 1550
rect 26855 1530 26865 1550
rect 26825 1515 26865 1530
rect 26880 1650 26920 1665
rect 26880 1630 26890 1650
rect 26910 1630 26920 1650
rect 26880 1600 26920 1630
rect 26880 1580 26890 1600
rect 26910 1580 26920 1600
rect 26880 1550 26920 1580
rect 26880 1530 26890 1550
rect 26910 1530 26920 1550
rect 26880 1515 26920 1530
rect 26935 1650 26975 1665
rect 26935 1630 26945 1650
rect 26965 1630 26975 1650
rect 26935 1600 26975 1630
rect 26935 1580 26945 1600
rect 26965 1580 26975 1600
rect 26935 1550 26975 1580
rect 26935 1530 26945 1550
rect 26965 1530 26975 1550
rect 26935 1515 26975 1530
rect 26990 1650 27030 1665
rect 27070 1650 27110 1665
rect 26990 1630 27000 1650
rect 27020 1630 27030 1650
rect 27070 1630 27080 1650
rect 27100 1630 27110 1650
rect 26990 1600 27030 1630
rect 27070 1600 27110 1630
rect 26990 1580 27000 1600
rect 27020 1580 27030 1600
rect 27070 1580 27080 1600
rect 27100 1580 27110 1600
rect 26990 1550 27030 1580
rect 27070 1550 27110 1580
rect 26990 1530 27000 1550
rect 27020 1530 27030 1550
rect 27070 1530 27080 1550
rect 27100 1530 27110 1550
rect 26990 1515 27030 1530
rect 27070 1515 27110 1530
rect 27125 1650 27165 1665
rect 27125 1630 27135 1650
rect 27155 1630 27165 1650
rect 27125 1600 27165 1630
rect 27125 1580 27135 1600
rect 27155 1580 27165 1600
rect 27125 1550 27165 1580
rect 27125 1530 27135 1550
rect 27155 1530 27165 1550
rect 27125 1515 27165 1530
rect 27180 1650 27220 1665
rect 27180 1630 27190 1650
rect 27210 1630 27220 1650
rect 27180 1600 27220 1630
rect 27180 1580 27190 1600
rect 27210 1580 27220 1600
rect 27180 1550 27220 1580
rect 27180 1530 27190 1550
rect 27210 1530 27220 1550
rect 27180 1515 27220 1530
rect 27235 1650 27275 1665
rect 27235 1630 27245 1650
rect 27265 1630 27275 1650
rect 27235 1600 27275 1630
rect 27235 1580 27245 1600
rect 27265 1580 27275 1600
rect 27235 1550 27275 1580
rect 27235 1530 27245 1550
rect 27265 1530 27275 1550
rect 27235 1515 27275 1530
rect 27290 1650 27330 1665
rect 27290 1630 27300 1650
rect 27320 1630 27330 1650
rect 27290 1600 27330 1630
rect 27290 1580 27300 1600
rect 27320 1580 27330 1600
rect 27290 1550 27330 1580
rect 27290 1530 27300 1550
rect 27320 1530 27330 1550
rect 27290 1515 27330 1530
rect 27345 1650 27385 1665
rect 27345 1630 27355 1650
rect 27375 1630 27385 1650
rect 27345 1600 27385 1630
rect 27345 1580 27355 1600
rect 27375 1580 27385 1600
rect 27345 1550 27385 1580
rect 27345 1530 27355 1550
rect 27375 1530 27385 1550
rect 27345 1515 27385 1530
rect 27400 1650 27440 1665
rect 27400 1630 27410 1650
rect 27430 1630 27440 1650
rect 27400 1600 27440 1630
rect 27400 1580 27410 1600
rect 27430 1580 27440 1600
rect 27400 1550 27440 1580
rect 27400 1530 27410 1550
rect 27430 1530 27440 1550
rect 27400 1515 27440 1530
rect 27455 1650 27495 1665
rect 27455 1630 27465 1650
rect 27485 1630 27495 1650
rect 27455 1600 27495 1630
rect 27455 1580 27465 1600
rect 27485 1580 27495 1600
rect 27455 1550 27495 1580
rect 27455 1530 27465 1550
rect 27485 1530 27495 1550
rect 27455 1515 27495 1530
rect 27510 1650 27550 1665
rect 27510 1630 27520 1650
rect 27540 1630 27550 1650
rect 27510 1600 27550 1630
rect 27510 1580 27520 1600
rect 27540 1580 27550 1600
rect 27510 1550 27550 1580
rect 27510 1530 27520 1550
rect 27540 1530 27550 1550
rect 27510 1515 27550 1530
rect 27565 1650 27605 1665
rect 27565 1630 27575 1650
rect 27595 1630 27605 1650
rect 27565 1600 27605 1630
rect 27565 1580 27575 1600
rect 27595 1580 27605 1600
rect 27565 1550 27605 1580
rect 27565 1530 27575 1550
rect 27595 1530 27605 1550
rect 27565 1515 27605 1530
rect 27620 1650 27660 1665
rect 27620 1630 27630 1650
rect 27650 1630 27660 1650
rect 27620 1600 27660 1630
rect 27620 1580 27630 1600
rect 27650 1580 27660 1600
rect 27620 1550 27660 1580
rect 27620 1530 27630 1550
rect 27650 1530 27660 1550
rect 27620 1515 27660 1530
rect 27675 1650 27715 1665
rect 27675 1630 27685 1650
rect 27705 1630 27715 1650
rect 27675 1600 27715 1630
rect 27675 1580 27685 1600
rect 27705 1580 27715 1600
rect 27675 1550 27715 1580
rect 27675 1530 27685 1550
rect 27705 1530 27715 1550
rect 27675 1515 27715 1530
rect 27730 1650 27770 1665
rect 27730 1630 27740 1650
rect 27760 1630 27770 1650
rect 27730 1600 27770 1630
rect 27730 1580 27740 1600
rect 27760 1580 27770 1600
rect 27730 1550 27770 1580
rect 27730 1530 27740 1550
rect 27760 1530 27770 1550
rect 27730 1515 27770 1530
rect 27895 1505 27935 1520
rect 27895 1485 27905 1505
rect 27925 1485 27935 1505
rect 27895 1455 27935 1485
rect 27895 1435 27905 1455
rect 27925 1435 27935 1455
rect 27895 1405 27935 1435
rect 27895 1385 27905 1405
rect 27925 1385 27935 1405
rect 27895 1370 27935 1385
rect 27950 1505 27990 1520
rect 27950 1485 27960 1505
rect 27980 1485 27990 1505
rect 27950 1455 27990 1485
rect 27950 1435 27960 1455
rect 27980 1435 27990 1455
rect 27950 1405 27990 1435
rect 27950 1385 27960 1405
rect 27980 1385 27990 1405
rect 27950 1370 27990 1385
rect 28005 1505 28045 1520
rect 28005 1485 28015 1505
rect 28035 1485 28045 1505
rect 28005 1455 28045 1485
rect 28005 1435 28015 1455
rect 28035 1435 28045 1455
rect 28005 1405 28045 1435
rect 28005 1385 28015 1405
rect 28035 1385 28045 1405
rect 28005 1370 28045 1385
rect 28060 1505 28100 1520
rect 28060 1485 28070 1505
rect 28090 1485 28100 1505
rect 28060 1455 28100 1485
rect 28060 1435 28070 1455
rect 28090 1435 28100 1455
rect 28060 1405 28100 1435
rect 28060 1385 28070 1405
rect 28090 1385 28100 1405
rect 28060 1370 28100 1385
rect 28115 1505 28155 1520
rect 28195 1505 28235 1520
rect 28115 1485 28125 1505
rect 28145 1485 28155 1505
rect 28195 1485 28205 1505
rect 28225 1485 28235 1505
rect 28115 1455 28155 1485
rect 28195 1455 28235 1485
rect 28115 1435 28125 1455
rect 28145 1435 28155 1455
rect 28195 1435 28205 1455
rect 28225 1435 28235 1455
rect 28115 1405 28155 1435
rect 28195 1405 28235 1435
rect 28115 1385 28125 1405
rect 28145 1385 28155 1405
rect 28195 1385 28205 1405
rect 28225 1385 28235 1405
rect 28115 1370 28155 1385
rect 28195 1370 28235 1385
rect 28250 1505 28290 1520
rect 28250 1485 28260 1505
rect 28280 1485 28290 1505
rect 28250 1455 28290 1485
rect 28250 1435 28260 1455
rect 28280 1435 28290 1455
rect 28250 1405 28290 1435
rect 28250 1385 28260 1405
rect 28280 1385 28290 1405
rect 28250 1370 28290 1385
rect 28305 1505 28345 1520
rect 28305 1485 28315 1505
rect 28335 1485 28345 1505
rect 28305 1455 28345 1485
rect 28305 1435 28315 1455
rect 28335 1435 28345 1455
rect 28305 1405 28345 1435
rect 28305 1385 28315 1405
rect 28335 1385 28345 1405
rect 28305 1370 28345 1385
rect 28360 1505 28400 1520
rect 28360 1485 28370 1505
rect 28390 1485 28400 1505
rect 28360 1455 28400 1485
rect 28360 1435 28370 1455
rect 28390 1435 28400 1455
rect 28360 1405 28400 1435
rect 28360 1385 28370 1405
rect 28390 1385 28400 1405
rect 28360 1370 28400 1385
rect 28415 1505 28455 1520
rect 28415 1485 28425 1505
rect 28445 1485 28455 1505
rect 28415 1455 28455 1485
rect 28415 1435 28425 1455
rect 28445 1435 28455 1455
rect 28415 1405 28455 1435
rect 28415 1385 28425 1405
rect 28445 1385 28455 1405
rect 28415 1370 28455 1385
rect 26205 1210 26245 1225
rect 26205 1190 26215 1210
rect 26235 1190 26245 1210
rect 26205 1160 26245 1190
rect 26205 1140 26215 1160
rect 26235 1140 26245 1160
rect 26205 1110 26245 1140
rect 26205 1090 26215 1110
rect 26235 1090 26245 1110
rect 26205 1060 26245 1090
rect 26205 1040 26215 1060
rect 26235 1040 26245 1060
rect 26205 1010 26245 1040
rect 26205 990 26215 1010
rect 26235 990 26245 1010
rect 26205 975 26245 990
rect 26260 1210 26300 1225
rect 26260 1190 26270 1210
rect 26290 1190 26300 1210
rect 26260 1160 26300 1190
rect 26260 1140 26270 1160
rect 26290 1140 26300 1160
rect 26260 1110 26300 1140
rect 26260 1090 26270 1110
rect 26290 1090 26300 1110
rect 26260 1060 26300 1090
rect 26260 1040 26270 1060
rect 26290 1040 26300 1060
rect 26260 1010 26300 1040
rect 26260 990 26270 1010
rect 26290 990 26300 1010
rect 26260 975 26300 990
rect 26315 1210 26355 1225
rect 26315 1190 26325 1210
rect 26345 1190 26355 1210
rect 26315 1160 26355 1190
rect 26315 1140 26325 1160
rect 26345 1140 26355 1160
rect 26315 1110 26355 1140
rect 26315 1090 26325 1110
rect 26345 1090 26355 1110
rect 26315 1060 26355 1090
rect 26315 1040 26325 1060
rect 26345 1040 26355 1060
rect 26315 1010 26355 1040
rect 26315 990 26325 1010
rect 26345 990 26355 1010
rect 26315 975 26355 990
rect 26370 1210 26410 1225
rect 26370 1190 26380 1210
rect 26400 1190 26410 1210
rect 26370 1160 26410 1190
rect 26370 1140 26380 1160
rect 26400 1140 26410 1160
rect 26370 1110 26410 1140
rect 26370 1090 26380 1110
rect 26400 1090 26410 1110
rect 26370 1060 26410 1090
rect 26370 1040 26380 1060
rect 26400 1040 26410 1060
rect 26370 1010 26410 1040
rect 26370 990 26380 1010
rect 26400 990 26410 1010
rect 26370 975 26410 990
rect 26425 1210 26465 1225
rect 26425 1190 26435 1210
rect 26455 1190 26465 1210
rect 26425 1160 26465 1190
rect 26425 1140 26435 1160
rect 26455 1140 26465 1160
rect 26425 1110 26465 1140
rect 26425 1090 26435 1110
rect 26455 1090 26465 1110
rect 26425 1060 26465 1090
rect 26425 1040 26435 1060
rect 26455 1040 26465 1060
rect 26425 1010 26465 1040
rect 26425 990 26435 1010
rect 26455 990 26465 1010
rect 26425 975 26465 990
rect 26480 1210 26520 1225
rect 26480 1190 26490 1210
rect 26510 1190 26520 1210
rect 26480 1160 26520 1190
rect 26480 1140 26490 1160
rect 26510 1140 26520 1160
rect 26480 1110 26520 1140
rect 26480 1090 26490 1110
rect 26510 1090 26520 1110
rect 26480 1060 26520 1090
rect 26480 1040 26490 1060
rect 26510 1040 26520 1060
rect 26480 1010 26520 1040
rect 26480 990 26490 1010
rect 26510 990 26520 1010
rect 26480 975 26520 990
rect 26535 1210 26575 1225
rect 26535 1190 26545 1210
rect 26565 1190 26575 1210
rect 26535 1160 26575 1190
rect 26535 1140 26545 1160
rect 26565 1140 26575 1160
rect 26535 1110 26575 1140
rect 26535 1090 26545 1110
rect 26565 1090 26575 1110
rect 26535 1060 26575 1090
rect 26535 1040 26545 1060
rect 26565 1040 26575 1060
rect 26535 1010 26575 1040
rect 26535 990 26545 1010
rect 26565 990 26575 1010
rect 26535 975 26575 990
rect 26590 1210 26630 1225
rect 26590 1190 26600 1210
rect 26620 1190 26630 1210
rect 26590 1160 26630 1190
rect 26590 1140 26600 1160
rect 26620 1140 26630 1160
rect 26590 1110 26630 1140
rect 26590 1090 26600 1110
rect 26620 1090 26630 1110
rect 26590 1060 26630 1090
rect 26590 1040 26600 1060
rect 26620 1040 26630 1060
rect 26590 1010 26630 1040
rect 26590 990 26600 1010
rect 26620 990 26630 1010
rect 26590 975 26630 990
rect 26645 1210 26685 1225
rect 26645 1190 26655 1210
rect 26675 1190 26685 1210
rect 26645 1160 26685 1190
rect 26645 1140 26655 1160
rect 26675 1140 26685 1160
rect 26645 1110 26685 1140
rect 26645 1090 26655 1110
rect 26675 1090 26685 1110
rect 26645 1060 26685 1090
rect 26645 1040 26655 1060
rect 26675 1040 26685 1060
rect 26645 1010 26685 1040
rect 26645 990 26655 1010
rect 26675 990 26685 1010
rect 26645 975 26685 990
rect 26700 1210 26740 1225
rect 26700 1190 26710 1210
rect 26730 1190 26740 1210
rect 26700 1160 26740 1190
rect 26700 1140 26710 1160
rect 26730 1140 26740 1160
rect 26700 1110 26740 1140
rect 26700 1090 26710 1110
rect 26730 1090 26740 1110
rect 26700 1060 26740 1090
rect 26700 1040 26710 1060
rect 26730 1040 26740 1060
rect 26700 1010 26740 1040
rect 26700 990 26710 1010
rect 26730 990 26740 1010
rect 26700 975 26740 990
rect 26755 1210 26795 1225
rect 26755 1190 26765 1210
rect 26785 1190 26795 1210
rect 26755 1160 26795 1190
rect 26755 1140 26765 1160
rect 26785 1140 26795 1160
rect 26755 1110 26795 1140
rect 26755 1090 26765 1110
rect 26785 1090 26795 1110
rect 26755 1060 26795 1090
rect 26755 1040 26765 1060
rect 26785 1040 26795 1060
rect 26755 1010 26795 1040
rect 26755 990 26765 1010
rect 26785 990 26795 1010
rect 26755 975 26795 990
rect 26810 1210 26850 1225
rect 26810 1190 26820 1210
rect 26840 1190 26850 1210
rect 26810 1160 26850 1190
rect 26810 1140 26820 1160
rect 26840 1140 26850 1160
rect 26810 1110 26850 1140
rect 26810 1090 26820 1110
rect 26840 1090 26850 1110
rect 26810 1060 26850 1090
rect 26810 1040 26820 1060
rect 26840 1040 26850 1060
rect 26810 1010 26850 1040
rect 26810 990 26820 1010
rect 26840 990 26850 1010
rect 26810 975 26850 990
rect 26865 1210 26905 1225
rect 26865 1190 26875 1210
rect 26895 1190 26905 1210
rect 26865 1160 26905 1190
rect 26865 1140 26875 1160
rect 26895 1140 26905 1160
rect 26865 1110 26905 1140
rect 26865 1090 26875 1110
rect 26895 1090 26905 1110
rect 26865 1060 26905 1090
rect 26865 1040 26875 1060
rect 26895 1040 26905 1060
rect 26865 1010 26905 1040
rect 26865 990 26875 1010
rect 26895 990 26905 1010
rect 26865 975 26905 990
rect 26920 1210 26960 1225
rect 26920 1190 26930 1210
rect 26950 1190 26960 1210
rect 26920 1160 26960 1190
rect 26920 1140 26930 1160
rect 26950 1140 26960 1160
rect 26920 1110 26960 1140
rect 26920 1090 26930 1110
rect 26950 1090 26960 1110
rect 26920 1060 26960 1090
rect 26920 1040 26930 1060
rect 26950 1040 26960 1060
rect 26920 1010 26960 1040
rect 26920 990 26930 1010
rect 26950 990 26960 1010
rect 26920 975 26960 990
rect 26975 1210 27015 1225
rect 26975 1190 26985 1210
rect 27005 1190 27015 1210
rect 26975 1160 27015 1190
rect 26975 1140 26985 1160
rect 27005 1140 27015 1160
rect 26975 1110 27015 1140
rect 26975 1090 26985 1110
rect 27005 1090 27015 1110
rect 26975 1060 27015 1090
rect 26975 1040 26985 1060
rect 27005 1040 27015 1060
rect 26975 1010 27015 1040
rect 26975 990 26985 1010
rect 27005 990 27015 1010
rect 26975 975 27015 990
rect 27030 1210 27070 1225
rect 27030 1190 27040 1210
rect 27060 1190 27070 1210
rect 27030 1160 27070 1190
rect 27030 1140 27040 1160
rect 27060 1140 27070 1160
rect 27030 1110 27070 1140
rect 27030 1090 27040 1110
rect 27060 1090 27070 1110
rect 27030 1060 27070 1090
rect 27030 1040 27040 1060
rect 27060 1040 27070 1060
rect 27030 1010 27070 1040
rect 27030 990 27040 1010
rect 27060 990 27070 1010
rect 27030 975 27070 990
rect 27085 1210 27125 1225
rect 27085 1190 27095 1210
rect 27115 1190 27125 1210
rect 27085 1160 27125 1190
rect 27085 1140 27095 1160
rect 27115 1140 27125 1160
rect 27085 1110 27125 1140
rect 27085 1090 27095 1110
rect 27115 1090 27125 1110
rect 27085 1060 27125 1090
rect 27085 1040 27095 1060
rect 27115 1040 27125 1060
rect 27085 1010 27125 1040
rect 27085 990 27095 1010
rect 27115 990 27125 1010
rect 27085 975 27125 990
rect 27140 1210 27180 1225
rect 27140 1190 27150 1210
rect 27170 1190 27180 1210
rect 27140 1160 27180 1190
rect 27140 1140 27150 1160
rect 27170 1140 27180 1160
rect 27140 1110 27180 1140
rect 27140 1090 27150 1110
rect 27170 1090 27180 1110
rect 27140 1060 27180 1090
rect 27140 1040 27150 1060
rect 27170 1040 27180 1060
rect 27140 1010 27180 1040
rect 27140 990 27150 1010
rect 27170 990 27180 1010
rect 27140 975 27180 990
rect 27195 1210 27235 1225
rect 27195 1190 27205 1210
rect 27225 1190 27235 1210
rect 27195 1160 27235 1190
rect 27195 1140 27205 1160
rect 27225 1140 27235 1160
rect 27195 1110 27235 1140
rect 27195 1090 27205 1110
rect 27225 1090 27235 1110
rect 27195 1060 27235 1090
rect 27195 1040 27205 1060
rect 27225 1040 27235 1060
rect 27195 1010 27235 1040
rect 27195 990 27205 1010
rect 27225 990 27235 1010
rect 27195 975 27235 990
rect 27250 1210 27290 1225
rect 27250 1190 27260 1210
rect 27280 1190 27290 1210
rect 27250 1160 27290 1190
rect 27250 1140 27260 1160
rect 27280 1140 27290 1160
rect 27250 1110 27290 1140
rect 27250 1090 27260 1110
rect 27280 1090 27290 1110
rect 27250 1060 27290 1090
rect 27250 1040 27260 1060
rect 27280 1040 27290 1060
rect 27250 1010 27290 1040
rect 27250 990 27260 1010
rect 27280 990 27290 1010
rect 27250 975 27290 990
rect 27305 1210 27345 1225
rect 27305 1190 27315 1210
rect 27335 1190 27345 1210
rect 27305 1160 27345 1190
rect 27305 1140 27315 1160
rect 27335 1140 27345 1160
rect 27305 1110 27345 1140
rect 27305 1090 27315 1110
rect 27335 1090 27345 1110
rect 27305 1060 27345 1090
rect 27305 1040 27315 1060
rect 27335 1040 27345 1060
rect 27305 1010 27345 1040
rect 27305 990 27315 1010
rect 27335 990 27345 1010
rect 27305 975 27345 990
rect 27360 1210 27400 1225
rect 27360 1190 27370 1210
rect 27390 1190 27400 1210
rect 27360 1160 27400 1190
rect 27360 1140 27370 1160
rect 27390 1140 27400 1160
rect 27360 1110 27400 1140
rect 27360 1090 27370 1110
rect 27390 1090 27400 1110
rect 27360 1060 27400 1090
rect 27360 1040 27370 1060
rect 27390 1040 27400 1060
rect 27360 1010 27400 1040
rect 27360 990 27370 1010
rect 27390 990 27400 1010
rect 27360 975 27400 990
rect 27415 1210 27455 1225
rect 27415 1190 27425 1210
rect 27445 1190 27455 1210
rect 27415 1160 27455 1190
rect 27415 1140 27425 1160
rect 27445 1140 27455 1160
rect 27415 1110 27455 1140
rect 27415 1090 27425 1110
rect 27445 1090 27455 1110
rect 27415 1060 27455 1090
rect 27415 1040 27425 1060
rect 27445 1040 27455 1060
rect 27415 1010 27455 1040
rect 27415 990 27425 1010
rect 27445 990 27455 1010
rect 27415 975 27455 990
rect 27470 1210 27510 1225
rect 27470 1190 27480 1210
rect 27500 1190 27510 1210
rect 27470 1160 27510 1190
rect 27470 1140 27480 1160
rect 27500 1140 27510 1160
rect 27470 1110 27510 1140
rect 27470 1090 27480 1110
rect 27500 1090 27510 1110
rect 27470 1060 27510 1090
rect 27470 1040 27480 1060
rect 27500 1040 27510 1060
rect 27470 1010 27510 1040
rect 27470 990 27480 1010
rect 27500 990 27510 1010
rect 27470 975 27510 990
rect 27525 1210 27565 1225
rect 27525 1190 27535 1210
rect 27555 1190 27565 1210
rect 27525 1160 27565 1190
rect 27525 1140 27535 1160
rect 27555 1140 27565 1160
rect 27525 1110 27565 1140
rect 27525 1090 27535 1110
rect 27555 1090 27565 1110
rect 27525 1060 27565 1090
rect 27525 1040 27535 1060
rect 27555 1040 27565 1060
rect 27525 1010 27565 1040
rect 27525 990 27535 1010
rect 27555 990 27565 1010
rect 27525 975 27565 990
rect 27580 1210 27620 1225
rect 27580 1190 27590 1210
rect 27610 1190 27620 1210
rect 27580 1160 27620 1190
rect 27580 1140 27590 1160
rect 27610 1140 27620 1160
rect 27580 1110 27620 1140
rect 27580 1090 27590 1110
rect 27610 1090 27620 1110
rect 27580 1060 27620 1090
rect 27580 1040 27590 1060
rect 27610 1040 27620 1060
rect 27580 1010 27620 1040
rect 28045 1165 28085 1180
rect 28045 1145 28055 1165
rect 28075 1145 28085 1165
rect 28045 1115 28085 1145
rect 28045 1095 28055 1115
rect 28075 1095 28085 1115
rect 28045 1065 28085 1095
rect 28045 1045 28055 1065
rect 28075 1045 28085 1065
rect 28045 1030 28085 1045
rect 28100 1165 28140 1180
rect 28100 1145 28110 1165
rect 28130 1145 28140 1165
rect 28100 1115 28140 1145
rect 28100 1095 28110 1115
rect 28130 1095 28140 1115
rect 28100 1065 28140 1095
rect 28100 1045 28110 1065
rect 28130 1045 28140 1065
rect 28100 1030 28140 1045
rect 28155 1165 28195 1180
rect 28155 1145 28165 1165
rect 28185 1145 28195 1165
rect 28155 1115 28195 1145
rect 28155 1095 28165 1115
rect 28185 1095 28195 1115
rect 28155 1065 28195 1095
rect 28155 1045 28165 1065
rect 28185 1045 28195 1065
rect 28155 1030 28195 1045
rect 28210 1165 28250 1180
rect 28210 1145 28220 1165
rect 28240 1145 28250 1165
rect 28210 1115 28250 1145
rect 28210 1095 28220 1115
rect 28240 1095 28250 1115
rect 28210 1065 28250 1095
rect 28210 1045 28220 1065
rect 28240 1045 28250 1065
rect 28210 1030 28250 1045
rect 28265 1165 28305 1180
rect 28265 1145 28275 1165
rect 28295 1145 28305 1165
rect 28265 1115 28305 1145
rect 28265 1095 28275 1115
rect 28295 1095 28305 1115
rect 28265 1065 28305 1095
rect 28265 1045 28275 1065
rect 28295 1045 28305 1065
rect 28265 1030 28305 1045
rect 27580 990 27590 1010
rect 27610 990 27620 1010
rect 27580 975 27620 990
rect 2995 865 3035 880
rect 2995 845 3005 865
rect 3025 845 3035 865
rect 2995 815 3035 845
rect 2995 795 3005 815
rect 3025 795 3035 815
rect 2995 780 3035 795
rect 3085 865 3125 880
rect 3085 845 3095 865
rect 3115 845 3125 865
rect 3085 815 3125 845
rect 3085 795 3095 815
rect 3115 795 3125 815
rect 3085 780 3125 795
rect 3175 865 3215 880
rect 3175 845 3185 865
rect 3205 845 3215 865
rect 3175 815 3215 845
rect 3175 795 3185 815
rect 3205 795 3215 815
rect 3175 780 3215 795
rect 3265 865 3305 880
rect 3265 845 3275 865
rect 3295 845 3305 865
rect 3265 815 3305 845
rect 3265 795 3275 815
rect 3295 795 3305 815
rect 3265 780 3305 795
rect 3355 865 3395 880
rect 3355 845 3365 865
rect 3385 845 3395 865
rect 3355 815 3395 845
rect 3355 795 3365 815
rect 3385 795 3395 815
rect 3355 780 3395 795
rect 3445 865 3485 880
rect 3445 845 3455 865
rect 3475 845 3485 865
rect 3445 815 3485 845
rect 3445 795 3455 815
rect 3475 795 3485 815
rect 3445 780 3485 795
rect 3535 865 3575 880
rect 3535 845 3545 865
rect 3565 845 3575 865
rect 3535 815 3575 845
rect 3535 795 3545 815
rect 3565 795 3575 815
rect 3535 780 3575 795
rect 3625 865 3665 880
rect 3625 845 3635 865
rect 3655 845 3665 865
rect 3625 815 3665 845
rect 3625 795 3635 815
rect 3655 795 3665 815
rect 3625 780 3665 795
rect 3715 865 3755 880
rect 3715 845 3725 865
rect 3745 845 3755 865
rect 3715 815 3755 845
rect 3715 795 3725 815
rect 3745 795 3755 815
rect 3715 780 3755 795
rect 3805 865 3845 880
rect 3805 845 3815 865
rect 3835 845 3845 865
rect 3805 815 3845 845
rect 3805 795 3815 815
rect 3835 795 3845 815
rect 3805 780 3845 795
rect 3895 865 3935 880
rect 3895 845 3905 865
rect 3925 845 3935 865
rect 3895 815 3935 845
rect 3895 795 3905 815
rect 3925 795 3935 815
rect 3895 780 3935 795
rect 3985 865 4025 880
rect 3985 845 3995 865
rect 4015 845 4025 865
rect 3985 815 4025 845
rect 3985 795 3995 815
rect 4015 795 4025 815
rect 3985 780 4025 795
rect 4075 865 4115 880
rect 4075 845 4085 865
rect 4105 845 4115 865
rect 4075 815 4115 845
rect 4075 795 4085 815
rect 4105 795 4115 815
rect 4075 780 4115 795
rect 4165 865 4205 880
rect 4165 845 4175 865
rect 4195 845 4205 865
rect 4165 815 4205 845
rect 4165 795 4175 815
rect 4195 795 4205 815
rect 4165 780 4205 795
rect 4255 865 4295 880
rect 4255 845 4265 865
rect 4285 845 4295 865
rect 4255 815 4295 845
rect 4255 795 4265 815
rect 4285 795 4295 815
rect 4255 780 4295 795
rect 4345 865 4385 880
rect 4345 845 4355 865
rect 4375 845 4385 865
rect 4345 815 4385 845
rect 4345 795 4355 815
rect 4375 795 4385 815
rect 4345 780 4385 795
rect 4435 865 4475 880
rect 4435 845 4445 865
rect 4465 845 4475 865
rect 4435 815 4475 845
rect 4435 795 4445 815
rect 4465 795 4475 815
rect 4435 780 4475 795
rect 4525 865 4565 880
rect 4525 845 4535 865
rect 4555 845 4565 865
rect 4525 815 4565 845
rect 4525 795 4535 815
rect 4555 795 4565 815
rect 4525 780 4565 795
rect 4615 865 4655 880
rect 4615 845 4625 865
rect 4645 845 4655 865
rect 4615 815 4655 845
rect 4615 795 4625 815
rect 4645 795 4655 815
rect 4615 780 4655 795
rect 4705 865 4745 880
rect 4705 845 4715 865
rect 4735 845 4745 865
rect 4705 815 4745 845
rect 4705 795 4715 815
rect 4735 795 4745 815
rect 4705 780 4745 795
rect 4795 865 4835 880
rect 4795 845 4805 865
rect 4825 845 4835 865
rect 4795 815 4835 845
rect 4795 795 4805 815
rect 4825 795 4835 815
rect 4795 780 4835 795
rect 4885 865 4925 880
rect 4885 845 4895 865
rect 4915 845 4925 865
rect 4885 815 4925 845
rect 4885 795 4895 815
rect 4915 795 4925 815
rect 4885 780 4925 795
rect 4975 865 5015 880
rect 4975 845 4985 865
rect 5005 845 5015 865
rect 4975 815 5015 845
rect 4975 795 4985 815
rect 5005 795 5015 815
rect 4975 780 5015 795
rect 11260 730 11300 745
rect 11260 710 11270 730
rect 11290 710 11300 730
rect 11260 680 11300 710
rect 11260 660 11270 680
rect 11290 660 11300 680
rect 11260 645 11300 660
rect 11490 730 11530 745
rect 11490 710 11500 730
rect 11520 710 11530 730
rect 11490 680 11530 710
rect 11880 735 11920 750
rect 11880 715 11890 735
rect 11910 715 11920 735
rect 11880 700 11920 715
rect 11935 735 11975 750
rect 11935 715 11945 735
rect 11965 715 11975 735
rect 11935 700 11975 715
rect 11990 735 12030 750
rect 11990 715 12000 735
rect 12020 715 12030 735
rect 11990 700 12030 715
rect 12045 735 12085 750
rect 12045 715 12055 735
rect 12075 715 12085 735
rect 12045 700 12085 715
rect 12100 735 12140 750
rect 12100 715 12110 735
rect 12130 715 12140 735
rect 12100 700 12140 715
rect 12155 735 12195 750
rect 12155 715 12165 735
rect 12185 715 12195 735
rect 12155 700 12195 715
rect 12210 735 12250 750
rect 12210 715 12220 735
rect 12240 715 12250 735
rect 12210 700 12250 715
rect 12265 735 12305 750
rect 12265 715 12275 735
rect 12295 715 12305 735
rect 12265 700 12305 715
rect 12320 735 12360 750
rect 12320 715 12330 735
rect 12350 715 12360 735
rect 12320 700 12360 715
rect 12375 735 12415 750
rect 12375 715 12385 735
rect 12405 715 12415 735
rect 12375 700 12415 715
rect 12430 735 12470 750
rect 12430 715 12440 735
rect 12460 715 12470 735
rect 12430 700 12470 715
rect 12485 735 12525 750
rect 12485 715 12495 735
rect 12515 715 12525 735
rect 12485 700 12525 715
rect 12540 735 12580 750
rect 12540 715 12550 735
rect 12570 715 12580 735
rect 12540 700 12580 715
rect 11490 660 11500 680
rect 11520 660 11530 680
rect 11490 645 11530 660
rect 10955 -1450 10980 -1420
rect 10820 -1485 10860 -1450
rect 10820 -1505 10830 -1485
rect 10850 -1505 10860 -1485
rect 10820 -1535 10860 -1505
rect 10820 -1555 10830 -1535
rect 10850 -1555 10860 -1535
rect 10820 -1585 10860 -1555
rect 10820 -1605 10830 -1585
rect 10850 -1605 10860 -1585
rect 10820 -1635 10860 -1605
rect 10820 -1655 10830 -1635
rect 10850 -1655 10860 -1635
rect 10820 -1685 10860 -1655
rect 10820 -1705 10830 -1685
rect 10850 -1705 10860 -1685
rect 10490 -1735 10530 -1707
rect 10490 -1755 10500 -1735
rect 10520 -1755 10530 -1735
rect 10490 -1770 10530 -1755
rect 10550 -1730 10590 -1707
rect 10550 -1750 10560 -1730
rect 10580 -1750 10590 -1730
rect 10550 -1770 10590 -1750
rect 10610 -1730 10650 -1707
rect 10610 -1750 10620 -1730
rect 10640 -1750 10650 -1730
rect 10610 -1770 10650 -1750
rect 10670 -1735 10710 -1707
rect 10670 -1755 10680 -1735
rect 10700 -1755 10710 -1735
rect 10670 -1770 10710 -1755
rect 10820 -1735 10860 -1705
rect 10820 -1755 10830 -1735
rect 10850 -1755 10860 -1735
rect 10820 -1770 10860 -1755
rect 10880 -1485 10920 -1450
rect 10880 -1505 10890 -1485
rect 10910 -1505 10920 -1485
rect 10880 -1535 10920 -1505
rect 10880 -1555 10890 -1535
rect 10910 -1555 10920 -1535
rect 10880 -1585 10920 -1555
rect 10880 -1605 10890 -1585
rect 10910 -1605 10920 -1585
rect 10880 -1635 10920 -1605
rect 10880 -1655 10890 -1635
rect 10910 -1655 10920 -1635
rect 10880 -1685 10920 -1655
rect 10880 -1705 10890 -1685
rect 10910 -1705 10920 -1685
rect 10880 -1735 10920 -1705
rect 10880 -1755 10890 -1735
rect 10910 -1755 10920 -1735
rect 10880 -1770 10920 -1755
rect 10940 -1485 10980 -1450
rect 10940 -1505 10950 -1485
rect 10970 -1505 10980 -1485
rect 10940 -1535 10980 -1505
rect 10940 -1555 10950 -1535
rect 10970 -1555 10980 -1535
rect 10940 -1585 10980 -1555
rect 10940 -1605 10950 -1585
rect 10970 -1605 10980 -1585
rect 10940 -1635 10980 -1605
rect 10940 -1655 10950 -1635
rect 10970 -1655 10980 -1635
rect 10940 -1685 10980 -1655
rect 10940 -1705 10950 -1685
rect 10970 -1705 10980 -1685
rect 10940 -1735 10980 -1705
rect 10940 -1755 10950 -1735
rect 10970 -1755 10980 -1735
rect 10940 -1770 10980 -1755
rect 11000 -1435 11040 -1420
rect 11000 -1455 11010 -1435
rect 11030 -1455 11040 -1435
rect 11000 -1485 11040 -1455
rect 11000 -1505 11010 -1485
rect 11030 -1505 11040 -1485
rect 11000 -1535 11040 -1505
rect 11000 -1555 11010 -1535
rect 11030 -1555 11040 -1535
rect 11000 -1585 11040 -1555
rect 11000 -1605 11010 -1585
rect 11030 -1605 11040 -1585
rect 11000 -1635 11040 -1605
rect 11000 -1655 11010 -1635
rect 11030 -1655 11040 -1635
rect 11000 -1685 11040 -1655
rect 11000 -1705 11010 -1685
rect 11030 -1705 11040 -1685
rect 11000 -1735 11040 -1705
rect 11000 -1755 11010 -1735
rect 11030 -1755 11040 -1735
rect 11000 -1770 11040 -1755
rect 11060 -1435 11100 -1420
rect 11060 -1455 11070 -1435
rect 11090 -1455 11100 -1435
rect 11060 -1485 11100 -1455
rect 11060 -1505 11070 -1485
rect 11090 -1505 11100 -1485
rect 11060 -1535 11100 -1505
rect 11060 -1555 11070 -1535
rect 11090 -1555 11100 -1535
rect 11060 -1585 11100 -1555
rect 11060 -1605 11070 -1585
rect 11090 -1605 11100 -1585
rect 11060 -1635 11100 -1605
rect 11060 -1655 11070 -1635
rect 11090 -1655 11100 -1635
rect 11060 -1685 11100 -1655
rect 11060 -1705 11070 -1685
rect 11090 -1705 11100 -1685
rect 11060 -1735 11100 -1705
rect 11060 -1755 11070 -1735
rect 11090 -1755 11100 -1735
rect 11060 -1770 11100 -1755
rect 11220 -1440 11260 -1425
rect 11220 -1460 11230 -1440
rect 11250 -1460 11260 -1440
rect 11220 -1490 11260 -1460
rect 11220 -1510 11230 -1490
rect 11250 -1510 11260 -1490
rect 11220 -1540 11260 -1510
rect 11220 -1560 11230 -1540
rect 11250 -1560 11260 -1540
rect 11220 -1590 11260 -1560
rect 11220 -1610 11230 -1590
rect 11250 -1610 11260 -1590
rect 11220 -1640 11260 -1610
rect 11220 -1660 11230 -1640
rect 11250 -1660 11260 -1640
rect 11220 -1690 11260 -1660
rect 11220 -1710 11230 -1690
rect 11250 -1710 11260 -1690
rect 11220 -1740 11260 -1710
rect 11220 -1760 11230 -1740
rect 11250 -1760 11260 -1740
rect 11220 -1790 11260 -1760
rect 11220 -1810 11230 -1790
rect 11250 -1810 11260 -1790
rect 11220 -1825 11260 -1810
rect 11280 -1440 11320 -1425
rect 11280 -1460 11290 -1440
rect 11310 -1460 11320 -1440
rect 11280 -1490 11320 -1460
rect 11280 -1510 11290 -1490
rect 11310 -1510 11320 -1490
rect 11280 -1540 11320 -1510
rect 11280 -1560 11290 -1540
rect 11310 -1560 11320 -1540
rect 11280 -1590 11320 -1560
rect 11280 -1610 11290 -1590
rect 11310 -1610 11320 -1590
rect 11280 -1640 11320 -1610
rect 11280 -1660 11290 -1640
rect 11310 -1660 11320 -1640
rect 11280 -1690 11320 -1660
rect 11280 -1710 11290 -1690
rect 11310 -1710 11320 -1690
rect 11280 -1740 11320 -1710
rect 11280 -1760 11290 -1740
rect 11310 -1760 11320 -1740
rect 11280 -1790 11320 -1760
rect 11280 -1810 11290 -1790
rect 11310 -1810 11320 -1790
rect 11280 -1825 11320 -1810
rect 11340 -1440 11380 -1425
rect 11340 -1460 11350 -1440
rect 11370 -1460 11380 -1440
rect 11340 -1490 11380 -1460
rect 11340 -1510 11350 -1490
rect 11370 -1510 11380 -1490
rect 11340 -1540 11380 -1510
rect 11340 -1560 11350 -1540
rect 11370 -1560 11380 -1540
rect 11340 -1590 11380 -1560
rect 11340 -1610 11350 -1590
rect 11370 -1610 11380 -1590
rect 11340 -1640 11380 -1610
rect 11340 -1660 11350 -1640
rect 11370 -1660 11380 -1640
rect 11340 -1690 11380 -1660
rect 11340 -1710 11350 -1690
rect 11370 -1710 11380 -1690
rect 11340 -1740 11380 -1710
rect 11340 -1760 11350 -1740
rect 11370 -1760 11380 -1740
rect 11340 -1790 11380 -1760
rect 11340 -1810 11350 -1790
rect 11370 -1810 11380 -1790
rect 11340 -1825 11380 -1810
rect 11400 -1440 11440 -1425
rect 11400 -1460 11410 -1440
rect 11430 -1460 11440 -1440
rect 11400 -1490 11440 -1460
rect 11400 -1510 11410 -1490
rect 11430 -1510 11440 -1490
rect 11400 -1540 11440 -1510
rect 11400 -1560 11410 -1540
rect 11430 -1560 11440 -1540
rect 11400 -1590 11440 -1560
rect 11400 -1610 11410 -1590
rect 11430 -1610 11440 -1590
rect 11400 -1640 11440 -1610
rect 11400 -1660 11410 -1640
rect 11430 -1660 11440 -1640
rect 11400 -1690 11440 -1660
rect 11400 -1710 11410 -1690
rect 11430 -1710 11440 -1690
rect 11400 -1740 11440 -1710
rect 11400 -1760 11410 -1740
rect 11430 -1760 11440 -1740
rect 11400 -1790 11440 -1760
rect 11400 -1810 11410 -1790
rect 11430 -1810 11440 -1790
rect 11400 -1825 11440 -1810
rect 11460 -1440 11500 -1425
rect 11460 -1460 11470 -1440
rect 11490 -1460 11500 -1440
rect 11460 -1490 11500 -1460
rect 11460 -1510 11470 -1490
rect 11490 -1510 11500 -1490
rect 11460 -1540 11500 -1510
rect 11460 -1560 11470 -1540
rect 11490 -1560 11500 -1540
rect 11460 -1590 11500 -1560
rect 11460 -1610 11470 -1590
rect 11490 -1610 11500 -1590
rect 11460 -1640 11500 -1610
rect 11460 -1660 11470 -1640
rect 11490 -1660 11500 -1640
rect 11460 -1690 11500 -1660
rect 11460 -1710 11470 -1690
rect 11490 -1710 11500 -1690
rect 11460 -1740 11500 -1710
rect 11460 -1760 11470 -1740
rect 11490 -1760 11500 -1740
rect 11460 -1790 11500 -1760
rect 11460 -1810 11470 -1790
rect 11490 -1810 11500 -1790
rect 11460 -1825 11500 -1810
rect 11520 -1440 11560 -1425
rect 11520 -1460 11530 -1440
rect 11550 -1460 11560 -1440
rect 11520 -1490 11560 -1460
rect 11520 -1510 11530 -1490
rect 11550 -1510 11560 -1490
rect 11520 -1540 11560 -1510
rect 11520 -1560 11530 -1540
rect 11550 -1560 11560 -1540
rect 11520 -1590 11560 -1560
rect 11520 -1610 11530 -1590
rect 11550 -1610 11560 -1590
rect 11520 -1640 11560 -1610
rect 11520 -1660 11530 -1640
rect 11550 -1660 11560 -1640
rect 11520 -1690 11560 -1660
rect 11520 -1710 11530 -1690
rect 11550 -1710 11560 -1690
rect 11520 -1740 11560 -1710
rect 11520 -1760 11530 -1740
rect 11550 -1760 11560 -1740
rect 11520 -1790 11560 -1760
rect 11520 -1810 11530 -1790
rect 11550 -1810 11560 -1790
rect 11520 -1825 11560 -1810
rect 11580 -1440 11620 -1425
rect 11580 -1460 11590 -1440
rect 11610 -1460 11620 -1440
rect 11580 -1490 11620 -1460
rect 11580 -1510 11590 -1490
rect 11610 -1510 11620 -1490
rect 11580 -1540 11620 -1510
rect 11580 -1560 11590 -1540
rect 11610 -1560 11620 -1540
rect 11580 -1590 11620 -1560
rect 11580 -1610 11590 -1590
rect 11610 -1610 11620 -1590
rect 11580 -1640 11620 -1610
rect 11580 -1660 11590 -1640
rect 11610 -1660 11620 -1640
rect 11580 -1690 11620 -1660
rect 11580 -1710 11590 -1690
rect 11610 -1710 11620 -1690
rect 11580 -1740 11620 -1710
rect 11580 -1760 11590 -1740
rect 11610 -1760 11620 -1740
rect 11580 -1790 11620 -1760
rect 11580 -1810 11590 -1790
rect 11610 -1810 11620 -1790
rect 11580 -1825 11620 -1810
rect 11640 -1440 11680 -1425
rect 11640 -1460 11650 -1440
rect 11670 -1460 11680 -1440
rect 11640 -1490 11680 -1460
rect 11640 -1510 11650 -1490
rect 11670 -1510 11680 -1490
rect 11640 -1540 11680 -1510
rect 11640 -1560 11650 -1540
rect 11670 -1560 11680 -1540
rect 11640 -1590 11680 -1560
rect 11640 -1610 11650 -1590
rect 11670 -1610 11680 -1590
rect 11640 -1640 11680 -1610
rect 11640 -1660 11650 -1640
rect 11670 -1660 11680 -1640
rect 11640 -1690 11680 -1660
rect 11640 -1710 11650 -1690
rect 11670 -1710 11680 -1690
rect 11640 -1740 11680 -1710
rect 11640 -1760 11650 -1740
rect 11670 -1760 11680 -1740
rect 11640 -1790 11680 -1760
rect 11640 -1810 11650 -1790
rect 11670 -1810 11680 -1790
rect 11640 -1825 11680 -1810
rect 11700 -1440 11740 -1425
rect 11700 -1460 11710 -1440
rect 11730 -1460 11740 -1440
rect 11700 -1490 11740 -1460
rect 11700 -1510 11710 -1490
rect 11730 -1510 11740 -1490
rect 11700 -1540 11740 -1510
rect 11700 -1560 11710 -1540
rect 11730 -1560 11740 -1540
rect 11700 -1590 11740 -1560
rect 11700 -1610 11710 -1590
rect 11730 -1610 11740 -1590
rect 11700 -1640 11740 -1610
rect 11700 -1660 11710 -1640
rect 11730 -1660 11740 -1640
rect 11700 -1690 11740 -1660
rect 11700 -1710 11710 -1690
rect 11730 -1710 11740 -1690
rect 11700 -1740 11740 -1710
rect 11700 -1760 11710 -1740
rect 11730 -1760 11740 -1740
rect 11700 -1790 11740 -1760
rect 11700 -1810 11710 -1790
rect 11730 -1810 11740 -1790
rect 11700 -1825 11740 -1810
rect 11760 -1440 11800 -1425
rect 11760 -1460 11770 -1440
rect 11790 -1460 11800 -1440
rect 11760 -1490 11800 -1460
rect 11760 -1510 11770 -1490
rect 11790 -1510 11800 -1490
rect 11760 -1540 11800 -1510
rect 11760 -1560 11770 -1540
rect 11790 -1560 11800 -1540
rect 11760 -1590 11800 -1560
rect 11760 -1610 11770 -1590
rect 11790 -1610 11800 -1590
rect 11760 -1640 11800 -1610
rect 11760 -1660 11770 -1640
rect 11790 -1660 11800 -1640
rect 11760 -1690 11800 -1660
rect 11760 -1710 11770 -1690
rect 11790 -1710 11800 -1690
rect 11760 -1740 11800 -1710
rect 11760 -1760 11770 -1740
rect 11790 -1760 11800 -1740
rect 11760 -1790 11800 -1760
rect 11760 -1810 11770 -1790
rect 11790 -1810 11800 -1790
rect 11760 -1825 11800 -1810
rect 11820 -1440 11860 -1425
rect 11820 -1460 11830 -1440
rect 11850 -1460 11860 -1440
rect 11820 -1490 11860 -1460
rect 11820 -1510 11830 -1490
rect 11850 -1510 11860 -1490
rect 11820 -1540 11860 -1510
rect 11820 -1560 11830 -1540
rect 11850 -1560 11860 -1540
rect 11820 -1590 11860 -1560
rect 11820 -1610 11830 -1590
rect 11850 -1610 11860 -1590
rect 11820 -1640 11860 -1610
rect 11820 -1660 11830 -1640
rect 11850 -1660 11860 -1640
rect 11820 -1690 11860 -1660
rect 11820 -1710 11830 -1690
rect 11850 -1710 11860 -1690
rect 11820 -1740 11860 -1710
rect 11820 -1760 11830 -1740
rect 11850 -1760 11860 -1740
rect 11820 -1790 11860 -1760
rect 11820 -1810 11830 -1790
rect 11850 -1810 11860 -1790
rect 11820 -1825 11860 -1810
rect 11880 -1440 11920 -1425
rect 11880 -1460 11890 -1440
rect 11910 -1460 11920 -1440
rect 11880 -1490 11920 -1460
rect 11880 -1510 11890 -1490
rect 11910 -1510 11920 -1490
rect 11880 -1540 11920 -1510
rect 11880 -1560 11890 -1540
rect 11910 -1560 11920 -1540
rect 11880 -1590 11920 -1560
rect 11880 -1610 11890 -1590
rect 11910 -1610 11920 -1590
rect 11880 -1640 11920 -1610
rect 11880 -1660 11890 -1640
rect 11910 -1660 11920 -1640
rect 11880 -1690 11920 -1660
rect 11880 -1710 11890 -1690
rect 11910 -1710 11920 -1690
rect 11880 -1740 11920 -1710
rect 11880 -1760 11890 -1740
rect 11910 -1760 11920 -1740
rect 11880 -1790 11920 -1760
rect 11880 -1810 11890 -1790
rect 11910 -1810 11920 -1790
rect 11880 -1825 11920 -1810
rect 11940 -1440 11980 -1425
rect 11940 -1460 11950 -1440
rect 11970 -1460 11980 -1440
rect 11940 -1490 11980 -1460
rect 11940 -1510 11950 -1490
rect 11970 -1510 11980 -1490
rect 11940 -1540 11980 -1510
rect 11940 -1560 11950 -1540
rect 11970 -1560 11980 -1540
rect 11940 -1590 11980 -1560
rect 11940 -1610 11950 -1590
rect 11970 -1610 11980 -1590
rect 11940 -1640 11980 -1610
rect 11940 -1660 11950 -1640
rect 11970 -1660 11980 -1640
rect 11940 -1690 11980 -1660
rect 11940 -1710 11950 -1690
rect 11970 -1710 11980 -1690
rect 11940 -1740 11980 -1710
rect 11940 -1760 11950 -1740
rect 11970 -1760 11980 -1740
rect 11940 -1790 11980 -1760
rect 11940 -1810 11950 -1790
rect 11970 -1810 11980 -1790
rect 11940 -1825 11980 -1810
rect 12000 -1440 12040 -1425
rect 12000 -1460 12010 -1440
rect 12030 -1460 12040 -1440
rect 12000 -1490 12040 -1460
rect 12000 -1510 12010 -1490
rect 12030 -1510 12040 -1490
rect 12000 -1540 12040 -1510
rect 12000 -1560 12010 -1540
rect 12030 -1560 12040 -1540
rect 12000 -1590 12040 -1560
rect 12000 -1610 12010 -1590
rect 12030 -1610 12040 -1590
rect 12000 -1640 12040 -1610
rect 12000 -1660 12010 -1640
rect 12030 -1660 12040 -1640
rect 12000 -1690 12040 -1660
rect 12000 -1710 12010 -1690
rect 12030 -1710 12040 -1690
rect 12000 -1740 12040 -1710
rect 12000 -1760 12010 -1740
rect 12030 -1760 12040 -1740
rect 12000 -1790 12040 -1760
rect 12000 -1810 12010 -1790
rect 12030 -1810 12040 -1790
rect 12000 -1825 12040 -1810
rect 12060 -1440 12100 -1425
rect 12060 -1460 12070 -1440
rect 12090 -1460 12100 -1440
rect 12060 -1490 12100 -1460
rect 12060 -1510 12070 -1490
rect 12090 -1510 12100 -1490
rect 12060 -1540 12100 -1510
rect 12060 -1560 12070 -1540
rect 12090 -1560 12100 -1540
rect 12060 -1590 12100 -1560
rect 12060 -1610 12070 -1590
rect 12090 -1610 12100 -1590
rect 12060 -1640 12100 -1610
rect 12060 -1660 12070 -1640
rect 12090 -1660 12100 -1640
rect 12060 -1690 12100 -1660
rect 12060 -1710 12070 -1690
rect 12090 -1710 12100 -1690
rect 12060 -1740 12100 -1710
rect 12060 -1760 12070 -1740
rect 12090 -1760 12100 -1740
rect 12060 -1790 12100 -1760
rect 12060 -1810 12070 -1790
rect 12090 -1810 12100 -1790
rect 12060 -1825 12100 -1810
rect 12120 -1440 12160 -1425
rect 12120 -1460 12130 -1440
rect 12150 -1460 12160 -1440
rect 12120 -1490 12160 -1460
rect 12120 -1510 12130 -1490
rect 12150 -1510 12160 -1490
rect 12120 -1540 12160 -1510
rect 12120 -1560 12130 -1540
rect 12150 -1560 12160 -1540
rect 12120 -1590 12160 -1560
rect 12120 -1610 12130 -1590
rect 12150 -1610 12160 -1590
rect 12120 -1640 12160 -1610
rect 12120 -1660 12130 -1640
rect 12150 -1660 12160 -1640
rect 12120 -1690 12160 -1660
rect 12120 -1710 12130 -1690
rect 12150 -1710 12160 -1690
rect 12120 -1740 12160 -1710
rect 12120 -1760 12130 -1740
rect 12150 -1760 12160 -1740
rect 12120 -1790 12160 -1760
rect 12120 -1810 12130 -1790
rect 12150 -1810 12160 -1790
rect 12120 -1825 12160 -1810
rect 12180 -1440 12220 -1425
rect 12180 -1460 12190 -1440
rect 12210 -1460 12220 -1440
rect 12180 -1490 12220 -1460
rect 12180 -1510 12190 -1490
rect 12210 -1510 12220 -1490
rect 12180 -1540 12220 -1510
rect 12180 -1560 12190 -1540
rect 12210 -1560 12220 -1540
rect 12180 -1590 12220 -1560
rect 12180 -1610 12190 -1590
rect 12210 -1610 12220 -1590
rect 12180 -1640 12220 -1610
rect 12180 -1660 12190 -1640
rect 12210 -1660 12220 -1640
rect 12180 -1690 12220 -1660
rect 12180 -1710 12190 -1690
rect 12210 -1710 12220 -1690
rect 12180 -1740 12220 -1710
rect 12180 -1760 12190 -1740
rect 12210 -1760 12220 -1740
rect 12180 -1790 12220 -1760
rect 12180 -1810 12190 -1790
rect 12210 -1810 12220 -1790
rect 12180 -1825 12220 -1810
rect 12240 -1440 12280 -1425
rect 12240 -1460 12250 -1440
rect 12270 -1460 12280 -1440
rect 12240 -1490 12280 -1460
rect 12240 -1510 12250 -1490
rect 12270 -1510 12280 -1490
rect 12240 -1540 12280 -1510
rect 12240 -1560 12250 -1540
rect 12270 -1560 12280 -1540
rect 12240 -1590 12280 -1560
rect 12240 -1610 12250 -1590
rect 12270 -1610 12280 -1590
rect 12240 -1640 12280 -1610
rect 12240 -1660 12250 -1640
rect 12270 -1660 12280 -1640
rect 12240 -1690 12280 -1660
rect 12240 -1710 12250 -1690
rect 12270 -1710 12280 -1690
rect 12240 -1740 12280 -1710
rect 12240 -1760 12250 -1740
rect 12270 -1760 12280 -1740
rect 12240 -1790 12280 -1760
rect 12240 -1810 12250 -1790
rect 12270 -1810 12280 -1790
rect 12240 -1825 12280 -1810
rect 12300 -1440 12340 -1425
rect 12300 -1460 12310 -1440
rect 12330 -1460 12340 -1440
rect 12300 -1490 12340 -1460
rect 12300 -1510 12310 -1490
rect 12330 -1510 12340 -1490
rect 12300 -1540 12340 -1510
rect 12300 -1560 12310 -1540
rect 12330 -1560 12340 -1540
rect 12300 -1590 12340 -1560
rect 12300 -1610 12310 -1590
rect 12330 -1610 12340 -1590
rect 12300 -1640 12340 -1610
rect 12300 -1660 12310 -1640
rect 12330 -1660 12340 -1640
rect 12300 -1690 12340 -1660
rect 12300 -1710 12310 -1690
rect 12330 -1710 12340 -1690
rect 12300 -1740 12340 -1710
rect 12300 -1760 12310 -1740
rect 12330 -1760 12340 -1740
rect 12300 -1790 12340 -1760
rect 12300 -1810 12310 -1790
rect 12330 -1810 12340 -1790
rect 12300 -1825 12340 -1810
rect 12360 -1440 12400 -1425
rect 12360 -1460 12370 -1440
rect 12390 -1460 12400 -1440
rect 12360 -1490 12400 -1460
rect 12360 -1510 12370 -1490
rect 12390 -1510 12400 -1490
rect 12360 -1540 12400 -1510
rect 12360 -1560 12370 -1540
rect 12390 -1560 12400 -1540
rect 12360 -1590 12400 -1560
rect 12360 -1610 12370 -1590
rect 12390 -1610 12400 -1590
rect 12360 -1640 12400 -1610
rect 12360 -1660 12370 -1640
rect 12390 -1660 12400 -1640
rect 12360 -1690 12400 -1660
rect 12360 -1710 12370 -1690
rect 12390 -1710 12400 -1690
rect 12360 -1740 12400 -1710
rect 12360 -1760 12370 -1740
rect 12390 -1760 12400 -1740
rect 12360 -1790 12400 -1760
rect 12360 -1810 12370 -1790
rect 12390 -1810 12400 -1790
rect 12360 -1825 12400 -1810
rect 12420 -1440 12460 -1425
rect 12420 -1460 12430 -1440
rect 12450 -1460 12460 -1440
rect 12420 -1490 12460 -1460
rect 12420 -1510 12430 -1490
rect 12450 -1510 12460 -1490
rect 12420 -1540 12460 -1510
rect 12420 -1560 12430 -1540
rect 12450 -1560 12460 -1540
rect 12420 -1590 12460 -1560
rect 12420 -1610 12430 -1590
rect 12450 -1610 12460 -1590
rect 12420 -1640 12460 -1610
rect 12420 -1660 12430 -1640
rect 12450 -1660 12460 -1640
rect 12420 -1690 12460 -1660
rect 12420 -1710 12430 -1690
rect 12450 -1710 12460 -1690
rect 12420 -1740 12460 -1710
rect 12420 -1760 12430 -1740
rect 12450 -1760 12460 -1740
rect 12420 -1790 12460 -1760
rect 12420 -1810 12430 -1790
rect 12450 -1810 12460 -1790
rect 12420 -1825 12460 -1810
rect 12480 -1440 12520 -1425
rect 12480 -1460 12490 -1440
rect 12510 -1460 12520 -1440
rect 12480 -1490 12520 -1460
rect 12480 -1510 12490 -1490
rect 12510 -1510 12520 -1490
rect 12480 -1540 12520 -1510
rect 12480 -1560 12490 -1540
rect 12510 -1560 12520 -1540
rect 12480 -1590 12520 -1560
rect 12480 -1610 12490 -1590
rect 12510 -1610 12520 -1590
rect 12480 -1640 12520 -1610
rect 12480 -1660 12490 -1640
rect 12510 -1660 12520 -1640
rect 12480 -1690 12520 -1660
rect 12480 -1710 12490 -1690
rect 12510 -1710 12520 -1690
rect 12480 -1740 12520 -1710
rect 12480 -1760 12490 -1740
rect 12510 -1760 12520 -1740
rect 12480 -1790 12520 -1760
rect 12480 -1810 12490 -1790
rect 12510 -1810 12520 -1790
rect 12480 -1825 12520 -1810
rect 12540 -1440 12580 -1425
rect 12540 -1460 12550 -1440
rect 12570 -1460 12580 -1440
rect 12540 -1490 12580 -1460
rect 12540 -1510 12550 -1490
rect 12570 -1510 12580 -1490
rect 12540 -1540 12580 -1510
rect 12540 -1560 12550 -1540
rect 12570 -1560 12580 -1540
rect 12540 -1590 12580 -1560
rect 12540 -1610 12550 -1590
rect 12570 -1610 12580 -1590
rect 12540 -1640 12580 -1610
rect 12540 -1660 12550 -1640
rect 12570 -1660 12580 -1640
rect 12540 -1690 12580 -1660
rect 12540 -1710 12550 -1690
rect 12570 -1710 12580 -1690
rect 12540 -1740 12580 -1710
rect 12540 -1760 12550 -1740
rect 12570 -1760 12580 -1740
rect 12540 -1790 12580 -1760
rect 12540 -1810 12550 -1790
rect 12570 -1810 12580 -1790
rect 12540 -1825 12580 -1810
rect 12895 -2030 12935 -2015
rect 12895 -2050 12905 -2030
rect 12925 -2050 12935 -2030
rect 12895 -2080 12935 -2050
rect 12895 -2100 12905 -2080
rect 12925 -2100 12935 -2080
rect 11220 -2120 11260 -2105
rect 11220 -2140 11230 -2120
rect 11250 -2140 11260 -2120
rect 11220 -2170 11260 -2140
rect 11220 -2190 11230 -2170
rect 11250 -2190 11260 -2170
rect 11220 -2220 11260 -2190
rect 11220 -2240 11230 -2220
rect 11250 -2240 11260 -2220
rect 11220 -2270 11260 -2240
rect 11220 -2290 11230 -2270
rect 11250 -2290 11260 -2270
rect 11220 -2320 11260 -2290
rect 11220 -2340 11230 -2320
rect 11250 -2340 11260 -2320
rect 11220 -2370 11260 -2340
rect 11220 -2390 11230 -2370
rect 11250 -2390 11260 -2370
rect 11220 -2420 11260 -2390
rect 11220 -2440 11230 -2420
rect 11250 -2440 11260 -2420
rect 11220 -2470 11260 -2440
rect 11220 -2490 11230 -2470
rect 11250 -2490 11260 -2470
rect 11220 -2505 11260 -2490
rect 11280 -2120 11320 -2105
rect 11280 -2140 11290 -2120
rect 11310 -2140 11320 -2120
rect 11280 -2170 11320 -2140
rect 11280 -2190 11290 -2170
rect 11310 -2190 11320 -2170
rect 11280 -2220 11320 -2190
rect 11280 -2240 11290 -2220
rect 11310 -2240 11320 -2220
rect 11280 -2270 11320 -2240
rect 11280 -2290 11290 -2270
rect 11310 -2290 11320 -2270
rect 11280 -2320 11320 -2290
rect 11280 -2340 11290 -2320
rect 11310 -2340 11320 -2320
rect 11280 -2370 11320 -2340
rect 11280 -2390 11290 -2370
rect 11310 -2390 11320 -2370
rect 11280 -2420 11320 -2390
rect 11280 -2440 11290 -2420
rect 11310 -2440 11320 -2420
rect 11280 -2470 11320 -2440
rect 11280 -2490 11290 -2470
rect 11310 -2490 11320 -2470
rect 11280 -2505 11320 -2490
rect 11340 -2120 11380 -2105
rect 11340 -2140 11350 -2120
rect 11370 -2140 11380 -2120
rect 11340 -2170 11380 -2140
rect 11340 -2190 11350 -2170
rect 11370 -2190 11380 -2170
rect 11340 -2220 11380 -2190
rect 11340 -2240 11350 -2220
rect 11370 -2240 11380 -2220
rect 11340 -2270 11380 -2240
rect 11340 -2290 11350 -2270
rect 11370 -2290 11380 -2270
rect 11340 -2320 11380 -2290
rect 11340 -2340 11350 -2320
rect 11370 -2340 11380 -2320
rect 11340 -2370 11380 -2340
rect 11340 -2390 11350 -2370
rect 11370 -2390 11380 -2370
rect 11340 -2420 11380 -2390
rect 11340 -2440 11350 -2420
rect 11370 -2440 11380 -2420
rect 11340 -2470 11380 -2440
rect 11340 -2490 11350 -2470
rect 11370 -2490 11380 -2470
rect 11340 -2505 11380 -2490
rect 11400 -2120 11440 -2105
rect 11400 -2140 11410 -2120
rect 11430 -2140 11440 -2120
rect 11400 -2170 11440 -2140
rect 11400 -2190 11410 -2170
rect 11430 -2190 11440 -2170
rect 11400 -2220 11440 -2190
rect 11400 -2240 11410 -2220
rect 11430 -2240 11440 -2220
rect 11400 -2270 11440 -2240
rect 11400 -2290 11410 -2270
rect 11430 -2290 11440 -2270
rect 11400 -2320 11440 -2290
rect 11400 -2340 11410 -2320
rect 11430 -2340 11440 -2320
rect 11400 -2370 11440 -2340
rect 11400 -2390 11410 -2370
rect 11430 -2390 11440 -2370
rect 11400 -2420 11440 -2390
rect 11400 -2440 11410 -2420
rect 11430 -2440 11440 -2420
rect 11400 -2470 11440 -2440
rect 11400 -2490 11410 -2470
rect 11430 -2490 11440 -2470
rect 11400 -2505 11440 -2490
rect 11460 -2120 11500 -2105
rect 11460 -2140 11470 -2120
rect 11490 -2140 11500 -2120
rect 11460 -2170 11500 -2140
rect 11460 -2190 11470 -2170
rect 11490 -2190 11500 -2170
rect 11460 -2220 11500 -2190
rect 11460 -2240 11470 -2220
rect 11490 -2240 11500 -2220
rect 11460 -2270 11500 -2240
rect 11460 -2290 11470 -2270
rect 11490 -2290 11500 -2270
rect 11460 -2320 11500 -2290
rect 11460 -2340 11470 -2320
rect 11490 -2340 11500 -2320
rect 11460 -2370 11500 -2340
rect 11460 -2390 11470 -2370
rect 11490 -2390 11500 -2370
rect 11460 -2420 11500 -2390
rect 11460 -2440 11470 -2420
rect 11490 -2440 11500 -2420
rect 11460 -2470 11500 -2440
rect 11460 -2490 11470 -2470
rect 11490 -2490 11500 -2470
rect 11460 -2505 11500 -2490
rect 11520 -2120 11560 -2105
rect 11520 -2140 11530 -2120
rect 11550 -2140 11560 -2120
rect 11520 -2170 11560 -2140
rect 11520 -2190 11530 -2170
rect 11550 -2190 11560 -2170
rect 11520 -2220 11560 -2190
rect 11520 -2240 11530 -2220
rect 11550 -2240 11560 -2220
rect 11520 -2270 11560 -2240
rect 11520 -2290 11530 -2270
rect 11550 -2290 11560 -2270
rect 11520 -2320 11560 -2290
rect 11520 -2340 11530 -2320
rect 11550 -2340 11560 -2320
rect 11520 -2370 11560 -2340
rect 11520 -2390 11530 -2370
rect 11550 -2390 11560 -2370
rect 11520 -2420 11560 -2390
rect 11520 -2440 11530 -2420
rect 11550 -2440 11560 -2420
rect 11520 -2470 11560 -2440
rect 11520 -2490 11530 -2470
rect 11550 -2490 11560 -2470
rect 11520 -2505 11560 -2490
rect 11580 -2120 11620 -2105
rect 11580 -2140 11590 -2120
rect 11610 -2140 11620 -2120
rect 11580 -2170 11620 -2140
rect 11580 -2190 11590 -2170
rect 11610 -2190 11620 -2170
rect 11580 -2220 11620 -2190
rect 11580 -2240 11590 -2220
rect 11610 -2240 11620 -2220
rect 11580 -2270 11620 -2240
rect 11580 -2290 11590 -2270
rect 11610 -2290 11620 -2270
rect 11580 -2320 11620 -2290
rect 11580 -2340 11590 -2320
rect 11610 -2340 11620 -2320
rect 11580 -2370 11620 -2340
rect 11580 -2390 11590 -2370
rect 11610 -2390 11620 -2370
rect 11580 -2420 11620 -2390
rect 11580 -2440 11590 -2420
rect 11610 -2440 11620 -2420
rect 11580 -2470 11620 -2440
rect 11580 -2490 11590 -2470
rect 11610 -2490 11620 -2470
rect 11580 -2505 11620 -2490
rect 11640 -2120 11680 -2105
rect 11640 -2140 11650 -2120
rect 11670 -2140 11680 -2120
rect 11640 -2170 11680 -2140
rect 11640 -2190 11650 -2170
rect 11670 -2190 11680 -2170
rect 11640 -2220 11680 -2190
rect 11640 -2240 11650 -2220
rect 11670 -2240 11680 -2220
rect 11640 -2270 11680 -2240
rect 11640 -2290 11650 -2270
rect 11670 -2290 11680 -2270
rect 11640 -2320 11680 -2290
rect 11640 -2340 11650 -2320
rect 11670 -2340 11680 -2320
rect 11640 -2370 11680 -2340
rect 11640 -2390 11650 -2370
rect 11670 -2390 11680 -2370
rect 11640 -2420 11680 -2390
rect 11640 -2440 11650 -2420
rect 11670 -2440 11680 -2420
rect 11640 -2470 11680 -2440
rect 11640 -2490 11650 -2470
rect 11670 -2490 11680 -2470
rect 11640 -2505 11680 -2490
rect 11700 -2120 11740 -2105
rect 11700 -2140 11710 -2120
rect 11730 -2140 11740 -2120
rect 11700 -2170 11740 -2140
rect 11700 -2190 11710 -2170
rect 11730 -2190 11740 -2170
rect 11700 -2220 11740 -2190
rect 11700 -2240 11710 -2220
rect 11730 -2240 11740 -2220
rect 11700 -2270 11740 -2240
rect 11700 -2290 11710 -2270
rect 11730 -2290 11740 -2270
rect 11700 -2320 11740 -2290
rect 11700 -2340 11710 -2320
rect 11730 -2340 11740 -2320
rect 11700 -2370 11740 -2340
rect 11700 -2390 11710 -2370
rect 11730 -2390 11740 -2370
rect 11700 -2420 11740 -2390
rect 11700 -2440 11710 -2420
rect 11730 -2440 11740 -2420
rect 11700 -2470 11740 -2440
rect 11700 -2490 11710 -2470
rect 11730 -2490 11740 -2470
rect 11700 -2505 11740 -2490
rect 11760 -2120 11800 -2105
rect 11760 -2140 11770 -2120
rect 11790 -2140 11800 -2120
rect 11760 -2170 11800 -2140
rect 11760 -2190 11770 -2170
rect 11790 -2190 11800 -2170
rect 11760 -2220 11800 -2190
rect 11760 -2240 11770 -2220
rect 11790 -2240 11800 -2220
rect 11760 -2270 11800 -2240
rect 11760 -2290 11770 -2270
rect 11790 -2290 11800 -2270
rect 11760 -2320 11800 -2290
rect 11760 -2340 11770 -2320
rect 11790 -2340 11800 -2320
rect 11760 -2370 11800 -2340
rect 11760 -2390 11770 -2370
rect 11790 -2390 11800 -2370
rect 11760 -2420 11800 -2390
rect 11760 -2440 11770 -2420
rect 11790 -2440 11800 -2420
rect 11760 -2470 11800 -2440
rect 11760 -2490 11770 -2470
rect 11790 -2490 11800 -2470
rect 11760 -2505 11800 -2490
rect 11820 -2120 11860 -2105
rect 11820 -2140 11830 -2120
rect 11850 -2140 11860 -2120
rect 11820 -2170 11860 -2140
rect 11820 -2190 11830 -2170
rect 11850 -2190 11860 -2170
rect 11820 -2220 11860 -2190
rect 11820 -2240 11830 -2220
rect 11850 -2240 11860 -2220
rect 11820 -2270 11860 -2240
rect 11820 -2290 11830 -2270
rect 11850 -2290 11860 -2270
rect 11820 -2320 11860 -2290
rect 11820 -2340 11830 -2320
rect 11850 -2340 11860 -2320
rect 11820 -2370 11860 -2340
rect 11820 -2390 11830 -2370
rect 11850 -2390 11860 -2370
rect 11820 -2420 11860 -2390
rect 11820 -2440 11830 -2420
rect 11850 -2440 11860 -2420
rect 11820 -2470 11860 -2440
rect 11820 -2490 11830 -2470
rect 11850 -2490 11860 -2470
rect 11820 -2505 11860 -2490
rect 11880 -2120 11920 -2105
rect 11880 -2140 11890 -2120
rect 11910 -2140 11920 -2120
rect 11880 -2170 11920 -2140
rect 11880 -2190 11890 -2170
rect 11910 -2190 11920 -2170
rect 11880 -2220 11920 -2190
rect 11880 -2240 11890 -2220
rect 11910 -2240 11920 -2220
rect 11880 -2270 11920 -2240
rect 11880 -2290 11890 -2270
rect 11910 -2290 11920 -2270
rect 11880 -2320 11920 -2290
rect 11880 -2340 11890 -2320
rect 11910 -2340 11920 -2320
rect 11880 -2370 11920 -2340
rect 11880 -2390 11890 -2370
rect 11910 -2390 11920 -2370
rect 11880 -2420 11920 -2390
rect 11880 -2440 11890 -2420
rect 11910 -2440 11920 -2420
rect 11880 -2470 11920 -2440
rect 11880 -2490 11890 -2470
rect 11910 -2490 11920 -2470
rect 11880 -2505 11920 -2490
rect 11940 -2120 11980 -2105
rect 11940 -2140 11950 -2120
rect 11970 -2140 11980 -2120
rect 11940 -2170 11980 -2140
rect 11940 -2190 11950 -2170
rect 11970 -2190 11980 -2170
rect 11940 -2220 11980 -2190
rect 11940 -2240 11950 -2220
rect 11970 -2240 11980 -2220
rect 11940 -2270 11980 -2240
rect 11940 -2290 11950 -2270
rect 11970 -2290 11980 -2270
rect 11940 -2320 11980 -2290
rect 11940 -2340 11950 -2320
rect 11970 -2340 11980 -2320
rect 11940 -2370 11980 -2340
rect 11940 -2390 11950 -2370
rect 11970 -2390 11980 -2370
rect 11940 -2420 11980 -2390
rect 11940 -2440 11950 -2420
rect 11970 -2440 11980 -2420
rect 11940 -2470 11980 -2440
rect 11940 -2490 11950 -2470
rect 11970 -2490 11980 -2470
rect 11940 -2505 11980 -2490
rect 12000 -2120 12040 -2105
rect 12000 -2140 12010 -2120
rect 12030 -2140 12040 -2120
rect 12000 -2170 12040 -2140
rect 12000 -2190 12010 -2170
rect 12030 -2190 12040 -2170
rect 12000 -2220 12040 -2190
rect 12000 -2240 12010 -2220
rect 12030 -2240 12040 -2220
rect 12000 -2270 12040 -2240
rect 12000 -2290 12010 -2270
rect 12030 -2290 12040 -2270
rect 12000 -2320 12040 -2290
rect 12000 -2340 12010 -2320
rect 12030 -2340 12040 -2320
rect 12000 -2370 12040 -2340
rect 12000 -2390 12010 -2370
rect 12030 -2390 12040 -2370
rect 12000 -2420 12040 -2390
rect 12000 -2440 12010 -2420
rect 12030 -2440 12040 -2420
rect 12000 -2470 12040 -2440
rect 12000 -2490 12010 -2470
rect 12030 -2490 12040 -2470
rect 12000 -2505 12040 -2490
rect 12060 -2120 12100 -2105
rect 12060 -2140 12070 -2120
rect 12090 -2140 12100 -2120
rect 12060 -2170 12100 -2140
rect 12060 -2190 12070 -2170
rect 12090 -2190 12100 -2170
rect 12060 -2220 12100 -2190
rect 12060 -2240 12070 -2220
rect 12090 -2240 12100 -2220
rect 12060 -2270 12100 -2240
rect 12060 -2290 12070 -2270
rect 12090 -2290 12100 -2270
rect 12060 -2320 12100 -2290
rect 12060 -2340 12070 -2320
rect 12090 -2340 12100 -2320
rect 12060 -2370 12100 -2340
rect 12060 -2390 12070 -2370
rect 12090 -2390 12100 -2370
rect 12060 -2420 12100 -2390
rect 12060 -2440 12070 -2420
rect 12090 -2440 12100 -2420
rect 12060 -2470 12100 -2440
rect 12060 -2490 12070 -2470
rect 12090 -2490 12100 -2470
rect 12060 -2505 12100 -2490
rect 12120 -2120 12160 -2105
rect 12120 -2140 12130 -2120
rect 12150 -2140 12160 -2120
rect 12120 -2170 12160 -2140
rect 12120 -2190 12130 -2170
rect 12150 -2190 12160 -2170
rect 12120 -2220 12160 -2190
rect 12120 -2240 12130 -2220
rect 12150 -2240 12160 -2220
rect 12120 -2270 12160 -2240
rect 12120 -2290 12130 -2270
rect 12150 -2290 12160 -2270
rect 12120 -2320 12160 -2290
rect 12120 -2340 12130 -2320
rect 12150 -2340 12160 -2320
rect 12120 -2370 12160 -2340
rect 12120 -2390 12130 -2370
rect 12150 -2390 12160 -2370
rect 12120 -2420 12160 -2390
rect 12120 -2440 12130 -2420
rect 12150 -2440 12160 -2420
rect 12120 -2470 12160 -2440
rect 12120 -2490 12130 -2470
rect 12150 -2490 12160 -2470
rect 12120 -2505 12160 -2490
rect 12180 -2120 12220 -2105
rect 12180 -2140 12190 -2120
rect 12210 -2140 12220 -2120
rect 12180 -2170 12220 -2140
rect 12180 -2190 12190 -2170
rect 12210 -2190 12220 -2170
rect 12180 -2220 12220 -2190
rect 12180 -2240 12190 -2220
rect 12210 -2240 12220 -2220
rect 12180 -2270 12220 -2240
rect 12180 -2290 12190 -2270
rect 12210 -2290 12220 -2270
rect 12180 -2320 12220 -2290
rect 12180 -2340 12190 -2320
rect 12210 -2340 12220 -2320
rect 12180 -2370 12220 -2340
rect 12180 -2390 12190 -2370
rect 12210 -2390 12220 -2370
rect 12180 -2420 12220 -2390
rect 12180 -2440 12190 -2420
rect 12210 -2440 12220 -2420
rect 12180 -2470 12220 -2440
rect 12180 -2490 12190 -2470
rect 12210 -2490 12220 -2470
rect 12180 -2505 12220 -2490
rect 12240 -2120 12280 -2105
rect 12240 -2140 12250 -2120
rect 12270 -2140 12280 -2120
rect 12240 -2170 12280 -2140
rect 12240 -2190 12250 -2170
rect 12270 -2190 12280 -2170
rect 12240 -2220 12280 -2190
rect 12240 -2240 12250 -2220
rect 12270 -2240 12280 -2220
rect 12240 -2270 12280 -2240
rect 12240 -2290 12250 -2270
rect 12270 -2290 12280 -2270
rect 12240 -2320 12280 -2290
rect 12240 -2340 12250 -2320
rect 12270 -2340 12280 -2320
rect 12240 -2370 12280 -2340
rect 12240 -2390 12250 -2370
rect 12270 -2390 12280 -2370
rect 12240 -2420 12280 -2390
rect 12240 -2440 12250 -2420
rect 12270 -2440 12280 -2420
rect 12240 -2470 12280 -2440
rect 12240 -2490 12250 -2470
rect 12270 -2490 12280 -2470
rect 12240 -2505 12280 -2490
rect 12300 -2120 12340 -2105
rect 12300 -2140 12310 -2120
rect 12330 -2140 12340 -2120
rect 12300 -2170 12340 -2140
rect 12300 -2190 12310 -2170
rect 12330 -2190 12340 -2170
rect 12300 -2220 12340 -2190
rect 12300 -2240 12310 -2220
rect 12330 -2240 12340 -2220
rect 12300 -2270 12340 -2240
rect 12300 -2290 12310 -2270
rect 12330 -2290 12340 -2270
rect 12300 -2320 12340 -2290
rect 12300 -2340 12310 -2320
rect 12330 -2340 12340 -2320
rect 12300 -2370 12340 -2340
rect 12300 -2390 12310 -2370
rect 12330 -2390 12340 -2370
rect 12300 -2420 12340 -2390
rect 12300 -2440 12310 -2420
rect 12330 -2440 12340 -2420
rect 12300 -2470 12340 -2440
rect 12300 -2490 12310 -2470
rect 12330 -2490 12340 -2470
rect 12300 -2505 12340 -2490
rect 12360 -2120 12400 -2105
rect 12360 -2140 12370 -2120
rect 12390 -2140 12400 -2120
rect 12360 -2170 12400 -2140
rect 12360 -2190 12370 -2170
rect 12390 -2190 12400 -2170
rect 12360 -2220 12400 -2190
rect 12360 -2240 12370 -2220
rect 12390 -2240 12400 -2220
rect 12360 -2270 12400 -2240
rect 12360 -2290 12370 -2270
rect 12390 -2290 12400 -2270
rect 12360 -2320 12400 -2290
rect 12360 -2340 12370 -2320
rect 12390 -2340 12400 -2320
rect 12360 -2370 12400 -2340
rect 12360 -2390 12370 -2370
rect 12390 -2390 12400 -2370
rect 12360 -2420 12400 -2390
rect 12360 -2440 12370 -2420
rect 12390 -2440 12400 -2420
rect 12360 -2470 12400 -2440
rect 12360 -2490 12370 -2470
rect 12390 -2490 12400 -2470
rect 12360 -2505 12400 -2490
rect 12420 -2120 12460 -2105
rect 12420 -2140 12430 -2120
rect 12450 -2140 12460 -2120
rect 12420 -2170 12460 -2140
rect 12420 -2190 12430 -2170
rect 12450 -2190 12460 -2170
rect 12420 -2220 12460 -2190
rect 12420 -2240 12430 -2220
rect 12450 -2240 12460 -2220
rect 12420 -2270 12460 -2240
rect 12420 -2290 12430 -2270
rect 12450 -2290 12460 -2270
rect 12420 -2320 12460 -2290
rect 12420 -2340 12430 -2320
rect 12450 -2340 12460 -2320
rect 12420 -2370 12460 -2340
rect 12420 -2390 12430 -2370
rect 12450 -2390 12460 -2370
rect 12420 -2420 12460 -2390
rect 12420 -2440 12430 -2420
rect 12450 -2440 12460 -2420
rect 12420 -2470 12460 -2440
rect 12420 -2490 12430 -2470
rect 12450 -2490 12460 -2470
rect 12420 -2505 12460 -2490
rect 12480 -2120 12520 -2105
rect 12480 -2140 12490 -2120
rect 12510 -2140 12520 -2120
rect 12480 -2170 12520 -2140
rect 12480 -2190 12490 -2170
rect 12510 -2190 12520 -2170
rect 12480 -2220 12520 -2190
rect 12480 -2240 12490 -2220
rect 12510 -2240 12520 -2220
rect 12480 -2270 12520 -2240
rect 12480 -2290 12490 -2270
rect 12510 -2290 12520 -2270
rect 12480 -2320 12520 -2290
rect 12480 -2340 12490 -2320
rect 12510 -2340 12520 -2320
rect 12480 -2370 12520 -2340
rect 12480 -2390 12490 -2370
rect 12510 -2390 12520 -2370
rect 12480 -2420 12520 -2390
rect 12480 -2440 12490 -2420
rect 12510 -2440 12520 -2420
rect 12480 -2470 12520 -2440
rect 12480 -2490 12490 -2470
rect 12510 -2490 12520 -2470
rect 12480 -2505 12520 -2490
rect 12540 -2120 12580 -2105
rect 12540 -2140 12550 -2120
rect 12570 -2140 12580 -2120
rect 12540 -2170 12580 -2140
rect 12540 -2190 12550 -2170
rect 12570 -2190 12580 -2170
rect 12540 -2220 12580 -2190
rect 12540 -2240 12550 -2220
rect 12570 -2240 12580 -2220
rect 12540 -2270 12580 -2240
rect 12540 -2290 12550 -2270
rect 12570 -2290 12580 -2270
rect 12540 -2320 12580 -2290
rect 12895 -2130 12935 -2100
rect 12895 -2150 12905 -2130
rect 12925 -2150 12935 -2130
rect 12895 -2180 12935 -2150
rect 12895 -2200 12905 -2180
rect 12925 -2200 12935 -2180
rect 12895 -2230 12935 -2200
rect 12895 -2250 12905 -2230
rect 12925 -2250 12935 -2230
rect 12895 -2280 12935 -2250
rect 12895 -2300 12905 -2280
rect 12925 -2300 12935 -2280
rect 12895 -2315 12935 -2300
rect 12950 -2030 12990 -2015
rect 12950 -2050 12960 -2030
rect 12980 -2050 12990 -2030
rect 12950 -2080 12990 -2050
rect 12950 -2100 12960 -2080
rect 12980 -2100 12990 -2080
rect 12950 -2130 12990 -2100
rect 12950 -2150 12960 -2130
rect 12980 -2150 12990 -2130
rect 12950 -2180 12990 -2150
rect 12950 -2200 12960 -2180
rect 12980 -2200 12990 -2180
rect 12950 -2230 12990 -2200
rect 12950 -2250 12960 -2230
rect 12980 -2250 12990 -2230
rect 12950 -2280 12990 -2250
rect 12950 -2300 12960 -2280
rect 12980 -2300 12990 -2280
rect 12950 -2315 12990 -2300
rect 13005 -2030 13045 -2015
rect 13005 -2050 13015 -2030
rect 13035 -2050 13045 -2030
rect 13005 -2080 13045 -2050
rect 13005 -2100 13015 -2080
rect 13035 -2100 13045 -2080
rect 13005 -2130 13045 -2100
rect 13005 -2150 13015 -2130
rect 13035 -2150 13045 -2130
rect 13005 -2180 13045 -2150
rect 13005 -2200 13015 -2180
rect 13035 -2200 13045 -2180
rect 13005 -2230 13045 -2200
rect 13005 -2250 13015 -2230
rect 13035 -2250 13045 -2230
rect 13005 -2280 13045 -2250
rect 13005 -2300 13015 -2280
rect 13035 -2300 13045 -2280
rect 13005 -2315 13045 -2300
rect 13060 -2030 13100 -2015
rect 13060 -2050 13070 -2030
rect 13090 -2050 13100 -2030
rect 13060 -2080 13100 -2050
rect 13060 -2100 13070 -2080
rect 13090 -2100 13100 -2080
rect 13060 -2130 13100 -2100
rect 13060 -2150 13070 -2130
rect 13090 -2150 13100 -2130
rect 13060 -2180 13100 -2150
rect 13060 -2200 13070 -2180
rect 13090 -2200 13100 -2180
rect 13060 -2230 13100 -2200
rect 13060 -2250 13070 -2230
rect 13090 -2250 13100 -2230
rect 13060 -2280 13100 -2250
rect 13060 -2300 13070 -2280
rect 13090 -2300 13100 -2280
rect 13060 -2315 13100 -2300
rect 13115 -2030 13155 -2015
rect 13115 -2050 13125 -2030
rect 13145 -2050 13155 -2030
rect 13115 -2080 13155 -2050
rect 13115 -2100 13125 -2080
rect 13145 -2100 13155 -2080
rect 13115 -2130 13155 -2100
rect 13115 -2150 13125 -2130
rect 13145 -2150 13155 -2130
rect 13115 -2180 13155 -2150
rect 13115 -2200 13125 -2180
rect 13145 -2200 13155 -2180
rect 13115 -2230 13155 -2200
rect 13115 -2250 13125 -2230
rect 13145 -2250 13155 -2230
rect 13115 -2280 13155 -2250
rect 13115 -2300 13125 -2280
rect 13145 -2300 13155 -2280
rect 13115 -2315 13155 -2300
rect 13170 -2030 13210 -2015
rect 13170 -2050 13180 -2030
rect 13200 -2050 13210 -2030
rect 13170 -2080 13210 -2050
rect 13170 -2100 13180 -2080
rect 13200 -2100 13210 -2080
rect 13170 -2130 13210 -2100
rect 13170 -2150 13180 -2130
rect 13200 -2150 13210 -2130
rect 13170 -2180 13210 -2150
rect 13170 -2200 13180 -2180
rect 13200 -2200 13210 -2180
rect 13170 -2230 13210 -2200
rect 13170 -2250 13180 -2230
rect 13200 -2250 13210 -2230
rect 13170 -2280 13210 -2250
rect 13170 -2300 13180 -2280
rect 13200 -2300 13210 -2280
rect 13170 -2315 13210 -2300
rect 13225 -2030 13265 -2015
rect 13225 -2050 13235 -2030
rect 13255 -2050 13265 -2030
rect 13225 -2080 13265 -2050
rect 13225 -2100 13235 -2080
rect 13255 -2100 13265 -2080
rect 13225 -2130 13265 -2100
rect 13225 -2150 13235 -2130
rect 13255 -2150 13265 -2130
rect 13225 -2180 13265 -2150
rect 13225 -2200 13235 -2180
rect 13255 -2200 13265 -2180
rect 13225 -2230 13265 -2200
rect 13225 -2250 13235 -2230
rect 13255 -2250 13265 -2230
rect 13225 -2280 13265 -2250
rect 13225 -2300 13235 -2280
rect 13255 -2300 13265 -2280
rect 13225 -2315 13265 -2300
rect 13280 -2030 13320 -2015
rect 13280 -2050 13290 -2030
rect 13310 -2050 13320 -2030
rect 13280 -2080 13320 -2050
rect 13280 -2100 13290 -2080
rect 13310 -2100 13320 -2080
rect 13280 -2130 13320 -2100
rect 13280 -2150 13290 -2130
rect 13310 -2150 13320 -2130
rect 13280 -2180 13320 -2150
rect 13280 -2200 13290 -2180
rect 13310 -2200 13320 -2180
rect 13280 -2230 13320 -2200
rect 13280 -2250 13290 -2230
rect 13310 -2250 13320 -2230
rect 13280 -2280 13320 -2250
rect 13280 -2300 13290 -2280
rect 13310 -2300 13320 -2280
rect 13280 -2315 13320 -2300
rect 13335 -2030 13375 -2015
rect 13335 -2050 13345 -2030
rect 13365 -2050 13375 -2030
rect 13335 -2080 13375 -2050
rect 13335 -2100 13345 -2080
rect 13365 -2100 13375 -2080
rect 13335 -2130 13375 -2100
rect 13335 -2150 13345 -2130
rect 13365 -2150 13375 -2130
rect 13335 -2180 13375 -2150
rect 13335 -2200 13345 -2180
rect 13365 -2200 13375 -2180
rect 13335 -2230 13375 -2200
rect 13335 -2250 13345 -2230
rect 13365 -2250 13375 -2230
rect 13335 -2280 13375 -2250
rect 13335 -2300 13345 -2280
rect 13365 -2300 13375 -2280
rect 13335 -2315 13375 -2300
rect 13390 -2030 13430 -2015
rect 13390 -2050 13400 -2030
rect 13420 -2050 13430 -2030
rect 13390 -2080 13430 -2050
rect 13390 -2100 13400 -2080
rect 13420 -2100 13430 -2080
rect 13390 -2130 13430 -2100
rect 13390 -2150 13400 -2130
rect 13420 -2150 13430 -2130
rect 13390 -2180 13430 -2150
rect 13390 -2200 13400 -2180
rect 13420 -2200 13430 -2180
rect 13390 -2230 13430 -2200
rect 13390 -2250 13400 -2230
rect 13420 -2250 13430 -2230
rect 13390 -2280 13430 -2250
rect 13390 -2300 13400 -2280
rect 13420 -2300 13430 -2280
rect 13390 -2315 13430 -2300
rect 13445 -2030 13485 -2015
rect 13445 -2050 13455 -2030
rect 13475 -2050 13485 -2030
rect 13445 -2080 13485 -2050
rect 13445 -2100 13455 -2080
rect 13475 -2100 13485 -2080
rect 13445 -2130 13485 -2100
rect 13445 -2150 13455 -2130
rect 13475 -2150 13485 -2130
rect 13445 -2180 13485 -2150
rect 13445 -2200 13455 -2180
rect 13475 -2200 13485 -2180
rect 13445 -2230 13485 -2200
rect 13445 -2250 13455 -2230
rect 13475 -2250 13485 -2230
rect 13445 -2280 13485 -2250
rect 13445 -2300 13455 -2280
rect 13475 -2300 13485 -2280
rect 13445 -2315 13485 -2300
rect 13500 -2030 13540 -2015
rect 13500 -2050 13510 -2030
rect 13530 -2050 13540 -2030
rect 13500 -2080 13540 -2050
rect 13500 -2100 13510 -2080
rect 13530 -2100 13540 -2080
rect 13500 -2130 13540 -2100
rect 13500 -2150 13510 -2130
rect 13530 -2150 13540 -2130
rect 13500 -2180 13540 -2150
rect 13500 -2200 13510 -2180
rect 13530 -2200 13540 -2180
rect 13500 -2230 13540 -2200
rect 13500 -2250 13510 -2230
rect 13530 -2250 13540 -2230
rect 13500 -2280 13540 -2250
rect 13500 -2300 13510 -2280
rect 13530 -2300 13540 -2280
rect 13500 -2315 13540 -2300
rect 13555 -2030 13595 -2015
rect 13555 -2050 13565 -2030
rect 13585 -2050 13595 -2030
rect 13555 -2080 13595 -2050
rect 13555 -2100 13565 -2080
rect 13585 -2100 13595 -2080
rect 13555 -2130 13595 -2100
rect 13555 -2150 13565 -2130
rect 13585 -2150 13595 -2130
rect 13555 -2180 13595 -2150
rect 13555 -2200 13565 -2180
rect 13585 -2200 13595 -2180
rect 13555 -2230 13595 -2200
rect 13555 -2250 13565 -2230
rect 13585 -2250 13595 -2230
rect 13555 -2280 13595 -2250
rect 13555 -2300 13565 -2280
rect 13585 -2300 13595 -2280
rect 13555 -2315 13595 -2300
rect 13610 -2030 13650 -2015
rect 13610 -2050 13620 -2030
rect 13640 -2050 13650 -2030
rect 13610 -2080 13650 -2050
rect 13610 -2100 13620 -2080
rect 13640 -2100 13650 -2080
rect 13610 -2130 13650 -2100
rect 13610 -2150 13620 -2130
rect 13640 -2150 13650 -2130
rect 13610 -2180 13650 -2150
rect 13610 -2200 13620 -2180
rect 13640 -2200 13650 -2180
rect 13610 -2230 13650 -2200
rect 13610 -2250 13620 -2230
rect 13640 -2250 13650 -2230
rect 13610 -2280 13650 -2250
rect 13610 -2300 13620 -2280
rect 13640 -2300 13650 -2280
rect 13610 -2315 13650 -2300
rect 13665 -2030 13705 -2015
rect 13665 -2050 13675 -2030
rect 13695 -2050 13705 -2030
rect 13665 -2080 13705 -2050
rect 13665 -2100 13675 -2080
rect 13695 -2100 13705 -2080
rect 13665 -2130 13705 -2100
rect 13665 -2150 13675 -2130
rect 13695 -2150 13705 -2130
rect 13665 -2180 13705 -2150
rect 13665 -2200 13675 -2180
rect 13695 -2200 13705 -2180
rect 13665 -2230 13705 -2200
rect 13665 -2250 13675 -2230
rect 13695 -2250 13705 -2230
rect 13665 -2280 13705 -2250
rect 13665 -2300 13675 -2280
rect 13695 -2300 13705 -2280
rect 13665 -2315 13705 -2300
rect 13720 -2030 13760 -2015
rect 13720 -2050 13730 -2030
rect 13750 -2050 13760 -2030
rect 13720 -2080 13760 -2050
rect 13720 -2100 13730 -2080
rect 13750 -2100 13760 -2080
rect 13720 -2130 13760 -2100
rect 13720 -2150 13730 -2130
rect 13750 -2150 13760 -2130
rect 13720 -2180 13760 -2150
rect 13720 -2200 13730 -2180
rect 13750 -2200 13760 -2180
rect 13720 -2230 13760 -2200
rect 13720 -2250 13730 -2230
rect 13750 -2250 13760 -2230
rect 13720 -2280 13760 -2250
rect 13720 -2300 13730 -2280
rect 13750 -2300 13760 -2280
rect 13720 -2315 13760 -2300
rect 13775 -2030 13815 -2015
rect 13775 -2050 13785 -2030
rect 13805 -2050 13815 -2030
rect 13775 -2080 13815 -2050
rect 13775 -2100 13785 -2080
rect 13805 -2100 13815 -2080
rect 13775 -2130 13815 -2100
rect 13775 -2150 13785 -2130
rect 13805 -2150 13815 -2130
rect 13775 -2180 13815 -2150
rect 13775 -2200 13785 -2180
rect 13805 -2200 13815 -2180
rect 13775 -2230 13815 -2200
rect 13775 -2250 13785 -2230
rect 13805 -2250 13815 -2230
rect 13775 -2280 13815 -2250
rect 13775 -2300 13785 -2280
rect 13805 -2300 13815 -2280
rect 13775 -2315 13815 -2300
rect 13830 -2030 13870 -2015
rect 13830 -2050 13840 -2030
rect 13860 -2050 13870 -2030
rect 13830 -2080 13870 -2050
rect 13830 -2100 13840 -2080
rect 13860 -2100 13870 -2080
rect 13830 -2130 13870 -2100
rect 13830 -2150 13840 -2130
rect 13860 -2150 13870 -2130
rect 13830 -2180 13870 -2150
rect 13830 -2200 13840 -2180
rect 13860 -2200 13870 -2180
rect 13830 -2230 13870 -2200
rect 13830 -2250 13840 -2230
rect 13860 -2250 13870 -2230
rect 13830 -2280 13870 -2250
rect 13830 -2300 13840 -2280
rect 13860 -2300 13870 -2280
rect 13830 -2315 13870 -2300
rect 13885 -2030 13925 -2015
rect 13885 -2050 13895 -2030
rect 13915 -2050 13925 -2030
rect 13885 -2080 13925 -2050
rect 13885 -2100 13895 -2080
rect 13915 -2100 13925 -2080
rect 13885 -2130 13925 -2100
rect 13885 -2150 13895 -2130
rect 13915 -2150 13925 -2130
rect 13885 -2180 13925 -2150
rect 13885 -2200 13895 -2180
rect 13915 -2200 13925 -2180
rect 13885 -2230 13925 -2200
rect 13885 -2250 13895 -2230
rect 13915 -2250 13925 -2230
rect 13885 -2280 13925 -2250
rect 13885 -2300 13895 -2280
rect 13915 -2300 13925 -2280
rect 13885 -2315 13925 -2300
rect 13940 -2030 13980 -2015
rect 13940 -2050 13950 -2030
rect 13970 -2050 13980 -2030
rect 13940 -2080 13980 -2050
rect 13940 -2100 13950 -2080
rect 13970 -2100 13980 -2080
rect 13940 -2130 13980 -2100
rect 13940 -2150 13950 -2130
rect 13970 -2150 13980 -2130
rect 13940 -2180 13980 -2150
rect 13940 -2200 13950 -2180
rect 13970 -2200 13980 -2180
rect 13940 -2230 13980 -2200
rect 13940 -2250 13950 -2230
rect 13970 -2250 13980 -2230
rect 13940 -2280 13980 -2250
rect 13940 -2300 13950 -2280
rect 13970 -2300 13980 -2280
rect 13940 -2315 13980 -2300
rect 13995 -2030 14035 -2015
rect 13995 -2050 14005 -2030
rect 14025 -2050 14035 -2030
rect 13995 -2080 14035 -2050
rect 13995 -2100 14005 -2080
rect 14025 -2100 14035 -2080
rect 13995 -2130 14035 -2100
rect 13995 -2150 14005 -2130
rect 14025 -2150 14035 -2130
rect 13995 -2180 14035 -2150
rect 13995 -2200 14005 -2180
rect 14025 -2200 14035 -2180
rect 13995 -2230 14035 -2200
rect 13995 -2250 14005 -2230
rect 14025 -2250 14035 -2230
rect 13995 -2280 14035 -2250
rect 13995 -2300 14005 -2280
rect 14025 -2300 14035 -2280
rect 13995 -2315 14035 -2300
rect 14050 -2030 14090 -2015
rect 14050 -2050 14060 -2030
rect 14080 -2050 14090 -2030
rect 14050 -2080 14090 -2050
rect 14050 -2100 14060 -2080
rect 14080 -2100 14090 -2080
rect 14050 -2130 14090 -2100
rect 14050 -2150 14060 -2130
rect 14080 -2150 14090 -2130
rect 14050 -2180 14090 -2150
rect 14050 -2200 14060 -2180
rect 14080 -2200 14090 -2180
rect 14050 -2230 14090 -2200
rect 14050 -2250 14060 -2230
rect 14080 -2250 14090 -2230
rect 14050 -2280 14090 -2250
rect 14050 -2300 14060 -2280
rect 14080 -2300 14090 -2280
rect 14050 -2315 14090 -2300
rect 14105 -2030 14145 -2015
rect 14105 -2050 14115 -2030
rect 14135 -2050 14145 -2030
rect 14105 -2080 14145 -2050
rect 14105 -2100 14115 -2080
rect 14135 -2100 14145 -2080
rect 14105 -2130 14145 -2100
rect 14105 -2150 14115 -2130
rect 14135 -2150 14145 -2130
rect 14105 -2180 14145 -2150
rect 14105 -2200 14115 -2180
rect 14135 -2200 14145 -2180
rect 14105 -2230 14145 -2200
rect 14105 -2250 14115 -2230
rect 14135 -2250 14145 -2230
rect 14105 -2280 14145 -2250
rect 14105 -2300 14115 -2280
rect 14135 -2300 14145 -2280
rect 14105 -2315 14145 -2300
rect 12540 -2340 12550 -2320
rect 12570 -2340 12580 -2320
rect 12540 -2370 12580 -2340
rect 12540 -2390 12550 -2370
rect 12570 -2390 12580 -2370
rect 12540 -2420 12580 -2390
rect 12540 -2440 12550 -2420
rect 12570 -2440 12580 -2420
rect 12540 -2470 12580 -2440
rect 12540 -2490 12550 -2470
rect 12570 -2490 12580 -2470
rect 12540 -2505 12580 -2490
rect 12895 -2460 12935 -2445
rect 12895 -2480 12905 -2460
rect 12925 -2480 12935 -2460
rect 12895 -2510 12935 -2480
rect 12895 -2530 12905 -2510
rect 12925 -2530 12935 -2510
rect 12895 -2545 12935 -2530
rect 12950 -2460 12990 -2445
rect 12950 -2480 12960 -2460
rect 12980 -2480 12990 -2460
rect 12950 -2510 12990 -2480
rect 12950 -2530 12960 -2510
rect 12980 -2530 12990 -2510
rect 12950 -2545 12990 -2530
rect 13005 -2460 13045 -2445
rect 13005 -2480 13015 -2460
rect 13035 -2480 13045 -2460
rect 13005 -2510 13045 -2480
rect 13005 -2530 13015 -2510
rect 13035 -2530 13045 -2510
rect 13005 -2545 13045 -2530
rect 13060 -2460 13100 -2445
rect 13060 -2480 13070 -2460
rect 13090 -2480 13100 -2460
rect 13060 -2510 13100 -2480
rect 13060 -2530 13070 -2510
rect 13090 -2530 13100 -2510
rect 13060 -2545 13100 -2530
rect 13115 -2460 13155 -2445
rect 13115 -2480 13125 -2460
rect 13145 -2480 13155 -2460
rect 13115 -2510 13155 -2480
rect 13115 -2530 13125 -2510
rect 13145 -2530 13155 -2510
rect 13115 -2545 13155 -2530
rect 13170 -2460 13210 -2445
rect 13170 -2480 13180 -2460
rect 13200 -2480 13210 -2460
rect 13170 -2510 13210 -2480
rect 13170 -2530 13180 -2510
rect 13200 -2530 13210 -2510
rect 13170 -2545 13210 -2530
rect 13225 -2460 13265 -2445
rect 13225 -2480 13235 -2460
rect 13255 -2480 13265 -2460
rect 13225 -2510 13265 -2480
rect 13225 -2530 13235 -2510
rect 13255 -2530 13265 -2510
rect 13225 -2545 13265 -2530
rect 13280 -2460 13320 -2445
rect 13280 -2480 13290 -2460
rect 13310 -2480 13320 -2460
rect 13280 -2510 13320 -2480
rect 13280 -2530 13290 -2510
rect 13310 -2530 13320 -2510
rect 13280 -2545 13320 -2530
rect 13335 -2460 13375 -2445
rect 13335 -2480 13345 -2460
rect 13365 -2480 13375 -2460
rect 13335 -2510 13375 -2480
rect 13335 -2530 13345 -2510
rect 13365 -2530 13375 -2510
rect 13335 -2545 13375 -2530
rect 13390 -2460 13430 -2445
rect 13390 -2480 13400 -2460
rect 13420 -2480 13430 -2460
rect 13390 -2510 13430 -2480
rect 13390 -2530 13400 -2510
rect 13420 -2530 13430 -2510
rect 13390 -2545 13430 -2530
rect 13445 -2460 13485 -2445
rect 13445 -2480 13455 -2460
rect 13475 -2480 13485 -2460
rect 13445 -2510 13485 -2480
rect 13445 -2530 13455 -2510
rect 13475 -2530 13485 -2510
rect 13445 -2545 13485 -2530
rect 13500 -2460 13540 -2445
rect 13500 -2480 13510 -2460
rect 13530 -2480 13540 -2460
rect 13500 -2510 13540 -2480
rect 13500 -2530 13510 -2510
rect 13530 -2530 13540 -2510
rect 13500 -2545 13540 -2530
rect 13555 -2460 13595 -2445
rect 13555 -2480 13565 -2460
rect 13585 -2480 13595 -2460
rect 13555 -2510 13595 -2480
rect 13555 -2530 13565 -2510
rect 13585 -2530 13595 -2510
rect 13555 -2545 13595 -2530
rect 13610 -2460 13650 -2445
rect 13610 -2480 13620 -2460
rect 13640 -2480 13650 -2460
rect 13610 -2510 13650 -2480
rect 13610 -2530 13620 -2510
rect 13640 -2530 13650 -2510
rect 13610 -2545 13650 -2530
rect 13665 -2460 13705 -2445
rect 13665 -2480 13675 -2460
rect 13695 -2480 13705 -2460
rect 13665 -2510 13705 -2480
rect 13665 -2530 13675 -2510
rect 13695 -2530 13705 -2510
rect 13665 -2545 13705 -2530
rect 13720 -2460 13760 -2445
rect 13720 -2480 13730 -2460
rect 13750 -2480 13760 -2460
rect 13720 -2510 13760 -2480
rect 13720 -2530 13730 -2510
rect 13750 -2530 13760 -2510
rect 13720 -2545 13760 -2530
rect 13775 -2460 13815 -2445
rect 13775 -2480 13785 -2460
rect 13805 -2480 13815 -2460
rect 13775 -2510 13815 -2480
rect 13775 -2530 13785 -2510
rect 13805 -2530 13815 -2510
rect 13775 -2545 13815 -2530
rect 13830 -2460 13870 -2445
rect 13830 -2480 13840 -2460
rect 13860 -2480 13870 -2460
rect 13830 -2510 13870 -2480
rect 13830 -2530 13840 -2510
rect 13860 -2530 13870 -2510
rect 13830 -2545 13870 -2530
rect 13885 -2460 13925 -2445
rect 13885 -2480 13895 -2460
rect 13915 -2480 13925 -2460
rect 13885 -2510 13925 -2480
rect 13885 -2530 13895 -2510
rect 13915 -2530 13925 -2510
rect 13885 -2545 13925 -2530
rect 13940 -2460 13980 -2445
rect 13940 -2480 13950 -2460
rect 13970 -2480 13980 -2460
rect 13940 -2510 13980 -2480
rect 13940 -2530 13950 -2510
rect 13970 -2530 13980 -2510
rect 13940 -2545 13980 -2530
rect 13995 -2460 14035 -2445
rect 13995 -2480 14005 -2460
rect 14025 -2480 14035 -2460
rect 13995 -2510 14035 -2480
rect 13995 -2530 14005 -2510
rect 14025 -2530 14035 -2510
rect 13995 -2545 14035 -2530
rect 14050 -2460 14090 -2445
rect 14050 -2480 14060 -2460
rect 14080 -2480 14090 -2460
rect 14050 -2510 14090 -2480
rect 14050 -2530 14060 -2510
rect 14080 -2530 14090 -2510
rect 14050 -2545 14090 -2530
rect 14105 -2460 14145 -2445
rect 14105 -2480 14115 -2460
rect 14135 -2480 14145 -2460
rect 14105 -2510 14145 -2480
rect 14105 -2530 14115 -2510
rect 14135 -2530 14145 -2510
rect 14105 -2545 14145 -2530
rect 12895 -2750 12935 -2735
rect 12895 -2770 12905 -2750
rect 12925 -2770 12935 -2750
rect 12895 -2800 12935 -2770
rect 12895 -2820 12905 -2800
rect 12925 -2820 12935 -2800
rect 12895 -2850 12935 -2820
rect 12895 -2870 12905 -2850
rect 12925 -2870 12935 -2850
rect 11275 -2885 11315 -2870
rect 11275 -2905 11285 -2885
rect 11305 -2905 11315 -2885
rect 11275 -2935 11315 -2905
rect 11275 -2955 11285 -2935
rect 11305 -2955 11315 -2935
rect 11275 -2985 11315 -2955
rect 11275 -3005 11285 -2985
rect 11305 -3005 11315 -2985
rect 11275 -3020 11315 -3005
rect 11330 -2885 11370 -2870
rect 11330 -2905 11340 -2885
rect 11360 -2905 11370 -2885
rect 11330 -2935 11370 -2905
rect 11330 -2955 11340 -2935
rect 11360 -2955 11370 -2935
rect 11330 -2985 11370 -2955
rect 11330 -3005 11340 -2985
rect 11360 -3005 11370 -2985
rect 11330 -3020 11370 -3005
rect 11385 -2885 11425 -2870
rect 11385 -2905 11395 -2885
rect 11415 -2905 11425 -2885
rect 11385 -2935 11425 -2905
rect 11385 -2955 11395 -2935
rect 11415 -2955 11425 -2935
rect 11385 -2985 11425 -2955
rect 11385 -3005 11395 -2985
rect 11415 -3005 11425 -2985
rect 11385 -3020 11425 -3005
rect 11440 -2885 11480 -2870
rect 11440 -2905 11450 -2885
rect 11470 -2905 11480 -2885
rect 11440 -2935 11480 -2905
rect 11440 -2955 11450 -2935
rect 11470 -2955 11480 -2935
rect 11440 -2985 11480 -2955
rect 11440 -3005 11450 -2985
rect 11470 -3005 11480 -2985
rect 11440 -3020 11480 -3005
rect 11495 -2885 11535 -2870
rect 11495 -2905 11505 -2885
rect 11525 -2905 11535 -2885
rect 11495 -2935 11535 -2905
rect 11495 -2955 11505 -2935
rect 11525 -2955 11535 -2935
rect 11495 -2985 11535 -2955
rect 11495 -3005 11505 -2985
rect 11525 -3005 11535 -2985
rect 11495 -3020 11535 -3005
rect 11550 -2885 11590 -2870
rect 11550 -2905 11560 -2885
rect 11580 -2905 11590 -2885
rect 11550 -2935 11590 -2905
rect 11550 -2955 11560 -2935
rect 11580 -2955 11590 -2935
rect 11550 -2985 11590 -2955
rect 11550 -3005 11560 -2985
rect 11580 -3005 11590 -2985
rect 11550 -3020 11590 -3005
rect 11605 -2885 11645 -2870
rect 11605 -2905 11615 -2885
rect 11635 -2905 11645 -2885
rect 11605 -2935 11645 -2905
rect 11605 -2955 11615 -2935
rect 11635 -2955 11645 -2935
rect 11605 -2985 11645 -2955
rect 11605 -3005 11615 -2985
rect 11635 -3005 11645 -2985
rect 11605 -3020 11645 -3005
rect 11660 -2885 11700 -2870
rect 11660 -2905 11670 -2885
rect 11690 -2905 11700 -2885
rect 11660 -2935 11700 -2905
rect 11660 -2955 11670 -2935
rect 11690 -2955 11700 -2935
rect 11660 -2985 11700 -2955
rect 11660 -3005 11670 -2985
rect 11690 -3005 11700 -2985
rect 11660 -3020 11700 -3005
rect 11715 -2885 11755 -2870
rect 11715 -2905 11725 -2885
rect 11745 -2905 11755 -2885
rect 11715 -2935 11755 -2905
rect 11715 -2955 11725 -2935
rect 11745 -2955 11755 -2935
rect 11715 -2985 11755 -2955
rect 11715 -3005 11725 -2985
rect 11745 -3005 11755 -2985
rect 11715 -3020 11755 -3005
rect 11770 -2885 11810 -2870
rect 11770 -2905 11780 -2885
rect 11800 -2905 11810 -2885
rect 11770 -2935 11810 -2905
rect 11770 -2955 11780 -2935
rect 11800 -2955 11810 -2935
rect 11770 -2985 11810 -2955
rect 11770 -3005 11780 -2985
rect 11800 -3005 11810 -2985
rect 11770 -3020 11810 -3005
rect 11825 -2885 11865 -2870
rect 11825 -2905 11835 -2885
rect 11855 -2905 11865 -2885
rect 11825 -2935 11865 -2905
rect 11825 -2955 11835 -2935
rect 11855 -2955 11865 -2935
rect 11825 -2985 11865 -2955
rect 11825 -3005 11835 -2985
rect 11855 -3005 11865 -2985
rect 11825 -3020 11865 -3005
rect 11880 -2885 11920 -2870
rect 11880 -2905 11890 -2885
rect 11910 -2905 11920 -2885
rect 11880 -2935 11920 -2905
rect 11880 -2955 11890 -2935
rect 11910 -2955 11920 -2935
rect 11880 -2985 11920 -2955
rect 11880 -3005 11890 -2985
rect 11910 -3005 11920 -2985
rect 11880 -3020 11920 -3005
rect 11935 -2885 11975 -2870
rect 11935 -2905 11945 -2885
rect 11965 -2905 11975 -2885
rect 11935 -2935 11975 -2905
rect 11935 -2955 11945 -2935
rect 11965 -2955 11975 -2935
rect 11935 -2985 11975 -2955
rect 11935 -3005 11945 -2985
rect 11965 -3005 11975 -2985
rect 11935 -3020 11975 -3005
rect 11990 -2885 12030 -2870
rect 11990 -2905 12000 -2885
rect 12020 -2905 12030 -2885
rect 11990 -2935 12030 -2905
rect 11990 -2955 12000 -2935
rect 12020 -2955 12030 -2935
rect 11990 -2985 12030 -2955
rect 11990 -3005 12000 -2985
rect 12020 -3005 12030 -2985
rect 11990 -3020 12030 -3005
rect 12045 -2885 12085 -2870
rect 12045 -2905 12055 -2885
rect 12075 -2905 12085 -2885
rect 12045 -2935 12085 -2905
rect 12045 -2955 12055 -2935
rect 12075 -2955 12085 -2935
rect 12045 -2985 12085 -2955
rect 12045 -3005 12055 -2985
rect 12075 -3005 12085 -2985
rect 12045 -3020 12085 -3005
rect 12100 -2885 12140 -2870
rect 12100 -2905 12110 -2885
rect 12130 -2905 12140 -2885
rect 12100 -2935 12140 -2905
rect 12100 -2955 12110 -2935
rect 12130 -2955 12140 -2935
rect 12100 -2985 12140 -2955
rect 12100 -3005 12110 -2985
rect 12130 -3005 12140 -2985
rect 12100 -3020 12140 -3005
rect 12155 -2885 12195 -2870
rect 12155 -2905 12165 -2885
rect 12185 -2905 12195 -2885
rect 12155 -2935 12195 -2905
rect 12155 -2955 12165 -2935
rect 12185 -2955 12195 -2935
rect 12155 -2985 12195 -2955
rect 12155 -3005 12165 -2985
rect 12185 -3005 12195 -2985
rect 12155 -3020 12195 -3005
rect 12210 -2885 12250 -2870
rect 12210 -2905 12220 -2885
rect 12240 -2905 12250 -2885
rect 12210 -2935 12250 -2905
rect 12210 -2955 12220 -2935
rect 12240 -2955 12250 -2935
rect 12210 -2985 12250 -2955
rect 12210 -3005 12220 -2985
rect 12240 -3005 12250 -2985
rect 12210 -3020 12250 -3005
rect 12265 -2885 12305 -2870
rect 12265 -2905 12275 -2885
rect 12295 -2905 12305 -2885
rect 12265 -2935 12305 -2905
rect 12265 -2955 12275 -2935
rect 12295 -2955 12305 -2935
rect 12265 -2985 12305 -2955
rect 12265 -3005 12275 -2985
rect 12295 -3005 12305 -2985
rect 12265 -3020 12305 -3005
rect 12320 -2885 12360 -2870
rect 12320 -2905 12330 -2885
rect 12350 -2905 12360 -2885
rect 12320 -2935 12360 -2905
rect 12320 -2955 12330 -2935
rect 12350 -2955 12360 -2935
rect 12320 -2985 12360 -2955
rect 12320 -3005 12330 -2985
rect 12350 -3005 12360 -2985
rect 12320 -3020 12360 -3005
rect 12375 -2885 12415 -2870
rect 12375 -2905 12385 -2885
rect 12405 -2905 12415 -2885
rect 12375 -2935 12415 -2905
rect 12375 -2955 12385 -2935
rect 12405 -2955 12415 -2935
rect 12375 -2985 12415 -2955
rect 12375 -3005 12385 -2985
rect 12405 -3005 12415 -2985
rect 12375 -3020 12415 -3005
rect 12430 -2885 12470 -2870
rect 12430 -2905 12440 -2885
rect 12460 -2905 12470 -2885
rect 12430 -2935 12470 -2905
rect 12430 -2955 12440 -2935
rect 12460 -2955 12470 -2935
rect 12430 -2985 12470 -2955
rect 12430 -3005 12440 -2985
rect 12460 -3005 12470 -2985
rect 12430 -3020 12470 -3005
rect 12485 -2885 12525 -2870
rect 12895 -2885 12935 -2870
rect 12950 -2750 12990 -2735
rect 12950 -2770 12960 -2750
rect 12980 -2770 12990 -2750
rect 12950 -2800 12990 -2770
rect 12950 -2820 12960 -2800
rect 12980 -2820 12990 -2800
rect 12950 -2850 12990 -2820
rect 12950 -2870 12960 -2850
rect 12980 -2870 12990 -2850
rect 12950 -2885 12990 -2870
rect 13005 -2750 13045 -2735
rect 13005 -2770 13015 -2750
rect 13035 -2770 13045 -2750
rect 13005 -2800 13045 -2770
rect 13005 -2820 13015 -2800
rect 13035 -2820 13045 -2800
rect 13005 -2850 13045 -2820
rect 13005 -2870 13015 -2850
rect 13035 -2870 13045 -2850
rect 13005 -2885 13045 -2870
rect 13060 -2750 13100 -2735
rect 13060 -2770 13070 -2750
rect 13090 -2770 13100 -2750
rect 13060 -2800 13100 -2770
rect 13060 -2820 13070 -2800
rect 13090 -2820 13100 -2800
rect 13060 -2850 13100 -2820
rect 13060 -2870 13070 -2850
rect 13090 -2870 13100 -2850
rect 13060 -2885 13100 -2870
rect 13115 -2750 13155 -2735
rect 13115 -2770 13125 -2750
rect 13145 -2770 13155 -2750
rect 13115 -2800 13155 -2770
rect 13115 -2820 13125 -2800
rect 13145 -2820 13155 -2800
rect 13115 -2850 13155 -2820
rect 13115 -2870 13125 -2850
rect 13145 -2870 13155 -2850
rect 13115 -2885 13155 -2870
rect 13170 -2750 13210 -2735
rect 13170 -2770 13180 -2750
rect 13200 -2770 13210 -2750
rect 13170 -2800 13210 -2770
rect 13170 -2820 13180 -2800
rect 13200 -2820 13210 -2800
rect 13170 -2850 13210 -2820
rect 13170 -2870 13180 -2850
rect 13200 -2870 13210 -2850
rect 13170 -2885 13210 -2870
rect 13225 -2750 13265 -2735
rect 13225 -2770 13235 -2750
rect 13255 -2770 13265 -2750
rect 13225 -2800 13265 -2770
rect 13225 -2820 13235 -2800
rect 13255 -2820 13265 -2800
rect 13225 -2850 13265 -2820
rect 13225 -2870 13235 -2850
rect 13255 -2870 13265 -2850
rect 13225 -2885 13265 -2870
rect 13280 -2750 13320 -2735
rect 13280 -2770 13290 -2750
rect 13310 -2770 13320 -2750
rect 13280 -2800 13320 -2770
rect 13280 -2820 13290 -2800
rect 13310 -2820 13320 -2800
rect 13280 -2850 13320 -2820
rect 13280 -2870 13290 -2850
rect 13310 -2870 13320 -2850
rect 13280 -2885 13320 -2870
rect 13335 -2750 13375 -2735
rect 13335 -2770 13345 -2750
rect 13365 -2770 13375 -2750
rect 13335 -2800 13375 -2770
rect 13335 -2820 13345 -2800
rect 13365 -2820 13375 -2800
rect 13335 -2850 13375 -2820
rect 13335 -2870 13345 -2850
rect 13365 -2870 13375 -2850
rect 13335 -2885 13375 -2870
rect 13390 -2750 13430 -2735
rect 13390 -2770 13400 -2750
rect 13420 -2770 13430 -2750
rect 13390 -2800 13430 -2770
rect 13390 -2820 13400 -2800
rect 13420 -2820 13430 -2800
rect 13390 -2850 13430 -2820
rect 13390 -2870 13400 -2850
rect 13420 -2870 13430 -2850
rect 13390 -2885 13430 -2870
rect 13445 -2750 13485 -2735
rect 13445 -2770 13455 -2750
rect 13475 -2770 13485 -2750
rect 13445 -2800 13485 -2770
rect 13445 -2820 13455 -2800
rect 13475 -2820 13485 -2800
rect 13445 -2850 13485 -2820
rect 13445 -2870 13455 -2850
rect 13475 -2870 13485 -2850
rect 13445 -2885 13485 -2870
rect 13500 -2750 13540 -2735
rect 13500 -2770 13510 -2750
rect 13530 -2770 13540 -2750
rect 13500 -2800 13540 -2770
rect 13500 -2820 13510 -2800
rect 13530 -2820 13540 -2800
rect 13500 -2850 13540 -2820
rect 13500 -2870 13510 -2850
rect 13530 -2870 13540 -2850
rect 13500 -2885 13540 -2870
rect 13555 -2750 13595 -2735
rect 13555 -2770 13565 -2750
rect 13585 -2770 13595 -2750
rect 13555 -2800 13595 -2770
rect 13555 -2820 13565 -2800
rect 13585 -2820 13595 -2800
rect 13555 -2850 13595 -2820
rect 13555 -2870 13565 -2850
rect 13585 -2870 13595 -2850
rect 13555 -2885 13595 -2870
rect 13610 -2750 13650 -2735
rect 13610 -2770 13620 -2750
rect 13640 -2770 13650 -2750
rect 13610 -2800 13650 -2770
rect 13610 -2820 13620 -2800
rect 13640 -2820 13650 -2800
rect 13610 -2850 13650 -2820
rect 13610 -2870 13620 -2850
rect 13640 -2870 13650 -2850
rect 13610 -2885 13650 -2870
rect 13665 -2750 13705 -2735
rect 13665 -2770 13675 -2750
rect 13695 -2770 13705 -2750
rect 13665 -2800 13705 -2770
rect 13665 -2820 13675 -2800
rect 13695 -2820 13705 -2800
rect 13665 -2850 13705 -2820
rect 13665 -2870 13675 -2850
rect 13695 -2870 13705 -2850
rect 13665 -2885 13705 -2870
rect 13720 -2750 13760 -2735
rect 13720 -2770 13730 -2750
rect 13750 -2770 13760 -2750
rect 13720 -2800 13760 -2770
rect 13720 -2820 13730 -2800
rect 13750 -2820 13760 -2800
rect 13720 -2850 13760 -2820
rect 13720 -2870 13730 -2850
rect 13750 -2870 13760 -2850
rect 13720 -2885 13760 -2870
rect 13775 -2750 13815 -2735
rect 13775 -2770 13785 -2750
rect 13805 -2770 13815 -2750
rect 13775 -2800 13815 -2770
rect 13775 -2820 13785 -2800
rect 13805 -2820 13815 -2800
rect 13775 -2850 13815 -2820
rect 13775 -2870 13785 -2850
rect 13805 -2870 13815 -2850
rect 13775 -2885 13815 -2870
rect 13830 -2750 13870 -2735
rect 13830 -2770 13840 -2750
rect 13860 -2770 13870 -2750
rect 13830 -2800 13870 -2770
rect 13830 -2820 13840 -2800
rect 13860 -2820 13870 -2800
rect 13830 -2850 13870 -2820
rect 13830 -2870 13840 -2850
rect 13860 -2870 13870 -2850
rect 13830 -2885 13870 -2870
rect 13885 -2750 13925 -2735
rect 13885 -2770 13895 -2750
rect 13915 -2770 13925 -2750
rect 13885 -2800 13925 -2770
rect 13885 -2820 13895 -2800
rect 13915 -2820 13925 -2800
rect 13885 -2850 13925 -2820
rect 13885 -2870 13895 -2850
rect 13915 -2870 13925 -2850
rect 13885 -2885 13925 -2870
rect 13940 -2750 13980 -2735
rect 13940 -2770 13950 -2750
rect 13970 -2770 13980 -2750
rect 13940 -2800 13980 -2770
rect 13940 -2820 13950 -2800
rect 13970 -2820 13980 -2800
rect 13940 -2850 13980 -2820
rect 13940 -2870 13950 -2850
rect 13970 -2870 13980 -2850
rect 13940 -2885 13980 -2870
rect 13995 -2750 14035 -2735
rect 13995 -2770 14005 -2750
rect 14025 -2770 14035 -2750
rect 13995 -2800 14035 -2770
rect 13995 -2820 14005 -2800
rect 14025 -2820 14035 -2800
rect 13995 -2850 14035 -2820
rect 13995 -2870 14005 -2850
rect 14025 -2870 14035 -2850
rect 13995 -2885 14035 -2870
rect 14050 -2750 14090 -2735
rect 14050 -2770 14060 -2750
rect 14080 -2770 14090 -2750
rect 14050 -2800 14090 -2770
rect 14050 -2820 14060 -2800
rect 14080 -2820 14090 -2800
rect 14050 -2850 14090 -2820
rect 14050 -2870 14060 -2850
rect 14080 -2870 14090 -2850
rect 14050 -2885 14090 -2870
rect 14105 -2750 14145 -2735
rect 14105 -2770 14115 -2750
rect 14135 -2770 14145 -2750
rect 14105 -2800 14145 -2770
rect 14105 -2820 14115 -2800
rect 14135 -2820 14145 -2800
rect 14105 -2850 14145 -2820
rect 14105 -2870 14115 -2850
rect 14135 -2870 14145 -2850
rect 14105 -2885 14145 -2870
rect 12485 -2905 12495 -2885
rect 12515 -2905 12525 -2885
rect 12485 -2935 12525 -2905
rect 12485 -2955 12495 -2935
rect 12515 -2955 12525 -2935
rect 12485 -2985 12525 -2955
rect 12485 -3005 12495 -2985
rect 12515 -3005 12525 -2985
rect 12485 -3020 12525 -3005
rect 12895 -3030 12935 -3015
rect 12895 -3050 12905 -3030
rect 12925 -3050 12935 -3030
rect 12895 -3075 12935 -3050
rect 12895 -3095 12905 -3075
rect 12925 -3095 12935 -3075
rect 12895 -3120 12935 -3095
rect 12895 -3140 12905 -3120
rect 12925 -3140 12935 -3120
rect 12895 -3170 12935 -3140
rect 12895 -3190 12905 -3170
rect 12925 -3190 12935 -3170
rect 12895 -3215 12935 -3190
rect 12895 -3235 12905 -3215
rect 12925 -3235 12935 -3215
rect 12895 -3260 12935 -3235
rect 12895 -3280 12905 -3260
rect 12925 -3280 12935 -3260
rect 12895 -3295 12935 -3280
rect 12995 -3030 13035 -3015
rect 12995 -3050 13005 -3030
rect 13025 -3050 13035 -3030
rect 12995 -3075 13035 -3050
rect 12995 -3095 13005 -3075
rect 13025 -3095 13035 -3075
rect 12995 -3120 13035 -3095
rect 12995 -3140 13005 -3120
rect 13025 -3140 13035 -3120
rect 12995 -3170 13035 -3140
rect 12995 -3190 13005 -3170
rect 13025 -3190 13035 -3170
rect 12995 -3215 13035 -3190
rect 12995 -3235 13005 -3215
rect 13025 -3235 13035 -3215
rect 12995 -3260 13035 -3235
rect 12995 -3280 13005 -3260
rect 13025 -3280 13035 -3260
rect 12995 -3295 13035 -3280
rect 13095 -3030 13135 -3015
rect 13095 -3050 13105 -3030
rect 13125 -3050 13135 -3030
rect 13095 -3075 13135 -3050
rect 13095 -3095 13105 -3075
rect 13125 -3095 13135 -3075
rect 13095 -3120 13135 -3095
rect 13095 -3140 13105 -3120
rect 13125 -3140 13135 -3120
rect 13095 -3170 13135 -3140
rect 13095 -3190 13105 -3170
rect 13125 -3190 13135 -3170
rect 13095 -3215 13135 -3190
rect 13095 -3235 13105 -3215
rect 13125 -3235 13135 -3215
rect 13095 -3260 13135 -3235
rect 13095 -3280 13105 -3260
rect 13125 -3280 13135 -3260
rect 13095 -3295 13135 -3280
rect 13195 -3030 13235 -3015
rect 13195 -3050 13205 -3030
rect 13225 -3050 13235 -3030
rect 13195 -3075 13235 -3050
rect 13195 -3095 13205 -3075
rect 13225 -3095 13235 -3075
rect 13195 -3120 13235 -3095
rect 13195 -3140 13205 -3120
rect 13225 -3140 13235 -3120
rect 13195 -3170 13235 -3140
rect 13195 -3190 13205 -3170
rect 13225 -3190 13235 -3170
rect 13195 -3215 13235 -3190
rect 13195 -3235 13205 -3215
rect 13225 -3235 13235 -3215
rect 13195 -3260 13235 -3235
rect 13195 -3280 13205 -3260
rect 13225 -3280 13235 -3260
rect 13195 -3295 13235 -3280
rect 13295 -3030 13335 -3015
rect 13295 -3050 13305 -3030
rect 13325 -3050 13335 -3030
rect 13295 -3075 13335 -3050
rect 13295 -3095 13305 -3075
rect 13325 -3095 13335 -3075
rect 13295 -3120 13335 -3095
rect 13295 -3140 13305 -3120
rect 13325 -3140 13335 -3120
rect 13295 -3170 13335 -3140
rect 13295 -3190 13305 -3170
rect 13325 -3190 13335 -3170
rect 13295 -3215 13335 -3190
rect 13295 -3235 13305 -3215
rect 13325 -3235 13335 -3215
rect 13295 -3260 13335 -3235
rect 13295 -3280 13305 -3260
rect 13325 -3280 13335 -3260
rect 13295 -3295 13335 -3280
rect 13395 -3030 13435 -3015
rect 13395 -3050 13405 -3030
rect 13425 -3050 13435 -3030
rect 13395 -3075 13435 -3050
rect 13395 -3095 13405 -3075
rect 13425 -3095 13435 -3075
rect 13395 -3120 13435 -3095
rect 13395 -3140 13405 -3120
rect 13425 -3140 13435 -3120
rect 13395 -3170 13435 -3140
rect 13395 -3190 13405 -3170
rect 13425 -3190 13435 -3170
rect 13395 -3215 13435 -3190
rect 13395 -3235 13405 -3215
rect 13425 -3235 13435 -3215
rect 13395 -3260 13435 -3235
rect 13395 -3280 13405 -3260
rect 13425 -3280 13435 -3260
rect 13395 -3295 13435 -3280
rect 13495 -3030 13535 -3015
rect 13495 -3050 13505 -3030
rect 13525 -3050 13535 -3030
rect 13495 -3075 13535 -3050
rect 13495 -3095 13505 -3075
rect 13525 -3095 13535 -3075
rect 13495 -3120 13535 -3095
rect 13495 -3140 13505 -3120
rect 13525 -3140 13535 -3120
rect 13495 -3170 13535 -3140
rect 13495 -3190 13505 -3170
rect 13525 -3190 13535 -3170
rect 13495 -3215 13535 -3190
rect 13495 -3235 13505 -3215
rect 13525 -3235 13535 -3215
rect 13495 -3260 13535 -3235
rect 13495 -3280 13505 -3260
rect 13525 -3280 13535 -3260
rect 13495 -3295 13535 -3280
rect 13595 -3030 13635 -3015
rect 13595 -3050 13605 -3030
rect 13625 -3050 13635 -3030
rect 13595 -3075 13635 -3050
rect 13595 -3095 13605 -3075
rect 13625 -3095 13635 -3075
rect 13595 -3120 13635 -3095
rect 13595 -3140 13605 -3120
rect 13625 -3140 13635 -3120
rect 13595 -3170 13635 -3140
rect 13595 -3190 13605 -3170
rect 13625 -3190 13635 -3170
rect 13595 -3215 13635 -3190
rect 13595 -3235 13605 -3215
rect 13625 -3235 13635 -3215
rect 13595 -3260 13635 -3235
rect 13595 -3280 13605 -3260
rect 13625 -3280 13635 -3260
rect 13595 -3295 13635 -3280
rect 13695 -3030 13735 -3015
rect 13695 -3050 13705 -3030
rect 13725 -3050 13735 -3030
rect 13695 -3075 13735 -3050
rect 13695 -3095 13705 -3075
rect 13725 -3095 13735 -3075
rect 13695 -3120 13735 -3095
rect 13695 -3140 13705 -3120
rect 13725 -3140 13735 -3120
rect 13695 -3170 13735 -3140
rect 13695 -3190 13705 -3170
rect 13725 -3190 13735 -3170
rect 13695 -3215 13735 -3190
rect 13695 -3235 13705 -3215
rect 13725 -3235 13735 -3215
rect 13695 -3260 13735 -3235
rect 13695 -3280 13705 -3260
rect 13725 -3280 13735 -3260
rect 13695 -3295 13735 -3280
rect 13795 -3030 13835 -3015
rect 13795 -3050 13805 -3030
rect 13825 -3050 13835 -3030
rect 13795 -3075 13835 -3050
rect 13795 -3095 13805 -3075
rect 13825 -3095 13835 -3075
rect 13795 -3120 13835 -3095
rect 13795 -3140 13805 -3120
rect 13825 -3140 13835 -3120
rect 13795 -3170 13835 -3140
rect 13795 -3190 13805 -3170
rect 13825 -3190 13835 -3170
rect 13795 -3215 13835 -3190
rect 13795 -3235 13805 -3215
rect 13825 -3235 13835 -3215
rect 13795 -3260 13835 -3235
rect 13795 -3280 13805 -3260
rect 13825 -3280 13835 -3260
rect 13795 -3295 13835 -3280
rect 13895 -3030 13935 -3015
rect 13895 -3050 13905 -3030
rect 13925 -3050 13935 -3030
rect 13895 -3075 13935 -3050
rect 13895 -3095 13905 -3075
rect 13925 -3095 13935 -3075
rect 13895 -3120 13935 -3095
rect 13895 -3140 13905 -3120
rect 13925 -3140 13935 -3120
rect 13895 -3170 13935 -3140
rect 13895 -3190 13905 -3170
rect 13925 -3190 13935 -3170
rect 13895 -3215 13935 -3190
rect 13895 -3235 13905 -3215
rect 13925 -3235 13935 -3215
rect 13895 -3260 13935 -3235
rect 13895 -3280 13905 -3260
rect 13925 -3280 13935 -3260
rect 13895 -3295 13935 -3280
rect 13995 -3030 14035 -3015
rect 13995 -3050 14005 -3030
rect 14025 -3050 14035 -3030
rect 13995 -3075 14035 -3050
rect 13995 -3095 14005 -3075
rect 14025 -3095 14035 -3075
rect 13995 -3120 14035 -3095
rect 13995 -3140 14005 -3120
rect 14025 -3140 14035 -3120
rect 13995 -3170 14035 -3140
rect 13995 -3190 14005 -3170
rect 14025 -3190 14035 -3170
rect 13995 -3215 14035 -3190
rect 13995 -3235 14005 -3215
rect 14025 -3235 14035 -3215
rect 13995 -3260 14035 -3235
rect 13995 -3280 14005 -3260
rect 14025 -3280 14035 -3260
rect 13995 -3295 14035 -3280
rect 14095 -3030 14135 -3015
rect 14095 -3050 14105 -3030
rect 14125 -3050 14135 -3030
rect 14095 -3075 14135 -3050
rect 14095 -3095 14105 -3075
rect 14125 -3095 14135 -3075
rect 14095 -3120 14135 -3095
rect 14095 -3140 14105 -3120
rect 14125 -3140 14135 -3120
rect 14095 -3170 14135 -3140
rect 14095 -3190 14105 -3170
rect 14125 -3190 14135 -3170
rect 14095 -3215 14135 -3190
rect 14095 -3235 14105 -3215
rect 14125 -3235 14135 -3215
rect 14095 -3260 14135 -3235
rect 14095 -3280 14105 -3260
rect 14125 -3280 14135 -3260
rect 14095 -3295 14135 -3280
rect 11030 -3350 11070 -3335
rect 11030 -3370 11040 -3350
rect 11060 -3370 11070 -3350
rect 11030 -3400 11070 -3370
rect 11030 -3420 11040 -3400
rect 11060 -3420 11070 -3400
rect 11030 -3450 11070 -3420
rect 11030 -3470 11040 -3450
rect 11060 -3470 11070 -3450
rect 11030 -3485 11070 -3470
rect 11085 -3350 11125 -3335
rect 11085 -3370 11095 -3350
rect 11115 -3370 11125 -3350
rect 11085 -3400 11125 -3370
rect 11085 -3420 11095 -3400
rect 11115 -3420 11125 -3400
rect 11085 -3450 11125 -3420
rect 11085 -3470 11095 -3450
rect 11115 -3470 11125 -3450
rect 11085 -3485 11125 -3470
rect 11140 -3350 11180 -3335
rect 11140 -3370 11150 -3350
rect 11170 -3370 11180 -3350
rect 11140 -3400 11180 -3370
rect 11140 -3420 11150 -3400
rect 11170 -3420 11180 -3400
rect 11140 -3450 11180 -3420
rect 11140 -3470 11150 -3450
rect 11170 -3470 11180 -3450
rect 11140 -3485 11180 -3470
rect 11195 -3350 11235 -3335
rect 11195 -3370 11205 -3350
rect 11225 -3370 11235 -3350
rect 11195 -3400 11235 -3370
rect 11195 -3420 11205 -3400
rect 11225 -3420 11235 -3400
rect 11195 -3450 11235 -3420
rect 11195 -3470 11205 -3450
rect 11225 -3470 11235 -3450
rect 11195 -3485 11235 -3470
rect 11250 -3350 11290 -3335
rect 11250 -3370 11260 -3350
rect 11280 -3370 11290 -3350
rect 11250 -3400 11290 -3370
rect 11250 -3420 11260 -3400
rect 11280 -3420 11290 -3400
rect 11250 -3450 11290 -3420
rect 11250 -3470 11260 -3450
rect 11280 -3470 11290 -3450
rect 11250 -3485 11290 -3470
rect 11305 -3350 11345 -3335
rect 11305 -3370 11315 -3350
rect 11335 -3370 11345 -3350
rect 11305 -3400 11345 -3370
rect 11305 -3420 11315 -3400
rect 11335 -3420 11345 -3400
rect 11305 -3450 11345 -3420
rect 11305 -3470 11315 -3450
rect 11335 -3470 11345 -3450
rect 11305 -3485 11345 -3470
rect 11360 -3350 11400 -3335
rect 11360 -3370 11370 -3350
rect 11390 -3370 11400 -3350
rect 11360 -3400 11400 -3370
rect 11360 -3420 11370 -3400
rect 11390 -3420 11400 -3400
rect 11360 -3450 11400 -3420
rect 11360 -3470 11370 -3450
rect 11390 -3470 11400 -3450
rect 11360 -3485 11400 -3470
rect 11415 -3350 11455 -3335
rect 11415 -3370 11425 -3350
rect 11445 -3370 11455 -3350
rect 11415 -3400 11455 -3370
rect 11415 -3420 11425 -3400
rect 11445 -3420 11455 -3400
rect 11415 -3450 11455 -3420
rect 11415 -3470 11425 -3450
rect 11445 -3470 11455 -3450
rect 11415 -3485 11455 -3470
rect 11470 -3350 11510 -3335
rect 11470 -3370 11480 -3350
rect 11500 -3370 11510 -3350
rect 11470 -3400 11510 -3370
rect 11470 -3420 11480 -3400
rect 11500 -3420 11510 -3400
rect 11470 -3450 11510 -3420
rect 11470 -3470 11480 -3450
rect 11500 -3470 11510 -3450
rect 11470 -3485 11510 -3470
rect 11525 -3350 11565 -3335
rect 11525 -3370 11535 -3350
rect 11555 -3370 11565 -3350
rect 11525 -3400 11565 -3370
rect 11525 -3420 11535 -3400
rect 11555 -3420 11565 -3400
rect 11525 -3450 11565 -3420
rect 11525 -3470 11535 -3450
rect 11555 -3470 11565 -3450
rect 11525 -3485 11565 -3470
rect 11580 -3350 11620 -3335
rect 11580 -3370 11590 -3350
rect 11610 -3370 11620 -3350
rect 11580 -3400 11620 -3370
rect 11580 -3420 11590 -3400
rect 11610 -3420 11620 -3400
rect 11580 -3450 11620 -3420
rect 11580 -3470 11590 -3450
rect 11610 -3470 11620 -3450
rect 11580 -3485 11620 -3470
rect 11635 -3350 11675 -3335
rect 11635 -3370 11645 -3350
rect 11665 -3370 11675 -3350
rect 11635 -3400 11675 -3370
rect 11635 -3420 11645 -3400
rect 11665 -3420 11675 -3400
rect 11635 -3450 11675 -3420
rect 11635 -3470 11645 -3450
rect 11665 -3470 11675 -3450
rect 11635 -3485 11675 -3470
rect 11690 -3350 11730 -3335
rect 11770 -3350 11810 -3335
rect 11690 -3370 11700 -3350
rect 11720 -3370 11730 -3350
rect 11770 -3370 11780 -3350
rect 11800 -3370 11810 -3350
rect 11690 -3400 11730 -3370
rect 11770 -3400 11810 -3370
rect 11690 -3420 11700 -3400
rect 11720 -3420 11730 -3400
rect 11770 -3420 11780 -3400
rect 11800 -3420 11810 -3400
rect 11690 -3450 11730 -3420
rect 11770 -3450 11810 -3420
rect 11690 -3470 11700 -3450
rect 11720 -3470 11730 -3450
rect 11770 -3470 11780 -3450
rect 11800 -3470 11810 -3450
rect 11690 -3485 11730 -3470
rect 11770 -3485 11810 -3470
rect 11825 -3350 11865 -3335
rect 11825 -3370 11835 -3350
rect 11855 -3370 11865 -3350
rect 11825 -3400 11865 -3370
rect 11825 -3420 11835 -3400
rect 11855 -3420 11865 -3400
rect 11825 -3450 11865 -3420
rect 11825 -3470 11835 -3450
rect 11855 -3470 11865 -3450
rect 11825 -3485 11865 -3470
rect 11880 -3350 11920 -3335
rect 11880 -3370 11890 -3350
rect 11910 -3370 11920 -3350
rect 11880 -3400 11920 -3370
rect 11880 -3420 11890 -3400
rect 11910 -3420 11920 -3400
rect 11880 -3450 11920 -3420
rect 11880 -3470 11890 -3450
rect 11910 -3470 11920 -3450
rect 11880 -3485 11920 -3470
rect 11935 -3350 11975 -3335
rect 11935 -3370 11945 -3350
rect 11965 -3370 11975 -3350
rect 11935 -3400 11975 -3370
rect 11935 -3420 11945 -3400
rect 11965 -3420 11975 -3400
rect 11935 -3450 11975 -3420
rect 11935 -3470 11945 -3450
rect 11965 -3470 11975 -3450
rect 11935 -3485 11975 -3470
rect 11990 -3350 12030 -3335
rect 12070 -3350 12110 -3335
rect 11990 -3370 12000 -3350
rect 12020 -3370 12030 -3350
rect 12070 -3370 12080 -3350
rect 12100 -3370 12110 -3350
rect 11990 -3400 12030 -3370
rect 12070 -3400 12110 -3370
rect 11990 -3420 12000 -3400
rect 12020 -3420 12030 -3400
rect 12070 -3420 12080 -3400
rect 12100 -3420 12110 -3400
rect 11990 -3450 12030 -3420
rect 12070 -3450 12110 -3420
rect 11990 -3470 12000 -3450
rect 12020 -3470 12030 -3450
rect 12070 -3470 12080 -3450
rect 12100 -3470 12110 -3450
rect 11990 -3485 12030 -3470
rect 12070 -3485 12110 -3470
rect 12125 -3350 12165 -3335
rect 12125 -3370 12135 -3350
rect 12155 -3370 12165 -3350
rect 12125 -3400 12165 -3370
rect 12125 -3420 12135 -3400
rect 12155 -3420 12165 -3400
rect 12125 -3450 12165 -3420
rect 12125 -3470 12135 -3450
rect 12155 -3470 12165 -3450
rect 12125 -3485 12165 -3470
rect 12180 -3350 12220 -3335
rect 12180 -3370 12190 -3350
rect 12210 -3370 12220 -3350
rect 12180 -3400 12220 -3370
rect 12180 -3420 12190 -3400
rect 12210 -3420 12220 -3400
rect 12180 -3450 12220 -3420
rect 12180 -3470 12190 -3450
rect 12210 -3470 12220 -3450
rect 12180 -3485 12220 -3470
rect 12235 -3350 12275 -3335
rect 12235 -3370 12245 -3350
rect 12265 -3370 12275 -3350
rect 12235 -3400 12275 -3370
rect 12235 -3420 12245 -3400
rect 12265 -3420 12275 -3400
rect 12235 -3450 12275 -3420
rect 12235 -3470 12245 -3450
rect 12265 -3470 12275 -3450
rect 12235 -3485 12275 -3470
rect 12290 -3350 12330 -3335
rect 12290 -3370 12300 -3350
rect 12320 -3370 12330 -3350
rect 12290 -3400 12330 -3370
rect 12290 -3420 12300 -3400
rect 12320 -3420 12330 -3400
rect 12290 -3450 12330 -3420
rect 12290 -3470 12300 -3450
rect 12320 -3470 12330 -3450
rect 12290 -3485 12330 -3470
rect 12345 -3350 12385 -3335
rect 12345 -3370 12355 -3350
rect 12375 -3370 12385 -3350
rect 12345 -3400 12385 -3370
rect 12345 -3420 12355 -3400
rect 12375 -3420 12385 -3400
rect 12345 -3450 12385 -3420
rect 12345 -3470 12355 -3450
rect 12375 -3470 12385 -3450
rect 12345 -3485 12385 -3470
rect 12400 -3350 12440 -3335
rect 12400 -3370 12410 -3350
rect 12430 -3370 12440 -3350
rect 12400 -3400 12440 -3370
rect 12400 -3420 12410 -3400
rect 12430 -3420 12440 -3400
rect 12400 -3450 12440 -3420
rect 12400 -3470 12410 -3450
rect 12430 -3470 12440 -3450
rect 12400 -3485 12440 -3470
rect 12455 -3350 12495 -3335
rect 12455 -3370 12465 -3350
rect 12485 -3370 12495 -3350
rect 12455 -3400 12495 -3370
rect 12455 -3420 12465 -3400
rect 12485 -3420 12495 -3400
rect 12455 -3450 12495 -3420
rect 12455 -3470 12465 -3450
rect 12485 -3470 12495 -3450
rect 12455 -3485 12495 -3470
rect 12510 -3350 12550 -3335
rect 12510 -3370 12520 -3350
rect 12540 -3370 12550 -3350
rect 12510 -3400 12550 -3370
rect 12510 -3420 12520 -3400
rect 12540 -3420 12550 -3400
rect 12510 -3450 12550 -3420
rect 12510 -3470 12520 -3450
rect 12540 -3470 12550 -3450
rect 12510 -3485 12550 -3470
rect 12565 -3350 12605 -3335
rect 12565 -3370 12575 -3350
rect 12595 -3370 12605 -3350
rect 12565 -3400 12605 -3370
rect 12565 -3420 12575 -3400
rect 12595 -3420 12605 -3400
rect 12565 -3450 12605 -3420
rect 12565 -3470 12575 -3450
rect 12595 -3470 12605 -3450
rect 12565 -3485 12605 -3470
rect 12620 -3350 12660 -3335
rect 12620 -3370 12630 -3350
rect 12650 -3370 12660 -3350
rect 12620 -3400 12660 -3370
rect 12620 -3420 12630 -3400
rect 12650 -3420 12660 -3400
rect 12620 -3450 12660 -3420
rect 12620 -3470 12630 -3450
rect 12650 -3470 12660 -3450
rect 12620 -3485 12660 -3470
rect 12675 -3350 12715 -3335
rect 12675 -3370 12685 -3350
rect 12705 -3370 12715 -3350
rect 12675 -3400 12715 -3370
rect 12675 -3420 12685 -3400
rect 12705 -3420 12715 -3400
rect 12675 -3450 12715 -3420
rect 12675 -3470 12685 -3450
rect 12705 -3470 12715 -3450
rect 12675 -3485 12715 -3470
rect 12730 -3350 12770 -3335
rect 12730 -3370 12740 -3350
rect 12760 -3370 12770 -3350
rect 12730 -3400 12770 -3370
rect 12730 -3420 12740 -3400
rect 12760 -3420 12770 -3400
rect 12730 -3450 12770 -3420
rect 12730 -3470 12740 -3450
rect 12760 -3470 12770 -3450
rect 12730 -3485 12770 -3470
rect 11205 -3830 11245 -3815
rect 11205 -3850 11215 -3830
rect 11235 -3850 11245 -3830
rect 11205 -3880 11245 -3850
rect 11205 -3900 11215 -3880
rect 11235 -3900 11245 -3880
rect 11205 -3930 11245 -3900
rect 11205 -3950 11215 -3930
rect 11235 -3950 11245 -3930
rect 11205 -3980 11245 -3950
rect 11205 -4000 11215 -3980
rect 11235 -4000 11245 -3980
rect 11205 -4030 11245 -4000
rect 11205 -4050 11215 -4030
rect 11235 -4050 11245 -4030
rect 11205 -4065 11245 -4050
rect 11260 -3830 11300 -3815
rect 11260 -3850 11270 -3830
rect 11290 -3850 11300 -3830
rect 11260 -3880 11300 -3850
rect 11260 -3900 11270 -3880
rect 11290 -3900 11300 -3880
rect 11260 -3930 11300 -3900
rect 11260 -3950 11270 -3930
rect 11290 -3950 11300 -3930
rect 11260 -3980 11300 -3950
rect 11260 -4000 11270 -3980
rect 11290 -4000 11300 -3980
rect 11260 -4030 11300 -4000
rect 11260 -4050 11270 -4030
rect 11290 -4050 11300 -4030
rect 11260 -4065 11300 -4050
rect 11315 -3830 11355 -3815
rect 11315 -3850 11325 -3830
rect 11345 -3850 11355 -3830
rect 11315 -3880 11355 -3850
rect 11315 -3900 11325 -3880
rect 11345 -3900 11355 -3880
rect 11315 -3930 11355 -3900
rect 11315 -3950 11325 -3930
rect 11345 -3950 11355 -3930
rect 11315 -3980 11355 -3950
rect 11315 -4000 11325 -3980
rect 11345 -4000 11355 -3980
rect 11315 -4030 11355 -4000
rect 11315 -4050 11325 -4030
rect 11345 -4050 11355 -4030
rect 11315 -4065 11355 -4050
rect 11370 -3830 11410 -3815
rect 11370 -3850 11380 -3830
rect 11400 -3850 11410 -3830
rect 11370 -3880 11410 -3850
rect 11370 -3900 11380 -3880
rect 11400 -3900 11410 -3880
rect 11370 -3930 11410 -3900
rect 11370 -3950 11380 -3930
rect 11400 -3950 11410 -3930
rect 11370 -3980 11410 -3950
rect 11370 -4000 11380 -3980
rect 11400 -4000 11410 -3980
rect 11370 -4030 11410 -4000
rect 11370 -4050 11380 -4030
rect 11400 -4050 11410 -4030
rect 11370 -4065 11410 -4050
rect 11425 -3830 11465 -3815
rect 11425 -3850 11435 -3830
rect 11455 -3850 11465 -3830
rect 11425 -3880 11465 -3850
rect 11425 -3900 11435 -3880
rect 11455 -3900 11465 -3880
rect 11425 -3930 11465 -3900
rect 11425 -3950 11435 -3930
rect 11455 -3950 11465 -3930
rect 11425 -3980 11465 -3950
rect 11425 -4000 11435 -3980
rect 11455 -4000 11465 -3980
rect 11425 -4030 11465 -4000
rect 11425 -4050 11435 -4030
rect 11455 -4050 11465 -4030
rect 11425 -4065 11465 -4050
rect 11480 -3830 11520 -3815
rect 11480 -3850 11490 -3830
rect 11510 -3850 11520 -3830
rect 11480 -3880 11520 -3850
rect 11480 -3900 11490 -3880
rect 11510 -3900 11520 -3880
rect 11480 -3930 11520 -3900
rect 11480 -3950 11490 -3930
rect 11510 -3950 11520 -3930
rect 11480 -3980 11520 -3950
rect 11480 -4000 11490 -3980
rect 11510 -4000 11520 -3980
rect 11480 -4030 11520 -4000
rect 11480 -4050 11490 -4030
rect 11510 -4050 11520 -4030
rect 11480 -4065 11520 -4050
rect 11535 -3830 11575 -3815
rect 11535 -3850 11545 -3830
rect 11565 -3850 11575 -3830
rect 11535 -3880 11575 -3850
rect 11535 -3900 11545 -3880
rect 11565 -3900 11575 -3880
rect 11535 -3930 11575 -3900
rect 11535 -3950 11545 -3930
rect 11565 -3950 11575 -3930
rect 11535 -3980 11575 -3950
rect 11535 -4000 11545 -3980
rect 11565 -4000 11575 -3980
rect 11535 -4030 11575 -4000
rect 11535 -4050 11545 -4030
rect 11565 -4050 11575 -4030
rect 11535 -4065 11575 -4050
rect 11590 -3830 11630 -3815
rect 11590 -3850 11600 -3830
rect 11620 -3850 11630 -3830
rect 11590 -3880 11630 -3850
rect 11590 -3900 11600 -3880
rect 11620 -3900 11630 -3880
rect 11590 -3930 11630 -3900
rect 11590 -3950 11600 -3930
rect 11620 -3950 11630 -3930
rect 11590 -3980 11630 -3950
rect 11590 -4000 11600 -3980
rect 11620 -4000 11630 -3980
rect 11590 -4030 11630 -4000
rect 11590 -4050 11600 -4030
rect 11620 -4050 11630 -4030
rect 11590 -4065 11630 -4050
rect 11645 -3830 11685 -3815
rect 11645 -3850 11655 -3830
rect 11675 -3850 11685 -3830
rect 11645 -3880 11685 -3850
rect 11645 -3900 11655 -3880
rect 11675 -3900 11685 -3880
rect 11645 -3930 11685 -3900
rect 11645 -3950 11655 -3930
rect 11675 -3950 11685 -3930
rect 11645 -3980 11685 -3950
rect 11645 -4000 11655 -3980
rect 11675 -4000 11685 -3980
rect 11645 -4030 11685 -4000
rect 11645 -4050 11655 -4030
rect 11675 -4050 11685 -4030
rect 11645 -4065 11685 -4050
rect 11700 -3830 11740 -3815
rect 11700 -3850 11710 -3830
rect 11730 -3850 11740 -3830
rect 11700 -3880 11740 -3850
rect 11700 -3900 11710 -3880
rect 11730 -3900 11740 -3880
rect 11700 -3930 11740 -3900
rect 11700 -3950 11710 -3930
rect 11730 -3950 11740 -3930
rect 11700 -3980 11740 -3950
rect 11700 -4000 11710 -3980
rect 11730 -4000 11740 -3980
rect 11700 -4030 11740 -4000
rect 11700 -4050 11710 -4030
rect 11730 -4050 11740 -4030
rect 11700 -4065 11740 -4050
rect 11755 -3830 11795 -3815
rect 11755 -3850 11765 -3830
rect 11785 -3850 11795 -3830
rect 11755 -3880 11795 -3850
rect 11755 -3900 11765 -3880
rect 11785 -3900 11795 -3880
rect 11755 -3930 11795 -3900
rect 11755 -3950 11765 -3930
rect 11785 -3950 11795 -3930
rect 11755 -3980 11795 -3950
rect 11755 -4000 11765 -3980
rect 11785 -4000 11795 -3980
rect 11755 -4030 11795 -4000
rect 11755 -4050 11765 -4030
rect 11785 -4050 11795 -4030
rect 11755 -4065 11795 -4050
rect 11810 -3830 11850 -3815
rect 11810 -3850 11820 -3830
rect 11840 -3850 11850 -3830
rect 11810 -3880 11850 -3850
rect 11810 -3900 11820 -3880
rect 11840 -3900 11850 -3880
rect 11810 -3930 11850 -3900
rect 11810 -3950 11820 -3930
rect 11840 -3950 11850 -3930
rect 11810 -3980 11850 -3950
rect 11810 -4000 11820 -3980
rect 11840 -4000 11850 -3980
rect 11810 -4030 11850 -4000
rect 11810 -4050 11820 -4030
rect 11840 -4050 11850 -4030
rect 11810 -4065 11850 -4050
rect 11865 -3830 11905 -3815
rect 11865 -3850 11875 -3830
rect 11895 -3850 11905 -3830
rect 11865 -3880 11905 -3850
rect 11865 -3900 11875 -3880
rect 11895 -3900 11905 -3880
rect 11865 -3930 11905 -3900
rect 11865 -3950 11875 -3930
rect 11895 -3950 11905 -3930
rect 11865 -3980 11905 -3950
rect 11865 -4000 11875 -3980
rect 11895 -4000 11905 -3980
rect 11865 -4030 11905 -4000
rect 11865 -4050 11875 -4030
rect 11895 -4050 11905 -4030
rect 11865 -4065 11905 -4050
rect 11920 -3830 11960 -3815
rect 11920 -3850 11930 -3830
rect 11950 -3850 11960 -3830
rect 11920 -3880 11960 -3850
rect 11920 -3900 11930 -3880
rect 11950 -3900 11960 -3880
rect 11920 -3930 11960 -3900
rect 11920 -3950 11930 -3930
rect 11950 -3950 11960 -3930
rect 11920 -3980 11960 -3950
rect 11920 -4000 11930 -3980
rect 11950 -4000 11960 -3980
rect 11920 -4030 11960 -4000
rect 11920 -4050 11930 -4030
rect 11950 -4050 11960 -4030
rect 11920 -4065 11960 -4050
rect 11975 -3830 12015 -3815
rect 11975 -3850 11985 -3830
rect 12005 -3850 12015 -3830
rect 11975 -3880 12015 -3850
rect 11975 -3900 11985 -3880
rect 12005 -3900 12015 -3880
rect 11975 -3930 12015 -3900
rect 11975 -3950 11985 -3930
rect 12005 -3950 12015 -3930
rect 11975 -3980 12015 -3950
rect 11975 -4000 11985 -3980
rect 12005 -4000 12015 -3980
rect 11975 -4030 12015 -4000
rect 11975 -4050 11985 -4030
rect 12005 -4050 12015 -4030
rect 11975 -4065 12015 -4050
rect 12030 -3830 12070 -3815
rect 12030 -3850 12040 -3830
rect 12060 -3850 12070 -3830
rect 12030 -3880 12070 -3850
rect 12030 -3900 12040 -3880
rect 12060 -3900 12070 -3880
rect 12030 -3930 12070 -3900
rect 12030 -3950 12040 -3930
rect 12060 -3950 12070 -3930
rect 12030 -3980 12070 -3950
rect 12030 -4000 12040 -3980
rect 12060 -4000 12070 -3980
rect 12030 -4030 12070 -4000
rect 12030 -4050 12040 -4030
rect 12060 -4050 12070 -4030
rect 12030 -4065 12070 -4050
rect 12085 -3830 12125 -3815
rect 12085 -3850 12095 -3830
rect 12115 -3850 12125 -3830
rect 12085 -3880 12125 -3850
rect 12085 -3900 12095 -3880
rect 12115 -3900 12125 -3880
rect 12085 -3930 12125 -3900
rect 12085 -3950 12095 -3930
rect 12115 -3950 12125 -3930
rect 12085 -3980 12125 -3950
rect 12085 -4000 12095 -3980
rect 12115 -4000 12125 -3980
rect 12085 -4030 12125 -4000
rect 12085 -4050 12095 -4030
rect 12115 -4050 12125 -4030
rect 12085 -4065 12125 -4050
rect 12140 -3830 12180 -3815
rect 12140 -3850 12150 -3830
rect 12170 -3850 12180 -3830
rect 12140 -3880 12180 -3850
rect 12140 -3900 12150 -3880
rect 12170 -3900 12180 -3880
rect 12140 -3930 12180 -3900
rect 12140 -3950 12150 -3930
rect 12170 -3950 12180 -3930
rect 12140 -3980 12180 -3950
rect 12140 -4000 12150 -3980
rect 12170 -4000 12180 -3980
rect 12140 -4030 12180 -4000
rect 12140 -4050 12150 -4030
rect 12170 -4050 12180 -4030
rect 12140 -4065 12180 -4050
rect 12195 -3830 12235 -3815
rect 12195 -3850 12205 -3830
rect 12225 -3850 12235 -3830
rect 12195 -3880 12235 -3850
rect 12195 -3900 12205 -3880
rect 12225 -3900 12235 -3880
rect 12195 -3930 12235 -3900
rect 12195 -3950 12205 -3930
rect 12225 -3950 12235 -3930
rect 12195 -3980 12235 -3950
rect 12195 -4000 12205 -3980
rect 12225 -4000 12235 -3980
rect 12195 -4030 12235 -4000
rect 12195 -4050 12205 -4030
rect 12225 -4050 12235 -4030
rect 12195 -4065 12235 -4050
rect 12250 -3830 12290 -3815
rect 12250 -3850 12260 -3830
rect 12280 -3850 12290 -3830
rect 12250 -3880 12290 -3850
rect 12250 -3900 12260 -3880
rect 12280 -3900 12290 -3880
rect 12250 -3930 12290 -3900
rect 12250 -3950 12260 -3930
rect 12280 -3950 12290 -3930
rect 12250 -3980 12290 -3950
rect 12250 -4000 12260 -3980
rect 12280 -4000 12290 -3980
rect 12250 -4030 12290 -4000
rect 12250 -4050 12260 -4030
rect 12280 -4050 12290 -4030
rect 12250 -4065 12290 -4050
rect 12305 -3830 12345 -3815
rect 12305 -3850 12315 -3830
rect 12335 -3850 12345 -3830
rect 12305 -3880 12345 -3850
rect 12305 -3900 12315 -3880
rect 12335 -3900 12345 -3880
rect 12305 -3930 12345 -3900
rect 12305 -3950 12315 -3930
rect 12335 -3950 12345 -3930
rect 12305 -3980 12345 -3950
rect 12305 -4000 12315 -3980
rect 12335 -4000 12345 -3980
rect 12305 -4030 12345 -4000
rect 12305 -4050 12315 -4030
rect 12335 -4050 12345 -4030
rect 12305 -4065 12345 -4050
rect 12360 -3830 12400 -3815
rect 12360 -3850 12370 -3830
rect 12390 -3850 12400 -3830
rect 12360 -3880 12400 -3850
rect 12360 -3900 12370 -3880
rect 12390 -3900 12400 -3880
rect 12360 -3930 12400 -3900
rect 12360 -3950 12370 -3930
rect 12390 -3950 12400 -3930
rect 12360 -3980 12400 -3950
rect 12360 -4000 12370 -3980
rect 12390 -4000 12400 -3980
rect 12360 -4030 12400 -4000
rect 12360 -4050 12370 -4030
rect 12390 -4050 12400 -4030
rect 12360 -4065 12400 -4050
rect 12415 -3830 12455 -3815
rect 12415 -3850 12425 -3830
rect 12445 -3850 12455 -3830
rect 12415 -3880 12455 -3850
rect 12415 -3900 12425 -3880
rect 12445 -3900 12455 -3880
rect 12415 -3930 12455 -3900
rect 12415 -3950 12425 -3930
rect 12445 -3950 12455 -3930
rect 12415 -3980 12455 -3950
rect 12415 -4000 12425 -3980
rect 12445 -4000 12455 -3980
rect 12415 -4030 12455 -4000
rect 12415 -4050 12425 -4030
rect 12445 -4050 12455 -4030
rect 12415 -4065 12455 -4050
rect 12470 -3830 12510 -3815
rect 12470 -3850 12480 -3830
rect 12500 -3850 12510 -3830
rect 12470 -3880 12510 -3850
rect 12470 -3900 12480 -3880
rect 12500 -3900 12510 -3880
rect 12470 -3930 12510 -3900
rect 12470 -3950 12480 -3930
rect 12500 -3950 12510 -3930
rect 12470 -3980 12510 -3950
rect 12470 -4000 12480 -3980
rect 12500 -4000 12510 -3980
rect 12470 -4030 12510 -4000
rect 12470 -4050 12480 -4030
rect 12500 -4050 12510 -4030
rect 12470 -4065 12510 -4050
rect 12525 -3830 12565 -3815
rect 12525 -3850 12535 -3830
rect 12555 -3850 12565 -3830
rect 12525 -3880 12565 -3850
rect 12525 -3900 12535 -3880
rect 12555 -3900 12565 -3880
rect 12525 -3930 12565 -3900
rect 12525 -3950 12535 -3930
rect 12555 -3950 12565 -3930
rect 12525 -3980 12565 -3950
rect 12525 -4000 12535 -3980
rect 12555 -4000 12565 -3980
rect 12525 -4030 12565 -4000
rect 12525 -4050 12535 -4030
rect 12555 -4050 12565 -4030
rect 12525 -4065 12565 -4050
rect 12580 -3830 12620 -3815
rect 12580 -3850 12590 -3830
rect 12610 -3850 12620 -3830
rect 12580 -3880 12620 -3850
rect 12580 -3900 12590 -3880
rect 12610 -3900 12620 -3880
rect 12580 -3930 12620 -3900
rect 12580 -3950 12590 -3930
rect 12610 -3950 12620 -3930
rect 12580 -3980 12620 -3950
rect 12580 -4000 12590 -3980
rect 12610 -4000 12620 -3980
rect 12580 -4030 12620 -4000
rect 12580 -4050 12590 -4030
rect 12610 -4050 12620 -4030
rect 12580 -4065 12620 -4050
<< pdiff >>
rect 2995 2915 3035 2930
rect 2995 2895 3005 2915
rect 3025 2895 3035 2915
rect 2995 2865 3035 2895
rect 2995 2845 3005 2865
rect 3025 2845 3035 2865
rect 2995 2830 3035 2845
rect 3085 2915 3125 2930
rect 3085 2895 3095 2915
rect 3115 2895 3125 2915
rect 3085 2865 3125 2895
rect 3085 2845 3095 2865
rect 3115 2845 3125 2865
rect 3085 2830 3125 2845
rect 3175 2915 3215 2930
rect 3175 2895 3185 2915
rect 3205 2895 3215 2915
rect 3175 2865 3215 2895
rect 3175 2845 3185 2865
rect 3205 2845 3215 2865
rect 3175 2830 3215 2845
rect 3265 2915 3305 2930
rect 3265 2895 3275 2915
rect 3295 2895 3305 2915
rect 3265 2865 3305 2895
rect 3265 2845 3275 2865
rect 3295 2845 3305 2865
rect 3265 2830 3305 2845
rect 3355 2915 3395 2930
rect 3355 2895 3365 2915
rect 3385 2895 3395 2915
rect 3355 2865 3395 2895
rect 3355 2845 3365 2865
rect 3385 2845 3395 2865
rect 3355 2830 3395 2845
rect 3445 2915 3485 2930
rect 3445 2895 3455 2915
rect 3475 2895 3485 2915
rect 3445 2865 3485 2895
rect 3445 2845 3455 2865
rect 3475 2845 3485 2865
rect 3445 2830 3485 2845
rect 3535 2915 3575 2930
rect 3535 2895 3545 2915
rect 3565 2895 3575 2915
rect 3535 2865 3575 2895
rect 3535 2845 3545 2865
rect 3565 2845 3575 2865
rect 3535 2830 3575 2845
rect 3625 2915 3665 2930
rect 3625 2895 3635 2915
rect 3655 2895 3665 2915
rect 3625 2865 3665 2895
rect 3625 2845 3635 2865
rect 3655 2845 3665 2865
rect 3625 2830 3665 2845
rect 3715 2915 3755 2930
rect 3715 2895 3725 2915
rect 3745 2895 3755 2915
rect 3715 2865 3755 2895
rect 3715 2845 3725 2865
rect 3745 2845 3755 2865
rect 3715 2830 3755 2845
rect 3805 2915 3845 2930
rect 3805 2895 3815 2915
rect 3835 2895 3845 2915
rect 3805 2865 3845 2895
rect 3805 2845 3815 2865
rect 3835 2845 3845 2865
rect 3805 2830 3845 2845
rect 3895 2915 3935 2930
rect 3895 2895 3905 2915
rect 3925 2895 3935 2915
rect 3895 2865 3935 2895
rect 3895 2845 3905 2865
rect 3925 2845 3935 2865
rect 3895 2830 3935 2845
rect 3985 2915 4025 2930
rect 3985 2895 3995 2915
rect 4015 2895 4025 2915
rect 3985 2865 4025 2895
rect 3985 2845 3995 2865
rect 4015 2845 4025 2865
rect 3985 2830 4025 2845
rect 4075 2915 4115 2930
rect 4075 2895 4085 2915
rect 4105 2895 4115 2915
rect 4075 2865 4115 2895
rect 4075 2845 4085 2865
rect 4105 2845 4115 2865
rect 4075 2830 4115 2845
rect 4165 2915 4205 2930
rect 4165 2895 4175 2915
rect 4195 2895 4205 2915
rect 4165 2865 4205 2895
rect 4165 2845 4175 2865
rect 4195 2845 4205 2865
rect 4165 2830 4205 2845
rect 4255 2915 4295 2930
rect 4255 2895 4265 2915
rect 4285 2895 4295 2915
rect 4255 2865 4295 2895
rect 4255 2845 4265 2865
rect 4285 2845 4295 2865
rect 4255 2830 4295 2845
rect 4345 2915 4385 2930
rect 4345 2895 4355 2915
rect 4375 2895 4385 2915
rect 4345 2865 4385 2895
rect 4345 2845 4355 2865
rect 4375 2845 4385 2865
rect 4345 2830 4385 2845
rect 4435 2915 4475 2930
rect 4435 2895 4445 2915
rect 4465 2895 4475 2915
rect 4435 2865 4475 2895
rect 4435 2845 4445 2865
rect 4465 2845 4475 2865
rect 4435 2830 4475 2845
rect 4525 2915 4565 2930
rect 4525 2895 4535 2915
rect 4555 2895 4565 2915
rect 4525 2865 4565 2895
rect 4525 2845 4535 2865
rect 4555 2845 4565 2865
rect 4525 2830 4565 2845
rect 4615 2915 4655 2930
rect 4615 2895 4625 2915
rect 4645 2895 4655 2915
rect 4615 2865 4655 2895
rect 4615 2845 4625 2865
rect 4645 2845 4655 2865
rect 4615 2830 4655 2845
rect 4705 2915 4745 2930
rect 4705 2895 4715 2915
rect 4735 2895 4745 2915
rect 4705 2865 4745 2895
rect 4705 2845 4715 2865
rect 4735 2845 4745 2865
rect 4705 2830 4745 2845
rect 4795 2915 4835 2930
rect 4795 2895 4805 2915
rect 4825 2895 4835 2915
rect 4795 2865 4835 2895
rect 4795 2845 4805 2865
rect 4825 2845 4835 2865
rect 4795 2830 4835 2845
rect 4885 2915 4925 2930
rect 4885 2895 4895 2915
rect 4915 2895 4925 2915
rect 4885 2865 4925 2895
rect 4885 2845 4895 2865
rect 4915 2845 4925 2865
rect 4885 2830 4925 2845
rect 4975 2915 5015 2930
rect 4975 2895 4985 2915
rect 5005 2895 5015 2915
rect 4975 2865 5015 2895
rect 4975 2845 4985 2865
rect 5005 2845 5015 2865
rect 4975 2830 5015 2845
rect 3175 2685 3215 2700
rect 3175 2665 3185 2685
rect 3205 2665 3215 2685
rect 3175 2635 3215 2665
rect 3175 2615 3185 2635
rect 3205 2615 3215 2635
rect 3175 2585 3215 2615
rect 3175 2565 3185 2585
rect 3205 2565 3215 2585
rect 3175 2535 3215 2565
rect 3175 2515 3185 2535
rect 3205 2515 3215 2535
rect 3175 2485 3215 2515
rect 3175 2465 3185 2485
rect 3205 2465 3215 2485
rect 3175 2435 3215 2465
rect 3175 2415 3185 2435
rect 3205 2415 3215 2435
rect 3175 2400 3215 2415
rect 3265 2685 3305 2700
rect 3265 2665 3275 2685
rect 3295 2665 3305 2685
rect 3265 2635 3305 2665
rect 3265 2615 3275 2635
rect 3295 2615 3305 2635
rect 3265 2585 3305 2615
rect 3265 2565 3275 2585
rect 3295 2565 3305 2585
rect 3265 2535 3305 2565
rect 3265 2515 3275 2535
rect 3295 2515 3305 2535
rect 3265 2485 3305 2515
rect 3265 2465 3275 2485
rect 3295 2465 3305 2485
rect 3265 2435 3305 2465
rect 3265 2415 3275 2435
rect 3295 2415 3305 2435
rect 3265 2400 3305 2415
rect 3355 2685 3395 2700
rect 3355 2665 3365 2685
rect 3385 2665 3395 2685
rect 3355 2635 3395 2665
rect 3355 2615 3365 2635
rect 3385 2615 3395 2635
rect 3355 2585 3395 2615
rect 3355 2565 3365 2585
rect 3385 2565 3395 2585
rect 3355 2535 3395 2565
rect 3355 2515 3365 2535
rect 3385 2515 3395 2535
rect 3355 2485 3395 2515
rect 3355 2465 3365 2485
rect 3385 2465 3395 2485
rect 3355 2435 3395 2465
rect 3355 2415 3365 2435
rect 3385 2415 3395 2435
rect 3355 2400 3395 2415
rect 3445 2685 3485 2700
rect 3445 2665 3455 2685
rect 3475 2665 3485 2685
rect 3445 2635 3485 2665
rect 3445 2615 3455 2635
rect 3475 2615 3485 2635
rect 3445 2585 3485 2615
rect 3445 2565 3455 2585
rect 3475 2565 3485 2585
rect 3445 2535 3485 2565
rect 3445 2515 3455 2535
rect 3475 2515 3485 2535
rect 3445 2485 3485 2515
rect 3445 2465 3455 2485
rect 3475 2465 3485 2485
rect 3445 2435 3485 2465
rect 3445 2415 3455 2435
rect 3475 2415 3485 2435
rect 3445 2400 3485 2415
rect 3535 2685 3575 2700
rect 3535 2665 3545 2685
rect 3565 2665 3575 2685
rect 3535 2635 3575 2665
rect 3535 2615 3545 2635
rect 3565 2615 3575 2635
rect 3535 2585 3575 2615
rect 3535 2565 3545 2585
rect 3565 2565 3575 2585
rect 3535 2535 3575 2565
rect 3535 2515 3545 2535
rect 3565 2515 3575 2535
rect 3535 2485 3575 2515
rect 3535 2465 3545 2485
rect 3565 2465 3575 2485
rect 3535 2435 3575 2465
rect 3535 2415 3545 2435
rect 3565 2415 3575 2435
rect 3535 2400 3575 2415
rect 3625 2685 3665 2700
rect 3625 2665 3635 2685
rect 3655 2665 3665 2685
rect 3625 2635 3665 2665
rect 3625 2615 3635 2635
rect 3655 2615 3665 2635
rect 3625 2585 3665 2615
rect 3625 2565 3635 2585
rect 3655 2565 3665 2585
rect 3625 2535 3665 2565
rect 3625 2515 3635 2535
rect 3655 2515 3665 2535
rect 3625 2485 3665 2515
rect 3625 2465 3635 2485
rect 3655 2465 3665 2485
rect 3625 2435 3665 2465
rect 3625 2415 3635 2435
rect 3655 2415 3665 2435
rect 3625 2400 3665 2415
rect 3715 2685 3755 2700
rect 3715 2665 3725 2685
rect 3745 2665 3755 2685
rect 3715 2635 3755 2665
rect 3715 2615 3725 2635
rect 3745 2615 3755 2635
rect 3715 2585 3755 2615
rect 3715 2565 3725 2585
rect 3745 2565 3755 2585
rect 3715 2535 3755 2565
rect 3715 2515 3725 2535
rect 3745 2515 3755 2535
rect 3715 2485 3755 2515
rect 3715 2465 3725 2485
rect 3745 2465 3755 2485
rect 3715 2435 3755 2465
rect 3715 2415 3725 2435
rect 3745 2415 3755 2435
rect 3715 2400 3755 2415
rect 3805 2685 3845 2700
rect 3805 2665 3815 2685
rect 3835 2665 3845 2685
rect 3805 2635 3845 2665
rect 3805 2615 3815 2635
rect 3835 2615 3845 2635
rect 3805 2585 3845 2615
rect 3805 2565 3815 2585
rect 3835 2565 3845 2585
rect 3805 2535 3845 2565
rect 3805 2515 3815 2535
rect 3835 2515 3845 2535
rect 3805 2485 3845 2515
rect 3805 2465 3815 2485
rect 3835 2465 3845 2485
rect 3805 2435 3845 2465
rect 3805 2415 3815 2435
rect 3835 2415 3845 2435
rect 3805 2400 3845 2415
rect 3895 2685 3935 2700
rect 3895 2665 3905 2685
rect 3925 2665 3935 2685
rect 3895 2635 3935 2665
rect 3895 2615 3905 2635
rect 3925 2615 3935 2635
rect 3895 2585 3935 2615
rect 3895 2565 3905 2585
rect 3925 2565 3935 2585
rect 3895 2535 3935 2565
rect 3895 2515 3905 2535
rect 3925 2515 3935 2535
rect 3895 2485 3935 2515
rect 3895 2465 3905 2485
rect 3925 2465 3935 2485
rect 3895 2435 3935 2465
rect 3895 2415 3905 2435
rect 3925 2415 3935 2435
rect 3895 2400 3935 2415
rect 3985 2685 4025 2700
rect 3985 2665 3995 2685
rect 4015 2665 4025 2685
rect 3985 2635 4025 2665
rect 3985 2615 3995 2635
rect 4015 2615 4025 2635
rect 3985 2585 4025 2615
rect 3985 2565 3995 2585
rect 4015 2565 4025 2585
rect 3985 2535 4025 2565
rect 3985 2515 3995 2535
rect 4015 2515 4025 2535
rect 3985 2485 4025 2515
rect 3985 2465 3995 2485
rect 4015 2465 4025 2485
rect 3985 2435 4025 2465
rect 3985 2415 3995 2435
rect 4015 2415 4025 2435
rect 3985 2400 4025 2415
rect 4075 2685 4115 2700
rect 4075 2665 4085 2685
rect 4105 2665 4115 2685
rect 4075 2635 4115 2665
rect 4075 2615 4085 2635
rect 4105 2615 4115 2635
rect 4075 2585 4115 2615
rect 4075 2565 4085 2585
rect 4105 2565 4115 2585
rect 4075 2535 4115 2565
rect 4075 2515 4085 2535
rect 4105 2515 4115 2535
rect 4075 2485 4115 2515
rect 4075 2465 4085 2485
rect 4105 2465 4115 2485
rect 4075 2435 4115 2465
rect 4075 2415 4085 2435
rect 4105 2415 4115 2435
rect 4075 2400 4115 2415
rect 4165 2685 4205 2700
rect 4165 2665 4175 2685
rect 4195 2665 4205 2685
rect 4165 2635 4205 2665
rect 4165 2615 4175 2635
rect 4195 2615 4205 2635
rect 4165 2585 4205 2615
rect 4165 2565 4175 2585
rect 4195 2565 4205 2585
rect 4165 2535 4205 2565
rect 4165 2515 4175 2535
rect 4195 2515 4205 2535
rect 4165 2485 4205 2515
rect 4165 2465 4175 2485
rect 4195 2465 4205 2485
rect 4165 2435 4205 2465
rect 4165 2415 4175 2435
rect 4195 2415 4205 2435
rect 4165 2400 4205 2415
rect 4255 2685 4295 2700
rect 4255 2665 4265 2685
rect 4285 2665 4295 2685
rect 4255 2635 4295 2665
rect 4255 2615 4265 2635
rect 4285 2615 4295 2635
rect 4255 2585 4295 2615
rect 4255 2565 4265 2585
rect 4285 2565 4295 2585
rect 4255 2535 4295 2565
rect 4255 2515 4265 2535
rect 4285 2515 4295 2535
rect 4255 2485 4295 2515
rect 4255 2465 4265 2485
rect 4285 2465 4295 2485
rect 4255 2435 4295 2465
rect 4255 2415 4265 2435
rect 4285 2415 4295 2435
rect 4255 2400 4295 2415
rect 4345 2685 4385 2700
rect 4345 2665 4355 2685
rect 4375 2665 4385 2685
rect 4345 2635 4385 2665
rect 4345 2615 4355 2635
rect 4375 2615 4385 2635
rect 4345 2585 4385 2615
rect 4345 2565 4355 2585
rect 4375 2565 4385 2585
rect 4345 2535 4385 2565
rect 4345 2515 4355 2535
rect 4375 2515 4385 2535
rect 4345 2485 4385 2515
rect 4345 2465 4355 2485
rect 4375 2465 4385 2485
rect 4345 2435 4385 2465
rect 4345 2415 4355 2435
rect 4375 2415 4385 2435
rect 4345 2400 4385 2415
rect 4435 2685 4475 2700
rect 4435 2665 4445 2685
rect 4465 2665 4475 2685
rect 4435 2635 4475 2665
rect 4435 2615 4445 2635
rect 4465 2615 4475 2635
rect 4435 2585 4475 2615
rect 4435 2565 4445 2585
rect 4465 2565 4475 2585
rect 4435 2535 4475 2565
rect 4435 2515 4445 2535
rect 4465 2515 4475 2535
rect 4435 2485 4475 2515
rect 4435 2465 4445 2485
rect 4465 2465 4475 2485
rect 4435 2435 4475 2465
rect 4435 2415 4445 2435
rect 4465 2415 4475 2435
rect 4435 2400 4475 2415
rect 4525 2685 4565 2700
rect 4525 2665 4535 2685
rect 4555 2665 4565 2685
rect 4525 2635 4565 2665
rect 4525 2615 4535 2635
rect 4555 2615 4565 2635
rect 4525 2585 4565 2615
rect 4525 2565 4535 2585
rect 4555 2565 4565 2585
rect 4525 2535 4565 2565
rect 4525 2515 4535 2535
rect 4555 2515 4565 2535
rect 4525 2485 4565 2515
rect 4525 2465 4535 2485
rect 4555 2465 4565 2485
rect 4525 2435 4565 2465
rect 4525 2415 4535 2435
rect 4555 2415 4565 2435
rect 4525 2400 4565 2415
rect 4615 2685 4655 2700
rect 4615 2665 4625 2685
rect 4645 2665 4655 2685
rect 4615 2635 4655 2665
rect 4615 2615 4625 2635
rect 4645 2615 4655 2635
rect 4615 2585 4655 2615
rect 4615 2565 4625 2585
rect 4645 2565 4655 2585
rect 4615 2535 4655 2565
rect 4615 2515 4625 2535
rect 4645 2515 4655 2535
rect 4615 2485 4655 2515
rect 4615 2465 4625 2485
rect 4645 2465 4655 2485
rect 4615 2435 4655 2465
rect 4615 2415 4625 2435
rect 4645 2415 4655 2435
rect 4615 2400 4655 2415
rect 4705 2685 4745 2700
rect 4705 2665 4715 2685
rect 4735 2665 4745 2685
rect 4705 2635 4745 2665
rect 4705 2615 4715 2635
rect 4735 2615 4745 2635
rect 4705 2585 4745 2615
rect 4705 2565 4715 2585
rect 4735 2565 4745 2585
rect 4705 2535 4745 2565
rect 4705 2515 4715 2535
rect 4735 2515 4745 2535
rect 4705 2485 4745 2515
rect 4705 2465 4715 2485
rect 4735 2465 4745 2485
rect 4705 2435 4745 2465
rect 4705 2415 4715 2435
rect 4735 2415 4745 2435
rect 4705 2400 4745 2415
rect 4795 2685 4835 2700
rect 4795 2665 4805 2685
rect 4825 2665 4835 2685
rect 4795 2635 4835 2665
rect 4795 2615 4805 2635
rect 4825 2615 4835 2635
rect 4795 2585 4835 2615
rect 4795 2565 4805 2585
rect 4825 2565 4835 2585
rect 4795 2535 4835 2565
rect 4795 2515 4805 2535
rect 4825 2515 4835 2535
rect 4795 2485 4835 2515
rect 4795 2465 4805 2485
rect 4825 2465 4835 2485
rect 4795 2435 4835 2465
rect 4795 2415 4805 2435
rect 4825 2415 4835 2435
rect 4795 2400 4835 2415
rect 2565 1985 2605 2000
rect 2565 1965 2575 1985
rect 2595 1965 2605 1985
rect 2565 1935 2605 1965
rect 2565 1915 2575 1935
rect 2595 1915 2605 1935
rect 2565 1900 2605 1915
rect 2620 1985 2660 2000
rect 2620 1965 2630 1985
rect 2650 1965 2660 1985
rect 2620 1935 2660 1965
rect 2620 1915 2630 1935
rect 2650 1915 2660 1935
rect 2620 1900 2660 1915
rect 2675 1985 2715 2000
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1900 2715 1915
rect 2745 1985 2785 2000
rect 2745 1965 2755 1985
rect 2775 1965 2785 1985
rect 2745 1935 2785 1965
rect 2745 1915 2755 1935
rect 2775 1915 2785 1935
rect 2745 1900 2785 1915
rect 2805 1985 2845 2000
rect 2805 1965 2815 1985
rect 2835 1965 2845 1985
rect 2805 1935 2845 1965
rect 2805 1915 2815 1935
rect 2835 1915 2845 1935
rect 2805 1900 2845 1915
rect 2865 1985 2905 2000
rect 2865 1965 2875 1985
rect 2895 1965 2905 1985
rect 2865 1935 2905 1965
rect 2865 1915 2875 1935
rect 2895 1915 2905 1935
rect 2865 1900 2905 1915
rect 2925 1985 2965 2000
rect 2925 1965 2935 1985
rect 2955 1965 2965 1985
rect 2925 1935 2965 1965
rect 2925 1915 2935 1935
rect 2955 1915 2965 1935
rect 2925 1900 2965 1915
rect 2985 1985 3025 2000
rect 2985 1965 2995 1985
rect 3015 1965 3025 1985
rect 2985 1935 3025 1965
rect 2985 1915 2995 1935
rect 3015 1915 3025 1935
rect 2985 1900 3025 1915
rect 3045 1985 3085 2000
rect 3045 1965 3055 1985
rect 3075 1965 3085 1985
rect 3045 1935 3085 1965
rect 3045 1915 3055 1935
rect 3075 1915 3085 1935
rect 3045 1900 3085 1915
rect 3105 1985 3145 2000
rect 3105 1965 3115 1985
rect 3135 1965 3145 1985
rect 3105 1935 3145 1965
rect 3105 1915 3115 1935
rect 3135 1915 3145 1935
rect 3105 1900 3145 1915
rect 3165 1985 3205 2000
rect 3165 1965 3175 1985
rect 3195 1965 3205 1985
rect 3165 1935 3205 1965
rect 3165 1915 3175 1935
rect 3195 1915 3205 1935
rect 3165 1900 3205 1915
rect 3225 1985 3265 2000
rect 3225 1965 3235 1985
rect 3255 1965 3265 1985
rect 3225 1935 3265 1965
rect 3225 1915 3235 1935
rect 3255 1915 3265 1935
rect 3225 1900 3265 1915
rect 3285 1985 3325 2000
rect 3285 1965 3295 1985
rect 3315 1965 3325 1985
rect 3285 1935 3325 1965
rect 3285 1915 3295 1935
rect 3315 1915 3325 1935
rect 3285 1900 3325 1915
rect 3345 1985 3385 2000
rect 3345 1965 3355 1985
rect 3375 1965 3385 1985
rect 3345 1935 3385 1965
rect 3345 1915 3355 1935
rect 3375 1915 3385 1935
rect 3345 1900 3385 1915
rect 3405 1985 3445 2000
rect 3405 1965 3415 1985
rect 3435 1965 3445 1985
rect 3405 1935 3445 1965
rect 3405 1915 3415 1935
rect 3435 1915 3445 1935
rect 3405 1900 3445 1915
rect 3465 1985 3505 2000
rect 3465 1965 3475 1985
rect 3495 1965 3505 1985
rect 3465 1935 3505 1965
rect 3465 1915 3475 1935
rect 3495 1915 3505 1935
rect 3465 1900 3505 1915
rect 3525 1985 3565 2000
rect 3525 1965 3535 1985
rect 3555 1965 3565 1985
rect 3525 1935 3565 1965
rect 3525 1915 3535 1935
rect 3555 1915 3565 1935
rect 3525 1900 3565 1915
rect 3585 1985 3625 2000
rect 3585 1965 3595 1985
rect 3615 1965 3625 1985
rect 3585 1935 3625 1965
rect 3585 1915 3595 1935
rect 3615 1915 3625 1935
rect 3585 1900 3625 1915
rect 3645 1985 3685 2000
rect 3645 1965 3655 1985
rect 3675 1965 3685 1985
rect 3645 1935 3685 1965
rect 3645 1915 3655 1935
rect 3675 1915 3685 1935
rect 3645 1900 3685 1915
rect 3705 1985 3745 2000
rect 3705 1965 3715 1985
rect 3735 1965 3745 1985
rect 3705 1935 3745 1965
rect 3705 1915 3715 1935
rect 3735 1915 3745 1935
rect 3705 1900 3745 1915
rect 3765 1985 3805 2000
rect 3765 1965 3775 1985
rect 3795 1965 3805 1985
rect 3765 1935 3805 1965
rect 3765 1915 3775 1935
rect 3795 1915 3805 1935
rect 3765 1900 3805 1915
rect 3825 1985 3865 2000
rect 3825 1965 3835 1985
rect 3855 1965 3865 1985
rect 3825 1935 3865 1965
rect 3825 1915 3835 1935
rect 3855 1915 3865 1935
rect 3825 1900 3865 1915
rect 3885 1985 3925 2000
rect 3885 1965 3895 1985
rect 3915 1965 3925 1985
rect 3885 1935 3925 1965
rect 3885 1915 3895 1935
rect 3915 1915 3925 1935
rect 3885 1900 3925 1915
rect 3945 1985 3985 2000
rect 4025 1985 4065 2000
rect 3945 1965 3955 1985
rect 3975 1965 3985 1985
rect 4025 1965 4035 1985
rect 4055 1965 4065 1985
rect 3945 1935 3985 1965
rect 4025 1935 4065 1965
rect 3945 1915 3955 1935
rect 3975 1915 3985 1935
rect 4025 1915 4035 1935
rect 4055 1915 4065 1935
rect 3945 1900 3985 1915
rect 4025 1900 4065 1915
rect 4085 1985 4125 2000
rect 4085 1965 4095 1985
rect 4115 1965 4125 1985
rect 4085 1935 4125 1965
rect 4085 1915 4095 1935
rect 4115 1915 4125 1935
rect 4085 1900 4125 1915
rect 4145 1985 4185 2000
rect 4145 1965 4155 1985
rect 4175 1965 4185 1985
rect 4145 1935 4185 1965
rect 4145 1915 4155 1935
rect 4175 1915 4185 1935
rect 4145 1900 4185 1915
rect 4205 1985 4245 2000
rect 4205 1965 4215 1985
rect 4235 1965 4245 1985
rect 4205 1935 4245 1965
rect 4205 1915 4215 1935
rect 4235 1915 4245 1935
rect 4205 1900 4245 1915
rect 4265 1985 4305 2000
rect 4265 1965 4275 1985
rect 4295 1965 4305 1985
rect 4265 1935 4305 1965
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1900 4305 1915
rect 4325 1985 4365 2000
rect 4325 1965 4335 1985
rect 4355 1965 4365 1985
rect 4325 1935 4365 1965
rect 4325 1915 4335 1935
rect 4355 1915 4365 1935
rect 4325 1900 4365 1915
rect 4385 1985 4425 2000
rect 4385 1965 4395 1985
rect 4415 1965 4425 1985
rect 4385 1935 4425 1965
rect 4385 1915 4395 1935
rect 4415 1915 4425 1935
rect 4385 1900 4425 1915
rect 4445 1985 4485 2000
rect 4445 1965 4455 1985
rect 4475 1965 4485 1985
rect 4445 1935 4485 1965
rect 4445 1915 4455 1935
rect 4475 1915 4485 1935
rect 4445 1900 4485 1915
rect 4505 1985 4545 2000
rect 4505 1965 4515 1985
rect 4535 1965 4545 1985
rect 4505 1935 4545 1965
rect 4505 1915 4515 1935
rect 4535 1915 4545 1935
rect 4505 1900 4545 1915
rect 4565 1985 4605 2000
rect 4565 1965 4575 1985
rect 4595 1965 4605 1985
rect 4565 1935 4605 1965
rect 4565 1915 4575 1935
rect 4595 1915 4605 1935
rect 4565 1900 4605 1915
rect 4625 1985 4665 2000
rect 4625 1965 4635 1985
rect 4655 1965 4665 1985
rect 4625 1935 4665 1965
rect 4625 1915 4635 1935
rect 4655 1915 4665 1935
rect 4625 1900 4665 1915
rect 4685 1985 4725 2000
rect 4685 1965 4695 1985
rect 4715 1965 4725 1985
rect 4685 1935 4725 1965
rect 4685 1915 4695 1935
rect 4715 1915 4725 1935
rect 4685 1900 4725 1915
rect 4745 1985 4785 2000
rect 4745 1965 4755 1985
rect 4775 1965 4785 1985
rect 4745 1935 4785 1965
rect 4745 1915 4755 1935
rect 4775 1915 4785 1935
rect 4745 1900 4785 1915
rect 4805 1985 4845 2000
rect 4805 1965 4815 1985
rect 4835 1965 4845 1985
rect 4805 1935 4845 1965
rect 4805 1915 4815 1935
rect 4835 1915 4845 1935
rect 4805 1900 4845 1915
rect 4865 1985 4905 2000
rect 4865 1965 4875 1985
rect 4895 1965 4905 1985
rect 4865 1935 4905 1965
rect 4865 1915 4875 1935
rect 4895 1915 4905 1935
rect 4865 1900 4905 1915
rect 4925 1985 4965 2000
rect 4925 1965 4935 1985
rect 4955 1965 4965 1985
rect 4925 1935 4965 1965
rect 4925 1915 4935 1935
rect 4955 1915 4965 1935
rect 4925 1900 4965 1915
rect 4985 1985 5025 2000
rect 4985 1965 4995 1985
rect 5015 1965 5025 1985
rect 4985 1935 5025 1965
rect 4985 1915 4995 1935
rect 5015 1915 5025 1935
rect 4985 1900 5025 1915
rect 5045 1985 5085 2000
rect 5045 1965 5055 1985
rect 5075 1965 5085 1985
rect 5045 1935 5085 1965
rect 5045 1915 5055 1935
rect 5075 1915 5085 1935
rect 5045 1900 5085 1915
rect 5105 1985 5145 2000
rect 5105 1965 5115 1985
rect 5135 1965 5145 1985
rect 5105 1935 5145 1965
rect 5105 1915 5115 1935
rect 5135 1915 5145 1935
rect 5105 1900 5145 1915
rect 5165 1985 5205 2000
rect 5165 1965 5175 1985
rect 5195 1965 5205 1985
rect 5165 1935 5205 1965
rect 5165 1915 5175 1935
rect 5195 1915 5205 1935
rect 5165 1900 5205 1915
rect 5225 1985 5265 2000
rect 5225 1965 5235 1985
rect 5255 1965 5265 1985
rect 5225 1935 5265 1965
rect 5225 1915 5235 1935
rect 5255 1915 5265 1935
rect 5225 1900 5265 1915
<< ndiffc >>
rect 11250 8895 11270 8915
rect 11310 8900 11330 8920
rect 11370 8900 11390 8920
rect 11430 8895 11450 8915
rect 11580 8910 11600 8930
rect 11640 8910 11660 8930
rect 11700 8910 11720 8930
rect 11760 8910 11780 8930
rect 11820 8910 11840 8930
rect 11880 8910 11900 8930
rect 11940 8910 11960 8930
rect 12090 8895 12110 8915
rect 12150 8895 12170 8915
rect 12210 8895 12230 8915
rect 12270 8895 12290 8915
rect 12330 8895 12350 8915
rect 12390 8895 12410 8915
rect 12450 8895 12470 8915
rect 12510 8895 12530 8915
rect 12570 8895 12590 8915
rect 10830 8495 10850 8515
rect 10830 8445 10850 8465
rect 10830 8395 10850 8415
rect 10830 8345 10850 8365
rect 10830 8295 10850 8315
rect 10500 8245 10520 8265
rect 10560 8250 10580 8270
rect 10620 8250 10640 8270
rect 10680 8245 10700 8265
rect 10830 8245 10850 8265
rect 10890 8495 10910 8515
rect 10890 8445 10910 8465
rect 10890 8395 10910 8415
rect 10890 8345 10910 8365
rect 10890 8295 10910 8315
rect 10890 8245 10910 8265
rect 10950 8495 10970 8515
rect 10950 8445 10970 8465
rect 10950 8395 10970 8415
rect 10950 8345 10970 8365
rect 10950 8295 10970 8315
rect 10950 8245 10970 8265
rect 11010 8545 11030 8565
rect 11010 8495 11030 8515
rect 11010 8445 11030 8465
rect 11010 8395 11030 8415
rect 11010 8345 11030 8365
rect 11010 8295 11030 8315
rect 11010 8245 11030 8265
rect 11070 8545 11090 8565
rect 11070 8495 11090 8515
rect 11070 8445 11090 8465
rect 11070 8395 11090 8415
rect 11070 8345 11090 8365
rect 11070 8295 11090 8315
rect 11070 8245 11090 8265
rect 11230 8540 11250 8560
rect 11230 8490 11250 8510
rect 11230 8440 11250 8460
rect 11230 8390 11250 8410
rect 11230 8340 11250 8360
rect 11230 8290 11250 8310
rect 11230 8240 11250 8260
rect 11230 8190 11250 8210
rect 11290 8540 11310 8560
rect 11290 8490 11310 8510
rect 11290 8440 11310 8460
rect 11290 8390 11310 8410
rect 11290 8340 11310 8360
rect 11290 8290 11310 8310
rect 11290 8240 11310 8260
rect 11290 8190 11310 8210
rect 11350 8540 11370 8560
rect 11350 8490 11370 8510
rect 11350 8440 11370 8460
rect 11350 8390 11370 8410
rect 11350 8340 11370 8360
rect 11350 8290 11370 8310
rect 11350 8240 11370 8260
rect 11350 8190 11370 8210
rect 11410 8540 11430 8560
rect 11410 8490 11430 8510
rect 11410 8440 11430 8460
rect 11410 8390 11430 8410
rect 11410 8340 11430 8360
rect 11410 8290 11430 8310
rect 11410 8240 11430 8260
rect 11410 8190 11430 8210
rect 11470 8540 11490 8560
rect 11470 8490 11490 8510
rect 11470 8440 11490 8460
rect 11470 8390 11490 8410
rect 11470 8340 11490 8360
rect 11470 8290 11490 8310
rect 11470 8240 11490 8260
rect 11470 8190 11490 8210
rect 11530 8540 11550 8560
rect 11530 8490 11550 8510
rect 11530 8440 11550 8460
rect 11530 8390 11550 8410
rect 11530 8340 11550 8360
rect 11530 8290 11550 8310
rect 11530 8240 11550 8260
rect 11530 8190 11550 8210
rect 11590 8540 11610 8560
rect 11590 8490 11610 8510
rect 11590 8440 11610 8460
rect 11590 8390 11610 8410
rect 11590 8340 11610 8360
rect 11590 8290 11610 8310
rect 11590 8240 11610 8260
rect 11590 8190 11610 8210
rect 11650 8540 11670 8560
rect 11650 8490 11670 8510
rect 11650 8440 11670 8460
rect 11650 8390 11670 8410
rect 11650 8340 11670 8360
rect 11650 8290 11670 8310
rect 11650 8240 11670 8260
rect 11650 8190 11670 8210
rect 11710 8540 11730 8560
rect 11710 8490 11730 8510
rect 11710 8440 11730 8460
rect 11710 8390 11730 8410
rect 11710 8340 11730 8360
rect 11710 8290 11730 8310
rect 11710 8240 11730 8260
rect 11710 8190 11730 8210
rect 11770 8540 11790 8560
rect 11770 8490 11790 8510
rect 11770 8440 11790 8460
rect 11770 8390 11790 8410
rect 11770 8340 11790 8360
rect 11770 8290 11790 8310
rect 11770 8240 11790 8260
rect 11770 8190 11790 8210
rect 11830 8540 11850 8560
rect 11830 8490 11850 8510
rect 11830 8440 11850 8460
rect 11830 8390 11850 8410
rect 11830 8340 11850 8360
rect 11830 8290 11850 8310
rect 11830 8240 11850 8260
rect 11830 8190 11850 8210
rect 11890 8540 11910 8560
rect 11890 8490 11910 8510
rect 11890 8440 11910 8460
rect 11890 8390 11910 8410
rect 11890 8340 11910 8360
rect 11890 8290 11910 8310
rect 11890 8240 11910 8260
rect 11890 8190 11910 8210
rect 11950 8540 11970 8560
rect 11950 8490 11970 8510
rect 11950 8440 11970 8460
rect 11950 8390 11970 8410
rect 11950 8340 11970 8360
rect 11950 8290 11970 8310
rect 11950 8240 11970 8260
rect 11950 8190 11970 8210
rect 12010 8540 12030 8560
rect 12010 8490 12030 8510
rect 12010 8440 12030 8460
rect 12010 8390 12030 8410
rect 12010 8340 12030 8360
rect 12010 8290 12030 8310
rect 12010 8240 12030 8260
rect 12010 8190 12030 8210
rect 12070 8540 12090 8560
rect 12070 8490 12090 8510
rect 12070 8440 12090 8460
rect 12070 8390 12090 8410
rect 12070 8340 12090 8360
rect 12070 8290 12090 8310
rect 12070 8240 12090 8260
rect 12070 8190 12090 8210
rect 12130 8540 12150 8560
rect 12130 8490 12150 8510
rect 12130 8440 12150 8460
rect 12130 8390 12150 8410
rect 12130 8340 12150 8360
rect 12130 8290 12150 8310
rect 12130 8240 12150 8260
rect 12130 8190 12150 8210
rect 12190 8540 12210 8560
rect 12190 8490 12210 8510
rect 12190 8440 12210 8460
rect 12190 8390 12210 8410
rect 12190 8340 12210 8360
rect 12190 8290 12210 8310
rect 12190 8240 12210 8260
rect 12190 8190 12210 8210
rect 12250 8540 12270 8560
rect 12250 8490 12270 8510
rect 12250 8440 12270 8460
rect 12250 8390 12270 8410
rect 12250 8340 12270 8360
rect 12250 8290 12270 8310
rect 12250 8240 12270 8260
rect 12250 8190 12270 8210
rect 12310 8540 12330 8560
rect 12310 8490 12330 8510
rect 12310 8440 12330 8460
rect 12310 8390 12330 8410
rect 12310 8340 12330 8360
rect 12310 8290 12330 8310
rect 12310 8240 12330 8260
rect 12310 8190 12330 8210
rect 12370 8540 12390 8560
rect 12370 8490 12390 8510
rect 12370 8440 12390 8460
rect 12370 8390 12390 8410
rect 12370 8340 12390 8360
rect 12370 8290 12390 8310
rect 12370 8240 12390 8260
rect 12370 8190 12390 8210
rect 12430 8540 12450 8560
rect 12430 8490 12450 8510
rect 12430 8440 12450 8460
rect 12430 8390 12450 8410
rect 12430 8340 12450 8360
rect 12430 8290 12450 8310
rect 12430 8240 12450 8260
rect 12430 8190 12450 8210
rect 12490 8540 12510 8560
rect 12490 8490 12510 8510
rect 12490 8440 12510 8460
rect 12490 8390 12510 8410
rect 12490 8340 12510 8360
rect 12490 8290 12510 8310
rect 12490 8240 12510 8260
rect 12490 8190 12510 8210
rect 12550 8540 12570 8560
rect 12550 8490 12570 8510
rect 12550 8440 12570 8460
rect 12550 8390 12570 8410
rect 12550 8340 12570 8360
rect 18330 8495 18350 8515
rect 18330 8445 18350 8465
rect 18330 8395 18350 8415
rect 12550 8290 12570 8310
rect 18330 8345 18350 8365
rect 18330 8295 18350 8315
rect 12550 8240 12570 8260
rect 18000 8245 18020 8265
rect 12550 8190 12570 8210
rect 12905 8205 12925 8225
rect 12905 8155 12925 8175
rect 12905 8105 12925 8125
rect 12905 8055 12925 8075
rect 12905 8005 12925 8025
rect 12905 7955 12925 7975
rect 12960 8205 12980 8225
rect 12960 8155 12980 8175
rect 12960 8105 12980 8125
rect 12960 8055 12980 8075
rect 12960 8005 12980 8025
rect 12960 7955 12980 7975
rect 13015 8205 13035 8225
rect 13015 8155 13035 8175
rect 13015 8105 13035 8125
rect 13015 8055 13035 8075
rect 13015 8005 13035 8025
rect 13015 7955 13035 7975
rect 13070 8205 13090 8225
rect 13070 8155 13090 8175
rect 13070 8105 13090 8125
rect 13070 8055 13090 8075
rect 13070 8005 13090 8025
rect 13070 7955 13090 7975
rect 13125 8205 13145 8225
rect 13125 8155 13145 8175
rect 13125 8105 13145 8125
rect 13125 8055 13145 8075
rect 13125 8005 13145 8025
rect 13125 7955 13145 7975
rect 13180 8205 13200 8225
rect 13180 8155 13200 8175
rect 13180 8105 13200 8125
rect 13180 8055 13200 8075
rect 13180 8005 13200 8025
rect 13180 7955 13200 7975
rect 13235 8205 13255 8225
rect 13235 8155 13255 8175
rect 13235 8105 13255 8125
rect 13235 8055 13255 8075
rect 13235 8005 13255 8025
rect 13235 7955 13255 7975
rect 13290 8205 13310 8225
rect 13290 8155 13310 8175
rect 13290 8105 13310 8125
rect 13290 8055 13310 8075
rect 13290 8005 13310 8025
rect 13290 7955 13310 7975
rect 13345 8205 13365 8225
rect 13345 8155 13365 8175
rect 13345 8105 13365 8125
rect 13345 8055 13365 8075
rect 13345 8005 13365 8025
rect 13345 7955 13365 7975
rect 13400 8205 13420 8225
rect 13400 8155 13420 8175
rect 13400 8105 13420 8125
rect 13400 8055 13420 8075
rect 13400 8005 13420 8025
rect 13400 7955 13420 7975
rect 13455 8205 13475 8225
rect 13455 8155 13475 8175
rect 13455 8105 13475 8125
rect 13455 8055 13475 8075
rect 13455 8005 13475 8025
rect 13455 7955 13475 7975
rect 13510 8205 13530 8225
rect 13510 8155 13530 8175
rect 13510 8105 13530 8125
rect 13510 8055 13530 8075
rect 13510 8005 13530 8025
rect 13510 7955 13530 7975
rect 13565 8205 13585 8225
rect 13565 8155 13585 8175
rect 13565 8105 13585 8125
rect 13565 8055 13585 8075
rect 13565 8005 13585 8025
rect 13565 7955 13585 7975
rect 13620 8205 13640 8225
rect 13620 8155 13640 8175
rect 13620 8105 13640 8125
rect 13620 8055 13640 8075
rect 13620 8005 13640 8025
rect 13620 7955 13640 7975
rect 13675 8205 13695 8225
rect 13675 8155 13695 8175
rect 13675 8105 13695 8125
rect 13675 8055 13695 8075
rect 13675 8005 13695 8025
rect 13675 7955 13695 7975
rect 13730 8205 13750 8225
rect 13730 8155 13750 8175
rect 13730 8105 13750 8125
rect 13730 8055 13750 8075
rect 13730 8005 13750 8025
rect 13730 7955 13750 7975
rect 13785 8205 13805 8225
rect 13785 8155 13805 8175
rect 13785 8105 13805 8125
rect 13785 8055 13805 8075
rect 13785 8005 13805 8025
rect 13785 7955 13805 7975
rect 13840 8205 13860 8225
rect 13840 8155 13860 8175
rect 13840 8105 13860 8125
rect 13840 8055 13860 8075
rect 13840 8005 13860 8025
rect 13840 7955 13860 7975
rect 13895 8205 13915 8225
rect 13895 8155 13915 8175
rect 13895 8105 13915 8125
rect 13895 8055 13915 8075
rect 13895 8005 13915 8025
rect 13895 7955 13915 7975
rect 13950 8205 13970 8225
rect 13950 8155 13970 8175
rect 13950 8105 13970 8125
rect 13950 8055 13970 8075
rect 13950 8005 13970 8025
rect 13950 7955 13970 7975
rect 14005 8205 14025 8225
rect 14005 8155 14025 8175
rect 14005 8105 14025 8125
rect 14005 8055 14025 8075
rect 14005 8005 14025 8025
rect 14005 7955 14025 7975
rect 14060 8205 14080 8225
rect 14060 8155 14080 8175
rect 14060 8105 14080 8125
rect 14060 8055 14080 8075
rect 14060 8005 14080 8025
rect 14060 7955 14080 7975
rect 18060 8250 18080 8270
rect 18120 8250 18140 8270
rect 18180 8245 18200 8265
rect 18330 8245 18350 8265
rect 18390 8495 18410 8515
rect 18390 8445 18410 8465
rect 18390 8395 18410 8415
rect 18390 8345 18410 8365
rect 18390 8295 18410 8315
rect 18390 8245 18410 8265
rect 18450 8495 18470 8515
rect 18450 8445 18470 8465
rect 18450 8395 18470 8415
rect 18450 8345 18470 8365
rect 18450 8295 18470 8315
rect 18450 8245 18470 8265
rect 18510 8545 18530 8565
rect 18510 8495 18530 8515
rect 18510 8445 18530 8465
rect 18510 8395 18530 8415
rect 18510 8345 18530 8365
rect 18510 8295 18530 8315
rect 18510 8245 18530 8265
rect 18570 8545 18590 8565
rect 18570 8495 18590 8515
rect 18570 8445 18590 8465
rect 18570 8395 18590 8415
rect 18570 8345 18590 8365
rect 18570 8295 18590 8315
rect 18570 8245 18590 8265
rect 18730 8540 18750 8560
rect 18730 8490 18750 8510
rect 18730 8440 18750 8460
rect 18730 8390 18750 8410
rect 18730 8340 18750 8360
rect 18730 8290 18750 8310
rect 18730 8240 18750 8260
rect 14115 8205 14135 8225
rect 18730 8190 18750 8210
rect 18790 8540 18810 8560
rect 18790 8490 18810 8510
rect 18790 8440 18810 8460
rect 18790 8390 18810 8410
rect 18790 8340 18810 8360
rect 18790 8290 18810 8310
rect 18790 8240 18810 8260
rect 18790 8190 18810 8210
rect 18850 8540 18870 8560
rect 18850 8490 18870 8510
rect 18850 8440 18870 8460
rect 18850 8390 18870 8410
rect 18850 8340 18870 8360
rect 18850 8290 18870 8310
rect 18850 8240 18870 8260
rect 18850 8190 18870 8210
rect 18910 8540 18930 8560
rect 18910 8490 18930 8510
rect 18910 8440 18930 8460
rect 18910 8390 18930 8410
rect 18910 8340 18930 8360
rect 18910 8290 18930 8310
rect 18910 8240 18930 8260
rect 18910 8190 18930 8210
rect 18970 8540 18990 8560
rect 18970 8490 18990 8510
rect 18970 8440 18990 8460
rect 18970 8390 18990 8410
rect 18970 8340 18990 8360
rect 18970 8290 18990 8310
rect 18970 8240 18990 8260
rect 18970 8190 18990 8210
rect 19030 8540 19050 8560
rect 19030 8490 19050 8510
rect 19030 8440 19050 8460
rect 19030 8390 19050 8410
rect 19030 8340 19050 8360
rect 19030 8290 19050 8310
rect 19030 8240 19050 8260
rect 19030 8190 19050 8210
rect 19090 8540 19110 8560
rect 19090 8490 19110 8510
rect 19090 8440 19110 8460
rect 19090 8390 19110 8410
rect 19090 8340 19110 8360
rect 19090 8290 19110 8310
rect 19090 8240 19110 8260
rect 19090 8190 19110 8210
rect 19150 8540 19170 8560
rect 19150 8490 19170 8510
rect 19150 8440 19170 8460
rect 19150 8390 19170 8410
rect 19150 8340 19170 8360
rect 19150 8290 19170 8310
rect 19150 8240 19170 8260
rect 19150 8190 19170 8210
rect 19210 8540 19230 8560
rect 19210 8490 19230 8510
rect 19210 8440 19230 8460
rect 19210 8390 19230 8410
rect 19210 8340 19230 8360
rect 19210 8290 19230 8310
rect 19210 8240 19230 8260
rect 19210 8190 19230 8210
rect 19270 8540 19290 8560
rect 19270 8490 19290 8510
rect 19270 8440 19290 8460
rect 19270 8390 19290 8410
rect 19270 8340 19290 8360
rect 19270 8290 19290 8310
rect 19270 8240 19290 8260
rect 19270 8190 19290 8210
rect 19330 8540 19350 8560
rect 19330 8490 19350 8510
rect 19330 8440 19350 8460
rect 19330 8390 19350 8410
rect 19330 8340 19350 8360
rect 19330 8290 19350 8310
rect 19330 8240 19350 8260
rect 19330 8190 19350 8210
rect 19390 8540 19410 8560
rect 19390 8490 19410 8510
rect 19390 8440 19410 8460
rect 19390 8390 19410 8410
rect 19390 8340 19410 8360
rect 19390 8290 19410 8310
rect 19390 8240 19410 8260
rect 19390 8190 19410 8210
rect 19450 8540 19470 8560
rect 19450 8490 19470 8510
rect 19450 8440 19470 8460
rect 19450 8390 19470 8410
rect 19450 8340 19470 8360
rect 19450 8290 19470 8310
rect 19450 8240 19470 8260
rect 19450 8190 19470 8210
rect 19510 8540 19530 8560
rect 19510 8490 19530 8510
rect 19510 8440 19530 8460
rect 19510 8390 19530 8410
rect 19510 8340 19530 8360
rect 19510 8290 19530 8310
rect 19510 8240 19530 8260
rect 19510 8190 19530 8210
rect 19570 8540 19590 8560
rect 19570 8490 19590 8510
rect 19570 8440 19590 8460
rect 19570 8390 19590 8410
rect 19570 8340 19590 8360
rect 19570 8290 19590 8310
rect 19570 8240 19590 8260
rect 19570 8190 19590 8210
rect 19630 8540 19650 8560
rect 19630 8490 19650 8510
rect 19630 8440 19650 8460
rect 19630 8390 19650 8410
rect 19630 8340 19650 8360
rect 19630 8290 19650 8310
rect 19630 8240 19650 8260
rect 19630 8190 19650 8210
rect 19690 8540 19710 8560
rect 19690 8490 19710 8510
rect 19690 8440 19710 8460
rect 19690 8390 19710 8410
rect 19690 8340 19710 8360
rect 19690 8290 19710 8310
rect 19690 8240 19710 8260
rect 19690 8190 19710 8210
rect 19750 8540 19770 8560
rect 19750 8490 19770 8510
rect 19750 8440 19770 8460
rect 19750 8390 19770 8410
rect 19750 8340 19770 8360
rect 19750 8290 19770 8310
rect 19750 8240 19770 8260
rect 19750 8190 19770 8210
rect 19810 8540 19830 8560
rect 19810 8490 19830 8510
rect 19810 8440 19830 8460
rect 19810 8390 19830 8410
rect 19810 8340 19830 8360
rect 19810 8290 19830 8310
rect 19810 8240 19830 8260
rect 19810 8190 19830 8210
rect 19870 8540 19890 8560
rect 19870 8490 19890 8510
rect 19870 8440 19890 8460
rect 19870 8390 19890 8410
rect 19870 8340 19890 8360
rect 19870 8290 19890 8310
rect 19870 8240 19890 8260
rect 19870 8190 19890 8210
rect 19930 8540 19950 8560
rect 19930 8490 19950 8510
rect 19930 8440 19950 8460
rect 19930 8390 19950 8410
rect 19930 8340 19950 8360
rect 19930 8290 19950 8310
rect 19930 8240 19950 8260
rect 19930 8190 19950 8210
rect 19990 8540 20010 8560
rect 19990 8490 20010 8510
rect 19990 8440 20010 8460
rect 19990 8390 20010 8410
rect 19990 8340 20010 8360
rect 19990 8290 20010 8310
rect 19990 8240 20010 8260
rect 19990 8190 20010 8210
rect 20050 8540 20070 8560
rect 20050 8490 20070 8510
rect 20050 8440 20070 8460
rect 20050 8390 20070 8410
rect 20050 8340 20070 8360
rect 20050 8290 20070 8310
rect 20050 8240 20070 8260
rect 20050 8190 20070 8210
rect 20400 8205 20420 8225
rect 14115 8155 14135 8175
rect 20400 8155 20420 8175
rect 14115 8105 14135 8125
rect 14115 8055 14135 8075
rect 14115 8005 14135 8025
rect 14115 7955 14135 7975
rect 20400 8105 20420 8125
rect 20400 8055 20420 8075
rect 20400 8005 20420 8025
rect 20400 7955 20420 7975
rect 11230 7860 11250 7880
rect 11230 7810 11250 7830
rect 11230 7760 11250 7780
rect 11230 7710 11250 7730
rect 11230 7660 11250 7680
rect 9690 7585 9710 7605
rect 9690 7535 9710 7555
rect 9745 7585 9765 7605
rect 9745 7535 9765 7555
rect 9800 7585 9820 7605
rect 9800 7535 9820 7555
rect 9855 7585 9875 7605
rect 9855 7535 9875 7555
rect 9910 7585 9930 7605
rect 9910 7535 9930 7555
rect 9965 7585 9985 7605
rect 9965 7535 9985 7555
rect 10020 7585 10040 7605
rect 10020 7535 10040 7555
rect 10075 7585 10095 7605
rect 10075 7535 10095 7555
rect 10130 7585 10150 7605
rect 10130 7535 10150 7555
rect 10185 7585 10205 7605
rect 10185 7535 10205 7555
rect 10240 7585 10260 7605
rect 10240 7535 10260 7555
rect 10295 7585 10315 7605
rect 10295 7535 10315 7555
rect 10350 7585 10370 7605
rect 10350 7535 10370 7555
rect 10405 7585 10425 7605
rect 10405 7535 10425 7555
rect 10460 7585 10480 7605
rect 10460 7535 10480 7555
rect 10515 7585 10535 7605
rect 10515 7535 10535 7555
rect 10570 7585 10590 7605
rect 10570 7535 10590 7555
rect 10625 7585 10645 7605
rect 10625 7535 10645 7555
rect 10680 7585 10700 7605
rect 10680 7535 10700 7555
rect 10735 7585 10755 7605
rect 10735 7535 10755 7555
rect 10790 7585 10810 7605
rect 10790 7535 10810 7555
rect 10845 7585 10865 7605
rect 10845 7535 10865 7555
rect 10900 7585 10920 7605
rect 10900 7535 10920 7555
rect 11230 7610 11250 7630
rect 11230 7560 11250 7580
rect 11230 7510 11250 7530
rect 11290 7860 11310 7880
rect 11290 7810 11310 7830
rect 11290 7760 11310 7780
rect 11290 7710 11310 7730
rect 11290 7660 11310 7680
rect 11290 7610 11310 7630
rect 11290 7560 11310 7580
rect 11290 7510 11310 7530
rect 11350 7860 11370 7880
rect 11350 7810 11370 7830
rect 11350 7760 11370 7780
rect 11350 7710 11370 7730
rect 11350 7660 11370 7680
rect 11350 7610 11370 7630
rect 11350 7560 11370 7580
rect 11350 7510 11370 7530
rect 11410 7860 11430 7880
rect 11410 7810 11430 7830
rect 11410 7760 11430 7780
rect 11410 7710 11430 7730
rect 11410 7660 11430 7680
rect 11410 7610 11430 7630
rect 11410 7560 11430 7580
rect 11410 7510 11430 7530
rect 11470 7860 11490 7880
rect 11470 7810 11490 7830
rect 11470 7760 11490 7780
rect 11470 7710 11490 7730
rect 11470 7660 11490 7680
rect 11470 7610 11490 7630
rect 11470 7560 11490 7580
rect 11470 7510 11490 7530
rect 11530 7860 11550 7880
rect 11530 7810 11550 7830
rect 11530 7760 11550 7780
rect 11530 7710 11550 7730
rect 11530 7660 11550 7680
rect 11530 7610 11550 7630
rect 11530 7560 11550 7580
rect 11530 7510 11550 7530
rect 11590 7860 11610 7880
rect 11590 7810 11610 7830
rect 11590 7760 11610 7780
rect 11590 7710 11610 7730
rect 11590 7660 11610 7680
rect 11590 7610 11610 7630
rect 11590 7560 11610 7580
rect 11590 7510 11610 7530
rect 11650 7860 11670 7880
rect 11650 7810 11670 7830
rect 11650 7760 11670 7780
rect 11650 7710 11670 7730
rect 11650 7660 11670 7680
rect 11650 7610 11670 7630
rect 11650 7560 11670 7580
rect 11650 7510 11670 7530
rect 11710 7860 11730 7880
rect 11710 7810 11730 7830
rect 11710 7760 11730 7780
rect 11710 7710 11730 7730
rect 11710 7660 11730 7680
rect 11710 7610 11730 7630
rect 11710 7560 11730 7580
rect 11710 7510 11730 7530
rect 11770 7860 11790 7880
rect 11770 7810 11790 7830
rect 11770 7760 11790 7780
rect 11770 7710 11790 7730
rect 11770 7660 11790 7680
rect 11770 7610 11790 7630
rect 11770 7560 11790 7580
rect 11770 7510 11790 7530
rect 11830 7860 11850 7880
rect 11830 7810 11850 7830
rect 11830 7760 11850 7780
rect 11830 7710 11850 7730
rect 11830 7660 11850 7680
rect 11830 7610 11850 7630
rect 11830 7560 11850 7580
rect 11830 7510 11850 7530
rect 11890 7860 11910 7880
rect 11890 7810 11910 7830
rect 11890 7760 11910 7780
rect 11890 7710 11910 7730
rect 11890 7660 11910 7680
rect 11890 7610 11910 7630
rect 11890 7560 11910 7580
rect 11890 7510 11910 7530
rect 11950 7860 11970 7880
rect 11950 7810 11970 7830
rect 11950 7760 11970 7780
rect 11950 7710 11970 7730
rect 11950 7660 11970 7680
rect 11950 7610 11970 7630
rect 11950 7560 11970 7580
rect 11950 7510 11970 7530
rect 12010 7860 12030 7880
rect 12010 7810 12030 7830
rect 12010 7760 12030 7780
rect 12010 7710 12030 7730
rect 12010 7660 12030 7680
rect 12010 7610 12030 7630
rect 12010 7560 12030 7580
rect 12010 7510 12030 7530
rect 12070 7860 12090 7880
rect 12070 7810 12090 7830
rect 12070 7760 12090 7780
rect 12070 7710 12090 7730
rect 12070 7660 12090 7680
rect 12070 7610 12090 7630
rect 12070 7560 12090 7580
rect 12070 7510 12090 7530
rect 12130 7860 12150 7880
rect 12130 7810 12150 7830
rect 12130 7760 12150 7780
rect 12130 7710 12150 7730
rect 12130 7660 12150 7680
rect 12130 7610 12150 7630
rect 12130 7560 12150 7580
rect 12130 7510 12150 7530
rect 12190 7860 12210 7880
rect 12190 7810 12210 7830
rect 12190 7760 12210 7780
rect 12190 7710 12210 7730
rect 12190 7660 12210 7680
rect 12190 7610 12210 7630
rect 12190 7560 12210 7580
rect 12190 7510 12210 7530
rect 12250 7860 12270 7880
rect 12250 7810 12270 7830
rect 12250 7760 12270 7780
rect 12250 7710 12270 7730
rect 12250 7660 12270 7680
rect 12250 7610 12270 7630
rect 12250 7560 12270 7580
rect 12250 7510 12270 7530
rect 12310 7860 12330 7880
rect 12310 7810 12330 7830
rect 12310 7760 12330 7780
rect 12310 7710 12330 7730
rect 12310 7660 12330 7680
rect 12310 7610 12330 7630
rect 12310 7560 12330 7580
rect 12310 7510 12330 7530
rect 12370 7860 12390 7880
rect 12370 7810 12390 7830
rect 12370 7760 12390 7780
rect 12370 7710 12390 7730
rect 12370 7660 12390 7680
rect 12370 7610 12390 7630
rect 12370 7560 12390 7580
rect 12370 7510 12390 7530
rect 12430 7860 12450 7880
rect 12430 7810 12450 7830
rect 12430 7760 12450 7780
rect 12430 7710 12450 7730
rect 12430 7660 12450 7680
rect 12430 7610 12450 7630
rect 12430 7560 12450 7580
rect 12430 7510 12450 7530
rect 12490 7860 12510 7880
rect 12490 7810 12510 7830
rect 12490 7760 12510 7780
rect 12490 7710 12510 7730
rect 12490 7660 12510 7680
rect 12490 7610 12510 7630
rect 12490 7560 12510 7580
rect 12490 7510 12510 7530
rect 20455 8205 20475 8225
rect 20455 8155 20475 8175
rect 20455 8105 20475 8125
rect 20455 8055 20475 8075
rect 20455 8005 20475 8025
rect 20455 7955 20475 7975
rect 20510 8205 20530 8225
rect 20510 8155 20530 8175
rect 20510 8105 20530 8125
rect 20510 8055 20530 8075
rect 20510 8005 20530 8025
rect 20510 7955 20530 7975
rect 20565 8205 20585 8225
rect 20565 8155 20585 8175
rect 20565 8105 20585 8125
rect 20565 8055 20585 8075
rect 20565 8005 20585 8025
rect 20565 7955 20585 7975
rect 20620 8205 20640 8225
rect 20620 8155 20640 8175
rect 20620 8105 20640 8125
rect 20620 8055 20640 8075
rect 20620 8005 20640 8025
rect 20620 7955 20640 7975
rect 20675 8205 20695 8225
rect 20675 8155 20695 8175
rect 20675 8105 20695 8125
rect 20675 8055 20695 8075
rect 20675 8005 20695 8025
rect 20675 7955 20695 7975
rect 20730 8205 20750 8225
rect 20730 8155 20750 8175
rect 20730 8105 20750 8125
rect 20730 8055 20750 8075
rect 20730 8005 20750 8025
rect 20730 7955 20750 7975
rect 20785 8205 20805 8225
rect 20785 8155 20805 8175
rect 20785 8105 20805 8125
rect 20785 8055 20805 8075
rect 20785 8005 20805 8025
rect 20785 7955 20805 7975
rect 20840 8205 20860 8225
rect 20840 8155 20860 8175
rect 20840 8105 20860 8125
rect 20840 8055 20860 8075
rect 20840 8005 20860 8025
rect 20840 7955 20860 7975
rect 20895 8205 20915 8225
rect 20895 8155 20915 8175
rect 20895 8105 20915 8125
rect 20895 8055 20915 8075
rect 20895 8005 20915 8025
rect 20895 7955 20915 7975
rect 20950 8205 20970 8225
rect 20950 8155 20970 8175
rect 20950 8105 20970 8125
rect 20950 8055 20970 8075
rect 20950 8005 20970 8025
rect 20950 7955 20970 7975
rect 21005 8205 21025 8225
rect 21005 8155 21025 8175
rect 21005 8105 21025 8125
rect 21005 8055 21025 8075
rect 21005 8005 21025 8025
rect 21005 7955 21025 7975
rect 21060 8205 21080 8225
rect 21060 8155 21080 8175
rect 21060 8105 21080 8125
rect 21060 8055 21080 8075
rect 21060 8005 21080 8025
rect 21060 7955 21080 7975
rect 21115 8205 21135 8225
rect 21115 8155 21135 8175
rect 21115 8105 21135 8125
rect 21115 8055 21135 8075
rect 21115 8005 21135 8025
rect 21115 7955 21135 7975
rect 21170 8205 21190 8225
rect 21170 8155 21190 8175
rect 21170 8105 21190 8125
rect 21170 8055 21190 8075
rect 21170 8005 21190 8025
rect 21170 7955 21190 7975
rect 21225 8205 21245 8225
rect 21225 8155 21245 8175
rect 21225 8105 21245 8125
rect 21225 8055 21245 8075
rect 21225 8005 21245 8025
rect 21225 7955 21245 7975
rect 21280 8205 21300 8225
rect 21280 8155 21300 8175
rect 21280 8105 21300 8125
rect 21280 8055 21300 8075
rect 21280 8005 21300 8025
rect 21280 7955 21300 7975
rect 21335 8205 21355 8225
rect 21335 8155 21355 8175
rect 21335 8105 21355 8125
rect 21335 8055 21355 8075
rect 21335 8005 21355 8025
rect 21335 7955 21355 7975
rect 21390 8205 21410 8225
rect 21390 8155 21410 8175
rect 21390 8105 21410 8125
rect 21390 8055 21410 8075
rect 21390 8005 21410 8025
rect 21390 7955 21410 7975
rect 21445 8205 21465 8225
rect 21445 8155 21465 8175
rect 21445 8105 21465 8125
rect 21445 8055 21465 8075
rect 21445 8005 21465 8025
rect 21445 7955 21465 7975
rect 21500 8205 21520 8225
rect 21500 8155 21520 8175
rect 21500 8105 21520 8125
rect 21500 8055 21520 8075
rect 21500 8005 21520 8025
rect 21500 7955 21520 7975
rect 21555 8205 21575 8225
rect 21555 8155 21575 8175
rect 21555 8105 21575 8125
rect 21555 8055 21575 8075
rect 21555 8005 21575 8025
rect 21555 7955 21575 7975
rect 21610 8205 21630 8225
rect 21610 8155 21630 8175
rect 21610 8105 21630 8125
rect 21610 8055 21630 8075
rect 21610 8005 21630 8025
rect 21610 7955 21630 7975
rect 12550 7860 12570 7880
rect 18730 7860 18750 7880
rect 12550 7810 12570 7830
rect 12550 7760 12570 7780
rect 12550 7710 12570 7730
rect 18730 7810 18750 7830
rect 18730 7760 18750 7780
rect 18730 7710 18750 7730
rect 12550 7660 12570 7680
rect 18730 7660 18750 7680
rect 12550 7610 12570 7630
rect 12550 7560 12570 7580
rect 12550 7510 12570 7530
rect 12905 7585 12925 7605
rect 12905 7535 12925 7555
rect 12960 7585 12980 7605
rect 12960 7535 12980 7555
rect 13015 7585 13035 7605
rect 13015 7535 13035 7555
rect 13070 7585 13090 7605
rect 13070 7535 13090 7555
rect 13125 7585 13145 7605
rect 13125 7535 13145 7555
rect 13180 7585 13200 7605
rect 13180 7535 13200 7555
rect 13235 7585 13255 7605
rect 13235 7535 13255 7555
rect 13290 7585 13310 7605
rect 13290 7535 13310 7555
rect 13345 7585 13365 7605
rect 13345 7535 13365 7555
rect 13400 7585 13420 7605
rect 13400 7535 13420 7555
rect 13455 7585 13475 7605
rect 13455 7535 13475 7555
rect 13510 7585 13530 7605
rect 13510 7535 13530 7555
rect 13565 7585 13585 7605
rect 13565 7535 13585 7555
rect 13620 7585 13640 7605
rect 13620 7535 13640 7555
rect 13675 7585 13695 7605
rect 13675 7535 13695 7555
rect 13730 7585 13750 7605
rect 13730 7535 13750 7555
rect 13785 7585 13805 7605
rect 13785 7535 13805 7555
rect 13840 7585 13860 7605
rect 13840 7535 13860 7555
rect 13895 7585 13915 7605
rect 13895 7535 13915 7555
rect 13950 7585 13970 7605
rect 13950 7535 13970 7555
rect 14005 7585 14025 7605
rect 14005 7535 14025 7555
rect 14060 7585 14080 7605
rect 14060 7535 14080 7555
rect 14115 7585 14135 7605
rect 14115 7535 14135 7555
rect 17190 7585 17210 7605
rect 17190 7535 17210 7555
rect 17245 7585 17265 7605
rect 17245 7535 17265 7555
rect 17300 7585 17320 7605
rect 17300 7535 17320 7555
rect 17355 7585 17375 7605
rect 17355 7535 17375 7555
rect 17410 7585 17430 7605
rect 17410 7535 17430 7555
rect 17465 7585 17485 7605
rect 17465 7535 17485 7555
rect 17520 7585 17540 7605
rect 17520 7535 17540 7555
rect 17575 7585 17595 7605
rect 17575 7535 17595 7555
rect 17630 7585 17650 7605
rect 17630 7535 17650 7555
rect 17685 7585 17705 7605
rect 17685 7535 17705 7555
rect 17740 7585 17760 7605
rect 17740 7535 17760 7555
rect 17795 7585 17815 7605
rect 17795 7535 17815 7555
rect 17850 7585 17870 7605
rect 17850 7535 17870 7555
rect 17905 7585 17925 7605
rect 17905 7535 17925 7555
rect 17960 7585 17980 7605
rect 17960 7535 17980 7555
rect 18015 7585 18035 7605
rect 18015 7535 18035 7555
rect 18070 7585 18090 7605
rect 18070 7535 18090 7555
rect 18125 7585 18145 7605
rect 18125 7535 18145 7555
rect 18180 7585 18200 7605
rect 18180 7535 18200 7555
rect 18235 7585 18255 7605
rect 18235 7535 18255 7555
rect 18290 7585 18310 7605
rect 18290 7535 18310 7555
rect 18345 7585 18365 7605
rect 18345 7535 18365 7555
rect 18400 7585 18420 7605
rect 18400 7535 18420 7555
rect 18730 7610 18750 7630
rect 18730 7560 18750 7580
rect 18730 7510 18750 7530
rect 18790 7860 18810 7880
rect 18790 7810 18810 7830
rect 18790 7760 18810 7780
rect 18790 7710 18810 7730
rect 18790 7660 18810 7680
rect 18790 7610 18810 7630
rect 18790 7560 18810 7580
rect 18790 7510 18810 7530
rect 18850 7860 18870 7880
rect 18850 7810 18870 7830
rect 18850 7760 18870 7780
rect 18850 7710 18870 7730
rect 18850 7660 18870 7680
rect 18850 7610 18870 7630
rect 18850 7560 18870 7580
rect 18850 7510 18870 7530
rect 18910 7860 18930 7880
rect 18910 7810 18930 7830
rect 18910 7760 18930 7780
rect 18910 7710 18930 7730
rect 18910 7660 18930 7680
rect 18910 7610 18930 7630
rect 18910 7560 18930 7580
rect 18910 7510 18930 7530
rect 18970 7860 18990 7880
rect 18970 7810 18990 7830
rect 18970 7760 18990 7780
rect 18970 7710 18990 7730
rect 18970 7660 18990 7680
rect 18970 7610 18990 7630
rect 18970 7560 18990 7580
rect 18970 7510 18990 7530
rect 19030 7860 19050 7880
rect 19030 7810 19050 7830
rect 19030 7760 19050 7780
rect 19030 7710 19050 7730
rect 19030 7660 19050 7680
rect 19030 7610 19050 7630
rect 19030 7560 19050 7580
rect 19030 7510 19050 7530
rect 19090 7860 19110 7880
rect 19090 7810 19110 7830
rect 19090 7760 19110 7780
rect 19090 7710 19110 7730
rect 19090 7660 19110 7680
rect 19090 7610 19110 7630
rect 19090 7560 19110 7580
rect 19090 7510 19110 7530
rect 19150 7860 19170 7880
rect 19150 7810 19170 7830
rect 19150 7760 19170 7780
rect 19150 7710 19170 7730
rect 19150 7660 19170 7680
rect 19150 7610 19170 7630
rect 19150 7560 19170 7580
rect 19150 7510 19170 7530
rect 19210 7860 19230 7880
rect 19210 7810 19230 7830
rect 19210 7760 19230 7780
rect 19210 7710 19230 7730
rect 19210 7660 19230 7680
rect 19210 7610 19230 7630
rect 19210 7560 19230 7580
rect 19210 7510 19230 7530
rect 19270 7860 19290 7880
rect 19270 7810 19290 7830
rect 19270 7760 19290 7780
rect 19270 7710 19290 7730
rect 19270 7660 19290 7680
rect 19270 7610 19290 7630
rect 19270 7560 19290 7580
rect 19270 7510 19290 7530
rect 19330 7860 19350 7880
rect 19330 7810 19350 7830
rect 19330 7760 19350 7780
rect 19330 7710 19350 7730
rect 19330 7660 19350 7680
rect 19330 7610 19350 7630
rect 19330 7560 19350 7580
rect 19330 7510 19350 7530
rect 19390 7860 19410 7880
rect 19390 7810 19410 7830
rect 19390 7760 19410 7780
rect 19390 7710 19410 7730
rect 19390 7660 19410 7680
rect 19390 7610 19410 7630
rect 19390 7560 19410 7580
rect 19390 7510 19410 7530
rect 19450 7860 19470 7880
rect 19450 7810 19470 7830
rect 19450 7760 19470 7780
rect 19450 7710 19470 7730
rect 19450 7660 19470 7680
rect 19450 7610 19470 7630
rect 19450 7560 19470 7580
rect 19450 7510 19470 7530
rect 19510 7860 19530 7880
rect 19510 7810 19530 7830
rect 19510 7760 19530 7780
rect 19510 7710 19530 7730
rect 19510 7660 19530 7680
rect 19510 7610 19530 7630
rect 19510 7560 19530 7580
rect 19510 7510 19530 7530
rect 19570 7860 19590 7880
rect 19570 7810 19590 7830
rect 19570 7760 19590 7780
rect 19570 7710 19590 7730
rect 19570 7660 19590 7680
rect 19570 7610 19590 7630
rect 19570 7560 19590 7580
rect 19570 7510 19590 7530
rect 19630 7860 19650 7880
rect 19630 7810 19650 7830
rect 19630 7760 19650 7780
rect 19630 7710 19650 7730
rect 19630 7660 19650 7680
rect 19630 7610 19650 7630
rect 19630 7560 19650 7580
rect 19630 7510 19650 7530
rect 19690 7860 19710 7880
rect 19690 7810 19710 7830
rect 19690 7760 19710 7780
rect 19690 7710 19710 7730
rect 19690 7660 19710 7680
rect 19690 7610 19710 7630
rect 19690 7560 19710 7580
rect 19690 7510 19710 7530
rect 19750 7860 19770 7880
rect 19750 7810 19770 7830
rect 19750 7760 19770 7780
rect 19750 7710 19770 7730
rect 19750 7660 19770 7680
rect 19750 7610 19770 7630
rect 19750 7560 19770 7580
rect 19750 7510 19770 7530
rect 19810 7860 19830 7880
rect 19810 7810 19830 7830
rect 19810 7760 19830 7780
rect 19810 7710 19830 7730
rect 19810 7660 19830 7680
rect 19810 7610 19830 7630
rect 19810 7560 19830 7580
rect 19810 7510 19830 7530
rect 19870 7860 19890 7880
rect 19870 7810 19890 7830
rect 19870 7760 19890 7780
rect 19870 7710 19890 7730
rect 19870 7660 19890 7680
rect 19870 7610 19890 7630
rect 19870 7560 19890 7580
rect 19870 7510 19890 7530
rect 19930 7860 19950 7880
rect 19930 7810 19950 7830
rect 19930 7760 19950 7780
rect 19930 7710 19950 7730
rect 19930 7660 19950 7680
rect 19930 7610 19950 7630
rect 19930 7560 19950 7580
rect 19930 7510 19950 7530
rect 19990 7860 20010 7880
rect 19990 7810 20010 7830
rect 19990 7760 20010 7780
rect 19990 7710 20010 7730
rect 19990 7660 20010 7680
rect 19990 7610 20010 7630
rect 19990 7560 20010 7580
rect 19990 7510 20010 7530
rect 20050 7860 20070 7880
rect 20050 7810 20070 7830
rect 20050 7760 20070 7780
rect 20050 7710 20070 7730
rect 20050 7660 20070 7680
rect 20050 7610 20070 7630
rect 20050 7560 20070 7580
rect 20050 7510 20070 7530
rect 20400 7585 20420 7605
rect 20400 7535 20420 7555
rect 20455 7585 20475 7605
rect 20455 7535 20475 7555
rect 20510 7585 20530 7605
rect 20510 7535 20530 7555
rect 20565 7585 20585 7605
rect 20565 7535 20585 7555
rect 20620 7585 20640 7605
rect 20620 7535 20640 7555
rect 20675 7585 20695 7605
rect 20675 7535 20695 7555
rect 20730 7585 20750 7605
rect 20730 7535 20750 7555
rect 20785 7585 20805 7605
rect 20785 7535 20805 7555
rect 20840 7585 20860 7605
rect 20840 7535 20860 7555
rect 20895 7585 20915 7605
rect 20895 7535 20915 7555
rect 20950 7585 20970 7605
rect 20950 7535 20970 7555
rect 21005 7585 21025 7605
rect 21005 7535 21025 7555
rect 21060 7585 21080 7605
rect 21060 7535 21080 7555
rect 21115 7585 21135 7605
rect 21115 7535 21135 7555
rect 21170 7585 21190 7605
rect 21170 7535 21190 7555
rect 21225 7585 21245 7605
rect 21225 7535 21245 7555
rect 21280 7585 21300 7605
rect 21280 7535 21300 7555
rect 21335 7585 21355 7605
rect 21335 7535 21355 7555
rect 21390 7585 21410 7605
rect 21390 7535 21410 7555
rect 21445 7585 21465 7605
rect 21445 7535 21465 7555
rect 21500 7585 21520 7605
rect 21500 7535 21520 7555
rect 21555 7585 21575 7605
rect 21555 7535 21575 7555
rect 21610 7585 21630 7605
rect 21610 7535 21630 7555
rect 9690 7135 9710 7155
rect 9690 7085 9710 7105
rect 9690 7035 9710 7055
rect 9745 7135 9765 7155
rect 9745 7085 9765 7105
rect 9745 7035 9765 7055
rect 9800 7135 9820 7155
rect 9800 7085 9820 7105
rect 9800 7035 9820 7055
rect 9855 7135 9875 7155
rect 9855 7085 9875 7105
rect 9855 7035 9875 7055
rect 9910 7135 9930 7155
rect 9910 7085 9930 7105
rect 9910 7035 9930 7055
rect 9965 7135 9985 7155
rect 9965 7085 9985 7105
rect 9965 7035 9985 7055
rect 10020 7135 10040 7155
rect 10020 7085 10040 7105
rect 10020 7035 10040 7055
rect 10075 7135 10095 7155
rect 10075 7085 10095 7105
rect 10075 7035 10095 7055
rect 10130 7135 10150 7155
rect 10130 7085 10150 7105
rect 10130 7035 10150 7055
rect 10185 7135 10205 7155
rect 10185 7085 10205 7105
rect 10185 7035 10205 7055
rect 10240 7135 10260 7155
rect 10240 7085 10260 7105
rect 10240 7035 10260 7055
rect 10295 7135 10315 7155
rect 10295 7085 10315 7105
rect 10295 7035 10315 7055
rect 10350 7135 10370 7155
rect 10350 7085 10370 7105
rect 10350 7035 10370 7055
rect 10405 7135 10425 7155
rect 10405 7085 10425 7105
rect 10405 7035 10425 7055
rect 10460 7135 10480 7155
rect 10460 7085 10480 7105
rect 10460 7035 10480 7055
rect 10515 7135 10535 7155
rect 10515 7085 10535 7105
rect 10515 7035 10535 7055
rect 10570 7135 10590 7155
rect 10570 7085 10590 7105
rect 10570 7035 10590 7055
rect 10625 7135 10645 7155
rect 10625 7085 10645 7105
rect 10625 7035 10645 7055
rect 10680 7135 10700 7155
rect 10680 7085 10700 7105
rect 10680 7035 10700 7055
rect 10735 7135 10755 7155
rect 10735 7085 10755 7105
rect 10735 7035 10755 7055
rect 10790 7135 10810 7155
rect 10790 7085 10810 7105
rect 10790 7035 10810 7055
rect 10845 7135 10865 7155
rect 10845 7085 10865 7105
rect 10845 7035 10865 7055
rect 10900 7135 10920 7155
rect 12905 7135 12925 7155
rect 10900 7085 10920 7105
rect 10900 7035 10920 7055
rect 11285 7095 11305 7115
rect 11285 7045 11305 7065
rect 11285 6995 11305 7015
rect 11340 7095 11360 7115
rect 11340 7045 11360 7065
rect 11340 6995 11360 7015
rect 11395 7095 11415 7115
rect 11395 7045 11415 7065
rect 11395 6995 11415 7015
rect 11450 7095 11470 7115
rect 11450 7045 11470 7065
rect 11450 6995 11470 7015
rect 11505 7095 11525 7115
rect 11505 7045 11525 7065
rect 11505 6995 11525 7015
rect 11560 7095 11580 7115
rect 11560 7045 11580 7065
rect 11560 6995 11580 7015
rect 11615 7095 11635 7115
rect 11615 7045 11635 7065
rect 11615 6995 11635 7015
rect 11670 7095 11690 7115
rect 11670 7045 11690 7065
rect 11670 6995 11690 7015
rect 11725 7095 11745 7115
rect 11725 7045 11745 7065
rect 11725 6995 11745 7015
rect 11780 7095 11800 7115
rect 11780 7045 11800 7065
rect 11780 6995 11800 7015
rect 11835 7095 11855 7115
rect 11835 7045 11855 7065
rect 11835 6995 11855 7015
rect 11890 7095 11910 7115
rect 11890 7045 11910 7065
rect 11890 6995 11910 7015
rect 11945 7095 11965 7115
rect 11945 7045 11965 7065
rect 11945 6995 11965 7015
rect 12000 7095 12020 7115
rect 12000 7045 12020 7065
rect 12000 6995 12020 7015
rect 12055 7095 12075 7115
rect 12055 7045 12075 7065
rect 12055 6995 12075 7015
rect 12110 7095 12130 7115
rect 12110 7045 12130 7065
rect 12110 6995 12130 7015
rect 12165 7095 12185 7115
rect 12165 7045 12185 7065
rect 12165 6995 12185 7015
rect 12220 7095 12240 7115
rect 12220 7045 12240 7065
rect 12220 6995 12240 7015
rect 12275 7095 12295 7115
rect 12275 7045 12295 7065
rect 12275 6995 12295 7015
rect 12330 7095 12350 7115
rect 12330 7045 12350 7065
rect 12330 6995 12350 7015
rect 12385 7095 12405 7115
rect 12385 7045 12405 7065
rect 12385 6995 12405 7015
rect 12440 7095 12460 7115
rect 12440 7045 12460 7065
rect 12440 6995 12460 7015
rect 12495 7095 12515 7115
rect 12495 7045 12515 7065
rect 12905 7085 12925 7105
rect 12905 7035 12925 7055
rect 12960 7135 12980 7155
rect 12960 7085 12980 7105
rect 12960 7035 12980 7055
rect 13015 7135 13035 7155
rect 13015 7085 13035 7105
rect 13015 7035 13035 7055
rect 13070 7135 13090 7155
rect 13070 7085 13090 7105
rect 13070 7035 13090 7055
rect 13125 7135 13145 7155
rect 13125 7085 13145 7105
rect 13125 7035 13145 7055
rect 13180 7135 13200 7155
rect 13180 7085 13200 7105
rect 13180 7035 13200 7055
rect 13235 7135 13255 7155
rect 13235 7085 13255 7105
rect 13235 7035 13255 7055
rect 13290 7135 13310 7155
rect 13290 7085 13310 7105
rect 13290 7035 13310 7055
rect 13345 7135 13365 7155
rect 13345 7085 13365 7105
rect 13345 7035 13365 7055
rect 13400 7135 13420 7155
rect 13400 7085 13420 7105
rect 13400 7035 13420 7055
rect 13455 7135 13475 7155
rect 13455 7085 13475 7105
rect 13455 7035 13475 7055
rect 13510 7135 13530 7155
rect 13510 7085 13530 7105
rect 13510 7035 13530 7055
rect 13565 7135 13585 7155
rect 13565 7085 13585 7105
rect 13565 7035 13585 7055
rect 13620 7135 13640 7155
rect 13620 7085 13640 7105
rect 13620 7035 13640 7055
rect 13675 7135 13695 7155
rect 13675 7085 13695 7105
rect 13675 7035 13695 7055
rect 13730 7135 13750 7155
rect 13730 7085 13750 7105
rect 13730 7035 13750 7055
rect 13785 7135 13805 7155
rect 13785 7085 13805 7105
rect 13785 7035 13805 7055
rect 13840 7135 13860 7155
rect 13840 7085 13860 7105
rect 13840 7035 13860 7055
rect 13895 7135 13915 7155
rect 13895 7085 13915 7105
rect 13895 7035 13915 7055
rect 13950 7135 13970 7155
rect 13950 7085 13970 7105
rect 13950 7035 13970 7055
rect 14005 7135 14025 7155
rect 14005 7085 14025 7105
rect 14005 7035 14025 7055
rect 14060 7135 14080 7155
rect 14060 7085 14080 7105
rect 14060 7035 14080 7055
rect 14115 7135 14135 7155
rect 14115 7085 14135 7105
rect 14115 7035 14135 7055
rect 17190 7135 17210 7155
rect 17190 7085 17210 7105
rect 17190 7035 17210 7055
rect 17245 7135 17265 7155
rect 17245 7085 17265 7105
rect 17245 7035 17265 7055
rect 17300 7135 17320 7155
rect 17300 7085 17320 7105
rect 17300 7035 17320 7055
rect 17355 7135 17375 7155
rect 17355 7085 17375 7105
rect 17355 7035 17375 7055
rect 17410 7135 17430 7155
rect 17410 7085 17430 7105
rect 17410 7035 17430 7055
rect 17465 7135 17485 7155
rect 17465 7085 17485 7105
rect 17465 7035 17485 7055
rect 17520 7135 17540 7155
rect 17520 7085 17540 7105
rect 17520 7035 17540 7055
rect 17575 7135 17595 7155
rect 17575 7085 17595 7105
rect 17575 7035 17595 7055
rect 17630 7135 17650 7155
rect 17630 7085 17650 7105
rect 17630 7035 17650 7055
rect 17685 7135 17705 7155
rect 17685 7085 17705 7105
rect 17685 7035 17705 7055
rect 17740 7135 17760 7155
rect 17740 7085 17760 7105
rect 17740 7035 17760 7055
rect 17795 7135 17815 7155
rect 17795 7085 17815 7105
rect 17795 7035 17815 7055
rect 17850 7135 17870 7155
rect 17850 7085 17870 7105
rect 17850 7035 17870 7055
rect 17905 7135 17925 7155
rect 17905 7085 17925 7105
rect 17905 7035 17925 7055
rect 17960 7135 17980 7155
rect 17960 7085 17980 7105
rect 17960 7035 17980 7055
rect 18015 7135 18035 7155
rect 18015 7085 18035 7105
rect 18015 7035 18035 7055
rect 18070 7135 18090 7155
rect 18070 7085 18090 7105
rect 18070 7035 18090 7055
rect 18125 7135 18145 7155
rect 18125 7085 18145 7105
rect 18125 7035 18145 7055
rect 18180 7135 18200 7155
rect 18180 7085 18200 7105
rect 18180 7035 18200 7055
rect 18235 7135 18255 7155
rect 18235 7085 18255 7105
rect 18235 7035 18255 7055
rect 18290 7135 18310 7155
rect 18290 7085 18310 7105
rect 18290 7035 18310 7055
rect 18345 7135 18365 7155
rect 18345 7085 18365 7105
rect 18345 7035 18365 7055
rect 18400 7135 18420 7155
rect 20400 7135 20420 7155
rect 18400 7085 18420 7105
rect 18400 7035 18420 7055
rect 18785 7095 18805 7115
rect 18785 7045 18805 7065
rect 12495 6995 12515 7015
rect 18785 6995 18805 7015
rect 18840 7095 18860 7115
rect 18840 7045 18860 7065
rect 18840 6995 18860 7015
rect 18895 7095 18915 7115
rect 18895 7045 18915 7065
rect 18895 6995 18915 7015
rect 18950 7095 18970 7115
rect 18950 7045 18970 7065
rect 18950 6995 18970 7015
rect 19005 7095 19025 7115
rect 19005 7045 19025 7065
rect 19005 6995 19025 7015
rect 19060 7095 19080 7115
rect 19060 7045 19080 7065
rect 19060 6995 19080 7015
rect 19115 7095 19135 7115
rect 19115 7045 19135 7065
rect 19115 6995 19135 7015
rect 19170 7095 19190 7115
rect 19170 7045 19190 7065
rect 19170 6995 19190 7015
rect 19225 7095 19245 7115
rect 19225 7045 19245 7065
rect 19225 6995 19245 7015
rect 19280 7095 19300 7115
rect 19280 7045 19300 7065
rect 19280 6995 19300 7015
rect 19335 7095 19355 7115
rect 19335 7045 19355 7065
rect 19335 6995 19355 7015
rect 19390 7095 19410 7115
rect 19390 7045 19410 7065
rect 19390 6995 19410 7015
rect 19445 7095 19465 7115
rect 19445 7045 19465 7065
rect 19445 6995 19465 7015
rect 19500 7095 19520 7115
rect 19500 7045 19520 7065
rect 19500 6995 19520 7015
rect 19555 7095 19575 7115
rect 19555 7045 19575 7065
rect 19555 6995 19575 7015
rect 19610 7095 19630 7115
rect 19610 7045 19630 7065
rect 19610 6995 19630 7015
rect 19665 7095 19685 7115
rect 19665 7045 19685 7065
rect 19665 6995 19685 7015
rect 19720 7095 19740 7115
rect 19720 7045 19740 7065
rect 19720 6995 19740 7015
rect 19775 7095 19795 7115
rect 19775 7045 19795 7065
rect 19775 6995 19795 7015
rect 19830 7095 19850 7115
rect 19830 7045 19850 7065
rect 19830 6995 19850 7015
rect 19885 7095 19905 7115
rect 19885 7045 19905 7065
rect 19885 6995 19905 7015
rect 19940 7095 19960 7115
rect 19940 7045 19960 7065
rect 19940 6995 19960 7015
rect 19995 7095 20015 7115
rect 19995 7045 20015 7065
rect 20400 7085 20420 7105
rect 20400 7035 20420 7055
rect 20455 7135 20475 7155
rect 20455 7085 20475 7105
rect 20455 7035 20475 7055
rect 20510 7135 20530 7155
rect 20510 7085 20530 7105
rect 20510 7035 20530 7055
rect 20565 7135 20585 7155
rect 20565 7085 20585 7105
rect 20565 7035 20585 7055
rect 20620 7135 20640 7155
rect 20620 7085 20640 7105
rect 20620 7035 20640 7055
rect 20675 7135 20695 7155
rect 20675 7085 20695 7105
rect 20675 7035 20695 7055
rect 20730 7135 20750 7155
rect 20730 7085 20750 7105
rect 20730 7035 20750 7055
rect 20785 7135 20805 7155
rect 20785 7085 20805 7105
rect 20785 7035 20805 7055
rect 20840 7135 20860 7155
rect 20840 7085 20860 7105
rect 20840 7035 20860 7055
rect 20895 7135 20915 7155
rect 20895 7085 20915 7105
rect 20895 7035 20915 7055
rect 20950 7135 20970 7155
rect 20950 7085 20970 7105
rect 20950 7035 20970 7055
rect 21005 7135 21025 7155
rect 21005 7085 21025 7105
rect 21005 7035 21025 7055
rect 21060 7135 21080 7155
rect 21060 7085 21080 7105
rect 21060 7035 21080 7055
rect 21115 7135 21135 7155
rect 21115 7085 21135 7105
rect 21115 7035 21135 7055
rect 21170 7135 21190 7155
rect 21170 7085 21190 7105
rect 21170 7035 21190 7055
rect 21225 7135 21245 7155
rect 21225 7085 21245 7105
rect 21225 7035 21245 7055
rect 21280 7135 21300 7155
rect 21280 7085 21300 7105
rect 21280 7035 21300 7055
rect 21335 7135 21355 7155
rect 21335 7085 21355 7105
rect 21335 7035 21355 7055
rect 21390 7135 21410 7155
rect 21390 7085 21410 7105
rect 21390 7035 21410 7055
rect 21445 7135 21465 7155
rect 21445 7085 21465 7105
rect 21445 7035 21465 7055
rect 21500 7135 21520 7155
rect 21500 7085 21520 7105
rect 21500 7035 21520 7055
rect 21555 7135 21575 7155
rect 21555 7085 21575 7105
rect 21555 7035 21575 7055
rect 21610 7135 21630 7155
rect 21610 7085 21630 7105
rect 21610 7035 21630 7055
rect 19995 6995 20015 7015
rect 20500 6820 20520 6840
rect 20500 6770 20520 6790
rect 20500 6720 20520 6740
rect 20555 6820 20575 6840
rect 20555 6770 20575 6790
rect 20555 6720 20575 6740
rect 20610 6820 20630 6840
rect 20610 6770 20630 6790
rect 20610 6720 20630 6740
rect 20665 6820 20685 6840
rect 20665 6770 20685 6790
rect 20665 6720 20685 6740
rect 20720 6820 20740 6840
rect 20720 6770 20740 6790
rect 20720 6720 20740 6740
rect 20775 6820 20795 6840
rect 20775 6770 20795 6790
rect 20775 6720 20795 6740
rect 20830 6820 20850 6840
rect 20830 6770 20850 6790
rect 20830 6720 20850 6740
rect 11040 6630 11060 6650
rect 11040 6580 11060 6600
rect 11040 6530 11060 6550
rect 11095 6630 11115 6650
rect 11095 6580 11115 6600
rect 11095 6530 11115 6550
rect 11150 6630 11170 6650
rect 11150 6580 11170 6600
rect 11150 6530 11170 6550
rect 11205 6630 11225 6650
rect 11205 6580 11225 6600
rect 11205 6530 11225 6550
rect 11260 6630 11280 6650
rect 11260 6580 11280 6600
rect 11260 6530 11280 6550
rect 11315 6630 11335 6650
rect 11315 6580 11335 6600
rect 11315 6530 11335 6550
rect 11370 6630 11390 6650
rect 11370 6580 11390 6600
rect 11370 6530 11390 6550
rect 11425 6630 11445 6650
rect 11425 6580 11445 6600
rect 11425 6530 11445 6550
rect 11480 6630 11500 6650
rect 11480 6580 11500 6600
rect 11480 6530 11500 6550
rect 11535 6630 11555 6650
rect 11535 6580 11555 6600
rect 11535 6530 11555 6550
rect 11590 6630 11610 6650
rect 11590 6580 11610 6600
rect 11590 6530 11610 6550
rect 11645 6630 11665 6650
rect 11645 6580 11665 6600
rect 11645 6530 11665 6550
rect 11700 6630 11720 6650
rect 11780 6630 11800 6650
rect 11700 6580 11720 6600
rect 11780 6580 11800 6600
rect 11700 6530 11720 6550
rect 11780 6530 11800 6550
rect 11835 6630 11855 6650
rect 11835 6580 11855 6600
rect 11835 6530 11855 6550
rect 11890 6630 11910 6650
rect 11890 6580 11910 6600
rect 11890 6530 11910 6550
rect 11945 6630 11965 6650
rect 11945 6580 11965 6600
rect 11945 6530 11965 6550
rect 12000 6630 12020 6650
rect 12080 6630 12100 6650
rect 12000 6580 12020 6600
rect 12080 6580 12100 6600
rect 12000 6530 12020 6550
rect 12080 6530 12100 6550
rect 12135 6630 12155 6650
rect 12135 6580 12155 6600
rect 12135 6530 12155 6550
rect 12190 6630 12210 6650
rect 12190 6580 12210 6600
rect 12190 6530 12210 6550
rect 12245 6630 12265 6650
rect 12245 6580 12265 6600
rect 12245 6530 12265 6550
rect 12300 6630 12320 6650
rect 12300 6580 12320 6600
rect 12300 6530 12320 6550
rect 12355 6630 12375 6650
rect 12355 6580 12375 6600
rect 12355 6530 12375 6550
rect 12410 6630 12430 6650
rect 12410 6580 12430 6600
rect 12410 6530 12430 6550
rect 12465 6630 12485 6650
rect 12465 6580 12485 6600
rect 12465 6530 12485 6550
rect 12520 6630 12540 6650
rect 12520 6580 12540 6600
rect 12520 6530 12540 6550
rect 12575 6630 12595 6650
rect 12575 6580 12595 6600
rect 12575 6530 12595 6550
rect 12630 6630 12650 6650
rect 12630 6580 12650 6600
rect 12630 6530 12650 6550
rect 12685 6630 12705 6650
rect 12685 6580 12705 6600
rect 12685 6530 12705 6550
rect 12740 6630 12760 6650
rect 12740 6580 12760 6600
rect 12740 6530 12760 6550
rect 18540 6630 18560 6650
rect 18540 6580 18560 6600
rect 18540 6530 18560 6550
rect 18595 6630 18615 6650
rect 18595 6580 18615 6600
rect 18595 6530 18615 6550
rect 18650 6630 18670 6650
rect 18650 6580 18670 6600
rect 18650 6530 18670 6550
rect 18705 6630 18725 6650
rect 18705 6580 18725 6600
rect 18705 6530 18725 6550
rect 18760 6630 18780 6650
rect 18760 6580 18780 6600
rect 18760 6530 18780 6550
rect 18815 6630 18835 6650
rect 18815 6580 18835 6600
rect 18815 6530 18835 6550
rect 18870 6630 18890 6650
rect 18870 6580 18890 6600
rect 18870 6530 18890 6550
rect 18925 6630 18945 6650
rect 18925 6580 18945 6600
rect 18925 6530 18945 6550
rect 18980 6630 19000 6650
rect 18980 6580 19000 6600
rect 18980 6530 19000 6550
rect 19035 6630 19055 6650
rect 19035 6580 19055 6600
rect 19035 6530 19055 6550
rect 19090 6630 19110 6650
rect 19090 6580 19110 6600
rect 19090 6530 19110 6550
rect 19145 6630 19165 6650
rect 19145 6580 19165 6600
rect 19145 6530 19165 6550
rect 19200 6630 19220 6650
rect 19280 6630 19300 6650
rect 19200 6580 19220 6600
rect 19280 6580 19300 6600
rect 19200 6530 19220 6550
rect 19280 6530 19300 6550
rect 19335 6630 19355 6650
rect 19335 6580 19355 6600
rect 19335 6530 19355 6550
rect 19390 6630 19410 6650
rect 19390 6580 19410 6600
rect 19390 6530 19410 6550
rect 19445 6630 19465 6650
rect 19445 6580 19465 6600
rect 19445 6530 19465 6550
rect 19500 6630 19520 6650
rect 19580 6630 19600 6650
rect 19500 6580 19520 6600
rect 19580 6580 19600 6600
rect 19500 6530 19520 6550
rect 19580 6530 19600 6550
rect 19635 6630 19655 6650
rect 19635 6580 19655 6600
rect 19635 6530 19655 6550
rect 19690 6630 19710 6650
rect 19690 6580 19710 6600
rect 19690 6530 19710 6550
rect 19745 6630 19765 6650
rect 19745 6580 19765 6600
rect 19745 6530 19765 6550
rect 19800 6630 19820 6650
rect 19800 6580 19820 6600
rect 19800 6530 19820 6550
rect 19855 6630 19875 6650
rect 19855 6580 19875 6600
rect 19855 6530 19875 6550
rect 19910 6630 19930 6650
rect 19910 6580 19930 6600
rect 19910 6530 19930 6550
rect 19965 6630 19985 6650
rect 19965 6580 19985 6600
rect 19965 6530 19985 6550
rect 20020 6630 20040 6650
rect 20020 6580 20040 6600
rect 20020 6530 20040 6550
rect 20075 6630 20095 6650
rect 20075 6580 20095 6600
rect 20075 6530 20095 6550
rect 20130 6630 20150 6650
rect 20130 6580 20150 6600
rect 20130 6530 20150 6550
rect 20185 6630 20205 6650
rect 20185 6580 20205 6600
rect 20185 6530 20205 6550
rect 20240 6630 20260 6650
rect 20240 6580 20260 6600
rect 20240 6530 20260 6550
rect 20405 6485 20425 6505
rect 20405 6435 20425 6455
rect 20405 6385 20425 6405
rect 20460 6485 20480 6505
rect 20460 6435 20480 6455
rect 20460 6385 20480 6405
rect 20515 6485 20535 6505
rect 20515 6435 20535 6455
rect 20515 6385 20535 6405
rect 20570 6485 20590 6505
rect 20570 6435 20590 6455
rect 20570 6385 20590 6405
rect 20625 6485 20645 6505
rect 20705 6485 20725 6505
rect 20625 6435 20645 6455
rect 20705 6435 20725 6455
rect 20625 6385 20645 6405
rect 20705 6385 20725 6405
rect 20760 6485 20780 6505
rect 20760 6435 20780 6455
rect 20760 6385 20780 6405
rect 20815 6485 20835 6505
rect 20815 6435 20835 6455
rect 20815 6385 20835 6405
rect 20870 6485 20890 6505
rect 20870 6435 20890 6455
rect 20870 6385 20890 6405
rect 20925 6485 20945 6505
rect 20925 6435 20945 6455
rect 20925 6385 20945 6405
rect 9675 6250 9695 6270
rect 9675 6205 9695 6225
rect 9675 6160 9695 6180
rect 9675 6110 9695 6130
rect 9675 6065 9695 6085
rect 9675 6020 9695 6040
rect 9775 6250 9795 6270
rect 9775 6205 9795 6225
rect 9775 6160 9795 6180
rect 9775 6110 9795 6130
rect 9775 6065 9795 6085
rect 9775 6020 9795 6040
rect 9875 6250 9895 6270
rect 9875 6205 9895 6225
rect 9875 6160 9895 6180
rect 9875 6110 9895 6130
rect 9875 6065 9895 6085
rect 9875 6020 9895 6040
rect 9975 6250 9995 6270
rect 9975 6205 9995 6225
rect 9975 6160 9995 6180
rect 9975 6110 9995 6130
rect 9975 6065 9995 6085
rect 9975 6020 9995 6040
rect 10075 6250 10095 6270
rect 10075 6205 10095 6225
rect 10075 6160 10095 6180
rect 10075 6110 10095 6130
rect 10075 6065 10095 6085
rect 10075 6020 10095 6040
rect 10175 6250 10195 6270
rect 10175 6205 10195 6225
rect 10175 6160 10195 6180
rect 10175 6110 10195 6130
rect 10175 6065 10195 6085
rect 10175 6020 10195 6040
rect 10275 6250 10295 6270
rect 10275 6205 10295 6225
rect 10275 6160 10295 6180
rect 10275 6110 10295 6130
rect 10275 6065 10295 6085
rect 10275 6020 10295 6040
rect 10375 6250 10395 6270
rect 10375 6205 10395 6225
rect 10375 6160 10395 6180
rect 10375 6110 10395 6130
rect 10375 6065 10395 6085
rect 10375 6020 10395 6040
rect 10475 6250 10495 6270
rect 10475 6205 10495 6225
rect 10475 6160 10495 6180
rect 10475 6110 10495 6130
rect 10475 6065 10495 6085
rect 10475 6020 10495 6040
rect 10575 6250 10595 6270
rect 10575 6205 10595 6225
rect 10575 6160 10595 6180
rect 10575 6110 10595 6130
rect 10575 6065 10595 6085
rect 10575 6020 10595 6040
rect 10675 6250 10695 6270
rect 10675 6205 10695 6225
rect 10675 6160 10695 6180
rect 10675 6110 10695 6130
rect 10675 6065 10695 6085
rect 10675 6020 10695 6040
rect 10775 6250 10795 6270
rect 10775 6205 10795 6225
rect 10775 6160 10795 6180
rect 10775 6110 10795 6130
rect 10775 6065 10795 6085
rect 10775 6020 10795 6040
rect 10875 6250 10895 6270
rect 10875 6205 10895 6225
rect 12905 6250 12925 6270
rect 12905 6205 12925 6225
rect 10875 6160 10895 6180
rect 10875 6110 10895 6130
rect 10875 6065 10895 6085
rect 10875 6020 10895 6040
rect 11215 6150 11235 6170
rect 11215 6100 11235 6120
rect 11215 6050 11235 6070
rect 11215 6000 11235 6020
rect 11215 5950 11235 5970
rect 11270 6150 11290 6170
rect 11270 6100 11290 6120
rect 11270 6050 11290 6070
rect 11270 6000 11290 6020
rect 11270 5950 11290 5970
rect 11325 6150 11345 6170
rect 11325 6100 11345 6120
rect 11325 6050 11345 6070
rect 11325 6000 11345 6020
rect 11325 5950 11345 5970
rect 11380 6150 11400 6170
rect 11380 6100 11400 6120
rect 11380 6050 11400 6070
rect 11380 6000 11400 6020
rect 11380 5950 11400 5970
rect 11435 6150 11455 6170
rect 11435 6100 11455 6120
rect 11435 6050 11455 6070
rect 11435 6000 11455 6020
rect 11435 5950 11455 5970
rect 11490 6150 11510 6170
rect 11490 6100 11510 6120
rect 11490 6050 11510 6070
rect 11490 6000 11510 6020
rect 11490 5950 11510 5970
rect 11545 6150 11565 6170
rect 11545 6100 11565 6120
rect 11545 6050 11565 6070
rect 11545 6000 11565 6020
rect 11545 5950 11565 5970
rect 11600 6150 11620 6170
rect 11600 6100 11620 6120
rect 11600 6050 11620 6070
rect 11600 6000 11620 6020
rect 11600 5950 11620 5970
rect 11655 6150 11675 6170
rect 11655 6100 11675 6120
rect 11655 6050 11675 6070
rect 11655 6000 11675 6020
rect 11655 5950 11675 5970
rect 11710 6150 11730 6170
rect 11710 6100 11730 6120
rect 11710 6050 11730 6070
rect 11710 6000 11730 6020
rect 11710 5950 11730 5970
rect 11765 6150 11785 6170
rect 11765 6100 11785 6120
rect 11765 6050 11785 6070
rect 11765 6000 11785 6020
rect 11765 5950 11785 5970
rect 11820 6150 11840 6170
rect 11820 6100 11840 6120
rect 11820 6050 11840 6070
rect 11820 6000 11840 6020
rect 11820 5950 11840 5970
rect 11875 6150 11895 6170
rect 11875 6100 11895 6120
rect 11875 6050 11895 6070
rect 11875 6000 11895 6020
rect 11875 5950 11895 5970
rect 11930 6150 11950 6170
rect 11930 6100 11950 6120
rect 11930 6050 11950 6070
rect 11930 6000 11950 6020
rect 11930 5950 11950 5970
rect 11985 6150 12005 6170
rect 11985 6100 12005 6120
rect 11985 6050 12005 6070
rect 11985 6000 12005 6020
rect 11985 5950 12005 5970
rect 12040 6150 12060 6170
rect 12040 6100 12060 6120
rect 12040 6050 12060 6070
rect 12040 6000 12060 6020
rect 12040 5950 12060 5970
rect 12095 6150 12115 6170
rect 12095 6100 12115 6120
rect 12095 6050 12115 6070
rect 12095 6000 12115 6020
rect 12095 5950 12115 5970
rect 12150 6150 12170 6170
rect 12150 6100 12170 6120
rect 12150 6050 12170 6070
rect 12150 6000 12170 6020
rect 12150 5950 12170 5970
rect 12205 6150 12225 6170
rect 12205 6100 12225 6120
rect 12205 6050 12225 6070
rect 12205 6000 12225 6020
rect 12205 5950 12225 5970
rect 12260 6150 12280 6170
rect 12260 6100 12280 6120
rect 12260 6050 12280 6070
rect 12260 6000 12280 6020
rect 12260 5950 12280 5970
rect 12315 6150 12335 6170
rect 12315 6100 12335 6120
rect 12315 6050 12335 6070
rect 12315 6000 12335 6020
rect 12315 5950 12335 5970
rect 12370 6150 12390 6170
rect 12370 6100 12390 6120
rect 12370 6050 12390 6070
rect 12370 6000 12390 6020
rect 12370 5950 12390 5970
rect 12425 6150 12445 6170
rect 12425 6100 12445 6120
rect 12425 6050 12445 6070
rect 12425 6000 12445 6020
rect 12425 5950 12445 5970
rect 12480 6150 12500 6170
rect 12480 6100 12500 6120
rect 12480 6050 12500 6070
rect 12480 6000 12500 6020
rect 12480 5950 12500 5970
rect 12535 6150 12555 6170
rect 12535 6100 12555 6120
rect 12535 6050 12555 6070
rect 12535 6000 12555 6020
rect 12535 5950 12555 5970
rect 12590 6150 12610 6170
rect 12590 6100 12610 6120
rect 12590 6050 12610 6070
rect 12590 6000 12610 6020
rect 12905 6160 12925 6180
rect 12905 6110 12925 6130
rect 12905 6065 12925 6085
rect 12905 6020 12925 6040
rect 13005 6250 13025 6270
rect 13005 6205 13025 6225
rect 13005 6160 13025 6180
rect 13005 6110 13025 6130
rect 13005 6065 13025 6085
rect 13005 6020 13025 6040
rect 13105 6250 13125 6270
rect 13105 6205 13125 6225
rect 13105 6160 13125 6180
rect 13105 6110 13125 6130
rect 13105 6065 13125 6085
rect 13105 6020 13125 6040
rect 13205 6250 13225 6270
rect 13205 6205 13225 6225
rect 13205 6160 13225 6180
rect 13205 6110 13225 6130
rect 13205 6065 13225 6085
rect 13205 6020 13225 6040
rect 13305 6250 13325 6270
rect 13305 6205 13325 6225
rect 13305 6160 13325 6180
rect 13305 6110 13325 6130
rect 13305 6065 13325 6085
rect 13305 6020 13325 6040
rect 13405 6250 13425 6270
rect 13405 6205 13425 6225
rect 13405 6160 13425 6180
rect 13405 6110 13425 6130
rect 13405 6065 13425 6085
rect 13405 6020 13425 6040
rect 13505 6250 13525 6270
rect 13505 6205 13525 6225
rect 13505 6160 13525 6180
rect 13505 6110 13525 6130
rect 13505 6065 13525 6085
rect 13505 6020 13525 6040
rect 13605 6250 13625 6270
rect 13605 6205 13625 6225
rect 13605 6160 13625 6180
rect 13605 6110 13625 6130
rect 13605 6065 13625 6085
rect 13605 6020 13625 6040
rect 13705 6250 13725 6270
rect 13705 6205 13725 6225
rect 13705 6160 13725 6180
rect 13705 6110 13725 6130
rect 13705 6065 13725 6085
rect 13705 6020 13725 6040
rect 13805 6250 13825 6270
rect 13805 6205 13825 6225
rect 13805 6160 13825 6180
rect 13805 6110 13825 6130
rect 13805 6065 13825 6085
rect 13805 6020 13825 6040
rect 13905 6250 13925 6270
rect 13905 6205 13925 6225
rect 13905 6160 13925 6180
rect 13905 6110 13925 6130
rect 13905 6065 13925 6085
rect 13905 6020 13925 6040
rect 14005 6250 14025 6270
rect 14005 6205 14025 6225
rect 14005 6160 14025 6180
rect 14005 6110 14025 6130
rect 14005 6065 14025 6085
rect 14005 6020 14025 6040
rect 14105 6250 14125 6270
rect 14105 6205 14125 6225
rect 14105 6160 14125 6180
rect 14105 6110 14125 6130
rect 14105 6065 14125 6085
rect 14105 6020 14125 6040
rect 18715 6190 18735 6210
rect 18715 6140 18735 6160
rect 18715 6090 18735 6110
rect 18715 6040 18735 6060
rect 12590 5950 12610 5970
rect 18715 5990 18735 6010
rect 18770 6190 18790 6210
rect 18770 6140 18790 6160
rect 18770 6090 18790 6110
rect 18770 6040 18790 6060
rect 18770 5990 18790 6010
rect 18825 6190 18845 6210
rect 18825 6140 18845 6160
rect 18825 6090 18845 6110
rect 18825 6040 18845 6060
rect 18825 5990 18845 6010
rect 18880 6190 18900 6210
rect 18880 6140 18900 6160
rect 18880 6090 18900 6110
rect 18880 6040 18900 6060
rect 18880 5990 18900 6010
rect 18935 6190 18955 6210
rect 18935 6140 18955 6160
rect 18935 6090 18955 6110
rect 18935 6040 18955 6060
rect 18935 5990 18955 6010
rect 18990 6190 19010 6210
rect 18990 6140 19010 6160
rect 18990 6090 19010 6110
rect 18990 6040 19010 6060
rect 18990 5990 19010 6010
rect 19045 6190 19065 6210
rect 19045 6140 19065 6160
rect 19045 6090 19065 6110
rect 19045 6040 19065 6060
rect 19045 5990 19065 6010
rect 19100 6190 19120 6210
rect 19100 6140 19120 6160
rect 19100 6090 19120 6110
rect 19100 6040 19120 6060
rect 19100 5990 19120 6010
rect 19155 6190 19175 6210
rect 19155 6140 19175 6160
rect 19155 6090 19175 6110
rect 19155 6040 19175 6060
rect 19155 5990 19175 6010
rect 19210 6190 19230 6210
rect 19210 6140 19230 6160
rect 19210 6090 19230 6110
rect 19210 6040 19230 6060
rect 19210 5990 19230 6010
rect 19265 6190 19285 6210
rect 19265 6140 19285 6160
rect 19265 6090 19285 6110
rect 19265 6040 19285 6060
rect 19265 5990 19285 6010
rect 19320 6190 19340 6210
rect 19320 6140 19340 6160
rect 19320 6090 19340 6110
rect 19320 6040 19340 6060
rect 19320 5990 19340 6010
rect 19375 6190 19395 6210
rect 19375 6140 19395 6160
rect 19375 6090 19395 6110
rect 19375 6040 19395 6060
rect 19375 5990 19395 6010
rect 19430 6190 19450 6210
rect 19430 6140 19450 6160
rect 19430 6090 19450 6110
rect 19430 6040 19450 6060
rect 19430 5990 19450 6010
rect 19485 6190 19505 6210
rect 19485 6140 19505 6160
rect 19485 6090 19505 6110
rect 19485 6040 19505 6060
rect 19485 5990 19505 6010
rect 19540 6190 19560 6210
rect 19540 6140 19560 6160
rect 19540 6090 19560 6110
rect 19540 6040 19560 6060
rect 19540 5990 19560 6010
rect 19595 6190 19615 6210
rect 19595 6140 19615 6160
rect 19595 6090 19615 6110
rect 19595 6040 19615 6060
rect 19595 5990 19615 6010
rect 19650 6190 19670 6210
rect 19650 6140 19670 6160
rect 19650 6090 19670 6110
rect 19650 6040 19670 6060
rect 19650 5990 19670 6010
rect 19705 6190 19725 6210
rect 19705 6140 19725 6160
rect 19705 6090 19725 6110
rect 19705 6040 19725 6060
rect 19705 5990 19725 6010
rect 19760 6190 19780 6210
rect 19760 6140 19780 6160
rect 19760 6090 19780 6110
rect 19760 6040 19780 6060
rect 19760 5990 19780 6010
rect 19815 6190 19835 6210
rect 19815 6140 19835 6160
rect 19815 6090 19835 6110
rect 19815 6040 19835 6060
rect 19815 5990 19835 6010
rect 19870 6190 19890 6210
rect 19870 6140 19890 6160
rect 19870 6090 19890 6110
rect 19870 6040 19890 6060
rect 19870 5990 19890 6010
rect 19925 6190 19945 6210
rect 19925 6140 19945 6160
rect 19925 6090 19945 6110
rect 19925 6040 19945 6060
rect 19925 5990 19945 6010
rect 19980 6190 20000 6210
rect 19980 6140 20000 6160
rect 19980 6090 20000 6110
rect 19980 6040 20000 6060
rect 19980 5990 20000 6010
rect 20035 6190 20055 6210
rect 20035 6140 20055 6160
rect 20035 6090 20055 6110
rect 20035 6040 20055 6060
rect 20035 5990 20055 6010
rect 20090 6190 20110 6210
rect 20090 6140 20110 6160
rect 20090 6090 20110 6110
rect 20090 6040 20110 6060
rect 20555 6145 20575 6165
rect 20555 6095 20575 6115
rect 20555 6045 20575 6065
rect 20610 6145 20630 6165
rect 20610 6095 20630 6115
rect 20610 6045 20630 6065
rect 20665 6145 20685 6165
rect 20665 6095 20685 6115
rect 20665 6045 20685 6065
rect 20720 6145 20740 6165
rect 20720 6095 20740 6115
rect 20720 6045 20740 6065
rect 20775 6145 20795 6165
rect 20775 6095 20795 6115
rect 20775 6045 20795 6065
rect 20090 5990 20110 6010
rect 11250 4355 11270 4375
rect 11310 4360 11330 4380
rect 11370 4360 11390 4380
rect 11430 4355 11450 4375
rect 11580 4370 11600 4390
rect 11640 4370 11660 4390
rect 11700 4370 11720 4390
rect 11760 4370 11780 4390
rect 11820 4370 11840 4390
rect 11880 4370 11900 4390
rect 11940 4370 11960 4390
rect 12090 4355 12110 4375
rect 12150 4355 12170 4375
rect 12210 4355 12230 4375
rect 12270 4355 12290 4375
rect 12330 4355 12350 4375
rect 12390 4355 12410 4375
rect 12450 4355 12470 4375
rect 12510 4355 12530 4375
rect 12570 4355 12590 4375
rect 11260 4120 11280 4140
rect 11315 4120 11335 4140
rect 11370 4120 11390 4140
rect 11425 4120 11445 4140
rect 11480 4120 11500 4140
rect 11535 4120 11555 4140
rect 11590 4120 11610 4140
rect 11645 4120 11665 4140
rect 11700 4120 11720 4140
rect 11755 4120 11775 4140
rect 11810 4120 11830 4140
rect 11865 4120 11885 4140
rect 11920 4120 11940 4140
rect 11975 4120 11995 4140
rect 12030 4120 12050 4140
rect 12085 4120 12105 4140
rect 12140 4120 12160 4140
rect 12195 4120 12215 4140
rect 12250 4120 12270 4140
rect 12305 4120 12325 4140
rect 12360 4120 12380 4140
rect 12415 4120 12435 4140
rect 12470 4120 12490 4140
rect 11205 3815 11225 3835
rect 11260 3815 11280 3835
rect 11315 3815 11335 3835
rect 11370 3815 11390 3835
rect 11425 3815 11445 3835
rect 11480 3815 11500 3835
rect 11535 3815 11555 3835
rect 11590 3815 11610 3835
rect 11645 3815 11665 3835
rect 11700 3815 11720 3835
rect 11755 3815 11775 3835
rect 11810 3815 11830 3835
rect 11865 3815 11885 3835
rect 11945 3815 11965 3835
rect 12000 3815 12020 3835
rect 12055 3815 12075 3835
rect 12110 3815 12130 3835
rect 12165 3815 12185 3835
rect 12220 3815 12240 3835
rect 12275 3815 12295 3835
rect 12330 3815 12350 3835
rect 12385 3815 12405 3835
rect 12440 3815 12460 3835
rect 12495 3815 12515 3835
rect 12550 3815 12570 3835
rect 12605 3815 12625 3835
rect 10165 3550 10185 3570
rect 10165 3500 10185 3520
rect 10165 3450 10185 3470
rect 10165 3400 10185 3420
rect 10165 3350 10185 3370
rect 10165 3300 10185 3320
rect 10165 3250 10185 3270
rect 10165 3200 10185 3220
rect 10165 3150 10185 3170
rect 10165 3100 10185 3120
rect 10165 3050 10185 3070
rect 10165 3000 10185 3020
rect 10220 3550 10240 3570
rect 10220 3500 10240 3520
rect 10220 3450 10240 3470
rect 10220 3400 10240 3420
rect 10220 3350 10240 3370
rect 10220 3300 10240 3320
rect 10220 3250 10240 3270
rect 10220 3200 10240 3220
rect 10220 3150 10240 3170
rect 10220 3100 10240 3120
rect 10220 3050 10240 3070
rect 10220 3000 10240 3020
rect 10275 3550 10295 3570
rect 10275 3500 10295 3520
rect 10275 3450 10295 3470
rect 10275 3400 10295 3420
rect 10275 3350 10295 3370
rect 10275 3300 10295 3320
rect 10275 3250 10295 3270
rect 10275 3200 10295 3220
rect 10275 3150 10295 3170
rect 10275 3100 10295 3120
rect 10275 3050 10295 3070
rect 10275 3000 10295 3020
rect 10330 3550 10350 3570
rect 10330 3500 10350 3520
rect 10330 3450 10350 3470
rect 10330 3400 10350 3420
rect 10330 3350 10350 3370
rect 10330 3300 10350 3320
rect 10330 3250 10350 3270
rect 10330 3200 10350 3220
rect 10330 3150 10350 3170
rect 10330 3100 10350 3120
rect 10330 3050 10350 3070
rect 10330 3000 10350 3020
rect 10385 3550 10405 3570
rect 10385 3500 10405 3520
rect 10385 3450 10405 3470
rect 10385 3400 10405 3420
rect 10385 3350 10405 3370
rect 10385 3300 10405 3320
rect 10385 3250 10405 3270
rect 10385 3200 10405 3220
rect 10385 3150 10405 3170
rect 10385 3100 10405 3120
rect 10385 3050 10405 3070
rect 10385 3000 10405 3020
rect 10440 3550 10460 3570
rect 10440 3500 10460 3520
rect 10440 3450 10460 3470
rect 10440 3400 10460 3420
rect 10440 3350 10460 3370
rect 10440 3300 10460 3320
rect 10440 3250 10460 3270
rect 10440 3200 10460 3220
rect 10440 3150 10460 3170
rect 10440 3100 10460 3120
rect 10440 3050 10460 3070
rect 10440 3000 10460 3020
rect 10495 3550 10515 3570
rect 10495 3500 10515 3520
rect 10495 3450 10515 3470
rect 10495 3400 10515 3420
rect 10495 3350 10515 3370
rect 10495 3300 10515 3320
rect 10495 3250 10515 3270
rect 10495 3200 10515 3220
rect 10495 3150 10515 3170
rect 10495 3100 10515 3120
rect 10495 3050 10515 3070
rect 10495 3000 10515 3020
rect 10550 3550 10570 3570
rect 10550 3500 10570 3520
rect 10550 3450 10570 3470
rect 10550 3400 10570 3420
rect 10550 3350 10570 3370
rect 10550 3300 10570 3320
rect 10550 3250 10570 3270
rect 10550 3200 10570 3220
rect 10550 3150 10570 3170
rect 10550 3100 10570 3120
rect 10550 3050 10570 3070
rect 10550 3000 10570 3020
rect 10605 3550 10625 3570
rect 10605 3500 10625 3520
rect 10605 3450 10625 3470
rect 10605 3400 10625 3420
rect 10605 3350 10625 3370
rect 10605 3300 10625 3320
rect 10605 3250 10625 3270
rect 10605 3200 10625 3220
rect 10605 3150 10625 3170
rect 10605 3100 10625 3120
rect 10605 3050 10625 3070
rect 10605 3000 10625 3020
rect 10660 3550 10680 3570
rect 10660 3500 10680 3520
rect 10660 3450 10680 3470
rect 10660 3400 10680 3420
rect 10660 3350 10680 3370
rect 10660 3300 10680 3320
rect 10660 3250 10680 3270
rect 10660 3200 10680 3220
rect 10660 3150 10680 3170
rect 10660 3100 10680 3120
rect 10660 3050 10680 3070
rect 10660 3000 10680 3020
rect 10715 3550 10735 3570
rect 10715 3500 10735 3520
rect 10715 3450 10735 3470
rect 10715 3400 10735 3420
rect 10715 3350 10735 3370
rect 10715 3300 10735 3320
rect 10715 3250 10735 3270
rect 10715 3200 10735 3220
rect 10715 3150 10735 3170
rect 10715 3100 10735 3120
rect 10715 3050 10735 3070
rect 10715 3000 10735 3020
rect 10770 3550 10790 3570
rect 10770 3500 10790 3520
rect 10770 3450 10790 3470
rect 10770 3400 10790 3420
rect 10770 3350 10790 3370
rect 10770 3300 10790 3320
rect 10770 3250 10790 3270
rect 10770 3200 10790 3220
rect 10770 3150 10790 3170
rect 10770 3100 10790 3120
rect 10770 3050 10790 3070
rect 10770 3000 10790 3020
rect 10825 3550 10845 3570
rect 10825 3500 10845 3520
rect 10825 3450 10845 3470
rect 10825 3400 10845 3420
rect 10825 3350 10845 3370
rect 10825 3300 10845 3320
rect 10825 3250 10845 3270
rect 10825 3200 10845 3220
rect 11230 3540 11250 3560
rect 11230 3490 11250 3510
rect 11230 3440 11250 3460
rect 11230 3390 11250 3410
rect 11230 3340 11250 3360
rect 11230 3290 11250 3310
rect 11230 3240 11250 3260
rect 11230 3190 11250 3210
rect 11290 3540 11310 3560
rect 11290 3490 11310 3510
rect 11290 3440 11310 3460
rect 11290 3390 11310 3410
rect 11290 3340 11310 3360
rect 11290 3290 11310 3310
rect 11290 3240 11310 3260
rect 11290 3190 11310 3210
rect 11350 3540 11370 3560
rect 11350 3490 11370 3510
rect 11350 3440 11370 3460
rect 11350 3390 11370 3410
rect 11350 3340 11370 3360
rect 11350 3290 11370 3310
rect 11350 3240 11370 3260
rect 11350 3190 11370 3210
rect 11410 3540 11430 3560
rect 11410 3490 11430 3510
rect 11410 3440 11430 3460
rect 11410 3390 11430 3410
rect 11410 3340 11430 3360
rect 11410 3290 11430 3310
rect 11410 3240 11430 3260
rect 11410 3190 11430 3210
rect 11470 3540 11490 3560
rect 11470 3490 11490 3510
rect 11470 3440 11490 3460
rect 11470 3390 11490 3410
rect 11470 3340 11490 3360
rect 11470 3290 11490 3310
rect 11470 3240 11490 3260
rect 11470 3190 11490 3210
rect 11530 3540 11550 3560
rect 11530 3490 11550 3510
rect 11530 3440 11550 3460
rect 11530 3390 11550 3410
rect 11530 3340 11550 3360
rect 11530 3290 11550 3310
rect 11530 3240 11550 3260
rect 11530 3190 11550 3210
rect 11590 3540 11610 3560
rect 11590 3490 11610 3510
rect 11590 3440 11610 3460
rect 11590 3390 11610 3410
rect 11590 3340 11610 3360
rect 11590 3290 11610 3310
rect 11590 3240 11610 3260
rect 11590 3190 11610 3210
rect 11650 3540 11670 3560
rect 11650 3490 11670 3510
rect 11650 3440 11670 3460
rect 11650 3390 11670 3410
rect 11650 3340 11670 3360
rect 11650 3290 11670 3310
rect 11650 3240 11670 3260
rect 11650 3190 11670 3210
rect 11710 3540 11730 3560
rect 11710 3490 11730 3510
rect 11710 3440 11730 3460
rect 11710 3390 11730 3410
rect 11710 3340 11730 3360
rect 11710 3290 11730 3310
rect 11710 3240 11730 3260
rect 11710 3190 11730 3210
rect 11770 3540 11790 3560
rect 11770 3490 11790 3510
rect 11770 3440 11790 3460
rect 11770 3390 11790 3410
rect 11770 3340 11790 3360
rect 11770 3290 11790 3310
rect 11770 3240 11790 3260
rect 11770 3190 11790 3210
rect 11830 3540 11850 3560
rect 11830 3490 11850 3510
rect 11830 3440 11850 3460
rect 11830 3390 11850 3410
rect 11830 3340 11850 3360
rect 11830 3290 11850 3310
rect 11830 3240 11850 3260
rect 11830 3190 11850 3210
rect 11890 3540 11910 3560
rect 11890 3490 11910 3510
rect 11890 3440 11910 3460
rect 11890 3390 11910 3410
rect 11890 3340 11910 3360
rect 11890 3290 11910 3310
rect 11890 3240 11910 3260
rect 11890 3190 11910 3210
rect 11950 3540 11970 3560
rect 11950 3490 11970 3510
rect 11950 3440 11970 3460
rect 11950 3390 11970 3410
rect 11950 3340 11970 3360
rect 11950 3290 11970 3310
rect 11950 3240 11970 3260
rect 11950 3190 11970 3210
rect 12010 3540 12030 3560
rect 12010 3490 12030 3510
rect 12010 3440 12030 3460
rect 12010 3390 12030 3410
rect 12010 3340 12030 3360
rect 12010 3290 12030 3310
rect 12010 3240 12030 3260
rect 12010 3190 12030 3210
rect 12070 3540 12090 3560
rect 12070 3490 12090 3510
rect 12070 3440 12090 3460
rect 12070 3390 12090 3410
rect 12070 3340 12090 3360
rect 12070 3290 12090 3310
rect 12070 3240 12090 3260
rect 12070 3190 12090 3210
rect 12130 3540 12150 3560
rect 12130 3490 12150 3510
rect 12130 3440 12150 3460
rect 12130 3390 12150 3410
rect 12130 3340 12150 3360
rect 12130 3290 12150 3310
rect 12130 3240 12150 3260
rect 12130 3190 12150 3210
rect 12190 3540 12210 3560
rect 12190 3490 12210 3510
rect 12190 3440 12210 3460
rect 12190 3390 12210 3410
rect 12190 3340 12210 3360
rect 12190 3290 12210 3310
rect 12190 3240 12210 3260
rect 12190 3190 12210 3210
rect 12250 3540 12270 3560
rect 12250 3490 12270 3510
rect 12250 3440 12270 3460
rect 12250 3390 12270 3410
rect 12250 3340 12270 3360
rect 12250 3290 12270 3310
rect 12250 3240 12270 3260
rect 12250 3190 12270 3210
rect 12310 3540 12330 3560
rect 12310 3490 12330 3510
rect 12310 3440 12330 3460
rect 12310 3390 12330 3410
rect 12310 3340 12330 3360
rect 12310 3290 12330 3310
rect 12310 3240 12330 3260
rect 12310 3190 12330 3210
rect 12370 3540 12390 3560
rect 12370 3490 12390 3510
rect 12370 3440 12390 3460
rect 12370 3390 12390 3410
rect 12370 3340 12390 3360
rect 12370 3290 12390 3310
rect 12370 3240 12390 3260
rect 12370 3190 12390 3210
rect 12430 3540 12450 3560
rect 12430 3490 12450 3510
rect 12430 3440 12450 3460
rect 12430 3390 12450 3410
rect 12430 3340 12450 3360
rect 12430 3290 12450 3310
rect 12430 3240 12450 3260
rect 12430 3190 12450 3210
rect 12490 3540 12510 3560
rect 12490 3490 12510 3510
rect 12490 3440 12510 3460
rect 12490 3390 12510 3410
rect 12490 3340 12510 3360
rect 12490 3290 12510 3310
rect 12490 3240 12510 3260
rect 12490 3190 12510 3210
rect 12550 3540 12570 3560
rect 12550 3490 12570 3510
rect 12550 3440 12570 3460
rect 12550 3390 12570 3410
rect 12550 3340 12570 3360
rect 12550 3290 12570 3310
rect 12550 3240 12570 3260
rect 12550 3190 12570 3210
rect 12955 3550 12975 3570
rect 12955 3500 12975 3520
rect 12955 3450 12975 3470
rect 12955 3400 12975 3420
rect 12955 3350 12975 3370
rect 12955 3300 12975 3320
rect 12955 3250 12975 3270
rect 12955 3200 12975 3220
rect 10825 3150 10845 3170
rect 12955 3150 12975 3170
rect 10825 3100 10845 3120
rect 10825 3050 10845 3070
rect 10825 3000 10845 3020
rect 12955 3100 12975 3120
rect 12955 3050 12975 3070
rect 12955 3000 12975 3020
rect 13010 3550 13030 3570
rect 13010 3500 13030 3520
rect 13010 3450 13030 3470
rect 13010 3400 13030 3420
rect 13010 3350 13030 3370
rect 13010 3300 13030 3320
rect 13010 3250 13030 3270
rect 13010 3200 13030 3220
rect 13010 3150 13030 3170
rect 13010 3100 13030 3120
rect 13010 3050 13030 3070
rect 13010 3000 13030 3020
rect 13065 3550 13085 3570
rect 13065 3500 13085 3520
rect 13065 3450 13085 3470
rect 13065 3400 13085 3420
rect 13065 3350 13085 3370
rect 13065 3300 13085 3320
rect 13065 3250 13085 3270
rect 13065 3200 13085 3220
rect 13065 3150 13085 3170
rect 13065 3100 13085 3120
rect 13065 3050 13085 3070
rect 13065 3000 13085 3020
rect 13120 3550 13140 3570
rect 13120 3500 13140 3520
rect 13120 3450 13140 3470
rect 13120 3400 13140 3420
rect 13120 3350 13140 3370
rect 13120 3300 13140 3320
rect 13120 3250 13140 3270
rect 13120 3200 13140 3220
rect 13120 3150 13140 3170
rect 13120 3100 13140 3120
rect 13120 3050 13140 3070
rect 13120 3000 13140 3020
rect 13175 3550 13195 3570
rect 13175 3500 13195 3520
rect 13175 3450 13195 3470
rect 13175 3400 13195 3420
rect 13175 3350 13195 3370
rect 13175 3300 13195 3320
rect 13175 3250 13195 3270
rect 13175 3200 13195 3220
rect 13175 3150 13195 3170
rect 13175 3100 13195 3120
rect 13175 3050 13195 3070
rect 13175 3000 13195 3020
rect 13230 3550 13250 3570
rect 13230 3500 13250 3520
rect 13230 3450 13250 3470
rect 13230 3400 13250 3420
rect 13230 3350 13250 3370
rect 13230 3300 13250 3320
rect 13230 3250 13250 3270
rect 13230 3200 13250 3220
rect 13230 3150 13250 3170
rect 13230 3100 13250 3120
rect 13230 3050 13250 3070
rect 13230 3000 13250 3020
rect 13285 3550 13305 3570
rect 13285 3500 13305 3520
rect 13285 3450 13305 3470
rect 13285 3400 13305 3420
rect 13285 3350 13305 3370
rect 13285 3300 13305 3320
rect 13285 3250 13305 3270
rect 13285 3200 13305 3220
rect 13285 3150 13305 3170
rect 13285 3100 13305 3120
rect 13285 3050 13305 3070
rect 13285 3000 13305 3020
rect 13340 3550 13360 3570
rect 13340 3500 13360 3520
rect 13340 3450 13360 3470
rect 13340 3400 13360 3420
rect 13340 3350 13360 3370
rect 13340 3300 13360 3320
rect 13340 3250 13360 3270
rect 13340 3200 13360 3220
rect 13340 3150 13360 3170
rect 13340 3100 13360 3120
rect 13340 3050 13360 3070
rect 13340 3000 13360 3020
rect 13395 3550 13415 3570
rect 13395 3500 13415 3520
rect 13395 3450 13415 3470
rect 13395 3400 13415 3420
rect 13395 3350 13415 3370
rect 13395 3300 13415 3320
rect 13395 3250 13415 3270
rect 13395 3200 13415 3220
rect 13395 3150 13415 3170
rect 13395 3100 13415 3120
rect 13395 3050 13415 3070
rect 13395 3000 13415 3020
rect 13450 3550 13470 3570
rect 13450 3500 13470 3520
rect 13450 3450 13470 3470
rect 13450 3400 13470 3420
rect 13450 3350 13470 3370
rect 13450 3300 13470 3320
rect 13450 3250 13470 3270
rect 13450 3200 13470 3220
rect 13450 3150 13470 3170
rect 13450 3100 13470 3120
rect 13450 3050 13470 3070
rect 13450 3000 13470 3020
rect 13505 3550 13525 3570
rect 13505 3500 13525 3520
rect 13505 3450 13525 3470
rect 13505 3400 13525 3420
rect 13505 3350 13525 3370
rect 13505 3300 13525 3320
rect 13505 3250 13525 3270
rect 13505 3200 13525 3220
rect 13505 3150 13525 3170
rect 13505 3100 13525 3120
rect 13505 3050 13525 3070
rect 13505 3000 13525 3020
rect 13560 3550 13580 3570
rect 13560 3500 13580 3520
rect 13560 3450 13580 3470
rect 13560 3400 13580 3420
rect 13560 3350 13580 3370
rect 13560 3300 13580 3320
rect 13560 3250 13580 3270
rect 13560 3200 13580 3220
rect 13560 3150 13580 3170
rect 13560 3100 13580 3120
rect 13560 3050 13580 3070
rect 13560 3000 13580 3020
rect 13615 3550 13635 3570
rect 13615 3500 13635 3520
rect 13615 3450 13635 3470
rect 13615 3400 13635 3420
rect 13615 3350 13635 3370
rect 13615 3300 13635 3320
rect 13615 3250 13635 3270
rect 13615 3200 13635 3220
rect 13615 3150 13635 3170
rect 13615 3100 13635 3120
rect 13615 3050 13635 3070
rect 13615 3000 13635 3020
rect 25830 3495 25850 3515
rect 25830 3445 25850 3465
rect 25830 3395 25850 3415
rect 25830 3345 25850 3365
rect 25830 3295 25850 3315
rect 25500 3245 25520 3265
rect 25560 3250 25580 3270
rect 25620 3250 25640 3270
rect 25680 3245 25700 3265
rect 25830 3245 25850 3265
rect 25890 3495 25910 3515
rect 25890 3445 25910 3465
rect 25890 3395 25910 3415
rect 25890 3345 25910 3365
rect 25890 3295 25910 3315
rect 25890 3245 25910 3265
rect 25950 3495 25970 3515
rect 25950 3445 25970 3465
rect 25950 3395 25970 3415
rect 25950 3345 25970 3365
rect 25950 3295 25970 3315
rect 25950 3245 25970 3265
rect 26010 3545 26030 3565
rect 26010 3495 26030 3515
rect 26010 3445 26030 3465
rect 26010 3395 26030 3415
rect 26010 3345 26030 3365
rect 26010 3295 26030 3315
rect 26010 3245 26030 3265
rect 26070 3545 26090 3565
rect 26070 3495 26090 3515
rect 26070 3445 26090 3465
rect 26070 3395 26090 3415
rect 26070 3345 26090 3365
rect 26070 3295 26090 3315
rect 26070 3245 26090 3265
rect 26230 3540 26250 3560
rect 26230 3490 26250 3510
rect 26230 3440 26250 3460
rect 26230 3390 26250 3410
rect 26230 3340 26250 3360
rect 26230 3290 26250 3310
rect 26230 3240 26250 3260
rect 26230 3190 26250 3210
rect 26290 3540 26310 3560
rect 26290 3490 26310 3510
rect 26290 3440 26310 3460
rect 26290 3390 26310 3410
rect 26290 3340 26310 3360
rect 26290 3290 26310 3310
rect 26290 3240 26310 3260
rect 26290 3190 26310 3210
rect 26350 3540 26370 3560
rect 26350 3490 26370 3510
rect 26350 3440 26370 3460
rect 26350 3390 26370 3410
rect 26350 3340 26370 3360
rect 26350 3290 26370 3310
rect 26350 3240 26370 3260
rect 26350 3190 26370 3210
rect 26410 3540 26430 3560
rect 26410 3490 26430 3510
rect 26410 3440 26430 3460
rect 26410 3390 26430 3410
rect 26410 3340 26430 3360
rect 26410 3290 26430 3310
rect 26410 3240 26430 3260
rect 26410 3190 26430 3210
rect 26470 3540 26490 3560
rect 26470 3490 26490 3510
rect 26470 3440 26490 3460
rect 26470 3390 26490 3410
rect 26470 3340 26490 3360
rect 26470 3290 26490 3310
rect 26470 3240 26490 3260
rect 26470 3190 26490 3210
rect 26530 3540 26550 3560
rect 26530 3490 26550 3510
rect 26530 3440 26550 3460
rect 26530 3390 26550 3410
rect 26530 3340 26550 3360
rect 26530 3290 26550 3310
rect 26530 3240 26550 3260
rect 26530 3190 26550 3210
rect 26590 3540 26610 3560
rect 26590 3490 26610 3510
rect 26590 3440 26610 3460
rect 26590 3390 26610 3410
rect 26590 3340 26610 3360
rect 26590 3290 26610 3310
rect 26590 3240 26610 3260
rect 26590 3190 26610 3210
rect 26650 3540 26670 3560
rect 26650 3490 26670 3510
rect 26650 3440 26670 3460
rect 26650 3390 26670 3410
rect 26650 3340 26670 3360
rect 26650 3290 26670 3310
rect 26650 3240 26670 3260
rect 26650 3190 26670 3210
rect 26710 3540 26730 3560
rect 26710 3490 26730 3510
rect 26710 3440 26730 3460
rect 26710 3390 26730 3410
rect 26710 3340 26730 3360
rect 26710 3290 26730 3310
rect 26710 3240 26730 3260
rect 26710 3190 26730 3210
rect 26770 3540 26790 3560
rect 26770 3490 26790 3510
rect 26770 3440 26790 3460
rect 26770 3390 26790 3410
rect 26770 3340 26790 3360
rect 26770 3290 26790 3310
rect 26770 3240 26790 3260
rect 26770 3190 26790 3210
rect 26830 3540 26850 3560
rect 26830 3490 26850 3510
rect 26830 3440 26850 3460
rect 26830 3390 26850 3410
rect 26830 3340 26850 3360
rect 26830 3290 26850 3310
rect 26830 3240 26850 3260
rect 26830 3190 26850 3210
rect 26890 3540 26910 3560
rect 26890 3490 26910 3510
rect 26890 3440 26910 3460
rect 26890 3390 26910 3410
rect 26890 3340 26910 3360
rect 26890 3290 26910 3310
rect 26890 3240 26910 3260
rect 26890 3190 26910 3210
rect 26950 3540 26970 3560
rect 26950 3490 26970 3510
rect 26950 3440 26970 3460
rect 26950 3390 26970 3410
rect 26950 3340 26970 3360
rect 26950 3290 26970 3310
rect 26950 3240 26970 3260
rect 26950 3190 26970 3210
rect 27010 3540 27030 3560
rect 27010 3490 27030 3510
rect 27010 3440 27030 3460
rect 27010 3390 27030 3410
rect 27010 3340 27030 3360
rect 27010 3290 27030 3310
rect 27010 3240 27030 3260
rect 27010 3190 27030 3210
rect 27070 3540 27090 3560
rect 27070 3490 27090 3510
rect 27070 3440 27090 3460
rect 27070 3390 27090 3410
rect 27070 3340 27090 3360
rect 27070 3290 27090 3310
rect 27070 3240 27090 3260
rect 27070 3190 27090 3210
rect 27130 3540 27150 3560
rect 27130 3490 27150 3510
rect 27130 3440 27150 3460
rect 27130 3390 27150 3410
rect 27130 3340 27150 3360
rect 27130 3290 27150 3310
rect 27130 3240 27150 3260
rect 27130 3190 27150 3210
rect 27190 3540 27210 3560
rect 27190 3490 27210 3510
rect 27190 3440 27210 3460
rect 27190 3390 27210 3410
rect 27190 3340 27210 3360
rect 27190 3290 27210 3310
rect 27190 3240 27210 3260
rect 27190 3190 27210 3210
rect 27250 3540 27270 3560
rect 27250 3490 27270 3510
rect 27250 3440 27270 3460
rect 27250 3390 27270 3410
rect 27250 3340 27270 3360
rect 27250 3290 27270 3310
rect 27250 3240 27270 3260
rect 27250 3190 27270 3210
rect 27310 3540 27330 3560
rect 27310 3490 27330 3510
rect 27310 3440 27330 3460
rect 27310 3390 27330 3410
rect 27310 3340 27330 3360
rect 27310 3290 27330 3310
rect 27310 3240 27330 3260
rect 27310 3190 27330 3210
rect 27370 3540 27390 3560
rect 27370 3490 27390 3510
rect 27370 3440 27390 3460
rect 27370 3390 27390 3410
rect 27370 3340 27390 3360
rect 27370 3290 27390 3310
rect 27370 3240 27390 3260
rect 27370 3190 27390 3210
rect 27430 3540 27450 3560
rect 27430 3490 27450 3510
rect 27430 3440 27450 3460
rect 27430 3390 27450 3410
rect 27430 3340 27450 3360
rect 27430 3290 27450 3310
rect 27430 3240 27450 3260
rect 27430 3190 27450 3210
rect 27490 3540 27510 3560
rect 27490 3490 27510 3510
rect 27490 3440 27510 3460
rect 27490 3390 27510 3410
rect 27490 3340 27510 3360
rect 27490 3290 27510 3310
rect 27490 3240 27510 3260
rect 27490 3190 27510 3210
rect 27550 3540 27570 3560
rect 27550 3490 27570 3510
rect 27550 3440 27570 3460
rect 27550 3390 27570 3410
rect 27550 3340 27570 3360
rect 27550 3290 27570 3310
rect 27550 3240 27570 3260
rect 27550 3190 27570 3210
rect 27900 3205 27920 3225
rect 27900 3155 27920 3175
rect 27900 3105 27920 3125
rect 27900 3055 27920 3075
rect 27900 3005 27920 3025
rect 27900 2955 27920 2975
rect 27955 3205 27975 3225
rect 27955 3155 27975 3175
rect 27955 3105 27975 3125
rect 27955 3055 27975 3075
rect 27955 3005 27975 3025
rect 27955 2955 27975 2975
rect 28010 3205 28030 3225
rect 28010 3155 28030 3175
rect 28010 3105 28030 3125
rect 28010 3055 28030 3075
rect 28010 3005 28030 3025
rect 28010 2955 28030 2975
rect 28065 3205 28085 3225
rect 28065 3155 28085 3175
rect 28065 3105 28085 3125
rect 28065 3055 28085 3075
rect 28065 3005 28085 3025
rect 28065 2955 28085 2975
rect 28120 3205 28140 3225
rect 28120 3155 28140 3175
rect 28120 3105 28140 3125
rect 28120 3055 28140 3075
rect 28120 3005 28140 3025
rect 28120 2955 28140 2975
rect 28175 3205 28195 3225
rect 28175 3155 28195 3175
rect 28175 3105 28195 3125
rect 28175 3055 28195 3075
rect 28175 3005 28195 3025
rect 28175 2955 28195 2975
rect 28230 3205 28250 3225
rect 28230 3155 28250 3175
rect 28230 3105 28250 3125
rect 28230 3055 28250 3075
rect 28230 3005 28250 3025
rect 28230 2955 28250 2975
rect 28285 3205 28305 3225
rect 28285 3155 28305 3175
rect 28285 3105 28305 3125
rect 28285 3055 28305 3075
rect 28285 3005 28305 3025
rect 28285 2955 28305 2975
rect 28340 3205 28360 3225
rect 28340 3155 28360 3175
rect 28340 3105 28360 3125
rect 28340 3055 28360 3075
rect 28340 3005 28360 3025
rect 28340 2955 28360 2975
rect 28395 3205 28415 3225
rect 28395 3155 28415 3175
rect 28395 3105 28415 3125
rect 28395 3055 28415 3075
rect 28395 3005 28415 3025
rect 28395 2955 28415 2975
rect 28450 3205 28470 3225
rect 28450 3155 28470 3175
rect 28450 3105 28470 3125
rect 28450 3055 28470 3075
rect 28450 3005 28470 3025
rect 28450 2955 28470 2975
rect 28505 3205 28525 3225
rect 28505 3155 28525 3175
rect 28505 3105 28525 3125
rect 28505 3055 28525 3075
rect 28505 3005 28525 3025
rect 28505 2955 28525 2975
rect 28560 3205 28580 3225
rect 28560 3155 28580 3175
rect 28560 3105 28580 3125
rect 28560 3055 28580 3075
rect 28560 3005 28580 3025
rect 28560 2955 28580 2975
rect 28615 3205 28635 3225
rect 28615 3155 28635 3175
rect 28615 3105 28635 3125
rect 28615 3055 28635 3075
rect 28615 3005 28635 3025
rect 28615 2955 28635 2975
rect 28670 3205 28690 3225
rect 28670 3155 28690 3175
rect 28670 3105 28690 3125
rect 28670 3055 28690 3075
rect 28670 3005 28690 3025
rect 28670 2955 28690 2975
rect 28725 3205 28745 3225
rect 28725 3155 28745 3175
rect 28725 3105 28745 3125
rect 28725 3055 28745 3075
rect 28725 3005 28745 3025
rect 28725 2955 28745 2975
rect 28780 3205 28800 3225
rect 28780 3155 28800 3175
rect 28780 3105 28800 3125
rect 28780 3055 28800 3075
rect 28780 3005 28800 3025
rect 28780 2955 28800 2975
rect 28835 3205 28855 3225
rect 28835 3155 28855 3175
rect 28835 3105 28855 3125
rect 28835 3055 28855 3075
rect 28835 3005 28855 3025
rect 28835 2955 28855 2975
rect 28890 3205 28910 3225
rect 28890 3155 28910 3175
rect 28890 3105 28910 3125
rect 28890 3055 28910 3075
rect 28890 3005 28910 3025
rect 28890 2955 28910 2975
rect 28945 3205 28965 3225
rect 28945 3155 28965 3175
rect 28945 3105 28965 3125
rect 28945 3055 28965 3075
rect 28945 3005 28965 3025
rect 28945 2955 28965 2975
rect 29000 3205 29020 3225
rect 29000 3155 29020 3175
rect 29000 3105 29020 3125
rect 29000 3055 29020 3075
rect 29000 3005 29020 3025
rect 29000 2955 29020 2975
rect 29055 3205 29075 3225
rect 29055 3155 29075 3175
rect 29055 3105 29075 3125
rect 29055 3055 29075 3075
rect 29055 3005 29075 3025
rect 29055 2955 29075 2975
rect 29110 3205 29130 3225
rect 29110 3155 29130 3175
rect 29110 3105 29130 3125
rect 29110 3055 29130 3075
rect 29110 3005 29130 3025
rect 29110 2955 29130 2975
rect 11230 2860 11250 2880
rect 11230 2810 11250 2830
rect 11230 2760 11250 2780
rect 11230 2710 11250 2730
rect 11230 2660 11250 2680
rect 10165 2620 10185 2640
rect 10165 2570 10185 2590
rect 10165 2520 10185 2540
rect 10165 2470 10185 2490
rect 10220 2620 10240 2640
rect 10220 2570 10240 2590
rect 10220 2520 10240 2540
rect 10220 2470 10240 2490
rect 10275 2620 10295 2640
rect 10275 2570 10295 2590
rect 10275 2520 10295 2540
rect 10275 2470 10295 2490
rect 10330 2620 10350 2640
rect 10330 2570 10350 2590
rect 10330 2520 10350 2540
rect 10330 2470 10350 2490
rect 10385 2620 10405 2640
rect 10385 2570 10405 2590
rect 10385 2520 10405 2540
rect 10385 2470 10405 2490
rect 10440 2620 10460 2640
rect 10440 2570 10460 2590
rect 10440 2520 10460 2540
rect 10440 2470 10460 2490
rect 10495 2620 10515 2640
rect 10495 2570 10515 2590
rect 10495 2520 10515 2540
rect 10495 2470 10515 2490
rect 10550 2620 10570 2640
rect 10550 2570 10570 2590
rect 10550 2520 10570 2540
rect 10550 2470 10570 2490
rect 10605 2620 10625 2640
rect 10605 2570 10625 2590
rect 10605 2520 10625 2540
rect 10605 2470 10625 2490
rect 10660 2620 10680 2640
rect 10660 2570 10680 2590
rect 10660 2520 10680 2540
rect 10660 2470 10680 2490
rect 10715 2620 10735 2640
rect 10715 2570 10735 2590
rect 10715 2520 10735 2540
rect 10715 2470 10735 2490
rect 10770 2620 10790 2640
rect 10770 2570 10790 2590
rect 10770 2520 10790 2540
rect 10770 2470 10790 2490
rect 10825 2620 10845 2640
rect 10825 2570 10845 2590
rect 10825 2520 10845 2540
rect 11230 2610 11250 2630
rect 11230 2560 11250 2580
rect 11230 2510 11250 2530
rect 11290 2860 11310 2880
rect 11290 2810 11310 2830
rect 11290 2760 11310 2780
rect 11290 2710 11310 2730
rect 11290 2660 11310 2680
rect 11290 2610 11310 2630
rect 11290 2560 11310 2580
rect 11290 2510 11310 2530
rect 11350 2860 11370 2880
rect 11350 2810 11370 2830
rect 11350 2760 11370 2780
rect 11350 2710 11370 2730
rect 11350 2660 11370 2680
rect 11350 2610 11370 2630
rect 11350 2560 11370 2580
rect 11350 2510 11370 2530
rect 11410 2860 11430 2880
rect 11410 2810 11430 2830
rect 11410 2760 11430 2780
rect 11410 2710 11430 2730
rect 11410 2660 11430 2680
rect 11410 2610 11430 2630
rect 11410 2560 11430 2580
rect 11410 2510 11430 2530
rect 11470 2860 11490 2880
rect 11470 2810 11490 2830
rect 11470 2760 11490 2780
rect 11470 2710 11490 2730
rect 11470 2660 11490 2680
rect 11470 2610 11490 2630
rect 11470 2560 11490 2580
rect 11470 2510 11490 2530
rect 11530 2860 11550 2880
rect 11530 2810 11550 2830
rect 11530 2760 11550 2780
rect 11530 2710 11550 2730
rect 11530 2660 11550 2680
rect 11530 2610 11550 2630
rect 11530 2560 11550 2580
rect 11530 2510 11550 2530
rect 11590 2860 11610 2880
rect 11590 2810 11610 2830
rect 11590 2760 11610 2780
rect 11590 2710 11610 2730
rect 11590 2660 11610 2680
rect 11590 2610 11610 2630
rect 11590 2560 11610 2580
rect 11590 2510 11610 2530
rect 11650 2860 11670 2880
rect 11650 2810 11670 2830
rect 11650 2760 11670 2780
rect 11650 2710 11670 2730
rect 11650 2660 11670 2680
rect 11650 2610 11670 2630
rect 11650 2560 11670 2580
rect 11650 2510 11670 2530
rect 11710 2860 11730 2880
rect 11710 2810 11730 2830
rect 11710 2760 11730 2780
rect 11710 2710 11730 2730
rect 11710 2660 11730 2680
rect 11710 2610 11730 2630
rect 11710 2560 11730 2580
rect 11710 2510 11730 2530
rect 11770 2860 11790 2880
rect 11770 2810 11790 2830
rect 11770 2760 11790 2780
rect 11770 2710 11790 2730
rect 11770 2660 11790 2680
rect 11770 2610 11790 2630
rect 11770 2560 11790 2580
rect 11770 2510 11790 2530
rect 11830 2860 11850 2880
rect 11830 2810 11850 2830
rect 11830 2760 11850 2780
rect 11830 2710 11850 2730
rect 11830 2660 11850 2680
rect 11830 2610 11850 2630
rect 11830 2560 11850 2580
rect 11830 2510 11850 2530
rect 11890 2860 11910 2880
rect 11890 2810 11910 2830
rect 11890 2760 11910 2780
rect 11890 2710 11910 2730
rect 11890 2660 11910 2680
rect 11890 2610 11910 2630
rect 11890 2560 11910 2580
rect 11890 2510 11910 2530
rect 11950 2860 11970 2880
rect 11950 2810 11970 2830
rect 11950 2760 11970 2780
rect 11950 2710 11970 2730
rect 11950 2660 11970 2680
rect 11950 2610 11970 2630
rect 11950 2560 11970 2580
rect 11950 2510 11970 2530
rect 12010 2860 12030 2880
rect 12010 2810 12030 2830
rect 12010 2760 12030 2780
rect 12010 2710 12030 2730
rect 12010 2660 12030 2680
rect 12010 2610 12030 2630
rect 12010 2560 12030 2580
rect 12010 2510 12030 2530
rect 12070 2860 12090 2880
rect 12070 2810 12090 2830
rect 12070 2760 12090 2780
rect 12070 2710 12090 2730
rect 12070 2660 12090 2680
rect 12070 2610 12090 2630
rect 12070 2560 12090 2580
rect 12070 2510 12090 2530
rect 12130 2860 12150 2880
rect 12130 2810 12150 2830
rect 12130 2760 12150 2780
rect 12130 2710 12150 2730
rect 12130 2660 12150 2680
rect 12130 2610 12150 2630
rect 12130 2560 12150 2580
rect 12130 2510 12150 2530
rect 12190 2860 12210 2880
rect 12190 2810 12210 2830
rect 12190 2760 12210 2780
rect 12190 2710 12210 2730
rect 12190 2660 12210 2680
rect 12190 2610 12210 2630
rect 12190 2560 12210 2580
rect 12190 2510 12210 2530
rect 12250 2860 12270 2880
rect 12250 2810 12270 2830
rect 12250 2760 12270 2780
rect 12250 2710 12270 2730
rect 12250 2660 12270 2680
rect 12250 2610 12270 2630
rect 12250 2560 12270 2580
rect 12250 2510 12270 2530
rect 12310 2860 12330 2880
rect 12310 2810 12330 2830
rect 12310 2760 12330 2780
rect 12310 2710 12330 2730
rect 12310 2660 12330 2680
rect 12310 2610 12330 2630
rect 12310 2560 12330 2580
rect 12310 2510 12330 2530
rect 12370 2860 12390 2880
rect 12370 2810 12390 2830
rect 12370 2760 12390 2780
rect 12370 2710 12390 2730
rect 12370 2660 12390 2680
rect 12370 2610 12390 2630
rect 12370 2560 12390 2580
rect 12370 2510 12390 2530
rect 12430 2860 12450 2880
rect 12430 2810 12450 2830
rect 12430 2760 12450 2780
rect 12430 2710 12450 2730
rect 12430 2660 12450 2680
rect 12430 2610 12450 2630
rect 12430 2560 12450 2580
rect 12430 2510 12450 2530
rect 12490 2860 12510 2880
rect 12490 2810 12510 2830
rect 12490 2760 12510 2780
rect 12490 2710 12510 2730
rect 12490 2660 12510 2680
rect 12490 2610 12510 2630
rect 12490 2560 12510 2580
rect 12490 2510 12510 2530
rect 12550 2860 12570 2880
rect 12550 2810 12570 2830
rect 12550 2760 12570 2780
rect 12550 2710 12570 2730
rect 12550 2660 12570 2680
rect 26230 2860 26250 2880
rect 26230 2810 26250 2830
rect 26230 2760 26250 2780
rect 26230 2710 26250 2730
rect 26230 2660 26250 2680
rect 12550 2610 12570 2630
rect 12550 2560 12570 2580
rect 12550 2510 12570 2530
rect 12955 2620 12975 2640
rect 12955 2570 12975 2590
rect 12955 2520 12975 2540
rect 10825 2470 10845 2490
rect 12955 2470 12975 2490
rect 13010 2620 13030 2640
rect 13010 2570 13030 2590
rect 13010 2520 13030 2540
rect 13010 2470 13030 2490
rect 13065 2620 13085 2640
rect 13065 2570 13085 2590
rect 13065 2520 13085 2540
rect 13065 2470 13085 2490
rect 13120 2620 13140 2640
rect 13120 2570 13140 2590
rect 13120 2520 13140 2540
rect 13120 2470 13140 2490
rect 13175 2620 13195 2640
rect 13175 2570 13195 2590
rect 13175 2520 13195 2540
rect 13175 2470 13195 2490
rect 13230 2620 13250 2640
rect 13230 2570 13250 2590
rect 13230 2520 13250 2540
rect 13230 2470 13250 2490
rect 13285 2620 13305 2640
rect 13285 2570 13305 2590
rect 13285 2520 13305 2540
rect 13285 2470 13305 2490
rect 13340 2620 13360 2640
rect 13340 2570 13360 2590
rect 13340 2520 13360 2540
rect 13340 2470 13360 2490
rect 13395 2620 13415 2640
rect 13395 2570 13415 2590
rect 13395 2520 13415 2540
rect 13395 2470 13415 2490
rect 13450 2620 13470 2640
rect 13450 2570 13470 2590
rect 13450 2520 13470 2540
rect 13450 2470 13470 2490
rect 13505 2620 13525 2640
rect 13505 2570 13525 2590
rect 13505 2520 13525 2540
rect 13505 2470 13525 2490
rect 13560 2620 13580 2640
rect 13560 2570 13580 2590
rect 13560 2520 13580 2540
rect 13560 2470 13580 2490
rect 13615 2620 13635 2640
rect 13615 2570 13635 2590
rect 13615 2520 13635 2540
rect 13615 2470 13635 2490
rect 10165 2230 10185 2250
rect 10165 2180 10185 2200
rect 10165 2130 10185 2150
rect 10165 2080 10185 2100
rect 10165 2030 10185 2050
rect 10165 1980 10185 2000
rect 10220 2230 10240 2250
rect 10220 2180 10240 2200
rect 10220 2130 10240 2150
rect 10220 2080 10240 2100
rect 10220 2030 10240 2050
rect 10220 1980 10240 2000
rect 10275 2230 10295 2250
rect 10275 2180 10295 2200
rect 10275 2130 10295 2150
rect 10275 2080 10295 2100
rect 10275 2030 10295 2050
rect 10275 1980 10295 2000
rect 10330 2230 10350 2250
rect 10330 2180 10350 2200
rect 10330 2130 10350 2150
rect 10330 2080 10350 2100
rect 10330 2030 10350 2050
rect 10330 1980 10350 2000
rect 10385 2230 10405 2250
rect 10385 2180 10405 2200
rect 10385 2130 10405 2150
rect 10385 2080 10405 2100
rect 10385 2030 10405 2050
rect 10385 1980 10405 2000
rect 10440 2230 10460 2250
rect 10440 2180 10460 2200
rect 10440 2130 10460 2150
rect 10440 2080 10460 2100
rect 10440 2030 10460 2050
rect 10440 1980 10460 2000
rect 10495 2230 10515 2250
rect 10495 2180 10515 2200
rect 10495 2130 10515 2150
rect 10495 2080 10515 2100
rect 10495 2030 10515 2050
rect 10495 1980 10515 2000
rect 10550 2230 10570 2250
rect 10550 2180 10570 2200
rect 10550 2130 10570 2150
rect 10550 2080 10570 2100
rect 10550 2030 10570 2050
rect 10550 1980 10570 2000
rect 10605 2230 10625 2250
rect 10605 2180 10625 2200
rect 10605 2130 10625 2150
rect 10605 2080 10625 2100
rect 10605 2030 10625 2050
rect 10605 1980 10625 2000
rect 10660 2230 10680 2250
rect 10660 2180 10680 2200
rect 10660 2130 10680 2150
rect 10660 2080 10680 2100
rect 10660 2030 10680 2050
rect 10660 1980 10680 2000
rect 10715 2230 10735 2250
rect 10715 2180 10735 2200
rect 10715 2130 10735 2150
rect 10715 2080 10735 2100
rect 10715 2030 10735 2050
rect 10715 1980 10735 2000
rect 10770 2230 10790 2250
rect 10770 2180 10790 2200
rect 10770 2130 10790 2150
rect 10770 2080 10790 2100
rect 10770 2030 10790 2050
rect 10770 1980 10790 2000
rect 10825 2230 10845 2250
rect 10825 2180 10845 2200
rect 12955 2230 12975 2250
rect 12955 2180 12975 2200
rect 10825 2130 10845 2150
rect 12955 2130 12975 2150
rect 10825 2080 10845 2100
rect 10825 2030 10845 2050
rect 10825 1980 10845 2000
rect 11285 2095 11305 2115
rect 11285 2045 11305 2065
rect 11285 1995 11305 2015
rect 11340 2095 11360 2115
rect 11340 2045 11360 2065
rect 11340 1995 11360 2015
rect 11395 2095 11415 2115
rect 11395 2045 11415 2065
rect 11395 1995 11415 2015
rect 11450 2095 11470 2115
rect 11450 2045 11470 2065
rect 11450 1995 11470 2015
rect 11505 2095 11525 2115
rect 11505 2045 11525 2065
rect 11505 1995 11525 2015
rect 11560 2095 11580 2115
rect 11560 2045 11580 2065
rect 11560 1995 11580 2015
rect 11615 2095 11635 2115
rect 11615 2045 11635 2065
rect 11615 1995 11635 2015
rect 11670 2095 11690 2115
rect 11670 2045 11690 2065
rect 11670 1995 11690 2015
rect 11725 2095 11745 2115
rect 11725 2045 11745 2065
rect 11725 1995 11745 2015
rect 11780 2095 11800 2115
rect 11780 2045 11800 2065
rect 11780 1995 11800 2015
rect 11835 2095 11855 2115
rect 11835 2045 11855 2065
rect 11835 1995 11855 2015
rect 11890 2095 11910 2115
rect 11890 2045 11910 2065
rect 11890 1995 11910 2015
rect 11945 2095 11965 2115
rect 11945 2045 11965 2065
rect 11945 1995 11965 2015
rect 12000 2095 12020 2115
rect 12000 2045 12020 2065
rect 12000 1995 12020 2015
rect 12055 2095 12075 2115
rect 12055 2045 12075 2065
rect 12055 1995 12075 2015
rect 12110 2095 12130 2115
rect 12110 2045 12130 2065
rect 12110 1995 12130 2015
rect 12165 2095 12185 2115
rect 12165 2045 12185 2065
rect 12165 1995 12185 2015
rect 12220 2095 12240 2115
rect 12220 2045 12240 2065
rect 12220 1995 12240 2015
rect 12275 2095 12295 2115
rect 12275 2045 12295 2065
rect 12275 1995 12295 2015
rect 12330 2095 12350 2115
rect 12330 2045 12350 2065
rect 12330 1995 12350 2015
rect 12385 2095 12405 2115
rect 12385 2045 12405 2065
rect 12385 1995 12405 2015
rect 12440 2095 12460 2115
rect 12440 2045 12460 2065
rect 12440 1995 12460 2015
rect 12495 2095 12515 2115
rect 12495 2045 12515 2065
rect 12495 1995 12515 2015
rect 12955 2080 12975 2100
rect 12955 2030 12975 2050
rect 12955 1980 12975 2000
rect 13010 2230 13030 2250
rect 13010 2180 13030 2200
rect 13010 2130 13030 2150
rect 13010 2080 13030 2100
rect 13010 2030 13030 2050
rect 13010 1980 13030 2000
rect 13065 2230 13085 2250
rect 13065 2180 13085 2200
rect 13065 2130 13085 2150
rect 13065 2080 13085 2100
rect 13065 2030 13085 2050
rect 13065 1980 13085 2000
rect 13120 2230 13140 2250
rect 13120 2180 13140 2200
rect 13120 2130 13140 2150
rect 13120 2080 13140 2100
rect 13120 2030 13140 2050
rect 13120 1980 13140 2000
rect 13175 2230 13195 2250
rect 13175 2180 13195 2200
rect 13175 2130 13195 2150
rect 13175 2080 13195 2100
rect 13175 2030 13195 2050
rect 13175 1980 13195 2000
rect 13230 2230 13250 2250
rect 13230 2180 13250 2200
rect 13230 2130 13250 2150
rect 13230 2080 13250 2100
rect 13230 2030 13250 2050
rect 13230 1980 13250 2000
rect 13285 2230 13305 2250
rect 13285 2180 13305 2200
rect 13285 2130 13305 2150
rect 13285 2080 13305 2100
rect 13285 2030 13305 2050
rect 13285 1980 13305 2000
rect 13340 2230 13360 2250
rect 13340 2180 13360 2200
rect 13340 2130 13360 2150
rect 13340 2080 13360 2100
rect 13340 2030 13360 2050
rect 13340 1980 13360 2000
rect 13395 2230 13415 2250
rect 13395 2180 13415 2200
rect 13395 2130 13415 2150
rect 13395 2080 13415 2100
rect 13395 2030 13415 2050
rect 13395 1980 13415 2000
rect 13450 2230 13470 2250
rect 13450 2180 13470 2200
rect 13450 2130 13470 2150
rect 13450 2080 13470 2100
rect 13450 2030 13470 2050
rect 13450 1980 13470 2000
rect 13505 2230 13525 2250
rect 13505 2180 13525 2200
rect 13505 2130 13525 2150
rect 13505 2080 13525 2100
rect 13505 2030 13525 2050
rect 13505 1980 13525 2000
rect 13560 2230 13580 2250
rect 13560 2180 13580 2200
rect 13560 2130 13580 2150
rect 13560 2080 13580 2100
rect 13560 2030 13580 2050
rect 13560 1980 13580 2000
rect 13615 2230 13635 2250
rect 13615 2180 13635 2200
rect 13615 2130 13635 2150
rect 13615 2080 13635 2100
rect 13615 2030 13635 2050
rect 24690 2585 24710 2605
rect 24690 2535 24710 2555
rect 24745 2585 24765 2605
rect 24745 2535 24765 2555
rect 24800 2585 24820 2605
rect 24800 2535 24820 2555
rect 24855 2585 24875 2605
rect 24855 2535 24875 2555
rect 24910 2585 24930 2605
rect 24910 2535 24930 2555
rect 24965 2585 24985 2605
rect 24965 2535 24985 2555
rect 25020 2585 25040 2605
rect 25020 2535 25040 2555
rect 25075 2585 25095 2605
rect 25075 2535 25095 2555
rect 25130 2585 25150 2605
rect 25130 2535 25150 2555
rect 25185 2585 25205 2605
rect 25185 2535 25205 2555
rect 25240 2585 25260 2605
rect 25240 2535 25260 2555
rect 25295 2585 25315 2605
rect 25295 2535 25315 2555
rect 25350 2585 25370 2605
rect 25350 2535 25370 2555
rect 25405 2585 25425 2605
rect 25405 2535 25425 2555
rect 25460 2585 25480 2605
rect 25460 2535 25480 2555
rect 25515 2585 25535 2605
rect 25515 2535 25535 2555
rect 25570 2585 25590 2605
rect 25570 2535 25590 2555
rect 25625 2585 25645 2605
rect 25625 2535 25645 2555
rect 25680 2585 25700 2605
rect 25680 2535 25700 2555
rect 25735 2585 25755 2605
rect 25735 2535 25755 2555
rect 25790 2585 25810 2605
rect 25790 2535 25810 2555
rect 25845 2585 25865 2605
rect 25845 2535 25865 2555
rect 25900 2585 25920 2605
rect 25900 2535 25920 2555
rect 26230 2610 26250 2630
rect 26230 2560 26250 2580
rect 26230 2510 26250 2530
rect 26290 2860 26310 2880
rect 26290 2810 26310 2830
rect 26290 2760 26310 2780
rect 26290 2710 26310 2730
rect 26290 2660 26310 2680
rect 26290 2610 26310 2630
rect 26290 2560 26310 2580
rect 26290 2510 26310 2530
rect 26350 2860 26370 2880
rect 26350 2810 26370 2830
rect 26350 2760 26370 2780
rect 26350 2710 26370 2730
rect 26350 2660 26370 2680
rect 26350 2610 26370 2630
rect 26350 2560 26370 2580
rect 26350 2510 26370 2530
rect 26410 2860 26430 2880
rect 26410 2810 26430 2830
rect 26410 2760 26430 2780
rect 26410 2710 26430 2730
rect 26410 2660 26430 2680
rect 26410 2610 26430 2630
rect 26410 2560 26430 2580
rect 26410 2510 26430 2530
rect 26470 2860 26490 2880
rect 26470 2810 26490 2830
rect 26470 2760 26490 2780
rect 26470 2710 26490 2730
rect 26470 2660 26490 2680
rect 26470 2610 26490 2630
rect 26470 2560 26490 2580
rect 26470 2510 26490 2530
rect 26530 2860 26550 2880
rect 26530 2810 26550 2830
rect 26530 2760 26550 2780
rect 26530 2710 26550 2730
rect 26530 2660 26550 2680
rect 26530 2610 26550 2630
rect 26530 2560 26550 2580
rect 26530 2510 26550 2530
rect 26590 2860 26610 2880
rect 26590 2810 26610 2830
rect 26590 2760 26610 2780
rect 26590 2710 26610 2730
rect 26590 2660 26610 2680
rect 26590 2610 26610 2630
rect 26590 2560 26610 2580
rect 26590 2510 26610 2530
rect 26650 2860 26670 2880
rect 26650 2810 26670 2830
rect 26650 2760 26670 2780
rect 26650 2710 26670 2730
rect 26650 2660 26670 2680
rect 26650 2610 26670 2630
rect 26650 2560 26670 2580
rect 26650 2510 26670 2530
rect 26710 2860 26730 2880
rect 26710 2810 26730 2830
rect 26710 2760 26730 2780
rect 26710 2710 26730 2730
rect 26710 2660 26730 2680
rect 26710 2610 26730 2630
rect 26710 2560 26730 2580
rect 26710 2510 26730 2530
rect 26770 2860 26790 2880
rect 26770 2810 26790 2830
rect 26770 2760 26790 2780
rect 26770 2710 26790 2730
rect 26770 2660 26790 2680
rect 26770 2610 26790 2630
rect 26770 2560 26790 2580
rect 26770 2510 26790 2530
rect 26830 2860 26850 2880
rect 26830 2810 26850 2830
rect 26830 2760 26850 2780
rect 26830 2710 26850 2730
rect 26830 2660 26850 2680
rect 26830 2610 26850 2630
rect 26830 2560 26850 2580
rect 26830 2510 26850 2530
rect 26890 2860 26910 2880
rect 26890 2810 26910 2830
rect 26890 2760 26910 2780
rect 26890 2710 26910 2730
rect 26890 2660 26910 2680
rect 26890 2610 26910 2630
rect 26890 2560 26910 2580
rect 26890 2510 26910 2530
rect 26950 2860 26970 2880
rect 26950 2810 26970 2830
rect 26950 2760 26970 2780
rect 26950 2710 26970 2730
rect 26950 2660 26970 2680
rect 26950 2610 26970 2630
rect 26950 2560 26970 2580
rect 26950 2510 26970 2530
rect 27010 2860 27030 2880
rect 27010 2810 27030 2830
rect 27010 2760 27030 2780
rect 27010 2710 27030 2730
rect 27010 2660 27030 2680
rect 27010 2610 27030 2630
rect 27010 2560 27030 2580
rect 27010 2510 27030 2530
rect 27070 2860 27090 2880
rect 27070 2810 27090 2830
rect 27070 2760 27090 2780
rect 27070 2710 27090 2730
rect 27070 2660 27090 2680
rect 27070 2610 27090 2630
rect 27070 2560 27090 2580
rect 27070 2510 27090 2530
rect 27130 2860 27150 2880
rect 27130 2810 27150 2830
rect 27130 2760 27150 2780
rect 27130 2710 27150 2730
rect 27130 2660 27150 2680
rect 27130 2610 27150 2630
rect 27130 2560 27150 2580
rect 27130 2510 27150 2530
rect 27190 2860 27210 2880
rect 27190 2810 27210 2830
rect 27190 2760 27210 2780
rect 27190 2710 27210 2730
rect 27190 2660 27210 2680
rect 27190 2610 27210 2630
rect 27190 2560 27210 2580
rect 27190 2510 27210 2530
rect 27250 2860 27270 2880
rect 27250 2810 27270 2830
rect 27250 2760 27270 2780
rect 27250 2710 27270 2730
rect 27250 2660 27270 2680
rect 27250 2610 27270 2630
rect 27250 2560 27270 2580
rect 27250 2510 27270 2530
rect 27310 2860 27330 2880
rect 27310 2810 27330 2830
rect 27310 2760 27330 2780
rect 27310 2710 27330 2730
rect 27310 2660 27330 2680
rect 27310 2610 27330 2630
rect 27310 2560 27330 2580
rect 27310 2510 27330 2530
rect 27370 2860 27390 2880
rect 27370 2810 27390 2830
rect 27370 2760 27390 2780
rect 27370 2710 27390 2730
rect 27370 2660 27390 2680
rect 27370 2610 27390 2630
rect 27370 2560 27390 2580
rect 27370 2510 27390 2530
rect 27430 2860 27450 2880
rect 27430 2810 27450 2830
rect 27430 2760 27450 2780
rect 27430 2710 27450 2730
rect 27430 2660 27450 2680
rect 27430 2610 27450 2630
rect 27430 2560 27450 2580
rect 27430 2510 27450 2530
rect 27490 2860 27510 2880
rect 27490 2810 27510 2830
rect 27490 2760 27510 2780
rect 27490 2710 27510 2730
rect 27490 2660 27510 2680
rect 27490 2610 27510 2630
rect 27490 2560 27510 2580
rect 27490 2510 27510 2530
rect 27550 2860 27570 2880
rect 27550 2810 27570 2830
rect 27550 2760 27570 2780
rect 27550 2710 27570 2730
rect 27550 2660 27570 2680
rect 27550 2610 27570 2630
rect 27550 2560 27570 2580
rect 27550 2510 27570 2530
rect 27900 2585 27920 2605
rect 27900 2535 27920 2555
rect 27955 2585 27975 2605
rect 27955 2535 27975 2555
rect 28010 2585 28030 2605
rect 28010 2535 28030 2555
rect 28065 2585 28085 2605
rect 28065 2535 28085 2555
rect 28120 2585 28140 2605
rect 28120 2535 28140 2555
rect 28175 2585 28195 2605
rect 28175 2535 28195 2555
rect 28230 2585 28250 2605
rect 28230 2535 28250 2555
rect 28285 2585 28305 2605
rect 28285 2535 28305 2555
rect 28340 2585 28360 2605
rect 28340 2535 28360 2555
rect 28395 2585 28415 2605
rect 28395 2535 28415 2555
rect 28450 2585 28470 2605
rect 28450 2535 28470 2555
rect 28505 2585 28525 2605
rect 28505 2535 28525 2555
rect 28560 2585 28580 2605
rect 28560 2535 28580 2555
rect 28615 2585 28635 2605
rect 28615 2535 28635 2555
rect 28670 2585 28690 2605
rect 28670 2535 28690 2555
rect 28725 2585 28745 2605
rect 28725 2535 28745 2555
rect 28780 2585 28800 2605
rect 28780 2535 28800 2555
rect 28835 2585 28855 2605
rect 28835 2535 28855 2555
rect 28890 2585 28910 2605
rect 28890 2535 28910 2555
rect 28945 2585 28965 2605
rect 28945 2535 28965 2555
rect 29000 2585 29020 2605
rect 29000 2535 29020 2555
rect 29055 2585 29075 2605
rect 29055 2535 29075 2555
rect 29110 2585 29130 2605
rect 29110 2535 29130 2555
rect 24690 2135 24710 2155
rect 24690 2085 24710 2105
rect 24690 2035 24710 2055
rect 24745 2135 24765 2155
rect 24745 2085 24765 2105
rect 24745 2035 24765 2055
rect 24800 2135 24820 2155
rect 24800 2085 24820 2105
rect 24800 2035 24820 2055
rect 24855 2135 24875 2155
rect 24855 2085 24875 2105
rect 24855 2035 24875 2055
rect 24910 2135 24930 2155
rect 24910 2085 24930 2105
rect 24910 2035 24930 2055
rect 24965 2135 24985 2155
rect 24965 2085 24985 2105
rect 24965 2035 24985 2055
rect 25020 2135 25040 2155
rect 25020 2085 25040 2105
rect 25020 2035 25040 2055
rect 25075 2135 25095 2155
rect 25075 2085 25095 2105
rect 25075 2035 25095 2055
rect 25130 2135 25150 2155
rect 25130 2085 25150 2105
rect 25130 2035 25150 2055
rect 25185 2135 25205 2155
rect 25185 2085 25205 2105
rect 25185 2035 25205 2055
rect 25240 2135 25260 2155
rect 25240 2085 25260 2105
rect 25240 2035 25260 2055
rect 25295 2135 25315 2155
rect 25295 2085 25315 2105
rect 25295 2035 25315 2055
rect 25350 2135 25370 2155
rect 25350 2085 25370 2105
rect 25350 2035 25370 2055
rect 25405 2135 25425 2155
rect 25405 2085 25425 2105
rect 25405 2035 25425 2055
rect 25460 2135 25480 2155
rect 25460 2085 25480 2105
rect 25460 2035 25480 2055
rect 25515 2135 25535 2155
rect 25515 2085 25535 2105
rect 25515 2035 25535 2055
rect 25570 2135 25590 2155
rect 25570 2085 25590 2105
rect 25570 2035 25590 2055
rect 25625 2135 25645 2155
rect 25625 2085 25645 2105
rect 25625 2035 25645 2055
rect 25680 2135 25700 2155
rect 25680 2085 25700 2105
rect 25680 2035 25700 2055
rect 25735 2135 25755 2155
rect 25735 2085 25755 2105
rect 25735 2035 25755 2055
rect 25790 2135 25810 2155
rect 25790 2085 25810 2105
rect 25790 2035 25810 2055
rect 25845 2135 25865 2155
rect 25845 2085 25865 2105
rect 25845 2035 25865 2055
rect 25900 2135 25920 2155
rect 27900 2135 27920 2155
rect 25900 2085 25920 2105
rect 25900 2035 25920 2055
rect 26285 2095 26305 2115
rect 26285 2045 26305 2065
rect 13615 1980 13635 2000
rect 26285 1995 26305 2015
rect 26340 2095 26360 2115
rect 26340 2045 26360 2065
rect 26340 1995 26360 2015
rect 26395 2095 26415 2115
rect 26395 2045 26415 2065
rect 26395 1995 26415 2015
rect 26450 2095 26470 2115
rect 26450 2045 26470 2065
rect 26450 1995 26470 2015
rect 26505 2095 26525 2115
rect 26505 2045 26525 2065
rect 26505 1995 26525 2015
rect 26560 2095 26580 2115
rect 26560 2045 26580 2065
rect 26560 1995 26580 2015
rect 26615 2095 26635 2115
rect 26615 2045 26635 2065
rect 26615 1995 26635 2015
rect 26670 2095 26690 2115
rect 26670 2045 26690 2065
rect 26670 1995 26690 2015
rect 26725 2095 26745 2115
rect 26725 2045 26745 2065
rect 26725 1995 26745 2015
rect 26780 2095 26800 2115
rect 26780 2045 26800 2065
rect 26780 1995 26800 2015
rect 26835 2095 26855 2115
rect 26835 2045 26855 2065
rect 26835 1995 26855 2015
rect 26890 2095 26910 2115
rect 26890 2045 26910 2065
rect 26890 1995 26910 2015
rect 26945 2095 26965 2115
rect 26945 2045 26965 2065
rect 26945 1995 26965 2015
rect 27000 2095 27020 2115
rect 27000 2045 27020 2065
rect 27000 1995 27020 2015
rect 27055 2095 27075 2115
rect 27055 2045 27075 2065
rect 27055 1995 27075 2015
rect 27110 2095 27130 2115
rect 27110 2045 27130 2065
rect 27110 1995 27130 2015
rect 27165 2095 27185 2115
rect 27165 2045 27185 2065
rect 27165 1995 27185 2015
rect 27220 2095 27240 2115
rect 27220 2045 27240 2065
rect 27220 1995 27240 2015
rect 27275 2095 27295 2115
rect 27275 2045 27295 2065
rect 27275 1995 27295 2015
rect 27330 2095 27350 2115
rect 27330 2045 27350 2065
rect 27330 1995 27350 2015
rect 27385 2095 27405 2115
rect 27385 2045 27405 2065
rect 27385 1995 27405 2015
rect 27440 2095 27460 2115
rect 27440 2045 27460 2065
rect 27440 1995 27460 2015
rect 27495 2095 27515 2115
rect 27495 2045 27515 2065
rect 27900 2085 27920 2105
rect 27900 2035 27920 2055
rect 27955 2135 27975 2155
rect 27955 2085 27975 2105
rect 27955 2035 27975 2055
rect 28010 2135 28030 2155
rect 28010 2085 28030 2105
rect 28010 2035 28030 2055
rect 28065 2135 28085 2155
rect 28065 2085 28085 2105
rect 28065 2035 28085 2055
rect 28120 2135 28140 2155
rect 28120 2085 28140 2105
rect 28120 2035 28140 2055
rect 28175 2135 28195 2155
rect 28175 2085 28195 2105
rect 28175 2035 28195 2055
rect 28230 2135 28250 2155
rect 28230 2085 28250 2105
rect 28230 2035 28250 2055
rect 28285 2135 28305 2155
rect 28285 2085 28305 2105
rect 28285 2035 28305 2055
rect 28340 2135 28360 2155
rect 28340 2085 28360 2105
rect 28340 2035 28360 2055
rect 28395 2135 28415 2155
rect 28395 2085 28415 2105
rect 28395 2035 28415 2055
rect 28450 2135 28470 2155
rect 28450 2085 28470 2105
rect 28450 2035 28470 2055
rect 28505 2135 28525 2155
rect 28505 2085 28525 2105
rect 28505 2035 28525 2055
rect 28560 2135 28580 2155
rect 28560 2085 28580 2105
rect 28560 2035 28580 2055
rect 28615 2135 28635 2155
rect 28615 2085 28635 2105
rect 28615 2035 28635 2055
rect 28670 2135 28690 2155
rect 28670 2085 28690 2105
rect 28670 2035 28690 2055
rect 28725 2135 28745 2155
rect 28725 2085 28745 2105
rect 28725 2035 28745 2055
rect 28780 2135 28800 2155
rect 28780 2085 28800 2105
rect 28780 2035 28800 2055
rect 28835 2135 28855 2155
rect 28835 2085 28855 2105
rect 28835 2035 28855 2055
rect 28890 2135 28910 2155
rect 28890 2085 28910 2105
rect 28890 2035 28910 2055
rect 28945 2135 28965 2155
rect 28945 2085 28965 2105
rect 28945 2035 28965 2055
rect 29000 2135 29020 2155
rect 29000 2085 29020 2105
rect 29000 2035 29020 2055
rect 29055 2135 29075 2155
rect 29055 2085 29075 2105
rect 29055 2035 29075 2055
rect 29110 2135 29130 2155
rect 29110 2085 29130 2105
rect 29110 2035 29130 2055
rect 27495 1995 27515 2015
rect 28000 1820 28020 1840
rect 28000 1770 28020 1790
rect 28000 1720 28020 1740
rect 28055 1820 28075 1840
rect 28055 1770 28075 1790
rect 28055 1720 28075 1740
rect 28110 1820 28130 1840
rect 28110 1770 28130 1790
rect 28110 1720 28130 1740
rect 28165 1820 28185 1840
rect 28165 1770 28185 1790
rect 28165 1720 28185 1740
rect 28220 1820 28240 1840
rect 28220 1770 28240 1790
rect 28220 1720 28240 1740
rect 28275 1820 28295 1840
rect 28275 1770 28295 1790
rect 28275 1720 28295 1740
rect 28330 1820 28350 1840
rect 28330 1770 28350 1790
rect 28330 1720 28350 1740
rect 3175 1630 3195 1650
rect 3235 1630 3255 1650
rect 3295 1630 3315 1650
rect 3355 1630 3375 1650
rect 3415 1630 3435 1650
rect 3475 1630 3495 1650
rect 3535 1630 3555 1650
rect 3595 1630 3615 1650
rect 3655 1630 3675 1650
rect 3715 1630 3735 1650
rect 3775 1630 3795 1650
rect 4215 1630 4235 1650
rect 4275 1630 4295 1650
rect 4335 1630 4355 1650
rect 4395 1630 4415 1650
rect 4455 1630 4475 1650
rect 4515 1630 4535 1650
rect 4575 1630 4595 1650
rect 4635 1630 4655 1650
rect 4695 1630 4715 1650
rect 4755 1630 4775 1650
rect 4815 1630 4835 1650
rect 10165 1620 10185 1640
rect 2845 1420 2865 1440
rect 2845 1370 2865 1390
rect 2845 1320 2865 1340
rect 2845 1270 2865 1290
rect 2845 1220 2865 1240
rect 3385 1420 3405 1440
rect 3385 1370 3405 1390
rect 3385 1320 3405 1340
rect 3385 1270 3405 1290
rect 3385 1220 3405 1240
rect 3925 1420 3945 1440
rect 3925 1370 3945 1390
rect 3925 1320 3945 1340
rect 3925 1270 3945 1290
rect 3925 1220 3945 1240
rect 4065 1420 4085 1440
rect 4065 1370 4085 1390
rect 4065 1320 4085 1340
rect 4065 1270 4085 1290
rect 4065 1220 4085 1240
rect 4605 1420 4625 1440
rect 4605 1370 4625 1390
rect 4605 1320 4625 1340
rect 4605 1270 4625 1290
rect 4605 1220 4625 1240
rect 5145 1420 5165 1440
rect 5145 1370 5165 1390
rect 5145 1320 5165 1340
rect 5145 1270 5165 1290
rect 5145 1220 5165 1240
rect 2955 1040 2975 1060
rect 2955 990 2975 1010
rect 3995 1040 4015 1060
rect 3995 990 4015 1010
rect 5035 1040 5055 1060
rect 5035 990 5055 1010
rect 10165 1570 10185 1590
rect 10165 1520 10185 1540
rect 10165 1470 10185 1490
rect 10165 1420 10185 1440
rect 10165 1370 10185 1390
rect 10165 1320 10185 1340
rect 10165 1270 10185 1290
rect 10165 1220 10185 1240
rect 10165 1170 10185 1190
rect 10165 1120 10185 1140
rect 10165 1070 10185 1090
rect 10165 1020 10185 1040
rect 10165 970 10185 990
rect 10265 1620 10285 1640
rect 10265 1570 10285 1590
rect 10265 1520 10285 1540
rect 10265 1470 10285 1490
rect 10265 1420 10285 1440
rect 10265 1370 10285 1390
rect 10265 1320 10285 1340
rect 10265 1270 10285 1290
rect 10265 1220 10285 1240
rect 10265 1170 10285 1190
rect 10265 1120 10285 1140
rect 10265 1070 10285 1090
rect 10265 1020 10285 1040
rect 10265 970 10285 990
rect 10365 1620 10385 1640
rect 10365 1570 10385 1590
rect 10365 1520 10385 1540
rect 10365 1470 10385 1490
rect 10365 1420 10385 1440
rect 10365 1370 10385 1390
rect 10365 1320 10385 1340
rect 10365 1270 10385 1290
rect 10365 1220 10385 1240
rect 10365 1170 10385 1190
rect 10365 1120 10385 1140
rect 10365 1070 10385 1090
rect 10365 1020 10385 1040
rect 10365 970 10385 990
rect 10465 1620 10485 1640
rect 10465 1570 10485 1590
rect 10465 1520 10485 1540
rect 10465 1470 10485 1490
rect 10465 1420 10485 1440
rect 10465 1370 10485 1390
rect 10465 1320 10485 1340
rect 10465 1270 10485 1290
rect 10465 1220 10485 1240
rect 10465 1170 10485 1190
rect 10465 1120 10485 1140
rect 10465 1070 10485 1090
rect 10465 1020 10485 1040
rect 10465 970 10485 990
rect 10565 1620 10585 1640
rect 10565 1570 10585 1590
rect 10565 1520 10585 1540
rect 10565 1470 10585 1490
rect 10565 1420 10585 1440
rect 10565 1370 10585 1390
rect 10565 1320 10585 1340
rect 10565 1270 10585 1290
rect 10565 1220 10585 1240
rect 10565 1170 10585 1190
rect 10565 1120 10585 1140
rect 10565 1070 10585 1090
rect 10565 1020 10585 1040
rect 10565 970 10585 990
rect 10665 1620 10685 1640
rect 10665 1570 10685 1590
rect 10665 1520 10685 1540
rect 10665 1470 10685 1490
rect 10665 1420 10685 1440
rect 10665 1370 10685 1390
rect 10665 1320 10685 1340
rect 10665 1270 10685 1290
rect 10665 1220 10685 1240
rect 10665 1170 10685 1190
rect 10665 1120 10685 1140
rect 10665 1070 10685 1090
rect 10665 1020 10685 1040
rect 10665 970 10685 990
rect 10765 1620 10785 1640
rect 10765 1570 10785 1590
rect 10765 1520 10785 1540
rect 11040 1630 11060 1650
rect 11040 1580 11060 1600
rect 11040 1530 11060 1550
rect 11095 1630 11115 1650
rect 11095 1580 11115 1600
rect 11095 1530 11115 1550
rect 11150 1630 11170 1650
rect 11150 1580 11170 1600
rect 11150 1530 11170 1550
rect 11205 1630 11225 1650
rect 11205 1580 11225 1600
rect 11205 1530 11225 1550
rect 11260 1630 11280 1650
rect 11260 1580 11280 1600
rect 11260 1530 11280 1550
rect 11315 1630 11335 1650
rect 11315 1580 11335 1600
rect 11315 1530 11335 1550
rect 11370 1630 11390 1650
rect 11370 1580 11390 1600
rect 11370 1530 11390 1550
rect 11425 1630 11445 1650
rect 11425 1580 11445 1600
rect 11425 1530 11445 1550
rect 11480 1630 11500 1650
rect 11480 1580 11500 1600
rect 11480 1530 11500 1550
rect 11535 1630 11555 1650
rect 11535 1580 11555 1600
rect 11535 1530 11555 1550
rect 11590 1630 11610 1650
rect 11590 1580 11610 1600
rect 11590 1530 11610 1550
rect 11645 1630 11665 1650
rect 11645 1580 11665 1600
rect 11645 1530 11665 1550
rect 11700 1630 11720 1650
rect 11780 1630 11800 1650
rect 11700 1580 11720 1600
rect 11780 1580 11800 1600
rect 11700 1530 11720 1550
rect 11780 1530 11800 1550
rect 11835 1630 11855 1650
rect 11835 1580 11855 1600
rect 11835 1530 11855 1550
rect 11890 1630 11910 1650
rect 11890 1580 11910 1600
rect 11890 1530 11910 1550
rect 11945 1630 11965 1650
rect 11945 1580 11965 1600
rect 11945 1530 11965 1550
rect 12000 1630 12020 1650
rect 12080 1630 12100 1650
rect 12000 1580 12020 1600
rect 12080 1580 12100 1600
rect 12000 1530 12020 1550
rect 12080 1530 12100 1550
rect 12135 1630 12155 1650
rect 12135 1580 12155 1600
rect 12135 1530 12155 1550
rect 12190 1630 12210 1650
rect 12190 1580 12210 1600
rect 12190 1530 12210 1550
rect 12245 1630 12265 1650
rect 12245 1580 12265 1600
rect 12245 1530 12265 1550
rect 12300 1630 12320 1650
rect 12300 1580 12320 1600
rect 12300 1530 12320 1550
rect 12355 1630 12375 1650
rect 12355 1580 12375 1600
rect 12355 1530 12375 1550
rect 12410 1630 12430 1650
rect 12410 1580 12430 1600
rect 12410 1530 12430 1550
rect 12465 1630 12485 1650
rect 12465 1580 12485 1600
rect 12465 1530 12485 1550
rect 12520 1630 12540 1650
rect 12520 1580 12540 1600
rect 12520 1530 12540 1550
rect 12575 1630 12595 1650
rect 12575 1580 12595 1600
rect 12575 1530 12595 1550
rect 12630 1630 12650 1650
rect 12630 1580 12650 1600
rect 12630 1530 12650 1550
rect 12685 1630 12705 1650
rect 12685 1580 12705 1600
rect 12685 1530 12705 1550
rect 12740 1630 12760 1650
rect 12740 1580 12760 1600
rect 12740 1530 12760 1550
rect 13015 1620 13035 1640
rect 13015 1570 13035 1590
rect 13015 1520 13035 1540
rect 10765 1470 10785 1490
rect 13015 1470 13035 1490
rect 10765 1420 10785 1440
rect 10765 1370 10785 1390
rect 10765 1320 10785 1340
rect 10765 1270 10785 1290
rect 13015 1420 13035 1440
rect 13015 1370 13035 1390
rect 13015 1320 13035 1340
rect 13015 1270 13035 1290
rect 10765 1220 10785 1240
rect 10765 1170 10785 1190
rect 13015 1220 13035 1240
rect 10765 1120 10785 1140
rect 10765 1070 10785 1090
rect 10765 1020 10785 1040
rect 10765 970 10785 990
rect 11215 1150 11235 1170
rect 11215 1100 11235 1120
rect 11215 1050 11235 1070
rect 11215 1000 11235 1020
rect 11215 950 11235 970
rect 11270 1150 11290 1170
rect 11270 1100 11290 1120
rect 11270 1050 11290 1070
rect 11270 1000 11290 1020
rect 11270 950 11290 970
rect 11325 1150 11345 1170
rect 11325 1100 11345 1120
rect 11325 1050 11345 1070
rect 11325 1000 11345 1020
rect 11325 950 11345 970
rect 11380 1150 11400 1170
rect 11380 1100 11400 1120
rect 11380 1050 11400 1070
rect 11380 1000 11400 1020
rect 11380 950 11400 970
rect 11435 1150 11455 1170
rect 11435 1100 11455 1120
rect 11435 1050 11455 1070
rect 11435 1000 11455 1020
rect 11435 950 11455 970
rect 11490 1150 11510 1170
rect 11490 1100 11510 1120
rect 11490 1050 11510 1070
rect 11490 1000 11510 1020
rect 11490 950 11510 970
rect 11545 1150 11565 1170
rect 11545 1100 11565 1120
rect 11545 1050 11565 1070
rect 11545 1000 11565 1020
rect 11545 950 11565 970
rect 11600 1150 11620 1170
rect 11600 1100 11620 1120
rect 11600 1050 11620 1070
rect 11600 1000 11620 1020
rect 11600 950 11620 970
rect 11655 1150 11675 1170
rect 11655 1100 11675 1120
rect 11655 1050 11675 1070
rect 11655 1000 11675 1020
rect 11655 950 11675 970
rect 11710 1150 11730 1170
rect 11710 1100 11730 1120
rect 11710 1050 11730 1070
rect 11710 1000 11730 1020
rect 11710 950 11730 970
rect 11765 1150 11785 1170
rect 11765 1100 11785 1120
rect 11765 1050 11785 1070
rect 11765 1000 11785 1020
rect 11765 950 11785 970
rect 11820 1150 11840 1170
rect 11820 1100 11840 1120
rect 11820 1050 11840 1070
rect 11820 1000 11840 1020
rect 11820 950 11840 970
rect 11875 1150 11895 1170
rect 11875 1100 11895 1120
rect 11875 1050 11895 1070
rect 11875 1000 11895 1020
rect 11875 950 11895 970
rect 11930 1150 11950 1170
rect 11930 1100 11950 1120
rect 11930 1050 11950 1070
rect 11930 1000 11950 1020
rect 11930 950 11950 970
rect 11985 1150 12005 1170
rect 11985 1100 12005 1120
rect 11985 1050 12005 1070
rect 11985 1000 12005 1020
rect 11985 950 12005 970
rect 12040 1150 12060 1170
rect 12040 1100 12060 1120
rect 12040 1050 12060 1070
rect 12040 1000 12060 1020
rect 12040 950 12060 970
rect 12095 1150 12115 1170
rect 12095 1100 12115 1120
rect 12095 1050 12115 1070
rect 12095 1000 12115 1020
rect 12095 950 12115 970
rect 12150 1150 12170 1170
rect 12150 1100 12170 1120
rect 12150 1050 12170 1070
rect 12150 1000 12170 1020
rect 12150 950 12170 970
rect 12205 1150 12225 1170
rect 12205 1100 12225 1120
rect 12205 1050 12225 1070
rect 12205 1000 12225 1020
rect 12205 950 12225 970
rect 12260 1150 12280 1170
rect 12260 1100 12280 1120
rect 12260 1050 12280 1070
rect 12260 1000 12280 1020
rect 12260 950 12280 970
rect 12315 1150 12335 1170
rect 12315 1100 12335 1120
rect 12315 1050 12335 1070
rect 12315 1000 12335 1020
rect 12315 950 12335 970
rect 12370 1150 12390 1170
rect 12370 1100 12390 1120
rect 12370 1050 12390 1070
rect 12370 1000 12390 1020
rect 12370 950 12390 970
rect 12425 1150 12445 1170
rect 12425 1100 12445 1120
rect 12425 1050 12445 1070
rect 12425 1000 12445 1020
rect 12425 950 12445 970
rect 12480 1150 12500 1170
rect 12480 1100 12500 1120
rect 12480 1050 12500 1070
rect 12480 1000 12500 1020
rect 12480 950 12500 970
rect 12535 1150 12555 1170
rect 12535 1100 12555 1120
rect 12535 1050 12555 1070
rect 12535 1000 12555 1020
rect 12535 950 12555 970
rect 12590 1150 12610 1170
rect 12590 1100 12610 1120
rect 12590 1050 12610 1070
rect 12590 1000 12610 1020
rect 12590 950 12610 970
rect 13015 1170 13035 1190
rect 13015 1120 13035 1140
rect 13015 1070 13035 1090
rect 13015 1020 13035 1040
rect 13015 970 13035 990
rect 13115 1620 13135 1640
rect 13115 1570 13135 1590
rect 13115 1520 13135 1540
rect 13115 1470 13135 1490
rect 13115 1420 13135 1440
rect 13115 1370 13135 1390
rect 13115 1320 13135 1340
rect 13115 1270 13135 1290
rect 13115 1220 13135 1240
rect 13115 1170 13135 1190
rect 13115 1120 13135 1140
rect 13115 1070 13135 1090
rect 13115 1020 13135 1040
rect 13115 970 13135 990
rect 13215 1620 13235 1640
rect 13215 1570 13235 1590
rect 13215 1520 13235 1540
rect 13215 1470 13235 1490
rect 13215 1420 13235 1440
rect 13215 1370 13235 1390
rect 13215 1320 13235 1340
rect 13215 1270 13235 1290
rect 13215 1220 13235 1240
rect 13215 1170 13235 1190
rect 13215 1120 13235 1140
rect 13215 1070 13235 1090
rect 13215 1020 13235 1040
rect 13215 970 13235 990
rect 13315 1620 13335 1640
rect 13315 1570 13335 1590
rect 13315 1520 13335 1540
rect 13315 1470 13335 1490
rect 13315 1420 13335 1440
rect 13315 1370 13335 1390
rect 13315 1320 13335 1340
rect 13315 1270 13335 1290
rect 13315 1220 13335 1240
rect 13315 1170 13335 1190
rect 13315 1120 13335 1140
rect 13315 1070 13335 1090
rect 13315 1020 13335 1040
rect 13315 970 13335 990
rect 13415 1620 13435 1640
rect 13415 1570 13435 1590
rect 13415 1520 13435 1540
rect 13415 1470 13435 1490
rect 13415 1420 13435 1440
rect 13415 1370 13435 1390
rect 13415 1320 13435 1340
rect 13415 1270 13435 1290
rect 13415 1220 13435 1240
rect 13415 1170 13435 1190
rect 13415 1120 13435 1140
rect 13415 1070 13435 1090
rect 13415 1020 13435 1040
rect 13415 970 13435 990
rect 13515 1620 13535 1640
rect 13515 1570 13535 1590
rect 13515 1520 13535 1540
rect 13515 1470 13535 1490
rect 13515 1420 13535 1440
rect 13515 1370 13535 1390
rect 13515 1320 13535 1340
rect 13515 1270 13535 1290
rect 13515 1220 13535 1240
rect 13515 1170 13535 1190
rect 13515 1120 13535 1140
rect 13515 1070 13535 1090
rect 13515 1020 13535 1040
rect 13515 970 13535 990
rect 13615 1620 13635 1640
rect 26040 1630 26060 1650
rect 13615 1570 13635 1590
rect 13615 1520 13635 1540
rect 13615 1470 13635 1490
rect 13615 1420 13635 1440
rect 13615 1370 13635 1390
rect 13615 1320 13635 1340
rect 13615 1270 13635 1290
rect 13615 1220 13635 1240
rect 13615 1170 13635 1190
rect 13615 1120 13635 1140
rect 13615 1070 13635 1090
rect 13615 1020 13635 1040
rect 13615 970 13635 990
rect 26040 1580 26060 1600
rect 26040 1530 26060 1550
rect 26095 1630 26115 1650
rect 26095 1580 26115 1600
rect 26095 1530 26115 1550
rect 26150 1630 26170 1650
rect 26150 1580 26170 1600
rect 26150 1530 26170 1550
rect 26205 1630 26225 1650
rect 26205 1580 26225 1600
rect 26205 1530 26225 1550
rect 26260 1630 26280 1650
rect 26260 1580 26280 1600
rect 26260 1530 26280 1550
rect 26315 1630 26335 1650
rect 26315 1580 26335 1600
rect 26315 1530 26335 1550
rect 26370 1630 26390 1650
rect 26370 1580 26390 1600
rect 26370 1530 26390 1550
rect 26425 1630 26445 1650
rect 26425 1580 26445 1600
rect 26425 1530 26445 1550
rect 26480 1630 26500 1650
rect 26480 1580 26500 1600
rect 26480 1530 26500 1550
rect 26535 1630 26555 1650
rect 26535 1580 26555 1600
rect 26535 1530 26555 1550
rect 26590 1630 26610 1650
rect 26590 1580 26610 1600
rect 26590 1530 26610 1550
rect 26645 1630 26665 1650
rect 26645 1580 26665 1600
rect 26645 1530 26665 1550
rect 26700 1630 26720 1650
rect 26780 1630 26800 1650
rect 26700 1580 26720 1600
rect 26780 1580 26800 1600
rect 26700 1530 26720 1550
rect 26780 1530 26800 1550
rect 26835 1630 26855 1650
rect 26835 1580 26855 1600
rect 26835 1530 26855 1550
rect 26890 1630 26910 1650
rect 26890 1580 26910 1600
rect 26890 1530 26910 1550
rect 26945 1630 26965 1650
rect 26945 1580 26965 1600
rect 26945 1530 26965 1550
rect 27000 1630 27020 1650
rect 27080 1630 27100 1650
rect 27000 1580 27020 1600
rect 27080 1580 27100 1600
rect 27000 1530 27020 1550
rect 27080 1530 27100 1550
rect 27135 1630 27155 1650
rect 27135 1580 27155 1600
rect 27135 1530 27155 1550
rect 27190 1630 27210 1650
rect 27190 1580 27210 1600
rect 27190 1530 27210 1550
rect 27245 1630 27265 1650
rect 27245 1580 27265 1600
rect 27245 1530 27265 1550
rect 27300 1630 27320 1650
rect 27300 1580 27320 1600
rect 27300 1530 27320 1550
rect 27355 1630 27375 1650
rect 27355 1580 27375 1600
rect 27355 1530 27375 1550
rect 27410 1630 27430 1650
rect 27410 1580 27430 1600
rect 27410 1530 27430 1550
rect 27465 1630 27485 1650
rect 27465 1580 27485 1600
rect 27465 1530 27485 1550
rect 27520 1630 27540 1650
rect 27520 1580 27540 1600
rect 27520 1530 27540 1550
rect 27575 1630 27595 1650
rect 27575 1580 27595 1600
rect 27575 1530 27595 1550
rect 27630 1630 27650 1650
rect 27630 1580 27650 1600
rect 27630 1530 27650 1550
rect 27685 1630 27705 1650
rect 27685 1580 27705 1600
rect 27685 1530 27705 1550
rect 27740 1630 27760 1650
rect 27740 1580 27760 1600
rect 27740 1530 27760 1550
rect 27905 1485 27925 1505
rect 27905 1435 27925 1455
rect 27905 1385 27925 1405
rect 27960 1485 27980 1505
rect 27960 1435 27980 1455
rect 27960 1385 27980 1405
rect 28015 1485 28035 1505
rect 28015 1435 28035 1455
rect 28015 1385 28035 1405
rect 28070 1485 28090 1505
rect 28070 1435 28090 1455
rect 28070 1385 28090 1405
rect 28125 1485 28145 1505
rect 28205 1485 28225 1505
rect 28125 1435 28145 1455
rect 28205 1435 28225 1455
rect 28125 1385 28145 1405
rect 28205 1385 28225 1405
rect 28260 1485 28280 1505
rect 28260 1435 28280 1455
rect 28260 1385 28280 1405
rect 28315 1485 28335 1505
rect 28315 1435 28335 1455
rect 28315 1385 28335 1405
rect 28370 1485 28390 1505
rect 28370 1435 28390 1455
rect 28370 1385 28390 1405
rect 28425 1485 28445 1505
rect 28425 1435 28445 1455
rect 28425 1385 28445 1405
rect 26215 1190 26235 1210
rect 26215 1140 26235 1160
rect 26215 1090 26235 1110
rect 26215 1040 26235 1060
rect 26215 990 26235 1010
rect 26270 1190 26290 1210
rect 26270 1140 26290 1160
rect 26270 1090 26290 1110
rect 26270 1040 26290 1060
rect 26270 990 26290 1010
rect 26325 1190 26345 1210
rect 26325 1140 26345 1160
rect 26325 1090 26345 1110
rect 26325 1040 26345 1060
rect 26325 990 26345 1010
rect 26380 1190 26400 1210
rect 26380 1140 26400 1160
rect 26380 1090 26400 1110
rect 26380 1040 26400 1060
rect 26380 990 26400 1010
rect 26435 1190 26455 1210
rect 26435 1140 26455 1160
rect 26435 1090 26455 1110
rect 26435 1040 26455 1060
rect 26435 990 26455 1010
rect 26490 1190 26510 1210
rect 26490 1140 26510 1160
rect 26490 1090 26510 1110
rect 26490 1040 26510 1060
rect 26490 990 26510 1010
rect 26545 1190 26565 1210
rect 26545 1140 26565 1160
rect 26545 1090 26565 1110
rect 26545 1040 26565 1060
rect 26545 990 26565 1010
rect 26600 1190 26620 1210
rect 26600 1140 26620 1160
rect 26600 1090 26620 1110
rect 26600 1040 26620 1060
rect 26600 990 26620 1010
rect 26655 1190 26675 1210
rect 26655 1140 26675 1160
rect 26655 1090 26675 1110
rect 26655 1040 26675 1060
rect 26655 990 26675 1010
rect 26710 1190 26730 1210
rect 26710 1140 26730 1160
rect 26710 1090 26730 1110
rect 26710 1040 26730 1060
rect 26710 990 26730 1010
rect 26765 1190 26785 1210
rect 26765 1140 26785 1160
rect 26765 1090 26785 1110
rect 26765 1040 26785 1060
rect 26765 990 26785 1010
rect 26820 1190 26840 1210
rect 26820 1140 26840 1160
rect 26820 1090 26840 1110
rect 26820 1040 26840 1060
rect 26820 990 26840 1010
rect 26875 1190 26895 1210
rect 26875 1140 26895 1160
rect 26875 1090 26895 1110
rect 26875 1040 26895 1060
rect 26875 990 26895 1010
rect 26930 1190 26950 1210
rect 26930 1140 26950 1160
rect 26930 1090 26950 1110
rect 26930 1040 26950 1060
rect 26930 990 26950 1010
rect 26985 1190 27005 1210
rect 26985 1140 27005 1160
rect 26985 1090 27005 1110
rect 26985 1040 27005 1060
rect 26985 990 27005 1010
rect 27040 1190 27060 1210
rect 27040 1140 27060 1160
rect 27040 1090 27060 1110
rect 27040 1040 27060 1060
rect 27040 990 27060 1010
rect 27095 1190 27115 1210
rect 27095 1140 27115 1160
rect 27095 1090 27115 1110
rect 27095 1040 27115 1060
rect 27095 990 27115 1010
rect 27150 1190 27170 1210
rect 27150 1140 27170 1160
rect 27150 1090 27170 1110
rect 27150 1040 27170 1060
rect 27150 990 27170 1010
rect 27205 1190 27225 1210
rect 27205 1140 27225 1160
rect 27205 1090 27225 1110
rect 27205 1040 27225 1060
rect 27205 990 27225 1010
rect 27260 1190 27280 1210
rect 27260 1140 27280 1160
rect 27260 1090 27280 1110
rect 27260 1040 27280 1060
rect 27260 990 27280 1010
rect 27315 1190 27335 1210
rect 27315 1140 27335 1160
rect 27315 1090 27335 1110
rect 27315 1040 27335 1060
rect 27315 990 27335 1010
rect 27370 1190 27390 1210
rect 27370 1140 27390 1160
rect 27370 1090 27390 1110
rect 27370 1040 27390 1060
rect 27370 990 27390 1010
rect 27425 1190 27445 1210
rect 27425 1140 27445 1160
rect 27425 1090 27445 1110
rect 27425 1040 27445 1060
rect 27425 990 27445 1010
rect 27480 1190 27500 1210
rect 27480 1140 27500 1160
rect 27480 1090 27500 1110
rect 27480 1040 27500 1060
rect 27480 990 27500 1010
rect 27535 1190 27555 1210
rect 27535 1140 27555 1160
rect 27535 1090 27555 1110
rect 27535 1040 27555 1060
rect 27535 990 27555 1010
rect 27590 1190 27610 1210
rect 27590 1140 27610 1160
rect 27590 1090 27610 1110
rect 27590 1040 27610 1060
rect 28055 1145 28075 1165
rect 28055 1095 28075 1115
rect 28055 1045 28075 1065
rect 28110 1145 28130 1165
rect 28110 1095 28130 1115
rect 28110 1045 28130 1065
rect 28165 1145 28185 1165
rect 28165 1095 28185 1115
rect 28165 1045 28185 1065
rect 28220 1145 28240 1165
rect 28220 1095 28240 1115
rect 28220 1045 28240 1065
rect 28275 1145 28295 1165
rect 28275 1095 28295 1115
rect 28275 1045 28295 1065
rect 27590 990 27610 1010
rect 3005 845 3025 865
rect 3005 795 3025 815
rect 3095 845 3115 865
rect 3095 795 3115 815
rect 3185 845 3205 865
rect 3185 795 3205 815
rect 3275 845 3295 865
rect 3275 795 3295 815
rect 3365 845 3385 865
rect 3365 795 3385 815
rect 3455 845 3475 865
rect 3455 795 3475 815
rect 3545 845 3565 865
rect 3545 795 3565 815
rect 3635 845 3655 865
rect 3635 795 3655 815
rect 3725 845 3745 865
rect 3725 795 3745 815
rect 3815 845 3835 865
rect 3815 795 3835 815
rect 3905 845 3925 865
rect 3905 795 3925 815
rect 3995 845 4015 865
rect 3995 795 4015 815
rect 4085 845 4105 865
rect 4085 795 4105 815
rect 4175 845 4195 865
rect 4175 795 4195 815
rect 4265 845 4285 865
rect 4265 795 4285 815
rect 4355 845 4375 865
rect 4355 795 4375 815
rect 4445 845 4465 865
rect 4445 795 4465 815
rect 4535 845 4555 865
rect 4535 795 4555 815
rect 4625 845 4645 865
rect 4625 795 4645 815
rect 4715 845 4735 865
rect 4715 795 4735 815
rect 4805 845 4825 865
rect 4805 795 4825 815
rect 4895 845 4915 865
rect 4895 795 4915 815
rect 4985 845 5005 865
rect 4985 795 5005 815
rect 11270 710 11290 730
rect 11270 660 11290 680
rect 11500 710 11520 730
rect 11890 715 11910 735
rect 11945 715 11965 735
rect 12000 715 12020 735
rect 12055 715 12075 735
rect 12110 715 12130 735
rect 12165 715 12185 735
rect 12220 715 12240 735
rect 12275 715 12295 735
rect 12330 715 12350 735
rect 12385 715 12405 735
rect 12440 715 12460 735
rect 12495 715 12515 735
rect 12550 715 12570 735
rect 11500 660 11520 680
rect 10830 -1505 10850 -1485
rect 10830 -1555 10850 -1535
rect 10830 -1605 10850 -1585
rect 10830 -1655 10850 -1635
rect 10830 -1705 10850 -1685
rect 10500 -1755 10520 -1735
rect 10560 -1750 10580 -1730
rect 10620 -1750 10640 -1730
rect 10680 -1755 10700 -1735
rect 10830 -1755 10850 -1735
rect 10890 -1505 10910 -1485
rect 10890 -1555 10910 -1535
rect 10890 -1605 10910 -1585
rect 10890 -1655 10910 -1635
rect 10890 -1705 10910 -1685
rect 10890 -1755 10910 -1735
rect 10950 -1505 10970 -1485
rect 10950 -1555 10970 -1535
rect 10950 -1605 10970 -1585
rect 10950 -1655 10970 -1635
rect 10950 -1705 10970 -1685
rect 10950 -1755 10970 -1735
rect 11010 -1455 11030 -1435
rect 11010 -1505 11030 -1485
rect 11010 -1555 11030 -1535
rect 11010 -1605 11030 -1585
rect 11010 -1655 11030 -1635
rect 11010 -1705 11030 -1685
rect 11010 -1755 11030 -1735
rect 11070 -1455 11090 -1435
rect 11070 -1505 11090 -1485
rect 11070 -1555 11090 -1535
rect 11070 -1605 11090 -1585
rect 11070 -1655 11090 -1635
rect 11070 -1705 11090 -1685
rect 11070 -1755 11090 -1735
rect 11230 -1460 11250 -1440
rect 11230 -1510 11250 -1490
rect 11230 -1560 11250 -1540
rect 11230 -1610 11250 -1590
rect 11230 -1660 11250 -1640
rect 11230 -1710 11250 -1690
rect 11230 -1760 11250 -1740
rect 11230 -1810 11250 -1790
rect 11290 -1460 11310 -1440
rect 11290 -1510 11310 -1490
rect 11290 -1560 11310 -1540
rect 11290 -1610 11310 -1590
rect 11290 -1660 11310 -1640
rect 11290 -1710 11310 -1690
rect 11290 -1760 11310 -1740
rect 11290 -1810 11310 -1790
rect 11350 -1460 11370 -1440
rect 11350 -1510 11370 -1490
rect 11350 -1560 11370 -1540
rect 11350 -1610 11370 -1590
rect 11350 -1660 11370 -1640
rect 11350 -1710 11370 -1690
rect 11350 -1760 11370 -1740
rect 11350 -1810 11370 -1790
rect 11410 -1460 11430 -1440
rect 11410 -1510 11430 -1490
rect 11410 -1560 11430 -1540
rect 11410 -1610 11430 -1590
rect 11410 -1660 11430 -1640
rect 11410 -1710 11430 -1690
rect 11410 -1760 11430 -1740
rect 11410 -1810 11430 -1790
rect 11470 -1460 11490 -1440
rect 11470 -1510 11490 -1490
rect 11470 -1560 11490 -1540
rect 11470 -1610 11490 -1590
rect 11470 -1660 11490 -1640
rect 11470 -1710 11490 -1690
rect 11470 -1760 11490 -1740
rect 11470 -1810 11490 -1790
rect 11530 -1460 11550 -1440
rect 11530 -1510 11550 -1490
rect 11530 -1560 11550 -1540
rect 11530 -1610 11550 -1590
rect 11530 -1660 11550 -1640
rect 11530 -1710 11550 -1690
rect 11530 -1760 11550 -1740
rect 11530 -1810 11550 -1790
rect 11590 -1460 11610 -1440
rect 11590 -1510 11610 -1490
rect 11590 -1560 11610 -1540
rect 11590 -1610 11610 -1590
rect 11590 -1660 11610 -1640
rect 11590 -1710 11610 -1690
rect 11590 -1760 11610 -1740
rect 11590 -1810 11610 -1790
rect 11650 -1460 11670 -1440
rect 11650 -1510 11670 -1490
rect 11650 -1560 11670 -1540
rect 11650 -1610 11670 -1590
rect 11650 -1660 11670 -1640
rect 11650 -1710 11670 -1690
rect 11650 -1760 11670 -1740
rect 11650 -1810 11670 -1790
rect 11710 -1460 11730 -1440
rect 11710 -1510 11730 -1490
rect 11710 -1560 11730 -1540
rect 11710 -1610 11730 -1590
rect 11710 -1660 11730 -1640
rect 11710 -1710 11730 -1690
rect 11710 -1760 11730 -1740
rect 11710 -1810 11730 -1790
rect 11770 -1460 11790 -1440
rect 11770 -1510 11790 -1490
rect 11770 -1560 11790 -1540
rect 11770 -1610 11790 -1590
rect 11770 -1660 11790 -1640
rect 11770 -1710 11790 -1690
rect 11770 -1760 11790 -1740
rect 11770 -1810 11790 -1790
rect 11830 -1460 11850 -1440
rect 11830 -1510 11850 -1490
rect 11830 -1560 11850 -1540
rect 11830 -1610 11850 -1590
rect 11830 -1660 11850 -1640
rect 11830 -1710 11850 -1690
rect 11830 -1760 11850 -1740
rect 11830 -1810 11850 -1790
rect 11890 -1460 11910 -1440
rect 11890 -1510 11910 -1490
rect 11890 -1560 11910 -1540
rect 11890 -1610 11910 -1590
rect 11890 -1660 11910 -1640
rect 11890 -1710 11910 -1690
rect 11890 -1760 11910 -1740
rect 11890 -1810 11910 -1790
rect 11950 -1460 11970 -1440
rect 11950 -1510 11970 -1490
rect 11950 -1560 11970 -1540
rect 11950 -1610 11970 -1590
rect 11950 -1660 11970 -1640
rect 11950 -1710 11970 -1690
rect 11950 -1760 11970 -1740
rect 11950 -1810 11970 -1790
rect 12010 -1460 12030 -1440
rect 12010 -1510 12030 -1490
rect 12010 -1560 12030 -1540
rect 12010 -1610 12030 -1590
rect 12010 -1660 12030 -1640
rect 12010 -1710 12030 -1690
rect 12010 -1760 12030 -1740
rect 12010 -1810 12030 -1790
rect 12070 -1460 12090 -1440
rect 12070 -1510 12090 -1490
rect 12070 -1560 12090 -1540
rect 12070 -1610 12090 -1590
rect 12070 -1660 12090 -1640
rect 12070 -1710 12090 -1690
rect 12070 -1760 12090 -1740
rect 12070 -1810 12090 -1790
rect 12130 -1460 12150 -1440
rect 12130 -1510 12150 -1490
rect 12130 -1560 12150 -1540
rect 12130 -1610 12150 -1590
rect 12130 -1660 12150 -1640
rect 12130 -1710 12150 -1690
rect 12130 -1760 12150 -1740
rect 12130 -1810 12150 -1790
rect 12190 -1460 12210 -1440
rect 12190 -1510 12210 -1490
rect 12190 -1560 12210 -1540
rect 12190 -1610 12210 -1590
rect 12190 -1660 12210 -1640
rect 12190 -1710 12210 -1690
rect 12190 -1760 12210 -1740
rect 12190 -1810 12210 -1790
rect 12250 -1460 12270 -1440
rect 12250 -1510 12270 -1490
rect 12250 -1560 12270 -1540
rect 12250 -1610 12270 -1590
rect 12250 -1660 12270 -1640
rect 12250 -1710 12270 -1690
rect 12250 -1760 12270 -1740
rect 12250 -1810 12270 -1790
rect 12310 -1460 12330 -1440
rect 12310 -1510 12330 -1490
rect 12310 -1560 12330 -1540
rect 12310 -1610 12330 -1590
rect 12310 -1660 12330 -1640
rect 12310 -1710 12330 -1690
rect 12310 -1760 12330 -1740
rect 12310 -1810 12330 -1790
rect 12370 -1460 12390 -1440
rect 12370 -1510 12390 -1490
rect 12370 -1560 12390 -1540
rect 12370 -1610 12390 -1590
rect 12370 -1660 12390 -1640
rect 12370 -1710 12390 -1690
rect 12370 -1760 12390 -1740
rect 12370 -1810 12390 -1790
rect 12430 -1460 12450 -1440
rect 12430 -1510 12450 -1490
rect 12430 -1560 12450 -1540
rect 12430 -1610 12450 -1590
rect 12430 -1660 12450 -1640
rect 12430 -1710 12450 -1690
rect 12430 -1760 12450 -1740
rect 12430 -1810 12450 -1790
rect 12490 -1460 12510 -1440
rect 12490 -1510 12510 -1490
rect 12490 -1560 12510 -1540
rect 12490 -1610 12510 -1590
rect 12490 -1660 12510 -1640
rect 12490 -1710 12510 -1690
rect 12490 -1760 12510 -1740
rect 12490 -1810 12510 -1790
rect 12550 -1460 12570 -1440
rect 12550 -1510 12570 -1490
rect 12550 -1560 12570 -1540
rect 12550 -1610 12570 -1590
rect 12550 -1660 12570 -1640
rect 12550 -1710 12570 -1690
rect 12550 -1760 12570 -1740
rect 12550 -1810 12570 -1790
rect 12905 -2050 12925 -2030
rect 12905 -2100 12925 -2080
rect 11230 -2140 11250 -2120
rect 11230 -2190 11250 -2170
rect 11230 -2240 11250 -2220
rect 11230 -2290 11250 -2270
rect 11230 -2340 11250 -2320
rect 11230 -2390 11250 -2370
rect 11230 -2440 11250 -2420
rect 11230 -2490 11250 -2470
rect 11290 -2140 11310 -2120
rect 11290 -2190 11310 -2170
rect 11290 -2240 11310 -2220
rect 11290 -2290 11310 -2270
rect 11290 -2340 11310 -2320
rect 11290 -2390 11310 -2370
rect 11290 -2440 11310 -2420
rect 11290 -2490 11310 -2470
rect 11350 -2140 11370 -2120
rect 11350 -2190 11370 -2170
rect 11350 -2240 11370 -2220
rect 11350 -2290 11370 -2270
rect 11350 -2340 11370 -2320
rect 11350 -2390 11370 -2370
rect 11350 -2440 11370 -2420
rect 11350 -2490 11370 -2470
rect 11410 -2140 11430 -2120
rect 11410 -2190 11430 -2170
rect 11410 -2240 11430 -2220
rect 11410 -2290 11430 -2270
rect 11410 -2340 11430 -2320
rect 11410 -2390 11430 -2370
rect 11410 -2440 11430 -2420
rect 11410 -2490 11430 -2470
rect 11470 -2140 11490 -2120
rect 11470 -2190 11490 -2170
rect 11470 -2240 11490 -2220
rect 11470 -2290 11490 -2270
rect 11470 -2340 11490 -2320
rect 11470 -2390 11490 -2370
rect 11470 -2440 11490 -2420
rect 11470 -2490 11490 -2470
rect 11530 -2140 11550 -2120
rect 11530 -2190 11550 -2170
rect 11530 -2240 11550 -2220
rect 11530 -2290 11550 -2270
rect 11530 -2340 11550 -2320
rect 11530 -2390 11550 -2370
rect 11530 -2440 11550 -2420
rect 11530 -2490 11550 -2470
rect 11590 -2140 11610 -2120
rect 11590 -2190 11610 -2170
rect 11590 -2240 11610 -2220
rect 11590 -2290 11610 -2270
rect 11590 -2340 11610 -2320
rect 11590 -2390 11610 -2370
rect 11590 -2440 11610 -2420
rect 11590 -2490 11610 -2470
rect 11650 -2140 11670 -2120
rect 11650 -2190 11670 -2170
rect 11650 -2240 11670 -2220
rect 11650 -2290 11670 -2270
rect 11650 -2340 11670 -2320
rect 11650 -2390 11670 -2370
rect 11650 -2440 11670 -2420
rect 11650 -2490 11670 -2470
rect 11710 -2140 11730 -2120
rect 11710 -2190 11730 -2170
rect 11710 -2240 11730 -2220
rect 11710 -2290 11730 -2270
rect 11710 -2340 11730 -2320
rect 11710 -2390 11730 -2370
rect 11710 -2440 11730 -2420
rect 11710 -2490 11730 -2470
rect 11770 -2140 11790 -2120
rect 11770 -2190 11790 -2170
rect 11770 -2240 11790 -2220
rect 11770 -2290 11790 -2270
rect 11770 -2340 11790 -2320
rect 11770 -2390 11790 -2370
rect 11770 -2440 11790 -2420
rect 11770 -2490 11790 -2470
rect 11830 -2140 11850 -2120
rect 11830 -2190 11850 -2170
rect 11830 -2240 11850 -2220
rect 11830 -2290 11850 -2270
rect 11830 -2340 11850 -2320
rect 11830 -2390 11850 -2370
rect 11830 -2440 11850 -2420
rect 11830 -2490 11850 -2470
rect 11890 -2140 11910 -2120
rect 11890 -2190 11910 -2170
rect 11890 -2240 11910 -2220
rect 11890 -2290 11910 -2270
rect 11890 -2340 11910 -2320
rect 11890 -2390 11910 -2370
rect 11890 -2440 11910 -2420
rect 11890 -2490 11910 -2470
rect 11950 -2140 11970 -2120
rect 11950 -2190 11970 -2170
rect 11950 -2240 11970 -2220
rect 11950 -2290 11970 -2270
rect 11950 -2340 11970 -2320
rect 11950 -2390 11970 -2370
rect 11950 -2440 11970 -2420
rect 11950 -2490 11970 -2470
rect 12010 -2140 12030 -2120
rect 12010 -2190 12030 -2170
rect 12010 -2240 12030 -2220
rect 12010 -2290 12030 -2270
rect 12010 -2340 12030 -2320
rect 12010 -2390 12030 -2370
rect 12010 -2440 12030 -2420
rect 12010 -2490 12030 -2470
rect 12070 -2140 12090 -2120
rect 12070 -2190 12090 -2170
rect 12070 -2240 12090 -2220
rect 12070 -2290 12090 -2270
rect 12070 -2340 12090 -2320
rect 12070 -2390 12090 -2370
rect 12070 -2440 12090 -2420
rect 12070 -2490 12090 -2470
rect 12130 -2140 12150 -2120
rect 12130 -2190 12150 -2170
rect 12130 -2240 12150 -2220
rect 12130 -2290 12150 -2270
rect 12130 -2340 12150 -2320
rect 12130 -2390 12150 -2370
rect 12130 -2440 12150 -2420
rect 12130 -2490 12150 -2470
rect 12190 -2140 12210 -2120
rect 12190 -2190 12210 -2170
rect 12190 -2240 12210 -2220
rect 12190 -2290 12210 -2270
rect 12190 -2340 12210 -2320
rect 12190 -2390 12210 -2370
rect 12190 -2440 12210 -2420
rect 12190 -2490 12210 -2470
rect 12250 -2140 12270 -2120
rect 12250 -2190 12270 -2170
rect 12250 -2240 12270 -2220
rect 12250 -2290 12270 -2270
rect 12250 -2340 12270 -2320
rect 12250 -2390 12270 -2370
rect 12250 -2440 12270 -2420
rect 12250 -2490 12270 -2470
rect 12310 -2140 12330 -2120
rect 12310 -2190 12330 -2170
rect 12310 -2240 12330 -2220
rect 12310 -2290 12330 -2270
rect 12310 -2340 12330 -2320
rect 12310 -2390 12330 -2370
rect 12310 -2440 12330 -2420
rect 12310 -2490 12330 -2470
rect 12370 -2140 12390 -2120
rect 12370 -2190 12390 -2170
rect 12370 -2240 12390 -2220
rect 12370 -2290 12390 -2270
rect 12370 -2340 12390 -2320
rect 12370 -2390 12390 -2370
rect 12370 -2440 12390 -2420
rect 12370 -2490 12390 -2470
rect 12430 -2140 12450 -2120
rect 12430 -2190 12450 -2170
rect 12430 -2240 12450 -2220
rect 12430 -2290 12450 -2270
rect 12430 -2340 12450 -2320
rect 12430 -2390 12450 -2370
rect 12430 -2440 12450 -2420
rect 12430 -2490 12450 -2470
rect 12490 -2140 12510 -2120
rect 12490 -2190 12510 -2170
rect 12490 -2240 12510 -2220
rect 12490 -2290 12510 -2270
rect 12490 -2340 12510 -2320
rect 12490 -2390 12510 -2370
rect 12490 -2440 12510 -2420
rect 12490 -2490 12510 -2470
rect 12550 -2140 12570 -2120
rect 12550 -2190 12570 -2170
rect 12550 -2240 12570 -2220
rect 12550 -2290 12570 -2270
rect 12905 -2150 12925 -2130
rect 12905 -2200 12925 -2180
rect 12905 -2250 12925 -2230
rect 12905 -2300 12925 -2280
rect 12960 -2050 12980 -2030
rect 12960 -2100 12980 -2080
rect 12960 -2150 12980 -2130
rect 12960 -2200 12980 -2180
rect 12960 -2250 12980 -2230
rect 12960 -2300 12980 -2280
rect 13015 -2050 13035 -2030
rect 13015 -2100 13035 -2080
rect 13015 -2150 13035 -2130
rect 13015 -2200 13035 -2180
rect 13015 -2250 13035 -2230
rect 13015 -2300 13035 -2280
rect 13070 -2050 13090 -2030
rect 13070 -2100 13090 -2080
rect 13070 -2150 13090 -2130
rect 13070 -2200 13090 -2180
rect 13070 -2250 13090 -2230
rect 13070 -2300 13090 -2280
rect 13125 -2050 13145 -2030
rect 13125 -2100 13145 -2080
rect 13125 -2150 13145 -2130
rect 13125 -2200 13145 -2180
rect 13125 -2250 13145 -2230
rect 13125 -2300 13145 -2280
rect 13180 -2050 13200 -2030
rect 13180 -2100 13200 -2080
rect 13180 -2150 13200 -2130
rect 13180 -2200 13200 -2180
rect 13180 -2250 13200 -2230
rect 13180 -2300 13200 -2280
rect 13235 -2050 13255 -2030
rect 13235 -2100 13255 -2080
rect 13235 -2150 13255 -2130
rect 13235 -2200 13255 -2180
rect 13235 -2250 13255 -2230
rect 13235 -2300 13255 -2280
rect 13290 -2050 13310 -2030
rect 13290 -2100 13310 -2080
rect 13290 -2150 13310 -2130
rect 13290 -2200 13310 -2180
rect 13290 -2250 13310 -2230
rect 13290 -2300 13310 -2280
rect 13345 -2050 13365 -2030
rect 13345 -2100 13365 -2080
rect 13345 -2150 13365 -2130
rect 13345 -2200 13365 -2180
rect 13345 -2250 13365 -2230
rect 13345 -2300 13365 -2280
rect 13400 -2050 13420 -2030
rect 13400 -2100 13420 -2080
rect 13400 -2150 13420 -2130
rect 13400 -2200 13420 -2180
rect 13400 -2250 13420 -2230
rect 13400 -2300 13420 -2280
rect 13455 -2050 13475 -2030
rect 13455 -2100 13475 -2080
rect 13455 -2150 13475 -2130
rect 13455 -2200 13475 -2180
rect 13455 -2250 13475 -2230
rect 13455 -2300 13475 -2280
rect 13510 -2050 13530 -2030
rect 13510 -2100 13530 -2080
rect 13510 -2150 13530 -2130
rect 13510 -2200 13530 -2180
rect 13510 -2250 13530 -2230
rect 13510 -2300 13530 -2280
rect 13565 -2050 13585 -2030
rect 13565 -2100 13585 -2080
rect 13565 -2150 13585 -2130
rect 13565 -2200 13585 -2180
rect 13565 -2250 13585 -2230
rect 13565 -2300 13585 -2280
rect 13620 -2050 13640 -2030
rect 13620 -2100 13640 -2080
rect 13620 -2150 13640 -2130
rect 13620 -2200 13640 -2180
rect 13620 -2250 13640 -2230
rect 13620 -2300 13640 -2280
rect 13675 -2050 13695 -2030
rect 13675 -2100 13695 -2080
rect 13675 -2150 13695 -2130
rect 13675 -2200 13695 -2180
rect 13675 -2250 13695 -2230
rect 13675 -2300 13695 -2280
rect 13730 -2050 13750 -2030
rect 13730 -2100 13750 -2080
rect 13730 -2150 13750 -2130
rect 13730 -2200 13750 -2180
rect 13730 -2250 13750 -2230
rect 13730 -2300 13750 -2280
rect 13785 -2050 13805 -2030
rect 13785 -2100 13805 -2080
rect 13785 -2150 13805 -2130
rect 13785 -2200 13805 -2180
rect 13785 -2250 13805 -2230
rect 13785 -2300 13805 -2280
rect 13840 -2050 13860 -2030
rect 13840 -2100 13860 -2080
rect 13840 -2150 13860 -2130
rect 13840 -2200 13860 -2180
rect 13840 -2250 13860 -2230
rect 13840 -2300 13860 -2280
rect 13895 -2050 13915 -2030
rect 13895 -2100 13915 -2080
rect 13895 -2150 13915 -2130
rect 13895 -2200 13915 -2180
rect 13895 -2250 13915 -2230
rect 13895 -2300 13915 -2280
rect 13950 -2050 13970 -2030
rect 13950 -2100 13970 -2080
rect 13950 -2150 13970 -2130
rect 13950 -2200 13970 -2180
rect 13950 -2250 13970 -2230
rect 13950 -2300 13970 -2280
rect 14005 -2050 14025 -2030
rect 14005 -2100 14025 -2080
rect 14005 -2150 14025 -2130
rect 14005 -2200 14025 -2180
rect 14005 -2250 14025 -2230
rect 14005 -2300 14025 -2280
rect 14060 -2050 14080 -2030
rect 14060 -2100 14080 -2080
rect 14060 -2150 14080 -2130
rect 14060 -2200 14080 -2180
rect 14060 -2250 14080 -2230
rect 14060 -2300 14080 -2280
rect 14115 -2050 14135 -2030
rect 14115 -2100 14135 -2080
rect 14115 -2150 14135 -2130
rect 14115 -2200 14135 -2180
rect 14115 -2250 14135 -2230
rect 14115 -2300 14135 -2280
rect 12550 -2340 12570 -2320
rect 12550 -2390 12570 -2370
rect 12550 -2440 12570 -2420
rect 12550 -2490 12570 -2470
rect 12905 -2480 12925 -2460
rect 12905 -2530 12925 -2510
rect 12960 -2480 12980 -2460
rect 12960 -2530 12980 -2510
rect 13015 -2480 13035 -2460
rect 13015 -2530 13035 -2510
rect 13070 -2480 13090 -2460
rect 13070 -2530 13090 -2510
rect 13125 -2480 13145 -2460
rect 13125 -2530 13145 -2510
rect 13180 -2480 13200 -2460
rect 13180 -2530 13200 -2510
rect 13235 -2480 13255 -2460
rect 13235 -2530 13255 -2510
rect 13290 -2480 13310 -2460
rect 13290 -2530 13310 -2510
rect 13345 -2480 13365 -2460
rect 13345 -2530 13365 -2510
rect 13400 -2480 13420 -2460
rect 13400 -2530 13420 -2510
rect 13455 -2480 13475 -2460
rect 13455 -2530 13475 -2510
rect 13510 -2480 13530 -2460
rect 13510 -2530 13530 -2510
rect 13565 -2480 13585 -2460
rect 13565 -2530 13585 -2510
rect 13620 -2480 13640 -2460
rect 13620 -2530 13640 -2510
rect 13675 -2480 13695 -2460
rect 13675 -2530 13695 -2510
rect 13730 -2480 13750 -2460
rect 13730 -2530 13750 -2510
rect 13785 -2480 13805 -2460
rect 13785 -2530 13805 -2510
rect 13840 -2480 13860 -2460
rect 13840 -2530 13860 -2510
rect 13895 -2480 13915 -2460
rect 13895 -2530 13915 -2510
rect 13950 -2480 13970 -2460
rect 13950 -2530 13970 -2510
rect 14005 -2480 14025 -2460
rect 14005 -2530 14025 -2510
rect 14060 -2480 14080 -2460
rect 14060 -2530 14080 -2510
rect 14115 -2480 14135 -2460
rect 14115 -2530 14135 -2510
rect 12905 -2770 12925 -2750
rect 12905 -2820 12925 -2800
rect 12905 -2870 12925 -2850
rect 11285 -2905 11305 -2885
rect 11285 -2955 11305 -2935
rect 11285 -3005 11305 -2985
rect 11340 -2905 11360 -2885
rect 11340 -2955 11360 -2935
rect 11340 -3005 11360 -2985
rect 11395 -2905 11415 -2885
rect 11395 -2955 11415 -2935
rect 11395 -3005 11415 -2985
rect 11450 -2905 11470 -2885
rect 11450 -2955 11470 -2935
rect 11450 -3005 11470 -2985
rect 11505 -2905 11525 -2885
rect 11505 -2955 11525 -2935
rect 11505 -3005 11525 -2985
rect 11560 -2905 11580 -2885
rect 11560 -2955 11580 -2935
rect 11560 -3005 11580 -2985
rect 11615 -2905 11635 -2885
rect 11615 -2955 11635 -2935
rect 11615 -3005 11635 -2985
rect 11670 -2905 11690 -2885
rect 11670 -2955 11690 -2935
rect 11670 -3005 11690 -2985
rect 11725 -2905 11745 -2885
rect 11725 -2955 11745 -2935
rect 11725 -3005 11745 -2985
rect 11780 -2905 11800 -2885
rect 11780 -2955 11800 -2935
rect 11780 -3005 11800 -2985
rect 11835 -2905 11855 -2885
rect 11835 -2955 11855 -2935
rect 11835 -3005 11855 -2985
rect 11890 -2905 11910 -2885
rect 11890 -2955 11910 -2935
rect 11890 -3005 11910 -2985
rect 11945 -2905 11965 -2885
rect 11945 -2955 11965 -2935
rect 11945 -3005 11965 -2985
rect 12000 -2905 12020 -2885
rect 12000 -2955 12020 -2935
rect 12000 -3005 12020 -2985
rect 12055 -2905 12075 -2885
rect 12055 -2955 12075 -2935
rect 12055 -3005 12075 -2985
rect 12110 -2905 12130 -2885
rect 12110 -2955 12130 -2935
rect 12110 -3005 12130 -2985
rect 12165 -2905 12185 -2885
rect 12165 -2955 12185 -2935
rect 12165 -3005 12185 -2985
rect 12220 -2905 12240 -2885
rect 12220 -2955 12240 -2935
rect 12220 -3005 12240 -2985
rect 12275 -2905 12295 -2885
rect 12275 -2955 12295 -2935
rect 12275 -3005 12295 -2985
rect 12330 -2905 12350 -2885
rect 12330 -2955 12350 -2935
rect 12330 -3005 12350 -2985
rect 12385 -2905 12405 -2885
rect 12385 -2955 12405 -2935
rect 12385 -3005 12405 -2985
rect 12440 -2905 12460 -2885
rect 12440 -2955 12460 -2935
rect 12440 -3005 12460 -2985
rect 12960 -2770 12980 -2750
rect 12960 -2820 12980 -2800
rect 12960 -2870 12980 -2850
rect 13015 -2770 13035 -2750
rect 13015 -2820 13035 -2800
rect 13015 -2870 13035 -2850
rect 13070 -2770 13090 -2750
rect 13070 -2820 13090 -2800
rect 13070 -2870 13090 -2850
rect 13125 -2770 13145 -2750
rect 13125 -2820 13145 -2800
rect 13125 -2870 13145 -2850
rect 13180 -2770 13200 -2750
rect 13180 -2820 13200 -2800
rect 13180 -2870 13200 -2850
rect 13235 -2770 13255 -2750
rect 13235 -2820 13255 -2800
rect 13235 -2870 13255 -2850
rect 13290 -2770 13310 -2750
rect 13290 -2820 13310 -2800
rect 13290 -2870 13310 -2850
rect 13345 -2770 13365 -2750
rect 13345 -2820 13365 -2800
rect 13345 -2870 13365 -2850
rect 13400 -2770 13420 -2750
rect 13400 -2820 13420 -2800
rect 13400 -2870 13420 -2850
rect 13455 -2770 13475 -2750
rect 13455 -2820 13475 -2800
rect 13455 -2870 13475 -2850
rect 13510 -2770 13530 -2750
rect 13510 -2820 13530 -2800
rect 13510 -2870 13530 -2850
rect 13565 -2770 13585 -2750
rect 13565 -2820 13585 -2800
rect 13565 -2870 13585 -2850
rect 13620 -2770 13640 -2750
rect 13620 -2820 13640 -2800
rect 13620 -2870 13640 -2850
rect 13675 -2770 13695 -2750
rect 13675 -2820 13695 -2800
rect 13675 -2870 13695 -2850
rect 13730 -2770 13750 -2750
rect 13730 -2820 13750 -2800
rect 13730 -2870 13750 -2850
rect 13785 -2770 13805 -2750
rect 13785 -2820 13805 -2800
rect 13785 -2870 13805 -2850
rect 13840 -2770 13860 -2750
rect 13840 -2820 13860 -2800
rect 13840 -2870 13860 -2850
rect 13895 -2770 13915 -2750
rect 13895 -2820 13915 -2800
rect 13895 -2870 13915 -2850
rect 13950 -2770 13970 -2750
rect 13950 -2820 13970 -2800
rect 13950 -2870 13970 -2850
rect 14005 -2770 14025 -2750
rect 14005 -2820 14025 -2800
rect 14005 -2870 14025 -2850
rect 14060 -2770 14080 -2750
rect 14060 -2820 14080 -2800
rect 14060 -2870 14080 -2850
rect 14115 -2770 14135 -2750
rect 14115 -2820 14135 -2800
rect 14115 -2870 14135 -2850
rect 12495 -2905 12515 -2885
rect 12495 -2955 12515 -2935
rect 12495 -3005 12515 -2985
rect 12905 -3050 12925 -3030
rect 12905 -3095 12925 -3075
rect 12905 -3140 12925 -3120
rect 12905 -3190 12925 -3170
rect 12905 -3235 12925 -3215
rect 12905 -3280 12925 -3260
rect 13005 -3050 13025 -3030
rect 13005 -3095 13025 -3075
rect 13005 -3140 13025 -3120
rect 13005 -3190 13025 -3170
rect 13005 -3235 13025 -3215
rect 13005 -3280 13025 -3260
rect 13105 -3050 13125 -3030
rect 13105 -3095 13125 -3075
rect 13105 -3140 13125 -3120
rect 13105 -3190 13125 -3170
rect 13105 -3235 13125 -3215
rect 13105 -3280 13125 -3260
rect 13205 -3050 13225 -3030
rect 13205 -3095 13225 -3075
rect 13205 -3140 13225 -3120
rect 13205 -3190 13225 -3170
rect 13205 -3235 13225 -3215
rect 13205 -3280 13225 -3260
rect 13305 -3050 13325 -3030
rect 13305 -3095 13325 -3075
rect 13305 -3140 13325 -3120
rect 13305 -3190 13325 -3170
rect 13305 -3235 13325 -3215
rect 13305 -3280 13325 -3260
rect 13405 -3050 13425 -3030
rect 13405 -3095 13425 -3075
rect 13405 -3140 13425 -3120
rect 13405 -3190 13425 -3170
rect 13405 -3235 13425 -3215
rect 13405 -3280 13425 -3260
rect 13505 -3050 13525 -3030
rect 13505 -3095 13525 -3075
rect 13505 -3140 13525 -3120
rect 13505 -3190 13525 -3170
rect 13505 -3235 13525 -3215
rect 13505 -3280 13525 -3260
rect 13605 -3050 13625 -3030
rect 13605 -3095 13625 -3075
rect 13605 -3140 13625 -3120
rect 13605 -3190 13625 -3170
rect 13605 -3235 13625 -3215
rect 13605 -3280 13625 -3260
rect 13705 -3050 13725 -3030
rect 13705 -3095 13725 -3075
rect 13705 -3140 13725 -3120
rect 13705 -3190 13725 -3170
rect 13705 -3235 13725 -3215
rect 13705 -3280 13725 -3260
rect 13805 -3050 13825 -3030
rect 13805 -3095 13825 -3075
rect 13805 -3140 13825 -3120
rect 13805 -3190 13825 -3170
rect 13805 -3235 13825 -3215
rect 13805 -3280 13825 -3260
rect 13905 -3050 13925 -3030
rect 13905 -3095 13925 -3075
rect 13905 -3140 13925 -3120
rect 13905 -3190 13925 -3170
rect 13905 -3235 13925 -3215
rect 13905 -3280 13925 -3260
rect 14005 -3050 14025 -3030
rect 14005 -3095 14025 -3075
rect 14005 -3140 14025 -3120
rect 14005 -3190 14025 -3170
rect 14005 -3235 14025 -3215
rect 14005 -3280 14025 -3260
rect 14105 -3050 14125 -3030
rect 14105 -3095 14125 -3075
rect 14105 -3140 14125 -3120
rect 14105 -3190 14125 -3170
rect 14105 -3235 14125 -3215
rect 14105 -3280 14125 -3260
rect 11040 -3370 11060 -3350
rect 11040 -3420 11060 -3400
rect 11040 -3470 11060 -3450
rect 11095 -3370 11115 -3350
rect 11095 -3420 11115 -3400
rect 11095 -3470 11115 -3450
rect 11150 -3370 11170 -3350
rect 11150 -3420 11170 -3400
rect 11150 -3470 11170 -3450
rect 11205 -3370 11225 -3350
rect 11205 -3420 11225 -3400
rect 11205 -3470 11225 -3450
rect 11260 -3370 11280 -3350
rect 11260 -3420 11280 -3400
rect 11260 -3470 11280 -3450
rect 11315 -3370 11335 -3350
rect 11315 -3420 11335 -3400
rect 11315 -3470 11335 -3450
rect 11370 -3370 11390 -3350
rect 11370 -3420 11390 -3400
rect 11370 -3470 11390 -3450
rect 11425 -3370 11445 -3350
rect 11425 -3420 11445 -3400
rect 11425 -3470 11445 -3450
rect 11480 -3370 11500 -3350
rect 11480 -3420 11500 -3400
rect 11480 -3470 11500 -3450
rect 11535 -3370 11555 -3350
rect 11535 -3420 11555 -3400
rect 11535 -3470 11555 -3450
rect 11590 -3370 11610 -3350
rect 11590 -3420 11610 -3400
rect 11590 -3470 11610 -3450
rect 11645 -3370 11665 -3350
rect 11645 -3420 11665 -3400
rect 11645 -3470 11665 -3450
rect 11700 -3370 11720 -3350
rect 11780 -3370 11800 -3350
rect 11700 -3420 11720 -3400
rect 11780 -3420 11800 -3400
rect 11700 -3470 11720 -3450
rect 11780 -3470 11800 -3450
rect 11835 -3370 11855 -3350
rect 11835 -3420 11855 -3400
rect 11835 -3470 11855 -3450
rect 11890 -3370 11910 -3350
rect 11890 -3420 11910 -3400
rect 11890 -3470 11910 -3450
rect 11945 -3370 11965 -3350
rect 11945 -3420 11965 -3400
rect 11945 -3470 11965 -3450
rect 12000 -3370 12020 -3350
rect 12080 -3370 12100 -3350
rect 12000 -3420 12020 -3400
rect 12080 -3420 12100 -3400
rect 12000 -3470 12020 -3450
rect 12080 -3470 12100 -3450
rect 12135 -3370 12155 -3350
rect 12135 -3420 12155 -3400
rect 12135 -3470 12155 -3450
rect 12190 -3370 12210 -3350
rect 12190 -3420 12210 -3400
rect 12190 -3470 12210 -3450
rect 12245 -3370 12265 -3350
rect 12245 -3420 12265 -3400
rect 12245 -3470 12265 -3450
rect 12300 -3370 12320 -3350
rect 12300 -3420 12320 -3400
rect 12300 -3470 12320 -3450
rect 12355 -3370 12375 -3350
rect 12355 -3420 12375 -3400
rect 12355 -3470 12375 -3450
rect 12410 -3370 12430 -3350
rect 12410 -3420 12430 -3400
rect 12410 -3470 12430 -3450
rect 12465 -3370 12485 -3350
rect 12465 -3420 12485 -3400
rect 12465 -3470 12485 -3450
rect 12520 -3370 12540 -3350
rect 12520 -3420 12540 -3400
rect 12520 -3470 12540 -3450
rect 12575 -3370 12595 -3350
rect 12575 -3420 12595 -3400
rect 12575 -3470 12595 -3450
rect 12630 -3370 12650 -3350
rect 12630 -3420 12650 -3400
rect 12630 -3470 12650 -3450
rect 12685 -3370 12705 -3350
rect 12685 -3420 12705 -3400
rect 12685 -3470 12705 -3450
rect 12740 -3370 12760 -3350
rect 12740 -3420 12760 -3400
rect 12740 -3470 12760 -3450
rect 11215 -3850 11235 -3830
rect 11215 -3900 11235 -3880
rect 11215 -3950 11235 -3930
rect 11215 -4000 11235 -3980
rect 11215 -4050 11235 -4030
rect 11270 -3850 11290 -3830
rect 11270 -3900 11290 -3880
rect 11270 -3950 11290 -3930
rect 11270 -4000 11290 -3980
rect 11270 -4050 11290 -4030
rect 11325 -3850 11345 -3830
rect 11325 -3900 11345 -3880
rect 11325 -3950 11345 -3930
rect 11325 -4000 11345 -3980
rect 11325 -4050 11345 -4030
rect 11380 -3850 11400 -3830
rect 11380 -3900 11400 -3880
rect 11380 -3950 11400 -3930
rect 11380 -4000 11400 -3980
rect 11380 -4050 11400 -4030
rect 11435 -3850 11455 -3830
rect 11435 -3900 11455 -3880
rect 11435 -3950 11455 -3930
rect 11435 -4000 11455 -3980
rect 11435 -4050 11455 -4030
rect 11490 -3850 11510 -3830
rect 11490 -3900 11510 -3880
rect 11490 -3950 11510 -3930
rect 11490 -4000 11510 -3980
rect 11490 -4050 11510 -4030
rect 11545 -3850 11565 -3830
rect 11545 -3900 11565 -3880
rect 11545 -3950 11565 -3930
rect 11545 -4000 11565 -3980
rect 11545 -4050 11565 -4030
rect 11600 -3850 11620 -3830
rect 11600 -3900 11620 -3880
rect 11600 -3950 11620 -3930
rect 11600 -4000 11620 -3980
rect 11600 -4050 11620 -4030
rect 11655 -3850 11675 -3830
rect 11655 -3900 11675 -3880
rect 11655 -3950 11675 -3930
rect 11655 -4000 11675 -3980
rect 11655 -4050 11675 -4030
rect 11710 -3850 11730 -3830
rect 11710 -3900 11730 -3880
rect 11710 -3950 11730 -3930
rect 11710 -4000 11730 -3980
rect 11710 -4050 11730 -4030
rect 11765 -3850 11785 -3830
rect 11765 -3900 11785 -3880
rect 11765 -3950 11785 -3930
rect 11765 -4000 11785 -3980
rect 11765 -4050 11785 -4030
rect 11820 -3850 11840 -3830
rect 11820 -3900 11840 -3880
rect 11820 -3950 11840 -3930
rect 11820 -4000 11840 -3980
rect 11820 -4050 11840 -4030
rect 11875 -3850 11895 -3830
rect 11875 -3900 11895 -3880
rect 11875 -3950 11895 -3930
rect 11875 -4000 11895 -3980
rect 11875 -4050 11895 -4030
rect 11930 -3850 11950 -3830
rect 11930 -3900 11950 -3880
rect 11930 -3950 11950 -3930
rect 11930 -4000 11950 -3980
rect 11930 -4050 11950 -4030
rect 11985 -3850 12005 -3830
rect 11985 -3900 12005 -3880
rect 11985 -3950 12005 -3930
rect 11985 -4000 12005 -3980
rect 11985 -4050 12005 -4030
rect 12040 -3850 12060 -3830
rect 12040 -3900 12060 -3880
rect 12040 -3950 12060 -3930
rect 12040 -4000 12060 -3980
rect 12040 -4050 12060 -4030
rect 12095 -3850 12115 -3830
rect 12095 -3900 12115 -3880
rect 12095 -3950 12115 -3930
rect 12095 -4000 12115 -3980
rect 12095 -4050 12115 -4030
rect 12150 -3850 12170 -3830
rect 12150 -3900 12170 -3880
rect 12150 -3950 12170 -3930
rect 12150 -4000 12170 -3980
rect 12150 -4050 12170 -4030
rect 12205 -3850 12225 -3830
rect 12205 -3900 12225 -3880
rect 12205 -3950 12225 -3930
rect 12205 -4000 12225 -3980
rect 12205 -4050 12225 -4030
rect 12260 -3850 12280 -3830
rect 12260 -3900 12280 -3880
rect 12260 -3950 12280 -3930
rect 12260 -4000 12280 -3980
rect 12260 -4050 12280 -4030
rect 12315 -3850 12335 -3830
rect 12315 -3900 12335 -3880
rect 12315 -3950 12335 -3930
rect 12315 -4000 12335 -3980
rect 12315 -4050 12335 -4030
rect 12370 -3850 12390 -3830
rect 12370 -3900 12390 -3880
rect 12370 -3950 12390 -3930
rect 12370 -4000 12390 -3980
rect 12370 -4050 12390 -4030
rect 12425 -3850 12445 -3830
rect 12425 -3900 12445 -3880
rect 12425 -3950 12445 -3930
rect 12425 -4000 12445 -3980
rect 12425 -4050 12445 -4030
rect 12480 -3850 12500 -3830
rect 12480 -3900 12500 -3880
rect 12480 -3950 12500 -3930
rect 12480 -4000 12500 -3980
rect 12480 -4050 12500 -4030
rect 12535 -3850 12555 -3830
rect 12535 -3900 12555 -3880
rect 12535 -3950 12555 -3930
rect 12535 -4000 12555 -3980
rect 12535 -4050 12555 -4030
rect 12590 -3850 12610 -3830
rect 12590 -3900 12610 -3880
rect 12590 -3950 12610 -3930
rect 12590 -4000 12610 -3980
rect 12590 -4050 12610 -4030
<< pdiffc >>
rect 3005 2895 3025 2915
rect 3005 2845 3025 2865
rect 3095 2895 3115 2915
rect 3095 2845 3115 2865
rect 3185 2895 3205 2915
rect 3185 2845 3205 2865
rect 3275 2895 3295 2915
rect 3275 2845 3295 2865
rect 3365 2895 3385 2915
rect 3365 2845 3385 2865
rect 3455 2895 3475 2915
rect 3455 2845 3475 2865
rect 3545 2895 3565 2915
rect 3545 2845 3565 2865
rect 3635 2895 3655 2915
rect 3635 2845 3655 2865
rect 3725 2895 3745 2915
rect 3725 2845 3745 2865
rect 3815 2895 3835 2915
rect 3815 2845 3835 2865
rect 3905 2895 3925 2915
rect 3905 2845 3925 2865
rect 3995 2895 4015 2915
rect 3995 2845 4015 2865
rect 4085 2895 4105 2915
rect 4085 2845 4105 2865
rect 4175 2895 4195 2915
rect 4175 2845 4195 2865
rect 4265 2895 4285 2915
rect 4265 2845 4285 2865
rect 4355 2895 4375 2915
rect 4355 2845 4375 2865
rect 4445 2895 4465 2915
rect 4445 2845 4465 2865
rect 4535 2895 4555 2915
rect 4535 2845 4555 2865
rect 4625 2895 4645 2915
rect 4625 2845 4645 2865
rect 4715 2895 4735 2915
rect 4715 2845 4735 2865
rect 4805 2895 4825 2915
rect 4805 2845 4825 2865
rect 4895 2895 4915 2915
rect 4895 2845 4915 2865
rect 4985 2895 5005 2915
rect 4985 2845 5005 2865
rect 3185 2665 3205 2685
rect 3185 2615 3205 2635
rect 3185 2565 3205 2585
rect 3185 2515 3205 2535
rect 3185 2465 3205 2485
rect 3185 2415 3205 2435
rect 3275 2665 3295 2685
rect 3275 2615 3295 2635
rect 3275 2565 3295 2585
rect 3275 2515 3295 2535
rect 3275 2465 3295 2485
rect 3275 2415 3295 2435
rect 3365 2665 3385 2685
rect 3365 2615 3385 2635
rect 3365 2565 3385 2585
rect 3365 2515 3385 2535
rect 3365 2465 3385 2485
rect 3365 2415 3385 2435
rect 3455 2665 3475 2685
rect 3455 2615 3475 2635
rect 3455 2565 3475 2585
rect 3455 2515 3475 2535
rect 3455 2465 3475 2485
rect 3455 2415 3475 2435
rect 3545 2665 3565 2685
rect 3545 2615 3565 2635
rect 3545 2565 3565 2585
rect 3545 2515 3565 2535
rect 3545 2465 3565 2485
rect 3545 2415 3565 2435
rect 3635 2665 3655 2685
rect 3635 2615 3655 2635
rect 3635 2565 3655 2585
rect 3635 2515 3655 2535
rect 3635 2465 3655 2485
rect 3635 2415 3655 2435
rect 3725 2665 3745 2685
rect 3725 2615 3745 2635
rect 3725 2565 3745 2585
rect 3725 2515 3745 2535
rect 3725 2465 3745 2485
rect 3725 2415 3745 2435
rect 3815 2665 3835 2685
rect 3815 2615 3835 2635
rect 3815 2565 3835 2585
rect 3815 2515 3835 2535
rect 3815 2465 3835 2485
rect 3815 2415 3835 2435
rect 3905 2665 3925 2685
rect 3905 2615 3925 2635
rect 3905 2565 3925 2585
rect 3905 2515 3925 2535
rect 3905 2465 3925 2485
rect 3905 2415 3925 2435
rect 3995 2665 4015 2685
rect 3995 2615 4015 2635
rect 3995 2565 4015 2585
rect 3995 2515 4015 2535
rect 3995 2465 4015 2485
rect 3995 2415 4015 2435
rect 4085 2665 4105 2685
rect 4085 2615 4105 2635
rect 4085 2565 4105 2585
rect 4085 2515 4105 2535
rect 4085 2465 4105 2485
rect 4085 2415 4105 2435
rect 4175 2665 4195 2685
rect 4175 2615 4195 2635
rect 4175 2565 4195 2585
rect 4175 2515 4195 2535
rect 4175 2465 4195 2485
rect 4175 2415 4195 2435
rect 4265 2665 4285 2685
rect 4265 2615 4285 2635
rect 4265 2565 4285 2585
rect 4265 2515 4285 2535
rect 4265 2465 4285 2485
rect 4265 2415 4285 2435
rect 4355 2665 4375 2685
rect 4355 2615 4375 2635
rect 4355 2565 4375 2585
rect 4355 2515 4375 2535
rect 4355 2465 4375 2485
rect 4355 2415 4375 2435
rect 4445 2665 4465 2685
rect 4445 2615 4465 2635
rect 4445 2565 4465 2585
rect 4445 2515 4465 2535
rect 4445 2465 4465 2485
rect 4445 2415 4465 2435
rect 4535 2665 4555 2685
rect 4535 2615 4555 2635
rect 4535 2565 4555 2585
rect 4535 2515 4555 2535
rect 4535 2465 4555 2485
rect 4535 2415 4555 2435
rect 4625 2665 4645 2685
rect 4625 2615 4645 2635
rect 4625 2565 4645 2585
rect 4625 2515 4645 2535
rect 4625 2465 4645 2485
rect 4625 2415 4645 2435
rect 4715 2665 4735 2685
rect 4715 2615 4735 2635
rect 4715 2565 4735 2585
rect 4715 2515 4735 2535
rect 4715 2465 4735 2485
rect 4715 2415 4735 2435
rect 4805 2665 4825 2685
rect 4805 2615 4825 2635
rect 4805 2565 4825 2585
rect 4805 2515 4825 2535
rect 4805 2465 4825 2485
rect 4805 2415 4825 2435
rect 2575 1965 2595 1985
rect 2575 1915 2595 1935
rect 2630 1965 2650 1985
rect 2630 1915 2650 1935
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2755 1965 2775 1985
rect 2755 1915 2775 1935
rect 2815 1965 2835 1985
rect 2815 1915 2835 1935
rect 2875 1965 2895 1985
rect 2875 1915 2895 1935
rect 2935 1965 2955 1985
rect 2935 1915 2955 1935
rect 2995 1965 3015 1985
rect 2995 1915 3015 1935
rect 3055 1965 3075 1985
rect 3055 1915 3075 1935
rect 3115 1965 3135 1985
rect 3115 1915 3135 1935
rect 3175 1965 3195 1985
rect 3175 1915 3195 1935
rect 3235 1965 3255 1985
rect 3235 1915 3255 1935
rect 3295 1965 3315 1985
rect 3295 1915 3315 1935
rect 3355 1965 3375 1985
rect 3355 1915 3375 1935
rect 3415 1965 3435 1985
rect 3415 1915 3435 1935
rect 3475 1965 3495 1985
rect 3475 1915 3495 1935
rect 3535 1965 3555 1985
rect 3535 1915 3555 1935
rect 3595 1965 3615 1985
rect 3595 1915 3615 1935
rect 3655 1965 3675 1985
rect 3655 1915 3675 1935
rect 3715 1965 3735 1985
rect 3715 1915 3735 1935
rect 3775 1965 3795 1985
rect 3775 1915 3795 1935
rect 3835 1965 3855 1985
rect 3835 1915 3855 1935
rect 3895 1965 3915 1985
rect 3895 1915 3915 1935
rect 3955 1965 3975 1985
rect 4035 1965 4055 1985
rect 3955 1915 3975 1935
rect 4035 1915 4055 1935
rect 4095 1965 4115 1985
rect 4095 1915 4115 1935
rect 4155 1965 4175 1985
rect 4155 1915 4175 1935
rect 4215 1965 4235 1985
rect 4215 1915 4235 1935
rect 4275 1965 4295 1985
rect 4275 1915 4295 1935
rect 4335 1965 4355 1985
rect 4335 1915 4355 1935
rect 4395 1965 4415 1985
rect 4395 1915 4415 1935
rect 4455 1965 4475 1985
rect 4455 1915 4475 1935
rect 4515 1965 4535 1985
rect 4515 1915 4535 1935
rect 4575 1965 4595 1985
rect 4575 1915 4595 1935
rect 4635 1965 4655 1985
rect 4635 1915 4655 1935
rect 4695 1965 4715 1985
rect 4695 1915 4715 1935
rect 4755 1965 4775 1985
rect 4755 1915 4775 1935
rect 4815 1965 4835 1985
rect 4815 1915 4835 1935
rect 4875 1965 4895 1985
rect 4875 1915 4895 1935
rect 4935 1965 4955 1985
rect 4935 1915 4955 1935
rect 4995 1965 5015 1985
rect 4995 1915 5015 1935
rect 5055 1965 5075 1985
rect 5055 1915 5075 1935
rect 5115 1965 5135 1985
rect 5115 1915 5135 1935
rect 5175 1965 5195 1985
rect 5175 1915 5195 1935
rect 5235 1965 5255 1985
rect 5235 1915 5255 1935
<< psubdiff >>
rect 11200 8915 11240 8943
rect 11200 8895 11210 8915
rect 11230 8895 11240 8915
rect 11200 8880 11240 8895
rect 11460 8915 11500 8943
rect 11460 8895 11470 8915
rect 11490 8895 11500 8915
rect 11460 8880 11500 8895
rect 11530 8930 11570 8960
rect 11530 8910 11540 8930
rect 11560 8910 11570 8930
rect 11530 8880 11570 8910
rect 11970 8930 12010 8960
rect 11970 8910 11980 8930
rect 12000 8910 12010 8930
rect 11970 8880 12010 8910
rect 12040 8915 12080 8935
rect 12040 8895 12050 8915
rect 12070 8895 12080 8915
rect 12040 8875 12080 8895
rect 12600 8915 12640 8935
rect 12600 8895 12610 8915
rect 12630 8895 12640 8915
rect 12600 8875 12640 8895
rect 10780 8515 10820 8550
rect 10780 8495 10790 8515
rect 10810 8495 10820 8515
rect 10780 8465 10820 8495
rect 10780 8445 10790 8465
rect 10810 8445 10820 8465
rect 10780 8415 10820 8445
rect 10780 8395 10790 8415
rect 10810 8395 10820 8415
rect 10780 8365 10820 8395
rect 10780 8345 10790 8365
rect 10810 8345 10820 8365
rect 10780 8315 10820 8345
rect 10780 8295 10790 8315
rect 10810 8295 10820 8315
rect 10450 8265 10490 8293
rect 10450 8245 10460 8265
rect 10480 8245 10490 8265
rect 10450 8230 10490 8245
rect 10710 8265 10750 8293
rect 10710 8245 10720 8265
rect 10740 8245 10750 8265
rect 10710 8230 10750 8245
rect 10780 8265 10820 8295
rect 10780 8245 10790 8265
rect 10810 8245 10820 8265
rect 10780 8230 10820 8245
rect 11100 8565 11140 8580
rect 11100 8545 11110 8565
rect 11130 8545 11140 8565
rect 11100 8515 11140 8545
rect 11100 8495 11110 8515
rect 11130 8495 11140 8515
rect 11100 8465 11140 8495
rect 11100 8445 11110 8465
rect 11130 8445 11140 8465
rect 11100 8415 11140 8445
rect 11100 8395 11110 8415
rect 11130 8395 11140 8415
rect 11100 8365 11140 8395
rect 11100 8345 11110 8365
rect 11130 8345 11140 8365
rect 11100 8315 11140 8345
rect 11100 8295 11110 8315
rect 11130 8295 11140 8315
rect 11100 8265 11140 8295
rect 11100 8245 11110 8265
rect 11130 8245 11140 8265
rect 11100 8230 11140 8245
rect 11180 8560 11220 8575
rect 11180 8540 11190 8560
rect 11210 8540 11220 8560
rect 11180 8510 11220 8540
rect 11180 8490 11190 8510
rect 11210 8490 11220 8510
rect 11180 8460 11220 8490
rect 11180 8440 11190 8460
rect 11210 8440 11220 8460
rect 11180 8410 11220 8440
rect 11180 8390 11190 8410
rect 11210 8390 11220 8410
rect 11180 8360 11220 8390
rect 11180 8340 11190 8360
rect 11210 8340 11220 8360
rect 11180 8310 11220 8340
rect 11180 8290 11190 8310
rect 11210 8290 11220 8310
rect 11180 8260 11220 8290
rect 11180 8240 11190 8260
rect 11210 8240 11220 8260
rect 11180 8210 11220 8240
rect 11180 8190 11190 8210
rect 11210 8190 11220 8210
rect 11180 8175 11220 8190
rect 12580 8560 12620 8575
rect 12580 8540 12590 8560
rect 12610 8540 12620 8560
rect 12580 8510 12620 8540
rect 12580 8490 12590 8510
rect 12610 8490 12620 8510
rect 12580 8460 12620 8490
rect 12580 8440 12590 8460
rect 12610 8440 12620 8460
rect 12580 8410 12620 8440
rect 12580 8390 12590 8410
rect 12610 8390 12620 8410
rect 12580 8360 12620 8390
rect 12580 8340 12590 8360
rect 12610 8340 12620 8360
rect 18280 8515 18320 8550
rect 18280 8495 18290 8515
rect 18310 8495 18320 8515
rect 18280 8465 18320 8495
rect 18280 8445 18290 8465
rect 18310 8445 18320 8465
rect 18280 8415 18320 8445
rect 18280 8395 18290 8415
rect 18310 8395 18320 8415
rect 18280 8365 18320 8395
rect 12580 8310 12620 8340
rect 12580 8290 12590 8310
rect 12610 8290 12620 8310
rect 18280 8345 18290 8365
rect 18310 8345 18320 8365
rect 18280 8315 18320 8345
rect 18280 8295 18290 8315
rect 18310 8295 18320 8315
rect 12580 8260 12620 8290
rect 12580 8240 12590 8260
rect 12610 8240 12620 8260
rect 17950 8265 17990 8293
rect 17950 8245 17960 8265
rect 17980 8245 17990 8265
rect 12580 8210 12620 8240
rect 12580 8190 12590 8210
rect 12610 8190 12620 8210
rect 12580 8175 12620 8190
rect 12855 8225 12895 8240
rect 12855 8205 12865 8225
rect 12885 8205 12895 8225
rect 12855 8175 12895 8205
rect 12855 8155 12865 8175
rect 12885 8155 12895 8175
rect 12855 8125 12895 8155
rect 12855 8105 12865 8125
rect 12885 8105 12895 8125
rect 12855 8075 12895 8105
rect 12855 8055 12865 8075
rect 12885 8055 12895 8075
rect 12855 8025 12895 8055
rect 12855 8005 12865 8025
rect 12885 8005 12895 8025
rect 12855 7975 12895 8005
rect 12855 7955 12865 7975
rect 12885 7955 12895 7975
rect 12855 7940 12895 7955
rect 14145 8225 14185 8240
rect 17950 8230 17990 8245
rect 18210 8265 18250 8293
rect 18210 8245 18220 8265
rect 18240 8245 18250 8265
rect 18210 8230 18250 8245
rect 18280 8265 18320 8295
rect 18280 8245 18290 8265
rect 18310 8245 18320 8265
rect 18280 8230 18320 8245
rect 18600 8565 18640 8580
rect 18600 8545 18610 8565
rect 18630 8545 18640 8565
rect 18600 8515 18640 8545
rect 18600 8495 18610 8515
rect 18630 8495 18640 8515
rect 18600 8465 18640 8495
rect 18600 8445 18610 8465
rect 18630 8445 18640 8465
rect 18600 8415 18640 8445
rect 18600 8395 18610 8415
rect 18630 8395 18640 8415
rect 18600 8365 18640 8395
rect 18600 8345 18610 8365
rect 18630 8345 18640 8365
rect 18600 8315 18640 8345
rect 18600 8295 18610 8315
rect 18630 8295 18640 8315
rect 18600 8265 18640 8295
rect 18600 8245 18610 8265
rect 18630 8245 18640 8265
rect 18600 8230 18640 8245
rect 18680 8560 18720 8575
rect 18680 8540 18690 8560
rect 18710 8540 18720 8560
rect 18680 8510 18720 8540
rect 18680 8490 18690 8510
rect 18710 8490 18720 8510
rect 18680 8460 18720 8490
rect 18680 8440 18690 8460
rect 18710 8440 18720 8460
rect 18680 8410 18720 8440
rect 18680 8390 18690 8410
rect 18710 8390 18720 8410
rect 18680 8360 18720 8390
rect 18680 8340 18690 8360
rect 18710 8340 18720 8360
rect 18680 8310 18720 8340
rect 18680 8290 18690 8310
rect 18710 8290 18720 8310
rect 18680 8260 18720 8290
rect 18680 8240 18690 8260
rect 18710 8240 18720 8260
rect 14145 8205 14155 8225
rect 14175 8205 14185 8225
rect 14145 8175 14185 8205
rect 18680 8210 18720 8240
rect 18680 8190 18690 8210
rect 18710 8190 18720 8210
rect 18680 8175 18720 8190
rect 20080 8560 20120 8575
rect 20080 8540 20090 8560
rect 20110 8540 20120 8560
rect 20080 8510 20120 8540
rect 20080 8490 20090 8510
rect 20110 8490 20120 8510
rect 20080 8460 20120 8490
rect 20080 8440 20090 8460
rect 20110 8440 20120 8460
rect 20080 8410 20120 8440
rect 20080 8390 20090 8410
rect 20110 8390 20120 8410
rect 20080 8360 20120 8390
rect 20080 8340 20090 8360
rect 20110 8340 20120 8360
rect 20080 8310 20120 8340
rect 20080 8290 20090 8310
rect 20110 8290 20120 8310
rect 20080 8260 20120 8290
rect 20080 8240 20090 8260
rect 20110 8240 20120 8260
rect 20080 8210 20120 8240
rect 20080 8190 20090 8210
rect 20110 8190 20120 8210
rect 20080 8175 20120 8190
rect 20350 8225 20390 8240
rect 20350 8205 20360 8225
rect 20380 8205 20390 8225
rect 20350 8175 20390 8205
rect 14145 8155 14155 8175
rect 14175 8155 14185 8175
rect 14145 8125 14185 8155
rect 20350 8155 20360 8175
rect 20380 8155 20390 8175
rect 14145 8105 14155 8125
rect 14175 8105 14185 8125
rect 20350 8125 20390 8155
rect 14145 8075 14185 8105
rect 14145 8055 14155 8075
rect 14175 8055 14185 8075
rect 14145 8025 14185 8055
rect 14145 8005 14155 8025
rect 14175 8005 14185 8025
rect 14145 7975 14185 8005
rect 14145 7955 14155 7975
rect 14175 7955 14185 7975
rect 14145 7940 14185 7955
rect 20350 8105 20360 8125
rect 20380 8105 20390 8125
rect 20350 8075 20390 8105
rect 20350 8055 20360 8075
rect 20380 8055 20390 8075
rect 20350 8025 20390 8055
rect 20350 8005 20360 8025
rect 20380 8005 20390 8025
rect 20350 7975 20390 8005
rect 20350 7955 20360 7975
rect 20380 7955 20390 7975
rect 11180 7880 11220 7895
rect 11180 7860 11190 7880
rect 11210 7860 11220 7880
rect 11180 7830 11220 7860
rect 11180 7810 11190 7830
rect 11210 7810 11220 7830
rect 11180 7780 11220 7810
rect 11180 7760 11190 7780
rect 11210 7760 11220 7780
rect 11180 7730 11220 7760
rect 11180 7710 11190 7730
rect 11210 7710 11220 7730
rect 11180 7680 11220 7710
rect 11180 7660 11190 7680
rect 11210 7660 11220 7680
rect 11180 7630 11220 7660
rect 9640 7605 9680 7620
rect 9640 7585 9650 7605
rect 9670 7585 9680 7605
rect 9640 7555 9680 7585
rect 9640 7535 9650 7555
rect 9670 7535 9680 7555
rect 9640 7520 9680 7535
rect 10930 7605 10970 7620
rect 10930 7585 10940 7605
rect 10960 7585 10970 7605
rect 10930 7555 10970 7585
rect 10930 7535 10940 7555
rect 10960 7535 10970 7555
rect 10930 7520 10970 7535
rect 11180 7610 11190 7630
rect 11210 7610 11220 7630
rect 11180 7580 11220 7610
rect 11180 7560 11190 7580
rect 11210 7560 11220 7580
rect 11180 7530 11220 7560
rect 11180 7510 11190 7530
rect 11210 7510 11220 7530
rect 11180 7495 11220 7510
rect 12580 7880 12620 7895
rect 20350 7940 20390 7955
rect 21640 8225 21680 8240
rect 21640 8205 21650 8225
rect 21670 8205 21680 8225
rect 21640 8175 21680 8205
rect 21640 8155 21650 8175
rect 21670 8155 21680 8175
rect 21640 8125 21680 8155
rect 21640 8105 21650 8125
rect 21670 8105 21680 8125
rect 21640 8075 21680 8105
rect 21640 8055 21650 8075
rect 21670 8055 21680 8075
rect 21640 8025 21680 8055
rect 21640 8005 21650 8025
rect 21670 8005 21680 8025
rect 21640 7975 21680 8005
rect 21640 7955 21650 7975
rect 21670 7955 21680 7975
rect 21640 7940 21680 7955
rect 12580 7860 12590 7880
rect 12610 7860 12620 7880
rect 12580 7830 12620 7860
rect 18680 7880 18720 7895
rect 18680 7860 18690 7880
rect 18710 7860 18720 7880
rect 12580 7810 12590 7830
rect 12610 7810 12620 7830
rect 12580 7780 12620 7810
rect 12580 7760 12590 7780
rect 12610 7760 12620 7780
rect 12580 7730 12620 7760
rect 12580 7710 12590 7730
rect 12610 7710 12620 7730
rect 12580 7680 12620 7710
rect 18680 7830 18720 7860
rect 18680 7810 18690 7830
rect 18710 7810 18720 7830
rect 18680 7780 18720 7810
rect 18680 7760 18690 7780
rect 18710 7760 18720 7780
rect 18680 7730 18720 7760
rect 18680 7710 18690 7730
rect 18710 7710 18720 7730
rect 12580 7660 12590 7680
rect 12610 7660 12620 7680
rect 12580 7630 12620 7660
rect 18680 7680 18720 7710
rect 18680 7660 18690 7680
rect 18710 7660 18720 7680
rect 12580 7610 12590 7630
rect 12610 7610 12620 7630
rect 18680 7630 18720 7660
rect 12580 7580 12620 7610
rect 12580 7560 12590 7580
rect 12610 7560 12620 7580
rect 12580 7530 12620 7560
rect 12580 7510 12590 7530
rect 12610 7510 12620 7530
rect 12855 7605 12895 7620
rect 12855 7585 12865 7605
rect 12885 7585 12895 7605
rect 12855 7555 12895 7585
rect 12855 7535 12865 7555
rect 12885 7535 12895 7555
rect 12855 7520 12895 7535
rect 14145 7605 14185 7620
rect 14145 7585 14155 7605
rect 14175 7585 14185 7605
rect 14145 7555 14185 7585
rect 14145 7535 14155 7555
rect 14175 7535 14185 7555
rect 14145 7520 14185 7535
rect 17140 7605 17180 7620
rect 17140 7585 17150 7605
rect 17170 7585 17180 7605
rect 17140 7555 17180 7585
rect 17140 7535 17150 7555
rect 17170 7535 17180 7555
rect 17140 7520 17180 7535
rect 18430 7605 18470 7620
rect 18430 7585 18440 7605
rect 18460 7585 18470 7605
rect 18430 7555 18470 7585
rect 18430 7535 18440 7555
rect 18460 7535 18470 7555
rect 18430 7520 18470 7535
rect 18680 7610 18690 7630
rect 18710 7610 18720 7630
rect 18680 7580 18720 7610
rect 18680 7560 18690 7580
rect 18710 7560 18720 7580
rect 18680 7530 18720 7560
rect 12580 7495 12620 7510
rect 18680 7510 18690 7530
rect 18710 7510 18720 7530
rect 18680 7495 18720 7510
rect 20080 7880 20120 7895
rect 20080 7860 20090 7880
rect 20110 7860 20120 7880
rect 20080 7830 20120 7860
rect 20080 7810 20090 7830
rect 20110 7810 20120 7830
rect 20080 7780 20120 7810
rect 20080 7760 20090 7780
rect 20110 7760 20120 7780
rect 20080 7730 20120 7760
rect 20080 7710 20090 7730
rect 20110 7710 20120 7730
rect 20080 7680 20120 7710
rect 20080 7660 20090 7680
rect 20110 7660 20120 7680
rect 20080 7630 20120 7660
rect 20080 7610 20090 7630
rect 20110 7610 20120 7630
rect 20080 7580 20120 7610
rect 20080 7560 20090 7580
rect 20110 7560 20120 7580
rect 20080 7530 20120 7560
rect 20080 7510 20090 7530
rect 20110 7510 20120 7530
rect 20350 7605 20390 7620
rect 20350 7585 20360 7605
rect 20380 7585 20390 7605
rect 20350 7555 20390 7585
rect 20350 7535 20360 7555
rect 20380 7535 20390 7555
rect 20350 7520 20390 7535
rect 21640 7605 21680 7620
rect 21640 7585 21650 7605
rect 21670 7585 21680 7605
rect 21640 7555 21680 7585
rect 21640 7535 21650 7555
rect 21670 7535 21680 7555
rect 21640 7520 21680 7535
rect 20080 7495 20120 7510
rect 9640 7155 9680 7170
rect 9640 7135 9650 7155
rect 9670 7135 9680 7155
rect 9640 7105 9680 7135
rect 9640 7085 9650 7105
rect 9670 7085 9680 7105
rect 9640 7055 9680 7085
rect 9640 7035 9650 7055
rect 9670 7035 9680 7055
rect 9640 7020 9680 7035
rect 10930 7155 10970 7170
rect 12855 7155 12895 7170
rect 10930 7135 10940 7155
rect 10960 7135 10970 7155
rect 10930 7105 10970 7135
rect 12855 7135 12865 7155
rect 12885 7135 12895 7155
rect 10930 7085 10940 7105
rect 10960 7085 10970 7105
rect 10930 7055 10970 7085
rect 10930 7035 10940 7055
rect 10960 7035 10970 7055
rect 10930 7020 10970 7035
rect 11235 7115 11275 7130
rect 11235 7095 11245 7115
rect 11265 7095 11275 7115
rect 11235 7065 11275 7095
rect 11235 7045 11245 7065
rect 11265 7045 11275 7065
rect 11235 7015 11275 7045
rect 11235 6995 11245 7015
rect 11265 6995 11275 7015
rect 11235 6980 11275 6995
rect 12525 7115 12565 7130
rect 12525 7095 12535 7115
rect 12555 7095 12565 7115
rect 12525 7065 12565 7095
rect 12525 7045 12535 7065
rect 12555 7045 12565 7065
rect 12525 7015 12565 7045
rect 12855 7105 12895 7135
rect 12855 7085 12865 7105
rect 12885 7085 12895 7105
rect 12855 7055 12895 7085
rect 12855 7035 12865 7055
rect 12885 7035 12895 7055
rect 12855 7020 12895 7035
rect 14145 7155 14185 7170
rect 14145 7135 14155 7155
rect 14175 7135 14185 7155
rect 14145 7105 14185 7135
rect 14145 7085 14155 7105
rect 14175 7085 14185 7105
rect 14145 7055 14185 7085
rect 14145 7035 14155 7055
rect 14175 7035 14185 7055
rect 14145 7020 14185 7035
rect 17140 7155 17180 7170
rect 17140 7135 17150 7155
rect 17170 7135 17180 7155
rect 17140 7105 17180 7135
rect 17140 7085 17150 7105
rect 17170 7085 17180 7105
rect 17140 7055 17180 7085
rect 17140 7035 17150 7055
rect 17170 7035 17180 7055
rect 17140 7020 17180 7035
rect 18430 7155 18470 7170
rect 20350 7155 20390 7170
rect 18430 7135 18440 7155
rect 18460 7135 18470 7155
rect 18430 7105 18470 7135
rect 20350 7135 20360 7155
rect 20380 7135 20390 7155
rect 18430 7085 18440 7105
rect 18460 7085 18470 7105
rect 18430 7055 18470 7085
rect 18430 7035 18440 7055
rect 18460 7035 18470 7055
rect 18430 7020 18470 7035
rect 18735 7115 18775 7130
rect 18735 7095 18745 7115
rect 18765 7095 18775 7115
rect 18735 7065 18775 7095
rect 18735 7045 18745 7065
rect 18765 7045 18775 7065
rect 12525 6995 12535 7015
rect 12555 6995 12565 7015
rect 18735 7015 18775 7045
rect 12525 6980 12565 6995
rect 18735 6995 18745 7015
rect 18765 6995 18775 7015
rect 18735 6980 18775 6995
rect 20025 7115 20065 7130
rect 20025 7095 20035 7115
rect 20055 7095 20065 7115
rect 20025 7065 20065 7095
rect 20025 7045 20035 7065
rect 20055 7045 20065 7065
rect 20025 7015 20065 7045
rect 20350 7105 20390 7135
rect 20350 7085 20360 7105
rect 20380 7085 20390 7105
rect 20350 7055 20390 7085
rect 20350 7035 20360 7055
rect 20380 7035 20390 7055
rect 20350 7020 20390 7035
rect 21640 7155 21680 7170
rect 21640 7135 21650 7155
rect 21670 7135 21680 7155
rect 21640 7105 21680 7135
rect 21640 7085 21650 7105
rect 21670 7085 21680 7105
rect 21640 7055 21680 7085
rect 21640 7035 21650 7055
rect 21670 7035 21680 7055
rect 21640 7020 21680 7035
rect 20025 6995 20035 7015
rect 20055 6995 20065 7015
rect 20025 6980 20065 6995
rect 20450 6840 20490 6855
rect 20450 6820 20460 6840
rect 20480 6820 20490 6840
rect 20450 6790 20490 6820
rect 20450 6770 20460 6790
rect 20480 6770 20490 6790
rect 20450 6740 20490 6770
rect 20450 6720 20460 6740
rect 20480 6720 20490 6740
rect 20450 6705 20490 6720
rect 20860 6840 20900 6855
rect 20860 6820 20870 6840
rect 20890 6820 20900 6840
rect 20860 6790 20900 6820
rect 20860 6770 20870 6790
rect 20890 6770 20900 6790
rect 20860 6740 20900 6770
rect 20860 6720 20870 6740
rect 20890 6720 20900 6740
rect 20860 6705 20900 6720
rect 10990 6650 11030 6665
rect 10990 6630 11000 6650
rect 11020 6630 11030 6650
rect 10990 6600 11030 6630
rect 10990 6580 11000 6600
rect 11020 6580 11030 6600
rect 10990 6550 11030 6580
rect 10990 6530 11000 6550
rect 11020 6530 11030 6550
rect 10990 6515 11030 6530
rect 11730 6650 11770 6665
rect 11730 6630 11740 6650
rect 11760 6630 11770 6650
rect 11730 6600 11770 6630
rect 11730 6580 11740 6600
rect 11760 6580 11770 6600
rect 11730 6550 11770 6580
rect 11730 6530 11740 6550
rect 11760 6530 11770 6550
rect 11730 6515 11770 6530
rect 12030 6650 12070 6665
rect 12030 6630 12040 6650
rect 12060 6630 12070 6650
rect 12030 6600 12070 6630
rect 12030 6580 12040 6600
rect 12060 6580 12070 6600
rect 12030 6550 12070 6580
rect 12030 6530 12040 6550
rect 12060 6530 12070 6550
rect 12030 6515 12070 6530
rect 12770 6650 12810 6665
rect 12770 6630 12780 6650
rect 12800 6630 12810 6650
rect 12770 6600 12810 6630
rect 12770 6580 12780 6600
rect 12800 6580 12810 6600
rect 12770 6550 12810 6580
rect 12770 6530 12780 6550
rect 12800 6530 12810 6550
rect 12770 6515 12810 6530
rect 18490 6650 18530 6665
rect 18490 6630 18500 6650
rect 18520 6630 18530 6650
rect 18490 6600 18530 6630
rect 18490 6580 18500 6600
rect 18520 6580 18530 6600
rect 18490 6550 18530 6580
rect 18490 6530 18500 6550
rect 18520 6530 18530 6550
rect 18490 6515 18530 6530
rect 19230 6650 19270 6665
rect 19230 6630 19240 6650
rect 19260 6630 19270 6650
rect 19230 6600 19270 6630
rect 19230 6580 19240 6600
rect 19260 6580 19270 6600
rect 19230 6550 19270 6580
rect 19230 6530 19240 6550
rect 19260 6530 19270 6550
rect 19230 6515 19270 6530
rect 19530 6650 19570 6665
rect 19530 6630 19540 6650
rect 19560 6630 19570 6650
rect 19530 6600 19570 6630
rect 19530 6580 19540 6600
rect 19560 6580 19570 6600
rect 19530 6550 19570 6580
rect 19530 6530 19540 6550
rect 19560 6530 19570 6550
rect 19530 6515 19570 6530
rect 20270 6650 20310 6665
rect 20270 6630 20280 6650
rect 20300 6630 20310 6650
rect 20270 6600 20310 6630
rect 20270 6580 20280 6600
rect 20300 6580 20310 6600
rect 20270 6550 20310 6580
rect 20270 6530 20280 6550
rect 20300 6530 20310 6550
rect 20270 6515 20310 6530
rect 20355 6505 20395 6520
rect 20355 6485 20365 6505
rect 20385 6485 20395 6505
rect 20355 6455 20395 6485
rect 20355 6435 20365 6455
rect 20385 6435 20395 6455
rect 20355 6405 20395 6435
rect 20355 6385 20365 6405
rect 20385 6385 20395 6405
rect 20355 6370 20395 6385
rect 20655 6505 20695 6520
rect 20655 6485 20665 6505
rect 20685 6485 20695 6505
rect 20655 6455 20695 6485
rect 20655 6435 20665 6455
rect 20685 6435 20695 6455
rect 20655 6405 20695 6435
rect 20655 6385 20665 6405
rect 20685 6385 20695 6405
rect 20655 6370 20695 6385
rect 20955 6505 20995 6520
rect 20955 6485 20965 6505
rect 20985 6485 20995 6505
rect 20955 6455 20995 6485
rect 20955 6435 20965 6455
rect 20985 6435 20995 6455
rect 20955 6405 20995 6435
rect 20955 6385 20965 6405
rect 20985 6385 20995 6405
rect 20955 6370 20995 6385
rect 9625 6270 9665 6285
rect 9625 6250 9635 6270
rect 9655 6250 9665 6270
rect 9625 6225 9665 6250
rect 9625 6205 9635 6225
rect 9655 6205 9665 6225
rect 9625 6180 9665 6205
rect 9625 6160 9635 6180
rect 9655 6160 9665 6180
rect 9625 6130 9665 6160
rect 9625 6110 9635 6130
rect 9655 6110 9665 6130
rect 9625 6085 9665 6110
rect 9625 6065 9635 6085
rect 9655 6065 9665 6085
rect 9625 6040 9665 6065
rect 9625 6020 9635 6040
rect 9655 6020 9665 6040
rect 9625 6005 9665 6020
rect 10905 6270 10945 6285
rect 10905 6250 10915 6270
rect 10935 6250 10945 6270
rect 12855 6270 12895 6285
rect 10905 6225 10945 6250
rect 10905 6205 10915 6225
rect 10935 6205 10945 6225
rect 10905 6180 10945 6205
rect 12855 6250 12865 6270
rect 12885 6250 12895 6270
rect 12855 6225 12895 6250
rect 12855 6205 12865 6225
rect 12885 6205 12895 6225
rect 10905 6160 10915 6180
rect 10935 6160 10945 6180
rect 10905 6130 10945 6160
rect 10905 6110 10915 6130
rect 10935 6110 10945 6130
rect 10905 6085 10945 6110
rect 10905 6065 10915 6085
rect 10935 6065 10945 6085
rect 10905 6040 10945 6065
rect 10905 6020 10915 6040
rect 10935 6020 10945 6040
rect 10905 6005 10945 6020
rect 11165 6170 11205 6185
rect 11165 6150 11175 6170
rect 11195 6150 11205 6170
rect 11165 6120 11205 6150
rect 11165 6100 11175 6120
rect 11195 6100 11205 6120
rect 11165 6070 11205 6100
rect 11165 6050 11175 6070
rect 11195 6050 11205 6070
rect 11165 6020 11205 6050
rect 11165 6000 11175 6020
rect 11195 6000 11205 6020
rect 11165 5970 11205 6000
rect 11165 5950 11175 5970
rect 11195 5950 11205 5970
rect 11165 5935 11205 5950
rect 12620 6170 12660 6185
rect 12620 6150 12630 6170
rect 12650 6150 12660 6170
rect 12620 6120 12660 6150
rect 12620 6100 12630 6120
rect 12650 6100 12660 6120
rect 12620 6070 12660 6100
rect 12620 6050 12630 6070
rect 12650 6050 12660 6070
rect 12620 6020 12660 6050
rect 12620 6000 12630 6020
rect 12650 6000 12660 6020
rect 12855 6180 12895 6205
rect 12855 6160 12865 6180
rect 12885 6160 12895 6180
rect 12855 6130 12895 6160
rect 12855 6110 12865 6130
rect 12885 6110 12895 6130
rect 12855 6085 12895 6110
rect 12855 6065 12865 6085
rect 12885 6065 12895 6085
rect 12855 6040 12895 6065
rect 12855 6020 12865 6040
rect 12885 6020 12895 6040
rect 12855 6005 12895 6020
rect 14135 6270 14175 6285
rect 14135 6250 14145 6270
rect 14165 6250 14175 6270
rect 14135 6225 14175 6250
rect 14135 6205 14145 6225
rect 14165 6205 14175 6225
rect 14135 6180 14175 6205
rect 14135 6160 14145 6180
rect 14165 6160 14175 6180
rect 14135 6130 14175 6160
rect 14135 6110 14145 6130
rect 14165 6110 14175 6130
rect 14135 6085 14175 6110
rect 14135 6065 14145 6085
rect 14165 6065 14175 6085
rect 14135 6040 14175 6065
rect 14135 6020 14145 6040
rect 14165 6020 14175 6040
rect 14135 6005 14175 6020
rect 18665 6210 18705 6225
rect 18665 6190 18675 6210
rect 18695 6190 18705 6210
rect 18665 6160 18705 6190
rect 18665 6140 18675 6160
rect 18695 6140 18705 6160
rect 18665 6110 18705 6140
rect 18665 6090 18675 6110
rect 18695 6090 18705 6110
rect 18665 6060 18705 6090
rect 18665 6040 18675 6060
rect 18695 6040 18705 6060
rect 18665 6010 18705 6040
rect 12620 5970 12660 6000
rect 12620 5950 12630 5970
rect 12650 5950 12660 5970
rect 18665 5990 18675 6010
rect 18695 5990 18705 6010
rect 18665 5975 18705 5990
rect 20120 6210 20160 6225
rect 20120 6190 20130 6210
rect 20150 6190 20160 6210
rect 20120 6160 20160 6190
rect 20120 6140 20130 6160
rect 20150 6140 20160 6160
rect 20120 6110 20160 6140
rect 20120 6090 20130 6110
rect 20150 6090 20160 6110
rect 20120 6060 20160 6090
rect 20120 6040 20130 6060
rect 20150 6040 20160 6060
rect 20120 6010 20160 6040
rect 20505 6165 20545 6180
rect 20505 6145 20515 6165
rect 20535 6145 20545 6165
rect 20505 6115 20545 6145
rect 20505 6095 20515 6115
rect 20535 6095 20545 6115
rect 20505 6065 20545 6095
rect 20505 6045 20515 6065
rect 20535 6045 20545 6065
rect 20505 6030 20545 6045
rect 20805 6165 20845 6180
rect 20805 6145 20815 6165
rect 20835 6145 20845 6165
rect 20805 6115 20845 6145
rect 20805 6095 20815 6115
rect 20835 6095 20845 6115
rect 20805 6065 20845 6095
rect 20805 6045 20815 6065
rect 20835 6045 20845 6065
rect 20805 6030 20845 6045
rect 20120 5990 20130 6010
rect 20150 5990 20160 6010
rect 20120 5975 20160 5990
rect 12620 5935 12660 5950
rect 11200 4375 11240 4403
rect 11200 4355 11210 4375
rect 11230 4355 11240 4375
rect 11200 4340 11240 4355
rect 11460 4375 11500 4403
rect 11460 4355 11470 4375
rect 11490 4355 11500 4375
rect 11460 4340 11500 4355
rect 11530 4390 11570 4420
rect 11530 4370 11540 4390
rect 11560 4370 11570 4390
rect 11530 4340 11570 4370
rect 11970 4390 12010 4420
rect 11970 4370 11980 4390
rect 12000 4370 12010 4390
rect 11970 4340 12010 4370
rect 12040 4375 12080 4395
rect 12040 4355 12050 4375
rect 12070 4355 12080 4375
rect 12040 4335 12080 4355
rect 12600 4375 12640 4395
rect 12600 4355 12610 4375
rect 12630 4355 12640 4375
rect 12600 4335 12640 4355
rect 11210 4140 11250 4155
rect 11210 4120 11220 4140
rect 11240 4120 11250 4140
rect 11210 4105 11250 4120
rect 12500 4140 12540 4155
rect 12500 4120 12510 4140
rect 12530 4120 12540 4140
rect 12500 4105 12540 4120
rect 11155 3835 11195 3850
rect 11155 3815 11165 3835
rect 11185 3815 11195 3835
rect 11155 3800 11195 3815
rect 11895 3835 11935 3850
rect 11895 3815 11905 3835
rect 11925 3815 11935 3835
rect 11895 3800 11935 3815
rect 12635 3835 12675 3850
rect 12635 3815 12645 3835
rect 12665 3815 12675 3835
rect 12635 3800 12675 3815
rect 10115 3570 10155 3585
rect 10115 3550 10125 3570
rect 10145 3550 10155 3570
rect 10115 3520 10155 3550
rect 10115 3500 10125 3520
rect 10145 3500 10155 3520
rect 10115 3470 10155 3500
rect 10115 3450 10125 3470
rect 10145 3450 10155 3470
rect 10115 3420 10155 3450
rect 10115 3400 10125 3420
rect 10145 3400 10155 3420
rect 10115 3370 10155 3400
rect 10115 3350 10125 3370
rect 10145 3350 10155 3370
rect 10115 3320 10155 3350
rect 10115 3300 10125 3320
rect 10145 3300 10155 3320
rect 10115 3270 10155 3300
rect 10115 3250 10125 3270
rect 10145 3250 10155 3270
rect 10115 3220 10155 3250
rect 10115 3200 10125 3220
rect 10145 3200 10155 3220
rect 10115 3170 10155 3200
rect 10115 3150 10125 3170
rect 10145 3150 10155 3170
rect 10115 3120 10155 3150
rect 10115 3100 10125 3120
rect 10145 3100 10155 3120
rect 10115 3070 10155 3100
rect 10115 3050 10125 3070
rect 10145 3050 10155 3070
rect 10115 3020 10155 3050
rect 10115 3000 10125 3020
rect 10145 3000 10155 3020
rect 10115 2985 10155 3000
rect 10855 3570 10895 3585
rect 10855 3550 10865 3570
rect 10885 3550 10895 3570
rect 10855 3520 10895 3550
rect 10855 3500 10865 3520
rect 10885 3500 10895 3520
rect 10855 3470 10895 3500
rect 10855 3450 10865 3470
rect 10885 3450 10895 3470
rect 10855 3420 10895 3450
rect 10855 3400 10865 3420
rect 10885 3400 10895 3420
rect 10855 3370 10895 3400
rect 10855 3350 10865 3370
rect 10885 3350 10895 3370
rect 10855 3320 10895 3350
rect 10855 3300 10865 3320
rect 10885 3300 10895 3320
rect 10855 3270 10895 3300
rect 10855 3250 10865 3270
rect 10885 3250 10895 3270
rect 10855 3220 10895 3250
rect 10855 3200 10865 3220
rect 10885 3200 10895 3220
rect 10855 3170 10895 3200
rect 11180 3560 11220 3575
rect 11180 3540 11190 3560
rect 11210 3540 11220 3560
rect 11180 3510 11220 3540
rect 11180 3490 11190 3510
rect 11210 3490 11220 3510
rect 11180 3460 11220 3490
rect 11180 3440 11190 3460
rect 11210 3440 11220 3460
rect 11180 3410 11220 3440
rect 11180 3390 11190 3410
rect 11210 3390 11220 3410
rect 11180 3360 11220 3390
rect 11180 3340 11190 3360
rect 11210 3340 11220 3360
rect 11180 3310 11220 3340
rect 11180 3290 11190 3310
rect 11210 3290 11220 3310
rect 11180 3260 11220 3290
rect 11180 3240 11190 3260
rect 11210 3240 11220 3260
rect 11180 3210 11220 3240
rect 11180 3190 11190 3210
rect 11210 3190 11220 3210
rect 11180 3175 11220 3190
rect 12580 3560 12620 3575
rect 12580 3540 12590 3560
rect 12610 3540 12620 3560
rect 12580 3510 12620 3540
rect 12580 3490 12590 3510
rect 12610 3490 12620 3510
rect 12580 3460 12620 3490
rect 12580 3440 12590 3460
rect 12610 3440 12620 3460
rect 12580 3410 12620 3440
rect 12580 3390 12590 3410
rect 12610 3390 12620 3410
rect 12580 3360 12620 3390
rect 12580 3340 12590 3360
rect 12610 3340 12620 3360
rect 12580 3310 12620 3340
rect 12580 3290 12590 3310
rect 12610 3290 12620 3310
rect 12580 3260 12620 3290
rect 12580 3240 12590 3260
rect 12610 3240 12620 3260
rect 12580 3210 12620 3240
rect 12580 3190 12590 3210
rect 12610 3190 12620 3210
rect 12580 3175 12620 3190
rect 12905 3570 12945 3585
rect 12905 3550 12915 3570
rect 12935 3550 12945 3570
rect 12905 3520 12945 3550
rect 12905 3500 12915 3520
rect 12935 3500 12945 3520
rect 12905 3470 12945 3500
rect 12905 3450 12915 3470
rect 12935 3450 12945 3470
rect 12905 3420 12945 3450
rect 12905 3400 12915 3420
rect 12935 3400 12945 3420
rect 12905 3370 12945 3400
rect 12905 3350 12915 3370
rect 12935 3350 12945 3370
rect 12905 3320 12945 3350
rect 12905 3300 12915 3320
rect 12935 3300 12945 3320
rect 12905 3270 12945 3300
rect 12905 3250 12915 3270
rect 12935 3250 12945 3270
rect 12905 3220 12945 3250
rect 12905 3200 12915 3220
rect 12935 3200 12945 3220
rect 10855 3150 10865 3170
rect 10885 3150 10895 3170
rect 12905 3170 12945 3200
rect 12905 3150 12915 3170
rect 12935 3150 12945 3170
rect 10855 3120 10895 3150
rect 12905 3120 12945 3150
rect 10855 3100 10865 3120
rect 10885 3100 10895 3120
rect 10855 3070 10895 3100
rect 10855 3050 10865 3070
rect 10885 3050 10895 3070
rect 10855 3020 10895 3050
rect 10855 3000 10865 3020
rect 10885 3000 10895 3020
rect 10855 2985 10895 3000
rect 12905 3100 12915 3120
rect 12935 3100 12945 3120
rect 12905 3070 12945 3100
rect 12905 3050 12915 3070
rect 12935 3050 12945 3070
rect 12905 3020 12945 3050
rect 12905 3000 12915 3020
rect 12935 3000 12945 3020
rect 12905 2985 12945 3000
rect 13645 3570 13685 3585
rect 13645 3550 13655 3570
rect 13675 3550 13685 3570
rect 13645 3520 13685 3550
rect 13645 3500 13655 3520
rect 13675 3500 13685 3520
rect 13645 3470 13685 3500
rect 13645 3450 13655 3470
rect 13675 3450 13685 3470
rect 13645 3420 13685 3450
rect 13645 3400 13655 3420
rect 13675 3400 13685 3420
rect 13645 3370 13685 3400
rect 13645 3350 13655 3370
rect 13675 3350 13685 3370
rect 13645 3320 13685 3350
rect 13645 3300 13655 3320
rect 13675 3300 13685 3320
rect 13645 3270 13685 3300
rect 13645 3250 13655 3270
rect 13675 3250 13685 3270
rect 13645 3220 13685 3250
rect 13645 3200 13655 3220
rect 13675 3200 13685 3220
rect 13645 3170 13685 3200
rect 13645 3150 13655 3170
rect 13675 3150 13685 3170
rect 13645 3120 13685 3150
rect 13645 3100 13655 3120
rect 13675 3100 13685 3120
rect 13645 3070 13685 3100
rect 13645 3050 13655 3070
rect 13675 3050 13685 3070
rect 13645 3020 13685 3050
rect 13645 3000 13655 3020
rect 13675 3000 13685 3020
rect 13645 2985 13685 3000
rect 25780 3515 25820 3550
rect 25780 3495 25790 3515
rect 25810 3495 25820 3515
rect 25780 3465 25820 3495
rect 25780 3445 25790 3465
rect 25810 3445 25820 3465
rect 25780 3415 25820 3445
rect 25780 3395 25790 3415
rect 25810 3395 25820 3415
rect 25780 3365 25820 3395
rect 25780 3345 25790 3365
rect 25810 3345 25820 3365
rect 25780 3315 25820 3345
rect 25780 3295 25790 3315
rect 25810 3295 25820 3315
rect 25450 3265 25490 3293
rect 25450 3245 25460 3265
rect 25480 3245 25490 3265
rect 25450 3230 25490 3245
rect 25710 3265 25750 3293
rect 25710 3245 25720 3265
rect 25740 3245 25750 3265
rect 25710 3230 25750 3245
rect 25780 3265 25820 3295
rect 25780 3245 25790 3265
rect 25810 3245 25820 3265
rect 25780 3230 25820 3245
rect 26100 3565 26140 3580
rect 26100 3545 26110 3565
rect 26130 3545 26140 3565
rect 26100 3515 26140 3545
rect 26100 3495 26110 3515
rect 26130 3495 26140 3515
rect 26100 3465 26140 3495
rect 26100 3445 26110 3465
rect 26130 3445 26140 3465
rect 26100 3415 26140 3445
rect 26100 3395 26110 3415
rect 26130 3395 26140 3415
rect 26100 3365 26140 3395
rect 26100 3345 26110 3365
rect 26130 3345 26140 3365
rect 26100 3315 26140 3345
rect 26100 3295 26110 3315
rect 26130 3295 26140 3315
rect 26100 3265 26140 3295
rect 26100 3245 26110 3265
rect 26130 3245 26140 3265
rect 26100 3230 26140 3245
rect 26180 3560 26220 3575
rect 26180 3540 26190 3560
rect 26210 3540 26220 3560
rect 26180 3510 26220 3540
rect 26180 3490 26190 3510
rect 26210 3490 26220 3510
rect 26180 3460 26220 3490
rect 26180 3440 26190 3460
rect 26210 3440 26220 3460
rect 26180 3410 26220 3440
rect 26180 3390 26190 3410
rect 26210 3390 26220 3410
rect 26180 3360 26220 3390
rect 26180 3340 26190 3360
rect 26210 3340 26220 3360
rect 26180 3310 26220 3340
rect 26180 3290 26190 3310
rect 26210 3290 26220 3310
rect 26180 3260 26220 3290
rect 26180 3240 26190 3260
rect 26210 3240 26220 3260
rect 26180 3210 26220 3240
rect 26180 3190 26190 3210
rect 26210 3190 26220 3210
rect 26180 3175 26220 3190
rect 27580 3560 27620 3575
rect 27580 3540 27590 3560
rect 27610 3540 27620 3560
rect 27580 3510 27620 3540
rect 27580 3490 27590 3510
rect 27610 3490 27620 3510
rect 27580 3460 27620 3490
rect 27580 3440 27590 3460
rect 27610 3440 27620 3460
rect 27580 3410 27620 3440
rect 27580 3390 27590 3410
rect 27610 3390 27620 3410
rect 27580 3360 27620 3390
rect 27580 3340 27590 3360
rect 27610 3340 27620 3360
rect 27580 3310 27620 3340
rect 27580 3290 27590 3310
rect 27610 3290 27620 3310
rect 27580 3260 27620 3290
rect 27580 3240 27590 3260
rect 27610 3240 27620 3260
rect 27580 3210 27620 3240
rect 27580 3190 27590 3210
rect 27610 3190 27620 3210
rect 27580 3175 27620 3190
rect 27850 3225 27890 3240
rect 27850 3205 27860 3225
rect 27880 3205 27890 3225
rect 27850 3175 27890 3205
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 27850 3155 27860 3175
rect 27880 3155 27890 3175
rect 27850 3125 27890 3155
rect 27850 3105 27860 3125
rect 27880 3105 27890 3125
rect 27850 3075 27890 3105
rect 27850 3055 27860 3075
rect 27880 3055 27890 3075
rect 27850 3025 27890 3055
rect 27850 3005 27860 3025
rect 27880 3005 27890 3025
rect 27850 2975 27890 3005
rect 27850 2955 27860 2975
rect 27880 2955 27890 2975
rect 27850 2940 27890 2955
rect 29140 3225 29180 3240
rect 29140 3205 29150 3225
rect 29170 3205 29180 3225
rect 29140 3175 29180 3205
rect 29140 3155 29150 3175
rect 29170 3155 29180 3175
rect 29140 3125 29180 3155
rect 29140 3105 29150 3125
rect 29170 3105 29180 3125
rect 29140 3075 29180 3105
rect 29140 3055 29150 3075
rect 29170 3055 29180 3075
rect 29140 3025 29180 3055
rect 29140 3005 29150 3025
rect 29170 3005 29180 3025
rect 29140 2975 29180 3005
rect 29140 2955 29150 2975
rect 29170 2955 29180 2975
rect 29140 2940 29180 2955
rect 11180 2880 11220 2895
rect 11180 2860 11190 2880
rect 11210 2860 11220 2880
rect 11180 2830 11220 2860
rect 11180 2810 11190 2830
rect 11210 2810 11220 2830
rect 11180 2780 11220 2810
rect 11180 2760 11190 2780
rect 11210 2760 11220 2780
rect 11180 2730 11220 2760
rect 11180 2710 11190 2730
rect 11210 2710 11220 2730
rect 11180 2680 11220 2710
rect 11180 2660 11190 2680
rect 11210 2660 11220 2680
rect 10115 2640 10155 2655
rect 10115 2620 10125 2640
rect 10145 2620 10155 2640
rect 10115 2590 10155 2620
rect 10115 2570 10125 2590
rect 10145 2570 10155 2590
rect 10115 2540 10155 2570
rect 10115 2520 10125 2540
rect 10145 2520 10155 2540
rect 10115 2490 10155 2520
rect 10115 2470 10125 2490
rect 10145 2470 10155 2490
rect 10115 2455 10155 2470
rect 10855 2640 10895 2655
rect 10855 2620 10865 2640
rect 10885 2620 10895 2640
rect 10855 2590 10895 2620
rect 10855 2570 10865 2590
rect 10885 2570 10895 2590
rect 10855 2540 10895 2570
rect 10855 2520 10865 2540
rect 10885 2520 10895 2540
rect 10855 2490 10895 2520
rect 11180 2630 11220 2660
rect 11180 2610 11190 2630
rect 11210 2610 11220 2630
rect 11180 2580 11220 2610
rect 11180 2560 11190 2580
rect 11210 2560 11220 2580
rect 11180 2530 11220 2560
rect 11180 2510 11190 2530
rect 11210 2510 11220 2530
rect 11180 2495 11220 2510
rect 12580 2880 12620 2895
rect 12580 2860 12590 2880
rect 12610 2860 12620 2880
rect 12580 2830 12620 2860
rect 12580 2810 12590 2830
rect 12610 2810 12620 2830
rect 12580 2780 12620 2810
rect 12580 2760 12590 2780
rect 12610 2760 12620 2780
rect 12580 2730 12620 2760
rect 12580 2710 12590 2730
rect 12610 2710 12620 2730
rect 12580 2680 12620 2710
rect 12580 2660 12590 2680
rect 12610 2660 12620 2680
rect 26180 2880 26220 2895
rect 26180 2860 26190 2880
rect 26210 2860 26220 2880
rect 26180 2830 26220 2860
rect 26180 2810 26190 2830
rect 26210 2810 26220 2830
rect 26180 2780 26220 2810
rect 26180 2760 26190 2780
rect 26210 2760 26220 2780
rect 26180 2730 26220 2760
rect 26180 2710 26190 2730
rect 26210 2710 26220 2730
rect 26180 2680 26220 2710
rect 12580 2630 12620 2660
rect 26180 2660 26190 2680
rect 26210 2660 26220 2680
rect 12580 2610 12590 2630
rect 12610 2610 12620 2630
rect 12580 2580 12620 2610
rect 12580 2560 12590 2580
rect 12610 2560 12620 2580
rect 12580 2530 12620 2560
rect 12580 2510 12590 2530
rect 12610 2510 12620 2530
rect 12580 2495 12620 2510
rect 12905 2640 12945 2655
rect 12905 2620 12915 2640
rect 12935 2620 12945 2640
rect 12905 2590 12945 2620
rect 12905 2570 12915 2590
rect 12935 2570 12945 2590
rect 12905 2540 12945 2570
rect 12905 2520 12915 2540
rect 12935 2520 12945 2540
rect 10855 2470 10865 2490
rect 10885 2470 10895 2490
rect 12905 2490 12945 2520
rect 12905 2470 12915 2490
rect 12935 2470 12945 2490
rect 10855 2455 10895 2470
rect 12905 2455 12945 2470
rect 13645 2640 13685 2655
rect 13645 2620 13655 2640
rect 13675 2620 13685 2640
rect 13645 2590 13685 2620
rect 13645 2570 13655 2590
rect 13675 2570 13685 2590
rect 13645 2540 13685 2570
rect 13645 2520 13655 2540
rect 13675 2520 13685 2540
rect 13645 2490 13685 2520
rect 13645 2470 13655 2490
rect 13675 2470 13685 2490
rect 13645 2455 13685 2470
rect 10115 2250 10155 2265
rect 10115 2230 10125 2250
rect 10145 2230 10155 2250
rect 10115 2200 10155 2230
rect 10115 2180 10125 2200
rect 10145 2180 10155 2200
rect 10115 2150 10155 2180
rect 10115 2130 10125 2150
rect 10145 2130 10155 2150
rect 10115 2100 10155 2130
rect 10115 2080 10125 2100
rect 10145 2080 10155 2100
rect 10115 2050 10155 2080
rect 10115 2030 10125 2050
rect 10145 2030 10155 2050
rect 10115 2000 10155 2030
rect 10115 1980 10125 2000
rect 10145 1980 10155 2000
rect 10115 1965 10155 1980
rect 10855 2250 10895 2265
rect 10855 2230 10865 2250
rect 10885 2230 10895 2250
rect 10855 2200 10895 2230
rect 10855 2180 10865 2200
rect 10885 2180 10895 2200
rect 12905 2250 12945 2265
rect 12905 2230 12915 2250
rect 12935 2230 12945 2250
rect 12905 2200 12945 2230
rect 10855 2150 10895 2180
rect 12905 2180 12915 2200
rect 12935 2180 12945 2200
rect 10855 2130 10865 2150
rect 10885 2130 10895 2150
rect 12905 2150 12945 2180
rect 12905 2130 12915 2150
rect 12935 2130 12945 2150
rect 10855 2100 10895 2130
rect 10855 2080 10865 2100
rect 10885 2080 10895 2100
rect 10855 2050 10895 2080
rect 10855 2030 10865 2050
rect 10885 2030 10895 2050
rect 10855 2000 10895 2030
rect 10855 1980 10865 2000
rect 10885 1980 10895 2000
rect 11235 2115 11275 2130
rect 11235 2095 11245 2115
rect 11265 2095 11275 2115
rect 11235 2065 11275 2095
rect 11235 2045 11245 2065
rect 11265 2045 11275 2065
rect 11235 2015 11275 2045
rect 11235 1995 11245 2015
rect 11265 1995 11275 2015
rect 11235 1980 11275 1995
rect 12525 2115 12565 2130
rect 12525 2095 12535 2115
rect 12555 2095 12565 2115
rect 12525 2065 12565 2095
rect 12525 2045 12535 2065
rect 12555 2045 12565 2065
rect 12525 2015 12565 2045
rect 12525 1995 12535 2015
rect 12555 1995 12565 2015
rect 12525 1980 12565 1995
rect 12905 2100 12945 2130
rect 12905 2080 12915 2100
rect 12935 2080 12945 2100
rect 12905 2050 12945 2080
rect 12905 2030 12915 2050
rect 12935 2030 12945 2050
rect 12905 2000 12945 2030
rect 12905 1980 12915 2000
rect 12935 1980 12945 2000
rect 10855 1965 10895 1980
rect 12905 1965 12945 1980
rect 13645 2250 13685 2265
rect 13645 2230 13655 2250
rect 13675 2230 13685 2250
rect 13645 2200 13685 2230
rect 13645 2180 13655 2200
rect 13675 2180 13685 2200
rect 13645 2150 13685 2180
rect 13645 2130 13655 2150
rect 13675 2130 13685 2150
rect 13645 2100 13685 2130
rect 13645 2080 13655 2100
rect 13675 2080 13685 2100
rect 13645 2050 13685 2080
rect 13645 2030 13655 2050
rect 13675 2030 13685 2050
rect 13645 2000 13685 2030
rect 26180 2630 26220 2660
rect 24640 2605 24680 2620
rect 24640 2585 24650 2605
rect 24670 2585 24680 2605
rect 24640 2555 24680 2585
rect 24640 2535 24650 2555
rect 24670 2535 24680 2555
rect 24640 2520 24680 2535
rect 25930 2605 25970 2620
rect 25930 2585 25940 2605
rect 25960 2585 25970 2605
rect 25930 2555 25970 2585
rect 25930 2535 25940 2555
rect 25960 2535 25970 2555
rect 25930 2520 25970 2535
rect 26180 2610 26190 2630
rect 26210 2610 26220 2630
rect 26180 2580 26220 2610
rect 26180 2560 26190 2580
rect 26210 2560 26220 2580
rect 26180 2530 26220 2560
rect 26180 2510 26190 2530
rect 26210 2510 26220 2530
rect 26180 2495 26220 2510
rect 27580 2880 27620 2895
rect 27580 2860 27590 2880
rect 27610 2860 27620 2880
rect 27580 2830 27620 2860
rect 27580 2810 27590 2830
rect 27610 2810 27620 2830
rect 27580 2780 27620 2810
rect 27580 2760 27590 2780
rect 27610 2760 27620 2780
rect 27580 2730 27620 2760
rect 27580 2710 27590 2730
rect 27610 2710 27620 2730
rect 27580 2680 27620 2710
rect 27580 2660 27590 2680
rect 27610 2660 27620 2680
rect 27580 2630 27620 2660
rect 27580 2610 27590 2630
rect 27610 2610 27620 2630
rect 27580 2580 27620 2610
rect 27580 2560 27590 2580
rect 27610 2560 27620 2580
rect 27580 2530 27620 2560
rect 27580 2510 27590 2530
rect 27610 2510 27620 2530
rect 27850 2605 27890 2620
rect 27850 2585 27860 2605
rect 27880 2585 27890 2605
rect 27850 2555 27890 2585
rect 27850 2535 27860 2555
rect 27880 2535 27890 2555
rect 27850 2520 27890 2535
rect 29140 2605 29180 2620
rect 29140 2585 29150 2605
rect 29170 2585 29180 2605
rect 29140 2555 29180 2585
rect 29140 2535 29150 2555
rect 29170 2535 29180 2555
rect 29140 2520 29180 2535
rect 27580 2495 27620 2510
rect 24640 2155 24680 2170
rect 24640 2135 24650 2155
rect 24670 2135 24680 2155
rect 24640 2105 24680 2135
rect 24640 2085 24650 2105
rect 24670 2085 24680 2105
rect 24640 2055 24680 2085
rect 24640 2035 24650 2055
rect 24670 2035 24680 2055
rect 24640 2020 24680 2035
rect 25930 2155 25970 2170
rect 27850 2155 27890 2170
rect 25930 2135 25940 2155
rect 25960 2135 25970 2155
rect 25930 2105 25970 2135
rect 27850 2135 27860 2155
rect 27880 2135 27890 2155
rect 25930 2085 25940 2105
rect 25960 2085 25970 2105
rect 25930 2055 25970 2085
rect 25930 2035 25940 2055
rect 25960 2035 25970 2055
rect 25930 2020 25970 2035
rect 26235 2115 26275 2130
rect 26235 2095 26245 2115
rect 26265 2095 26275 2115
rect 26235 2065 26275 2095
rect 26235 2045 26245 2065
rect 26265 2045 26275 2065
rect 26235 2015 26275 2045
rect 13645 1980 13655 2000
rect 13675 1980 13685 2000
rect 26235 1995 26245 2015
rect 26265 1995 26275 2015
rect 26235 1980 26275 1995
rect 27525 2115 27565 2130
rect 27525 2095 27535 2115
rect 27555 2095 27565 2115
rect 27525 2065 27565 2095
rect 27525 2045 27535 2065
rect 27555 2045 27565 2065
rect 27525 2015 27565 2045
rect 27850 2105 27890 2135
rect 27850 2085 27860 2105
rect 27880 2085 27890 2105
rect 27850 2055 27890 2085
rect 27850 2035 27860 2055
rect 27880 2035 27890 2055
rect 27850 2020 27890 2035
rect 29140 2155 29180 2170
rect 29140 2135 29150 2155
rect 29170 2135 29180 2155
rect 29140 2105 29180 2135
rect 29140 2085 29150 2105
rect 29170 2085 29180 2105
rect 29140 2055 29180 2085
rect 29140 2035 29150 2055
rect 29170 2035 29180 2055
rect 29140 2020 29180 2035
rect 27525 1995 27535 2015
rect 27555 1995 27565 2015
rect 27525 1980 27565 1995
rect 13645 1965 13685 1980
rect 27950 1840 27990 1855
rect 27950 1820 27960 1840
rect 27980 1820 27990 1840
rect 27950 1790 27990 1820
rect 27950 1770 27960 1790
rect 27980 1770 27990 1790
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect 27950 1740 27990 1770
rect 27950 1720 27960 1740
rect 27980 1720 27990 1740
rect -50 1680 100 1695
rect 27950 1705 27990 1720
rect 28360 1840 28400 1855
rect 28360 1820 28370 1840
rect 28390 1820 28400 1840
rect 28360 1790 28400 1820
rect 28360 1770 28370 1790
rect 28390 1770 28400 1790
rect 28360 1740 28400 1770
rect 28360 1720 28370 1740
rect 28390 1720 28400 1740
rect 28360 1705 28400 1720
rect 3980 1650 4030 1665
rect 3980 1630 3995 1650
rect 4015 1630 4030 1650
rect 3980 1615 4030 1630
rect 10115 1640 10155 1655
rect 10115 1620 10125 1640
rect 10145 1620 10155 1640
rect 5065 1060 5105 1075
rect 5065 1040 5075 1060
rect 5095 1040 5105 1060
rect 5065 1010 5105 1040
rect 5065 990 5075 1010
rect 5095 990 5105 1010
rect 5065 975 5105 990
rect 10115 1590 10155 1620
rect 10115 1570 10125 1590
rect 10145 1570 10155 1590
rect 10115 1540 10155 1570
rect 10115 1520 10125 1540
rect 10145 1520 10155 1540
rect 10115 1490 10155 1520
rect 10115 1470 10125 1490
rect 10145 1470 10155 1490
rect 10115 1440 10155 1470
rect 10115 1420 10125 1440
rect 10145 1420 10155 1440
rect 10115 1390 10155 1420
rect 10115 1370 10125 1390
rect 10145 1370 10155 1390
rect 10115 1340 10155 1370
rect 10115 1320 10125 1340
rect 10145 1320 10155 1340
rect 10115 1290 10155 1320
rect 10115 1270 10125 1290
rect 10145 1270 10155 1290
rect 10115 1240 10155 1270
rect 10115 1220 10125 1240
rect 10145 1220 10155 1240
rect 10115 1190 10155 1220
rect 10115 1170 10125 1190
rect 10145 1170 10155 1190
rect 10115 1140 10155 1170
rect 10115 1120 10125 1140
rect 10145 1120 10155 1140
rect 10115 1090 10155 1120
rect 10115 1070 10125 1090
rect 10145 1070 10155 1090
rect 10115 1040 10155 1070
rect 10115 1020 10125 1040
rect 10145 1020 10155 1040
rect 10115 990 10155 1020
rect 10115 970 10125 990
rect 10145 970 10155 990
rect 10115 955 10155 970
rect 10795 1640 10835 1655
rect 10795 1620 10805 1640
rect 10825 1620 10835 1640
rect 10795 1590 10835 1620
rect 10795 1570 10805 1590
rect 10825 1570 10835 1590
rect 10795 1540 10835 1570
rect 10795 1520 10805 1540
rect 10825 1520 10835 1540
rect 10795 1490 10835 1520
rect 10990 1650 11030 1665
rect 10990 1630 11000 1650
rect 11020 1630 11030 1650
rect 10990 1600 11030 1630
rect 10990 1580 11000 1600
rect 11020 1580 11030 1600
rect 10990 1550 11030 1580
rect 10990 1530 11000 1550
rect 11020 1530 11030 1550
rect 10990 1515 11030 1530
rect 11730 1650 11770 1665
rect 11730 1630 11740 1650
rect 11760 1630 11770 1650
rect 11730 1600 11770 1630
rect 11730 1580 11740 1600
rect 11760 1580 11770 1600
rect 11730 1550 11770 1580
rect 11730 1530 11740 1550
rect 11760 1530 11770 1550
rect 11730 1515 11770 1530
rect 12030 1650 12070 1665
rect 12030 1630 12040 1650
rect 12060 1630 12070 1650
rect 12030 1600 12070 1630
rect 12030 1580 12040 1600
rect 12060 1580 12070 1600
rect 12030 1550 12070 1580
rect 12030 1530 12040 1550
rect 12060 1530 12070 1550
rect 12030 1515 12070 1530
rect 12770 1650 12810 1665
rect 12770 1630 12780 1650
rect 12800 1630 12810 1650
rect 12770 1600 12810 1630
rect 12770 1580 12780 1600
rect 12800 1580 12810 1600
rect 12770 1550 12810 1580
rect 12770 1530 12780 1550
rect 12800 1530 12810 1550
rect 12770 1515 12810 1530
rect 12965 1640 13005 1655
rect 12965 1620 12975 1640
rect 12995 1620 13005 1640
rect 12965 1590 13005 1620
rect 12965 1570 12975 1590
rect 12995 1570 13005 1590
rect 12965 1540 13005 1570
rect 12965 1520 12975 1540
rect 12995 1520 13005 1540
rect 10795 1470 10805 1490
rect 10825 1470 10835 1490
rect 10795 1440 10835 1470
rect 12965 1490 13005 1520
rect 12965 1470 12975 1490
rect 12995 1470 13005 1490
rect 10795 1420 10805 1440
rect 10825 1420 10835 1440
rect 10795 1390 10835 1420
rect 10795 1370 10805 1390
rect 10825 1370 10835 1390
rect 10795 1340 10835 1370
rect 10795 1320 10805 1340
rect 10825 1320 10835 1340
rect 10795 1290 10835 1320
rect 10795 1270 10805 1290
rect 10825 1270 10835 1290
rect 10795 1240 10835 1270
rect 12965 1440 13005 1470
rect 12965 1420 12975 1440
rect 12995 1420 13005 1440
rect 12965 1390 13005 1420
rect 12965 1370 12975 1390
rect 12995 1370 13005 1390
rect 12965 1340 13005 1370
rect 12965 1320 12975 1340
rect 12995 1320 13005 1340
rect 12965 1290 13005 1320
rect 12965 1270 12975 1290
rect 12995 1270 13005 1290
rect 10795 1220 10805 1240
rect 10825 1220 10835 1240
rect 10795 1190 10835 1220
rect 10795 1170 10805 1190
rect 10825 1170 10835 1190
rect 12965 1240 13005 1270
rect 12965 1220 12975 1240
rect 12995 1220 13005 1240
rect 12965 1190 13005 1220
rect 10795 1140 10835 1170
rect 10795 1120 10805 1140
rect 10825 1120 10835 1140
rect 10795 1090 10835 1120
rect 10795 1070 10805 1090
rect 10825 1070 10835 1090
rect 10795 1040 10835 1070
rect 10795 1020 10805 1040
rect 10825 1020 10835 1040
rect 10795 990 10835 1020
rect 10795 970 10805 990
rect 10825 970 10835 990
rect 10795 955 10835 970
rect 11165 1170 11205 1185
rect 11165 1150 11175 1170
rect 11195 1150 11205 1170
rect 11165 1120 11205 1150
rect 11165 1100 11175 1120
rect 11195 1100 11205 1120
rect 11165 1070 11205 1100
rect 11165 1050 11175 1070
rect 11195 1050 11205 1070
rect 11165 1020 11205 1050
rect 11165 1000 11175 1020
rect 11195 1000 11205 1020
rect 11165 970 11205 1000
rect 11165 950 11175 970
rect 11195 950 11205 970
rect 11165 935 11205 950
rect 12620 1170 12660 1185
rect 12620 1150 12630 1170
rect 12650 1150 12660 1170
rect 12620 1120 12660 1150
rect 12620 1100 12630 1120
rect 12650 1100 12660 1120
rect 12620 1070 12660 1100
rect 12620 1050 12630 1070
rect 12650 1050 12660 1070
rect 12620 1020 12660 1050
rect 12620 1000 12630 1020
rect 12650 1000 12660 1020
rect 12620 970 12660 1000
rect 12620 950 12630 970
rect 12650 950 12660 970
rect 12965 1170 12975 1190
rect 12995 1170 13005 1190
rect 12965 1140 13005 1170
rect 12965 1120 12975 1140
rect 12995 1120 13005 1140
rect 12965 1090 13005 1120
rect 12965 1070 12975 1090
rect 12995 1070 13005 1090
rect 12965 1040 13005 1070
rect 12965 1020 12975 1040
rect 12995 1020 13005 1040
rect 12965 990 13005 1020
rect 12965 970 12975 990
rect 12995 970 13005 990
rect 12965 955 13005 970
rect 13645 1640 13685 1655
rect 13645 1620 13655 1640
rect 13675 1620 13685 1640
rect 13645 1590 13685 1620
rect 25990 1650 26030 1665
rect 25990 1630 26000 1650
rect 26020 1630 26030 1650
rect 13645 1570 13655 1590
rect 13675 1570 13685 1590
rect 13645 1540 13685 1570
rect 13645 1520 13655 1540
rect 13675 1520 13685 1540
rect 13645 1490 13685 1520
rect 13645 1470 13655 1490
rect 13675 1470 13685 1490
rect 13645 1440 13685 1470
rect 13645 1420 13655 1440
rect 13675 1420 13685 1440
rect 13645 1390 13685 1420
rect 13645 1370 13655 1390
rect 13675 1370 13685 1390
rect 13645 1340 13685 1370
rect 13645 1320 13655 1340
rect 13675 1320 13685 1340
rect 13645 1290 13685 1320
rect 13645 1270 13655 1290
rect 13675 1270 13685 1290
rect 13645 1240 13685 1270
rect 13645 1220 13655 1240
rect 13675 1220 13685 1240
rect 13645 1190 13685 1220
rect 13645 1170 13655 1190
rect 13675 1170 13685 1190
rect 13645 1140 13685 1170
rect 13645 1120 13655 1140
rect 13675 1120 13685 1140
rect 13645 1090 13685 1120
rect 13645 1070 13655 1090
rect 13675 1070 13685 1090
rect 13645 1040 13685 1070
rect 13645 1020 13655 1040
rect 13675 1020 13685 1040
rect 13645 990 13685 1020
rect 13645 970 13655 990
rect 13675 970 13685 990
rect 13645 955 13685 970
rect 12620 935 12660 950
rect 25990 1600 26030 1630
rect 25990 1580 26000 1600
rect 26020 1580 26030 1600
rect 25990 1550 26030 1580
rect 25990 1530 26000 1550
rect 26020 1530 26030 1550
rect 25990 1515 26030 1530
rect 26730 1650 26770 1665
rect 26730 1630 26740 1650
rect 26760 1630 26770 1650
rect 26730 1600 26770 1630
rect 26730 1580 26740 1600
rect 26760 1580 26770 1600
rect 26730 1550 26770 1580
rect 26730 1530 26740 1550
rect 26760 1530 26770 1550
rect 26730 1515 26770 1530
rect 27030 1650 27070 1665
rect 27030 1630 27040 1650
rect 27060 1630 27070 1650
rect 27030 1600 27070 1630
rect 27030 1580 27040 1600
rect 27060 1580 27070 1600
rect 27030 1550 27070 1580
rect 27030 1530 27040 1550
rect 27060 1530 27070 1550
rect 27030 1515 27070 1530
rect 27770 1650 27810 1665
rect 27770 1630 27780 1650
rect 27800 1630 27810 1650
rect 27770 1600 27810 1630
rect 27770 1580 27780 1600
rect 27800 1580 27810 1600
rect 27770 1550 27810 1580
rect 27770 1530 27780 1550
rect 27800 1530 27810 1550
rect 27770 1515 27810 1530
rect 27855 1505 27895 1520
rect 27855 1485 27865 1505
rect 27885 1485 27895 1505
rect 27855 1455 27895 1485
rect 27855 1435 27865 1455
rect 27885 1435 27895 1455
rect 27855 1405 27895 1435
rect 27855 1385 27865 1405
rect 27885 1385 27895 1405
rect 27855 1370 27895 1385
rect 28155 1505 28195 1520
rect 28155 1485 28165 1505
rect 28185 1485 28195 1505
rect 28155 1455 28195 1485
rect 28155 1435 28165 1455
rect 28185 1435 28195 1455
rect 28155 1405 28195 1435
rect 28155 1385 28165 1405
rect 28185 1385 28195 1405
rect 28155 1370 28195 1385
rect 28455 1505 28495 1520
rect 28455 1485 28465 1505
rect 28485 1485 28495 1505
rect 28455 1455 28495 1485
rect 28455 1435 28465 1455
rect 28485 1435 28495 1455
rect 28455 1405 28495 1435
rect 28455 1385 28465 1405
rect 28485 1385 28495 1405
rect 28455 1370 28495 1385
rect 26165 1210 26205 1225
rect 26165 1190 26175 1210
rect 26195 1190 26205 1210
rect 26165 1160 26205 1190
rect 26165 1140 26175 1160
rect 26195 1140 26205 1160
rect 26165 1110 26205 1140
rect 26165 1090 26175 1110
rect 26195 1090 26205 1110
rect 26165 1060 26205 1090
rect 26165 1040 26175 1060
rect 26195 1040 26205 1060
rect 26165 1010 26205 1040
rect 26165 990 26175 1010
rect 26195 990 26205 1010
rect 26165 975 26205 990
rect 27620 1210 27660 1225
rect 27620 1190 27630 1210
rect 27650 1190 27660 1210
rect 27620 1160 27660 1190
rect 27620 1140 27630 1160
rect 27650 1140 27660 1160
rect 27620 1110 27660 1140
rect 27620 1090 27630 1110
rect 27650 1090 27660 1110
rect 27620 1060 27660 1090
rect 27620 1040 27630 1060
rect 27650 1040 27660 1060
rect 27620 1010 27660 1040
rect 28005 1165 28045 1180
rect 28005 1145 28015 1165
rect 28035 1145 28045 1165
rect 28005 1115 28045 1145
rect 28005 1095 28015 1115
rect 28035 1095 28045 1115
rect 28005 1065 28045 1095
rect 28005 1045 28015 1065
rect 28035 1045 28045 1065
rect 28005 1030 28045 1045
rect 28305 1165 28345 1180
rect 28305 1145 28315 1165
rect 28335 1145 28345 1165
rect 28305 1115 28345 1145
rect 28305 1095 28315 1115
rect 28335 1095 28345 1115
rect 28305 1065 28345 1095
rect 28305 1045 28315 1065
rect 28335 1045 28345 1065
rect 28305 1030 28345 1045
rect 27620 990 27630 1010
rect 27650 990 27660 1010
rect 27620 975 27660 990
rect 2955 865 2995 880
rect 2955 845 2965 865
rect 2985 845 2995 865
rect 2955 815 2995 845
rect 2955 795 2965 815
rect 2985 795 2995 815
rect 2955 780 2995 795
rect 5015 865 5055 880
rect 5015 845 5025 865
rect 5045 845 5055 865
rect 5015 815 5055 845
rect 5015 795 5025 815
rect 5045 795 5055 815
rect 5015 780 5055 795
rect 11840 735 11880 750
rect 11840 715 11850 735
rect 11870 715 11880 735
rect 11840 700 11880 715
rect 12580 735 12620 750
rect 12580 715 12590 735
rect 12610 715 12620 735
rect 12580 700 12620 715
rect 10780 -1485 10820 -1450
rect 10780 -1505 10790 -1485
rect 10810 -1505 10820 -1485
rect 10780 -1535 10820 -1505
rect 10780 -1555 10790 -1535
rect 10810 -1555 10820 -1535
rect 10780 -1585 10820 -1555
rect 10780 -1605 10790 -1585
rect 10810 -1605 10820 -1585
rect 10780 -1635 10820 -1605
rect 10780 -1655 10790 -1635
rect 10810 -1655 10820 -1635
rect 10780 -1685 10820 -1655
rect 10780 -1705 10790 -1685
rect 10810 -1705 10820 -1685
rect 10450 -1735 10490 -1707
rect 10450 -1755 10460 -1735
rect 10480 -1755 10490 -1735
rect 10450 -1770 10490 -1755
rect 10710 -1735 10750 -1707
rect 10710 -1755 10720 -1735
rect 10740 -1755 10750 -1735
rect 10710 -1770 10750 -1755
rect 10780 -1735 10820 -1705
rect 10780 -1755 10790 -1735
rect 10810 -1755 10820 -1735
rect 10780 -1770 10820 -1755
rect 11100 -1435 11140 -1420
rect 11100 -1455 11110 -1435
rect 11130 -1455 11140 -1435
rect 11100 -1485 11140 -1455
rect 11100 -1505 11110 -1485
rect 11130 -1505 11140 -1485
rect 11100 -1535 11140 -1505
rect 11100 -1555 11110 -1535
rect 11130 -1555 11140 -1535
rect 11100 -1585 11140 -1555
rect 11100 -1605 11110 -1585
rect 11130 -1605 11140 -1585
rect 11100 -1635 11140 -1605
rect 11100 -1655 11110 -1635
rect 11130 -1655 11140 -1635
rect 11100 -1685 11140 -1655
rect 11100 -1705 11110 -1685
rect 11130 -1705 11140 -1685
rect 11100 -1735 11140 -1705
rect 11100 -1755 11110 -1735
rect 11130 -1755 11140 -1735
rect 11100 -1770 11140 -1755
rect 11180 -1440 11220 -1425
rect 11180 -1460 11190 -1440
rect 11210 -1460 11220 -1440
rect 11180 -1490 11220 -1460
rect 11180 -1510 11190 -1490
rect 11210 -1510 11220 -1490
rect 11180 -1540 11220 -1510
rect 11180 -1560 11190 -1540
rect 11210 -1560 11220 -1540
rect 11180 -1590 11220 -1560
rect 11180 -1610 11190 -1590
rect 11210 -1610 11220 -1590
rect 11180 -1640 11220 -1610
rect 11180 -1660 11190 -1640
rect 11210 -1660 11220 -1640
rect 11180 -1690 11220 -1660
rect 11180 -1710 11190 -1690
rect 11210 -1710 11220 -1690
rect 11180 -1740 11220 -1710
rect 11180 -1760 11190 -1740
rect 11210 -1760 11220 -1740
rect 11180 -1790 11220 -1760
rect 11180 -1810 11190 -1790
rect 11210 -1810 11220 -1790
rect 11180 -1825 11220 -1810
rect 12580 -1440 12620 -1425
rect 12580 -1460 12590 -1440
rect 12610 -1460 12620 -1440
rect 12580 -1490 12620 -1460
rect 12580 -1510 12590 -1490
rect 12610 -1510 12620 -1490
rect 12580 -1540 12620 -1510
rect 12580 -1560 12590 -1540
rect 12610 -1560 12620 -1540
rect 12580 -1590 12620 -1560
rect 12580 -1610 12590 -1590
rect 12610 -1610 12620 -1590
rect 12580 -1640 12620 -1610
rect 12580 -1660 12590 -1640
rect 12610 -1660 12620 -1640
rect 12580 -1690 12620 -1660
rect 12580 -1710 12590 -1690
rect 12610 -1710 12620 -1690
rect 12580 -1740 12620 -1710
rect 12580 -1760 12590 -1740
rect 12610 -1760 12620 -1740
rect 12580 -1790 12620 -1760
rect 12580 -1810 12590 -1790
rect 12610 -1810 12620 -1790
rect 12580 -1825 12620 -1810
rect 12855 -2030 12895 -2015
rect 12855 -2050 12865 -2030
rect 12885 -2050 12895 -2030
rect 12855 -2080 12895 -2050
rect 12855 -2100 12865 -2080
rect 12885 -2100 12895 -2080
rect 11180 -2120 11220 -2105
rect 11180 -2140 11190 -2120
rect 11210 -2140 11220 -2120
rect 11180 -2170 11220 -2140
rect 11180 -2190 11190 -2170
rect 11210 -2190 11220 -2170
rect 11180 -2220 11220 -2190
rect 11180 -2240 11190 -2220
rect 11210 -2240 11220 -2220
rect 11180 -2270 11220 -2240
rect 11180 -2290 11190 -2270
rect 11210 -2290 11220 -2270
rect 11180 -2320 11220 -2290
rect 11180 -2340 11190 -2320
rect 11210 -2340 11220 -2320
rect 11180 -2370 11220 -2340
rect 11180 -2390 11190 -2370
rect 11210 -2390 11220 -2370
rect 11180 -2420 11220 -2390
rect 11180 -2440 11190 -2420
rect 11210 -2440 11220 -2420
rect 11180 -2470 11220 -2440
rect 11180 -2490 11190 -2470
rect 11210 -2490 11220 -2470
rect 11180 -2505 11220 -2490
rect 12580 -2120 12620 -2105
rect 12580 -2140 12590 -2120
rect 12610 -2140 12620 -2120
rect 12580 -2170 12620 -2140
rect 12580 -2190 12590 -2170
rect 12610 -2190 12620 -2170
rect 12580 -2220 12620 -2190
rect 12580 -2240 12590 -2220
rect 12610 -2240 12620 -2220
rect 12580 -2270 12620 -2240
rect 12580 -2290 12590 -2270
rect 12610 -2290 12620 -2270
rect 12580 -2320 12620 -2290
rect 12855 -2130 12895 -2100
rect 12855 -2150 12865 -2130
rect 12885 -2150 12895 -2130
rect 12855 -2180 12895 -2150
rect 12855 -2200 12865 -2180
rect 12885 -2200 12895 -2180
rect 12855 -2230 12895 -2200
rect 12855 -2250 12865 -2230
rect 12885 -2250 12895 -2230
rect 12855 -2280 12895 -2250
rect 12855 -2300 12865 -2280
rect 12885 -2300 12895 -2280
rect 12855 -2315 12895 -2300
rect 14145 -2030 14185 -2015
rect 14145 -2050 14155 -2030
rect 14175 -2050 14185 -2030
rect 14145 -2080 14185 -2050
rect 14145 -2100 14155 -2080
rect 14175 -2100 14185 -2080
rect 14145 -2130 14185 -2100
rect 14145 -2150 14155 -2130
rect 14175 -2150 14185 -2130
rect 14145 -2180 14185 -2150
rect 14145 -2200 14155 -2180
rect 14175 -2200 14185 -2180
rect 14145 -2230 14185 -2200
rect 14145 -2250 14155 -2230
rect 14175 -2250 14185 -2230
rect 14145 -2280 14185 -2250
rect 14145 -2300 14155 -2280
rect 14175 -2300 14185 -2280
rect 14145 -2315 14185 -2300
rect 12580 -2340 12590 -2320
rect 12610 -2340 12620 -2320
rect 12580 -2370 12620 -2340
rect 12580 -2390 12590 -2370
rect 12610 -2390 12620 -2370
rect 12580 -2420 12620 -2390
rect 12580 -2440 12590 -2420
rect 12610 -2440 12620 -2420
rect 12580 -2470 12620 -2440
rect 12580 -2490 12590 -2470
rect 12610 -2490 12620 -2470
rect 12580 -2505 12620 -2490
rect 12855 -2460 12895 -2445
rect 12855 -2480 12865 -2460
rect 12885 -2480 12895 -2460
rect 12855 -2510 12895 -2480
rect 12855 -2530 12865 -2510
rect 12885 -2530 12895 -2510
rect 12855 -2545 12895 -2530
rect 14145 -2460 14185 -2445
rect 14145 -2480 14155 -2460
rect 14175 -2480 14185 -2460
rect 14145 -2510 14185 -2480
rect 14145 -2530 14155 -2510
rect 14175 -2530 14185 -2510
rect 14145 -2545 14185 -2530
rect 12855 -2750 12895 -2735
rect 12855 -2770 12865 -2750
rect 12885 -2770 12895 -2750
rect 12855 -2800 12895 -2770
rect 12855 -2820 12865 -2800
rect 12885 -2820 12895 -2800
rect 12855 -2850 12895 -2820
rect 12855 -2870 12865 -2850
rect 12885 -2870 12895 -2850
rect 11235 -2885 11275 -2870
rect 11235 -2905 11245 -2885
rect 11265 -2905 11275 -2885
rect 11235 -2935 11275 -2905
rect 11235 -2955 11245 -2935
rect 11265 -2955 11275 -2935
rect 11235 -2985 11275 -2955
rect 11235 -3005 11245 -2985
rect 11265 -3005 11275 -2985
rect 11235 -3020 11275 -3005
rect 12525 -2885 12565 -2870
rect 12855 -2885 12895 -2870
rect 14145 -2750 14185 -2735
rect 14145 -2770 14155 -2750
rect 14175 -2770 14185 -2750
rect 14145 -2800 14185 -2770
rect 14145 -2820 14155 -2800
rect 14175 -2820 14185 -2800
rect 14145 -2850 14185 -2820
rect 14145 -2870 14155 -2850
rect 14175 -2870 14185 -2850
rect 14145 -2885 14185 -2870
rect 12525 -2905 12535 -2885
rect 12555 -2905 12565 -2885
rect 12525 -2935 12565 -2905
rect 12525 -2955 12535 -2935
rect 12555 -2955 12565 -2935
rect 12525 -2985 12565 -2955
rect 12525 -3005 12535 -2985
rect 12555 -3005 12565 -2985
rect 12525 -3020 12565 -3005
rect 12855 -3030 12895 -3015
rect 12855 -3050 12865 -3030
rect 12885 -3050 12895 -3030
rect 12855 -3075 12895 -3050
rect 12855 -3095 12865 -3075
rect 12885 -3095 12895 -3075
rect 12855 -3120 12895 -3095
rect 12855 -3140 12865 -3120
rect 12885 -3140 12895 -3120
rect 12855 -3170 12895 -3140
rect 12855 -3190 12865 -3170
rect 12885 -3190 12895 -3170
rect 12855 -3215 12895 -3190
rect 12855 -3235 12865 -3215
rect 12885 -3235 12895 -3215
rect 12855 -3260 12895 -3235
rect 12855 -3280 12865 -3260
rect 12885 -3280 12895 -3260
rect 12855 -3295 12895 -3280
rect 14135 -3030 14175 -3015
rect 14135 -3050 14145 -3030
rect 14165 -3050 14175 -3030
rect 14135 -3075 14175 -3050
rect 14135 -3095 14145 -3075
rect 14165 -3095 14175 -3075
rect 14135 -3120 14175 -3095
rect 14135 -3140 14145 -3120
rect 14165 -3140 14175 -3120
rect 14135 -3170 14175 -3140
rect 14135 -3190 14145 -3170
rect 14165 -3190 14175 -3170
rect 14135 -3215 14175 -3190
rect 14135 -3235 14145 -3215
rect 14165 -3235 14175 -3215
rect 14135 -3260 14175 -3235
rect 14135 -3280 14145 -3260
rect 14165 -3280 14175 -3260
rect 14135 -3295 14175 -3280
rect 10990 -3350 11030 -3335
rect 10990 -3370 11000 -3350
rect 11020 -3370 11030 -3350
rect 10990 -3400 11030 -3370
rect 10990 -3420 11000 -3400
rect 11020 -3420 11030 -3400
rect 10990 -3450 11030 -3420
rect 10990 -3470 11000 -3450
rect 11020 -3470 11030 -3450
rect 10990 -3485 11030 -3470
rect 11730 -3350 11770 -3335
rect 11730 -3370 11740 -3350
rect 11760 -3370 11770 -3350
rect 11730 -3400 11770 -3370
rect 11730 -3420 11740 -3400
rect 11760 -3420 11770 -3400
rect 11730 -3450 11770 -3420
rect 11730 -3470 11740 -3450
rect 11760 -3470 11770 -3450
rect 11730 -3485 11770 -3470
rect 12030 -3350 12070 -3335
rect 12030 -3370 12040 -3350
rect 12060 -3370 12070 -3350
rect 12030 -3400 12070 -3370
rect 12030 -3420 12040 -3400
rect 12060 -3420 12070 -3400
rect 12030 -3450 12070 -3420
rect 12030 -3470 12040 -3450
rect 12060 -3470 12070 -3450
rect 12030 -3485 12070 -3470
rect 12770 -3350 12810 -3335
rect 12770 -3370 12780 -3350
rect 12800 -3370 12810 -3350
rect 12770 -3400 12810 -3370
rect 12770 -3420 12780 -3400
rect 12800 -3420 12810 -3400
rect 12770 -3450 12810 -3420
rect 12770 -3470 12780 -3450
rect 12800 -3470 12810 -3450
rect 12770 -3485 12810 -3470
rect 11165 -3830 11205 -3815
rect 11165 -3850 11175 -3830
rect 11195 -3850 11205 -3830
rect 11165 -3880 11205 -3850
rect 11165 -3900 11175 -3880
rect 11195 -3900 11205 -3880
rect 11165 -3930 11205 -3900
rect 11165 -3950 11175 -3930
rect 11195 -3950 11205 -3930
rect 11165 -3980 11205 -3950
rect 11165 -4000 11175 -3980
rect 11195 -4000 11205 -3980
rect 11165 -4030 11205 -4000
rect 11165 -4050 11175 -4030
rect 11195 -4050 11205 -4030
rect 11165 -4065 11205 -4050
rect 12620 -3830 12660 -3815
rect 12620 -3850 12630 -3830
rect 12650 -3850 12660 -3830
rect 12620 -3880 12660 -3850
rect 12620 -3900 12630 -3880
rect 12650 -3900 12660 -3880
rect 12620 -3930 12660 -3900
rect 12620 -3950 12630 -3930
rect 12650 -3950 12660 -3930
rect 12620 -3980 12660 -3950
rect 12620 -4000 12630 -3980
rect 12650 -4000 12660 -3980
rect 12620 -4030 12660 -4000
rect 12620 -4050 12630 -4030
rect 12650 -4050 12660 -4030
rect 12620 -4065 12660 -4050
<< nsubdiff >>
rect 2955 2915 2995 2930
rect 2955 2895 2965 2915
rect 2985 2895 2995 2915
rect 2955 2865 2995 2895
rect 2955 2845 2965 2865
rect 2985 2845 2995 2865
rect 2955 2830 2995 2845
rect 5015 2915 5055 2930
rect 5015 2895 5025 2915
rect 5045 2895 5055 2915
rect 5015 2865 5055 2895
rect 5015 2845 5025 2865
rect 5045 2845 5055 2865
rect 5015 2830 5055 2845
rect 3135 2685 3175 2700
rect 3135 2665 3145 2685
rect 3165 2665 3175 2685
rect 3135 2635 3175 2665
rect 3135 2615 3145 2635
rect 3165 2615 3175 2635
rect 3135 2585 3175 2615
rect 3135 2565 3145 2585
rect 3165 2565 3175 2585
rect 3135 2535 3175 2565
rect 3135 2515 3145 2535
rect 3165 2515 3175 2535
rect 3135 2485 3175 2515
rect 3135 2465 3145 2485
rect 3165 2465 3175 2485
rect 3135 2435 3175 2465
rect 3135 2415 3145 2435
rect 3165 2415 3175 2435
rect 3135 2400 3175 2415
rect 4835 2685 4875 2700
rect 4835 2665 4845 2685
rect 4865 2665 4875 2685
rect 4835 2635 4875 2665
rect 4835 2615 4845 2635
rect 4865 2615 4875 2635
rect 4835 2585 4875 2615
rect 4835 2565 4845 2585
rect 4865 2565 4875 2585
rect 4835 2535 4875 2565
rect 4835 2515 4845 2535
rect 4865 2515 4875 2535
rect 4835 2485 4875 2515
rect 4835 2465 4845 2485
rect 4865 2465 4875 2485
rect 4835 2435 4875 2465
rect 4835 2415 4845 2435
rect 4865 2415 4875 2435
rect 4835 2400 4875 2415
rect 3985 1985 4025 2000
rect 3985 1965 3995 1985
rect 4015 1965 4025 1985
rect 3985 1935 4025 1965
rect 3985 1915 3995 1935
rect 4015 1915 4025 1935
rect 3985 1900 4025 1915
<< psubdiffcont >>
rect 11210 8895 11230 8915
rect 11470 8895 11490 8915
rect 11540 8910 11560 8930
rect 11980 8910 12000 8930
rect 12050 8895 12070 8915
rect 12610 8895 12630 8915
rect 10790 8495 10810 8515
rect 10790 8445 10810 8465
rect 10790 8395 10810 8415
rect 10790 8345 10810 8365
rect 10790 8295 10810 8315
rect 10460 8245 10480 8265
rect 10720 8245 10740 8265
rect 10790 8245 10810 8265
rect 11110 8545 11130 8565
rect 11110 8495 11130 8515
rect 11110 8445 11130 8465
rect 11110 8395 11130 8415
rect 11110 8345 11130 8365
rect 11110 8295 11130 8315
rect 11110 8245 11130 8265
rect 11190 8540 11210 8560
rect 11190 8490 11210 8510
rect 11190 8440 11210 8460
rect 11190 8390 11210 8410
rect 11190 8340 11210 8360
rect 11190 8290 11210 8310
rect 11190 8240 11210 8260
rect 11190 8190 11210 8210
rect 12590 8540 12610 8560
rect 12590 8490 12610 8510
rect 12590 8440 12610 8460
rect 12590 8390 12610 8410
rect 12590 8340 12610 8360
rect 18290 8495 18310 8515
rect 18290 8445 18310 8465
rect 18290 8395 18310 8415
rect 12590 8290 12610 8310
rect 18290 8345 18310 8365
rect 18290 8295 18310 8315
rect 12590 8240 12610 8260
rect 17960 8245 17980 8265
rect 12590 8190 12610 8210
rect 12865 8205 12885 8225
rect 12865 8155 12885 8175
rect 12865 8105 12885 8125
rect 12865 8055 12885 8075
rect 12865 8005 12885 8025
rect 12865 7955 12885 7975
rect 18220 8245 18240 8265
rect 18290 8245 18310 8265
rect 18610 8545 18630 8565
rect 18610 8495 18630 8515
rect 18610 8445 18630 8465
rect 18610 8395 18630 8415
rect 18610 8345 18630 8365
rect 18610 8295 18630 8315
rect 18610 8245 18630 8265
rect 18690 8540 18710 8560
rect 18690 8490 18710 8510
rect 18690 8440 18710 8460
rect 18690 8390 18710 8410
rect 18690 8340 18710 8360
rect 18690 8290 18710 8310
rect 18690 8240 18710 8260
rect 14155 8205 14175 8225
rect 18690 8190 18710 8210
rect 20090 8540 20110 8560
rect 20090 8490 20110 8510
rect 20090 8440 20110 8460
rect 20090 8390 20110 8410
rect 20090 8340 20110 8360
rect 20090 8290 20110 8310
rect 20090 8240 20110 8260
rect 20090 8190 20110 8210
rect 20360 8205 20380 8225
rect 14155 8155 14175 8175
rect 20360 8155 20380 8175
rect 14155 8105 14175 8125
rect 14155 8055 14175 8075
rect 14155 8005 14175 8025
rect 14155 7955 14175 7975
rect 20360 8105 20380 8125
rect 20360 8055 20380 8075
rect 20360 8005 20380 8025
rect 20360 7955 20380 7975
rect 11190 7860 11210 7880
rect 11190 7810 11210 7830
rect 11190 7760 11210 7780
rect 11190 7710 11210 7730
rect 11190 7660 11210 7680
rect 9650 7585 9670 7605
rect 9650 7535 9670 7555
rect 10940 7585 10960 7605
rect 10940 7535 10960 7555
rect 11190 7610 11210 7630
rect 11190 7560 11210 7580
rect 11190 7510 11210 7530
rect 21650 8205 21670 8225
rect 21650 8155 21670 8175
rect 21650 8105 21670 8125
rect 21650 8055 21670 8075
rect 21650 8005 21670 8025
rect 21650 7955 21670 7975
rect 12590 7860 12610 7880
rect 18690 7860 18710 7880
rect 12590 7810 12610 7830
rect 12590 7760 12610 7780
rect 12590 7710 12610 7730
rect 18690 7810 18710 7830
rect 18690 7760 18710 7780
rect 18690 7710 18710 7730
rect 12590 7660 12610 7680
rect 18690 7660 18710 7680
rect 12590 7610 12610 7630
rect 12590 7560 12610 7580
rect 12590 7510 12610 7530
rect 12865 7585 12885 7605
rect 12865 7535 12885 7555
rect 14155 7585 14175 7605
rect 14155 7535 14175 7555
rect 17150 7585 17170 7605
rect 17150 7535 17170 7555
rect 18440 7585 18460 7605
rect 18440 7535 18460 7555
rect 18690 7610 18710 7630
rect 18690 7560 18710 7580
rect 18690 7510 18710 7530
rect 20090 7860 20110 7880
rect 20090 7810 20110 7830
rect 20090 7760 20110 7780
rect 20090 7710 20110 7730
rect 20090 7660 20110 7680
rect 20090 7610 20110 7630
rect 20090 7560 20110 7580
rect 20090 7510 20110 7530
rect 20360 7585 20380 7605
rect 20360 7535 20380 7555
rect 21650 7585 21670 7605
rect 21650 7535 21670 7555
rect 9650 7135 9670 7155
rect 9650 7085 9670 7105
rect 9650 7035 9670 7055
rect 10940 7135 10960 7155
rect 12865 7135 12885 7155
rect 10940 7085 10960 7105
rect 10940 7035 10960 7055
rect 11245 7095 11265 7115
rect 11245 7045 11265 7065
rect 11245 6995 11265 7015
rect 12535 7095 12555 7115
rect 12535 7045 12555 7065
rect 12865 7085 12885 7105
rect 12865 7035 12885 7055
rect 14155 7135 14175 7155
rect 14155 7085 14175 7105
rect 14155 7035 14175 7055
rect 17150 7135 17170 7155
rect 17150 7085 17170 7105
rect 17150 7035 17170 7055
rect 18440 7135 18460 7155
rect 20360 7135 20380 7155
rect 18440 7085 18460 7105
rect 18440 7035 18460 7055
rect 18745 7095 18765 7115
rect 18745 7045 18765 7065
rect 12535 6995 12555 7015
rect 18745 6995 18765 7015
rect 20035 7095 20055 7115
rect 20035 7045 20055 7065
rect 20360 7085 20380 7105
rect 20360 7035 20380 7055
rect 21650 7135 21670 7155
rect 21650 7085 21670 7105
rect 21650 7035 21670 7055
rect 20035 6995 20055 7015
rect 20460 6820 20480 6840
rect 20460 6770 20480 6790
rect 20460 6720 20480 6740
rect 20870 6820 20890 6840
rect 20870 6770 20890 6790
rect 20870 6720 20890 6740
rect 11000 6630 11020 6650
rect 11000 6580 11020 6600
rect 11000 6530 11020 6550
rect 11740 6630 11760 6650
rect 11740 6580 11760 6600
rect 11740 6530 11760 6550
rect 12040 6630 12060 6650
rect 12040 6580 12060 6600
rect 12040 6530 12060 6550
rect 12780 6630 12800 6650
rect 12780 6580 12800 6600
rect 12780 6530 12800 6550
rect 18500 6630 18520 6650
rect 18500 6580 18520 6600
rect 18500 6530 18520 6550
rect 19240 6630 19260 6650
rect 19240 6580 19260 6600
rect 19240 6530 19260 6550
rect 19540 6630 19560 6650
rect 19540 6580 19560 6600
rect 19540 6530 19560 6550
rect 20280 6630 20300 6650
rect 20280 6580 20300 6600
rect 20280 6530 20300 6550
rect 20365 6485 20385 6505
rect 20365 6435 20385 6455
rect 20365 6385 20385 6405
rect 20665 6485 20685 6505
rect 20665 6435 20685 6455
rect 20665 6385 20685 6405
rect 20965 6485 20985 6505
rect 20965 6435 20985 6455
rect 20965 6385 20985 6405
rect 9635 6250 9655 6270
rect 9635 6205 9655 6225
rect 9635 6160 9655 6180
rect 9635 6110 9655 6130
rect 9635 6065 9655 6085
rect 9635 6020 9655 6040
rect 10915 6250 10935 6270
rect 10915 6205 10935 6225
rect 12865 6250 12885 6270
rect 12865 6205 12885 6225
rect 10915 6160 10935 6180
rect 10915 6110 10935 6130
rect 10915 6065 10935 6085
rect 10915 6020 10935 6040
rect 11175 6150 11195 6170
rect 11175 6100 11195 6120
rect 11175 6050 11195 6070
rect 11175 6000 11195 6020
rect 11175 5950 11195 5970
rect 12630 6150 12650 6170
rect 12630 6100 12650 6120
rect 12630 6050 12650 6070
rect 12630 6000 12650 6020
rect 12865 6160 12885 6180
rect 12865 6110 12885 6130
rect 12865 6065 12885 6085
rect 12865 6020 12885 6040
rect 14145 6250 14165 6270
rect 14145 6205 14165 6225
rect 14145 6160 14165 6180
rect 14145 6110 14165 6130
rect 14145 6065 14165 6085
rect 14145 6020 14165 6040
rect 18675 6190 18695 6210
rect 18675 6140 18695 6160
rect 18675 6090 18695 6110
rect 18675 6040 18695 6060
rect 12630 5950 12650 5970
rect 18675 5990 18695 6010
rect 20130 6190 20150 6210
rect 20130 6140 20150 6160
rect 20130 6090 20150 6110
rect 20130 6040 20150 6060
rect 20515 6145 20535 6165
rect 20515 6095 20535 6115
rect 20515 6045 20535 6065
rect 20815 6145 20835 6165
rect 20815 6095 20835 6115
rect 20815 6045 20835 6065
rect 20130 5990 20150 6010
rect 11210 4355 11230 4375
rect 11470 4355 11490 4375
rect 11540 4370 11560 4390
rect 11980 4370 12000 4390
rect 12050 4355 12070 4375
rect 12610 4355 12630 4375
rect 11220 4120 11240 4140
rect 12510 4120 12530 4140
rect 11165 3815 11185 3835
rect 11905 3815 11925 3835
rect 12645 3815 12665 3835
rect 10125 3550 10145 3570
rect 10125 3500 10145 3520
rect 10125 3450 10145 3470
rect 10125 3400 10145 3420
rect 10125 3350 10145 3370
rect 10125 3300 10145 3320
rect 10125 3250 10145 3270
rect 10125 3200 10145 3220
rect 10125 3150 10145 3170
rect 10125 3100 10145 3120
rect 10125 3050 10145 3070
rect 10125 3000 10145 3020
rect 10865 3550 10885 3570
rect 10865 3500 10885 3520
rect 10865 3450 10885 3470
rect 10865 3400 10885 3420
rect 10865 3350 10885 3370
rect 10865 3300 10885 3320
rect 10865 3250 10885 3270
rect 10865 3200 10885 3220
rect 11190 3540 11210 3560
rect 11190 3490 11210 3510
rect 11190 3440 11210 3460
rect 11190 3390 11210 3410
rect 11190 3340 11210 3360
rect 11190 3290 11210 3310
rect 11190 3240 11210 3260
rect 11190 3190 11210 3210
rect 12590 3540 12610 3560
rect 12590 3490 12610 3510
rect 12590 3440 12610 3460
rect 12590 3390 12610 3410
rect 12590 3340 12610 3360
rect 12590 3290 12610 3310
rect 12590 3240 12610 3260
rect 12590 3190 12610 3210
rect 12915 3550 12935 3570
rect 12915 3500 12935 3520
rect 12915 3450 12935 3470
rect 12915 3400 12935 3420
rect 12915 3350 12935 3370
rect 12915 3300 12935 3320
rect 12915 3250 12935 3270
rect 12915 3200 12935 3220
rect 10865 3150 10885 3170
rect 12915 3150 12935 3170
rect 10865 3100 10885 3120
rect 10865 3050 10885 3070
rect 10865 3000 10885 3020
rect 12915 3100 12935 3120
rect 12915 3050 12935 3070
rect 12915 3000 12935 3020
rect 13655 3550 13675 3570
rect 13655 3500 13675 3520
rect 13655 3450 13675 3470
rect 13655 3400 13675 3420
rect 13655 3350 13675 3370
rect 13655 3300 13675 3320
rect 13655 3250 13675 3270
rect 13655 3200 13675 3220
rect 13655 3150 13675 3170
rect 13655 3100 13675 3120
rect 13655 3050 13675 3070
rect 13655 3000 13675 3020
rect 25790 3495 25810 3515
rect 25790 3445 25810 3465
rect 25790 3395 25810 3415
rect 25790 3345 25810 3365
rect 25790 3295 25810 3315
rect 25460 3245 25480 3265
rect 25720 3245 25740 3265
rect 25790 3245 25810 3265
rect 26110 3545 26130 3565
rect 26110 3495 26130 3515
rect 26110 3445 26130 3465
rect 26110 3395 26130 3415
rect 26110 3345 26130 3365
rect 26110 3295 26130 3315
rect 26110 3245 26130 3265
rect 26190 3540 26210 3560
rect 26190 3490 26210 3510
rect 26190 3440 26210 3460
rect 26190 3390 26210 3410
rect 26190 3340 26210 3360
rect 26190 3290 26210 3310
rect 26190 3240 26210 3260
rect 26190 3190 26210 3210
rect 27590 3540 27610 3560
rect 27590 3490 27610 3510
rect 27590 3440 27610 3460
rect 27590 3390 27610 3410
rect 27590 3340 27610 3360
rect 27590 3290 27610 3310
rect 27590 3240 27610 3260
rect 27590 3190 27610 3210
rect 27860 3205 27880 3225
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 27860 3155 27880 3175
rect 27860 3105 27880 3125
rect 27860 3055 27880 3075
rect 27860 3005 27880 3025
rect 27860 2955 27880 2975
rect 29150 3205 29170 3225
rect 29150 3155 29170 3175
rect 29150 3105 29170 3125
rect 29150 3055 29170 3075
rect 29150 3005 29170 3025
rect 29150 2955 29170 2975
rect 11190 2860 11210 2880
rect 11190 2810 11210 2830
rect 11190 2760 11210 2780
rect 11190 2710 11210 2730
rect 11190 2660 11210 2680
rect 10125 2620 10145 2640
rect 10125 2570 10145 2590
rect 10125 2520 10145 2540
rect 10125 2470 10145 2490
rect 10865 2620 10885 2640
rect 10865 2570 10885 2590
rect 10865 2520 10885 2540
rect 11190 2610 11210 2630
rect 11190 2560 11210 2580
rect 11190 2510 11210 2530
rect 12590 2860 12610 2880
rect 12590 2810 12610 2830
rect 12590 2760 12610 2780
rect 12590 2710 12610 2730
rect 12590 2660 12610 2680
rect 26190 2860 26210 2880
rect 26190 2810 26210 2830
rect 26190 2760 26210 2780
rect 26190 2710 26210 2730
rect 26190 2660 26210 2680
rect 12590 2610 12610 2630
rect 12590 2560 12610 2580
rect 12590 2510 12610 2530
rect 12915 2620 12935 2640
rect 12915 2570 12935 2590
rect 12915 2520 12935 2540
rect 10865 2470 10885 2490
rect 12915 2470 12935 2490
rect 13655 2620 13675 2640
rect 13655 2570 13675 2590
rect 13655 2520 13675 2540
rect 13655 2470 13675 2490
rect 10125 2230 10145 2250
rect 10125 2180 10145 2200
rect 10125 2130 10145 2150
rect 10125 2080 10145 2100
rect 10125 2030 10145 2050
rect 10125 1980 10145 2000
rect 10865 2230 10885 2250
rect 10865 2180 10885 2200
rect 12915 2230 12935 2250
rect 12915 2180 12935 2200
rect 10865 2130 10885 2150
rect 12915 2130 12935 2150
rect 10865 2080 10885 2100
rect 10865 2030 10885 2050
rect 10865 1980 10885 2000
rect 11245 2095 11265 2115
rect 11245 2045 11265 2065
rect 11245 1995 11265 2015
rect 12535 2095 12555 2115
rect 12535 2045 12555 2065
rect 12535 1995 12555 2015
rect 12915 2080 12935 2100
rect 12915 2030 12935 2050
rect 12915 1980 12935 2000
rect 13655 2230 13675 2250
rect 13655 2180 13675 2200
rect 13655 2130 13675 2150
rect 13655 2080 13675 2100
rect 13655 2030 13675 2050
rect 24650 2585 24670 2605
rect 24650 2535 24670 2555
rect 25940 2585 25960 2605
rect 25940 2535 25960 2555
rect 26190 2610 26210 2630
rect 26190 2560 26210 2580
rect 26190 2510 26210 2530
rect 27590 2860 27610 2880
rect 27590 2810 27610 2830
rect 27590 2760 27610 2780
rect 27590 2710 27610 2730
rect 27590 2660 27610 2680
rect 27590 2610 27610 2630
rect 27590 2560 27610 2580
rect 27590 2510 27610 2530
rect 27860 2585 27880 2605
rect 27860 2535 27880 2555
rect 29150 2585 29170 2605
rect 29150 2535 29170 2555
rect 24650 2135 24670 2155
rect 24650 2085 24670 2105
rect 24650 2035 24670 2055
rect 25940 2135 25960 2155
rect 27860 2135 27880 2155
rect 25940 2085 25960 2105
rect 25940 2035 25960 2055
rect 26245 2095 26265 2115
rect 26245 2045 26265 2065
rect 13655 1980 13675 2000
rect 26245 1995 26265 2015
rect 27535 2095 27555 2115
rect 27535 2045 27555 2065
rect 27860 2085 27880 2105
rect 27860 2035 27880 2055
rect 29150 2135 29170 2155
rect 29150 2085 29170 2105
rect 29150 2035 29170 2055
rect 27535 1995 27555 2015
rect 27960 1820 27980 1840
rect 27960 1770 27980 1790
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 27960 1720 27980 1740
rect 28370 1820 28390 1840
rect 28370 1770 28390 1790
rect 28370 1720 28390 1740
rect 3995 1630 4015 1650
rect 10125 1620 10145 1640
rect 5075 1040 5095 1060
rect 5075 990 5095 1010
rect 10125 1570 10145 1590
rect 10125 1520 10145 1540
rect 10125 1470 10145 1490
rect 10125 1420 10145 1440
rect 10125 1370 10145 1390
rect 10125 1320 10145 1340
rect 10125 1270 10145 1290
rect 10125 1220 10145 1240
rect 10125 1170 10145 1190
rect 10125 1120 10145 1140
rect 10125 1070 10145 1090
rect 10125 1020 10145 1040
rect 10125 970 10145 990
rect 10805 1620 10825 1640
rect 10805 1570 10825 1590
rect 10805 1520 10825 1540
rect 11000 1630 11020 1650
rect 11000 1580 11020 1600
rect 11000 1530 11020 1550
rect 11740 1630 11760 1650
rect 11740 1580 11760 1600
rect 11740 1530 11760 1550
rect 12040 1630 12060 1650
rect 12040 1580 12060 1600
rect 12040 1530 12060 1550
rect 12780 1630 12800 1650
rect 12780 1580 12800 1600
rect 12780 1530 12800 1550
rect 12975 1620 12995 1640
rect 12975 1570 12995 1590
rect 12975 1520 12995 1540
rect 10805 1470 10825 1490
rect 12975 1470 12995 1490
rect 10805 1420 10825 1440
rect 10805 1370 10825 1390
rect 10805 1320 10825 1340
rect 10805 1270 10825 1290
rect 12975 1420 12995 1440
rect 12975 1370 12995 1390
rect 12975 1320 12995 1340
rect 12975 1270 12995 1290
rect 10805 1220 10825 1240
rect 10805 1170 10825 1190
rect 12975 1220 12995 1240
rect 10805 1120 10825 1140
rect 10805 1070 10825 1090
rect 10805 1020 10825 1040
rect 10805 970 10825 990
rect 11175 1150 11195 1170
rect 11175 1100 11195 1120
rect 11175 1050 11195 1070
rect 11175 1000 11195 1020
rect 11175 950 11195 970
rect 12630 1150 12650 1170
rect 12630 1100 12650 1120
rect 12630 1050 12650 1070
rect 12630 1000 12650 1020
rect 12630 950 12650 970
rect 12975 1170 12995 1190
rect 12975 1120 12995 1140
rect 12975 1070 12995 1090
rect 12975 1020 12995 1040
rect 12975 970 12995 990
rect 13655 1620 13675 1640
rect 26000 1630 26020 1650
rect 13655 1570 13675 1590
rect 13655 1520 13675 1540
rect 13655 1470 13675 1490
rect 13655 1420 13675 1440
rect 13655 1370 13675 1390
rect 13655 1320 13675 1340
rect 13655 1270 13675 1290
rect 13655 1220 13675 1240
rect 13655 1170 13675 1190
rect 13655 1120 13675 1140
rect 13655 1070 13675 1090
rect 13655 1020 13675 1040
rect 13655 970 13675 990
rect 26000 1580 26020 1600
rect 26000 1530 26020 1550
rect 26740 1630 26760 1650
rect 26740 1580 26760 1600
rect 26740 1530 26760 1550
rect 27040 1630 27060 1650
rect 27040 1580 27060 1600
rect 27040 1530 27060 1550
rect 27780 1630 27800 1650
rect 27780 1580 27800 1600
rect 27780 1530 27800 1550
rect 27865 1485 27885 1505
rect 27865 1435 27885 1455
rect 27865 1385 27885 1405
rect 28165 1485 28185 1505
rect 28165 1435 28185 1455
rect 28165 1385 28185 1405
rect 28465 1485 28485 1505
rect 28465 1435 28485 1455
rect 28465 1385 28485 1405
rect 26175 1190 26195 1210
rect 26175 1140 26195 1160
rect 26175 1090 26195 1110
rect 26175 1040 26195 1060
rect 26175 990 26195 1010
rect 27630 1190 27650 1210
rect 27630 1140 27650 1160
rect 27630 1090 27650 1110
rect 27630 1040 27650 1060
rect 28015 1145 28035 1165
rect 28015 1095 28035 1115
rect 28015 1045 28035 1065
rect 28315 1145 28335 1165
rect 28315 1095 28335 1115
rect 28315 1045 28335 1065
rect 27630 990 27650 1010
rect 2965 845 2985 865
rect 2965 795 2985 815
rect 5025 845 5045 865
rect 5025 795 5045 815
rect 11850 715 11870 735
rect 12590 715 12610 735
rect 10790 -1505 10810 -1485
rect 10790 -1555 10810 -1535
rect 10790 -1605 10810 -1585
rect 10790 -1655 10810 -1635
rect 10790 -1705 10810 -1685
rect 10460 -1755 10480 -1735
rect 10720 -1755 10740 -1735
rect 10790 -1755 10810 -1735
rect 11110 -1455 11130 -1435
rect 11110 -1505 11130 -1485
rect 11110 -1555 11130 -1535
rect 11110 -1605 11130 -1585
rect 11110 -1655 11130 -1635
rect 11110 -1705 11130 -1685
rect 11110 -1755 11130 -1735
rect 11190 -1460 11210 -1440
rect 11190 -1510 11210 -1490
rect 11190 -1560 11210 -1540
rect 11190 -1610 11210 -1590
rect 11190 -1660 11210 -1640
rect 11190 -1710 11210 -1690
rect 11190 -1760 11210 -1740
rect 11190 -1810 11210 -1790
rect 12590 -1460 12610 -1440
rect 12590 -1510 12610 -1490
rect 12590 -1560 12610 -1540
rect 12590 -1610 12610 -1590
rect 12590 -1660 12610 -1640
rect 12590 -1710 12610 -1690
rect 12590 -1760 12610 -1740
rect 12590 -1810 12610 -1790
rect 12865 -2050 12885 -2030
rect 12865 -2100 12885 -2080
rect 11190 -2140 11210 -2120
rect 11190 -2190 11210 -2170
rect 11190 -2240 11210 -2220
rect 11190 -2290 11210 -2270
rect 11190 -2340 11210 -2320
rect 11190 -2390 11210 -2370
rect 11190 -2440 11210 -2420
rect 11190 -2490 11210 -2470
rect 12590 -2140 12610 -2120
rect 12590 -2190 12610 -2170
rect 12590 -2240 12610 -2220
rect 12590 -2290 12610 -2270
rect 12865 -2150 12885 -2130
rect 12865 -2200 12885 -2180
rect 12865 -2250 12885 -2230
rect 12865 -2300 12885 -2280
rect 14155 -2050 14175 -2030
rect 14155 -2100 14175 -2080
rect 14155 -2150 14175 -2130
rect 14155 -2200 14175 -2180
rect 14155 -2250 14175 -2230
rect 14155 -2300 14175 -2280
rect 12590 -2340 12610 -2320
rect 12590 -2390 12610 -2370
rect 12590 -2440 12610 -2420
rect 12590 -2490 12610 -2470
rect 12865 -2480 12885 -2460
rect 12865 -2530 12885 -2510
rect 14155 -2480 14175 -2460
rect 14155 -2530 14175 -2510
rect 12865 -2770 12885 -2750
rect 12865 -2820 12885 -2800
rect 12865 -2870 12885 -2850
rect 11245 -2905 11265 -2885
rect 11245 -2955 11265 -2935
rect 11245 -3005 11265 -2985
rect 14155 -2770 14175 -2750
rect 14155 -2820 14175 -2800
rect 14155 -2870 14175 -2850
rect 12535 -2905 12555 -2885
rect 12535 -2955 12555 -2935
rect 12535 -3005 12555 -2985
rect 12865 -3050 12885 -3030
rect 12865 -3095 12885 -3075
rect 12865 -3140 12885 -3120
rect 12865 -3190 12885 -3170
rect 12865 -3235 12885 -3215
rect 12865 -3280 12885 -3260
rect 14145 -3050 14165 -3030
rect 14145 -3095 14165 -3075
rect 14145 -3140 14165 -3120
rect 14145 -3190 14165 -3170
rect 14145 -3235 14165 -3215
rect 14145 -3280 14165 -3260
rect 11000 -3370 11020 -3350
rect 11000 -3420 11020 -3400
rect 11000 -3470 11020 -3450
rect 11740 -3370 11760 -3350
rect 11740 -3420 11760 -3400
rect 11740 -3470 11760 -3450
rect 12040 -3370 12060 -3350
rect 12040 -3420 12060 -3400
rect 12040 -3470 12060 -3450
rect 12780 -3370 12800 -3350
rect 12780 -3420 12800 -3400
rect 12780 -3470 12800 -3450
rect 11175 -3850 11195 -3830
rect 11175 -3900 11195 -3880
rect 11175 -3950 11195 -3930
rect 11175 -4000 11195 -3980
rect 11175 -4050 11195 -4030
rect 12630 -3850 12650 -3830
rect 12630 -3900 12650 -3880
rect 12630 -3950 12650 -3930
rect 12630 -4000 12650 -3980
rect 12630 -4050 12650 -4030
<< nsubdiffcont >>
rect 2965 2895 2985 2915
rect 2965 2845 2985 2865
rect 5025 2895 5045 2915
rect 5025 2845 5045 2865
rect 3145 2665 3165 2685
rect 3145 2615 3165 2635
rect 3145 2565 3165 2585
rect 3145 2515 3165 2535
rect 3145 2465 3165 2485
rect 3145 2415 3165 2435
rect 4845 2665 4865 2685
rect 4845 2615 4865 2635
rect 4845 2565 4865 2585
rect 4845 2515 4865 2535
rect 4845 2465 4865 2485
rect 4845 2415 4865 2435
rect 3995 1965 4015 1985
rect 3995 1915 4015 1935
<< poly >>
rect 11632 9050 11668 9060
rect 11632 9030 11640 9050
rect 11660 9030 11668 9050
rect 11632 9020 11668 9030
rect 11752 9050 11788 9060
rect 11752 9030 11760 9050
rect 11780 9030 11788 9050
rect 11752 9020 11788 9030
rect 11872 9050 11908 9060
rect 11872 9030 11880 9050
rect 11900 9030 11908 9050
rect 11872 9020 11908 9030
rect 11570 9005 11610 9015
rect 11200 8990 11240 9000
rect 11200 8970 11210 8990
rect 11230 8970 11240 8990
rect 11460 8990 11500 9000
rect 11460 8970 11470 8990
rect 11490 8970 11500 8990
rect 11570 8985 11580 9005
rect 11600 8990 11610 9005
rect 11930 9005 11970 9015
rect 11930 8990 11940 9005
rect 11600 8985 11630 8990
rect 11570 8975 11630 8985
rect 11910 8985 11940 8990
rect 11960 8985 11970 9005
rect 11910 8975 11970 8985
rect 11200 8955 11300 8970
rect 11280 8943 11300 8955
rect 11340 8943 11360 8958
rect 11400 8955 11500 8970
rect 11610 8960 11630 8975
rect 11670 8960 11690 8975
rect 11730 8960 11750 8975
rect 11790 8960 11810 8975
rect 11850 8960 11870 8975
rect 11910 8960 11930 8975
rect 11400 8943 11420 8955
rect 12120 8935 12140 8950
rect 12180 8935 12200 8950
rect 12240 8935 12260 8950
rect 12300 8935 12320 8950
rect 12360 8935 12380 8950
rect 12420 8935 12440 8950
rect 12480 8935 12500 8950
rect 12540 8935 12560 8950
rect 11280 8865 11300 8880
rect 11340 8865 11360 8880
rect 11400 8865 11420 8880
rect 11610 8865 11630 8880
rect 11670 8870 11690 8880
rect 11730 8870 11750 8880
rect 11790 8870 11810 8880
rect 11850 8870 11870 8880
rect 11330 8855 11370 8865
rect 11670 8855 11870 8870
rect 11910 8865 11930 8880
rect 12120 8865 12140 8875
rect 12180 8865 12200 8875
rect 12240 8865 12260 8875
rect 12300 8865 12320 8875
rect 12360 8865 12380 8875
rect 12420 8865 12440 8875
rect 12480 8865 12500 8875
rect 12540 8865 12560 8875
rect 11330 8835 11340 8855
rect 11360 8835 11370 8855
rect 11330 8825 11370 8835
rect 11750 8850 11790 8855
rect 12120 8850 12560 8865
rect 11750 8830 11760 8850
rect 11780 8830 11790 8850
rect 11750 8820 11790 8830
rect 12203 8830 12211 8850
rect 12229 8830 12237 8850
rect 12203 8820 12237 8830
rect 11180 8620 11220 8630
rect 10905 8605 10945 8615
rect 10905 8585 10915 8605
rect 10935 8585 10945 8605
rect 11180 8600 11190 8620
rect 11210 8600 11220 8620
rect 12580 8620 12620 8630
rect 12580 8600 12590 8620
rect 12610 8600 12620 8620
rect 18680 8620 18720 8630
rect 10905 8575 10945 8585
rect 10980 8580 11000 8595
rect 11040 8580 11060 8595
rect 11180 8585 11280 8600
rect 10860 8550 10880 8565
rect 10920 8550 10940 8575
rect 10450 8340 10490 8350
rect 10450 8320 10460 8340
rect 10480 8320 10490 8340
rect 10710 8340 10750 8350
rect 10710 8320 10720 8340
rect 10740 8320 10750 8340
rect 10450 8305 10550 8320
rect 10530 8293 10550 8305
rect 10590 8293 10610 8308
rect 10650 8305 10750 8320
rect 10650 8293 10670 8305
rect 11260 8575 11280 8585
rect 11320 8575 11340 8590
rect 11380 8575 11400 8590
rect 11440 8575 11460 8590
rect 11500 8575 11520 8590
rect 11560 8575 11580 8590
rect 11620 8575 11640 8590
rect 11680 8575 11700 8590
rect 11740 8575 11760 8590
rect 11800 8575 11820 8590
rect 11860 8575 11880 8590
rect 11920 8575 11940 8590
rect 11980 8575 12000 8590
rect 12040 8575 12060 8590
rect 12100 8575 12120 8590
rect 12160 8575 12180 8590
rect 12220 8575 12240 8590
rect 12280 8575 12300 8590
rect 12340 8575 12360 8590
rect 12400 8575 12420 8590
rect 12460 8575 12480 8590
rect 12520 8585 12620 8600
rect 18405 8605 18445 8615
rect 18405 8585 18415 8605
rect 18435 8585 18445 8605
rect 18680 8600 18690 8620
rect 18710 8600 18720 8620
rect 20080 8620 20120 8630
rect 20080 8600 20090 8620
rect 20110 8600 20120 8620
rect 12520 8575 12540 8585
rect 18405 8575 18445 8585
rect 18480 8580 18500 8595
rect 18540 8580 18560 8595
rect 18680 8585 18780 8600
rect 10530 8215 10550 8230
rect 10590 8215 10610 8230
rect 10650 8215 10670 8230
rect 10860 8220 10880 8230
rect 10580 8205 10620 8215
rect 10580 8185 10590 8205
rect 10610 8185 10620 8205
rect 10580 8175 10620 8185
rect 10780 8205 10880 8220
rect 10920 8215 10940 8230
rect 10905 8205 10940 8215
rect 10780 8185 10790 8205
rect 10810 8185 10820 8205
rect 10780 8175 10820 8185
rect 10905 8185 10910 8205
rect 10930 8185 10940 8205
rect 10905 8175 10940 8185
rect 10980 8215 11000 8230
rect 11040 8220 11060 8230
rect 10980 8205 11015 8215
rect 11040 8205 11140 8220
rect 10980 8185 10990 8205
rect 11010 8185 11015 8205
rect 10980 8175 11015 8185
rect 11100 8185 11110 8205
rect 11130 8185 11140 8205
rect 11100 8175 11140 8185
rect 18360 8550 18380 8565
rect 18420 8550 18440 8575
rect 17950 8340 17990 8350
rect 17950 8320 17960 8340
rect 17980 8320 17990 8340
rect 18210 8340 18250 8350
rect 18210 8320 18220 8340
rect 18240 8320 18250 8340
rect 17950 8305 18050 8320
rect 18030 8293 18050 8305
rect 18090 8293 18110 8308
rect 18150 8305 18250 8320
rect 18150 8293 18170 8305
rect 12935 8240 12950 8255
rect 12990 8240 13005 8255
rect 13045 8240 13060 8255
rect 13100 8240 13115 8255
rect 13155 8240 13170 8255
rect 13210 8240 13225 8255
rect 13265 8240 13280 8255
rect 13320 8240 13335 8255
rect 13375 8240 13390 8255
rect 13430 8240 13445 8255
rect 13485 8240 13500 8255
rect 13540 8240 13555 8255
rect 13595 8240 13610 8255
rect 13650 8240 13665 8255
rect 13705 8240 13720 8255
rect 13760 8240 13775 8255
rect 13815 8240 13830 8255
rect 13870 8240 13885 8255
rect 13925 8240 13940 8255
rect 13980 8240 13995 8255
rect 14035 8240 14050 8255
rect 14090 8240 14105 8255
rect 11260 8160 11280 8175
rect 11320 8165 11340 8175
rect 11380 8165 11400 8175
rect 11440 8165 11460 8175
rect 11500 8165 11520 8175
rect 11560 8165 11580 8175
rect 11620 8165 11640 8175
rect 11680 8165 11700 8175
rect 11740 8165 11760 8175
rect 11800 8165 11820 8175
rect 11860 8165 11880 8175
rect 11920 8165 11940 8175
rect 11980 8165 12000 8175
rect 12040 8165 12060 8175
rect 12100 8165 12120 8175
rect 12160 8165 12180 8175
rect 12220 8165 12240 8175
rect 12280 8165 12300 8175
rect 12340 8165 12360 8175
rect 12400 8165 12420 8175
rect 12460 8165 12480 8175
rect 11320 8150 12480 8165
rect 12520 8160 12540 8175
rect 11823 8130 11831 8150
rect 11849 8130 11857 8150
rect 11823 8120 11857 8130
rect 11180 7940 11220 7950
rect 11180 7920 11190 7940
rect 11210 7920 11220 7940
rect 12580 7940 12620 7950
rect 18760 8575 18780 8585
rect 18820 8575 18840 8590
rect 18880 8575 18900 8590
rect 18940 8575 18960 8590
rect 19000 8575 19020 8590
rect 19060 8575 19080 8590
rect 19120 8575 19140 8590
rect 19180 8575 19200 8590
rect 19240 8575 19260 8590
rect 19300 8575 19320 8590
rect 19360 8575 19380 8590
rect 19420 8575 19440 8590
rect 19480 8575 19500 8590
rect 19540 8575 19560 8590
rect 19600 8575 19620 8590
rect 19660 8575 19680 8590
rect 19720 8575 19740 8590
rect 19780 8575 19800 8590
rect 19840 8575 19860 8590
rect 19900 8575 19920 8590
rect 19960 8575 19980 8590
rect 20020 8585 20120 8600
rect 20020 8575 20040 8585
rect 18030 8215 18050 8230
rect 18090 8215 18110 8230
rect 18150 8215 18170 8230
rect 18360 8220 18380 8230
rect 18080 8205 18120 8215
rect 18080 8185 18090 8205
rect 18110 8185 18120 8205
rect 18080 8175 18120 8185
rect 18280 8205 18380 8220
rect 18420 8215 18440 8230
rect 18405 8205 18440 8215
rect 18280 8185 18290 8205
rect 18310 8185 18320 8205
rect 18280 8175 18320 8185
rect 18405 8185 18410 8205
rect 18430 8185 18440 8205
rect 18405 8175 18440 8185
rect 18480 8215 18500 8230
rect 18540 8220 18560 8230
rect 18480 8205 18515 8215
rect 18540 8205 18640 8220
rect 18480 8185 18490 8205
rect 18510 8185 18515 8205
rect 18480 8175 18515 8185
rect 18600 8185 18610 8205
rect 18630 8185 18640 8205
rect 18600 8175 18640 8185
rect 20430 8240 20445 8255
rect 20485 8240 20500 8255
rect 20540 8240 20555 8255
rect 20595 8240 20610 8255
rect 20650 8240 20665 8255
rect 20705 8240 20720 8255
rect 20760 8240 20775 8255
rect 20815 8240 20830 8255
rect 20870 8240 20885 8255
rect 20925 8240 20940 8255
rect 20980 8240 20995 8255
rect 21035 8240 21050 8255
rect 21090 8240 21105 8255
rect 21145 8240 21160 8255
rect 21200 8240 21215 8255
rect 21255 8240 21270 8255
rect 21310 8240 21325 8255
rect 21365 8240 21380 8255
rect 21420 8240 21435 8255
rect 21475 8240 21490 8255
rect 21530 8240 21545 8255
rect 21585 8240 21600 8255
rect 18760 8160 18780 8175
rect 18820 8165 18840 8175
rect 18880 8165 18900 8175
rect 18940 8165 18960 8175
rect 19000 8165 19020 8175
rect 19060 8165 19080 8175
rect 19120 8165 19140 8175
rect 19180 8165 19200 8175
rect 19240 8165 19260 8175
rect 19300 8165 19320 8175
rect 19360 8165 19380 8175
rect 19420 8165 19440 8175
rect 19480 8165 19500 8175
rect 19540 8165 19560 8175
rect 19600 8165 19620 8175
rect 19660 8165 19680 8175
rect 19720 8165 19740 8175
rect 19780 8165 19800 8175
rect 19840 8165 19860 8175
rect 19900 8165 19920 8175
rect 19960 8165 19980 8175
rect 18820 8150 19980 8165
rect 20020 8160 20040 8175
rect 19323 8130 19331 8150
rect 19349 8130 19357 8150
rect 19323 8120 19357 8130
rect 18680 7940 18720 7950
rect 12580 7920 12590 7940
rect 12610 7920 12620 7940
rect 12935 7930 12950 7940
rect 11180 7905 11280 7920
rect 11260 7895 11280 7905
rect 11320 7895 11340 7910
rect 11380 7895 11400 7910
rect 11440 7895 11460 7910
rect 11500 7895 11520 7910
rect 11560 7895 11580 7910
rect 11620 7895 11640 7910
rect 11680 7895 11700 7910
rect 11740 7895 11760 7910
rect 11800 7895 11820 7910
rect 11860 7895 11880 7910
rect 11920 7895 11940 7910
rect 11980 7895 12000 7910
rect 12040 7895 12060 7910
rect 12100 7895 12120 7910
rect 12160 7895 12180 7910
rect 12220 7895 12240 7910
rect 12280 7895 12300 7910
rect 12340 7895 12360 7910
rect 12400 7895 12420 7910
rect 12460 7895 12480 7910
rect 12520 7905 12620 7920
rect 12855 7915 12950 7930
rect 12990 7930 13005 7940
rect 13045 7930 13060 7940
rect 13100 7930 13115 7940
rect 13155 7930 13170 7940
rect 13210 7930 13225 7940
rect 13265 7930 13280 7940
rect 13320 7930 13335 7940
rect 13375 7930 13390 7940
rect 13430 7930 13445 7940
rect 13485 7930 13500 7940
rect 13540 7930 13555 7940
rect 13595 7930 13610 7940
rect 13650 7930 13665 7940
rect 13705 7930 13720 7940
rect 13760 7930 13775 7940
rect 13815 7930 13830 7940
rect 13870 7930 13885 7940
rect 13925 7930 13940 7940
rect 13980 7930 13995 7940
rect 14035 7930 14050 7940
rect 12990 7915 14050 7930
rect 14090 7930 14105 7940
rect 14090 7915 14185 7930
rect 12520 7895 12540 7905
rect 12855 7895 12865 7915
rect 12885 7895 12895 7915
rect 9720 7620 9735 7635
rect 9775 7620 9790 7635
rect 9830 7620 9845 7635
rect 9885 7620 9900 7635
rect 9940 7620 9955 7635
rect 9995 7620 10010 7635
rect 10050 7620 10065 7635
rect 10105 7620 10120 7635
rect 10160 7620 10175 7635
rect 10215 7620 10230 7635
rect 10270 7620 10285 7635
rect 10325 7620 10340 7635
rect 10380 7620 10395 7635
rect 10435 7620 10450 7635
rect 10490 7620 10505 7635
rect 10545 7620 10560 7635
rect 10600 7620 10615 7635
rect 10655 7620 10670 7635
rect 10710 7620 10725 7635
rect 10765 7620 10780 7635
rect 10820 7620 10835 7635
rect 10875 7620 10890 7635
rect 9720 7510 9735 7520
rect 9640 7495 9735 7510
rect 9775 7510 9790 7520
rect 9830 7510 9845 7520
rect 9885 7510 9900 7520
rect 9940 7510 9955 7520
rect 9995 7510 10010 7520
rect 10050 7510 10065 7520
rect 10105 7510 10120 7520
rect 10160 7510 10175 7520
rect 10215 7510 10230 7520
rect 10270 7510 10285 7520
rect 10325 7510 10340 7520
rect 10380 7510 10395 7520
rect 10435 7510 10450 7520
rect 10490 7510 10505 7520
rect 10545 7510 10560 7520
rect 10600 7510 10615 7520
rect 10655 7510 10670 7520
rect 10710 7510 10725 7520
rect 10765 7510 10780 7520
rect 10820 7510 10835 7520
rect 9775 7495 10835 7510
rect 10875 7510 10890 7520
rect 10875 7495 10970 7510
rect 12855 7885 12895 7895
rect 13063 7895 13071 7915
rect 13089 7895 13097 7915
rect 13063 7885 13097 7895
rect 14145 7895 14155 7915
rect 14175 7895 14185 7915
rect 18680 7920 18690 7940
rect 18710 7920 18720 7940
rect 20080 7940 20120 7950
rect 20080 7920 20090 7940
rect 20110 7920 20120 7940
rect 20430 7930 20445 7940
rect 18680 7905 18780 7920
rect 18760 7895 18780 7905
rect 18820 7895 18840 7910
rect 18880 7895 18900 7910
rect 18940 7895 18960 7910
rect 19000 7895 19020 7910
rect 19060 7895 19080 7910
rect 19120 7895 19140 7910
rect 19180 7895 19200 7910
rect 19240 7895 19260 7910
rect 19300 7895 19320 7910
rect 19360 7895 19380 7910
rect 19420 7895 19440 7910
rect 19480 7895 19500 7910
rect 19540 7895 19560 7910
rect 19600 7895 19620 7910
rect 19660 7895 19680 7910
rect 19720 7895 19740 7910
rect 19780 7895 19800 7910
rect 19840 7895 19860 7910
rect 19900 7895 19920 7910
rect 19960 7895 19980 7910
rect 20020 7905 20120 7920
rect 20350 7915 20445 7930
rect 20485 7930 20500 7940
rect 20540 7930 20555 7940
rect 20595 7930 20610 7940
rect 20650 7930 20665 7940
rect 20705 7930 20720 7940
rect 20760 7930 20775 7940
rect 20815 7930 20830 7940
rect 20870 7930 20885 7940
rect 20925 7930 20940 7940
rect 20980 7930 20995 7940
rect 21035 7930 21050 7940
rect 21090 7930 21105 7940
rect 21145 7930 21160 7940
rect 21200 7930 21215 7940
rect 21255 7930 21270 7940
rect 21310 7930 21325 7940
rect 21365 7930 21380 7940
rect 21420 7930 21435 7940
rect 21475 7930 21490 7940
rect 21530 7930 21545 7940
rect 20485 7915 21545 7930
rect 21585 7930 21600 7940
rect 21585 7915 21680 7930
rect 20020 7895 20040 7905
rect 20350 7895 20360 7915
rect 20380 7895 20390 7915
rect 14145 7885 14185 7895
rect 12935 7620 12950 7635
rect 12990 7620 13005 7635
rect 13045 7620 13060 7635
rect 13100 7620 13115 7635
rect 13155 7620 13170 7635
rect 13210 7620 13225 7635
rect 13265 7620 13280 7635
rect 13320 7620 13335 7635
rect 13375 7620 13390 7635
rect 13430 7620 13445 7635
rect 13485 7620 13500 7635
rect 13540 7620 13555 7635
rect 13595 7620 13610 7635
rect 13650 7620 13665 7635
rect 13705 7620 13720 7635
rect 13760 7620 13775 7635
rect 13815 7620 13830 7635
rect 13870 7620 13885 7635
rect 13925 7620 13940 7635
rect 13980 7620 13995 7635
rect 14035 7620 14050 7635
rect 14090 7620 14105 7635
rect 17220 7620 17235 7635
rect 17275 7620 17290 7635
rect 17330 7620 17345 7635
rect 17385 7620 17400 7635
rect 17440 7620 17455 7635
rect 17495 7620 17510 7635
rect 17550 7620 17565 7635
rect 17605 7620 17620 7635
rect 17660 7620 17675 7635
rect 17715 7620 17730 7635
rect 17770 7620 17785 7635
rect 17825 7620 17840 7635
rect 17880 7620 17895 7635
rect 17935 7620 17950 7635
rect 17990 7620 18005 7635
rect 18045 7620 18060 7635
rect 18100 7620 18115 7635
rect 18155 7620 18170 7635
rect 18210 7620 18225 7635
rect 18265 7620 18280 7635
rect 18320 7620 18335 7635
rect 18375 7620 18390 7635
rect 12935 7510 12950 7520
rect 12855 7495 12950 7510
rect 12990 7510 13005 7520
rect 13045 7510 13060 7520
rect 13100 7510 13115 7520
rect 13155 7510 13170 7520
rect 13210 7510 13225 7520
rect 13265 7510 13280 7520
rect 13320 7510 13335 7520
rect 13375 7510 13390 7520
rect 13430 7510 13445 7520
rect 13485 7510 13500 7520
rect 13540 7510 13555 7520
rect 13595 7510 13610 7520
rect 13650 7510 13665 7520
rect 13705 7510 13720 7520
rect 13760 7510 13775 7520
rect 13815 7510 13830 7520
rect 13870 7510 13885 7520
rect 13925 7510 13940 7520
rect 13980 7510 13995 7520
rect 14035 7510 14050 7520
rect 12990 7495 14050 7510
rect 14090 7510 14105 7520
rect 17220 7510 17235 7520
rect 14090 7495 14185 7510
rect 9640 7475 9650 7495
rect 9670 7475 9680 7495
rect 9640 7465 9680 7475
rect 10820 7445 10835 7495
rect 10930 7475 10940 7495
rect 10960 7475 10970 7495
rect 11260 7480 11280 7495
rect 11320 7485 11340 7495
rect 11380 7485 11400 7495
rect 11440 7485 11460 7495
rect 11500 7485 11520 7495
rect 11560 7485 11580 7495
rect 11620 7485 11640 7495
rect 11680 7485 11700 7495
rect 11740 7485 11760 7495
rect 11800 7485 11820 7495
rect 11860 7485 11880 7495
rect 11920 7485 11940 7495
rect 11980 7485 12000 7495
rect 12040 7485 12060 7495
rect 12100 7485 12120 7495
rect 12160 7485 12180 7495
rect 12220 7485 12240 7495
rect 12280 7485 12300 7495
rect 12340 7485 12360 7495
rect 12400 7485 12420 7495
rect 12460 7485 12480 7495
rect 10930 7465 10970 7475
rect 11320 7470 12480 7485
rect 12520 7480 12540 7495
rect 12855 7475 12865 7495
rect 12885 7475 12895 7495
rect 11823 7450 11831 7470
rect 11849 7450 11857 7470
rect 12855 7465 12895 7475
rect 10813 7435 10847 7445
rect 11823 7440 11857 7450
rect 12990 7445 13005 7495
rect 14145 7475 14155 7495
rect 14175 7475 14185 7495
rect 14145 7465 14185 7475
rect 17140 7495 17235 7510
rect 17275 7510 17290 7520
rect 17330 7510 17345 7520
rect 17385 7510 17400 7520
rect 17440 7510 17455 7520
rect 17495 7510 17510 7520
rect 17550 7510 17565 7520
rect 17605 7510 17620 7520
rect 17660 7510 17675 7520
rect 17715 7510 17730 7520
rect 17770 7510 17785 7520
rect 17825 7510 17840 7520
rect 17880 7510 17895 7520
rect 17935 7510 17950 7520
rect 17990 7510 18005 7520
rect 18045 7510 18060 7520
rect 18100 7510 18115 7520
rect 18155 7510 18170 7520
rect 18210 7510 18225 7520
rect 18265 7510 18280 7520
rect 18320 7510 18335 7520
rect 17275 7495 18335 7510
rect 18375 7510 18390 7520
rect 18375 7495 18470 7510
rect 20350 7885 20390 7895
rect 20558 7895 20566 7915
rect 20584 7895 20592 7915
rect 20558 7885 20592 7895
rect 21640 7895 21650 7915
rect 21670 7895 21680 7915
rect 21640 7885 21680 7895
rect 20430 7620 20445 7635
rect 20485 7620 20500 7635
rect 20540 7620 20555 7635
rect 20595 7620 20610 7635
rect 20650 7620 20665 7635
rect 20705 7620 20720 7635
rect 20760 7620 20775 7635
rect 20815 7620 20830 7635
rect 20870 7620 20885 7635
rect 20925 7620 20940 7635
rect 20980 7620 20995 7635
rect 21035 7620 21050 7635
rect 21090 7620 21105 7635
rect 21145 7620 21160 7635
rect 21200 7620 21215 7635
rect 21255 7620 21270 7635
rect 21310 7620 21325 7635
rect 21365 7620 21380 7635
rect 21420 7620 21435 7635
rect 21475 7620 21490 7635
rect 21530 7620 21545 7635
rect 21585 7620 21600 7635
rect 20430 7510 20445 7520
rect 20350 7495 20445 7510
rect 20485 7510 20500 7520
rect 20540 7510 20555 7520
rect 20595 7510 20610 7520
rect 20650 7510 20665 7520
rect 20705 7510 20720 7520
rect 20760 7510 20775 7520
rect 20815 7510 20830 7520
rect 20870 7510 20885 7520
rect 20925 7510 20940 7520
rect 20980 7510 20995 7520
rect 21035 7510 21050 7520
rect 21090 7510 21105 7520
rect 21145 7510 21160 7520
rect 21200 7510 21215 7520
rect 21255 7510 21270 7520
rect 21310 7510 21325 7520
rect 21365 7510 21380 7520
rect 21420 7510 21435 7520
rect 21475 7510 21490 7520
rect 21530 7510 21545 7520
rect 20485 7495 21545 7510
rect 21585 7510 21600 7520
rect 21585 7495 21680 7510
rect 17140 7475 17150 7495
rect 17170 7475 17180 7495
rect 17140 7465 17180 7475
rect 18320 7445 18335 7495
rect 18430 7475 18440 7495
rect 18460 7475 18470 7495
rect 18760 7480 18780 7495
rect 18820 7485 18840 7495
rect 18880 7485 18900 7495
rect 18940 7485 18960 7495
rect 19000 7485 19020 7495
rect 19060 7485 19080 7495
rect 19120 7485 19140 7495
rect 19180 7485 19200 7495
rect 19240 7485 19260 7495
rect 19300 7485 19320 7495
rect 19360 7485 19380 7495
rect 19420 7485 19440 7495
rect 19480 7485 19500 7495
rect 19540 7485 19560 7495
rect 19600 7485 19620 7495
rect 19660 7485 19680 7495
rect 19720 7485 19740 7495
rect 19780 7485 19800 7495
rect 19840 7485 19860 7495
rect 19900 7485 19920 7495
rect 19960 7485 19980 7495
rect 18430 7465 18470 7475
rect 18820 7470 19980 7485
rect 20020 7480 20040 7495
rect 20350 7475 20360 7495
rect 20380 7475 20390 7495
rect 19323 7450 19331 7470
rect 19349 7450 19357 7470
rect 20350 7465 20390 7475
rect 10813 7415 10821 7435
rect 10839 7415 10847 7435
rect 10813 7405 10847 7415
rect 12978 7435 13012 7445
rect 12978 7415 12986 7435
rect 13004 7415 13012 7435
rect 12978 7405 13012 7415
rect 18313 7435 18347 7445
rect 19323 7440 19357 7450
rect 20485 7445 20500 7495
rect 21640 7475 21650 7495
rect 21670 7475 21680 7495
rect 21640 7465 21680 7475
rect 18313 7415 18321 7435
rect 18339 7415 18347 7435
rect 18313 7405 18347 7415
rect 20473 7435 20507 7445
rect 20473 7415 20481 7435
rect 20499 7415 20507 7435
rect 20473 7405 20507 7415
rect 10813 7275 10847 7285
rect 10813 7255 10821 7275
rect 10839 7255 10847 7275
rect 10813 7245 10847 7255
rect 12978 7275 13012 7285
rect 12978 7255 12986 7275
rect 13004 7255 13012 7275
rect 12978 7245 13012 7255
rect 18313 7275 18347 7285
rect 18313 7255 18321 7275
rect 18339 7255 18347 7275
rect 18313 7245 18347 7255
rect 20473 7275 20507 7285
rect 20473 7255 20481 7275
rect 20499 7255 20507 7275
rect 20473 7245 20507 7255
rect 9640 7215 9680 7225
rect 9640 7195 9650 7215
rect 9670 7195 9680 7215
rect 10820 7195 10835 7245
rect 10930 7215 10970 7225
rect 10930 7195 10940 7215
rect 10960 7195 10970 7215
rect 9640 7180 9735 7195
rect 9720 7170 9735 7180
rect 9775 7180 10835 7195
rect 9775 7170 9790 7180
rect 9830 7170 9845 7180
rect 9885 7170 9900 7180
rect 9940 7170 9955 7180
rect 9995 7170 10010 7180
rect 10050 7170 10065 7180
rect 10105 7170 10120 7180
rect 10160 7170 10175 7180
rect 10215 7170 10230 7180
rect 10270 7170 10285 7180
rect 10325 7170 10340 7180
rect 10380 7170 10395 7180
rect 10435 7170 10450 7180
rect 10490 7170 10505 7180
rect 10545 7170 10560 7180
rect 10600 7170 10615 7180
rect 10655 7170 10670 7180
rect 10710 7170 10725 7180
rect 10765 7170 10780 7180
rect 10820 7170 10835 7180
rect 10875 7180 10970 7195
rect 12855 7215 12895 7225
rect 12855 7195 12865 7215
rect 12885 7195 12895 7215
rect 12990 7195 13005 7245
rect 14145 7215 14185 7225
rect 14145 7195 14155 7215
rect 14175 7195 14185 7215
rect 12855 7180 12950 7195
rect 10875 7170 10890 7180
rect 12935 7170 12950 7180
rect 12990 7180 14050 7195
rect 12990 7170 13005 7180
rect 13045 7170 13060 7180
rect 13100 7170 13115 7180
rect 13155 7170 13170 7180
rect 13210 7170 13225 7180
rect 13265 7170 13280 7180
rect 13320 7170 13335 7180
rect 13375 7170 13390 7180
rect 13430 7170 13445 7180
rect 13485 7170 13500 7180
rect 13540 7170 13555 7180
rect 13595 7170 13610 7180
rect 13650 7170 13665 7180
rect 13705 7170 13720 7180
rect 13760 7170 13775 7180
rect 13815 7170 13830 7180
rect 13870 7170 13885 7180
rect 13925 7170 13940 7180
rect 13980 7170 13995 7180
rect 14035 7170 14050 7180
rect 14090 7180 14185 7195
rect 17140 7215 17180 7225
rect 17140 7195 17150 7215
rect 17170 7195 17180 7215
rect 18320 7195 18335 7245
rect 18430 7215 18470 7225
rect 18430 7195 18440 7215
rect 18460 7195 18470 7215
rect 17140 7180 17235 7195
rect 14090 7170 14105 7180
rect 17220 7170 17235 7180
rect 17275 7180 18335 7195
rect 17275 7170 17290 7180
rect 17330 7170 17345 7180
rect 17385 7170 17400 7180
rect 17440 7170 17455 7180
rect 17495 7170 17510 7180
rect 17550 7170 17565 7180
rect 17605 7170 17620 7180
rect 17660 7170 17675 7180
rect 17715 7170 17730 7180
rect 17770 7170 17785 7180
rect 17825 7170 17840 7180
rect 17880 7170 17895 7180
rect 17935 7170 17950 7180
rect 17990 7170 18005 7180
rect 18045 7170 18060 7180
rect 18100 7170 18115 7180
rect 18155 7170 18170 7180
rect 18210 7170 18225 7180
rect 18265 7170 18280 7180
rect 18320 7170 18335 7180
rect 18375 7180 18470 7195
rect 20350 7215 20390 7225
rect 20350 7195 20360 7215
rect 20380 7195 20390 7215
rect 20485 7195 20500 7245
rect 21640 7215 21680 7225
rect 21640 7195 21650 7215
rect 21670 7195 21680 7215
rect 20350 7180 20445 7195
rect 18375 7170 18390 7180
rect 20430 7170 20445 7180
rect 20485 7180 21545 7195
rect 20485 7170 20500 7180
rect 20540 7170 20555 7180
rect 20595 7170 20610 7180
rect 20650 7170 20665 7180
rect 20705 7170 20720 7180
rect 20760 7170 20775 7180
rect 20815 7170 20830 7180
rect 20870 7170 20885 7180
rect 20925 7170 20940 7180
rect 20980 7170 20995 7180
rect 21035 7170 21050 7180
rect 21090 7170 21105 7180
rect 21145 7170 21160 7180
rect 21200 7170 21215 7180
rect 21255 7170 21270 7180
rect 21310 7170 21325 7180
rect 21365 7170 21380 7180
rect 21420 7170 21435 7180
rect 21475 7170 21490 7180
rect 21530 7170 21545 7180
rect 21585 7180 21680 7195
rect 21585 7170 21600 7180
rect 11315 7130 11330 7145
rect 11370 7140 12430 7155
rect 11370 7130 11385 7140
rect 11425 7130 11440 7140
rect 11480 7130 11495 7140
rect 11535 7130 11550 7140
rect 11590 7130 11605 7140
rect 11645 7130 11660 7140
rect 11700 7130 11715 7140
rect 11755 7130 11770 7140
rect 11810 7130 11825 7140
rect 11865 7130 11880 7140
rect 11920 7130 11935 7140
rect 11975 7130 11990 7140
rect 12030 7130 12045 7140
rect 12085 7130 12100 7140
rect 12140 7130 12155 7140
rect 12195 7130 12210 7140
rect 12250 7130 12265 7140
rect 12305 7130 12320 7140
rect 12360 7130 12375 7140
rect 12415 7130 12430 7140
rect 12470 7130 12485 7145
rect 9720 7005 9735 7020
rect 9775 7005 9790 7020
rect 9830 7005 9845 7020
rect 9885 7005 9900 7020
rect 9940 7005 9955 7020
rect 9995 7005 10010 7020
rect 10050 7005 10065 7020
rect 10105 7005 10120 7020
rect 10160 7005 10175 7020
rect 10215 7005 10230 7020
rect 10270 7005 10285 7020
rect 10325 7005 10340 7020
rect 10380 7005 10395 7020
rect 10435 7005 10450 7020
rect 10490 7005 10505 7020
rect 10545 7005 10560 7020
rect 10600 7005 10615 7020
rect 10655 7005 10670 7020
rect 10710 7005 10725 7020
rect 10765 7005 10780 7020
rect 10820 7005 10835 7020
rect 10875 7005 10890 7020
rect 18815 7130 18830 7145
rect 18870 7140 19930 7155
rect 18870 7130 18885 7140
rect 18925 7130 18940 7140
rect 18980 7130 18995 7140
rect 19035 7130 19050 7140
rect 19090 7130 19105 7140
rect 19145 7130 19160 7140
rect 19200 7130 19215 7140
rect 19255 7130 19270 7140
rect 19310 7130 19325 7140
rect 19365 7130 19380 7140
rect 19420 7130 19435 7140
rect 19475 7130 19490 7140
rect 19530 7130 19545 7140
rect 19585 7130 19600 7140
rect 19640 7130 19655 7140
rect 19695 7130 19710 7140
rect 19750 7130 19765 7140
rect 19805 7130 19820 7140
rect 19860 7130 19875 7140
rect 19915 7130 19930 7140
rect 19970 7130 19985 7145
rect 12935 7005 12950 7020
rect 12990 7005 13005 7020
rect 13045 7005 13060 7020
rect 13100 7005 13115 7020
rect 13155 7005 13170 7020
rect 13210 7005 13225 7020
rect 13265 7005 13280 7020
rect 13320 7005 13335 7020
rect 13375 7005 13390 7020
rect 13430 7005 13445 7020
rect 13485 7005 13500 7020
rect 13540 7005 13555 7020
rect 13595 7005 13610 7020
rect 13650 7005 13665 7020
rect 13705 7005 13720 7020
rect 13760 7005 13775 7020
rect 13815 7005 13830 7020
rect 13870 7005 13885 7020
rect 13925 7005 13940 7020
rect 13980 7005 13995 7020
rect 14035 7005 14050 7020
rect 14090 7005 14105 7020
rect 17220 7005 17235 7020
rect 17275 7005 17290 7020
rect 17330 7005 17345 7020
rect 17385 7005 17400 7020
rect 17440 7005 17455 7020
rect 17495 7005 17510 7020
rect 17550 7005 17565 7020
rect 17605 7005 17620 7020
rect 17660 7005 17675 7020
rect 17715 7005 17730 7020
rect 17770 7005 17785 7020
rect 17825 7005 17840 7020
rect 17880 7005 17895 7020
rect 17935 7005 17950 7020
rect 17990 7005 18005 7020
rect 18045 7005 18060 7020
rect 18100 7005 18115 7020
rect 18155 7005 18170 7020
rect 18210 7005 18225 7020
rect 18265 7005 18280 7020
rect 18320 7005 18335 7020
rect 18375 7005 18390 7020
rect 20430 7005 20445 7020
rect 20485 7005 20500 7020
rect 20540 7005 20555 7020
rect 20595 7005 20610 7020
rect 20650 7005 20665 7020
rect 20705 7005 20720 7020
rect 20760 7005 20775 7020
rect 20815 7005 20830 7020
rect 20870 7005 20885 7020
rect 20925 7005 20940 7020
rect 20980 7005 20995 7020
rect 21035 7005 21050 7020
rect 21090 7005 21105 7020
rect 21145 7005 21160 7020
rect 21200 7005 21215 7020
rect 21255 7005 21270 7020
rect 21310 7005 21325 7020
rect 21365 7005 21380 7020
rect 21420 7005 21435 7020
rect 21475 7005 21490 7020
rect 21530 7005 21545 7020
rect 21585 7005 21600 7020
rect 11315 6970 11330 6980
rect 11235 6955 11330 6970
rect 11370 6965 11385 6980
rect 11425 6965 11440 6980
rect 11480 6965 11495 6980
rect 11535 6965 11550 6980
rect 11590 6965 11605 6980
rect 11645 6965 11660 6980
rect 11700 6965 11715 6980
rect 11755 6965 11770 6980
rect 11810 6965 11825 6980
rect 11865 6965 11880 6980
rect 11920 6965 11935 6980
rect 11975 6965 11990 6980
rect 12030 6965 12045 6980
rect 12085 6965 12100 6980
rect 12140 6965 12155 6980
rect 12195 6965 12210 6980
rect 12250 6965 12265 6980
rect 12305 6965 12320 6980
rect 12360 6965 12375 6980
rect 12415 6965 12430 6980
rect 12470 6970 12485 6980
rect 18815 6970 18830 6980
rect 12470 6955 12565 6970
rect 11235 6935 11245 6955
rect 11265 6935 11275 6955
rect 11235 6925 11275 6935
rect 12525 6935 12535 6955
rect 12555 6935 12565 6955
rect 12525 6925 12565 6935
rect 18735 6955 18830 6970
rect 18870 6965 18885 6980
rect 18925 6965 18940 6980
rect 18980 6965 18995 6980
rect 19035 6965 19050 6980
rect 19090 6965 19105 6980
rect 19145 6965 19160 6980
rect 19200 6965 19215 6980
rect 19255 6965 19270 6980
rect 19310 6965 19325 6980
rect 19365 6965 19380 6980
rect 19420 6965 19435 6980
rect 19475 6965 19490 6980
rect 19530 6965 19545 6980
rect 19585 6965 19600 6980
rect 19640 6965 19655 6980
rect 19695 6965 19710 6980
rect 19750 6965 19765 6980
rect 19805 6965 19820 6980
rect 19860 6965 19875 6980
rect 19915 6965 19930 6980
rect 19970 6970 19985 6980
rect 19970 6955 20065 6970
rect 18735 6935 18745 6955
rect 18765 6935 18775 6955
rect 18735 6925 18775 6935
rect 20025 6935 20035 6955
rect 20055 6935 20065 6955
rect 20025 6925 20065 6935
rect 20450 6900 20490 6910
rect 20450 6880 20460 6900
rect 20480 6880 20490 6900
rect 20860 6900 20900 6910
rect 20860 6880 20870 6900
rect 20890 6880 20900 6900
rect 20450 6865 20545 6880
rect 20530 6855 20545 6865
rect 20585 6855 20600 6870
rect 20640 6855 20655 6870
rect 20695 6855 20710 6870
rect 20750 6855 20765 6870
rect 20805 6865 20900 6880
rect 20805 6855 20820 6865
rect 11237 6710 11269 6720
rect 11237 6690 11243 6710
rect 11260 6690 11269 6710
rect 11457 6710 11489 6720
rect 11457 6690 11463 6710
rect 11480 6690 11489 6710
rect 11180 6680 11269 6690
rect 11400 6680 11489 6690
rect 11601 6710 11635 6720
rect 11601 6690 11610 6710
rect 11627 6690 11635 6710
rect 11867 6710 11899 6720
rect 11867 6695 11876 6710
rect 11601 6680 11635 6690
rect 11865 6690 11876 6695
rect 11893 6690 11899 6710
rect 12277 6710 12309 6720
rect 12277 6690 12283 6710
rect 12300 6690 12309 6710
rect 12497 6710 12529 6720
rect 12497 6690 12503 6710
rect 12520 6690 12529 6710
rect 11865 6680 11899 6690
rect 12220 6680 12309 6690
rect 12440 6680 12529 6690
rect 12641 6710 12675 6720
rect 12641 6690 12650 6710
rect 12667 6690 12675 6710
rect 18737 6710 18769 6720
rect 18737 6690 18743 6710
rect 18760 6690 18769 6710
rect 18957 6710 18989 6720
rect 18957 6690 18963 6710
rect 18980 6690 18989 6710
rect 12641 6680 12675 6690
rect 18680 6680 18769 6690
rect 18900 6680 18989 6690
rect 19101 6710 19135 6720
rect 19101 6690 19110 6710
rect 19127 6690 19135 6710
rect 19367 6710 19399 6720
rect 19367 6695 19376 6710
rect 19101 6680 19135 6690
rect 19365 6690 19376 6695
rect 19393 6690 19399 6710
rect 19777 6710 19809 6720
rect 19777 6690 19783 6710
rect 19800 6690 19809 6710
rect 19997 6710 20029 6720
rect 19997 6690 20003 6710
rect 20020 6690 20029 6710
rect 19365 6680 19399 6690
rect 19720 6680 19809 6690
rect 19940 6680 20029 6690
rect 20141 6710 20175 6720
rect 20141 6690 20150 6710
rect 20167 6690 20175 6710
rect 20530 6690 20545 6705
rect 20585 6695 20600 6705
rect 20640 6695 20655 6705
rect 20695 6695 20710 6705
rect 20750 6695 20765 6705
rect 20141 6680 20175 6690
rect 20585 6685 20765 6695
rect 20805 6690 20820 6705
rect 20566 6680 20765 6685
rect 11070 6665 11085 6680
rect 11125 6665 11140 6680
rect 11180 6675 11250 6680
rect 11180 6665 11195 6675
rect 11235 6665 11250 6675
rect 11290 6665 11305 6680
rect 11345 6665 11360 6680
rect 11400 6675 11470 6680
rect 11400 6665 11415 6675
rect 11455 6665 11470 6675
rect 11510 6665 11525 6680
rect 11565 6665 11580 6680
rect 11620 6665 11635 6680
rect 11675 6665 11690 6680
rect 11810 6665 11825 6680
rect 11865 6665 11880 6680
rect 11920 6665 11935 6680
rect 11975 6665 11990 6680
rect 12110 6665 12125 6680
rect 12165 6665 12180 6680
rect 12220 6675 12290 6680
rect 12220 6665 12235 6675
rect 12275 6665 12290 6675
rect 12330 6665 12345 6680
rect 12385 6665 12400 6680
rect 12440 6675 12510 6680
rect 12440 6665 12455 6675
rect 12495 6665 12510 6675
rect 12550 6665 12565 6680
rect 12605 6665 12620 6680
rect 12660 6665 12675 6680
rect 12715 6665 12730 6680
rect 18570 6665 18585 6680
rect 18625 6665 18640 6680
rect 18680 6675 18750 6680
rect 18680 6665 18695 6675
rect 18735 6665 18750 6675
rect 18790 6665 18805 6680
rect 18845 6665 18860 6680
rect 18900 6675 18970 6680
rect 18900 6665 18915 6675
rect 18955 6665 18970 6675
rect 19010 6665 19025 6680
rect 19065 6665 19080 6680
rect 19120 6665 19135 6680
rect 19175 6665 19190 6680
rect 19310 6665 19325 6680
rect 19365 6665 19380 6680
rect 19420 6665 19435 6680
rect 19475 6665 19490 6680
rect 19610 6665 19625 6680
rect 19665 6665 19680 6680
rect 19720 6675 19790 6680
rect 19720 6665 19735 6675
rect 19775 6665 19790 6675
rect 19830 6665 19845 6680
rect 19885 6665 19900 6680
rect 19940 6675 20010 6680
rect 19940 6665 19955 6675
rect 19995 6665 20010 6675
rect 20050 6665 20065 6680
rect 20105 6665 20120 6680
rect 20160 6665 20175 6680
rect 20215 6665 20230 6680
rect 20566 6675 20600 6680
rect 20566 6655 20571 6675
rect 20591 6670 20600 6675
rect 20591 6655 20598 6670
rect 20566 6645 20598 6655
rect 20471 6565 20503 6575
rect 20471 6545 20476 6565
rect 20496 6550 20503 6565
rect 20847 6565 20879 6575
rect 20847 6550 20854 6565
rect 20496 6545 20505 6550
rect 20471 6535 20505 6545
rect 20845 6545 20854 6550
rect 20874 6545 20879 6565
rect 20845 6535 20879 6545
rect 20435 6520 20450 6535
rect 20490 6520 20505 6535
rect 20545 6520 20560 6535
rect 20600 6520 20615 6535
rect 20735 6520 20750 6535
rect 20790 6520 20805 6535
rect 20845 6520 20860 6535
rect 20900 6520 20915 6535
rect 11070 6505 11085 6515
rect 10990 6490 11085 6505
rect 11125 6500 11140 6515
rect 11180 6500 11195 6515
rect 11235 6500 11250 6515
rect 11290 6505 11305 6515
rect 11345 6505 11360 6515
rect 11106 6490 11140 6500
rect 11290 6490 11360 6505
rect 11400 6500 11415 6515
rect 11455 6500 11470 6515
rect 11510 6505 11525 6515
rect 11565 6505 11580 6515
rect 11510 6490 11580 6505
rect 11620 6500 11635 6515
rect 11675 6505 11690 6515
rect 11810 6505 11825 6515
rect 11675 6490 11825 6505
rect 11865 6500 11880 6515
rect 11920 6500 11935 6515
rect 11975 6505 11990 6515
rect 12110 6505 12125 6515
rect 11920 6490 11954 6500
rect 11975 6490 12125 6505
rect 12165 6500 12180 6515
rect 12220 6500 12235 6515
rect 12275 6500 12290 6515
rect 12330 6505 12345 6515
rect 12385 6505 12400 6515
rect 12146 6490 12180 6500
rect 12330 6490 12400 6505
rect 12440 6500 12455 6515
rect 12495 6500 12510 6515
rect 12550 6505 12565 6515
rect 12605 6505 12620 6515
rect 12550 6490 12620 6505
rect 12660 6500 12675 6515
rect 12715 6505 12730 6515
rect 18570 6505 18585 6515
rect 12715 6490 12810 6505
rect 10990 6470 11000 6490
rect 11020 6470 11030 6490
rect 10990 6460 11030 6470
rect 11106 6470 11112 6490
rect 11129 6470 11138 6490
rect 11106 6460 11138 6470
rect 11305 6470 11315 6490
rect 11335 6470 11345 6490
rect 11305 6460 11345 6470
rect 11525 6470 11535 6490
rect 11555 6470 11565 6490
rect 11525 6460 11565 6470
rect 11730 6470 11740 6490
rect 11760 6470 11770 6490
rect 11730 6460 11770 6470
rect 11922 6470 11928 6490
rect 11945 6470 11954 6490
rect 11922 6460 11954 6470
rect 12030 6470 12040 6490
rect 12060 6470 12070 6490
rect 12030 6460 12070 6470
rect 12146 6470 12152 6490
rect 12169 6470 12178 6490
rect 12146 6460 12178 6470
rect 12345 6470 12355 6490
rect 12375 6470 12385 6490
rect 12345 6460 12385 6470
rect 12565 6470 12575 6490
rect 12595 6470 12605 6490
rect 12565 6460 12605 6470
rect 12770 6470 12780 6490
rect 12800 6470 12810 6490
rect 12770 6460 12810 6470
rect 18490 6490 18585 6505
rect 18625 6500 18640 6515
rect 18680 6500 18695 6515
rect 18735 6500 18750 6515
rect 18790 6505 18805 6515
rect 18845 6505 18860 6515
rect 18606 6490 18640 6500
rect 18790 6490 18860 6505
rect 18900 6500 18915 6515
rect 18955 6500 18970 6515
rect 19010 6505 19025 6515
rect 19065 6505 19080 6515
rect 19010 6490 19080 6505
rect 19120 6500 19135 6515
rect 19175 6505 19190 6515
rect 19310 6505 19325 6515
rect 19175 6490 19325 6505
rect 19365 6500 19380 6515
rect 19420 6500 19435 6515
rect 19475 6505 19490 6515
rect 19610 6505 19625 6515
rect 19420 6490 19454 6500
rect 19475 6490 19625 6505
rect 19665 6500 19680 6515
rect 19720 6500 19735 6515
rect 19775 6500 19790 6515
rect 19830 6505 19845 6515
rect 19885 6505 19900 6515
rect 19646 6490 19680 6500
rect 19830 6490 19900 6505
rect 19940 6500 19955 6515
rect 19995 6500 20010 6515
rect 20050 6505 20065 6515
rect 20105 6505 20120 6515
rect 20050 6490 20120 6505
rect 20160 6500 20175 6515
rect 20215 6505 20230 6515
rect 20215 6490 20310 6505
rect 18490 6470 18500 6490
rect 18520 6470 18530 6490
rect 18490 6460 18530 6470
rect 18606 6470 18612 6490
rect 18629 6470 18638 6490
rect 18606 6460 18638 6470
rect 18805 6470 18815 6490
rect 18835 6470 18845 6490
rect 18805 6460 18845 6470
rect 19025 6470 19035 6490
rect 19055 6470 19065 6490
rect 19025 6460 19065 6470
rect 19230 6470 19240 6490
rect 19260 6470 19270 6490
rect 19230 6460 19270 6470
rect 19422 6470 19428 6490
rect 19445 6470 19454 6490
rect 19422 6460 19454 6470
rect 19530 6470 19540 6490
rect 19560 6470 19570 6490
rect 19530 6460 19570 6470
rect 19646 6470 19652 6490
rect 19669 6470 19678 6490
rect 19646 6460 19678 6470
rect 19845 6470 19855 6490
rect 19875 6470 19885 6490
rect 19845 6460 19885 6470
rect 20065 6470 20075 6490
rect 20095 6470 20105 6490
rect 20065 6460 20105 6470
rect 20270 6470 20280 6490
rect 20300 6470 20310 6490
rect 20270 6460 20310 6470
rect 20435 6360 20450 6370
rect 20355 6345 20450 6360
rect 20490 6355 20505 6370
rect 20545 6355 20560 6370
rect 20526 6345 20560 6355
rect 20600 6360 20615 6370
rect 20735 6360 20750 6370
rect 20600 6345 20750 6360
rect 20790 6355 20805 6370
rect 20845 6355 20860 6370
rect 20900 6360 20915 6370
rect 20790 6345 20824 6355
rect 20900 6345 20995 6360
rect 10668 6330 10702 6340
rect 10668 6310 10676 6330
rect 10694 6310 10702 6330
rect 13098 6330 13132 6340
rect 13098 6310 13106 6330
rect 13124 6310 13132 6330
rect 20355 6325 20365 6345
rect 20385 6325 20395 6345
rect 20355 6315 20395 6325
rect 20526 6325 20533 6345
rect 20553 6340 20560 6345
rect 20553 6325 20558 6340
rect 20526 6315 20558 6325
rect 20655 6325 20665 6345
rect 20685 6325 20695 6345
rect 20790 6340 20797 6345
rect 20655 6315 20695 6325
rect 20792 6325 20797 6340
rect 20817 6325 20824 6345
rect 20792 6315 20824 6325
rect 20955 6325 20965 6345
rect 20985 6325 20995 6345
rect 20955 6315 20995 6325
rect 9705 6285 9765 6300
rect 9805 6295 10765 6310
rect 9805 6285 9865 6295
rect 9905 6285 9965 6295
rect 10005 6285 10065 6295
rect 10105 6285 10165 6295
rect 10205 6285 10265 6295
rect 10305 6285 10365 6295
rect 10405 6285 10465 6295
rect 10505 6285 10565 6295
rect 10605 6285 10665 6295
rect 10705 6285 10765 6295
rect 10805 6285 10865 6300
rect 12935 6285 12995 6300
rect 13035 6295 13995 6310
rect 13035 6285 13095 6295
rect 13135 6285 13195 6295
rect 13235 6285 13295 6295
rect 13335 6285 13395 6295
rect 13435 6285 13495 6295
rect 13535 6285 13595 6295
rect 13635 6285 13695 6295
rect 13735 6285 13795 6295
rect 13835 6285 13895 6295
rect 13935 6285 13995 6295
rect 14035 6285 14095 6300
rect 20095 6285 20135 6295
rect 12595 6245 12635 6255
rect 12595 6240 12605 6245
rect 11815 6230 11845 6240
rect 11815 6210 11820 6230
rect 11840 6210 11845 6230
rect 12510 6225 12605 6240
rect 12625 6225 12635 6245
rect 11245 6185 11260 6200
rect 11300 6195 12360 6210
rect 11300 6185 11315 6195
rect 11355 6185 11370 6195
rect 11410 6185 11425 6195
rect 11465 6185 11480 6195
rect 11520 6185 11535 6195
rect 11575 6185 11590 6195
rect 11630 6185 11645 6195
rect 11685 6185 11700 6195
rect 11740 6185 11755 6195
rect 11795 6185 11810 6195
rect 11850 6185 11865 6195
rect 11905 6185 11920 6195
rect 11960 6185 11975 6195
rect 12015 6185 12030 6195
rect 12070 6185 12085 6195
rect 12125 6185 12140 6195
rect 12180 6185 12195 6195
rect 12235 6185 12250 6195
rect 12290 6185 12305 6195
rect 12345 6185 12360 6195
rect 12400 6195 12470 6210
rect 12400 6185 12415 6195
rect 12455 6185 12470 6195
rect 12510 6185 12525 6225
rect 12595 6215 12635 6225
rect 12565 6185 12580 6200
rect 9705 5995 9765 6005
rect 9625 5980 9765 5995
rect 9805 5990 9865 6005
rect 9905 5990 9965 6005
rect 10005 5990 10065 6005
rect 10105 5990 10165 6005
rect 10205 5990 10265 6005
rect 10305 5990 10365 6005
rect 10405 5990 10465 6005
rect 10505 5990 10565 6005
rect 10605 5990 10665 6005
rect 10705 5990 10765 6005
rect 10805 5995 10865 6005
rect 10805 5980 10945 5995
rect 9625 5960 9635 5980
rect 9655 5960 9665 5980
rect 9625 5950 9665 5960
rect 10905 5960 10915 5980
rect 10935 5960 10945 5980
rect 10905 5950 10945 5960
rect 20095 6280 20105 6285
rect 19315 6270 19345 6280
rect 19315 6250 19320 6270
rect 19340 6250 19345 6270
rect 20010 6265 20105 6280
rect 20125 6265 20135 6285
rect 18745 6225 18760 6240
rect 18800 6235 19860 6250
rect 18800 6225 18815 6235
rect 18855 6225 18870 6235
rect 18910 6225 18925 6235
rect 18965 6225 18980 6235
rect 19020 6225 19035 6235
rect 19075 6225 19090 6235
rect 19130 6225 19145 6235
rect 19185 6225 19200 6235
rect 19240 6225 19255 6235
rect 19295 6225 19310 6235
rect 19350 6225 19365 6235
rect 19405 6225 19420 6235
rect 19460 6225 19475 6235
rect 19515 6225 19530 6235
rect 19570 6225 19585 6235
rect 19625 6225 19640 6235
rect 19680 6225 19695 6235
rect 19735 6225 19750 6235
rect 19790 6225 19805 6235
rect 19845 6225 19860 6235
rect 19900 6235 19970 6250
rect 19900 6225 19915 6235
rect 19955 6225 19970 6235
rect 20010 6225 20025 6265
rect 20095 6255 20135 6265
rect 20065 6225 20080 6240
rect 12935 5995 12995 6005
rect 12855 5980 12995 5995
rect 13035 5990 13095 6005
rect 13135 5990 13195 6005
rect 13235 5990 13295 6005
rect 13335 5990 13395 6005
rect 13435 5990 13495 6005
rect 13535 5990 13595 6005
rect 13635 5990 13695 6005
rect 13735 5990 13795 6005
rect 13835 5990 13895 6005
rect 13935 5990 13995 6005
rect 14035 5995 14095 6005
rect 14035 5980 14175 5995
rect 12855 5960 12865 5980
rect 12885 5960 12895 5980
rect 12855 5950 12895 5960
rect 14135 5960 14145 5980
rect 14165 5960 14175 5980
rect 20585 6180 20600 6195
rect 20640 6180 20655 6195
rect 20695 6180 20710 6195
rect 20750 6180 20765 6195
rect 20585 6020 20600 6030
rect 20505 6005 20600 6020
rect 20640 6020 20655 6030
rect 20695 6020 20710 6030
rect 20640 6015 20710 6020
rect 20750 6020 20765 6030
rect 20640 6005 20725 6015
rect 20750 6005 20845 6020
rect 20505 5985 20515 6005
rect 20535 5985 20545 6005
rect 20505 5975 20545 5985
rect 20685 5985 20695 6005
rect 20715 5985 20725 6005
rect 20685 5975 20725 5985
rect 20805 5985 20815 6005
rect 20835 5985 20845 6005
rect 20805 5975 20845 5985
rect 18745 5960 18760 5975
rect 18800 5960 18815 5975
rect 18855 5960 18870 5975
rect 18910 5960 18925 5975
rect 18965 5960 18980 5975
rect 19020 5960 19035 5975
rect 19075 5960 19090 5975
rect 19130 5960 19145 5975
rect 19185 5960 19200 5975
rect 19240 5960 19255 5975
rect 19295 5960 19310 5975
rect 19350 5960 19365 5975
rect 19405 5960 19420 5975
rect 19460 5960 19475 5975
rect 19515 5960 19530 5975
rect 19570 5960 19585 5975
rect 19625 5960 19640 5975
rect 19680 5960 19695 5975
rect 19735 5960 19750 5975
rect 19790 5960 19805 5975
rect 19845 5960 19860 5975
rect 19900 5960 19915 5975
rect 19955 5960 19970 5975
rect 20010 5960 20025 5975
rect 20065 5960 20080 5975
rect 14135 5950 14175 5960
rect 18665 5950 18760 5960
rect 11245 5920 11260 5935
rect 11300 5920 11315 5935
rect 11355 5920 11370 5935
rect 11410 5920 11425 5935
rect 11465 5920 11480 5935
rect 11520 5920 11535 5935
rect 11575 5920 11590 5935
rect 11630 5920 11645 5935
rect 11685 5920 11700 5935
rect 11740 5920 11755 5935
rect 11795 5920 11810 5935
rect 11850 5920 11865 5935
rect 11905 5920 11920 5935
rect 11960 5920 11975 5935
rect 12015 5920 12030 5935
rect 12070 5920 12085 5935
rect 12125 5920 12140 5935
rect 12180 5920 12195 5935
rect 12235 5920 12250 5935
rect 12290 5920 12305 5935
rect 12345 5920 12360 5935
rect 12400 5920 12415 5935
rect 12455 5920 12470 5935
rect 12510 5920 12525 5935
rect 12565 5920 12580 5935
rect 18665 5930 18675 5950
rect 18695 5945 18760 5950
rect 20065 5950 20160 5960
rect 20065 5945 20130 5950
rect 18695 5930 18705 5945
rect 18665 5920 18705 5930
rect 20120 5930 20130 5945
rect 20150 5930 20160 5950
rect 20120 5920 20160 5930
rect 11165 5910 11260 5920
rect 11165 5890 11175 5910
rect 11195 5905 11260 5910
rect 12565 5910 12660 5920
rect 12565 5905 12630 5910
rect 11195 5890 11205 5905
rect 11165 5880 11205 5890
rect 12620 5890 12630 5905
rect 12650 5890 12660 5910
rect 12620 5880 12660 5890
rect 11632 4510 11668 4520
rect 11632 4490 11640 4510
rect 11660 4490 11668 4510
rect 11632 4480 11668 4490
rect 11752 4510 11788 4520
rect 11752 4490 11760 4510
rect 11780 4490 11788 4510
rect 11752 4480 11788 4490
rect 11872 4510 11908 4520
rect 11872 4490 11880 4510
rect 11900 4490 11908 4510
rect 11872 4480 11908 4490
rect 11570 4465 11610 4475
rect 11200 4450 11240 4460
rect 11200 4430 11210 4450
rect 11230 4430 11240 4450
rect 11460 4450 11500 4460
rect 11460 4430 11470 4450
rect 11490 4430 11500 4450
rect 11570 4445 11580 4465
rect 11600 4450 11610 4465
rect 11930 4465 11970 4475
rect 11930 4450 11940 4465
rect 11600 4445 11630 4450
rect 11570 4435 11630 4445
rect 11910 4445 11940 4450
rect 11960 4445 11970 4465
rect 11910 4435 11970 4445
rect 11200 4415 11300 4430
rect 11280 4403 11300 4415
rect 11340 4403 11360 4418
rect 11400 4415 11500 4430
rect 11610 4420 11630 4435
rect 11670 4420 11690 4435
rect 11730 4420 11750 4435
rect 11790 4420 11810 4435
rect 11850 4420 11870 4435
rect 11910 4420 11930 4435
rect 11400 4403 11420 4415
rect 12120 4395 12140 4410
rect 12180 4395 12200 4410
rect 12240 4395 12260 4410
rect 12300 4395 12320 4410
rect 12360 4395 12380 4410
rect 12420 4395 12440 4410
rect 12480 4395 12500 4410
rect 12540 4395 12560 4410
rect 11280 4325 11300 4340
rect 11340 4325 11360 4340
rect 11400 4325 11420 4340
rect 11610 4325 11630 4340
rect 11670 4330 11690 4340
rect 11730 4330 11750 4340
rect 11790 4330 11810 4340
rect 11850 4330 11870 4340
rect 11330 4315 11370 4325
rect 11670 4315 11870 4330
rect 11910 4325 11930 4340
rect 12120 4325 12140 4335
rect 12180 4325 12200 4335
rect 12240 4325 12260 4335
rect 12300 4325 12320 4335
rect 12360 4325 12380 4335
rect 12420 4325 12440 4335
rect 12480 4325 12500 4335
rect 12540 4325 12560 4335
rect 11330 4295 11340 4315
rect 11360 4295 11370 4315
rect 11330 4285 11370 4295
rect 11750 4310 11790 4315
rect 12120 4310 12560 4325
rect 11750 4290 11760 4310
rect 11780 4290 11790 4310
rect 11750 4280 11790 4290
rect 12203 4290 12211 4310
rect 12229 4290 12237 4310
rect 12203 4280 12237 4290
rect 11210 4200 11250 4210
rect 11210 4180 11220 4200
rect 11240 4180 11250 4200
rect 12500 4200 12540 4210
rect 12500 4180 12510 4200
rect 12530 4180 12540 4200
rect 11210 4165 11305 4180
rect 11290 4155 11305 4165
rect 11345 4155 11360 4170
rect 11400 4155 11415 4170
rect 11455 4155 11470 4170
rect 11510 4155 11525 4170
rect 11565 4155 11580 4170
rect 11620 4155 11635 4170
rect 11675 4155 11690 4170
rect 11730 4155 11745 4170
rect 11785 4155 11800 4170
rect 11840 4155 11855 4170
rect 11895 4155 11910 4170
rect 11950 4155 11965 4170
rect 12005 4155 12020 4170
rect 12060 4155 12075 4170
rect 12115 4155 12130 4170
rect 12170 4155 12185 4170
rect 12225 4155 12240 4170
rect 12280 4155 12295 4170
rect 12335 4155 12350 4170
rect 12390 4155 12405 4170
rect 12445 4165 12540 4180
rect 12445 4155 12460 4165
rect 11290 4090 11305 4105
rect 11345 4095 11360 4105
rect 11400 4095 11415 4105
rect 11455 4095 11470 4105
rect 11510 4095 11525 4105
rect 11565 4095 11580 4105
rect 11620 4095 11635 4105
rect 11675 4095 11690 4105
rect 11730 4095 11745 4105
rect 11785 4095 11800 4105
rect 11840 4095 11855 4105
rect 11895 4095 11910 4105
rect 11950 4095 11965 4105
rect 12005 4095 12020 4105
rect 12060 4095 12075 4105
rect 12115 4095 12130 4105
rect 12170 4095 12185 4105
rect 12225 4095 12240 4105
rect 12280 4095 12295 4105
rect 12335 4095 12350 4105
rect 12390 4095 12405 4105
rect 11345 4080 12405 4095
rect 12445 4090 12460 4105
rect 11362 4060 11370 4080
rect 11390 4060 11398 4080
rect 11362 4050 11398 4060
rect 11155 3895 11195 3905
rect 11155 3875 11165 3895
rect 11185 3875 11195 3895
rect 11271 3895 11303 3905
rect 11271 3875 11277 3895
rect 11294 3875 11303 3895
rect 11470 3895 11510 3905
rect 11470 3875 11480 3895
rect 11500 3875 11510 3895
rect 11690 3895 11730 3905
rect 11690 3875 11700 3895
rect 11720 3875 11730 3895
rect 11895 3895 11935 3905
rect 11895 3875 11905 3895
rect 11925 3875 11935 3895
rect 12011 3895 12043 3905
rect 12011 3875 12017 3895
rect 12034 3875 12043 3895
rect 12210 3895 12250 3905
rect 12210 3875 12220 3895
rect 12240 3875 12250 3895
rect 12430 3895 12470 3905
rect 12430 3875 12440 3895
rect 12460 3875 12470 3895
rect 12635 3895 12675 3905
rect 12635 3875 12645 3895
rect 12665 3875 12675 3895
rect 11155 3860 11250 3875
rect 11271 3865 11305 3875
rect 11235 3850 11250 3860
rect 11290 3850 11305 3865
rect 11345 3850 11360 3865
rect 11400 3850 11415 3865
rect 11455 3860 11525 3875
rect 11455 3850 11470 3860
rect 11510 3850 11525 3860
rect 11565 3850 11580 3865
rect 11620 3850 11635 3865
rect 11675 3860 11745 3875
rect 11675 3850 11690 3860
rect 11730 3850 11745 3860
rect 11785 3850 11800 3865
rect 11840 3860 11990 3875
rect 12011 3865 12045 3875
rect 11840 3850 11855 3860
rect 11975 3850 11990 3860
rect 12030 3850 12045 3865
rect 12085 3850 12100 3865
rect 12140 3850 12155 3865
rect 12195 3860 12265 3875
rect 12195 3850 12210 3860
rect 12250 3850 12265 3860
rect 12305 3850 12320 3865
rect 12360 3850 12375 3865
rect 12415 3860 12485 3875
rect 12415 3850 12430 3860
rect 12470 3850 12485 3860
rect 12525 3850 12540 3865
rect 12580 3860 12675 3875
rect 12580 3850 12595 3860
rect 11235 3785 11250 3800
rect 11290 3785 11305 3800
rect 11345 3790 11360 3800
rect 11400 3790 11415 3800
rect 11345 3785 11415 3790
rect 11455 3785 11470 3800
rect 11510 3785 11525 3800
rect 11565 3790 11580 3800
rect 11620 3790 11635 3800
rect 11565 3785 11635 3790
rect 11675 3785 11690 3800
rect 11730 3785 11745 3800
rect 11785 3785 11800 3800
rect 11840 3785 11855 3800
rect 11975 3785 11990 3800
rect 12030 3785 12045 3800
rect 12085 3790 12100 3800
rect 12140 3790 12155 3800
rect 12085 3785 12155 3790
rect 12195 3785 12210 3800
rect 12250 3785 12265 3800
rect 12305 3790 12320 3800
rect 12360 3790 12375 3800
rect 12305 3785 12375 3790
rect 12415 3785 12430 3800
rect 12470 3785 12485 3800
rect 12525 3785 12540 3800
rect 12580 3785 12595 3800
rect 11345 3775 11434 3785
rect 11565 3775 11654 3785
rect 11402 3755 11408 3775
rect 11425 3755 11434 3775
rect 11402 3745 11434 3755
rect 11622 3755 11628 3775
rect 11645 3755 11654 3775
rect 11622 3745 11654 3755
rect 11766 3775 11800 3785
rect 12085 3775 12174 3785
rect 12305 3775 12394 3785
rect 11766 3755 11775 3775
rect 11792 3755 11800 3775
rect 11766 3745 11800 3755
rect 12142 3755 12148 3775
rect 12165 3755 12174 3775
rect 12142 3745 12174 3755
rect 12362 3755 12368 3775
rect 12385 3755 12394 3775
rect 12362 3745 12394 3755
rect 12506 3775 12540 3785
rect 12506 3755 12515 3775
rect 12532 3755 12540 3775
rect 12506 3745 12540 3755
rect 11180 3620 11220 3630
rect 11180 3600 11190 3620
rect 11210 3600 11220 3620
rect 12580 3620 12620 3630
rect 12580 3600 12590 3620
rect 12610 3600 12620 3620
rect 26180 3620 26220 3630
rect 25905 3605 25945 3615
rect 10195 3585 10210 3600
rect 10250 3585 10265 3600
rect 10305 3585 10320 3600
rect 10360 3585 10375 3600
rect 10415 3585 10430 3600
rect 10470 3585 10485 3600
rect 10525 3585 10540 3600
rect 10580 3585 10595 3600
rect 10635 3585 10650 3600
rect 10690 3585 10705 3600
rect 10745 3585 10760 3600
rect 10800 3585 10815 3600
rect 11180 3585 11280 3600
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 3035 2930 3085 2945
rect 3125 2930 3175 2945
rect 3215 2930 3265 2945
rect 3305 2930 3355 2945
rect 3395 2930 3445 2945
rect 3485 2930 3535 2945
rect 3575 2930 3625 2945
rect 3665 2930 3715 2945
rect 3755 2930 3805 2945
rect 3845 2930 3895 2945
rect 3935 2930 3985 2945
rect 4025 2930 4075 2945
rect 4115 2930 4165 2945
rect 4205 2930 4255 2945
rect 4295 2930 4345 2945
rect 4385 2930 4435 2945
rect 4475 2930 4525 2945
rect 4565 2930 4615 2945
rect 4655 2930 4705 2945
rect 4745 2930 4795 2945
rect 4835 2930 4885 2945
rect 4925 2930 4975 2945
rect 11260 3575 11280 3585
rect 11320 3575 11340 3590
rect 11380 3575 11400 3590
rect 11440 3575 11460 3590
rect 11500 3575 11520 3590
rect 11560 3575 11580 3590
rect 11620 3575 11640 3590
rect 11680 3575 11700 3590
rect 11740 3575 11760 3590
rect 11800 3575 11820 3590
rect 11860 3575 11880 3590
rect 11920 3575 11940 3590
rect 11980 3575 12000 3590
rect 12040 3575 12060 3590
rect 12100 3575 12120 3590
rect 12160 3575 12180 3590
rect 12220 3575 12240 3590
rect 12280 3575 12300 3590
rect 12340 3575 12360 3590
rect 12400 3575 12420 3590
rect 12460 3575 12480 3590
rect 12520 3585 12620 3600
rect 12985 3585 13000 3600
rect 13040 3585 13055 3600
rect 13095 3585 13110 3600
rect 13150 3585 13165 3600
rect 13205 3585 13220 3600
rect 13260 3585 13275 3600
rect 13315 3585 13330 3600
rect 13370 3585 13385 3600
rect 13425 3585 13440 3600
rect 13480 3585 13495 3600
rect 13535 3585 13550 3600
rect 13590 3585 13605 3600
rect 25905 3585 25915 3605
rect 25935 3585 25945 3605
rect 26180 3600 26190 3620
rect 26210 3600 26220 3620
rect 27580 3620 27620 3630
rect 27580 3600 27590 3620
rect 27610 3600 27620 3620
rect 12520 3575 12540 3585
rect 11260 3160 11280 3175
rect 11320 3165 11340 3175
rect 11380 3165 11400 3175
rect 11440 3165 11460 3175
rect 11500 3165 11520 3175
rect 11560 3165 11580 3175
rect 11620 3165 11640 3175
rect 11680 3165 11700 3175
rect 11740 3165 11760 3175
rect 11800 3165 11820 3175
rect 11860 3165 11880 3175
rect 11920 3165 11940 3175
rect 11980 3165 12000 3175
rect 12040 3165 12060 3175
rect 12100 3165 12120 3175
rect 12160 3165 12180 3175
rect 12220 3165 12240 3175
rect 12280 3165 12300 3175
rect 12340 3165 12360 3175
rect 12400 3165 12420 3175
rect 12460 3165 12480 3175
rect 11320 3150 12480 3165
rect 12520 3160 12540 3175
rect 11823 3130 11831 3150
rect 11849 3130 11857 3150
rect 11823 3120 11857 3130
rect 25905 3575 25945 3585
rect 25980 3580 26000 3595
rect 26040 3580 26060 3595
rect 26180 3585 26280 3600
rect 25860 3550 25880 3565
rect 25920 3550 25940 3575
rect 25450 3340 25490 3350
rect 25450 3320 25460 3340
rect 25480 3320 25490 3340
rect 25710 3340 25750 3350
rect 25710 3320 25720 3340
rect 25740 3320 25750 3340
rect 25450 3305 25550 3320
rect 25530 3293 25550 3305
rect 25590 3293 25610 3308
rect 25650 3305 25750 3320
rect 25650 3293 25670 3305
rect 26260 3575 26280 3585
rect 26320 3575 26340 3590
rect 26380 3575 26400 3590
rect 26440 3575 26460 3590
rect 26500 3575 26520 3590
rect 26560 3575 26580 3590
rect 26620 3575 26640 3590
rect 26680 3575 26700 3590
rect 26740 3575 26760 3590
rect 26800 3575 26820 3590
rect 26860 3575 26880 3590
rect 26920 3575 26940 3590
rect 26980 3575 27000 3590
rect 27040 3575 27060 3590
rect 27100 3575 27120 3590
rect 27160 3575 27180 3590
rect 27220 3575 27240 3590
rect 27280 3575 27300 3590
rect 27340 3575 27360 3590
rect 27400 3575 27420 3590
rect 27460 3575 27480 3590
rect 27520 3585 27620 3600
rect 27520 3575 27540 3585
rect 25530 3215 25550 3230
rect 25590 3215 25610 3230
rect 25650 3215 25670 3230
rect 25860 3220 25880 3230
rect 25580 3205 25620 3215
rect 25580 3185 25590 3205
rect 25610 3185 25620 3205
rect 25580 3175 25620 3185
rect 25780 3205 25880 3220
rect 25920 3215 25940 3230
rect 25905 3205 25940 3215
rect 25780 3185 25790 3205
rect 25810 3185 25820 3205
rect 25780 3175 25820 3185
rect 25905 3185 25910 3205
rect 25930 3185 25940 3205
rect 25905 3175 25940 3185
rect 25980 3215 26000 3230
rect 26040 3220 26060 3230
rect 25980 3205 26015 3215
rect 26040 3205 26140 3220
rect 25980 3185 25990 3205
rect 26010 3185 26015 3205
rect 25980 3175 26015 3185
rect 26100 3185 26110 3205
rect 26130 3185 26140 3205
rect 26100 3175 26140 3185
rect 27930 3240 27945 3255
rect 27985 3240 28000 3255
rect 28040 3240 28055 3255
rect 28095 3240 28110 3255
rect 28150 3240 28165 3255
rect 28205 3240 28220 3255
rect 28260 3240 28275 3255
rect 28315 3240 28330 3255
rect 28370 3240 28385 3255
rect 28425 3240 28440 3255
rect 28480 3240 28495 3255
rect 28535 3240 28550 3255
rect 28590 3240 28605 3255
rect 28645 3240 28660 3255
rect 28700 3240 28715 3255
rect 28755 3240 28770 3255
rect 28810 3240 28825 3255
rect 28865 3240 28880 3255
rect 28920 3240 28935 3255
rect 28975 3240 28990 3255
rect 29030 3240 29045 3255
rect 29085 3240 29100 3255
rect 26260 3160 26280 3175
rect 26320 3165 26340 3175
rect 26380 3165 26400 3175
rect 26440 3165 26460 3175
rect 26500 3165 26520 3175
rect 26560 3165 26580 3175
rect 26620 3165 26640 3175
rect 26680 3165 26700 3175
rect 26740 3165 26760 3175
rect 26800 3165 26820 3175
rect 26860 3165 26880 3175
rect 26920 3165 26940 3175
rect 26980 3165 27000 3175
rect 27040 3165 27060 3175
rect 27100 3165 27120 3175
rect 27160 3165 27180 3175
rect 27220 3165 27240 3175
rect 27280 3165 27300 3175
rect 27340 3165 27360 3175
rect 27400 3165 27420 3175
rect 27460 3165 27480 3175
rect 10195 2975 10210 2985
rect 10115 2960 10210 2975
rect 10250 2975 10265 2985
rect 10305 2975 10320 2985
rect 10360 2975 10375 2985
rect 10415 2975 10430 2985
rect 10470 2975 10485 2985
rect 10525 2975 10540 2985
rect 10580 2975 10595 2985
rect 10635 2975 10650 2985
rect 10690 2975 10705 2985
rect 10745 2975 10760 2985
rect 10250 2960 10760 2975
rect 10800 2975 10815 2985
rect 12985 2975 13000 2985
rect 10800 2960 10895 2975
rect 10115 2940 10125 2960
rect 10145 2940 10155 2960
rect 10115 2930 10155 2940
rect 10653 2940 10661 2960
rect 10679 2940 10687 2960
rect 10653 2930 10687 2940
rect 10855 2940 10865 2960
rect 10885 2940 10895 2960
rect 12905 2960 13000 2975
rect 13040 2975 13055 2985
rect 13095 2975 13110 2985
rect 13150 2975 13165 2985
rect 13205 2975 13220 2985
rect 13260 2975 13275 2985
rect 13315 2975 13330 2985
rect 13370 2975 13385 2985
rect 13425 2975 13440 2985
rect 13480 2975 13495 2985
rect 13535 2975 13550 2985
rect 13040 2960 13550 2975
rect 13590 2975 13605 2985
rect 13590 2960 13685 2975
rect 10855 2930 10895 2940
rect 11180 2940 11220 2950
rect 11180 2920 11190 2940
rect 11210 2920 11220 2940
rect 12580 2940 12620 2950
rect 12580 2920 12590 2940
rect 12610 2920 12620 2940
rect 12905 2940 12915 2960
rect 12935 2940 12945 2960
rect 12905 2930 12945 2940
rect 13113 2940 13121 2960
rect 13139 2940 13147 2960
rect 13113 2930 13147 2940
rect 13645 2940 13655 2960
rect 13675 2940 13685 2960
rect 26320 3150 27480 3165
rect 27520 3160 27540 3175
rect 26823 3130 26831 3150
rect 26849 3130 26857 3150
rect 26823 3120 26857 3130
rect 26180 2940 26220 2950
rect 13645 2930 13685 2940
rect 11180 2905 11280 2920
rect 11260 2895 11280 2905
rect 11320 2895 11340 2910
rect 11380 2895 11400 2910
rect 11440 2895 11460 2910
rect 11500 2895 11520 2910
rect 11560 2895 11580 2910
rect 11620 2895 11640 2910
rect 11680 2895 11700 2910
rect 11740 2895 11760 2910
rect 11800 2895 11820 2910
rect 11860 2895 11880 2910
rect 11920 2895 11940 2910
rect 11980 2895 12000 2910
rect 12040 2895 12060 2910
rect 12100 2895 12120 2910
rect 12160 2895 12180 2910
rect 12220 2895 12240 2910
rect 12280 2895 12300 2910
rect 12340 2895 12360 2910
rect 12400 2895 12420 2910
rect 12460 2895 12480 2910
rect 12520 2905 12620 2920
rect 26180 2920 26190 2940
rect 26210 2920 26220 2940
rect 27580 2940 27620 2950
rect 27580 2920 27590 2940
rect 27610 2920 27620 2940
rect 27930 2930 27945 2940
rect 26180 2905 26280 2920
rect 12520 2895 12540 2905
rect 26260 2895 26280 2905
rect 26320 2895 26340 2910
rect 26380 2895 26400 2910
rect 26440 2895 26460 2910
rect 26500 2895 26520 2910
rect 26560 2895 26580 2910
rect 26620 2895 26640 2910
rect 26680 2895 26700 2910
rect 26740 2895 26760 2910
rect 26800 2895 26820 2910
rect 26860 2895 26880 2910
rect 26920 2895 26940 2910
rect 26980 2895 27000 2910
rect 27040 2895 27060 2910
rect 27100 2895 27120 2910
rect 27160 2895 27180 2910
rect 27220 2895 27240 2910
rect 27280 2895 27300 2910
rect 27340 2895 27360 2910
rect 27400 2895 27420 2910
rect 27460 2895 27480 2910
rect 27520 2905 27620 2920
rect 27850 2915 27945 2930
rect 27985 2930 28000 2940
rect 28040 2930 28055 2940
rect 28095 2930 28110 2940
rect 28150 2930 28165 2940
rect 28205 2930 28220 2940
rect 28260 2930 28275 2940
rect 28315 2930 28330 2940
rect 28370 2930 28385 2940
rect 28425 2930 28440 2940
rect 28480 2930 28495 2940
rect 28535 2930 28550 2940
rect 28590 2930 28605 2940
rect 28645 2930 28660 2940
rect 28700 2930 28715 2940
rect 28755 2930 28770 2940
rect 28810 2930 28825 2940
rect 28865 2930 28880 2940
rect 28920 2930 28935 2940
rect 28975 2930 28990 2940
rect 29030 2930 29045 2940
rect 27985 2915 29045 2930
rect 29085 2930 29100 2940
rect 29085 2915 29180 2930
rect 27520 2895 27540 2905
rect 27850 2895 27860 2915
rect 27880 2895 27890 2915
rect 3035 2815 3085 2830
rect 2995 2805 3085 2815
rect 3125 2820 3175 2830
rect 3215 2820 3265 2830
rect 3305 2820 3355 2830
rect 3395 2820 3445 2830
rect 3485 2820 3535 2830
rect 3575 2820 3625 2830
rect 3665 2820 3715 2830
rect 3755 2820 3805 2830
rect 3845 2820 3895 2830
rect 3935 2820 3985 2830
rect 4025 2820 4075 2830
rect 4115 2820 4165 2830
rect 4205 2820 4255 2830
rect 4295 2820 4345 2830
rect 4385 2820 4435 2830
rect 4475 2820 4525 2830
rect 4565 2820 4615 2830
rect 4655 2820 4705 2830
rect 4745 2820 4795 2830
rect 4835 2820 4885 2830
rect 3125 2805 4885 2820
rect 4925 2815 4975 2830
rect 4925 2805 5015 2815
rect 2995 2785 3005 2805
rect 3025 2800 3085 2805
rect 4925 2800 4985 2805
rect 3025 2785 3035 2800
rect 2995 2775 3035 2785
rect 4975 2785 4985 2800
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2730 3215 2745
rect 4795 2745 4835 2755
rect 4795 2730 4805 2745
rect 3205 2725 3265 2730
rect 3175 2715 3265 2725
rect 4745 2725 4805 2730
rect 4825 2725 4835 2745
rect 4745 2715 4835 2725
rect 3215 2700 3265 2715
rect 3305 2700 3355 2715
rect 3395 2700 3445 2715
rect 3485 2700 3535 2715
rect 3575 2700 3625 2715
rect 3665 2700 3715 2715
rect 3755 2700 3805 2715
rect 3845 2700 3895 2715
rect 3935 2700 3985 2715
rect 4025 2700 4075 2715
rect 4115 2700 4165 2715
rect 4205 2700 4255 2715
rect 4295 2700 4345 2715
rect 4385 2700 4435 2715
rect 4475 2700 4525 2715
rect 4565 2700 4615 2715
rect 4655 2700 4705 2715
rect 4745 2700 4795 2715
rect 10195 2655 10210 2670
rect 10250 2655 10265 2670
rect 10305 2655 10320 2670
rect 10360 2655 10375 2670
rect 10415 2655 10430 2670
rect 10470 2655 10485 2670
rect 10525 2655 10540 2670
rect 10580 2655 10595 2670
rect 10635 2655 10650 2670
rect 10690 2655 10705 2670
rect 10745 2655 10760 2670
rect 10800 2655 10815 2670
rect 3215 2385 3265 2400
rect 3305 2390 3355 2400
rect 3395 2390 3445 2400
rect 3485 2390 3535 2400
rect 3575 2390 3625 2400
rect 3665 2390 3715 2400
rect 3755 2390 3805 2400
rect 3845 2390 3895 2400
rect 3935 2390 3985 2400
rect 4025 2390 4075 2400
rect 4115 2390 4165 2400
rect 4205 2390 4255 2400
rect 4295 2390 4345 2400
rect 4385 2390 4435 2400
rect 4475 2390 4525 2400
rect 4565 2390 4615 2400
rect 4655 2390 4705 2400
rect 3305 2375 4705 2390
rect 4745 2385 4795 2400
rect 3355 2370 3395 2375
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 3355 2340 3395 2350
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 2605 2000 2620 2015
rect 2660 2000 2675 2015
rect 2785 2000 2805 2015
rect 2845 2000 2865 2015
rect 2905 2000 2925 2015
rect 2965 2000 2985 2015
rect 3025 2000 3045 2015
rect 3085 2000 3105 2015
rect 3145 2000 3165 2015
rect 3205 2000 3225 2015
rect 3265 2000 3285 2015
rect 3325 2000 3345 2015
rect 3385 2000 3405 2015
rect 3445 2000 3465 2015
rect 3505 2000 3525 2015
rect 3565 2000 3585 2015
rect 3625 2000 3645 2015
rect 3685 2000 3705 2015
rect 3745 2000 3765 2015
rect 3805 2000 3825 2015
rect 3865 2000 3885 2015
rect 3925 2000 3945 2015
rect 4065 2000 4085 2015
rect 4125 2000 4145 2015
rect 4185 2000 4205 2015
rect 4245 2000 4265 2015
rect 4305 2000 4325 2015
rect 4365 2000 4385 2015
rect 4425 2000 4445 2015
rect 4485 2000 4505 2015
rect 4545 2000 4565 2015
rect 4605 2000 4625 2015
rect 4665 2000 4685 2015
rect 4725 2000 4745 2015
rect 4785 2000 4805 2015
rect 4845 2000 4865 2015
rect 4905 2000 4925 2015
rect 4965 2000 4985 2015
rect 5025 2000 5045 2015
rect 5085 2000 5105 2015
rect 5145 2000 5165 2015
rect 5205 2000 5225 2015
rect 12985 2655 13000 2670
rect 13040 2655 13055 2670
rect 13095 2655 13110 2670
rect 13150 2655 13165 2670
rect 13205 2655 13220 2670
rect 13260 2655 13275 2670
rect 13315 2655 13330 2670
rect 13370 2655 13385 2670
rect 13425 2655 13440 2670
rect 13480 2655 13495 2670
rect 13535 2655 13550 2670
rect 13590 2655 13605 2670
rect 11260 2480 11280 2495
rect 11320 2485 11340 2495
rect 11380 2485 11400 2495
rect 11440 2485 11460 2495
rect 11500 2485 11520 2495
rect 11560 2485 11580 2495
rect 11620 2485 11640 2495
rect 11680 2485 11700 2495
rect 11740 2485 11760 2495
rect 11800 2485 11820 2495
rect 11860 2485 11880 2495
rect 11920 2485 11940 2495
rect 11980 2485 12000 2495
rect 12040 2485 12060 2495
rect 12100 2485 12120 2495
rect 12160 2485 12180 2495
rect 12220 2485 12240 2495
rect 12280 2485 12300 2495
rect 12340 2485 12360 2495
rect 12400 2485 12420 2495
rect 12460 2485 12480 2495
rect 11320 2470 12480 2485
rect 12520 2480 12540 2495
rect 10195 2445 10210 2455
rect 10115 2430 10210 2445
rect 10250 2445 10265 2455
rect 10305 2445 10320 2455
rect 10360 2445 10375 2455
rect 10415 2445 10430 2455
rect 10470 2445 10485 2455
rect 10525 2445 10540 2455
rect 10580 2445 10595 2455
rect 10635 2445 10650 2455
rect 10690 2445 10705 2455
rect 10745 2445 10760 2455
rect 10250 2430 10760 2445
rect 10800 2445 10815 2455
rect 11823 2450 11831 2470
rect 11849 2450 11857 2470
rect 10800 2430 10895 2445
rect 11823 2440 11857 2450
rect 12985 2445 13000 2455
rect 10115 2410 10125 2430
rect 10145 2410 10155 2430
rect 10115 2400 10155 2410
rect 10745 2395 10760 2430
rect 10855 2410 10865 2430
rect 10885 2410 10895 2430
rect 10855 2400 10895 2410
rect 12905 2430 13000 2445
rect 13040 2445 13055 2455
rect 13095 2445 13110 2455
rect 13150 2445 13165 2455
rect 13205 2445 13220 2455
rect 13260 2445 13275 2455
rect 13315 2445 13330 2455
rect 13370 2445 13385 2455
rect 13425 2445 13440 2455
rect 13480 2445 13495 2455
rect 13535 2445 13550 2455
rect 13040 2430 13550 2445
rect 13590 2445 13605 2455
rect 13590 2430 13685 2445
rect 12905 2410 12915 2430
rect 12935 2410 12945 2430
rect 12905 2400 12945 2410
rect 10745 2385 10805 2395
rect 10745 2365 10775 2385
rect 10795 2365 10805 2385
rect 13040 2380 13055 2430
rect 13645 2410 13655 2430
rect 13675 2410 13685 2430
rect 13645 2400 13685 2410
rect 10745 2355 10805 2365
rect 13025 2370 13065 2380
rect 10115 2310 10155 2320
rect 10115 2290 10125 2310
rect 10145 2290 10155 2310
rect 10745 2290 10760 2355
rect 13025 2350 13035 2370
rect 13055 2350 13065 2370
rect 13025 2340 13065 2350
rect 10855 2310 10895 2320
rect 10855 2290 10865 2310
rect 10885 2290 10895 2310
rect 10115 2275 10210 2290
rect 10195 2265 10210 2275
rect 10250 2275 10760 2290
rect 10250 2265 10265 2275
rect 10305 2265 10320 2275
rect 10360 2265 10375 2275
rect 10415 2265 10430 2275
rect 10470 2265 10485 2275
rect 10525 2265 10540 2275
rect 10580 2265 10595 2275
rect 10635 2265 10650 2275
rect 10690 2265 10705 2275
rect 10745 2265 10760 2275
rect 10800 2275 10895 2290
rect 12905 2310 12945 2320
rect 12905 2290 12915 2310
rect 12935 2290 12945 2310
rect 13040 2290 13055 2340
rect 13645 2310 13685 2320
rect 13645 2290 13655 2310
rect 13675 2290 13685 2310
rect 12905 2275 13000 2290
rect 10800 2265 10815 2275
rect 12985 2265 13000 2275
rect 13040 2275 13550 2290
rect 13040 2265 13055 2275
rect 13095 2265 13110 2275
rect 13150 2265 13165 2275
rect 13205 2265 13220 2275
rect 13260 2265 13275 2275
rect 13315 2265 13330 2275
rect 13370 2265 13385 2275
rect 13425 2265 13440 2275
rect 13480 2265 13495 2275
rect 13535 2265 13550 2275
rect 13590 2275 13685 2290
rect 13590 2265 13605 2275
rect 11828 2175 11862 2185
rect 11828 2155 11836 2175
rect 11854 2155 11862 2175
rect 11315 2130 11330 2145
rect 11370 2140 12430 2155
rect 11370 2130 11385 2140
rect 11425 2130 11440 2140
rect 11480 2130 11495 2140
rect 11535 2130 11550 2140
rect 11590 2130 11605 2140
rect 11645 2130 11660 2140
rect 11700 2130 11715 2140
rect 11755 2130 11770 2140
rect 11810 2130 11825 2140
rect 11865 2130 11880 2140
rect 11920 2130 11935 2140
rect 11975 2130 11990 2140
rect 12030 2130 12045 2140
rect 12085 2130 12100 2140
rect 12140 2130 12155 2140
rect 12195 2130 12210 2140
rect 12250 2130 12265 2140
rect 12305 2130 12320 2140
rect 12360 2130 12375 2140
rect 12415 2130 12430 2140
rect 12470 2130 12485 2145
rect 11315 1970 11330 1980
rect 10195 1950 10210 1965
rect 10250 1950 10265 1965
rect 10305 1950 10320 1965
rect 10360 1950 10375 1965
rect 10415 1950 10430 1965
rect 10470 1950 10485 1965
rect 10525 1950 10540 1965
rect 10580 1950 10595 1965
rect 10635 1950 10650 1965
rect 10690 1950 10705 1965
rect 10745 1950 10760 1965
rect 10800 1950 10815 1965
rect 11235 1955 11330 1970
rect 11370 1965 11385 1980
rect 11425 1965 11440 1980
rect 11480 1965 11495 1980
rect 11535 1965 11550 1980
rect 11590 1965 11605 1980
rect 11645 1965 11660 1980
rect 11700 1965 11715 1980
rect 11755 1965 11770 1980
rect 11810 1965 11825 1980
rect 11865 1965 11880 1980
rect 11920 1965 11935 1980
rect 11975 1965 11990 1980
rect 12030 1965 12045 1980
rect 12085 1965 12100 1980
rect 12140 1965 12155 1980
rect 12195 1965 12210 1980
rect 12250 1965 12265 1980
rect 12305 1965 12320 1980
rect 12360 1965 12375 1980
rect 12415 1965 12430 1980
rect 12470 1970 12485 1980
rect 12470 1955 12565 1970
rect 24720 2620 24735 2635
rect 24775 2620 24790 2635
rect 24830 2620 24845 2635
rect 24885 2620 24900 2635
rect 24940 2620 24955 2635
rect 24995 2620 25010 2635
rect 25050 2620 25065 2635
rect 25105 2620 25120 2635
rect 25160 2620 25175 2635
rect 25215 2620 25230 2635
rect 25270 2620 25285 2635
rect 25325 2620 25340 2635
rect 25380 2620 25395 2635
rect 25435 2620 25450 2635
rect 25490 2620 25505 2635
rect 25545 2620 25560 2635
rect 25600 2620 25615 2635
rect 25655 2620 25670 2635
rect 25710 2620 25725 2635
rect 25765 2620 25780 2635
rect 25820 2620 25835 2635
rect 25875 2620 25890 2635
rect 24720 2510 24735 2520
rect 24640 2495 24735 2510
rect 24775 2510 24790 2520
rect 24830 2510 24845 2520
rect 24885 2510 24900 2520
rect 24940 2510 24955 2520
rect 24995 2510 25010 2520
rect 25050 2510 25065 2520
rect 25105 2510 25120 2520
rect 25160 2510 25175 2520
rect 25215 2510 25230 2520
rect 25270 2510 25285 2520
rect 25325 2510 25340 2520
rect 25380 2510 25395 2520
rect 25435 2510 25450 2520
rect 25490 2510 25505 2520
rect 25545 2510 25560 2520
rect 25600 2510 25615 2520
rect 25655 2510 25670 2520
rect 25710 2510 25725 2520
rect 25765 2510 25780 2520
rect 25820 2510 25835 2520
rect 24775 2495 25835 2510
rect 25875 2510 25890 2520
rect 25875 2495 25970 2510
rect 27850 2885 27890 2895
rect 28058 2895 28066 2915
rect 28084 2895 28092 2915
rect 28058 2885 28092 2895
rect 29140 2895 29150 2915
rect 29170 2895 29180 2915
rect 29140 2885 29180 2895
rect 27930 2620 27945 2635
rect 27985 2620 28000 2635
rect 28040 2620 28055 2635
rect 28095 2620 28110 2635
rect 28150 2620 28165 2635
rect 28205 2620 28220 2635
rect 28260 2620 28275 2635
rect 28315 2620 28330 2635
rect 28370 2620 28385 2635
rect 28425 2620 28440 2635
rect 28480 2620 28495 2635
rect 28535 2620 28550 2635
rect 28590 2620 28605 2635
rect 28645 2620 28660 2635
rect 28700 2620 28715 2635
rect 28755 2620 28770 2635
rect 28810 2620 28825 2635
rect 28865 2620 28880 2635
rect 28920 2620 28935 2635
rect 28975 2620 28990 2635
rect 29030 2620 29045 2635
rect 29085 2620 29100 2635
rect 27930 2510 27945 2520
rect 27850 2495 27945 2510
rect 27985 2510 28000 2520
rect 28040 2510 28055 2520
rect 28095 2510 28110 2520
rect 28150 2510 28165 2520
rect 28205 2510 28220 2520
rect 28260 2510 28275 2520
rect 28315 2510 28330 2520
rect 28370 2510 28385 2520
rect 28425 2510 28440 2520
rect 28480 2510 28495 2520
rect 28535 2510 28550 2520
rect 28590 2510 28605 2520
rect 28645 2510 28660 2520
rect 28700 2510 28715 2520
rect 28755 2510 28770 2520
rect 28810 2510 28825 2520
rect 28865 2510 28880 2520
rect 28920 2510 28935 2520
rect 28975 2510 28990 2520
rect 29030 2510 29045 2520
rect 27985 2495 29045 2510
rect 29085 2510 29100 2520
rect 29085 2495 29180 2510
rect 24640 2475 24650 2495
rect 24670 2475 24680 2495
rect 24640 2465 24680 2475
rect 25820 2445 25835 2495
rect 25930 2475 25940 2495
rect 25960 2475 25970 2495
rect 26260 2480 26280 2495
rect 26320 2485 26340 2495
rect 26380 2485 26400 2495
rect 26440 2485 26460 2495
rect 26500 2485 26520 2495
rect 26560 2485 26580 2495
rect 26620 2485 26640 2495
rect 26680 2485 26700 2495
rect 26740 2485 26760 2495
rect 26800 2485 26820 2495
rect 26860 2485 26880 2495
rect 26920 2485 26940 2495
rect 26980 2485 27000 2495
rect 27040 2485 27060 2495
rect 27100 2485 27120 2495
rect 27160 2485 27180 2495
rect 27220 2485 27240 2495
rect 27280 2485 27300 2495
rect 27340 2485 27360 2495
rect 27400 2485 27420 2495
rect 27460 2485 27480 2495
rect 25930 2465 25970 2475
rect 26320 2470 27480 2485
rect 27520 2480 27540 2495
rect 27850 2475 27860 2495
rect 27880 2475 27890 2495
rect 26823 2450 26831 2470
rect 26849 2450 26857 2470
rect 27850 2465 27890 2475
rect 25813 2435 25847 2445
rect 26823 2440 26857 2450
rect 27985 2445 28000 2495
rect 29140 2475 29150 2495
rect 29170 2475 29180 2495
rect 29140 2465 29180 2475
rect 25813 2415 25821 2435
rect 25839 2415 25847 2435
rect 25813 2405 25847 2415
rect 27973 2435 28007 2445
rect 27973 2415 27981 2435
rect 27999 2415 28007 2435
rect 27973 2405 28007 2415
rect 25813 2275 25847 2285
rect 25813 2255 25821 2275
rect 25839 2255 25847 2275
rect 25813 2245 25847 2255
rect 27973 2275 28007 2285
rect 27973 2255 27981 2275
rect 27999 2255 28007 2275
rect 27973 2245 28007 2255
rect 24640 2215 24680 2225
rect 24640 2195 24650 2215
rect 24670 2195 24680 2215
rect 25820 2195 25835 2245
rect 25930 2215 25970 2225
rect 25930 2195 25940 2215
rect 25960 2195 25970 2215
rect 24640 2180 24735 2195
rect 24720 2170 24735 2180
rect 24775 2180 25835 2195
rect 24775 2170 24790 2180
rect 24830 2170 24845 2180
rect 24885 2170 24900 2180
rect 24940 2170 24955 2180
rect 24995 2170 25010 2180
rect 25050 2170 25065 2180
rect 25105 2170 25120 2180
rect 25160 2170 25175 2180
rect 25215 2170 25230 2180
rect 25270 2170 25285 2180
rect 25325 2170 25340 2180
rect 25380 2170 25395 2180
rect 25435 2170 25450 2180
rect 25490 2170 25505 2180
rect 25545 2170 25560 2180
rect 25600 2170 25615 2180
rect 25655 2170 25670 2180
rect 25710 2170 25725 2180
rect 25765 2170 25780 2180
rect 25820 2170 25835 2180
rect 25875 2180 25970 2195
rect 27850 2215 27890 2225
rect 27850 2195 27860 2215
rect 27880 2195 27890 2215
rect 27985 2195 28000 2245
rect 29140 2215 29180 2225
rect 29140 2195 29150 2215
rect 29170 2195 29180 2215
rect 27850 2180 27945 2195
rect 25875 2170 25890 2180
rect 27930 2170 27945 2180
rect 27985 2180 29045 2195
rect 27985 2170 28000 2180
rect 28040 2170 28055 2180
rect 28095 2170 28110 2180
rect 28150 2170 28165 2180
rect 28205 2170 28220 2180
rect 28260 2170 28275 2180
rect 28315 2170 28330 2180
rect 28370 2170 28385 2180
rect 28425 2170 28440 2180
rect 28480 2170 28495 2180
rect 28535 2170 28550 2180
rect 28590 2170 28605 2180
rect 28645 2170 28660 2180
rect 28700 2170 28715 2180
rect 28755 2170 28770 2180
rect 28810 2170 28825 2180
rect 28865 2170 28880 2180
rect 28920 2170 28935 2180
rect 28975 2170 28990 2180
rect 29030 2170 29045 2180
rect 29085 2180 29180 2195
rect 29085 2170 29100 2180
rect 26315 2130 26330 2145
rect 26370 2140 27430 2155
rect 26370 2130 26385 2140
rect 26425 2130 26440 2140
rect 26480 2130 26495 2140
rect 26535 2130 26550 2140
rect 26590 2130 26605 2140
rect 26645 2130 26660 2140
rect 26700 2130 26715 2140
rect 26755 2130 26770 2140
rect 26810 2130 26825 2140
rect 26865 2130 26880 2140
rect 26920 2130 26935 2140
rect 26975 2130 26990 2140
rect 27030 2130 27045 2140
rect 27085 2130 27100 2140
rect 27140 2130 27155 2140
rect 27195 2130 27210 2140
rect 27250 2130 27265 2140
rect 27305 2130 27320 2140
rect 27360 2130 27375 2140
rect 27415 2130 27430 2140
rect 27470 2130 27485 2145
rect 24720 2005 24735 2020
rect 24775 2005 24790 2020
rect 24830 2005 24845 2020
rect 24885 2005 24900 2020
rect 24940 2005 24955 2020
rect 24995 2005 25010 2020
rect 25050 2005 25065 2020
rect 25105 2005 25120 2020
rect 25160 2005 25175 2020
rect 25215 2005 25230 2020
rect 25270 2005 25285 2020
rect 25325 2005 25340 2020
rect 25380 2005 25395 2020
rect 25435 2005 25450 2020
rect 25490 2005 25505 2020
rect 25545 2005 25560 2020
rect 25600 2005 25615 2020
rect 25655 2005 25670 2020
rect 25710 2005 25725 2020
rect 25765 2005 25780 2020
rect 25820 2005 25835 2020
rect 25875 2005 25890 2020
rect 27930 2005 27945 2020
rect 27985 2005 28000 2020
rect 28040 2005 28055 2020
rect 28095 2005 28110 2020
rect 28150 2005 28165 2020
rect 28205 2005 28220 2020
rect 28260 2005 28275 2020
rect 28315 2005 28330 2020
rect 28370 2005 28385 2020
rect 28425 2005 28440 2020
rect 28480 2005 28495 2020
rect 28535 2005 28550 2020
rect 28590 2005 28605 2020
rect 28645 2005 28660 2020
rect 28700 2005 28715 2020
rect 28755 2005 28770 2020
rect 28810 2005 28825 2020
rect 28865 2005 28880 2020
rect 28920 2005 28935 2020
rect 28975 2005 28990 2020
rect 29030 2005 29045 2020
rect 29085 2005 29100 2020
rect 26315 1970 26330 1980
rect 11235 1935 11245 1955
rect 11265 1935 11275 1955
rect 11235 1925 11275 1935
rect 12525 1935 12535 1955
rect 12555 1935 12565 1955
rect 12985 1950 13000 1965
rect 13040 1950 13055 1965
rect 13095 1950 13110 1965
rect 13150 1950 13165 1965
rect 13205 1950 13220 1965
rect 13260 1950 13275 1965
rect 13315 1950 13330 1965
rect 13370 1950 13385 1965
rect 13425 1950 13440 1965
rect 13480 1950 13495 1965
rect 13535 1950 13550 1965
rect 13590 1950 13605 1965
rect 26235 1955 26330 1970
rect 26370 1965 26385 1980
rect 26425 1965 26440 1980
rect 26480 1965 26495 1980
rect 26535 1965 26550 1980
rect 26590 1965 26605 1980
rect 26645 1965 26660 1980
rect 26700 1965 26715 1980
rect 26755 1965 26770 1980
rect 26810 1965 26825 1980
rect 26865 1965 26880 1980
rect 26920 1965 26935 1980
rect 26975 1965 26990 1980
rect 27030 1965 27045 1980
rect 27085 1965 27100 1980
rect 27140 1965 27155 1980
rect 27195 1965 27210 1980
rect 27250 1965 27265 1980
rect 27305 1965 27320 1980
rect 27360 1965 27375 1980
rect 27415 1965 27430 1980
rect 27470 1970 27485 1980
rect 27470 1955 27565 1970
rect 12525 1925 12565 1935
rect 26235 1935 26245 1955
rect 26265 1935 26275 1955
rect 26235 1925 26275 1935
rect 27525 1935 27535 1955
rect 27555 1935 27565 1955
rect 27525 1925 27565 1935
rect 27950 1900 27990 1910
rect 2605 1890 2620 1900
rect 2660 1890 2675 1900
rect 2605 1875 2675 1890
rect 2785 1885 2805 1900
rect 2845 1885 2865 1900
rect 2905 1890 2925 1900
rect 2965 1890 2985 1900
rect 3025 1890 3045 1900
rect 3085 1890 3105 1900
rect 2765 1875 2805 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2765 1855 2775 1875
rect 2795 1855 2805 1875
rect 2765 1845 2805 1855
rect 2835 1875 2875 1885
rect 2905 1875 3105 1890
rect 3145 1890 3165 1900
rect 3205 1890 3225 1900
rect 3145 1875 3225 1890
rect 3265 1890 3285 1900
rect 3325 1890 3345 1900
rect 3385 1890 3405 1900
rect 3445 1890 3465 1900
rect 3265 1875 3465 1890
rect 3505 1890 3525 1900
rect 3565 1890 3585 1900
rect 3505 1875 3585 1890
rect 3625 1890 3645 1900
rect 3685 1890 3705 1900
rect 3745 1890 3765 1900
rect 3805 1890 3825 1900
rect 3625 1875 3825 1890
rect 3865 1885 3885 1900
rect 3925 1890 3945 1900
rect 4065 1890 4085 1900
rect 3855 1875 3895 1885
rect 3925 1875 4085 1890
rect 4125 1885 4145 1900
rect 4185 1890 4205 1900
rect 4245 1890 4265 1900
rect 4305 1890 4325 1900
rect 4365 1890 4385 1900
rect 4115 1875 4155 1885
rect 4185 1875 4385 1890
rect 4425 1890 4445 1900
rect 4485 1890 4505 1900
rect 4425 1875 4505 1890
rect 4545 1890 4565 1900
rect 4605 1890 4625 1900
rect 4665 1890 4685 1900
rect 4725 1890 4745 1900
rect 4545 1875 4745 1890
rect 4785 1890 4805 1900
rect 4845 1890 4865 1900
rect 4785 1875 4865 1890
rect 4905 1890 4925 1900
rect 4965 1890 4985 1900
rect 5025 1890 5045 1900
rect 5085 1890 5105 1900
rect 4905 1875 5105 1890
rect 5145 1885 5165 1900
rect 5205 1885 5225 1900
rect 5135 1875 5175 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1875
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5245 1885
rect 5205 1855 5215 1875
rect 5235 1855 5245 1875
rect 27950 1880 27960 1900
rect 27980 1880 27990 1900
rect 28360 1900 28400 1910
rect 28360 1880 28370 1900
rect 28390 1880 28400 1900
rect 27950 1865 28045 1880
rect 28030 1855 28045 1865
rect 28085 1855 28100 1870
rect 28140 1855 28155 1870
rect 28195 1855 28210 1870
rect 28250 1855 28265 1870
rect 28305 1865 28400 1880
rect 28305 1855 28320 1865
rect 5205 1845 5245 1855
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1720 3265 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1720 4785 1735
rect 3225 1705 3765 1720
rect 3205 1665 3225 1680
rect 3265 1665 3285 1705
rect 3325 1665 3345 1705
rect 3385 1665 3405 1680
rect 3445 1665 3465 1680
rect 3505 1665 3525 1705
rect 3565 1665 3585 1705
rect 3625 1665 3645 1680
rect 3685 1665 3705 1680
rect 3745 1665 3765 1705
rect 4245 1705 4785 1720
rect 11237 1710 11269 1720
rect 4245 1665 4265 1705
rect 4305 1665 4325 1680
rect 4365 1665 4385 1680
rect 4425 1665 4445 1705
rect 4485 1665 4505 1705
rect 4545 1665 4565 1680
rect 4605 1665 4625 1680
rect 4665 1665 4685 1705
rect 4725 1665 4745 1705
rect 10558 1700 10592 1710
rect 10558 1680 10566 1700
rect 10584 1680 10592 1700
rect 11237 1690 11243 1710
rect 11260 1690 11269 1710
rect 11457 1710 11489 1720
rect 11457 1690 11463 1710
rect 11480 1690 11489 1710
rect 11180 1680 11269 1690
rect 11400 1680 11489 1690
rect 11601 1710 11635 1720
rect 11601 1690 11610 1710
rect 11627 1690 11635 1710
rect 11867 1710 11899 1720
rect 11867 1695 11876 1710
rect 11601 1680 11635 1690
rect 11865 1690 11876 1695
rect 11893 1690 11899 1710
rect 12277 1710 12309 1720
rect 12277 1690 12283 1710
rect 12300 1690 12309 1710
rect 12497 1710 12529 1720
rect 12497 1690 12503 1710
rect 12520 1690 12529 1710
rect 11865 1680 11899 1690
rect 12220 1680 12309 1690
rect 12440 1680 12529 1690
rect 12641 1710 12675 1720
rect 26237 1710 26269 1720
rect 12641 1690 12650 1710
rect 12667 1690 12675 1710
rect 12641 1680 12675 1690
rect 13208 1700 13242 1710
rect 13208 1680 13216 1700
rect 13234 1680 13242 1700
rect 26237 1690 26243 1710
rect 26260 1690 26269 1710
rect 26457 1710 26489 1720
rect 26457 1690 26463 1710
rect 26480 1690 26489 1710
rect 26180 1680 26269 1690
rect 26400 1680 26489 1690
rect 26601 1710 26635 1720
rect 26601 1690 26610 1710
rect 26627 1690 26635 1710
rect 26867 1710 26899 1720
rect 26867 1695 26876 1710
rect 26601 1680 26635 1690
rect 26865 1690 26876 1695
rect 26893 1690 26899 1710
rect 27277 1710 27309 1720
rect 27277 1690 27283 1710
rect 27300 1690 27309 1710
rect 27497 1710 27529 1720
rect 27497 1690 27503 1710
rect 27520 1690 27529 1710
rect 26865 1680 26899 1690
rect 27220 1680 27309 1690
rect 27440 1680 27529 1690
rect 27641 1710 27675 1720
rect 27641 1690 27650 1710
rect 27667 1690 27675 1710
rect 28030 1690 28045 1705
rect 28085 1695 28100 1705
rect 28140 1695 28155 1705
rect 28195 1695 28210 1705
rect 28250 1695 28265 1705
rect 27641 1680 27675 1690
rect 28085 1685 28265 1695
rect 28305 1690 28320 1705
rect 28066 1680 28265 1685
rect 4785 1665 4805 1680
rect 10195 1655 10255 1670
rect 10295 1665 10655 1680
rect 10295 1655 10355 1665
rect 10395 1655 10455 1665
rect 10495 1655 10555 1665
rect 10595 1655 10655 1665
rect 10695 1655 10755 1670
rect 11070 1665 11085 1680
rect 11125 1665 11140 1680
rect 11180 1675 11250 1680
rect 11180 1665 11195 1675
rect 11235 1665 11250 1675
rect 11290 1665 11305 1680
rect 11345 1665 11360 1680
rect 11400 1675 11470 1680
rect 11400 1665 11415 1675
rect 11455 1665 11470 1675
rect 11510 1665 11525 1680
rect 11565 1665 11580 1680
rect 11620 1665 11635 1680
rect 11675 1665 11690 1680
rect 11810 1665 11825 1680
rect 11865 1665 11880 1680
rect 11920 1665 11935 1680
rect 11975 1665 11990 1680
rect 12110 1665 12125 1680
rect 12165 1665 12180 1680
rect 12220 1675 12290 1680
rect 12220 1665 12235 1675
rect 12275 1665 12290 1675
rect 12330 1665 12345 1680
rect 12385 1665 12400 1680
rect 12440 1675 12510 1680
rect 12440 1665 12455 1675
rect 12495 1665 12510 1675
rect 12550 1665 12565 1680
rect 12605 1665 12620 1680
rect 12660 1665 12675 1680
rect 12715 1665 12730 1680
rect 3205 1600 3225 1615
rect 3265 1600 3285 1615
rect 3325 1600 3345 1615
rect 3165 1590 3225 1600
rect 3165 1570 3175 1590
rect 3195 1575 3225 1590
rect 3385 1575 3405 1615
rect 3445 1575 3465 1615
rect 3505 1600 3525 1615
rect 3565 1600 3585 1615
rect 3625 1575 3645 1615
rect 3685 1575 3705 1615
rect 3745 1600 3765 1615
rect 4245 1600 4265 1615
rect 3195 1570 3705 1575
rect 3165 1560 3705 1570
rect 4305 1575 4325 1615
rect 4365 1575 4385 1615
rect 4425 1600 4445 1615
rect 4485 1600 4505 1615
rect 4545 1575 4565 1615
rect 4605 1575 4625 1615
rect 4665 1600 4685 1615
rect 4725 1600 4745 1615
rect 4785 1600 4805 1615
rect 4785 1590 4845 1600
rect 4785 1575 4815 1590
rect 4305 1570 4815 1575
rect 4835 1570 4845 1590
rect 4305 1560 4845 1570
rect 2925 1495 2965 1505
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1470 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1470 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1470 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1470 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1470 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1470 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 3765 1470 3805 1475
rect 4205 1495 4245 1505
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1470 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1470 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1470 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1470 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1470 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1470 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1470 5085 1475
rect 2875 1455 3375 1470
rect 3415 1455 3915 1470
rect 4095 1455 4595 1470
rect 4635 1455 5135 1470
rect 2875 1190 3375 1205
rect 3415 1190 3915 1205
rect 4095 1190 4595 1205
rect 4635 1190 5135 1205
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2985 1075 3985 1090
rect 4025 1075 5025 1090
rect 2985 960 3985 975
rect 4025 960 5025 975
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 13045 1655 13105 1670
rect 13145 1665 13505 1680
rect 13145 1655 13205 1665
rect 13245 1655 13305 1665
rect 13345 1655 13405 1665
rect 13445 1655 13505 1665
rect 13545 1655 13605 1670
rect 26070 1665 26085 1680
rect 26125 1665 26140 1680
rect 26180 1675 26250 1680
rect 26180 1665 26195 1675
rect 26235 1665 26250 1675
rect 26290 1665 26305 1680
rect 26345 1665 26360 1680
rect 26400 1675 26470 1680
rect 26400 1665 26415 1675
rect 26455 1665 26470 1675
rect 26510 1665 26525 1680
rect 26565 1665 26580 1680
rect 26620 1665 26635 1680
rect 26675 1665 26690 1680
rect 26810 1665 26825 1680
rect 26865 1665 26880 1680
rect 26920 1665 26935 1680
rect 26975 1665 26990 1680
rect 27110 1665 27125 1680
rect 27165 1665 27180 1680
rect 27220 1675 27290 1680
rect 27220 1665 27235 1675
rect 27275 1665 27290 1675
rect 27330 1665 27345 1680
rect 27385 1665 27400 1680
rect 27440 1675 27510 1680
rect 27440 1665 27455 1675
rect 27495 1665 27510 1675
rect 27550 1665 27565 1680
rect 27605 1665 27620 1680
rect 27660 1665 27675 1680
rect 27715 1665 27730 1680
rect 28066 1675 28100 1680
rect 11070 1505 11085 1515
rect 10990 1490 11085 1505
rect 11125 1500 11140 1515
rect 11180 1500 11195 1515
rect 11235 1500 11250 1515
rect 11290 1505 11305 1515
rect 11345 1505 11360 1515
rect 11106 1490 11140 1500
rect 11290 1490 11360 1505
rect 11400 1500 11415 1515
rect 11455 1500 11470 1515
rect 11510 1505 11525 1515
rect 11565 1505 11580 1515
rect 11510 1490 11580 1505
rect 11620 1500 11635 1515
rect 11675 1505 11690 1515
rect 11810 1505 11825 1515
rect 11675 1490 11825 1505
rect 11865 1500 11880 1515
rect 11920 1500 11935 1515
rect 11975 1505 11990 1515
rect 12110 1505 12125 1515
rect 11920 1490 11954 1500
rect 11975 1490 12125 1505
rect 12165 1500 12180 1515
rect 12220 1500 12235 1515
rect 12275 1500 12290 1515
rect 12330 1505 12345 1515
rect 12385 1505 12400 1515
rect 12146 1490 12180 1500
rect 12330 1490 12400 1505
rect 12440 1500 12455 1515
rect 12495 1500 12510 1515
rect 12550 1505 12565 1515
rect 12605 1505 12620 1515
rect 12550 1490 12620 1505
rect 12660 1500 12675 1515
rect 12715 1505 12730 1515
rect 12715 1490 12810 1505
rect 10990 1470 11000 1490
rect 11020 1470 11030 1490
rect 10990 1460 11030 1470
rect 11106 1470 11112 1490
rect 11129 1470 11138 1490
rect 11106 1460 11138 1470
rect 11305 1470 11315 1490
rect 11335 1470 11345 1490
rect 11305 1460 11345 1470
rect 11525 1470 11535 1490
rect 11555 1470 11565 1490
rect 11525 1460 11565 1470
rect 11730 1470 11740 1490
rect 11760 1470 11770 1490
rect 11730 1460 11770 1470
rect 11922 1470 11928 1490
rect 11945 1470 11954 1490
rect 11922 1460 11954 1470
rect 12030 1470 12040 1490
rect 12060 1470 12070 1490
rect 12030 1460 12070 1470
rect 12146 1470 12152 1490
rect 12169 1470 12178 1490
rect 12146 1460 12178 1470
rect 12345 1470 12355 1490
rect 12375 1470 12385 1490
rect 12345 1460 12385 1470
rect 12565 1470 12575 1490
rect 12595 1470 12605 1490
rect 12565 1460 12605 1470
rect 12770 1470 12780 1490
rect 12800 1470 12810 1490
rect 12770 1460 12810 1470
rect 12595 1245 12635 1255
rect 12595 1240 12605 1245
rect 11815 1230 11845 1240
rect 11815 1210 11820 1230
rect 11840 1210 11845 1230
rect 12510 1225 12605 1240
rect 12625 1225 12635 1245
rect 11245 1185 11260 1200
rect 11300 1195 12360 1210
rect 11300 1185 11315 1195
rect 11355 1185 11370 1195
rect 11410 1185 11425 1195
rect 11465 1185 11480 1195
rect 11520 1185 11535 1195
rect 11575 1185 11590 1195
rect 11630 1185 11645 1195
rect 11685 1185 11700 1195
rect 11740 1185 11755 1195
rect 11795 1185 11810 1195
rect 11850 1185 11865 1195
rect 11905 1185 11920 1195
rect 11960 1185 11975 1195
rect 12015 1185 12030 1195
rect 12070 1185 12085 1195
rect 12125 1185 12140 1195
rect 12180 1185 12195 1195
rect 12235 1185 12250 1195
rect 12290 1185 12305 1195
rect 12345 1185 12360 1195
rect 12400 1195 12470 1210
rect 12400 1185 12415 1195
rect 12455 1185 12470 1195
rect 12510 1185 12525 1225
rect 12595 1215 12635 1225
rect 12565 1185 12580 1200
rect 10195 945 10255 955
rect 10115 930 10255 945
rect 10295 940 10355 955
rect 10395 940 10455 955
rect 10495 940 10555 955
rect 10595 940 10655 955
rect 10695 945 10755 955
rect 10695 930 10835 945
rect 13045 945 13105 955
rect 10115 910 10125 930
rect 10145 910 10155 930
rect 2995 890 3085 905
rect 3035 880 3085 890
rect 3125 890 4885 905
rect 3125 880 3175 890
rect 3215 880 3265 890
rect 3305 880 3355 890
rect 3395 880 3445 890
rect 3485 880 3535 890
rect 3575 880 3625 890
rect 3665 880 3715 890
rect 3755 880 3805 890
rect 3845 880 3895 890
rect 3935 880 3985 890
rect 4025 880 4075 890
rect 4115 880 4165 890
rect 4205 880 4255 890
rect 4295 880 4345 890
rect 4385 880 4435 890
rect 4475 880 4525 890
rect 4565 880 4615 890
rect 4655 880 4705 890
rect 4745 880 4795 890
rect 4835 880 4885 890
rect 4925 890 5015 905
rect 10115 900 10155 910
rect 10795 910 10805 930
rect 10825 910 10835 930
rect 11245 920 11260 935
rect 11300 920 11315 935
rect 11355 920 11370 935
rect 11410 920 11425 935
rect 11465 920 11480 935
rect 11520 920 11535 935
rect 11575 920 11590 935
rect 11630 920 11645 935
rect 11685 920 11700 935
rect 11740 920 11755 935
rect 11795 920 11810 935
rect 11850 920 11865 935
rect 11905 920 11920 935
rect 11960 920 11975 935
rect 12015 920 12030 935
rect 12070 920 12085 935
rect 12125 920 12140 935
rect 12180 920 12195 935
rect 12235 920 12250 935
rect 12290 920 12305 935
rect 12345 920 12360 935
rect 12400 920 12415 935
rect 12455 920 12470 935
rect 12510 920 12525 935
rect 12565 920 12580 935
rect 12965 930 13105 945
rect 13145 940 13205 955
rect 13245 940 13305 955
rect 13345 940 13405 955
rect 13445 940 13505 955
rect 13545 945 13605 955
rect 13545 930 13685 945
rect 10795 900 10835 910
rect 11165 910 11260 920
rect 11165 890 11175 910
rect 11195 905 11260 910
rect 12565 910 12660 920
rect 12565 905 12630 910
rect 11195 890 11205 905
rect 4925 880 4975 890
rect 11165 880 11205 890
rect 12620 890 12630 905
rect 12650 890 12660 910
rect 12965 910 12975 930
rect 12995 910 13005 930
rect 12965 900 13005 910
rect 13645 910 13655 930
rect 13675 910 13685 930
rect 28066 1655 28071 1675
rect 28091 1670 28100 1675
rect 28091 1655 28098 1670
rect 28066 1645 28098 1655
rect 27971 1565 28003 1575
rect 27971 1545 27976 1565
rect 27996 1550 28003 1565
rect 28347 1565 28379 1575
rect 28347 1550 28354 1565
rect 27996 1545 28005 1550
rect 27971 1535 28005 1545
rect 28345 1545 28354 1550
rect 28374 1545 28379 1565
rect 28345 1535 28379 1545
rect 27935 1520 27950 1535
rect 27990 1520 28005 1535
rect 28045 1520 28060 1535
rect 28100 1520 28115 1535
rect 28235 1520 28250 1535
rect 28290 1520 28305 1535
rect 28345 1520 28360 1535
rect 28400 1520 28415 1535
rect 26070 1505 26085 1515
rect 25990 1490 26085 1505
rect 26125 1500 26140 1515
rect 26180 1500 26195 1515
rect 26235 1500 26250 1515
rect 26290 1505 26305 1515
rect 26345 1505 26360 1515
rect 26106 1490 26140 1500
rect 26290 1490 26360 1505
rect 26400 1500 26415 1515
rect 26455 1500 26470 1515
rect 26510 1505 26525 1515
rect 26565 1505 26580 1515
rect 26510 1490 26580 1505
rect 26620 1500 26635 1515
rect 26675 1505 26690 1515
rect 26810 1505 26825 1515
rect 26675 1490 26825 1505
rect 26865 1500 26880 1515
rect 26920 1500 26935 1515
rect 26975 1505 26990 1515
rect 27110 1505 27125 1515
rect 26920 1490 26954 1500
rect 26975 1490 27125 1505
rect 27165 1500 27180 1515
rect 27220 1500 27235 1515
rect 27275 1500 27290 1515
rect 27330 1505 27345 1515
rect 27385 1505 27400 1515
rect 27146 1490 27180 1500
rect 27330 1490 27400 1505
rect 27440 1500 27455 1515
rect 27495 1500 27510 1515
rect 27550 1505 27565 1515
rect 27605 1505 27620 1515
rect 27550 1490 27620 1505
rect 27660 1500 27675 1515
rect 27715 1505 27730 1515
rect 27715 1490 27810 1505
rect 25990 1470 26000 1490
rect 26020 1470 26030 1490
rect 25990 1460 26030 1470
rect 26106 1470 26112 1490
rect 26129 1470 26138 1490
rect 26106 1460 26138 1470
rect 26305 1470 26315 1490
rect 26335 1470 26345 1490
rect 26305 1460 26345 1470
rect 26525 1470 26535 1490
rect 26555 1470 26565 1490
rect 26525 1460 26565 1470
rect 26730 1470 26740 1490
rect 26760 1470 26770 1490
rect 26730 1460 26770 1470
rect 26922 1470 26928 1490
rect 26945 1470 26954 1490
rect 26922 1460 26954 1470
rect 27030 1470 27040 1490
rect 27060 1470 27070 1490
rect 27030 1460 27070 1470
rect 27146 1470 27152 1490
rect 27169 1470 27178 1490
rect 27146 1460 27178 1470
rect 27345 1470 27355 1490
rect 27375 1470 27385 1490
rect 27345 1460 27385 1470
rect 27565 1470 27575 1490
rect 27595 1470 27605 1490
rect 27565 1460 27605 1470
rect 27770 1470 27780 1490
rect 27800 1470 27810 1490
rect 27770 1460 27810 1470
rect 27935 1360 27950 1370
rect 27855 1345 27950 1360
rect 27990 1355 28005 1370
rect 28045 1355 28060 1370
rect 28026 1345 28060 1355
rect 28100 1360 28115 1370
rect 28235 1360 28250 1370
rect 28100 1345 28250 1360
rect 28290 1355 28305 1370
rect 28345 1355 28360 1370
rect 28400 1360 28415 1370
rect 28290 1345 28324 1355
rect 28400 1345 28495 1360
rect 27855 1325 27865 1345
rect 27885 1325 27895 1345
rect 27855 1315 27895 1325
rect 28026 1325 28033 1345
rect 28053 1340 28060 1345
rect 28053 1325 28058 1340
rect 28026 1315 28058 1325
rect 28155 1325 28165 1345
rect 28185 1325 28195 1345
rect 28290 1340 28297 1345
rect 28155 1315 28195 1325
rect 28292 1325 28297 1340
rect 28317 1325 28324 1345
rect 28292 1315 28324 1325
rect 28455 1325 28465 1345
rect 28485 1325 28495 1345
rect 28455 1315 28495 1325
rect 27595 1285 27635 1295
rect 27595 1280 27605 1285
rect 26815 1270 26845 1280
rect 26815 1250 26820 1270
rect 26840 1250 26845 1270
rect 27510 1265 27605 1280
rect 27625 1265 27635 1285
rect 26245 1225 26260 1240
rect 26300 1235 27360 1250
rect 26300 1225 26315 1235
rect 26355 1225 26370 1235
rect 26410 1225 26425 1235
rect 26465 1225 26480 1235
rect 26520 1225 26535 1235
rect 26575 1225 26590 1235
rect 26630 1225 26645 1235
rect 26685 1225 26700 1235
rect 26740 1225 26755 1235
rect 26795 1225 26810 1235
rect 26850 1225 26865 1235
rect 26905 1225 26920 1235
rect 26960 1225 26975 1235
rect 27015 1225 27030 1235
rect 27070 1225 27085 1235
rect 27125 1225 27140 1235
rect 27180 1225 27195 1235
rect 27235 1225 27250 1235
rect 27290 1225 27305 1235
rect 27345 1225 27360 1235
rect 27400 1235 27470 1250
rect 27400 1225 27415 1235
rect 27455 1225 27470 1235
rect 27510 1225 27525 1265
rect 27595 1255 27635 1265
rect 27565 1225 27580 1240
rect 28085 1180 28100 1195
rect 28140 1180 28155 1195
rect 28195 1180 28210 1195
rect 28250 1180 28265 1195
rect 28085 1020 28100 1030
rect 28005 1005 28100 1020
rect 28140 1020 28155 1030
rect 28195 1020 28210 1030
rect 28140 1015 28210 1020
rect 28250 1020 28265 1030
rect 28140 1005 28225 1015
rect 28250 1005 28345 1020
rect 28005 985 28015 1005
rect 28035 985 28045 1005
rect 28005 975 28045 985
rect 28185 985 28195 1005
rect 28215 985 28225 1005
rect 28185 975 28225 985
rect 28305 985 28315 1005
rect 28335 985 28345 1005
rect 28305 975 28345 985
rect 26245 960 26260 975
rect 26300 960 26315 975
rect 26355 960 26370 975
rect 26410 960 26425 975
rect 26465 960 26480 975
rect 26520 960 26535 975
rect 26575 960 26590 975
rect 26630 960 26645 975
rect 26685 960 26700 975
rect 26740 960 26755 975
rect 26795 960 26810 975
rect 26850 960 26865 975
rect 26905 960 26920 975
rect 26960 960 26975 975
rect 27015 960 27030 975
rect 27070 960 27085 975
rect 27125 960 27140 975
rect 27180 960 27195 975
rect 27235 960 27250 975
rect 27290 960 27305 975
rect 27345 960 27360 975
rect 27400 960 27415 975
rect 27455 960 27470 975
rect 27510 960 27525 975
rect 27565 960 27580 975
rect 26165 950 26260 960
rect 26165 930 26175 950
rect 26195 945 26260 950
rect 27565 950 27660 960
rect 27565 945 27630 950
rect 26195 930 26205 945
rect 26165 920 26205 930
rect 27620 930 27630 945
rect 27650 930 27660 950
rect 27620 920 27660 930
rect 13645 900 13685 910
rect 12620 880 12660 890
rect 11305 790 11345 800
rect 3035 765 3085 780
rect 3125 755 3175 780
rect 3215 765 3265 780
rect 3305 765 3355 780
rect 3395 765 3445 780
rect 3485 765 3535 780
rect 3575 765 3625 780
rect 3665 765 3715 780
rect 3755 765 3805 780
rect 3845 765 3895 780
rect 3935 765 3985 780
rect 4025 765 4075 780
rect 4115 765 4165 780
rect 4205 765 4255 780
rect 4295 765 4345 780
rect 4385 765 4435 780
rect 4475 765 4525 780
rect 4565 765 4615 780
rect 4655 765 4705 780
rect 4745 765 4795 780
rect 4835 765 4885 780
rect 4925 765 4975 780
rect 11305 770 11315 790
rect 11335 770 11345 790
rect 11305 760 11345 770
rect 11375 790 11415 800
rect 11375 770 11385 790
rect 11405 770 11415 790
rect 11375 760 11415 770
rect 11445 790 11485 800
rect 11445 770 11455 790
rect 11475 770 11485 790
rect 11935 795 11975 805
rect 11935 775 11945 795
rect 11965 775 11975 795
rect 12155 795 12195 805
rect 12155 775 12165 795
rect 12185 775 12195 795
rect 12375 795 12415 805
rect 12375 775 12385 795
rect 12405 775 12415 795
rect 11445 760 11485 770
rect 11920 760 12485 775
rect 3125 750 3140 755
rect 3130 735 3140 750
rect 3160 750 3175 755
rect 3160 735 3170 750
rect 11300 745 11490 760
rect 11920 750 11935 760
rect 11975 750 11990 760
rect 12030 750 12045 760
rect 12085 750 12100 760
rect 12140 750 12155 760
rect 12195 750 12210 760
rect 12250 750 12265 760
rect 12305 750 12320 760
rect 12360 750 12375 760
rect 12415 750 12430 760
rect 12470 750 12485 760
rect 12525 750 12540 765
rect 3130 725 3170 735
rect 11920 690 11935 700
rect 11840 675 11935 690
rect 11975 685 11990 700
rect 12030 685 12045 700
rect 12085 685 12100 700
rect 12140 685 12155 700
rect 12195 685 12210 700
rect 12250 685 12265 700
rect 12305 685 12320 700
rect 12360 685 12375 700
rect 12415 685 12430 700
rect 12470 685 12485 700
rect 12525 690 12540 700
rect 12525 675 12620 690
rect 11840 655 11850 675
rect 11870 655 11880 675
rect 11840 645 11880 655
rect 12580 655 12590 675
rect 12610 655 12620 675
rect 12580 645 12620 655
rect 11300 630 11490 645
rect 11180 -1380 11220 -1370
rect 10905 -1395 10945 -1385
rect 10905 -1415 10915 -1395
rect 10935 -1415 10945 -1395
rect 11180 -1400 11190 -1380
rect 11210 -1400 11220 -1380
rect 12580 -1380 12620 -1370
rect 12580 -1400 12590 -1380
rect 12610 -1400 12620 -1380
rect 10905 -1425 10945 -1415
rect 10980 -1420 11000 -1405
rect 11040 -1420 11060 -1405
rect 11180 -1415 11280 -1400
rect 10860 -1450 10880 -1435
rect 10920 -1450 10940 -1425
rect 10450 -1660 10490 -1650
rect 10450 -1680 10460 -1660
rect 10480 -1680 10490 -1660
rect 10710 -1660 10750 -1650
rect 10710 -1680 10720 -1660
rect 10740 -1680 10750 -1660
rect 10450 -1695 10550 -1680
rect 10530 -1707 10550 -1695
rect 10590 -1707 10610 -1692
rect 10650 -1695 10750 -1680
rect 10650 -1707 10670 -1695
rect 11260 -1425 11280 -1415
rect 11320 -1425 11340 -1410
rect 11380 -1425 11400 -1410
rect 11440 -1425 11460 -1410
rect 11500 -1425 11520 -1410
rect 11560 -1425 11580 -1410
rect 11620 -1425 11640 -1410
rect 11680 -1425 11700 -1410
rect 11740 -1425 11760 -1410
rect 11800 -1425 11820 -1410
rect 11860 -1425 11880 -1410
rect 11920 -1425 11940 -1410
rect 11980 -1425 12000 -1410
rect 12040 -1425 12060 -1410
rect 12100 -1425 12120 -1410
rect 12160 -1425 12180 -1410
rect 12220 -1425 12240 -1410
rect 12280 -1425 12300 -1410
rect 12340 -1425 12360 -1410
rect 12400 -1425 12420 -1410
rect 12460 -1425 12480 -1410
rect 12520 -1415 12620 -1400
rect 12520 -1425 12540 -1415
rect 10530 -1785 10550 -1770
rect 10590 -1785 10610 -1770
rect 10650 -1785 10670 -1770
rect 10860 -1780 10880 -1770
rect 10580 -1795 10620 -1785
rect 10580 -1815 10590 -1795
rect 10610 -1815 10620 -1795
rect 10580 -1825 10620 -1815
rect 10780 -1795 10880 -1780
rect 10920 -1785 10940 -1770
rect 10905 -1795 10940 -1785
rect 10780 -1815 10790 -1795
rect 10810 -1815 10820 -1795
rect 10780 -1825 10820 -1815
rect 10905 -1815 10910 -1795
rect 10930 -1815 10940 -1795
rect 10905 -1825 10940 -1815
rect 10980 -1785 11000 -1770
rect 11040 -1780 11060 -1770
rect 10980 -1795 11015 -1785
rect 11040 -1795 11140 -1780
rect 10980 -1815 10990 -1795
rect 11010 -1815 11015 -1795
rect 10980 -1825 11015 -1815
rect 11100 -1815 11110 -1795
rect 11130 -1815 11140 -1795
rect 11100 -1825 11140 -1815
rect 11260 -1840 11280 -1825
rect 11320 -1835 11340 -1825
rect 11380 -1835 11400 -1825
rect 11440 -1835 11460 -1825
rect 11500 -1835 11520 -1825
rect 11560 -1835 11580 -1825
rect 11620 -1835 11640 -1825
rect 11680 -1835 11700 -1825
rect 11740 -1835 11760 -1825
rect 11800 -1835 11820 -1825
rect 11860 -1835 11880 -1825
rect 11920 -1835 11940 -1825
rect 11980 -1835 12000 -1825
rect 12040 -1835 12060 -1825
rect 12100 -1835 12120 -1825
rect 12160 -1835 12180 -1825
rect 12220 -1835 12240 -1825
rect 12280 -1835 12300 -1825
rect 12340 -1835 12360 -1825
rect 12400 -1835 12420 -1825
rect 12460 -1835 12480 -1825
rect 11320 -1850 12480 -1835
rect 12520 -1840 12540 -1825
rect 11823 -1870 11831 -1850
rect 11849 -1870 11857 -1850
rect 11823 -1880 11857 -1870
rect 12935 -2015 12950 -2000
rect 12990 -2015 13005 -2000
rect 13045 -2015 13060 -2000
rect 13100 -2015 13115 -2000
rect 13155 -2015 13170 -2000
rect 13210 -2015 13225 -2000
rect 13265 -2015 13280 -2000
rect 13320 -2015 13335 -2000
rect 13375 -2015 13390 -2000
rect 13430 -2015 13445 -2000
rect 13485 -2015 13500 -2000
rect 13540 -2015 13555 -2000
rect 13595 -2015 13610 -2000
rect 13650 -2015 13665 -2000
rect 13705 -2015 13720 -2000
rect 13760 -2015 13775 -2000
rect 13815 -2015 13830 -2000
rect 13870 -2015 13885 -2000
rect 13925 -2015 13940 -2000
rect 13980 -2015 13995 -2000
rect 14035 -2015 14050 -2000
rect 14090 -2015 14105 -2000
rect 11180 -2060 11220 -2050
rect 11180 -2080 11190 -2060
rect 11210 -2080 11220 -2060
rect 12580 -2060 12620 -2050
rect 12580 -2080 12590 -2060
rect 12610 -2080 12620 -2060
rect 11180 -2095 11280 -2080
rect 11260 -2105 11280 -2095
rect 11320 -2105 11340 -2090
rect 11380 -2105 11400 -2090
rect 11440 -2105 11460 -2090
rect 11500 -2105 11520 -2090
rect 11560 -2105 11580 -2090
rect 11620 -2105 11640 -2090
rect 11680 -2105 11700 -2090
rect 11740 -2105 11760 -2090
rect 11800 -2105 11820 -2090
rect 11860 -2105 11880 -2090
rect 11920 -2105 11940 -2090
rect 11980 -2105 12000 -2090
rect 12040 -2105 12060 -2090
rect 12100 -2105 12120 -2090
rect 12160 -2105 12180 -2090
rect 12220 -2105 12240 -2090
rect 12280 -2105 12300 -2090
rect 12340 -2105 12360 -2090
rect 12400 -2105 12420 -2090
rect 12460 -2105 12480 -2090
rect 12520 -2095 12620 -2080
rect 12520 -2105 12540 -2095
rect 12935 -2325 12950 -2315
rect 12855 -2340 12950 -2325
rect 12990 -2325 13005 -2315
rect 13045 -2325 13060 -2315
rect 13100 -2325 13115 -2315
rect 13155 -2325 13170 -2315
rect 13210 -2325 13225 -2315
rect 13265 -2325 13280 -2315
rect 13320 -2325 13335 -2315
rect 13375 -2325 13390 -2315
rect 13430 -2325 13445 -2315
rect 13485 -2325 13500 -2315
rect 13540 -2325 13555 -2315
rect 13595 -2325 13610 -2315
rect 13650 -2325 13665 -2315
rect 13705 -2325 13720 -2315
rect 13760 -2325 13775 -2315
rect 13815 -2325 13830 -2315
rect 13870 -2325 13885 -2315
rect 13925 -2325 13940 -2315
rect 13980 -2325 13995 -2315
rect 14035 -2325 14050 -2315
rect 12990 -2340 14050 -2325
rect 14090 -2325 14105 -2315
rect 14090 -2340 14185 -2325
rect 12855 -2360 12865 -2340
rect 12885 -2360 12895 -2340
rect 12855 -2370 12895 -2360
rect 13063 -2360 13071 -2340
rect 13089 -2360 13097 -2340
rect 13063 -2370 13097 -2360
rect 14145 -2360 14155 -2340
rect 14175 -2360 14185 -2340
rect 14145 -2370 14185 -2360
rect 12935 -2445 12950 -2430
rect 12990 -2445 13005 -2430
rect 13045 -2445 13060 -2430
rect 13100 -2445 13115 -2430
rect 13155 -2445 13170 -2430
rect 13210 -2445 13225 -2430
rect 13265 -2445 13280 -2430
rect 13320 -2445 13335 -2430
rect 13375 -2445 13390 -2430
rect 13430 -2445 13445 -2430
rect 13485 -2445 13500 -2430
rect 13540 -2445 13555 -2430
rect 13595 -2445 13610 -2430
rect 13650 -2445 13665 -2430
rect 13705 -2445 13720 -2430
rect 13760 -2445 13775 -2430
rect 13815 -2445 13830 -2430
rect 13870 -2445 13885 -2430
rect 13925 -2445 13940 -2430
rect 13980 -2445 13995 -2430
rect 14035 -2445 14050 -2430
rect 14090 -2445 14105 -2430
rect 11260 -2520 11280 -2505
rect 11320 -2515 11340 -2505
rect 11380 -2515 11400 -2505
rect 11440 -2515 11460 -2505
rect 11500 -2515 11520 -2505
rect 11560 -2515 11580 -2505
rect 11620 -2515 11640 -2505
rect 11680 -2515 11700 -2505
rect 11740 -2515 11760 -2505
rect 11800 -2515 11820 -2505
rect 11860 -2515 11880 -2505
rect 11920 -2515 11940 -2505
rect 11980 -2515 12000 -2505
rect 12040 -2515 12060 -2505
rect 12100 -2515 12120 -2505
rect 12160 -2515 12180 -2505
rect 12220 -2515 12240 -2505
rect 12280 -2515 12300 -2505
rect 12340 -2515 12360 -2505
rect 12400 -2515 12420 -2505
rect 12460 -2515 12480 -2505
rect 11320 -2530 12480 -2515
rect 12520 -2520 12540 -2505
rect 11823 -2550 11831 -2530
rect 11849 -2550 11857 -2530
rect 11823 -2560 11857 -2550
rect 12935 -2555 12950 -2545
rect 12855 -2570 12950 -2555
rect 12990 -2555 13005 -2545
rect 13045 -2555 13060 -2545
rect 13100 -2555 13115 -2545
rect 13155 -2555 13170 -2545
rect 13210 -2555 13225 -2545
rect 13265 -2555 13280 -2545
rect 13320 -2555 13335 -2545
rect 13375 -2555 13390 -2545
rect 13430 -2555 13445 -2545
rect 13485 -2555 13500 -2545
rect 13540 -2555 13555 -2545
rect 13595 -2555 13610 -2545
rect 13650 -2555 13665 -2545
rect 13705 -2555 13720 -2545
rect 13760 -2555 13775 -2545
rect 13815 -2555 13830 -2545
rect 13870 -2555 13885 -2545
rect 13925 -2555 13940 -2545
rect 13980 -2555 13995 -2545
rect 14035 -2555 14050 -2545
rect 12990 -2570 14050 -2555
rect 14090 -2555 14105 -2545
rect 14090 -2570 14185 -2555
rect 12855 -2590 12865 -2570
rect 12885 -2590 12895 -2570
rect 12855 -2600 12895 -2590
rect 12990 -2620 13005 -2570
rect 14145 -2590 14155 -2570
rect 14175 -2590 14185 -2570
rect 14145 -2600 14185 -2590
rect 12975 -2630 13015 -2620
rect 12975 -2650 12985 -2630
rect 13005 -2650 13015 -2630
rect 12975 -2660 13015 -2650
rect 12855 -2690 12895 -2680
rect 12855 -2710 12865 -2690
rect 12885 -2710 12895 -2690
rect 12990 -2710 13005 -2660
rect 14145 -2690 14185 -2680
rect 14145 -2710 14155 -2690
rect 14175 -2710 14185 -2690
rect 12855 -2725 12950 -2710
rect 12935 -2735 12950 -2725
rect 12990 -2725 14050 -2710
rect 12990 -2735 13005 -2725
rect 13045 -2735 13060 -2725
rect 13100 -2735 13115 -2725
rect 13155 -2735 13170 -2725
rect 13210 -2735 13225 -2725
rect 13265 -2735 13280 -2725
rect 13320 -2735 13335 -2725
rect 13375 -2735 13390 -2725
rect 13430 -2735 13445 -2725
rect 13485 -2735 13500 -2725
rect 13540 -2735 13555 -2725
rect 13595 -2735 13610 -2725
rect 13650 -2735 13665 -2725
rect 13705 -2735 13720 -2725
rect 13760 -2735 13775 -2725
rect 13815 -2735 13830 -2725
rect 13870 -2735 13885 -2725
rect 13925 -2735 13940 -2725
rect 13980 -2735 13995 -2725
rect 14035 -2735 14050 -2725
rect 14090 -2725 14185 -2710
rect 14090 -2735 14105 -2725
rect 11315 -2870 11330 -2855
rect 11370 -2860 12430 -2845
rect 11370 -2870 11385 -2860
rect 11425 -2870 11440 -2860
rect 11480 -2870 11495 -2860
rect 11535 -2870 11550 -2860
rect 11590 -2870 11605 -2860
rect 11645 -2870 11660 -2860
rect 11700 -2870 11715 -2860
rect 11755 -2870 11770 -2860
rect 11810 -2870 11825 -2860
rect 11865 -2870 11880 -2860
rect 11920 -2870 11935 -2860
rect 11975 -2870 11990 -2860
rect 12030 -2870 12045 -2860
rect 12085 -2870 12100 -2860
rect 12140 -2870 12155 -2860
rect 12195 -2870 12210 -2860
rect 12250 -2870 12265 -2860
rect 12305 -2870 12320 -2860
rect 12360 -2870 12375 -2860
rect 12415 -2870 12430 -2860
rect 12470 -2870 12485 -2855
rect 12935 -2900 12950 -2885
rect 12990 -2900 13005 -2885
rect 13045 -2900 13060 -2885
rect 13100 -2900 13115 -2885
rect 13155 -2900 13170 -2885
rect 13210 -2900 13225 -2885
rect 13265 -2900 13280 -2885
rect 13320 -2900 13335 -2885
rect 13375 -2900 13390 -2885
rect 13430 -2900 13445 -2885
rect 13485 -2900 13500 -2885
rect 13540 -2900 13555 -2885
rect 13595 -2900 13610 -2885
rect 13650 -2900 13665 -2885
rect 13705 -2900 13720 -2885
rect 13760 -2900 13775 -2885
rect 13815 -2900 13830 -2885
rect 13870 -2900 13885 -2885
rect 13925 -2900 13940 -2885
rect 13980 -2900 13995 -2885
rect 14035 -2900 14050 -2885
rect 14090 -2900 14105 -2885
rect 13098 -2970 13132 -2960
rect 13098 -2990 13106 -2970
rect 13124 -2990 13132 -2970
rect 12935 -3015 12995 -3000
rect 13035 -3005 13995 -2990
rect 13035 -3015 13095 -3005
rect 13135 -3015 13195 -3005
rect 13235 -3015 13295 -3005
rect 13335 -3015 13395 -3005
rect 13435 -3015 13495 -3005
rect 13535 -3015 13595 -3005
rect 13635 -3015 13695 -3005
rect 13735 -3015 13795 -3005
rect 13835 -3015 13895 -3005
rect 13935 -3015 13995 -3005
rect 14035 -3015 14095 -3000
rect 11315 -3030 11330 -3020
rect 11235 -3045 11330 -3030
rect 11370 -3035 11385 -3020
rect 11425 -3035 11440 -3020
rect 11480 -3035 11495 -3020
rect 11535 -3035 11550 -3020
rect 11590 -3035 11605 -3020
rect 11645 -3035 11660 -3020
rect 11700 -3035 11715 -3020
rect 11755 -3035 11770 -3020
rect 11810 -3035 11825 -3020
rect 11865 -3035 11880 -3020
rect 11920 -3035 11935 -3020
rect 11975 -3035 11990 -3020
rect 12030 -3035 12045 -3020
rect 12085 -3035 12100 -3020
rect 12140 -3035 12155 -3020
rect 12195 -3035 12210 -3020
rect 12250 -3035 12265 -3020
rect 12305 -3035 12320 -3020
rect 12360 -3035 12375 -3020
rect 12415 -3035 12430 -3020
rect 12470 -3030 12485 -3020
rect 12470 -3045 12565 -3030
rect 11235 -3065 11245 -3045
rect 11265 -3065 11275 -3045
rect 11235 -3075 11275 -3065
rect 12525 -3065 12535 -3045
rect 12555 -3065 12565 -3045
rect 12525 -3075 12565 -3065
rect 11237 -3290 11269 -3280
rect 11237 -3310 11243 -3290
rect 11260 -3310 11269 -3290
rect 11457 -3290 11489 -3280
rect 11457 -3310 11463 -3290
rect 11480 -3310 11489 -3290
rect 11180 -3320 11269 -3310
rect 11400 -3320 11489 -3310
rect 11601 -3290 11635 -3280
rect 11601 -3310 11610 -3290
rect 11627 -3310 11635 -3290
rect 11867 -3290 11899 -3280
rect 11867 -3305 11876 -3290
rect 11601 -3320 11635 -3310
rect 11865 -3310 11876 -3305
rect 11893 -3310 11899 -3290
rect 12277 -3290 12309 -3280
rect 12277 -3310 12283 -3290
rect 12300 -3310 12309 -3290
rect 12497 -3290 12529 -3280
rect 12497 -3310 12503 -3290
rect 12520 -3310 12529 -3290
rect 11865 -3320 11899 -3310
rect 12220 -3320 12309 -3310
rect 12440 -3320 12529 -3310
rect 12641 -3290 12675 -3280
rect 12641 -3310 12650 -3290
rect 12667 -3310 12675 -3290
rect 12935 -3305 12995 -3295
rect 12641 -3320 12675 -3310
rect 12855 -3320 12995 -3305
rect 13035 -3310 13095 -3295
rect 13135 -3310 13195 -3295
rect 13235 -3310 13295 -3295
rect 13335 -3310 13395 -3295
rect 13435 -3310 13495 -3295
rect 13535 -3310 13595 -3295
rect 13635 -3310 13695 -3295
rect 13735 -3310 13795 -3295
rect 13835 -3310 13895 -3295
rect 13935 -3310 13995 -3295
rect 14035 -3305 14095 -3295
rect 14035 -3320 14175 -3305
rect 11070 -3335 11085 -3320
rect 11125 -3335 11140 -3320
rect 11180 -3325 11250 -3320
rect 11180 -3335 11195 -3325
rect 11235 -3335 11250 -3325
rect 11290 -3335 11305 -3320
rect 11345 -3335 11360 -3320
rect 11400 -3325 11470 -3320
rect 11400 -3335 11415 -3325
rect 11455 -3335 11470 -3325
rect 11510 -3335 11525 -3320
rect 11565 -3335 11580 -3320
rect 11620 -3335 11635 -3320
rect 11675 -3335 11690 -3320
rect 11810 -3335 11825 -3320
rect 11865 -3335 11880 -3320
rect 11920 -3335 11935 -3320
rect 11975 -3335 11990 -3320
rect 12110 -3335 12125 -3320
rect 12165 -3335 12180 -3320
rect 12220 -3325 12290 -3320
rect 12220 -3335 12235 -3325
rect 12275 -3335 12290 -3325
rect 12330 -3335 12345 -3320
rect 12385 -3335 12400 -3320
rect 12440 -3325 12510 -3320
rect 12440 -3335 12455 -3325
rect 12495 -3335 12510 -3325
rect 12550 -3335 12565 -3320
rect 12605 -3335 12620 -3320
rect 12660 -3335 12675 -3320
rect 12715 -3335 12730 -3320
rect 12855 -3340 12865 -3320
rect 12885 -3340 12895 -3320
rect 12855 -3350 12895 -3340
rect 14135 -3340 14145 -3320
rect 14165 -3340 14175 -3320
rect 14135 -3350 14175 -3340
rect 11070 -3495 11085 -3485
rect 10990 -3510 11085 -3495
rect 11125 -3500 11140 -3485
rect 11180 -3500 11195 -3485
rect 11235 -3500 11250 -3485
rect 11290 -3495 11305 -3485
rect 11345 -3495 11360 -3485
rect 11106 -3510 11140 -3500
rect 11290 -3510 11360 -3495
rect 11400 -3500 11415 -3485
rect 11455 -3500 11470 -3485
rect 11510 -3495 11525 -3485
rect 11565 -3495 11580 -3485
rect 11510 -3510 11580 -3495
rect 11620 -3500 11635 -3485
rect 11675 -3495 11690 -3485
rect 11810 -3495 11825 -3485
rect 11675 -3510 11825 -3495
rect 11865 -3500 11880 -3485
rect 11920 -3500 11935 -3485
rect 11975 -3495 11990 -3485
rect 12110 -3495 12125 -3485
rect 11920 -3510 11954 -3500
rect 11975 -3510 12125 -3495
rect 12165 -3500 12180 -3485
rect 12220 -3500 12235 -3485
rect 12275 -3500 12290 -3485
rect 12330 -3495 12345 -3485
rect 12385 -3495 12400 -3485
rect 12146 -3510 12180 -3500
rect 12330 -3510 12400 -3495
rect 12440 -3500 12455 -3485
rect 12495 -3500 12510 -3485
rect 12550 -3495 12565 -3485
rect 12605 -3495 12620 -3485
rect 12550 -3510 12620 -3495
rect 12660 -3500 12675 -3485
rect 12715 -3495 12730 -3485
rect 12715 -3510 12810 -3495
rect 10990 -3530 11000 -3510
rect 11020 -3530 11030 -3510
rect 10990 -3540 11030 -3530
rect 11106 -3530 11112 -3510
rect 11129 -3530 11138 -3510
rect 11106 -3540 11138 -3530
rect 11305 -3530 11315 -3510
rect 11335 -3530 11345 -3510
rect 11305 -3540 11345 -3530
rect 11525 -3530 11535 -3510
rect 11555 -3530 11565 -3510
rect 11525 -3540 11565 -3530
rect 11730 -3530 11740 -3510
rect 11760 -3530 11770 -3510
rect 11730 -3540 11770 -3530
rect 11922 -3530 11928 -3510
rect 11945 -3530 11954 -3510
rect 11922 -3540 11954 -3530
rect 12030 -3530 12040 -3510
rect 12060 -3530 12070 -3510
rect 12030 -3540 12070 -3530
rect 12146 -3530 12152 -3510
rect 12169 -3530 12178 -3510
rect 12146 -3540 12178 -3530
rect 12345 -3530 12355 -3510
rect 12375 -3530 12385 -3510
rect 12345 -3540 12385 -3530
rect 12565 -3530 12575 -3510
rect 12595 -3530 12605 -3510
rect 12565 -3540 12605 -3530
rect 12770 -3530 12780 -3510
rect 12800 -3530 12810 -3510
rect 12770 -3540 12810 -3530
rect 12595 -3755 12635 -3745
rect 12595 -3760 12605 -3755
rect 11815 -3770 11845 -3760
rect 11815 -3790 11820 -3770
rect 11840 -3790 11845 -3770
rect 12510 -3775 12605 -3760
rect 12625 -3775 12635 -3755
rect 11245 -3815 11260 -3800
rect 11300 -3805 12360 -3790
rect 11300 -3815 11315 -3805
rect 11355 -3815 11370 -3805
rect 11410 -3815 11425 -3805
rect 11465 -3815 11480 -3805
rect 11520 -3815 11535 -3805
rect 11575 -3815 11590 -3805
rect 11630 -3815 11645 -3805
rect 11685 -3815 11700 -3805
rect 11740 -3815 11755 -3805
rect 11795 -3815 11810 -3805
rect 11850 -3815 11865 -3805
rect 11905 -3815 11920 -3805
rect 11960 -3815 11975 -3805
rect 12015 -3815 12030 -3805
rect 12070 -3815 12085 -3805
rect 12125 -3815 12140 -3805
rect 12180 -3815 12195 -3805
rect 12235 -3815 12250 -3805
rect 12290 -3815 12305 -3805
rect 12345 -3815 12360 -3805
rect 12400 -3805 12470 -3790
rect 12400 -3815 12415 -3805
rect 12455 -3815 12470 -3805
rect 12510 -3815 12525 -3775
rect 12595 -3785 12635 -3775
rect 12565 -3815 12580 -3800
rect 11245 -4080 11260 -4065
rect 11300 -4080 11315 -4065
rect 11355 -4080 11370 -4065
rect 11410 -4080 11425 -4065
rect 11465 -4080 11480 -4065
rect 11520 -4080 11535 -4065
rect 11575 -4080 11590 -4065
rect 11630 -4080 11645 -4065
rect 11685 -4080 11700 -4065
rect 11740 -4080 11755 -4065
rect 11795 -4080 11810 -4065
rect 11850 -4080 11865 -4065
rect 11905 -4080 11920 -4065
rect 11960 -4080 11975 -4065
rect 12015 -4080 12030 -4065
rect 12070 -4080 12085 -4065
rect 12125 -4080 12140 -4065
rect 12180 -4080 12195 -4065
rect 12235 -4080 12250 -4065
rect 12290 -4080 12305 -4065
rect 12345 -4080 12360 -4065
rect 12400 -4080 12415 -4065
rect 12455 -4080 12470 -4065
rect 12510 -4080 12525 -4065
rect 12565 -4080 12580 -4065
rect 11165 -4090 11260 -4080
rect 11165 -4110 11175 -4090
rect 11195 -4095 11260 -4090
rect 12565 -4090 12660 -4080
rect 12565 -4095 12630 -4090
rect 11195 -4110 11205 -4095
rect 11165 -4120 11205 -4110
rect 12620 -4110 12630 -4095
rect 12650 -4110 12660 -4090
rect 12620 -4120 12660 -4110
<< polycont >>
rect 11640 9030 11660 9050
rect 11760 9030 11780 9050
rect 11880 9030 11900 9050
rect 11210 8970 11230 8990
rect 11470 8970 11490 8990
rect 11580 8985 11600 9005
rect 11940 8985 11960 9005
rect 11340 8835 11360 8855
rect 11760 8830 11780 8850
rect 12211 8830 12229 8850
rect 10915 8585 10935 8605
rect 11190 8600 11210 8620
rect 12590 8600 12610 8620
rect 10460 8320 10480 8340
rect 10720 8320 10740 8340
rect 18415 8585 18435 8605
rect 18690 8600 18710 8620
rect 20090 8600 20110 8620
rect 10590 8185 10610 8205
rect 10790 8185 10810 8205
rect 10910 8185 10930 8205
rect 10990 8185 11010 8205
rect 11110 8185 11130 8205
rect 17960 8320 17980 8340
rect 18220 8320 18240 8340
rect 11831 8130 11849 8150
rect 11190 7920 11210 7940
rect 18090 8185 18110 8205
rect 18290 8185 18310 8205
rect 18410 8185 18430 8205
rect 18490 8185 18510 8205
rect 18610 8185 18630 8205
rect 19331 8130 19349 8150
rect 12590 7920 12610 7940
rect 12865 7895 12885 7915
rect 13071 7895 13089 7915
rect 14155 7895 14175 7915
rect 18690 7920 18710 7940
rect 20090 7920 20110 7940
rect 20360 7895 20380 7915
rect 9650 7475 9670 7495
rect 10940 7475 10960 7495
rect 12865 7475 12885 7495
rect 11831 7450 11849 7470
rect 14155 7475 14175 7495
rect 20566 7895 20584 7915
rect 21650 7895 21670 7915
rect 17150 7475 17170 7495
rect 18440 7475 18460 7495
rect 20360 7475 20380 7495
rect 19331 7450 19349 7470
rect 10821 7415 10839 7435
rect 12986 7415 13004 7435
rect 21650 7475 21670 7495
rect 18321 7415 18339 7435
rect 20481 7415 20499 7435
rect 10821 7255 10839 7275
rect 12986 7255 13004 7275
rect 18321 7255 18339 7275
rect 20481 7255 20499 7275
rect 9650 7195 9670 7215
rect 10940 7195 10960 7215
rect 12865 7195 12885 7215
rect 14155 7195 14175 7215
rect 17150 7195 17170 7215
rect 18440 7195 18460 7215
rect 20360 7195 20380 7215
rect 21650 7195 21670 7215
rect 11245 6935 11265 6955
rect 12535 6935 12555 6955
rect 18745 6935 18765 6955
rect 20035 6935 20055 6955
rect 20460 6880 20480 6900
rect 20870 6880 20890 6900
rect 11243 6690 11260 6710
rect 11463 6690 11480 6710
rect 11610 6690 11627 6710
rect 11876 6690 11893 6710
rect 12283 6690 12300 6710
rect 12503 6690 12520 6710
rect 12650 6690 12667 6710
rect 18743 6690 18760 6710
rect 18963 6690 18980 6710
rect 19110 6690 19127 6710
rect 19376 6690 19393 6710
rect 19783 6690 19800 6710
rect 20003 6690 20020 6710
rect 20150 6690 20167 6710
rect 20571 6655 20591 6675
rect 20476 6545 20496 6565
rect 20854 6545 20874 6565
rect 11000 6470 11020 6490
rect 11112 6470 11129 6490
rect 11315 6470 11335 6490
rect 11535 6470 11555 6490
rect 11740 6470 11760 6490
rect 11928 6470 11945 6490
rect 12040 6470 12060 6490
rect 12152 6470 12169 6490
rect 12355 6470 12375 6490
rect 12575 6470 12595 6490
rect 12780 6470 12800 6490
rect 18500 6470 18520 6490
rect 18612 6470 18629 6490
rect 18815 6470 18835 6490
rect 19035 6470 19055 6490
rect 19240 6470 19260 6490
rect 19428 6470 19445 6490
rect 19540 6470 19560 6490
rect 19652 6470 19669 6490
rect 19855 6470 19875 6490
rect 20075 6470 20095 6490
rect 20280 6470 20300 6490
rect 10676 6310 10694 6330
rect 13106 6310 13124 6330
rect 20365 6325 20385 6345
rect 20533 6325 20553 6345
rect 20665 6325 20685 6345
rect 20797 6325 20817 6345
rect 20965 6325 20985 6345
rect 11820 6210 11840 6230
rect 12605 6225 12625 6245
rect 9635 5960 9655 5980
rect 10915 5960 10935 5980
rect 19320 6250 19340 6270
rect 20105 6265 20125 6285
rect 12865 5960 12885 5980
rect 14145 5960 14165 5980
rect 20515 5985 20535 6005
rect 20695 5985 20715 6005
rect 20815 5985 20835 6005
rect 18675 5930 18695 5950
rect 20130 5930 20150 5950
rect 11175 5890 11195 5910
rect 12630 5890 12650 5910
rect 11640 4490 11660 4510
rect 11760 4490 11780 4510
rect 11880 4490 11900 4510
rect 11210 4430 11230 4450
rect 11470 4430 11490 4450
rect 11580 4445 11600 4465
rect 11940 4445 11960 4465
rect 11340 4295 11360 4315
rect 11760 4290 11780 4310
rect 12211 4290 12229 4310
rect 11220 4180 11240 4200
rect 12510 4180 12530 4200
rect 11370 4060 11390 4080
rect 11165 3875 11185 3895
rect 11277 3875 11294 3895
rect 11480 3875 11500 3895
rect 11700 3875 11720 3895
rect 11905 3875 11925 3895
rect 12017 3875 12034 3895
rect 12220 3875 12240 3895
rect 12440 3875 12460 3895
rect 12645 3875 12665 3895
rect 11408 3755 11425 3775
rect 11628 3755 11645 3775
rect 11775 3755 11792 3775
rect 12148 3755 12165 3775
rect 12368 3755 12385 3775
rect 12515 3755 12532 3775
rect 11190 3600 11210 3620
rect 12590 3600 12610 3620
rect 3145 2955 3165 2975
rect 4845 2955 4865 2975
rect 25915 3585 25935 3605
rect 26190 3600 26210 3620
rect 27590 3600 27610 3620
rect 11831 3130 11849 3150
rect 25460 3320 25480 3340
rect 25720 3320 25740 3340
rect 25590 3185 25610 3205
rect 25790 3185 25810 3205
rect 25910 3185 25930 3205
rect 25990 3185 26010 3205
rect 26110 3185 26130 3205
rect 10125 2940 10145 2960
rect 10661 2940 10679 2960
rect 10865 2940 10885 2960
rect 11190 2920 11210 2940
rect 12590 2920 12610 2940
rect 12915 2940 12935 2960
rect 13121 2940 13139 2960
rect 13655 2940 13675 2960
rect 26831 3130 26849 3150
rect 26190 2920 26210 2940
rect 27590 2920 27610 2940
rect 27860 2895 27880 2915
rect 3005 2785 3025 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 4805 2725 4825 2745
rect 3365 2350 3385 2370
rect 3895 2355 3915 2375
rect 11831 2450 11849 2470
rect 10125 2410 10145 2430
rect 10865 2410 10885 2430
rect 12915 2410 12935 2430
rect 10775 2365 10795 2385
rect 13655 2410 13675 2430
rect 10125 2290 10145 2310
rect 13035 2350 13055 2370
rect 10865 2290 10885 2310
rect 12915 2290 12935 2310
rect 13655 2290 13675 2310
rect 11836 2155 11854 2175
rect 28066 2895 28084 2915
rect 29150 2895 29170 2915
rect 24650 2475 24670 2495
rect 25940 2475 25960 2495
rect 27860 2475 27880 2495
rect 26831 2450 26849 2470
rect 29150 2475 29170 2495
rect 25821 2415 25839 2435
rect 27981 2415 27999 2435
rect 25821 2255 25839 2275
rect 27981 2255 27999 2275
rect 24650 2195 24670 2215
rect 25940 2195 25960 2215
rect 27860 2195 27880 2215
rect 29150 2195 29170 2215
rect 11245 1935 11265 1955
rect 12535 1935 12555 1955
rect 26245 1935 26265 1955
rect 27535 1935 27555 1955
rect 2630 1855 2650 1875
rect 2775 1855 2795 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3865 1855 3885 1875
rect 3995 1850 4015 1870
rect 4125 1855 4145 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 5215 1855 5235 1875
rect 27960 1880 27980 1900
rect 28370 1880 28390 1900
rect 3235 1735 3255 1755
rect 4755 1735 4775 1755
rect 10566 1680 10584 1700
rect 11243 1690 11260 1710
rect 11463 1690 11480 1710
rect 11610 1690 11627 1710
rect 11876 1690 11893 1710
rect 12283 1690 12300 1710
rect 12503 1690 12520 1710
rect 12650 1690 12667 1710
rect 13216 1680 13234 1700
rect 26243 1690 26260 1710
rect 26463 1690 26480 1710
rect 26610 1690 26627 1710
rect 26876 1690 26893 1710
rect 27283 1690 27300 1710
rect 27503 1690 27520 1710
rect 27650 1690 27667 1710
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 3005 905 3025 925
rect 4985 905 5005 925
rect 11000 1470 11020 1490
rect 11112 1470 11129 1490
rect 11315 1470 11335 1490
rect 11535 1470 11555 1490
rect 11740 1470 11760 1490
rect 11928 1470 11945 1490
rect 12040 1470 12060 1490
rect 12152 1470 12169 1490
rect 12355 1470 12375 1490
rect 12575 1470 12595 1490
rect 12780 1470 12800 1490
rect 11820 1210 11840 1230
rect 12605 1225 12625 1245
rect 10125 910 10145 930
rect 10805 910 10825 930
rect 11175 890 11195 910
rect 12630 890 12650 910
rect 12975 910 12995 930
rect 13655 910 13675 930
rect 28071 1655 28091 1675
rect 27976 1545 27996 1565
rect 28354 1545 28374 1565
rect 26000 1470 26020 1490
rect 26112 1470 26129 1490
rect 26315 1470 26335 1490
rect 26535 1470 26555 1490
rect 26740 1470 26760 1490
rect 26928 1470 26945 1490
rect 27040 1470 27060 1490
rect 27152 1470 27169 1490
rect 27355 1470 27375 1490
rect 27575 1470 27595 1490
rect 27780 1470 27800 1490
rect 27865 1325 27885 1345
rect 28033 1325 28053 1345
rect 28165 1325 28185 1345
rect 28297 1325 28317 1345
rect 28465 1325 28485 1345
rect 26820 1250 26840 1270
rect 27605 1265 27625 1285
rect 28015 985 28035 1005
rect 28195 985 28215 1005
rect 28315 985 28335 1005
rect 26175 930 26195 950
rect 27630 930 27650 950
rect 11315 770 11335 790
rect 11385 770 11405 790
rect 11455 770 11475 790
rect 11945 775 11965 795
rect 12165 775 12185 795
rect 12385 775 12405 795
rect 3140 735 3160 755
rect 11850 655 11870 675
rect 12590 655 12610 675
rect 10915 -1415 10935 -1395
rect 11190 -1400 11210 -1380
rect 12590 -1400 12610 -1380
rect 10460 -1680 10480 -1660
rect 10720 -1680 10740 -1660
rect 10590 -1815 10610 -1795
rect 10790 -1815 10810 -1795
rect 10910 -1815 10930 -1795
rect 10990 -1815 11010 -1795
rect 11110 -1815 11130 -1795
rect 11831 -1870 11849 -1850
rect 11190 -2080 11210 -2060
rect 12590 -2080 12610 -2060
rect 12865 -2360 12885 -2340
rect 13071 -2360 13089 -2340
rect 14155 -2360 14175 -2340
rect 11831 -2550 11849 -2530
rect 12865 -2590 12885 -2570
rect 14155 -2590 14175 -2570
rect 12985 -2650 13005 -2630
rect 12865 -2710 12885 -2690
rect 14155 -2710 14175 -2690
rect 13106 -2990 13124 -2970
rect 11245 -3065 11265 -3045
rect 12535 -3065 12555 -3045
rect 11243 -3310 11260 -3290
rect 11463 -3310 11480 -3290
rect 11610 -3310 11627 -3290
rect 11876 -3310 11893 -3290
rect 12283 -3310 12300 -3290
rect 12503 -3310 12520 -3290
rect 12650 -3310 12667 -3290
rect 12865 -3340 12885 -3320
rect 14145 -3340 14165 -3320
rect 11000 -3530 11020 -3510
rect 11112 -3530 11129 -3510
rect 11315 -3530 11335 -3510
rect 11535 -3530 11555 -3510
rect 11740 -3530 11760 -3510
rect 11928 -3530 11945 -3510
rect 12040 -3530 12060 -3510
rect 12152 -3530 12169 -3510
rect 12355 -3530 12375 -3510
rect 12575 -3530 12595 -3510
rect 12780 -3530 12800 -3510
rect 11820 -3790 11840 -3770
rect 12605 -3775 12625 -3755
rect 11175 -4110 11195 -4090
rect 12630 -4110 12650 -4090
<< xpolycontact >>
rect 13100 7695 13320 7836
rect 13460 7695 13680 7836
rect 20595 7695 20815 7836
rect 20955 7695 21175 7836
rect 9845 7345 10065 7380
rect 10415 7345 10635 7380
rect 13190 7345 13410 7380
rect 13760 7345 13980 7380
rect 17345 7345 17565 7380
rect 17915 7345 18135 7380
rect 20685 7345 20905 7380
rect 21255 7345 21475 7380
rect 9845 7285 10065 7320
rect 10415 7285 10635 7320
rect 13190 7285 13410 7320
rect 13760 7285 13980 7320
rect 17345 7285 17565 7320
rect 17915 7285 18135 7320
rect 20685 7285 20905 7320
rect 21255 7285 21475 7320
rect 9805 6410 10025 6445
rect 10550 6410 10770 6445
rect 13030 6410 13250 6445
rect 13775 6410 13995 6445
rect 9899 3300 10040 3520
rect 91 3170 311 3205
rect 925 3170 1145 3205
rect 1306 3165 1526 3200
rect 2110 3165 2330 3200
rect 91 3110 311 3145
rect 925 3110 1145 3145
rect 1306 3105 1526 3140
rect 2110 3105 2330 3140
rect 91 3030 311 3065
rect 895 3030 1115 3065
rect 1306 3045 1526 3080
rect 2110 3045 2330 3080
rect 91 2970 311 3005
rect 895 2970 1115 3005
rect 1306 2985 1526 3020
rect 2110 2985 2330 3020
rect 1306 2925 1526 2960
rect 2110 2925 2330 2960
rect 9899 2940 10040 3160
rect 13760 3300 13901 3520
rect 1306 2865 1526 2900
rect 2110 2865 2330 2900
rect 96 2820 315 2855
rect 504 2820 724 2855
rect 1306 2805 1526 2840
rect 1740 2805 1960 2840
rect 13760 2940 13901 3160
rect 96 2760 315 2795
rect 504 2760 724 2795
rect 9790 2405 9825 2625
rect 9790 2010 9825 2230
rect 9850 2405 9885 2625
rect 9850 2010 9885 2230
rect 9910 2405 9945 2625
rect 9910 2010 9945 2230
rect 9970 2405 10005 2625
rect 13795 2405 13830 2625
rect 9970 2010 10005 2230
rect 13795 2010 13830 2230
rect 13855 2405 13890 2625
rect 13855 2010 13890 2230
rect 13915 2405 13950 2625
rect 13915 2010 13950 2230
rect 13975 2405 14010 2625
rect 28095 2695 28315 2836
rect 28455 2695 28675 2836
rect 24845 2345 25065 2380
rect 25415 2345 25635 2380
rect 28185 2345 28405 2380
rect 28755 2345 28975 2380
rect 24845 2285 25065 2320
rect 25415 2285 25635 2320
rect 28185 2285 28405 2320
rect 28755 2285 28975 2320
rect 13975 2010 14010 2230
rect 9970 1385 10005 1605
rect 9970 910 10005 1130
rect 10030 1385 10065 1605
rect 10030 910 10065 1130
rect 13735 1385 13770 1605
rect 13735 910 13770 1130
rect 13795 1385 13830 1605
rect 13795 910 13830 1130
<< ppolyres >>
rect 13320 7695 13460 7836
rect 20815 7695 20955 7836
rect 9899 3160 10040 3300
rect 13760 3160 13901 3300
rect 315 2820 504 2855
rect 315 2760 504 2795
rect 28315 2695 28455 2836
<< xpolyres >>
rect 10065 7345 10415 7380
rect 13410 7345 13760 7380
rect 17565 7345 17915 7380
rect 20905 7345 21255 7380
rect 10065 7285 10415 7320
rect 13410 7285 13760 7320
rect 17565 7285 17915 7320
rect 20905 7285 21255 7320
rect 10025 6410 10550 6445
rect 13250 6410 13775 6445
rect 311 3170 925 3205
rect 1526 3165 2110 3200
rect 311 3110 925 3145
rect 1526 3105 2110 3140
rect 311 3030 895 3065
rect 1526 3045 2110 3080
rect 311 2970 895 3005
rect 1526 2985 2110 3020
rect 1526 2925 2110 2960
rect 1526 2865 2110 2900
rect 1526 2805 1740 2840
rect 9790 2230 9825 2405
rect 9850 2230 9885 2405
rect 9910 2230 9945 2405
rect 9970 2230 10005 2405
rect 13795 2230 13830 2405
rect 13855 2230 13890 2405
rect 13915 2230 13950 2405
rect 13975 2230 14010 2405
rect 25065 2345 25415 2380
rect 28405 2345 28755 2380
rect 25065 2285 25415 2320
rect 28405 2285 28755 2320
rect 9970 1130 10005 1385
rect 10030 1130 10065 1385
rect 13735 1130 13770 1385
rect 13795 1130 13830 1385
<< locali >>
rect 11632 9050 11668 9060
rect 11632 9030 11640 9050
rect 11660 9030 11668 9050
rect 11632 9020 11668 9030
rect 11752 9050 11788 9060
rect 11752 9030 11760 9050
rect 11780 9030 11788 9050
rect 11752 9020 11788 9030
rect 11872 9050 11908 9060
rect 11872 9030 11880 9050
rect 11900 9030 11908 9050
rect 11872 9020 11908 9030
rect 11570 9005 11610 9015
rect 11200 8990 11240 9000
rect 11200 8970 11210 8990
rect 11230 8970 11240 8990
rect 11200 8960 11240 8970
rect 11460 8990 11500 9000
rect 11460 8970 11470 8990
rect 11490 8970 11500 8990
rect 11570 8985 11580 9005
rect 11600 8985 11610 9005
rect 11570 8975 11610 8985
rect 11460 8960 11500 8970
rect 11210 8938 11230 8960
rect 11470 8938 11490 8960
rect 11580 8955 11600 8975
rect 11640 8955 11660 9020
rect 11690 9005 11730 9015
rect 11690 8985 11700 9005
rect 11720 8985 11730 9005
rect 11690 8975 11730 8985
rect 11700 8955 11720 8975
rect 11760 8955 11780 9020
rect 11810 9005 11850 9015
rect 11810 8985 11820 9005
rect 11840 8985 11850 9005
rect 11810 8975 11850 8985
rect 11820 8955 11840 8975
rect 11880 8955 11900 9020
rect 11930 9005 11970 9015
rect 11930 8985 11940 9005
rect 11960 8985 11970 9005
rect 11930 8975 11970 8985
rect 12080 8980 12120 8990
rect 11940 8955 11960 8975
rect 12080 8960 12090 8980
rect 12110 8960 12120 8980
rect 11205 8915 11275 8938
rect 11205 8895 11210 8915
rect 11230 8895 11250 8915
rect 11270 8895 11275 8915
rect 11205 8885 11275 8895
rect 11305 8920 11335 8938
rect 11305 8900 11310 8920
rect 11330 8900 11335 8920
rect 11305 8885 11335 8900
rect 11365 8920 11395 8938
rect 11365 8900 11370 8920
rect 11390 8900 11395 8920
rect 11365 8885 11395 8900
rect 11425 8915 11495 8938
rect 11425 8895 11430 8915
rect 11450 8895 11470 8915
rect 11490 8895 11495 8915
rect 11425 8885 11495 8895
rect 11535 8930 11605 8955
rect 11535 8910 11540 8930
rect 11560 8910 11580 8930
rect 11600 8910 11605 8930
rect 11535 8885 11605 8910
rect 11635 8930 11665 8955
rect 11635 8910 11640 8930
rect 11660 8910 11665 8930
rect 11635 8885 11665 8910
rect 11695 8930 11725 8955
rect 11695 8910 11700 8930
rect 11720 8910 11725 8930
rect 11695 8885 11725 8910
rect 11755 8930 11785 8955
rect 11755 8910 11760 8930
rect 11780 8910 11785 8930
rect 11755 8885 11785 8910
rect 11815 8930 11845 8955
rect 11815 8910 11820 8930
rect 11840 8910 11845 8930
rect 11815 8885 11845 8910
rect 11875 8930 11905 8955
rect 11875 8910 11880 8930
rect 11900 8910 11905 8930
rect 11875 8885 11905 8910
rect 11935 8930 12005 8955
rect 12080 8950 12120 8960
rect 12200 8980 12240 8990
rect 12200 8960 12210 8980
rect 12230 8960 12240 8980
rect 12200 8950 12240 8960
rect 12320 8980 12360 8990
rect 12320 8960 12330 8980
rect 12350 8960 12360 8980
rect 12320 8950 12360 8960
rect 12440 8980 12480 8990
rect 12440 8960 12450 8980
rect 12470 8960 12480 8980
rect 12440 8950 12480 8960
rect 12560 8980 12600 8990
rect 12560 8960 12570 8980
rect 12590 8960 12600 8980
rect 12560 8950 12600 8960
rect 12090 8930 12110 8950
rect 12210 8930 12230 8950
rect 12330 8930 12350 8950
rect 12450 8930 12470 8950
rect 12570 8930 12590 8950
rect 11935 8910 11940 8930
rect 11960 8910 11980 8930
rect 12000 8910 12005 8930
rect 11935 8885 12005 8910
rect 12045 8915 12115 8930
rect 12045 8895 12050 8915
rect 12070 8895 12090 8915
rect 12110 8895 12115 8915
rect 11370 8865 11390 8885
rect 12045 8880 12115 8895
rect 12145 8915 12175 8930
rect 12145 8895 12150 8915
rect 12170 8895 12175 8915
rect 12145 8880 12175 8895
rect 12205 8915 12235 8930
rect 12205 8895 12210 8915
rect 12230 8895 12235 8915
rect 12205 8880 12235 8895
rect 12265 8915 12295 8930
rect 12265 8895 12270 8915
rect 12290 8895 12295 8915
rect 12265 8880 12295 8895
rect 12325 8915 12355 8930
rect 12325 8895 12330 8915
rect 12350 8895 12355 8915
rect 12325 8880 12355 8895
rect 12385 8915 12415 8930
rect 12385 8895 12390 8915
rect 12410 8895 12415 8915
rect 12385 8880 12415 8895
rect 12445 8915 12475 8930
rect 12445 8895 12450 8915
rect 12470 8895 12475 8915
rect 12445 8880 12475 8895
rect 12505 8915 12535 8930
rect 12505 8895 12510 8915
rect 12530 8895 12535 8915
rect 12505 8880 12535 8895
rect 12565 8915 12635 8930
rect 12565 8895 12570 8915
rect 12590 8895 12610 8915
rect 12630 8895 12635 8915
rect 12565 8880 12635 8895
rect 11330 8860 11390 8865
rect 12150 8860 12170 8880
rect 12270 8860 12290 8880
rect 12390 8860 12410 8880
rect 12510 8860 12530 8880
rect 11330 8835 11340 8860
rect 11360 8845 11390 8860
rect 11750 8850 11790 8860
rect 11360 8835 11370 8845
rect 11330 8825 11370 8835
rect 11750 8830 11760 8850
rect 11780 8830 11790 8850
rect 11750 8820 11790 8830
rect 12140 8850 12180 8860
rect 12140 8830 12150 8850
rect 12170 8830 12180 8850
rect 12140 8820 12180 8830
rect 12203 8850 12237 8860
rect 12203 8830 12211 8850
rect 12229 8830 12237 8850
rect 12203 8820 12237 8830
rect 12260 8850 12300 8860
rect 12260 8830 12270 8850
rect 12290 8830 12300 8850
rect 12260 8820 12300 8830
rect 12380 8850 12420 8860
rect 12380 8830 12390 8850
rect 12410 8830 12420 8850
rect 12380 8820 12420 8830
rect 12500 8850 12540 8860
rect 12500 8830 12510 8850
rect 12530 8830 12540 8850
rect 12500 8820 12540 8830
rect 11180 8620 11220 8630
rect 10905 8605 11030 8615
rect 10905 8585 10915 8605
rect 10935 8595 11030 8605
rect 10935 8585 10945 8595
rect 10905 8575 10945 8585
rect 11010 8575 11030 8595
rect 11180 8600 11190 8620
rect 11210 8600 11220 8620
rect 11180 8590 11220 8600
rect 11340 8620 11380 8630
rect 11340 8600 11350 8620
rect 11370 8600 11380 8620
rect 11340 8590 11380 8600
rect 11460 8620 11500 8630
rect 11460 8600 11470 8620
rect 11490 8600 11500 8620
rect 11460 8590 11500 8600
rect 11580 8620 11620 8630
rect 11580 8600 11590 8620
rect 11610 8600 11620 8620
rect 11580 8590 11620 8600
rect 11700 8620 11740 8630
rect 11700 8600 11710 8620
rect 11730 8600 11740 8620
rect 11700 8590 11740 8600
rect 11820 8620 11860 8630
rect 11820 8600 11830 8620
rect 11850 8600 11860 8620
rect 11820 8590 11860 8600
rect 11940 8620 11980 8630
rect 11940 8600 11950 8620
rect 11970 8600 11980 8620
rect 11940 8590 11980 8600
rect 12060 8620 12100 8630
rect 12060 8600 12070 8620
rect 12090 8600 12100 8620
rect 12060 8590 12100 8600
rect 12180 8620 12220 8630
rect 12180 8600 12190 8620
rect 12210 8600 12220 8620
rect 12180 8590 12220 8600
rect 12300 8620 12340 8630
rect 12300 8600 12310 8620
rect 12330 8600 12340 8620
rect 12300 8590 12340 8600
rect 12420 8620 12460 8630
rect 12420 8600 12430 8620
rect 12450 8600 12460 8620
rect 12420 8590 12460 8600
rect 12580 8620 12620 8630
rect 12580 8600 12590 8620
rect 12610 8600 12620 8620
rect 18680 8620 18720 8630
rect 12580 8590 12620 8600
rect 18405 8605 18530 8615
rect 11005 8565 11035 8575
rect 11005 8545 11010 8565
rect 11030 8545 11035 8565
rect 10785 8515 10855 8545
rect 10785 8495 10790 8515
rect 10810 8495 10830 8515
rect 10850 8495 10855 8515
rect 10785 8465 10855 8495
rect 10785 8445 10790 8465
rect 10810 8445 10830 8465
rect 10850 8445 10855 8465
rect 10785 8415 10855 8445
rect 10785 8395 10790 8415
rect 10810 8395 10830 8415
rect 10850 8395 10855 8415
rect 10785 8365 10855 8395
rect 10450 8340 10490 8350
rect 10450 8320 10460 8340
rect 10480 8320 10490 8340
rect 10450 8310 10490 8320
rect 10710 8340 10750 8350
rect 10710 8320 10720 8340
rect 10740 8320 10750 8340
rect 10710 8310 10750 8320
rect 10785 8345 10790 8365
rect 10810 8345 10830 8365
rect 10850 8345 10855 8365
rect 10785 8315 10855 8345
rect 10460 8288 10480 8310
rect 10720 8288 10740 8310
rect 10785 8295 10790 8315
rect 10810 8295 10830 8315
rect 10850 8295 10855 8315
rect 10455 8265 10525 8288
rect 10455 8245 10460 8265
rect 10480 8245 10500 8265
rect 10520 8245 10525 8265
rect 10455 8235 10525 8245
rect 10555 8270 10585 8288
rect 10555 8250 10560 8270
rect 10580 8250 10585 8270
rect 10555 8235 10585 8250
rect 10615 8270 10645 8288
rect 10615 8250 10620 8270
rect 10640 8250 10645 8270
rect 10615 8235 10645 8250
rect 10675 8265 10745 8288
rect 10675 8245 10680 8265
rect 10700 8245 10720 8265
rect 10740 8245 10745 8265
rect 10675 8235 10745 8245
rect 10785 8265 10855 8295
rect 10785 8245 10790 8265
rect 10810 8245 10830 8265
rect 10850 8245 10855 8265
rect 10785 8235 10855 8245
rect 10885 8515 10915 8545
rect 10885 8495 10890 8515
rect 10910 8495 10915 8515
rect 10885 8465 10915 8495
rect 10885 8445 10890 8465
rect 10910 8445 10915 8465
rect 10885 8415 10915 8445
rect 10885 8395 10890 8415
rect 10910 8395 10915 8415
rect 10885 8365 10915 8395
rect 10885 8345 10890 8365
rect 10910 8345 10915 8365
rect 10885 8315 10915 8345
rect 10885 8295 10890 8315
rect 10910 8295 10915 8315
rect 10885 8265 10915 8295
rect 10885 8245 10890 8265
rect 10910 8245 10915 8265
rect 10885 8235 10915 8245
rect 10945 8515 10975 8545
rect 10945 8495 10950 8515
rect 10970 8495 10975 8515
rect 10945 8465 10975 8495
rect 10945 8445 10950 8465
rect 10970 8445 10975 8465
rect 10945 8415 10975 8445
rect 10945 8395 10950 8415
rect 10970 8395 10975 8415
rect 10945 8365 10975 8395
rect 10945 8345 10950 8365
rect 10970 8345 10975 8365
rect 10945 8315 10975 8345
rect 10945 8295 10950 8315
rect 10970 8295 10975 8315
rect 10945 8265 10975 8295
rect 10945 8245 10950 8265
rect 10970 8245 10975 8265
rect 10945 8235 10975 8245
rect 11005 8515 11035 8545
rect 11005 8495 11010 8515
rect 11030 8495 11035 8515
rect 11005 8465 11035 8495
rect 11005 8445 11010 8465
rect 11030 8445 11035 8465
rect 11005 8415 11035 8445
rect 11005 8395 11010 8415
rect 11030 8395 11035 8415
rect 11005 8365 11035 8395
rect 11005 8345 11010 8365
rect 11030 8345 11035 8365
rect 11005 8315 11035 8345
rect 11005 8295 11010 8315
rect 11030 8295 11035 8315
rect 11005 8265 11035 8295
rect 11005 8245 11010 8265
rect 11030 8245 11035 8265
rect 11005 8235 11035 8245
rect 11065 8565 11135 8575
rect 11190 8570 11210 8590
rect 11350 8570 11370 8590
rect 11470 8570 11490 8590
rect 11590 8570 11610 8590
rect 11710 8570 11730 8590
rect 11830 8570 11850 8590
rect 11950 8570 11970 8590
rect 12070 8570 12090 8590
rect 12190 8570 12210 8590
rect 12310 8570 12330 8590
rect 12430 8570 12450 8590
rect 12590 8570 12610 8590
rect 18405 8585 18415 8605
rect 18435 8595 18530 8605
rect 18435 8585 18445 8595
rect 18405 8575 18445 8585
rect 18510 8575 18530 8595
rect 18680 8600 18690 8620
rect 18710 8600 18720 8620
rect 18680 8590 18720 8600
rect 18840 8620 18880 8630
rect 18840 8600 18850 8620
rect 18870 8600 18880 8620
rect 18840 8590 18880 8600
rect 18960 8620 19000 8630
rect 18960 8600 18970 8620
rect 18990 8600 19000 8620
rect 18960 8590 19000 8600
rect 19080 8620 19120 8630
rect 19080 8600 19090 8620
rect 19110 8600 19120 8620
rect 19080 8590 19120 8600
rect 19200 8620 19240 8630
rect 19200 8600 19210 8620
rect 19230 8600 19240 8620
rect 19200 8590 19240 8600
rect 19320 8620 19360 8630
rect 19320 8600 19330 8620
rect 19350 8600 19360 8620
rect 19320 8590 19360 8600
rect 19440 8620 19480 8630
rect 19440 8600 19450 8620
rect 19470 8600 19480 8620
rect 19440 8590 19480 8600
rect 19560 8620 19600 8630
rect 19560 8600 19570 8620
rect 19590 8600 19600 8620
rect 19560 8590 19600 8600
rect 19680 8620 19720 8630
rect 19680 8600 19690 8620
rect 19710 8600 19720 8620
rect 19680 8590 19720 8600
rect 19800 8620 19840 8630
rect 19800 8600 19810 8620
rect 19830 8600 19840 8620
rect 19800 8590 19840 8600
rect 19920 8620 19960 8630
rect 19920 8600 19930 8620
rect 19950 8600 19960 8620
rect 19920 8590 19960 8600
rect 20080 8620 20120 8630
rect 20080 8600 20090 8620
rect 20110 8600 20120 8620
rect 20080 8590 20120 8600
rect 11065 8545 11070 8565
rect 11090 8545 11110 8565
rect 11130 8545 11135 8565
rect 11065 8515 11135 8545
rect 11065 8495 11070 8515
rect 11090 8495 11110 8515
rect 11130 8495 11135 8515
rect 11065 8465 11135 8495
rect 11065 8445 11070 8465
rect 11090 8445 11110 8465
rect 11130 8445 11135 8465
rect 11065 8415 11135 8445
rect 11065 8395 11070 8415
rect 11090 8395 11110 8415
rect 11130 8395 11135 8415
rect 11065 8365 11135 8395
rect 11065 8345 11070 8365
rect 11090 8345 11110 8365
rect 11130 8345 11135 8365
rect 11065 8315 11135 8345
rect 11065 8295 11070 8315
rect 11090 8295 11110 8315
rect 11130 8295 11135 8315
rect 11065 8265 11135 8295
rect 11065 8245 11070 8265
rect 11090 8245 11110 8265
rect 11130 8245 11135 8265
rect 11065 8235 11135 8245
rect 11185 8560 11255 8570
rect 11185 8540 11190 8560
rect 11210 8540 11230 8560
rect 11250 8540 11255 8560
rect 11185 8510 11255 8540
rect 11185 8490 11190 8510
rect 11210 8490 11230 8510
rect 11250 8490 11255 8510
rect 11185 8460 11255 8490
rect 11185 8440 11190 8460
rect 11210 8440 11230 8460
rect 11250 8440 11255 8460
rect 11185 8410 11255 8440
rect 11185 8390 11190 8410
rect 11210 8390 11230 8410
rect 11250 8390 11255 8410
rect 11185 8360 11255 8390
rect 11185 8340 11190 8360
rect 11210 8340 11230 8360
rect 11250 8340 11255 8360
rect 11185 8310 11255 8340
rect 11185 8290 11190 8310
rect 11210 8290 11230 8310
rect 11250 8290 11255 8310
rect 11185 8260 11255 8290
rect 11185 8240 11190 8260
rect 11210 8240 11230 8260
rect 11250 8240 11255 8260
rect 10620 8215 10640 8235
rect 10790 8215 10810 8235
rect 11110 8215 11130 8235
rect 10580 8205 10640 8215
rect 10580 8185 10590 8205
rect 10610 8195 10640 8205
rect 10780 8205 10820 8215
rect 10610 8185 10620 8195
rect 10580 8175 10620 8185
rect 10780 8185 10790 8205
rect 10810 8185 10820 8205
rect 10780 8175 10820 8185
rect 10905 8205 10940 8215
rect 10905 8185 10910 8205
rect 10930 8185 10940 8205
rect 10905 8175 10940 8185
rect 10980 8205 11015 8215
rect 10980 8185 10990 8205
rect 11010 8185 11015 8205
rect 10980 8175 11015 8185
rect 11100 8205 11140 8215
rect 11100 8185 11110 8205
rect 11130 8185 11140 8205
rect 11100 8175 11140 8185
rect 11185 8210 11255 8240
rect 11185 8190 11190 8210
rect 11210 8190 11230 8210
rect 11250 8190 11255 8210
rect 11185 8180 11255 8190
rect 11285 8560 11315 8570
rect 11285 8540 11290 8560
rect 11310 8540 11315 8560
rect 11285 8510 11315 8540
rect 11285 8490 11290 8510
rect 11310 8490 11315 8510
rect 11285 8460 11315 8490
rect 11285 8440 11290 8460
rect 11310 8440 11315 8460
rect 11285 8410 11315 8440
rect 11285 8390 11290 8410
rect 11310 8390 11315 8410
rect 11285 8360 11315 8390
rect 11285 8340 11290 8360
rect 11310 8340 11315 8360
rect 11285 8310 11315 8340
rect 11285 8290 11290 8310
rect 11310 8290 11315 8310
rect 11285 8260 11315 8290
rect 11285 8240 11290 8260
rect 11310 8240 11315 8260
rect 11285 8210 11315 8240
rect 11285 8190 11290 8210
rect 11310 8190 11315 8210
rect 11285 8180 11315 8190
rect 11345 8560 11375 8570
rect 11345 8540 11350 8560
rect 11370 8540 11375 8560
rect 11345 8510 11375 8540
rect 11345 8490 11350 8510
rect 11370 8490 11375 8510
rect 11345 8460 11375 8490
rect 11345 8440 11350 8460
rect 11370 8440 11375 8460
rect 11345 8410 11375 8440
rect 11345 8390 11350 8410
rect 11370 8390 11375 8410
rect 11345 8360 11375 8390
rect 11345 8340 11350 8360
rect 11370 8340 11375 8360
rect 11345 8310 11375 8340
rect 11345 8290 11350 8310
rect 11370 8290 11375 8310
rect 11345 8260 11375 8290
rect 11345 8240 11350 8260
rect 11370 8240 11375 8260
rect 11345 8210 11375 8240
rect 11345 8190 11350 8210
rect 11370 8190 11375 8210
rect 11345 8180 11375 8190
rect 11405 8560 11435 8570
rect 11405 8540 11410 8560
rect 11430 8540 11435 8560
rect 11405 8510 11435 8540
rect 11405 8490 11410 8510
rect 11430 8490 11435 8510
rect 11405 8460 11435 8490
rect 11405 8440 11410 8460
rect 11430 8440 11435 8460
rect 11405 8410 11435 8440
rect 11405 8390 11410 8410
rect 11430 8390 11435 8410
rect 11405 8360 11435 8390
rect 11405 8340 11410 8360
rect 11430 8340 11435 8360
rect 11405 8310 11435 8340
rect 11405 8290 11410 8310
rect 11430 8290 11435 8310
rect 11405 8260 11435 8290
rect 11405 8240 11410 8260
rect 11430 8240 11435 8260
rect 11405 8210 11435 8240
rect 11405 8190 11410 8210
rect 11430 8190 11435 8210
rect 11405 8180 11435 8190
rect 11465 8560 11495 8570
rect 11465 8540 11470 8560
rect 11490 8540 11495 8560
rect 11465 8510 11495 8540
rect 11465 8490 11470 8510
rect 11490 8490 11495 8510
rect 11465 8460 11495 8490
rect 11465 8440 11470 8460
rect 11490 8440 11495 8460
rect 11465 8410 11495 8440
rect 11465 8390 11470 8410
rect 11490 8390 11495 8410
rect 11465 8360 11495 8390
rect 11465 8340 11470 8360
rect 11490 8340 11495 8360
rect 11465 8310 11495 8340
rect 11465 8290 11470 8310
rect 11490 8290 11495 8310
rect 11465 8260 11495 8290
rect 11465 8240 11470 8260
rect 11490 8240 11495 8260
rect 11465 8210 11495 8240
rect 11465 8190 11470 8210
rect 11490 8190 11495 8210
rect 11465 8180 11495 8190
rect 11525 8560 11555 8570
rect 11525 8540 11530 8560
rect 11550 8540 11555 8560
rect 11525 8510 11555 8540
rect 11525 8490 11530 8510
rect 11550 8490 11555 8510
rect 11525 8460 11555 8490
rect 11525 8440 11530 8460
rect 11550 8440 11555 8460
rect 11525 8410 11555 8440
rect 11525 8390 11530 8410
rect 11550 8390 11555 8410
rect 11525 8360 11555 8390
rect 11525 8340 11530 8360
rect 11550 8340 11555 8360
rect 11525 8310 11555 8340
rect 11525 8290 11530 8310
rect 11550 8290 11555 8310
rect 11525 8260 11555 8290
rect 11525 8240 11530 8260
rect 11550 8240 11555 8260
rect 11525 8210 11555 8240
rect 11525 8190 11530 8210
rect 11550 8190 11555 8210
rect 11525 8180 11555 8190
rect 11585 8560 11615 8570
rect 11585 8540 11590 8560
rect 11610 8540 11615 8560
rect 11585 8510 11615 8540
rect 11585 8490 11590 8510
rect 11610 8490 11615 8510
rect 11585 8460 11615 8490
rect 11585 8440 11590 8460
rect 11610 8440 11615 8460
rect 11585 8410 11615 8440
rect 11585 8390 11590 8410
rect 11610 8390 11615 8410
rect 11585 8360 11615 8390
rect 11585 8340 11590 8360
rect 11610 8340 11615 8360
rect 11585 8310 11615 8340
rect 11585 8290 11590 8310
rect 11610 8290 11615 8310
rect 11585 8260 11615 8290
rect 11585 8240 11590 8260
rect 11610 8240 11615 8260
rect 11585 8210 11615 8240
rect 11585 8190 11590 8210
rect 11610 8190 11615 8210
rect 11585 8180 11615 8190
rect 11645 8560 11675 8570
rect 11645 8540 11650 8560
rect 11670 8540 11675 8560
rect 11645 8510 11675 8540
rect 11645 8490 11650 8510
rect 11670 8490 11675 8510
rect 11645 8460 11675 8490
rect 11645 8440 11650 8460
rect 11670 8440 11675 8460
rect 11645 8410 11675 8440
rect 11645 8390 11650 8410
rect 11670 8390 11675 8410
rect 11645 8360 11675 8390
rect 11645 8340 11650 8360
rect 11670 8340 11675 8360
rect 11645 8310 11675 8340
rect 11645 8290 11650 8310
rect 11670 8290 11675 8310
rect 11645 8260 11675 8290
rect 11645 8240 11650 8260
rect 11670 8240 11675 8260
rect 11645 8210 11675 8240
rect 11645 8190 11650 8210
rect 11670 8190 11675 8210
rect 11645 8180 11675 8190
rect 11705 8560 11735 8570
rect 11705 8540 11710 8560
rect 11730 8540 11735 8560
rect 11705 8510 11735 8540
rect 11705 8490 11710 8510
rect 11730 8490 11735 8510
rect 11705 8460 11735 8490
rect 11705 8440 11710 8460
rect 11730 8440 11735 8460
rect 11705 8410 11735 8440
rect 11705 8390 11710 8410
rect 11730 8390 11735 8410
rect 11705 8360 11735 8390
rect 11705 8340 11710 8360
rect 11730 8340 11735 8360
rect 11705 8310 11735 8340
rect 11705 8290 11710 8310
rect 11730 8290 11735 8310
rect 11705 8260 11735 8290
rect 11705 8240 11710 8260
rect 11730 8240 11735 8260
rect 11705 8210 11735 8240
rect 11705 8190 11710 8210
rect 11730 8190 11735 8210
rect 11705 8180 11735 8190
rect 11765 8560 11795 8570
rect 11765 8540 11770 8560
rect 11790 8540 11795 8560
rect 11765 8510 11795 8540
rect 11765 8490 11770 8510
rect 11790 8490 11795 8510
rect 11765 8460 11795 8490
rect 11765 8440 11770 8460
rect 11790 8440 11795 8460
rect 11765 8410 11795 8440
rect 11765 8390 11770 8410
rect 11790 8390 11795 8410
rect 11765 8360 11795 8390
rect 11765 8340 11770 8360
rect 11790 8340 11795 8360
rect 11765 8310 11795 8340
rect 11765 8290 11770 8310
rect 11790 8290 11795 8310
rect 11765 8260 11795 8290
rect 11765 8240 11770 8260
rect 11790 8240 11795 8260
rect 11765 8210 11795 8240
rect 11765 8190 11770 8210
rect 11790 8190 11795 8210
rect 11765 8180 11795 8190
rect 11825 8560 11855 8570
rect 11825 8540 11830 8560
rect 11850 8540 11855 8560
rect 11825 8510 11855 8540
rect 11825 8490 11830 8510
rect 11850 8490 11855 8510
rect 11825 8460 11855 8490
rect 11825 8440 11830 8460
rect 11850 8440 11855 8460
rect 11825 8410 11855 8440
rect 11825 8390 11830 8410
rect 11850 8390 11855 8410
rect 11825 8360 11855 8390
rect 11825 8340 11830 8360
rect 11850 8340 11855 8360
rect 11825 8310 11855 8340
rect 11825 8290 11830 8310
rect 11850 8290 11855 8310
rect 11825 8260 11855 8290
rect 11825 8240 11830 8260
rect 11850 8240 11855 8260
rect 11825 8210 11855 8240
rect 11825 8190 11830 8210
rect 11850 8190 11855 8210
rect 11825 8180 11855 8190
rect 11885 8560 11915 8570
rect 11885 8540 11890 8560
rect 11910 8540 11915 8560
rect 11885 8510 11915 8540
rect 11885 8490 11890 8510
rect 11910 8490 11915 8510
rect 11885 8460 11915 8490
rect 11885 8440 11890 8460
rect 11910 8440 11915 8460
rect 11885 8410 11915 8440
rect 11885 8390 11890 8410
rect 11910 8390 11915 8410
rect 11885 8360 11915 8390
rect 11885 8340 11890 8360
rect 11910 8340 11915 8360
rect 11885 8310 11915 8340
rect 11885 8290 11890 8310
rect 11910 8290 11915 8310
rect 11885 8260 11915 8290
rect 11885 8240 11890 8260
rect 11910 8240 11915 8260
rect 11885 8210 11915 8240
rect 11885 8190 11890 8210
rect 11910 8190 11915 8210
rect 11885 8180 11915 8190
rect 11945 8560 11975 8570
rect 11945 8540 11950 8560
rect 11970 8540 11975 8560
rect 11945 8510 11975 8540
rect 11945 8490 11950 8510
rect 11970 8490 11975 8510
rect 11945 8460 11975 8490
rect 11945 8440 11950 8460
rect 11970 8440 11975 8460
rect 11945 8410 11975 8440
rect 11945 8390 11950 8410
rect 11970 8390 11975 8410
rect 11945 8360 11975 8390
rect 11945 8340 11950 8360
rect 11970 8340 11975 8360
rect 11945 8310 11975 8340
rect 11945 8290 11950 8310
rect 11970 8290 11975 8310
rect 11945 8260 11975 8290
rect 11945 8240 11950 8260
rect 11970 8240 11975 8260
rect 11945 8210 11975 8240
rect 11945 8190 11950 8210
rect 11970 8190 11975 8210
rect 11945 8180 11975 8190
rect 12005 8560 12035 8570
rect 12005 8540 12010 8560
rect 12030 8540 12035 8560
rect 12005 8510 12035 8540
rect 12005 8490 12010 8510
rect 12030 8490 12035 8510
rect 12005 8460 12035 8490
rect 12005 8440 12010 8460
rect 12030 8440 12035 8460
rect 12005 8410 12035 8440
rect 12005 8390 12010 8410
rect 12030 8390 12035 8410
rect 12005 8360 12035 8390
rect 12005 8340 12010 8360
rect 12030 8340 12035 8360
rect 12005 8310 12035 8340
rect 12005 8290 12010 8310
rect 12030 8290 12035 8310
rect 12005 8260 12035 8290
rect 12005 8240 12010 8260
rect 12030 8240 12035 8260
rect 12005 8210 12035 8240
rect 12005 8190 12010 8210
rect 12030 8190 12035 8210
rect 12005 8180 12035 8190
rect 12065 8560 12095 8570
rect 12065 8540 12070 8560
rect 12090 8540 12095 8560
rect 12065 8510 12095 8540
rect 12065 8490 12070 8510
rect 12090 8490 12095 8510
rect 12065 8460 12095 8490
rect 12065 8440 12070 8460
rect 12090 8440 12095 8460
rect 12065 8410 12095 8440
rect 12065 8390 12070 8410
rect 12090 8390 12095 8410
rect 12065 8360 12095 8390
rect 12065 8340 12070 8360
rect 12090 8340 12095 8360
rect 12065 8310 12095 8340
rect 12065 8290 12070 8310
rect 12090 8290 12095 8310
rect 12065 8260 12095 8290
rect 12065 8240 12070 8260
rect 12090 8240 12095 8260
rect 12065 8210 12095 8240
rect 12065 8190 12070 8210
rect 12090 8190 12095 8210
rect 12065 8180 12095 8190
rect 12125 8560 12155 8570
rect 12125 8540 12130 8560
rect 12150 8540 12155 8560
rect 12125 8510 12155 8540
rect 12125 8490 12130 8510
rect 12150 8490 12155 8510
rect 12125 8460 12155 8490
rect 12125 8440 12130 8460
rect 12150 8440 12155 8460
rect 12125 8410 12155 8440
rect 12125 8390 12130 8410
rect 12150 8390 12155 8410
rect 12125 8360 12155 8390
rect 12125 8340 12130 8360
rect 12150 8340 12155 8360
rect 12125 8310 12155 8340
rect 12125 8290 12130 8310
rect 12150 8290 12155 8310
rect 12125 8260 12155 8290
rect 12125 8240 12130 8260
rect 12150 8240 12155 8260
rect 12125 8210 12155 8240
rect 12125 8190 12130 8210
rect 12150 8190 12155 8210
rect 12125 8180 12155 8190
rect 12185 8560 12215 8570
rect 12185 8540 12190 8560
rect 12210 8540 12215 8560
rect 12185 8510 12215 8540
rect 12185 8490 12190 8510
rect 12210 8490 12215 8510
rect 12185 8460 12215 8490
rect 12185 8440 12190 8460
rect 12210 8440 12215 8460
rect 12185 8410 12215 8440
rect 12185 8390 12190 8410
rect 12210 8390 12215 8410
rect 12185 8360 12215 8390
rect 12185 8340 12190 8360
rect 12210 8340 12215 8360
rect 12185 8310 12215 8340
rect 12185 8290 12190 8310
rect 12210 8290 12215 8310
rect 12185 8260 12215 8290
rect 12185 8240 12190 8260
rect 12210 8240 12215 8260
rect 12185 8210 12215 8240
rect 12185 8190 12190 8210
rect 12210 8190 12215 8210
rect 12185 8180 12215 8190
rect 12245 8560 12275 8570
rect 12245 8540 12250 8560
rect 12270 8540 12275 8560
rect 12245 8510 12275 8540
rect 12245 8490 12250 8510
rect 12270 8490 12275 8510
rect 12245 8460 12275 8490
rect 12245 8440 12250 8460
rect 12270 8440 12275 8460
rect 12245 8410 12275 8440
rect 12245 8390 12250 8410
rect 12270 8390 12275 8410
rect 12245 8360 12275 8390
rect 12245 8340 12250 8360
rect 12270 8340 12275 8360
rect 12245 8310 12275 8340
rect 12245 8290 12250 8310
rect 12270 8290 12275 8310
rect 12245 8260 12275 8290
rect 12245 8240 12250 8260
rect 12270 8240 12275 8260
rect 12245 8210 12275 8240
rect 12245 8190 12250 8210
rect 12270 8190 12275 8210
rect 12245 8180 12275 8190
rect 12305 8560 12335 8570
rect 12305 8540 12310 8560
rect 12330 8540 12335 8560
rect 12305 8510 12335 8540
rect 12305 8490 12310 8510
rect 12330 8490 12335 8510
rect 12305 8460 12335 8490
rect 12305 8440 12310 8460
rect 12330 8440 12335 8460
rect 12305 8410 12335 8440
rect 12305 8390 12310 8410
rect 12330 8390 12335 8410
rect 12305 8360 12335 8390
rect 12305 8340 12310 8360
rect 12330 8340 12335 8360
rect 12305 8310 12335 8340
rect 12305 8290 12310 8310
rect 12330 8290 12335 8310
rect 12305 8260 12335 8290
rect 12305 8240 12310 8260
rect 12330 8240 12335 8260
rect 12305 8210 12335 8240
rect 12305 8190 12310 8210
rect 12330 8190 12335 8210
rect 12305 8180 12335 8190
rect 12365 8560 12395 8570
rect 12365 8540 12370 8560
rect 12390 8540 12395 8560
rect 12365 8510 12395 8540
rect 12365 8490 12370 8510
rect 12390 8490 12395 8510
rect 12365 8460 12395 8490
rect 12365 8440 12370 8460
rect 12390 8440 12395 8460
rect 12365 8410 12395 8440
rect 12365 8390 12370 8410
rect 12390 8390 12395 8410
rect 12365 8360 12395 8390
rect 12365 8340 12370 8360
rect 12390 8340 12395 8360
rect 12365 8310 12395 8340
rect 12365 8290 12370 8310
rect 12390 8290 12395 8310
rect 12365 8260 12395 8290
rect 12365 8240 12370 8260
rect 12390 8240 12395 8260
rect 12365 8210 12395 8240
rect 12365 8190 12370 8210
rect 12390 8190 12395 8210
rect 12365 8180 12395 8190
rect 12425 8560 12455 8570
rect 12425 8540 12430 8560
rect 12450 8540 12455 8560
rect 12425 8510 12455 8540
rect 12425 8490 12430 8510
rect 12450 8490 12455 8510
rect 12425 8460 12455 8490
rect 12425 8440 12430 8460
rect 12450 8440 12455 8460
rect 12425 8410 12455 8440
rect 12425 8390 12430 8410
rect 12450 8390 12455 8410
rect 12425 8360 12455 8390
rect 12425 8340 12430 8360
rect 12450 8340 12455 8360
rect 12425 8310 12455 8340
rect 12425 8290 12430 8310
rect 12450 8290 12455 8310
rect 12425 8260 12455 8290
rect 12425 8240 12430 8260
rect 12450 8240 12455 8260
rect 12425 8210 12455 8240
rect 12425 8190 12430 8210
rect 12450 8190 12455 8210
rect 12425 8180 12455 8190
rect 12485 8560 12515 8570
rect 12485 8540 12490 8560
rect 12510 8540 12515 8560
rect 12485 8510 12515 8540
rect 12485 8490 12490 8510
rect 12510 8490 12515 8510
rect 12485 8460 12515 8490
rect 12485 8440 12490 8460
rect 12510 8440 12515 8460
rect 12485 8410 12515 8440
rect 12485 8390 12490 8410
rect 12510 8390 12515 8410
rect 12485 8360 12515 8390
rect 12485 8340 12490 8360
rect 12510 8340 12515 8360
rect 12485 8310 12515 8340
rect 12485 8290 12490 8310
rect 12510 8290 12515 8310
rect 12485 8260 12515 8290
rect 12485 8240 12490 8260
rect 12510 8240 12515 8260
rect 12485 8210 12515 8240
rect 12485 8190 12490 8210
rect 12510 8190 12515 8210
rect 12485 8180 12515 8190
rect 12545 8560 12615 8570
rect 12545 8540 12550 8560
rect 12570 8540 12590 8560
rect 12610 8540 12615 8560
rect 18505 8565 18535 8575
rect 18505 8545 18510 8565
rect 18530 8545 18535 8565
rect 12545 8510 12615 8540
rect 12545 8490 12550 8510
rect 12570 8490 12590 8510
rect 12610 8490 12615 8510
rect 12545 8460 12615 8490
rect 12545 8440 12550 8460
rect 12570 8440 12590 8460
rect 12610 8440 12615 8460
rect 12545 8410 12615 8440
rect 12545 8390 12550 8410
rect 12570 8390 12590 8410
rect 12610 8390 12615 8410
rect 12545 8360 12615 8390
rect 12545 8340 12550 8360
rect 12570 8340 12590 8360
rect 12610 8340 12615 8360
rect 18285 8515 18355 8545
rect 18285 8495 18290 8515
rect 18310 8495 18330 8515
rect 18350 8495 18355 8515
rect 18285 8465 18355 8495
rect 18285 8445 18290 8465
rect 18310 8445 18330 8465
rect 18350 8445 18355 8465
rect 18285 8415 18355 8445
rect 18285 8395 18290 8415
rect 18310 8395 18330 8415
rect 18350 8395 18355 8415
rect 18285 8365 18355 8395
rect 12545 8310 12615 8340
rect 17950 8340 17990 8350
rect 17950 8320 17960 8340
rect 17980 8320 17990 8340
rect 17950 8310 17990 8320
rect 18210 8340 18250 8350
rect 18210 8320 18220 8340
rect 18240 8320 18250 8340
rect 18210 8310 18250 8320
rect 18285 8345 18290 8365
rect 18310 8345 18330 8365
rect 18350 8345 18355 8365
rect 18285 8315 18355 8345
rect 12545 8290 12550 8310
rect 12570 8290 12590 8310
rect 12610 8290 12615 8310
rect 12545 8260 12615 8290
rect 12545 8240 12550 8260
rect 12570 8240 12590 8260
rect 12610 8240 12615 8260
rect 12950 8285 12990 8295
rect 12950 8265 12960 8285
rect 12980 8265 12990 8285
rect 12950 8255 12990 8265
rect 13060 8285 13100 8295
rect 13060 8265 13070 8285
rect 13090 8265 13100 8285
rect 13060 8255 13100 8265
rect 13170 8285 13210 8295
rect 13170 8265 13180 8285
rect 13200 8265 13210 8285
rect 13170 8255 13210 8265
rect 13280 8285 13320 8295
rect 13280 8265 13290 8285
rect 13310 8265 13320 8285
rect 13280 8255 13320 8265
rect 13390 8285 13430 8295
rect 13390 8265 13400 8285
rect 13420 8265 13430 8285
rect 13390 8255 13430 8265
rect 13500 8285 13540 8295
rect 13500 8265 13510 8285
rect 13530 8265 13540 8285
rect 13500 8255 13540 8265
rect 13610 8285 13650 8295
rect 13610 8265 13620 8285
rect 13640 8265 13650 8285
rect 13610 8255 13650 8265
rect 13720 8285 13760 8295
rect 13720 8265 13730 8285
rect 13750 8265 13760 8285
rect 13720 8255 13760 8265
rect 13830 8285 13870 8295
rect 13830 8265 13840 8285
rect 13860 8265 13870 8285
rect 13830 8255 13870 8265
rect 13940 8285 13980 8295
rect 13940 8265 13950 8285
rect 13970 8265 13980 8285
rect 13940 8255 13980 8265
rect 14050 8285 14090 8295
rect 17960 8288 17980 8310
rect 18220 8288 18240 8310
rect 18285 8295 18290 8315
rect 18310 8295 18330 8315
rect 18350 8295 18355 8315
rect 14050 8265 14060 8285
rect 14080 8265 14090 8285
rect 14050 8255 14090 8265
rect 17955 8265 18025 8288
rect 12545 8210 12615 8240
rect 12960 8235 12980 8255
rect 13070 8235 13090 8255
rect 13180 8235 13200 8255
rect 13290 8235 13310 8255
rect 13400 8235 13420 8255
rect 13510 8235 13530 8255
rect 13620 8235 13640 8255
rect 13730 8235 13750 8255
rect 13840 8235 13860 8255
rect 13950 8235 13970 8255
rect 14060 8235 14080 8255
rect 17955 8245 17960 8265
rect 17980 8245 18000 8265
rect 18020 8245 18025 8265
rect 17955 8235 18025 8245
rect 18055 8270 18085 8288
rect 18055 8250 18060 8270
rect 18080 8250 18085 8270
rect 18055 8235 18085 8250
rect 18115 8270 18145 8288
rect 18115 8250 18120 8270
rect 18140 8250 18145 8270
rect 18115 8235 18145 8250
rect 18175 8265 18245 8288
rect 18175 8245 18180 8265
rect 18200 8245 18220 8265
rect 18240 8245 18245 8265
rect 18175 8235 18245 8245
rect 18285 8265 18355 8295
rect 18285 8245 18290 8265
rect 18310 8245 18330 8265
rect 18350 8245 18355 8265
rect 18285 8235 18355 8245
rect 18385 8515 18415 8545
rect 18385 8495 18390 8515
rect 18410 8495 18415 8515
rect 18385 8465 18415 8495
rect 18385 8445 18390 8465
rect 18410 8445 18415 8465
rect 18385 8415 18415 8445
rect 18385 8395 18390 8415
rect 18410 8395 18415 8415
rect 18385 8365 18415 8395
rect 18385 8345 18390 8365
rect 18410 8345 18415 8365
rect 18385 8315 18415 8345
rect 18385 8295 18390 8315
rect 18410 8295 18415 8315
rect 18385 8265 18415 8295
rect 18385 8245 18390 8265
rect 18410 8245 18415 8265
rect 18385 8235 18415 8245
rect 18445 8515 18475 8545
rect 18445 8495 18450 8515
rect 18470 8495 18475 8515
rect 18445 8465 18475 8495
rect 18445 8445 18450 8465
rect 18470 8445 18475 8465
rect 18445 8415 18475 8445
rect 18445 8395 18450 8415
rect 18470 8395 18475 8415
rect 18445 8365 18475 8395
rect 18445 8345 18450 8365
rect 18470 8345 18475 8365
rect 18445 8315 18475 8345
rect 18445 8295 18450 8315
rect 18470 8295 18475 8315
rect 18445 8265 18475 8295
rect 18445 8245 18450 8265
rect 18470 8245 18475 8265
rect 18445 8235 18475 8245
rect 18505 8515 18535 8545
rect 18505 8495 18510 8515
rect 18530 8495 18535 8515
rect 18505 8465 18535 8495
rect 18505 8445 18510 8465
rect 18530 8445 18535 8465
rect 18505 8415 18535 8445
rect 18505 8395 18510 8415
rect 18530 8395 18535 8415
rect 18505 8365 18535 8395
rect 18505 8345 18510 8365
rect 18530 8345 18535 8365
rect 18505 8315 18535 8345
rect 18505 8295 18510 8315
rect 18530 8295 18535 8315
rect 18505 8265 18535 8295
rect 18505 8245 18510 8265
rect 18530 8245 18535 8265
rect 18505 8235 18535 8245
rect 18565 8565 18635 8575
rect 18690 8570 18710 8590
rect 18850 8570 18870 8590
rect 18970 8570 18990 8590
rect 19090 8570 19110 8590
rect 19210 8570 19230 8590
rect 19330 8570 19350 8590
rect 19450 8570 19470 8590
rect 19570 8570 19590 8590
rect 19690 8570 19710 8590
rect 19810 8570 19830 8590
rect 19930 8570 19950 8590
rect 20090 8570 20110 8590
rect 18565 8545 18570 8565
rect 18590 8545 18610 8565
rect 18630 8545 18635 8565
rect 18565 8515 18635 8545
rect 18565 8495 18570 8515
rect 18590 8495 18610 8515
rect 18630 8495 18635 8515
rect 18565 8465 18635 8495
rect 18565 8445 18570 8465
rect 18590 8445 18610 8465
rect 18630 8445 18635 8465
rect 18565 8415 18635 8445
rect 18565 8395 18570 8415
rect 18590 8395 18610 8415
rect 18630 8395 18635 8415
rect 18565 8365 18635 8395
rect 18565 8345 18570 8365
rect 18590 8345 18610 8365
rect 18630 8345 18635 8365
rect 18565 8315 18635 8345
rect 18565 8295 18570 8315
rect 18590 8295 18610 8315
rect 18630 8295 18635 8315
rect 18565 8265 18635 8295
rect 18565 8245 18570 8265
rect 18590 8245 18610 8265
rect 18630 8245 18635 8265
rect 18565 8235 18635 8245
rect 18685 8560 18755 8570
rect 18685 8540 18690 8560
rect 18710 8540 18730 8560
rect 18750 8540 18755 8560
rect 18685 8510 18755 8540
rect 18685 8490 18690 8510
rect 18710 8490 18730 8510
rect 18750 8490 18755 8510
rect 18685 8460 18755 8490
rect 18685 8440 18690 8460
rect 18710 8440 18730 8460
rect 18750 8440 18755 8460
rect 18685 8410 18755 8440
rect 18685 8390 18690 8410
rect 18710 8390 18730 8410
rect 18750 8390 18755 8410
rect 18685 8360 18755 8390
rect 18685 8340 18690 8360
rect 18710 8340 18730 8360
rect 18750 8340 18755 8360
rect 18685 8310 18755 8340
rect 18685 8290 18690 8310
rect 18710 8290 18730 8310
rect 18750 8290 18755 8310
rect 18685 8260 18755 8290
rect 18685 8240 18690 8260
rect 18710 8240 18730 8260
rect 18750 8240 18755 8260
rect 12545 8190 12550 8210
rect 12570 8190 12590 8210
rect 12610 8190 12615 8210
rect 12545 8180 12615 8190
rect 12860 8225 12930 8235
rect 12860 8205 12865 8225
rect 12885 8205 12905 8225
rect 12925 8205 12930 8225
rect 11290 8160 11310 8180
rect 11410 8160 11430 8180
rect 11530 8160 11550 8180
rect 11650 8160 11670 8180
rect 11770 8160 11790 8180
rect 11890 8160 11910 8180
rect 12010 8160 12030 8180
rect 12130 8160 12150 8180
rect 12250 8160 12270 8180
rect 12370 8160 12390 8180
rect 12490 8160 12510 8180
rect 12860 8175 12930 8205
rect 11280 8150 11320 8160
rect 11280 8130 11290 8150
rect 11310 8130 11320 8150
rect 11280 8120 11320 8130
rect 11400 8150 11440 8160
rect 11400 8130 11410 8150
rect 11430 8130 11440 8150
rect 11400 8120 11440 8130
rect 11520 8150 11560 8160
rect 11520 8130 11530 8150
rect 11550 8130 11560 8150
rect 11520 8120 11560 8130
rect 11640 8150 11680 8160
rect 11640 8130 11650 8150
rect 11670 8130 11680 8150
rect 11640 8120 11680 8130
rect 11760 8150 11800 8160
rect 11760 8130 11770 8150
rect 11790 8130 11800 8150
rect 11760 8120 11800 8130
rect 11823 8150 11857 8160
rect 11823 8130 11831 8150
rect 11849 8130 11857 8150
rect 11823 8120 11857 8130
rect 11880 8150 11920 8160
rect 11880 8130 11890 8150
rect 11910 8130 11920 8150
rect 11880 8120 11920 8130
rect 12000 8150 12040 8160
rect 12000 8130 12010 8150
rect 12030 8130 12040 8150
rect 12000 8120 12040 8130
rect 12120 8150 12160 8160
rect 12120 8130 12130 8150
rect 12150 8130 12160 8150
rect 12120 8120 12160 8130
rect 12240 8150 12280 8160
rect 12240 8130 12250 8150
rect 12270 8130 12280 8150
rect 12240 8120 12280 8130
rect 12360 8150 12400 8160
rect 12360 8130 12370 8150
rect 12390 8130 12400 8150
rect 12360 8120 12400 8130
rect 12480 8150 12520 8160
rect 12480 8130 12490 8150
rect 12510 8130 12520 8150
rect 12480 8120 12520 8130
rect 12860 8155 12865 8175
rect 12885 8155 12905 8175
rect 12925 8155 12930 8175
rect 12860 8125 12930 8155
rect 12860 8105 12865 8125
rect 12885 8105 12905 8125
rect 12925 8105 12930 8125
rect 12860 8075 12930 8105
rect 12860 8055 12865 8075
rect 12885 8055 12905 8075
rect 12925 8055 12930 8075
rect 12860 8025 12930 8055
rect 12860 8005 12865 8025
rect 12885 8005 12905 8025
rect 12925 8005 12930 8025
rect 12860 7975 12930 8005
rect 12860 7955 12865 7975
rect 12885 7955 12905 7975
rect 12925 7955 12930 7975
rect 11180 7940 11220 7950
rect 11180 7920 11190 7940
rect 11210 7920 11220 7940
rect 11180 7910 11220 7920
rect 11340 7940 11380 7950
rect 11340 7920 11350 7940
rect 11370 7920 11380 7940
rect 11340 7910 11380 7920
rect 11460 7940 11500 7950
rect 11460 7920 11470 7940
rect 11490 7920 11500 7940
rect 11460 7910 11500 7920
rect 11580 7940 11620 7950
rect 11580 7920 11590 7940
rect 11610 7920 11620 7940
rect 11580 7910 11620 7920
rect 11700 7940 11740 7950
rect 11700 7920 11710 7940
rect 11730 7920 11740 7940
rect 11700 7910 11740 7920
rect 11820 7940 11860 7950
rect 11820 7920 11830 7940
rect 11850 7920 11860 7940
rect 11820 7910 11860 7920
rect 11940 7940 11980 7950
rect 11940 7920 11950 7940
rect 11970 7920 11980 7940
rect 11940 7910 11980 7920
rect 12060 7940 12100 7950
rect 12060 7920 12070 7940
rect 12090 7920 12100 7940
rect 12060 7910 12100 7920
rect 12180 7940 12220 7950
rect 12180 7920 12190 7940
rect 12210 7920 12220 7940
rect 12180 7910 12220 7920
rect 12300 7940 12340 7950
rect 12300 7920 12310 7940
rect 12330 7920 12340 7940
rect 12300 7910 12340 7920
rect 12420 7940 12460 7950
rect 12420 7920 12430 7940
rect 12450 7920 12460 7940
rect 12420 7910 12460 7920
rect 12480 7910 12520 7950
rect 12580 7940 12620 7950
rect 12860 7945 12930 7955
rect 12955 8225 12985 8235
rect 12955 8205 12960 8225
rect 12980 8205 12985 8225
rect 12955 8175 12985 8205
rect 12955 8155 12960 8175
rect 12980 8155 12985 8175
rect 12955 8125 12985 8155
rect 12955 8105 12960 8125
rect 12980 8105 12985 8125
rect 12955 8075 12985 8105
rect 12955 8055 12960 8075
rect 12980 8055 12985 8075
rect 12955 8025 12985 8055
rect 12955 8005 12960 8025
rect 12980 8005 12985 8025
rect 12955 7975 12985 8005
rect 12955 7955 12960 7975
rect 12980 7955 12985 7975
rect 12955 7945 12985 7955
rect 13010 8225 13040 8235
rect 13010 8205 13015 8225
rect 13035 8205 13040 8225
rect 13010 8175 13040 8205
rect 13010 8155 13015 8175
rect 13035 8155 13040 8175
rect 13010 8125 13040 8155
rect 13010 8105 13015 8125
rect 13035 8105 13040 8125
rect 13010 8075 13040 8105
rect 13010 8055 13015 8075
rect 13035 8055 13040 8075
rect 13010 8025 13040 8055
rect 13010 8005 13015 8025
rect 13035 8005 13040 8025
rect 13010 7975 13040 8005
rect 13010 7955 13015 7975
rect 13035 7955 13040 7975
rect 13010 7945 13040 7955
rect 13065 8225 13095 8235
rect 13065 8205 13070 8225
rect 13090 8205 13095 8225
rect 13065 8175 13095 8205
rect 13065 8155 13070 8175
rect 13090 8155 13095 8175
rect 13065 8125 13095 8155
rect 13065 8105 13070 8125
rect 13090 8105 13095 8125
rect 13065 8075 13095 8105
rect 13065 8055 13070 8075
rect 13090 8055 13095 8075
rect 13065 8025 13095 8055
rect 13065 8005 13070 8025
rect 13090 8005 13095 8025
rect 13065 7975 13095 8005
rect 13065 7955 13070 7975
rect 13090 7955 13095 7975
rect 13065 7945 13095 7955
rect 13120 8225 13150 8235
rect 13120 8205 13125 8225
rect 13145 8205 13150 8225
rect 13120 8175 13150 8205
rect 13120 8155 13125 8175
rect 13145 8155 13150 8175
rect 13120 8125 13150 8155
rect 13120 8105 13125 8125
rect 13145 8105 13150 8125
rect 13120 8075 13150 8105
rect 13120 8055 13125 8075
rect 13145 8055 13150 8075
rect 13120 8025 13150 8055
rect 13120 8005 13125 8025
rect 13145 8005 13150 8025
rect 13120 7975 13150 8005
rect 13120 7955 13125 7975
rect 13145 7955 13150 7975
rect 13120 7945 13150 7955
rect 13175 8225 13205 8235
rect 13175 8205 13180 8225
rect 13200 8205 13205 8225
rect 13175 8175 13205 8205
rect 13175 8155 13180 8175
rect 13200 8155 13205 8175
rect 13175 8125 13205 8155
rect 13175 8105 13180 8125
rect 13200 8105 13205 8125
rect 13175 8075 13205 8105
rect 13175 8055 13180 8075
rect 13200 8055 13205 8075
rect 13175 8025 13205 8055
rect 13175 8005 13180 8025
rect 13200 8005 13205 8025
rect 13175 7975 13205 8005
rect 13175 7955 13180 7975
rect 13200 7955 13205 7975
rect 13175 7945 13205 7955
rect 13230 8225 13260 8235
rect 13230 8205 13235 8225
rect 13255 8205 13260 8225
rect 13230 8175 13260 8205
rect 13230 8155 13235 8175
rect 13255 8155 13260 8175
rect 13230 8125 13260 8155
rect 13230 8105 13235 8125
rect 13255 8105 13260 8125
rect 13230 8075 13260 8105
rect 13230 8055 13235 8075
rect 13255 8055 13260 8075
rect 13230 8025 13260 8055
rect 13230 8005 13235 8025
rect 13255 8005 13260 8025
rect 13230 7975 13260 8005
rect 13230 7955 13235 7975
rect 13255 7955 13260 7975
rect 13230 7945 13260 7955
rect 13285 8225 13315 8235
rect 13285 8205 13290 8225
rect 13310 8205 13315 8225
rect 13285 8175 13315 8205
rect 13285 8155 13290 8175
rect 13310 8155 13315 8175
rect 13285 8125 13315 8155
rect 13285 8105 13290 8125
rect 13310 8105 13315 8125
rect 13285 8075 13315 8105
rect 13285 8055 13290 8075
rect 13310 8055 13315 8075
rect 13285 8025 13315 8055
rect 13285 8005 13290 8025
rect 13310 8005 13315 8025
rect 13285 7975 13315 8005
rect 13285 7955 13290 7975
rect 13310 7955 13315 7975
rect 13285 7945 13315 7955
rect 13340 8225 13370 8235
rect 13340 8205 13345 8225
rect 13365 8205 13370 8225
rect 13340 8175 13370 8205
rect 13340 8155 13345 8175
rect 13365 8155 13370 8175
rect 13340 8125 13370 8155
rect 13340 8105 13345 8125
rect 13365 8105 13370 8125
rect 13340 8075 13370 8105
rect 13340 8055 13345 8075
rect 13365 8055 13370 8075
rect 13340 8025 13370 8055
rect 13340 8005 13345 8025
rect 13365 8005 13370 8025
rect 13340 7975 13370 8005
rect 13340 7955 13345 7975
rect 13365 7955 13370 7975
rect 13340 7945 13370 7955
rect 13395 8225 13425 8235
rect 13395 8205 13400 8225
rect 13420 8205 13425 8225
rect 13395 8175 13425 8205
rect 13395 8155 13400 8175
rect 13420 8155 13425 8175
rect 13395 8125 13425 8155
rect 13395 8105 13400 8125
rect 13420 8105 13425 8125
rect 13395 8075 13425 8105
rect 13395 8055 13400 8075
rect 13420 8055 13425 8075
rect 13395 8025 13425 8055
rect 13395 8005 13400 8025
rect 13420 8005 13425 8025
rect 13395 7975 13425 8005
rect 13395 7955 13400 7975
rect 13420 7955 13425 7975
rect 13395 7945 13425 7955
rect 13450 8225 13480 8235
rect 13450 8205 13455 8225
rect 13475 8205 13480 8225
rect 13450 8175 13480 8205
rect 13450 8155 13455 8175
rect 13475 8155 13480 8175
rect 13450 8125 13480 8155
rect 13450 8105 13455 8125
rect 13475 8105 13480 8125
rect 13450 8075 13480 8105
rect 13450 8055 13455 8075
rect 13475 8055 13480 8075
rect 13450 8025 13480 8055
rect 13450 8005 13455 8025
rect 13475 8005 13480 8025
rect 13450 7975 13480 8005
rect 13450 7955 13455 7975
rect 13475 7955 13480 7975
rect 13450 7945 13480 7955
rect 13505 8225 13535 8235
rect 13505 8205 13510 8225
rect 13530 8205 13535 8225
rect 13505 8175 13535 8205
rect 13505 8155 13510 8175
rect 13530 8155 13535 8175
rect 13505 8125 13535 8155
rect 13505 8105 13510 8125
rect 13530 8105 13535 8125
rect 13505 8075 13535 8105
rect 13505 8055 13510 8075
rect 13530 8055 13535 8075
rect 13505 8025 13535 8055
rect 13505 8005 13510 8025
rect 13530 8005 13535 8025
rect 13505 7975 13535 8005
rect 13505 7955 13510 7975
rect 13530 7955 13535 7975
rect 13505 7945 13535 7955
rect 13560 8225 13590 8235
rect 13560 8205 13565 8225
rect 13585 8205 13590 8225
rect 13560 8175 13590 8205
rect 13560 8155 13565 8175
rect 13585 8155 13590 8175
rect 13560 8125 13590 8155
rect 13560 8105 13565 8125
rect 13585 8105 13590 8125
rect 13560 8075 13590 8105
rect 13560 8055 13565 8075
rect 13585 8055 13590 8075
rect 13560 8025 13590 8055
rect 13560 8005 13565 8025
rect 13585 8005 13590 8025
rect 13560 7975 13590 8005
rect 13560 7955 13565 7975
rect 13585 7955 13590 7975
rect 13560 7945 13590 7955
rect 13615 8225 13645 8235
rect 13615 8205 13620 8225
rect 13640 8205 13645 8225
rect 13615 8175 13645 8205
rect 13615 8155 13620 8175
rect 13640 8155 13645 8175
rect 13615 8125 13645 8155
rect 13615 8105 13620 8125
rect 13640 8105 13645 8125
rect 13615 8075 13645 8105
rect 13615 8055 13620 8075
rect 13640 8055 13645 8075
rect 13615 8025 13645 8055
rect 13615 8005 13620 8025
rect 13640 8005 13645 8025
rect 13615 7975 13645 8005
rect 13615 7955 13620 7975
rect 13640 7955 13645 7975
rect 13615 7945 13645 7955
rect 13670 8225 13700 8235
rect 13670 8205 13675 8225
rect 13695 8205 13700 8225
rect 13670 8175 13700 8205
rect 13670 8155 13675 8175
rect 13695 8155 13700 8175
rect 13670 8125 13700 8155
rect 13670 8105 13675 8125
rect 13695 8105 13700 8125
rect 13670 8075 13700 8105
rect 13670 8055 13675 8075
rect 13695 8055 13700 8075
rect 13670 8025 13700 8055
rect 13670 8005 13675 8025
rect 13695 8005 13700 8025
rect 13670 7975 13700 8005
rect 13670 7955 13675 7975
rect 13695 7955 13700 7975
rect 13670 7945 13700 7955
rect 13725 8225 13755 8235
rect 13725 8205 13730 8225
rect 13750 8205 13755 8225
rect 13725 8175 13755 8205
rect 13725 8155 13730 8175
rect 13750 8155 13755 8175
rect 13725 8125 13755 8155
rect 13725 8105 13730 8125
rect 13750 8105 13755 8125
rect 13725 8075 13755 8105
rect 13725 8055 13730 8075
rect 13750 8055 13755 8075
rect 13725 8025 13755 8055
rect 13725 8005 13730 8025
rect 13750 8005 13755 8025
rect 13725 7975 13755 8005
rect 13725 7955 13730 7975
rect 13750 7955 13755 7975
rect 13725 7945 13755 7955
rect 13780 8225 13810 8235
rect 13780 8205 13785 8225
rect 13805 8205 13810 8225
rect 13780 8175 13810 8205
rect 13780 8155 13785 8175
rect 13805 8155 13810 8175
rect 13780 8125 13810 8155
rect 13780 8105 13785 8125
rect 13805 8105 13810 8125
rect 13780 8075 13810 8105
rect 13780 8055 13785 8075
rect 13805 8055 13810 8075
rect 13780 8025 13810 8055
rect 13780 8005 13785 8025
rect 13805 8005 13810 8025
rect 13780 7975 13810 8005
rect 13780 7955 13785 7975
rect 13805 7955 13810 7975
rect 13780 7945 13810 7955
rect 13835 8225 13865 8235
rect 13835 8205 13840 8225
rect 13860 8205 13865 8225
rect 13835 8175 13865 8205
rect 13835 8155 13840 8175
rect 13860 8155 13865 8175
rect 13835 8125 13865 8155
rect 13835 8105 13840 8125
rect 13860 8105 13865 8125
rect 13835 8075 13865 8105
rect 13835 8055 13840 8075
rect 13860 8055 13865 8075
rect 13835 8025 13865 8055
rect 13835 8005 13840 8025
rect 13860 8005 13865 8025
rect 13835 7975 13865 8005
rect 13835 7955 13840 7975
rect 13860 7955 13865 7975
rect 13835 7945 13865 7955
rect 13890 8225 13920 8235
rect 13890 8205 13895 8225
rect 13915 8205 13920 8225
rect 13890 8175 13920 8205
rect 13890 8155 13895 8175
rect 13915 8155 13920 8175
rect 13890 8125 13920 8155
rect 13890 8105 13895 8125
rect 13915 8105 13920 8125
rect 13890 8075 13920 8105
rect 13890 8055 13895 8075
rect 13915 8055 13920 8075
rect 13890 8025 13920 8055
rect 13890 8005 13895 8025
rect 13915 8005 13920 8025
rect 13890 7975 13920 8005
rect 13890 7955 13895 7975
rect 13915 7955 13920 7975
rect 13890 7945 13920 7955
rect 13945 8225 13975 8235
rect 13945 8205 13950 8225
rect 13970 8205 13975 8225
rect 13945 8175 13975 8205
rect 13945 8155 13950 8175
rect 13970 8155 13975 8175
rect 13945 8125 13975 8155
rect 13945 8105 13950 8125
rect 13970 8105 13975 8125
rect 13945 8075 13975 8105
rect 13945 8055 13950 8075
rect 13970 8055 13975 8075
rect 13945 8025 13975 8055
rect 13945 8005 13950 8025
rect 13970 8005 13975 8025
rect 13945 7975 13975 8005
rect 13945 7955 13950 7975
rect 13970 7955 13975 7975
rect 13945 7945 13975 7955
rect 14000 8225 14030 8235
rect 14000 8205 14005 8225
rect 14025 8205 14030 8225
rect 14000 8175 14030 8205
rect 14000 8155 14005 8175
rect 14025 8155 14030 8175
rect 14000 8125 14030 8155
rect 14000 8105 14005 8125
rect 14025 8105 14030 8125
rect 14000 8075 14030 8105
rect 14000 8055 14005 8075
rect 14025 8055 14030 8075
rect 14000 8025 14030 8055
rect 14000 8005 14005 8025
rect 14025 8005 14030 8025
rect 14000 7975 14030 8005
rect 14000 7955 14005 7975
rect 14025 7955 14030 7975
rect 14000 7945 14030 7955
rect 14055 8225 14085 8235
rect 14055 8205 14060 8225
rect 14080 8205 14085 8225
rect 14055 8175 14085 8205
rect 14055 8155 14060 8175
rect 14080 8155 14085 8175
rect 14055 8125 14085 8155
rect 14055 8105 14060 8125
rect 14080 8105 14085 8125
rect 14055 8075 14085 8105
rect 14055 8055 14060 8075
rect 14080 8055 14085 8075
rect 14055 8025 14085 8055
rect 14055 8005 14060 8025
rect 14080 8005 14085 8025
rect 14055 7975 14085 8005
rect 14055 7955 14060 7975
rect 14080 7955 14085 7975
rect 14055 7945 14085 7955
rect 14110 8225 14180 8235
rect 14110 8205 14115 8225
rect 14135 8205 14155 8225
rect 14175 8205 14180 8225
rect 18120 8215 18140 8235
rect 18290 8215 18310 8235
rect 18610 8215 18630 8235
rect 14110 8175 14180 8205
rect 18080 8205 18140 8215
rect 18080 8185 18090 8205
rect 18110 8195 18140 8205
rect 18280 8205 18320 8215
rect 18110 8185 18120 8195
rect 18080 8175 18120 8185
rect 18280 8185 18290 8205
rect 18310 8185 18320 8205
rect 18280 8175 18320 8185
rect 18405 8205 18440 8215
rect 18405 8185 18410 8205
rect 18430 8185 18440 8205
rect 18405 8175 18440 8185
rect 18480 8205 18515 8215
rect 18480 8185 18490 8205
rect 18510 8185 18515 8205
rect 18480 8175 18515 8185
rect 18600 8205 18640 8215
rect 18600 8185 18610 8205
rect 18630 8185 18640 8205
rect 18600 8175 18640 8185
rect 18685 8210 18755 8240
rect 18685 8190 18690 8210
rect 18710 8190 18730 8210
rect 18750 8190 18755 8210
rect 18685 8180 18755 8190
rect 18785 8560 18815 8570
rect 18785 8540 18790 8560
rect 18810 8540 18815 8560
rect 18785 8510 18815 8540
rect 18785 8490 18790 8510
rect 18810 8490 18815 8510
rect 18785 8460 18815 8490
rect 18785 8440 18790 8460
rect 18810 8440 18815 8460
rect 18785 8410 18815 8440
rect 18785 8390 18790 8410
rect 18810 8390 18815 8410
rect 18785 8360 18815 8390
rect 18785 8340 18790 8360
rect 18810 8340 18815 8360
rect 18785 8310 18815 8340
rect 18785 8290 18790 8310
rect 18810 8290 18815 8310
rect 18785 8260 18815 8290
rect 18785 8240 18790 8260
rect 18810 8240 18815 8260
rect 18785 8210 18815 8240
rect 18785 8190 18790 8210
rect 18810 8190 18815 8210
rect 18785 8180 18815 8190
rect 18845 8560 18875 8570
rect 18845 8540 18850 8560
rect 18870 8540 18875 8560
rect 18845 8510 18875 8540
rect 18845 8490 18850 8510
rect 18870 8490 18875 8510
rect 18845 8460 18875 8490
rect 18845 8440 18850 8460
rect 18870 8440 18875 8460
rect 18845 8410 18875 8440
rect 18845 8390 18850 8410
rect 18870 8390 18875 8410
rect 18845 8360 18875 8390
rect 18845 8340 18850 8360
rect 18870 8340 18875 8360
rect 18845 8310 18875 8340
rect 18845 8290 18850 8310
rect 18870 8290 18875 8310
rect 18845 8260 18875 8290
rect 18845 8240 18850 8260
rect 18870 8240 18875 8260
rect 18845 8210 18875 8240
rect 18845 8190 18850 8210
rect 18870 8190 18875 8210
rect 18845 8180 18875 8190
rect 18905 8560 18935 8570
rect 18905 8540 18910 8560
rect 18930 8540 18935 8560
rect 18905 8510 18935 8540
rect 18905 8490 18910 8510
rect 18930 8490 18935 8510
rect 18905 8460 18935 8490
rect 18905 8440 18910 8460
rect 18930 8440 18935 8460
rect 18905 8410 18935 8440
rect 18905 8390 18910 8410
rect 18930 8390 18935 8410
rect 18905 8360 18935 8390
rect 18905 8340 18910 8360
rect 18930 8340 18935 8360
rect 18905 8310 18935 8340
rect 18905 8290 18910 8310
rect 18930 8290 18935 8310
rect 18905 8260 18935 8290
rect 18905 8240 18910 8260
rect 18930 8240 18935 8260
rect 18905 8210 18935 8240
rect 18905 8190 18910 8210
rect 18930 8190 18935 8210
rect 18905 8180 18935 8190
rect 18965 8560 18995 8570
rect 18965 8540 18970 8560
rect 18990 8540 18995 8560
rect 18965 8510 18995 8540
rect 18965 8490 18970 8510
rect 18990 8490 18995 8510
rect 18965 8460 18995 8490
rect 18965 8440 18970 8460
rect 18990 8440 18995 8460
rect 18965 8410 18995 8440
rect 18965 8390 18970 8410
rect 18990 8390 18995 8410
rect 18965 8360 18995 8390
rect 18965 8340 18970 8360
rect 18990 8340 18995 8360
rect 18965 8310 18995 8340
rect 18965 8290 18970 8310
rect 18990 8290 18995 8310
rect 18965 8260 18995 8290
rect 18965 8240 18970 8260
rect 18990 8240 18995 8260
rect 18965 8210 18995 8240
rect 18965 8190 18970 8210
rect 18990 8190 18995 8210
rect 18965 8180 18995 8190
rect 19025 8560 19055 8570
rect 19025 8540 19030 8560
rect 19050 8540 19055 8560
rect 19025 8510 19055 8540
rect 19025 8490 19030 8510
rect 19050 8490 19055 8510
rect 19025 8460 19055 8490
rect 19025 8440 19030 8460
rect 19050 8440 19055 8460
rect 19025 8410 19055 8440
rect 19025 8390 19030 8410
rect 19050 8390 19055 8410
rect 19025 8360 19055 8390
rect 19025 8340 19030 8360
rect 19050 8340 19055 8360
rect 19025 8310 19055 8340
rect 19025 8290 19030 8310
rect 19050 8290 19055 8310
rect 19025 8260 19055 8290
rect 19025 8240 19030 8260
rect 19050 8240 19055 8260
rect 19025 8210 19055 8240
rect 19025 8190 19030 8210
rect 19050 8190 19055 8210
rect 19025 8180 19055 8190
rect 19085 8560 19115 8570
rect 19085 8540 19090 8560
rect 19110 8540 19115 8560
rect 19085 8510 19115 8540
rect 19085 8490 19090 8510
rect 19110 8490 19115 8510
rect 19085 8460 19115 8490
rect 19085 8440 19090 8460
rect 19110 8440 19115 8460
rect 19085 8410 19115 8440
rect 19085 8390 19090 8410
rect 19110 8390 19115 8410
rect 19085 8360 19115 8390
rect 19085 8340 19090 8360
rect 19110 8340 19115 8360
rect 19085 8310 19115 8340
rect 19085 8290 19090 8310
rect 19110 8290 19115 8310
rect 19085 8260 19115 8290
rect 19085 8240 19090 8260
rect 19110 8240 19115 8260
rect 19085 8210 19115 8240
rect 19085 8190 19090 8210
rect 19110 8190 19115 8210
rect 19085 8180 19115 8190
rect 19145 8560 19175 8570
rect 19145 8540 19150 8560
rect 19170 8540 19175 8560
rect 19145 8510 19175 8540
rect 19145 8490 19150 8510
rect 19170 8490 19175 8510
rect 19145 8460 19175 8490
rect 19145 8440 19150 8460
rect 19170 8440 19175 8460
rect 19145 8410 19175 8440
rect 19145 8390 19150 8410
rect 19170 8390 19175 8410
rect 19145 8360 19175 8390
rect 19145 8340 19150 8360
rect 19170 8340 19175 8360
rect 19145 8310 19175 8340
rect 19145 8290 19150 8310
rect 19170 8290 19175 8310
rect 19145 8260 19175 8290
rect 19145 8240 19150 8260
rect 19170 8240 19175 8260
rect 19145 8210 19175 8240
rect 19145 8190 19150 8210
rect 19170 8190 19175 8210
rect 19145 8180 19175 8190
rect 19205 8560 19235 8570
rect 19205 8540 19210 8560
rect 19230 8540 19235 8560
rect 19205 8510 19235 8540
rect 19205 8490 19210 8510
rect 19230 8490 19235 8510
rect 19205 8460 19235 8490
rect 19205 8440 19210 8460
rect 19230 8440 19235 8460
rect 19205 8410 19235 8440
rect 19205 8390 19210 8410
rect 19230 8390 19235 8410
rect 19205 8360 19235 8390
rect 19205 8340 19210 8360
rect 19230 8340 19235 8360
rect 19205 8310 19235 8340
rect 19205 8290 19210 8310
rect 19230 8290 19235 8310
rect 19205 8260 19235 8290
rect 19205 8240 19210 8260
rect 19230 8240 19235 8260
rect 19205 8210 19235 8240
rect 19205 8190 19210 8210
rect 19230 8190 19235 8210
rect 19205 8180 19235 8190
rect 19265 8560 19295 8570
rect 19265 8540 19270 8560
rect 19290 8540 19295 8560
rect 19265 8510 19295 8540
rect 19265 8490 19270 8510
rect 19290 8490 19295 8510
rect 19265 8460 19295 8490
rect 19265 8440 19270 8460
rect 19290 8440 19295 8460
rect 19265 8410 19295 8440
rect 19265 8390 19270 8410
rect 19290 8390 19295 8410
rect 19265 8360 19295 8390
rect 19265 8340 19270 8360
rect 19290 8340 19295 8360
rect 19265 8310 19295 8340
rect 19265 8290 19270 8310
rect 19290 8290 19295 8310
rect 19265 8260 19295 8290
rect 19265 8240 19270 8260
rect 19290 8240 19295 8260
rect 19265 8210 19295 8240
rect 19265 8190 19270 8210
rect 19290 8190 19295 8210
rect 19265 8180 19295 8190
rect 19325 8560 19355 8570
rect 19325 8540 19330 8560
rect 19350 8540 19355 8560
rect 19325 8510 19355 8540
rect 19325 8490 19330 8510
rect 19350 8490 19355 8510
rect 19325 8460 19355 8490
rect 19325 8440 19330 8460
rect 19350 8440 19355 8460
rect 19325 8410 19355 8440
rect 19325 8390 19330 8410
rect 19350 8390 19355 8410
rect 19325 8360 19355 8390
rect 19325 8340 19330 8360
rect 19350 8340 19355 8360
rect 19325 8310 19355 8340
rect 19325 8290 19330 8310
rect 19350 8290 19355 8310
rect 19325 8260 19355 8290
rect 19325 8240 19330 8260
rect 19350 8240 19355 8260
rect 19325 8210 19355 8240
rect 19325 8190 19330 8210
rect 19350 8190 19355 8210
rect 19325 8180 19355 8190
rect 19385 8560 19415 8570
rect 19385 8540 19390 8560
rect 19410 8540 19415 8560
rect 19385 8510 19415 8540
rect 19385 8490 19390 8510
rect 19410 8490 19415 8510
rect 19385 8460 19415 8490
rect 19385 8440 19390 8460
rect 19410 8440 19415 8460
rect 19385 8410 19415 8440
rect 19385 8390 19390 8410
rect 19410 8390 19415 8410
rect 19385 8360 19415 8390
rect 19385 8340 19390 8360
rect 19410 8340 19415 8360
rect 19385 8310 19415 8340
rect 19385 8290 19390 8310
rect 19410 8290 19415 8310
rect 19385 8260 19415 8290
rect 19385 8240 19390 8260
rect 19410 8240 19415 8260
rect 19385 8210 19415 8240
rect 19385 8190 19390 8210
rect 19410 8190 19415 8210
rect 19385 8180 19415 8190
rect 19445 8560 19475 8570
rect 19445 8540 19450 8560
rect 19470 8540 19475 8560
rect 19445 8510 19475 8540
rect 19445 8490 19450 8510
rect 19470 8490 19475 8510
rect 19445 8460 19475 8490
rect 19445 8440 19450 8460
rect 19470 8440 19475 8460
rect 19445 8410 19475 8440
rect 19445 8390 19450 8410
rect 19470 8390 19475 8410
rect 19445 8360 19475 8390
rect 19445 8340 19450 8360
rect 19470 8340 19475 8360
rect 19445 8310 19475 8340
rect 19445 8290 19450 8310
rect 19470 8290 19475 8310
rect 19445 8260 19475 8290
rect 19445 8240 19450 8260
rect 19470 8240 19475 8260
rect 19445 8210 19475 8240
rect 19445 8190 19450 8210
rect 19470 8190 19475 8210
rect 19445 8180 19475 8190
rect 19505 8560 19535 8570
rect 19505 8540 19510 8560
rect 19530 8540 19535 8560
rect 19505 8510 19535 8540
rect 19505 8490 19510 8510
rect 19530 8490 19535 8510
rect 19505 8460 19535 8490
rect 19505 8440 19510 8460
rect 19530 8440 19535 8460
rect 19505 8410 19535 8440
rect 19505 8390 19510 8410
rect 19530 8390 19535 8410
rect 19505 8360 19535 8390
rect 19505 8340 19510 8360
rect 19530 8340 19535 8360
rect 19505 8310 19535 8340
rect 19505 8290 19510 8310
rect 19530 8290 19535 8310
rect 19505 8260 19535 8290
rect 19505 8240 19510 8260
rect 19530 8240 19535 8260
rect 19505 8210 19535 8240
rect 19505 8190 19510 8210
rect 19530 8190 19535 8210
rect 19505 8180 19535 8190
rect 19565 8560 19595 8570
rect 19565 8540 19570 8560
rect 19590 8540 19595 8560
rect 19565 8510 19595 8540
rect 19565 8490 19570 8510
rect 19590 8490 19595 8510
rect 19565 8460 19595 8490
rect 19565 8440 19570 8460
rect 19590 8440 19595 8460
rect 19565 8410 19595 8440
rect 19565 8390 19570 8410
rect 19590 8390 19595 8410
rect 19565 8360 19595 8390
rect 19565 8340 19570 8360
rect 19590 8340 19595 8360
rect 19565 8310 19595 8340
rect 19565 8290 19570 8310
rect 19590 8290 19595 8310
rect 19565 8260 19595 8290
rect 19565 8240 19570 8260
rect 19590 8240 19595 8260
rect 19565 8210 19595 8240
rect 19565 8190 19570 8210
rect 19590 8190 19595 8210
rect 19565 8180 19595 8190
rect 19625 8560 19655 8570
rect 19625 8540 19630 8560
rect 19650 8540 19655 8560
rect 19625 8510 19655 8540
rect 19625 8490 19630 8510
rect 19650 8490 19655 8510
rect 19625 8460 19655 8490
rect 19625 8440 19630 8460
rect 19650 8440 19655 8460
rect 19625 8410 19655 8440
rect 19625 8390 19630 8410
rect 19650 8390 19655 8410
rect 19625 8360 19655 8390
rect 19625 8340 19630 8360
rect 19650 8340 19655 8360
rect 19625 8310 19655 8340
rect 19625 8290 19630 8310
rect 19650 8290 19655 8310
rect 19625 8260 19655 8290
rect 19625 8240 19630 8260
rect 19650 8240 19655 8260
rect 19625 8210 19655 8240
rect 19625 8190 19630 8210
rect 19650 8190 19655 8210
rect 19625 8180 19655 8190
rect 19685 8560 19715 8570
rect 19685 8540 19690 8560
rect 19710 8540 19715 8560
rect 19685 8510 19715 8540
rect 19685 8490 19690 8510
rect 19710 8490 19715 8510
rect 19685 8460 19715 8490
rect 19685 8440 19690 8460
rect 19710 8440 19715 8460
rect 19685 8410 19715 8440
rect 19685 8390 19690 8410
rect 19710 8390 19715 8410
rect 19685 8360 19715 8390
rect 19685 8340 19690 8360
rect 19710 8340 19715 8360
rect 19685 8310 19715 8340
rect 19685 8290 19690 8310
rect 19710 8290 19715 8310
rect 19685 8260 19715 8290
rect 19685 8240 19690 8260
rect 19710 8240 19715 8260
rect 19685 8210 19715 8240
rect 19685 8190 19690 8210
rect 19710 8190 19715 8210
rect 19685 8180 19715 8190
rect 19745 8560 19775 8570
rect 19745 8540 19750 8560
rect 19770 8540 19775 8560
rect 19745 8510 19775 8540
rect 19745 8490 19750 8510
rect 19770 8490 19775 8510
rect 19745 8460 19775 8490
rect 19745 8440 19750 8460
rect 19770 8440 19775 8460
rect 19745 8410 19775 8440
rect 19745 8390 19750 8410
rect 19770 8390 19775 8410
rect 19745 8360 19775 8390
rect 19745 8340 19750 8360
rect 19770 8340 19775 8360
rect 19745 8310 19775 8340
rect 19745 8290 19750 8310
rect 19770 8290 19775 8310
rect 19745 8260 19775 8290
rect 19745 8240 19750 8260
rect 19770 8240 19775 8260
rect 19745 8210 19775 8240
rect 19745 8190 19750 8210
rect 19770 8190 19775 8210
rect 19745 8180 19775 8190
rect 19805 8560 19835 8570
rect 19805 8540 19810 8560
rect 19830 8540 19835 8560
rect 19805 8510 19835 8540
rect 19805 8490 19810 8510
rect 19830 8490 19835 8510
rect 19805 8460 19835 8490
rect 19805 8440 19810 8460
rect 19830 8440 19835 8460
rect 19805 8410 19835 8440
rect 19805 8390 19810 8410
rect 19830 8390 19835 8410
rect 19805 8360 19835 8390
rect 19805 8340 19810 8360
rect 19830 8340 19835 8360
rect 19805 8310 19835 8340
rect 19805 8290 19810 8310
rect 19830 8290 19835 8310
rect 19805 8260 19835 8290
rect 19805 8240 19810 8260
rect 19830 8240 19835 8260
rect 19805 8210 19835 8240
rect 19805 8190 19810 8210
rect 19830 8190 19835 8210
rect 19805 8180 19835 8190
rect 19865 8560 19895 8570
rect 19865 8540 19870 8560
rect 19890 8540 19895 8560
rect 19865 8510 19895 8540
rect 19865 8490 19870 8510
rect 19890 8490 19895 8510
rect 19865 8460 19895 8490
rect 19865 8440 19870 8460
rect 19890 8440 19895 8460
rect 19865 8410 19895 8440
rect 19865 8390 19870 8410
rect 19890 8390 19895 8410
rect 19865 8360 19895 8390
rect 19865 8340 19870 8360
rect 19890 8340 19895 8360
rect 19865 8310 19895 8340
rect 19865 8290 19870 8310
rect 19890 8290 19895 8310
rect 19865 8260 19895 8290
rect 19865 8240 19870 8260
rect 19890 8240 19895 8260
rect 19865 8210 19895 8240
rect 19865 8190 19870 8210
rect 19890 8190 19895 8210
rect 19865 8180 19895 8190
rect 19925 8560 19955 8570
rect 19925 8540 19930 8560
rect 19950 8540 19955 8560
rect 19925 8510 19955 8540
rect 19925 8490 19930 8510
rect 19950 8490 19955 8510
rect 19925 8460 19955 8490
rect 19925 8440 19930 8460
rect 19950 8440 19955 8460
rect 19925 8410 19955 8440
rect 19925 8390 19930 8410
rect 19950 8390 19955 8410
rect 19925 8360 19955 8390
rect 19925 8340 19930 8360
rect 19950 8340 19955 8360
rect 19925 8310 19955 8340
rect 19925 8290 19930 8310
rect 19950 8290 19955 8310
rect 19925 8260 19955 8290
rect 19925 8240 19930 8260
rect 19950 8240 19955 8260
rect 19925 8210 19955 8240
rect 19925 8190 19930 8210
rect 19950 8190 19955 8210
rect 19925 8180 19955 8190
rect 19985 8560 20015 8570
rect 19985 8540 19990 8560
rect 20010 8540 20015 8560
rect 19985 8510 20015 8540
rect 19985 8490 19990 8510
rect 20010 8490 20015 8510
rect 19985 8460 20015 8490
rect 19985 8440 19990 8460
rect 20010 8440 20015 8460
rect 19985 8410 20015 8440
rect 19985 8390 19990 8410
rect 20010 8390 20015 8410
rect 19985 8360 20015 8390
rect 19985 8340 19990 8360
rect 20010 8340 20015 8360
rect 19985 8310 20015 8340
rect 19985 8290 19990 8310
rect 20010 8290 20015 8310
rect 19985 8260 20015 8290
rect 19985 8240 19990 8260
rect 20010 8240 20015 8260
rect 19985 8210 20015 8240
rect 19985 8190 19990 8210
rect 20010 8190 20015 8210
rect 19985 8180 20015 8190
rect 20045 8560 20115 8570
rect 20045 8540 20050 8560
rect 20070 8540 20090 8560
rect 20110 8540 20115 8560
rect 20045 8510 20115 8540
rect 20045 8490 20050 8510
rect 20070 8490 20090 8510
rect 20110 8490 20115 8510
rect 20045 8460 20115 8490
rect 20045 8440 20050 8460
rect 20070 8440 20090 8460
rect 20110 8440 20115 8460
rect 20045 8410 20115 8440
rect 20045 8390 20050 8410
rect 20070 8390 20090 8410
rect 20110 8390 20115 8410
rect 20045 8360 20115 8390
rect 20045 8340 20050 8360
rect 20070 8340 20090 8360
rect 20110 8340 20115 8360
rect 20045 8310 20115 8340
rect 20045 8290 20050 8310
rect 20070 8290 20090 8310
rect 20110 8290 20115 8310
rect 20045 8260 20115 8290
rect 20045 8240 20050 8260
rect 20070 8240 20090 8260
rect 20110 8240 20115 8260
rect 20445 8285 20485 8295
rect 20445 8265 20455 8285
rect 20475 8265 20485 8285
rect 20445 8255 20485 8265
rect 20555 8285 20595 8295
rect 20555 8265 20565 8285
rect 20585 8265 20595 8285
rect 20555 8255 20595 8265
rect 20665 8285 20705 8295
rect 20665 8265 20675 8285
rect 20695 8265 20705 8285
rect 20665 8255 20705 8265
rect 20775 8285 20815 8295
rect 20775 8265 20785 8285
rect 20805 8265 20815 8285
rect 20775 8255 20815 8265
rect 20885 8285 20925 8295
rect 20885 8265 20895 8285
rect 20915 8265 20925 8285
rect 20885 8255 20925 8265
rect 20995 8285 21035 8295
rect 20995 8265 21005 8285
rect 21025 8265 21035 8285
rect 20995 8255 21035 8265
rect 21105 8285 21145 8295
rect 21105 8265 21115 8285
rect 21135 8265 21145 8285
rect 21105 8255 21145 8265
rect 21215 8285 21255 8295
rect 21215 8265 21225 8285
rect 21245 8265 21255 8285
rect 21215 8255 21255 8265
rect 21325 8285 21365 8295
rect 21325 8265 21335 8285
rect 21355 8265 21365 8285
rect 21325 8255 21365 8265
rect 21435 8285 21475 8295
rect 21435 8265 21445 8285
rect 21465 8265 21475 8285
rect 21435 8255 21475 8265
rect 21545 8285 21585 8295
rect 21545 8265 21555 8285
rect 21575 8265 21585 8285
rect 21545 8255 21585 8265
rect 20045 8210 20115 8240
rect 20455 8235 20475 8255
rect 20565 8235 20585 8255
rect 20675 8235 20695 8255
rect 20785 8235 20805 8255
rect 20895 8235 20915 8255
rect 21005 8235 21025 8255
rect 21115 8235 21135 8255
rect 21225 8235 21245 8255
rect 21335 8235 21355 8255
rect 21445 8235 21465 8255
rect 21555 8235 21575 8255
rect 20045 8190 20050 8210
rect 20070 8190 20090 8210
rect 20110 8190 20115 8210
rect 20045 8180 20115 8190
rect 20355 8225 20425 8235
rect 20355 8205 20360 8225
rect 20380 8205 20400 8225
rect 20420 8205 20425 8225
rect 14110 8155 14115 8175
rect 14135 8155 14155 8175
rect 14175 8155 14180 8175
rect 18790 8160 18810 8180
rect 18910 8160 18930 8180
rect 19030 8160 19050 8180
rect 19150 8160 19170 8180
rect 19270 8160 19290 8180
rect 19390 8160 19410 8180
rect 19510 8160 19530 8180
rect 19630 8160 19650 8180
rect 19750 8160 19770 8180
rect 19870 8160 19890 8180
rect 19990 8160 20010 8180
rect 20355 8175 20425 8205
rect 14110 8125 14180 8155
rect 14110 8105 14115 8125
rect 14135 8105 14155 8125
rect 14175 8105 14180 8125
rect 18780 8150 18820 8160
rect 18780 8130 18790 8150
rect 18810 8130 18820 8150
rect 18780 8120 18820 8130
rect 18900 8150 18940 8160
rect 18900 8130 18910 8150
rect 18930 8130 18940 8150
rect 18900 8120 18940 8130
rect 19020 8150 19060 8160
rect 19020 8130 19030 8150
rect 19050 8130 19060 8150
rect 19020 8120 19060 8130
rect 19140 8150 19180 8160
rect 19140 8130 19150 8150
rect 19170 8130 19180 8150
rect 19140 8120 19180 8130
rect 19260 8150 19300 8160
rect 19260 8130 19270 8150
rect 19290 8130 19300 8150
rect 19260 8120 19300 8130
rect 19323 8150 19357 8160
rect 19323 8130 19331 8150
rect 19349 8130 19357 8150
rect 19323 8120 19357 8130
rect 19380 8150 19420 8160
rect 19380 8130 19390 8150
rect 19410 8130 19420 8150
rect 19380 8120 19420 8130
rect 19500 8150 19540 8160
rect 19500 8130 19510 8150
rect 19530 8130 19540 8150
rect 19500 8120 19540 8130
rect 19620 8150 19660 8160
rect 19620 8130 19630 8150
rect 19650 8130 19660 8150
rect 19620 8120 19660 8130
rect 19740 8150 19780 8160
rect 19740 8130 19750 8150
rect 19770 8130 19780 8150
rect 19740 8120 19780 8130
rect 19860 8150 19900 8160
rect 19860 8130 19870 8150
rect 19890 8130 19900 8150
rect 19860 8120 19900 8130
rect 19980 8150 20020 8160
rect 19980 8130 19990 8150
rect 20010 8130 20020 8150
rect 19980 8120 20020 8130
rect 20355 8155 20360 8175
rect 20380 8155 20400 8175
rect 20420 8155 20425 8175
rect 20355 8125 20425 8155
rect 14110 8075 14180 8105
rect 14110 8055 14115 8075
rect 14135 8055 14155 8075
rect 14175 8055 14180 8075
rect 14110 8025 14180 8055
rect 14110 8005 14115 8025
rect 14135 8005 14155 8025
rect 14175 8005 14180 8025
rect 14110 7975 14180 8005
rect 14110 7955 14115 7975
rect 14135 7955 14155 7975
rect 14175 7955 14180 7975
rect 14110 7945 14180 7955
rect 20355 8105 20360 8125
rect 20380 8105 20400 8125
rect 20420 8105 20425 8125
rect 20355 8075 20425 8105
rect 20355 8055 20360 8075
rect 20380 8055 20400 8075
rect 20420 8055 20425 8075
rect 20355 8025 20425 8055
rect 20355 8005 20360 8025
rect 20380 8005 20400 8025
rect 20420 8005 20425 8025
rect 20355 7975 20425 8005
rect 20355 7955 20360 7975
rect 20380 7955 20400 7975
rect 20420 7955 20425 7975
rect 12580 7920 12590 7940
rect 12610 7920 12620 7940
rect 12865 7925 12885 7945
rect 13015 7925 13035 7945
rect 13125 7925 13145 7945
rect 13235 7925 13255 7945
rect 13345 7925 13365 7945
rect 13455 7925 13475 7945
rect 13565 7925 13585 7945
rect 13675 7925 13695 7945
rect 13785 7925 13805 7945
rect 13895 7925 13915 7945
rect 14005 7925 14025 7945
rect 14155 7925 14175 7945
rect 18680 7940 18720 7950
rect 12580 7910 12620 7920
rect 12855 7915 12895 7925
rect 11190 7890 11210 7910
rect 11350 7890 11370 7910
rect 11470 7890 11490 7910
rect 11590 7890 11610 7910
rect 11710 7890 11730 7910
rect 11830 7890 11850 7910
rect 11950 7890 11970 7910
rect 12070 7890 12090 7910
rect 12190 7890 12210 7910
rect 12310 7890 12330 7910
rect 12430 7890 12450 7910
rect 12590 7890 12610 7910
rect 12855 7895 12865 7915
rect 12885 7895 12895 7915
rect 11185 7880 11255 7890
rect 11185 7860 11190 7880
rect 11210 7860 11230 7880
rect 11250 7860 11255 7880
rect 11185 7830 11255 7860
rect 11185 7810 11190 7830
rect 11210 7810 11230 7830
rect 11250 7810 11255 7830
rect 11185 7780 11255 7810
rect 11185 7760 11190 7780
rect 11210 7760 11230 7780
rect 11250 7760 11255 7780
rect 11185 7730 11255 7760
rect 11185 7710 11190 7730
rect 11210 7710 11230 7730
rect 11250 7710 11255 7730
rect 11185 7680 11255 7710
rect 9735 7665 9775 7675
rect 9735 7645 9745 7665
rect 9765 7645 9775 7665
rect 9735 7635 9775 7645
rect 9845 7665 9885 7675
rect 9845 7645 9855 7665
rect 9875 7645 9885 7665
rect 9845 7635 9885 7645
rect 9955 7665 9995 7675
rect 9955 7645 9965 7665
rect 9985 7645 9995 7665
rect 9955 7635 9995 7645
rect 10065 7665 10105 7675
rect 10065 7645 10075 7665
rect 10095 7645 10105 7665
rect 10065 7635 10105 7645
rect 10175 7665 10215 7675
rect 10175 7645 10185 7665
rect 10205 7645 10215 7665
rect 10175 7635 10215 7645
rect 10285 7665 10325 7675
rect 10285 7645 10295 7665
rect 10315 7645 10325 7665
rect 10285 7635 10325 7645
rect 10395 7665 10435 7675
rect 10395 7645 10405 7665
rect 10425 7645 10435 7665
rect 10395 7635 10435 7645
rect 10505 7665 10545 7675
rect 10505 7645 10515 7665
rect 10535 7645 10545 7665
rect 10505 7635 10545 7645
rect 10615 7665 10655 7675
rect 10615 7645 10625 7665
rect 10645 7645 10655 7665
rect 10615 7635 10655 7645
rect 10725 7665 10765 7675
rect 10725 7645 10735 7665
rect 10755 7645 10765 7665
rect 10725 7635 10765 7645
rect 10835 7665 10875 7675
rect 10835 7645 10845 7665
rect 10865 7645 10875 7665
rect 10835 7635 10875 7645
rect 11185 7660 11190 7680
rect 11210 7660 11230 7680
rect 11250 7660 11255 7680
rect 9745 7615 9765 7635
rect 9855 7615 9875 7635
rect 9965 7615 9985 7635
rect 10075 7615 10095 7635
rect 10185 7615 10205 7635
rect 10295 7615 10315 7635
rect 10405 7615 10425 7635
rect 10515 7615 10535 7635
rect 10625 7615 10645 7635
rect 10735 7615 10755 7635
rect 10845 7615 10865 7635
rect 11185 7630 11255 7660
rect 9645 7605 9715 7615
rect 9645 7585 9650 7605
rect 9670 7585 9690 7605
rect 9710 7585 9715 7605
rect 9645 7555 9715 7585
rect 9645 7535 9650 7555
rect 9670 7535 9690 7555
rect 9710 7535 9715 7555
rect 9645 7525 9715 7535
rect 9740 7605 9770 7615
rect 9740 7585 9745 7605
rect 9765 7585 9770 7605
rect 9740 7555 9770 7585
rect 9740 7535 9745 7555
rect 9765 7535 9770 7555
rect 9740 7525 9770 7535
rect 9795 7605 9825 7615
rect 9795 7585 9800 7605
rect 9820 7585 9825 7605
rect 9795 7555 9825 7585
rect 9795 7535 9800 7555
rect 9820 7535 9825 7555
rect 9795 7525 9825 7535
rect 9850 7605 9880 7615
rect 9850 7585 9855 7605
rect 9875 7585 9880 7605
rect 9850 7555 9880 7585
rect 9850 7535 9855 7555
rect 9875 7535 9880 7555
rect 9850 7525 9880 7535
rect 9905 7605 9935 7615
rect 9905 7585 9910 7605
rect 9930 7585 9935 7605
rect 9905 7555 9935 7585
rect 9905 7535 9910 7555
rect 9930 7535 9935 7555
rect 9905 7525 9935 7535
rect 9960 7605 9990 7615
rect 9960 7585 9965 7605
rect 9985 7585 9990 7605
rect 9960 7555 9990 7585
rect 9960 7535 9965 7555
rect 9985 7535 9990 7555
rect 9960 7525 9990 7535
rect 10015 7605 10045 7615
rect 10015 7585 10020 7605
rect 10040 7585 10045 7605
rect 10015 7555 10045 7585
rect 10015 7535 10020 7555
rect 10040 7535 10045 7555
rect 10015 7525 10045 7535
rect 10070 7605 10100 7615
rect 10070 7585 10075 7605
rect 10095 7585 10100 7605
rect 10070 7555 10100 7585
rect 10070 7535 10075 7555
rect 10095 7535 10100 7555
rect 10070 7525 10100 7535
rect 10125 7605 10155 7615
rect 10125 7585 10130 7605
rect 10150 7585 10155 7605
rect 10125 7555 10155 7585
rect 10125 7535 10130 7555
rect 10150 7535 10155 7555
rect 10125 7525 10155 7535
rect 10180 7605 10210 7615
rect 10180 7585 10185 7605
rect 10205 7585 10210 7605
rect 10180 7555 10210 7585
rect 10180 7535 10185 7555
rect 10205 7535 10210 7555
rect 10180 7525 10210 7535
rect 10235 7605 10265 7615
rect 10235 7585 10240 7605
rect 10260 7585 10265 7605
rect 10235 7555 10265 7585
rect 10235 7535 10240 7555
rect 10260 7535 10265 7555
rect 10235 7525 10265 7535
rect 10290 7605 10320 7615
rect 10290 7585 10295 7605
rect 10315 7585 10320 7605
rect 10290 7555 10320 7585
rect 10290 7535 10295 7555
rect 10315 7535 10320 7555
rect 10290 7525 10320 7535
rect 10345 7605 10375 7615
rect 10345 7585 10350 7605
rect 10370 7585 10375 7605
rect 10345 7555 10375 7585
rect 10345 7535 10350 7555
rect 10370 7535 10375 7555
rect 10345 7525 10375 7535
rect 10400 7605 10430 7615
rect 10400 7585 10405 7605
rect 10425 7585 10430 7605
rect 10400 7555 10430 7585
rect 10400 7535 10405 7555
rect 10425 7535 10430 7555
rect 10400 7525 10430 7535
rect 10455 7605 10485 7615
rect 10455 7585 10460 7605
rect 10480 7585 10485 7605
rect 10455 7555 10485 7585
rect 10455 7535 10460 7555
rect 10480 7535 10485 7555
rect 10455 7525 10485 7535
rect 10510 7605 10540 7615
rect 10510 7585 10515 7605
rect 10535 7585 10540 7605
rect 10510 7555 10540 7585
rect 10510 7535 10515 7555
rect 10535 7535 10540 7555
rect 10510 7525 10540 7535
rect 10565 7605 10595 7615
rect 10565 7585 10570 7605
rect 10590 7585 10595 7605
rect 10565 7555 10595 7585
rect 10565 7535 10570 7555
rect 10590 7535 10595 7555
rect 10565 7525 10595 7535
rect 10620 7605 10650 7615
rect 10620 7585 10625 7605
rect 10645 7585 10650 7605
rect 10620 7555 10650 7585
rect 10620 7535 10625 7555
rect 10645 7535 10650 7555
rect 10620 7525 10650 7535
rect 10675 7605 10705 7615
rect 10675 7585 10680 7605
rect 10700 7585 10705 7605
rect 10675 7555 10705 7585
rect 10675 7535 10680 7555
rect 10700 7535 10705 7555
rect 10675 7525 10705 7535
rect 10730 7605 10760 7615
rect 10730 7585 10735 7605
rect 10755 7585 10760 7605
rect 10730 7555 10760 7585
rect 10730 7535 10735 7555
rect 10755 7535 10760 7555
rect 10730 7525 10760 7535
rect 10785 7605 10815 7615
rect 10785 7585 10790 7605
rect 10810 7585 10815 7605
rect 10785 7555 10815 7585
rect 10785 7535 10790 7555
rect 10810 7535 10815 7555
rect 10785 7525 10815 7535
rect 10840 7605 10870 7615
rect 10840 7585 10845 7605
rect 10865 7585 10870 7605
rect 10840 7555 10870 7585
rect 10840 7535 10845 7555
rect 10865 7535 10870 7555
rect 10840 7525 10870 7535
rect 10895 7605 10965 7615
rect 10895 7585 10900 7605
rect 10920 7585 10940 7605
rect 10960 7585 10965 7605
rect 10895 7555 10965 7585
rect 10895 7535 10900 7555
rect 10920 7535 10940 7555
rect 10960 7535 10965 7555
rect 10895 7525 10965 7535
rect 11185 7610 11190 7630
rect 11210 7610 11230 7630
rect 11250 7610 11255 7630
rect 11185 7580 11255 7610
rect 11185 7560 11190 7580
rect 11210 7560 11230 7580
rect 11250 7560 11255 7580
rect 11185 7530 11255 7560
rect 9650 7505 9670 7525
rect 9800 7505 9820 7525
rect 9910 7505 9930 7525
rect 10020 7505 10040 7525
rect 10130 7505 10150 7525
rect 10240 7505 10260 7525
rect 10350 7505 10370 7525
rect 10460 7505 10480 7525
rect 10570 7505 10590 7525
rect 10680 7505 10700 7525
rect 10790 7505 10810 7525
rect 10940 7505 10960 7525
rect 11185 7510 11190 7530
rect 11210 7510 11230 7530
rect 11250 7510 11255 7530
rect 9640 7495 9680 7505
rect 9640 7475 9650 7495
rect 9670 7475 9680 7495
rect 9640 7465 9680 7475
rect 9790 7495 9830 7505
rect 9790 7475 9800 7495
rect 9820 7475 9830 7495
rect 9790 7465 9830 7475
rect 9900 7495 9940 7505
rect 9900 7475 9910 7495
rect 9930 7475 9940 7495
rect 9900 7465 9940 7475
rect 10010 7495 10050 7505
rect 10010 7475 10020 7495
rect 10040 7475 10050 7495
rect 10010 7465 10050 7475
rect 10120 7495 10160 7505
rect 10120 7475 10130 7495
rect 10150 7475 10160 7495
rect 10120 7465 10160 7475
rect 10230 7495 10270 7505
rect 10230 7475 10240 7495
rect 10260 7475 10270 7495
rect 10230 7465 10270 7475
rect 10340 7495 10380 7505
rect 10340 7475 10350 7495
rect 10370 7475 10380 7495
rect 10340 7465 10380 7475
rect 10450 7495 10490 7505
rect 10450 7475 10460 7495
rect 10480 7475 10490 7495
rect 10450 7465 10490 7475
rect 10560 7495 10600 7505
rect 10560 7475 10570 7495
rect 10590 7475 10600 7495
rect 10560 7465 10600 7475
rect 10670 7495 10710 7505
rect 10670 7475 10680 7495
rect 10700 7475 10710 7495
rect 10670 7465 10710 7475
rect 10780 7495 10820 7505
rect 10780 7475 10790 7495
rect 10810 7475 10820 7495
rect 10780 7465 10820 7475
rect 10930 7495 10970 7505
rect 11185 7500 11255 7510
rect 11285 7880 11315 7890
rect 11285 7860 11290 7880
rect 11310 7860 11315 7880
rect 11285 7830 11315 7860
rect 11285 7810 11290 7830
rect 11310 7810 11315 7830
rect 11285 7780 11315 7810
rect 11285 7760 11290 7780
rect 11310 7760 11315 7780
rect 11285 7730 11315 7760
rect 11285 7710 11290 7730
rect 11310 7710 11315 7730
rect 11285 7680 11315 7710
rect 11285 7660 11290 7680
rect 11310 7660 11315 7680
rect 11285 7630 11315 7660
rect 11285 7610 11290 7630
rect 11310 7610 11315 7630
rect 11285 7580 11315 7610
rect 11285 7560 11290 7580
rect 11310 7560 11315 7580
rect 11285 7530 11315 7560
rect 11285 7510 11290 7530
rect 11310 7510 11315 7530
rect 11285 7500 11315 7510
rect 11345 7880 11375 7890
rect 11345 7860 11350 7880
rect 11370 7860 11375 7880
rect 11345 7830 11375 7860
rect 11345 7810 11350 7830
rect 11370 7810 11375 7830
rect 11345 7780 11375 7810
rect 11345 7760 11350 7780
rect 11370 7760 11375 7780
rect 11345 7730 11375 7760
rect 11345 7710 11350 7730
rect 11370 7710 11375 7730
rect 11345 7680 11375 7710
rect 11345 7660 11350 7680
rect 11370 7660 11375 7680
rect 11345 7630 11375 7660
rect 11345 7610 11350 7630
rect 11370 7610 11375 7630
rect 11345 7580 11375 7610
rect 11345 7560 11350 7580
rect 11370 7560 11375 7580
rect 11345 7530 11375 7560
rect 11345 7510 11350 7530
rect 11370 7510 11375 7530
rect 11345 7500 11375 7510
rect 11405 7880 11435 7890
rect 11405 7860 11410 7880
rect 11430 7860 11435 7880
rect 11405 7830 11435 7860
rect 11405 7810 11410 7830
rect 11430 7810 11435 7830
rect 11405 7780 11435 7810
rect 11405 7760 11410 7780
rect 11430 7760 11435 7780
rect 11405 7730 11435 7760
rect 11405 7710 11410 7730
rect 11430 7710 11435 7730
rect 11405 7680 11435 7710
rect 11405 7660 11410 7680
rect 11430 7660 11435 7680
rect 11405 7630 11435 7660
rect 11405 7610 11410 7630
rect 11430 7610 11435 7630
rect 11405 7580 11435 7610
rect 11405 7560 11410 7580
rect 11430 7560 11435 7580
rect 11405 7530 11435 7560
rect 11405 7510 11410 7530
rect 11430 7510 11435 7530
rect 11405 7500 11435 7510
rect 11465 7880 11495 7890
rect 11465 7860 11470 7880
rect 11490 7860 11495 7880
rect 11465 7830 11495 7860
rect 11465 7810 11470 7830
rect 11490 7810 11495 7830
rect 11465 7780 11495 7810
rect 11465 7760 11470 7780
rect 11490 7760 11495 7780
rect 11465 7730 11495 7760
rect 11465 7710 11470 7730
rect 11490 7710 11495 7730
rect 11465 7680 11495 7710
rect 11465 7660 11470 7680
rect 11490 7660 11495 7680
rect 11465 7630 11495 7660
rect 11465 7610 11470 7630
rect 11490 7610 11495 7630
rect 11465 7580 11495 7610
rect 11465 7560 11470 7580
rect 11490 7560 11495 7580
rect 11465 7530 11495 7560
rect 11465 7510 11470 7530
rect 11490 7510 11495 7530
rect 11465 7500 11495 7510
rect 11525 7880 11555 7890
rect 11525 7860 11530 7880
rect 11550 7860 11555 7880
rect 11525 7830 11555 7860
rect 11525 7810 11530 7830
rect 11550 7810 11555 7830
rect 11525 7780 11555 7810
rect 11525 7760 11530 7780
rect 11550 7760 11555 7780
rect 11525 7730 11555 7760
rect 11525 7710 11530 7730
rect 11550 7710 11555 7730
rect 11525 7680 11555 7710
rect 11525 7660 11530 7680
rect 11550 7660 11555 7680
rect 11525 7630 11555 7660
rect 11525 7610 11530 7630
rect 11550 7610 11555 7630
rect 11525 7580 11555 7610
rect 11525 7560 11530 7580
rect 11550 7560 11555 7580
rect 11525 7530 11555 7560
rect 11525 7510 11530 7530
rect 11550 7510 11555 7530
rect 11525 7500 11555 7510
rect 11585 7880 11615 7890
rect 11585 7860 11590 7880
rect 11610 7860 11615 7880
rect 11585 7830 11615 7860
rect 11585 7810 11590 7830
rect 11610 7810 11615 7830
rect 11585 7780 11615 7810
rect 11585 7760 11590 7780
rect 11610 7760 11615 7780
rect 11585 7730 11615 7760
rect 11585 7710 11590 7730
rect 11610 7710 11615 7730
rect 11585 7680 11615 7710
rect 11585 7660 11590 7680
rect 11610 7660 11615 7680
rect 11585 7630 11615 7660
rect 11585 7610 11590 7630
rect 11610 7610 11615 7630
rect 11585 7580 11615 7610
rect 11585 7560 11590 7580
rect 11610 7560 11615 7580
rect 11585 7530 11615 7560
rect 11585 7510 11590 7530
rect 11610 7510 11615 7530
rect 11585 7500 11615 7510
rect 11645 7880 11675 7890
rect 11645 7860 11650 7880
rect 11670 7860 11675 7880
rect 11645 7830 11675 7860
rect 11645 7810 11650 7830
rect 11670 7810 11675 7830
rect 11645 7780 11675 7810
rect 11645 7760 11650 7780
rect 11670 7760 11675 7780
rect 11645 7730 11675 7760
rect 11645 7710 11650 7730
rect 11670 7710 11675 7730
rect 11645 7680 11675 7710
rect 11645 7660 11650 7680
rect 11670 7660 11675 7680
rect 11645 7630 11675 7660
rect 11645 7610 11650 7630
rect 11670 7610 11675 7630
rect 11645 7580 11675 7610
rect 11645 7560 11650 7580
rect 11670 7560 11675 7580
rect 11645 7530 11675 7560
rect 11645 7510 11650 7530
rect 11670 7510 11675 7530
rect 11645 7500 11675 7510
rect 11705 7880 11735 7890
rect 11705 7860 11710 7880
rect 11730 7860 11735 7880
rect 11705 7830 11735 7860
rect 11705 7810 11710 7830
rect 11730 7810 11735 7830
rect 11705 7780 11735 7810
rect 11705 7760 11710 7780
rect 11730 7760 11735 7780
rect 11705 7730 11735 7760
rect 11705 7710 11710 7730
rect 11730 7710 11735 7730
rect 11705 7680 11735 7710
rect 11705 7660 11710 7680
rect 11730 7660 11735 7680
rect 11705 7630 11735 7660
rect 11705 7610 11710 7630
rect 11730 7610 11735 7630
rect 11705 7580 11735 7610
rect 11705 7560 11710 7580
rect 11730 7560 11735 7580
rect 11705 7530 11735 7560
rect 11705 7510 11710 7530
rect 11730 7510 11735 7530
rect 11705 7500 11735 7510
rect 11765 7880 11795 7890
rect 11765 7860 11770 7880
rect 11790 7860 11795 7880
rect 11765 7830 11795 7860
rect 11765 7810 11770 7830
rect 11790 7810 11795 7830
rect 11765 7780 11795 7810
rect 11765 7760 11770 7780
rect 11790 7760 11795 7780
rect 11765 7730 11795 7760
rect 11765 7710 11770 7730
rect 11790 7710 11795 7730
rect 11765 7680 11795 7710
rect 11765 7660 11770 7680
rect 11790 7660 11795 7680
rect 11765 7630 11795 7660
rect 11765 7610 11770 7630
rect 11790 7610 11795 7630
rect 11765 7580 11795 7610
rect 11765 7560 11770 7580
rect 11790 7560 11795 7580
rect 11765 7530 11795 7560
rect 11765 7510 11770 7530
rect 11790 7510 11795 7530
rect 11765 7500 11795 7510
rect 11825 7880 11855 7890
rect 11825 7860 11830 7880
rect 11850 7860 11855 7880
rect 11825 7830 11855 7860
rect 11825 7810 11830 7830
rect 11850 7810 11855 7830
rect 11825 7780 11855 7810
rect 11825 7760 11830 7780
rect 11850 7760 11855 7780
rect 11825 7730 11855 7760
rect 11825 7710 11830 7730
rect 11850 7710 11855 7730
rect 11825 7680 11855 7710
rect 11825 7660 11830 7680
rect 11850 7660 11855 7680
rect 11825 7630 11855 7660
rect 11825 7610 11830 7630
rect 11850 7610 11855 7630
rect 11825 7580 11855 7610
rect 11825 7560 11830 7580
rect 11850 7560 11855 7580
rect 11825 7530 11855 7560
rect 11825 7510 11830 7530
rect 11850 7510 11855 7530
rect 11825 7500 11855 7510
rect 11885 7880 11915 7890
rect 11885 7860 11890 7880
rect 11910 7860 11915 7880
rect 11885 7830 11915 7860
rect 11885 7810 11890 7830
rect 11910 7810 11915 7830
rect 11885 7780 11915 7810
rect 11885 7760 11890 7780
rect 11910 7760 11915 7780
rect 11885 7730 11915 7760
rect 11885 7710 11890 7730
rect 11910 7710 11915 7730
rect 11885 7680 11915 7710
rect 11885 7660 11890 7680
rect 11910 7660 11915 7680
rect 11885 7630 11915 7660
rect 11885 7610 11890 7630
rect 11910 7610 11915 7630
rect 11885 7580 11915 7610
rect 11885 7560 11890 7580
rect 11910 7560 11915 7580
rect 11885 7530 11915 7560
rect 11885 7510 11890 7530
rect 11910 7510 11915 7530
rect 11885 7500 11915 7510
rect 11945 7880 11975 7890
rect 11945 7860 11950 7880
rect 11970 7860 11975 7880
rect 11945 7830 11975 7860
rect 11945 7810 11950 7830
rect 11970 7810 11975 7830
rect 11945 7780 11975 7810
rect 11945 7760 11950 7780
rect 11970 7760 11975 7780
rect 11945 7730 11975 7760
rect 11945 7710 11950 7730
rect 11970 7710 11975 7730
rect 11945 7680 11975 7710
rect 11945 7660 11950 7680
rect 11970 7660 11975 7680
rect 11945 7630 11975 7660
rect 11945 7610 11950 7630
rect 11970 7610 11975 7630
rect 11945 7580 11975 7610
rect 11945 7560 11950 7580
rect 11970 7560 11975 7580
rect 11945 7530 11975 7560
rect 11945 7510 11950 7530
rect 11970 7510 11975 7530
rect 11945 7500 11975 7510
rect 12005 7880 12035 7890
rect 12005 7860 12010 7880
rect 12030 7860 12035 7880
rect 12005 7830 12035 7860
rect 12005 7810 12010 7830
rect 12030 7810 12035 7830
rect 12005 7780 12035 7810
rect 12005 7760 12010 7780
rect 12030 7760 12035 7780
rect 12005 7730 12035 7760
rect 12005 7710 12010 7730
rect 12030 7710 12035 7730
rect 12005 7680 12035 7710
rect 12005 7660 12010 7680
rect 12030 7660 12035 7680
rect 12005 7630 12035 7660
rect 12005 7610 12010 7630
rect 12030 7610 12035 7630
rect 12005 7580 12035 7610
rect 12005 7560 12010 7580
rect 12030 7560 12035 7580
rect 12005 7530 12035 7560
rect 12005 7510 12010 7530
rect 12030 7510 12035 7530
rect 12005 7500 12035 7510
rect 12065 7880 12095 7890
rect 12065 7860 12070 7880
rect 12090 7860 12095 7880
rect 12065 7830 12095 7860
rect 12065 7810 12070 7830
rect 12090 7810 12095 7830
rect 12065 7780 12095 7810
rect 12065 7760 12070 7780
rect 12090 7760 12095 7780
rect 12065 7730 12095 7760
rect 12065 7710 12070 7730
rect 12090 7710 12095 7730
rect 12065 7680 12095 7710
rect 12065 7660 12070 7680
rect 12090 7660 12095 7680
rect 12065 7630 12095 7660
rect 12065 7610 12070 7630
rect 12090 7610 12095 7630
rect 12065 7580 12095 7610
rect 12065 7560 12070 7580
rect 12090 7560 12095 7580
rect 12065 7530 12095 7560
rect 12065 7510 12070 7530
rect 12090 7510 12095 7530
rect 12065 7500 12095 7510
rect 12125 7880 12155 7890
rect 12125 7860 12130 7880
rect 12150 7860 12155 7880
rect 12125 7830 12155 7860
rect 12125 7810 12130 7830
rect 12150 7810 12155 7830
rect 12125 7780 12155 7810
rect 12125 7760 12130 7780
rect 12150 7760 12155 7780
rect 12125 7730 12155 7760
rect 12125 7710 12130 7730
rect 12150 7710 12155 7730
rect 12125 7680 12155 7710
rect 12125 7660 12130 7680
rect 12150 7660 12155 7680
rect 12125 7630 12155 7660
rect 12125 7610 12130 7630
rect 12150 7610 12155 7630
rect 12125 7580 12155 7610
rect 12125 7560 12130 7580
rect 12150 7560 12155 7580
rect 12125 7530 12155 7560
rect 12125 7510 12130 7530
rect 12150 7510 12155 7530
rect 12125 7500 12155 7510
rect 12185 7880 12215 7890
rect 12185 7860 12190 7880
rect 12210 7860 12215 7880
rect 12185 7830 12215 7860
rect 12185 7810 12190 7830
rect 12210 7810 12215 7830
rect 12185 7780 12215 7810
rect 12185 7760 12190 7780
rect 12210 7760 12215 7780
rect 12185 7730 12215 7760
rect 12185 7710 12190 7730
rect 12210 7710 12215 7730
rect 12185 7680 12215 7710
rect 12185 7660 12190 7680
rect 12210 7660 12215 7680
rect 12185 7630 12215 7660
rect 12185 7610 12190 7630
rect 12210 7610 12215 7630
rect 12185 7580 12215 7610
rect 12185 7560 12190 7580
rect 12210 7560 12215 7580
rect 12185 7530 12215 7560
rect 12185 7510 12190 7530
rect 12210 7510 12215 7530
rect 12185 7500 12215 7510
rect 12245 7880 12275 7890
rect 12245 7860 12250 7880
rect 12270 7860 12275 7880
rect 12245 7830 12275 7860
rect 12245 7810 12250 7830
rect 12270 7810 12275 7830
rect 12245 7780 12275 7810
rect 12245 7760 12250 7780
rect 12270 7760 12275 7780
rect 12245 7730 12275 7760
rect 12245 7710 12250 7730
rect 12270 7710 12275 7730
rect 12245 7680 12275 7710
rect 12245 7660 12250 7680
rect 12270 7660 12275 7680
rect 12245 7630 12275 7660
rect 12245 7610 12250 7630
rect 12270 7610 12275 7630
rect 12245 7580 12275 7610
rect 12245 7560 12250 7580
rect 12270 7560 12275 7580
rect 12245 7530 12275 7560
rect 12245 7510 12250 7530
rect 12270 7510 12275 7530
rect 12245 7500 12275 7510
rect 12305 7880 12335 7890
rect 12305 7860 12310 7880
rect 12330 7860 12335 7880
rect 12305 7830 12335 7860
rect 12305 7810 12310 7830
rect 12330 7810 12335 7830
rect 12305 7780 12335 7810
rect 12305 7760 12310 7780
rect 12330 7760 12335 7780
rect 12305 7730 12335 7760
rect 12305 7710 12310 7730
rect 12330 7710 12335 7730
rect 12305 7680 12335 7710
rect 12305 7660 12310 7680
rect 12330 7660 12335 7680
rect 12305 7630 12335 7660
rect 12305 7610 12310 7630
rect 12330 7610 12335 7630
rect 12305 7580 12335 7610
rect 12305 7560 12310 7580
rect 12330 7560 12335 7580
rect 12305 7530 12335 7560
rect 12305 7510 12310 7530
rect 12330 7510 12335 7530
rect 12305 7500 12335 7510
rect 12365 7880 12395 7890
rect 12365 7860 12370 7880
rect 12390 7860 12395 7880
rect 12365 7830 12395 7860
rect 12365 7810 12370 7830
rect 12390 7810 12395 7830
rect 12365 7780 12395 7810
rect 12365 7760 12370 7780
rect 12390 7760 12395 7780
rect 12365 7730 12395 7760
rect 12365 7710 12370 7730
rect 12390 7710 12395 7730
rect 12365 7680 12395 7710
rect 12365 7660 12370 7680
rect 12390 7660 12395 7680
rect 12365 7630 12395 7660
rect 12365 7610 12370 7630
rect 12390 7610 12395 7630
rect 12365 7580 12395 7610
rect 12365 7560 12370 7580
rect 12390 7560 12395 7580
rect 12365 7530 12395 7560
rect 12365 7510 12370 7530
rect 12390 7510 12395 7530
rect 12365 7500 12395 7510
rect 12425 7880 12455 7890
rect 12425 7860 12430 7880
rect 12450 7860 12455 7880
rect 12425 7830 12455 7860
rect 12425 7810 12430 7830
rect 12450 7810 12455 7830
rect 12425 7780 12455 7810
rect 12425 7760 12430 7780
rect 12450 7760 12455 7780
rect 12425 7730 12455 7760
rect 12425 7710 12430 7730
rect 12450 7710 12455 7730
rect 12425 7680 12455 7710
rect 12425 7660 12430 7680
rect 12450 7660 12455 7680
rect 12425 7630 12455 7660
rect 12425 7610 12430 7630
rect 12450 7610 12455 7630
rect 12425 7580 12455 7610
rect 12425 7560 12430 7580
rect 12450 7560 12455 7580
rect 12425 7530 12455 7560
rect 12425 7510 12430 7530
rect 12450 7510 12455 7530
rect 12425 7500 12455 7510
rect 12485 7880 12515 7890
rect 12485 7860 12490 7880
rect 12510 7860 12515 7880
rect 12485 7830 12515 7860
rect 12485 7810 12490 7830
rect 12510 7810 12515 7830
rect 12485 7780 12515 7810
rect 12485 7760 12490 7780
rect 12510 7760 12515 7780
rect 12485 7730 12515 7760
rect 12485 7710 12490 7730
rect 12510 7710 12515 7730
rect 12485 7680 12515 7710
rect 12485 7660 12490 7680
rect 12510 7660 12515 7680
rect 12485 7630 12515 7660
rect 12485 7610 12490 7630
rect 12510 7610 12515 7630
rect 12485 7580 12515 7610
rect 12485 7560 12490 7580
rect 12510 7560 12515 7580
rect 12485 7530 12515 7560
rect 12485 7510 12490 7530
rect 12510 7510 12515 7530
rect 12485 7500 12515 7510
rect 12545 7880 12615 7890
rect 12855 7885 12895 7895
rect 13005 7915 13045 7925
rect 13005 7895 13015 7915
rect 13035 7895 13045 7915
rect 13005 7885 13045 7895
rect 13063 7915 13097 7925
rect 13063 7895 13071 7915
rect 13089 7895 13097 7915
rect 13063 7885 13097 7895
rect 13115 7915 13155 7925
rect 13115 7895 13125 7915
rect 13145 7895 13155 7915
rect 13115 7885 13155 7895
rect 13225 7915 13265 7925
rect 13225 7895 13235 7915
rect 13255 7895 13265 7915
rect 13225 7885 13265 7895
rect 13335 7915 13375 7925
rect 13335 7895 13345 7915
rect 13365 7895 13375 7915
rect 13335 7885 13375 7895
rect 13445 7915 13485 7925
rect 13445 7895 13455 7915
rect 13475 7895 13485 7915
rect 13445 7885 13485 7895
rect 13555 7915 13595 7925
rect 13555 7895 13565 7915
rect 13585 7895 13595 7915
rect 13555 7885 13595 7895
rect 13665 7915 13705 7925
rect 13665 7895 13675 7915
rect 13695 7895 13705 7915
rect 13665 7885 13705 7895
rect 13775 7915 13815 7925
rect 13775 7895 13785 7915
rect 13805 7895 13815 7915
rect 13775 7885 13815 7895
rect 13885 7915 13925 7925
rect 13885 7895 13895 7915
rect 13915 7895 13925 7915
rect 13885 7885 13925 7895
rect 13995 7915 14035 7925
rect 13995 7895 14005 7915
rect 14025 7895 14035 7915
rect 13995 7885 14035 7895
rect 14145 7915 14185 7925
rect 14145 7895 14155 7915
rect 14175 7895 14185 7915
rect 18680 7920 18690 7940
rect 18710 7920 18720 7940
rect 18680 7910 18720 7920
rect 18840 7940 18880 7950
rect 18840 7920 18850 7940
rect 18870 7920 18880 7940
rect 18840 7910 18880 7920
rect 18960 7940 19000 7950
rect 18960 7920 18970 7940
rect 18990 7920 19000 7940
rect 18960 7910 19000 7920
rect 19080 7940 19120 7950
rect 19080 7920 19090 7940
rect 19110 7920 19120 7940
rect 19080 7910 19120 7920
rect 19200 7940 19240 7950
rect 19200 7920 19210 7940
rect 19230 7920 19240 7940
rect 19200 7910 19240 7920
rect 19320 7940 19360 7950
rect 19320 7920 19330 7940
rect 19350 7920 19360 7940
rect 19320 7910 19360 7920
rect 19440 7940 19480 7950
rect 19440 7920 19450 7940
rect 19470 7920 19480 7940
rect 19440 7910 19480 7920
rect 19560 7940 19600 7950
rect 19560 7920 19570 7940
rect 19590 7920 19600 7940
rect 19560 7910 19600 7920
rect 19680 7940 19720 7950
rect 19680 7920 19690 7940
rect 19710 7920 19720 7940
rect 19680 7910 19720 7920
rect 19800 7940 19840 7950
rect 19800 7920 19810 7940
rect 19830 7920 19840 7940
rect 19800 7910 19840 7920
rect 19920 7940 19960 7950
rect 19920 7920 19930 7940
rect 19950 7920 19960 7940
rect 19920 7910 19960 7920
rect 19980 7910 20020 7950
rect 20080 7940 20120 7950
rect 20355 7945 20425 7955
rect 20450 8225 20480 8235
rect 20450 8205 20455 8225
rect 20475 8205 20480 8225
rect 20450 8175 20480 8205
rect 20450 8155 20455 8175
rect 20475 8155 20480 8175
rect 20450 8125 20480 8155
rect 20450 8105 20455 8125
rect 20475 8105 20480 8125
rect 20450 8075 20480 8105
rect 20450 8055 20455 8075
rect 20475 8055 20480 8075
rect 20450 8025 20480 8055
rect 20450 8005 20455 8025
rect 20475 8005 20480 8025
rect 20450 7975 20480 8005
rect 20450 7955 20455 7975
rect 20475 7955 20480 7975
rect 20450 7945 20480 7955
rect 20505 8225 20535 8235
rect 20505 8205 20510 8225
rect 20530 8205 20535 8225
rect 20505 8175 20535 8205
rect 20505 8155 20510 8175
rect 20530 8155 20535 8175
rect 20505 8125 20535 8155
rect 20505 8105 20510 8125
rect 20530 8105 20535 8125
rect 20505 8075 20535 8105
rect 20505 8055 20510 8075
rect 20530 8055 20535 8075
rect 20505 8025 20535 8055
rect 20505 8005 20510 8025
rect 20530 8005 20535 8025
rect 20505 7975 20535 8005
rect 20505 7955 20510 7975
rect 20530 7955 20535 7975
rect 20505 7945 20535 7955
rect 20560 8225 20590 8235
rect 20560 8205 20565 8225
rect 20585 8205 20590 8225
rect 20560 8175 20590 8205
rect 20560 8155 20565 8175
rect 20585 8155 20590 8175
rect 20560 8125 20590 8155
rect 20560 8105 20565 8125
rect 20585 8105 20590 8125
rect 20560 8075 20590 8105
rect 20560 8055 20565 8075
rect 20585 8055 20590 8075
rect 20560 8025 20590 8055
rect 20560 8005 20565 8025
rect 20585 8005 20590 8025
rect 20560 7975 20590 8005
rect 20560 7955 20565 7975
rect 20585 7955 20590 7975
rect 20560 7945 20590 7955
rect 20615 8225 20645 8235
rect 20615 8205 20620 8225
rect 20640 8205 20645 8225
rect 20615 8175 20645 8205
rect 20615 8155 20620 8175
rect 20640 8155 20645 8175
rect 20615 8125 20645 8155
rect 20615 8105 20620 8125
rect 20640 8105 20645 8125
rect 20615 8075 20645 8105
rect 20615 8055 20620 8075
rect 20640 8055 20645 8075
rect 20615 8025 20645 8055
rect 20615 8005 20620 8025
rect 20640 8005 20645 8025
rect 20615 7975 20645 8005
rect 20615 7955 20620 7975
rect 20640 7955 20645 7975
rect 20615 7945 20645 7955
rect 20670 8225 20700 8235
rect 20670 8205 20675 8225
rect 20695 8205 20700 8225
rect 20670 8175 20700 8205
rect 20670 8155 20675 8175
rect 20695 8155 20700 8175
rect 20670 8125 20700 8155
rect 20670 8105 20675 8125
rect 20695 8105 20700 8125
rect 20670 8075 20700 8105
rect 20670 8055 20675 8075
rect 20695 8055 20700 8075
rect 20670 8025 20700 8055
rect 20670 8005 20675 8025
rect 20695 8005 20700 8025
rect 20670 7975 20700 8005
rect 20670 7955 20675 7975
rect 20695 7955 20700 7975
rect 20670 7945 20700 7955
rect 20725 8225 20755 8235
rect 20725 8205 20730 8225
rect 20750 8205 20755 8225
rect 20725 8175 20755 8205
rect 20725 8155 20730 8175
rect 20750 8155 20755 8175
rect 20725 8125 20755 8155
rect 20725 8105 20730 8125
rect 20750 8105 20755 8125
rect 20725 8075 20755 8105
rect 20725 8055 20730 8075
rect 20750 8055 20755 8075
rect 20725 8025 20755 8055
rect 20725 8005 20730 8025
rect 20750 8005 20755 8025
rect 20725 7975 20755 8005
rect 20725 7955 20730 7975
rect 20750 7955 20755 7975
rect 20725 7945 20755 7955
rect 20780 8225 20810 8235
rect 20780 8205 20785 8225
rect 20805 8205 20810 8225
rect 20780 8175 20810 8205
rect 20780 8155 20785 8175
rect 20805 8155 20810 8175
rect 20780 8125 20810 8155
rect 20780 8105 20785 8125
rect 20805 8105 20810 8125
rect 20780 8075 20810 8105
rect 20780 8055 20785 8075
rect 20805 8055 20810 8075
rect 20780 8025 20810 8055
rect 20780 8005 20785 8025
rect 20805 8005 20810 8025
rect 20780 7975 20810 8005
rect 20780 7955 20785 7975
rect 20805 7955 20810 7975
rect 20780 7945 20810 7955
rect 20835 8225 20865 8235
rect 20835 8205 20840 8225
rect 20860 8205 20865 8225
rect 20835 8175 20865 8205
rect 20835 8155 20840 8175
rect 20860 8155 20865 8175
rect 20835 8125 20865 8155
rect 20835 8105 20840 8125
rect 20860 8105 20865 8125
rect 20835 8075 20865 8105
rect 20835 8055 20840 8075
rect 20860 8055 20865 8075
rect 20835 8025 20865 8055
rect 20835 8005 20840 8025
rect 20860 8005 20865 8025
rect 20835 7975 20865 8005
rect 20835 7955 20840 7975
rect 20860 7955 20865 7975
rect 20835 7945 20865 7955
rect 20890 8225 20920 8235
rect 20890 8205 20895 8225
rect 20915 8205 20920 8225
rect 20890 8175 20920 8205
rect 20890 8155 20895 8175
rect 20915 8155 20920 8175
rect 20890 8125 20920 8155
rect 20890 8105 20895 8125
rect 20915 8105 20920 8125
rect 20890 8075 20920 8105
rect 20890 8055 20895 8075
rect 20915 8055 20920 8075
rect 20890 8025 20920 8055
rect 20890 8005 20895 8025
rect 20915 8005 20920 8025
rect 20890 7975 20920 8005
rect 20890 7955 20895 7975
rect 20915 7955 20920 7975
rect 20890 7945 20920 7955
rect 20945 8225 20975 8235
rect 20945 8205 20950 8225
rect 20970 8205 20975 8225
rect 20945 8175 20975 8205
rect 20945 8155 20950 8175
rect 20970 8155 20975 8175
rect 20945 8125 20975 8155
rect 20945 8105 20950 8125
rect 20970 8105 20975 8125
rect 20945 8075 20975 8105
rect 20945 8055 20950 8075
rect 20970 8055 20975 8075
rect 20945 8025 20975 8055
rect 20945 8005 20950 8025
rect 20970 8005 20975 8025
rect 20945 7975 20975 8005
rect 20945 7955 20950 7975
rect 20970 7955 20975 7975
rect 20945 7945 20975 7955
rect 21000 8225 21030 8235
rect 21000 8205 21005 8225
rect 21025 8205 21030 8225
rect 21000 8175 21030 8205
rect 21000 8155 21005 8175
rect 21025 8155 21030 8175
rect 21000 8125 21030 8155
rect 21000 8105 21005 8125
rect 21025 8105 21030 8125
rect 21000 8075 21030 8105
rect 21000 8055 21005 8075
rect 21025 8055 21030 8075
rect 21000 8025 21030 8055
rect 21000 8005 21005 8025
rect 21025 8005 21030 8025
rect 21000 7975 21030 8005
rect 21000 7955 21005 7975
rect 21025 7955 21030 7975
rect 21000 7945 21030 7955
rect 21055 8225 21085 8235
rect 21055 8205 21060 8225
rect 21080 8205 21085 8225
rect 21055 8175 21085 8205
rect 21055 8155 21060 8175
rect 21080 8155 21085 8175
rect 21055 8125 21085 8155
rect 21055 8105 21060 8125
rect 21080 8105 21085 8125
rect 21055 8075 21085 8105
rect 21055 8055 21060 8075
rect 21080 8055 21085 8075
rect 21055 8025 21085 8055
rect 21055 8005 21060 8025
rect 21080 8005 21085 8025
rect 21055 7975 21085 8005
rect 21055 7955 21060 7975
rect 21080 7955 21085 7975
rect 21055 7945 21085 7955
rect 21110 8225 21140 8235
rect 21110 8205 21115 8225
rect 21135 8205 21140 8225
rect 21110 8175 21140 8205
rect 21110 8155 21115 8175
rect 21135 8155 21140 8175
rect 21110 8125 21140 8155
rect 21110 8105 21115 8125
rect 21135 8105 21140 8125
rect 21110 8075 21140 8105
rect 21110 8055 21115 8075
rect 21135 8055 21140 8075
rect 21110 8025 21140 8055
rect 21110 8005 21115 8025
rect 21135 8005 21140 8025
rect 21110 7975 21140 8005
rect 21110 7955 21115 7975
rect 21135 7955 21140 7975
rect 21110 7945 21140 7955
rect 21165 8225 21195 8235
rect 21165 8205 21170 8225
rect 21190 8205 21195 8225
rect 21165 8175 21195 8205
rect 21165 8155 21170 8175
rect 21190 8155 21195 8175
rect 21165 8125 21195 8155
rect 21165 8105 21170 8125
rect 21190 8105 21195 8125
rect 21165 8075 21195 8105
rect 21165 8055 21170 8075
rect 21190 8055 21195 8075
rect 21165 8025 21195 8055
rect 21165 8005 21170 8025
rect 21190 8005 21195 8025
rect 21165 7975 21195 8005
rect 21165 7955 21170 7975
rect 21190 7955 21195 7975
rect 21165 7945 21195 7955
rect 21220 8225 21250 8235
rect 21220 8205 21225 8225
rect 21245 8205 21250 8225
rect 21220 8175 21250 8205
rect 21220 8155 21225 8175
rect 21245 8155 21250 8175
rect 21220 8125 21250 8155
rect 21220 8105 21225 8125
rect 21245 8105 21250 8125
rect 21220 8075 21250 8105
rect 21220 8055 21225 8075
rect 21245 8055 21250 8075
rect 21220 8025 21250 8055
rect 21220 8005 21225 8025
rect 21245 8005 21250 8025
rect 21220 7975 21250 8005
rect 21220 7955 21225 7975
rect 21245 7955 21250 7975
rect 21220 7945 21250 7955
rect 21275 8225 21305 8235
rect 21275 8205 21280 8225
rect 21300 8205 21305 8225
rect 21275 8175 21305 8205
rect 21275 8155 21280 8175
rect 21300 8155 21305 8175
rect 21275 8125 21305 8155
rect 21275 8105 21280 8125
rect 21300 8105 21305 8125
rect 21275 8075 21305 8105
rect 21275 8055 21280 8075
rect 21300 8055 21305 8075
rect 21275 8025 21305 8055
rect 21275 8005 21280 8025
rect 21300 8005 21305 8025
rect 21275 7975 21305 8005
rect 21275 7955 21280 7975
rect 21300 7955 21305 7975
rect 21275 7945 21305 7955
rect 21330 8225 21360 8235
rect 21330 8205 21335 8225
rect 21355 8205 21360 8225
rect 21330 8175 21360 8205
rect 21330 8155 21335 8175
rect 21355 8155 21360 8175
rect 21330 8125 21360 8155
rect 21330 8105 21335 8125
rect 21355 8105 21360 8125
rect 21330 8075 21360 8105
rect 21330 8055 21335 8075
rect 21355 8055 21360 8075
rect 21330 8025 21360 8055
rect 21330 8005 21335 8025
rect 21355 8005 21360 8025
rect 21330 7975 21360 8005
rect 21330 7955 21335 7975
rect 21355 7955 21360 7975
rect 21330 7945 21360 7955
rect 21385 8225 21415 8235
rect 21385 8205 21390 8225
rect 21410 8205 21415 8225
rect 21385 8175 21415 8205
rect 21385 8155 21390 8175
rect 21410 8155 21415 8175
rect 21385 8125 21415 8155
rect 21385 8105 21390 8125
rect 21410 8105 21415 8125
rect 21385 8075 21415 8105
rect 21385 8055 21390 8075
rect 21410 8055 21415 8075
rect 21385 8025 21415 8055
rect 21385 8005 21390 8025
rect 21410 8005 21415 8025
rect 21385 7975 21415 8005
rect 21385 7955 21390 7975
rect 21410 7955 21415 7975
rect 21385 7945 21415 7955
rect 21440 8225 21470 8235
rect 21440 8205 21445 8225
rect 21465 8205 21470 8225
rect 21440 8175 21470 8205
rect 21440 8155 21445 8175
rect 21465 8155 21470 8175
rect 21440 8125 21470 8155
rect 21440 8105 21445 8125
rect 21465 8105 21470 8125
rect 21440 8075 21470 8105
rect 21440 8055 21445 8075
rect 21465 8055 21470 8075
rect 21440 8025 21470 8055
rect 21440 8005 21445 8025
rect 21465 8005 21470 8025
rect 21440 7975 21470 8005
rect 21440 7955 21445 7975
rect 21465 7955 21470 7975
rect 21440 7945 21470 7955
rect 21495 8225 21525 8235
rect 21495 8205 21500 8225
rect 21520 8205 21525 8225
rect 21495 8175 21525 8205
rect 21495 8155 21500 8175
rect 21520 8155 21525 8175
rect 21495 8125 21525 8155
rect 21495 8105 21500 8125
rect 21520 8105 21525 8125
rect 21495 8075 21525 8105
rect 21495 8055 21500 8075
rect 21520 8055 21525 8075
rect 21495 8025 21525 8055
rect 21495 8005 21500 8025
rect 21520 8005 21525 8025
rect 21495 7975 21525 8005
rect 21495 7955 21500 7975
rect 21520 7955 21525 7975
rect 21495 7945 21525 7955
rect 21550 8225 21580 8235
rect 21550 8205 21555 8225
rect 21575 8205 21580 8225
rect 21550 8175 21580 8205
rect 21550 8155 21555 8175
rect 21575 8155 21580 8175
rect 21550 8125 21580 8155
rect 21550 8105 21555 8125
rect 21575 8105 21580 8125
rect 21550 8075 21580 8105
rect 21550 8055 21555 8075
rect 21575 8055 21580 8075
rect 21550 8025 21580 8055
rect 21550 8005 21555 8025
rect 21575 8005 21580 8025
rect 21550 7975 21580 8005
rect 21550 7955 21555 7975
rect 21575 7955 21580 7975
rect 21550 7945 21580 7955
rect 21605 8225 21675 8235
rect 21605 8205 21610 8225
rect 21630 8205 21650 8225
rect 21670 8205 21675 8225
rect 21605 8175 21675 8205
rect 21605 8155 21610 8175
rect 21630 8155 21650 8175
rect 21670 8155 21675 8175
rect 21605 8125 21675 8155
rect 21605 8105 21610 8125
rect 21630 8105 21650 8125
rect 21670 8105 21675 8125
rect 21605 8075 21675 8105
rect 21605 8055 21610 8075
rect 21630 8055 21650 8075
rect 21670 8055 21675 8075
rect 21605 8025 21675 8055
rect 21605 8005 21610 8025
rect 21630 8005 21650 8025
rect 21670 8005 21675 8025
rect 21605 7975 21675 8005
rect 21605 7955 21610 7975
rect 21630 7955 21650 7975
rect 21670 7955 21675 7975
rect 21605 7945 21675 7955
rect 20080 7920 20090 7940
rect 20110 7920 20120 7940
rect 20360 7925 20380 7945
rect 20510 7925 20530 7945
rect 20620 7925 20640 7945
rect 20730 7925 20750 7945
rect 20840 7925 20860 7945
rect 20950 7925 20970 7945
rect 21060 7925 21080 7945
rect 21170 7925 21190 7945
rect 21280 7925 21300 7945
rect 21390 7925 21410 7945
rect 21500 7925 21520 7945
rect 21650 7925 21670 7945
rect 20080 7910 20120 7920
rect 20350 7915 20390 7925
rect 14145 7885 14185 7895
rect 18690 7890 18710 7910
rect 18850 7890 18870 7910
rect 18970 7890 18990 7910
rect 19090 7890 19110 7910
rect 19210 7890 19230 7910
rect 19330 7890 19350 7910
rect 19450 7890 19470 7910
rect 19570 7890 19590 7910
rect 19690 7890 19710 7910
rect 19810 7890 19830 7910
rect 19930 7890 19950 7910
rect 20090 7890 20110 7910
rect 20350 7895 20360 7915
rect 20380 7895 20390 7915
rect 12545 7860 12550 7880
rect 12570 7860 12590 7880
rect 12610 7860 12615 7880
rect 12545 7830 12615 7860
rect 18685 7880 18755 7890
rect 18685 7860 18690 7880
rect 18710 7860 18730 7880
rect 18750 7860 18755 7880
rect 12545 7810 12550 7830
rect 12570 7810 12590 7830
rect 12610 7810 12615 7830
rect 12545 7780 12615 7810
rect 12545 7760 12550 7780
rect 12570 7760 12590 7780
rect 12610 7760 12615 7780
rect 12545 7730 12615 7760
rect 12545 7710 12550 7730
rect 12570 7710 12590 7730
rect 12610 7710 12615 7730
rect 12545 7680 12615 7710
rect 13060 7695 13100 7836
rect 13680 7695 13720 7836
rect 18685 7830 18755 7860
rect 18685 7810 18690 7830
rect 18710 7810 18730 7830
rect 18750 7810 18755 7830
rect 18685 7780 18755 7810
rect 18685 7760 18690 7780
rect 18710 7760 18730 7780
rect 18750 7760 18755 7780
rect 18685 7730 18755 7760
rect 18685 7710 18690 7730
rect 18710 7710 18730 7730
rect 18750 7710 18755 7730
rect 12545 7660 12550 7680
rect 12570 7660 12590 7680
rect 12610 7660 12615 7680
rect 18685 7680 18755 7710
rect 12545 7630 12615 7660
rect 12950 7665 12990 7675
rect 12950 7645 12960 7665
rect 12980 7645 12990 7665
rect 12950 7635 12990 7645
rect 13060 7665 13100 7675
rect 13060 7645 13070 7665
rect 13090 7645 13100 7665
rect 13060 7635 13100 7645
rect 13170 7665 13210 7675
rect 13170 7645 13180 7665
rect 13200 7645 13210 7665
rect 13170 7635 13210 7645
rect 13280 7665 13320 7675
rect 13280 7645 13290 7665
rect 13310 7645 13320 7665
rect 13280 7635 13320 7645
rect 13390 7665 13430 7675
rect 13390 7645 13400 7665
rect 13420 7645 13430 7665
rect 13390 7635 13430 7645
rect 13500 7665 13540 7675
rect 13500 7645 13510 7665
rect 13530 7645 13540 7665
rect 13500 7635 13540 7645
rect 13610 7665 13650 7675
rect 13610 7645 13620 7665
rect 13640 7645 13650 7665
rect 13610 7635 13650 7645
rect 13720 7665 13760 7675
rect 13720 7645 13730 7665
rect 13750 7645 13760 7665
rect 13720 7635 13760 7645
rect 13830 7665 13870 7675
rect 13830 7645 13840 7665
rect 13860 7645 13870 7665
rect 13830 7635 13870 7645
rect 13940 7665 13980 7675
rect 13940 7645 13950 7665
rect 13970 7645 13980 7665
rect 13940 7635 13980 7645
rect 14050 7665 14090 7675
rect 14050 7645 14060 7665
rect 14080 7645 14090 7665
rect 14050 7635 14090 7645
rect 17235 7665 17275 7675
rect 17235 7645 17245 7665
rect 17265 7645 17275 7665
rect 17235 7635 17275 7645
rect 17345 7665 17385 7675
rect 17345 7645 17355 7665
rect 17375 7645 17385 7665
rect 17345 7635 17385 7645
rect 17455 7665 17495 7675
rect 17455 7645 17465 7665
rect 17485 7645 17495 7665
rect 17455 7635 17495 7645
rect 17565 7665 17605 7675
rect 17565 7645 17575 7665
rect 17595 7645 17605 7665
rect 17565 7635 17605 7645
rect 17675 7665 17715 7675
rect 17675 7645 17685 7665
rect 17705 7645 17715 7665
rect 17675 7635 17715 7645
rect 17785 7665 17825 7675
rect 17785 7645 17795 7665
rect 17815 7645 17825 7665
rect 17785 7635 17825 7645
rect 17895 7665 17935 7675
rect 17895 7645 17905 7665
rect 17925 7645 17935 7665
rect 17895 7635 17935 7645
rect 18005 7665 18045 7675
rect 18005 7645 18015 7665
rect 18035 7645 18045 7665
rect 18005 7635 18045 7645
rect 18115 7665 18155 7675
rect 18115 7645 18125 7665
rect 18145 7645 18155 7665
rect 18115 7635 18155 7645
rect 18225 7665 18265 7675
rect 18225 7645 18235 7665
rect 18255 7645 18265 7665
rect 18225 7635 18265 7645
rect 18335 7665 18375 7675
rect 18335 7645 18345 7665
rect 18365 7645 18375 7665
rect 18335 7635 18375 7645
rect 18685 7660 18690 7680
rect 18710 7660 18730 7680
rect 18750 7660 18755 7680
rect 12545 7610 12550 7630
rect 12570 7610 12590 7630
rect 12610 7610 12615 7630
rect 12960 7615 12980 7635
rect 13070 7615 13090 7635
rect 13180 7615 13200 7635
rect 13290 7615 13310 7635
rect 13400 7615 13420 7635
rect 13510 7615 13530 7635
rect 13620 7615 13640 7635
rect 13730 7615 13750 7635
rect 13840 7615 13860 7635
rect 13950 7615 13970 7635
rect 14060 7615 14080 7635
rect 17245 7615 17265 7635
rect 17355 7615 17375 7635
rect 17465 7615 17485 7635
rect 17575 7615 17595 7635
rect 17685 7615 17705 7635
rect 17795 7615 17815 7635
rect 17905 7615 17925 7635
rect 18015 7615 18035 7635
rect 18125 7615 18145 7635
rect 18235 7615 18255 7635
rect 18345 7615 18365 7635
rect 18685 7630 18755 7660
rect 12545 7580 12615 7610
rect 12545 7560 12550 7580
rect 12570 7560 12590 7580
rect 12610 7560 12615 7580
rect 12545 7530 12615 7560
rect 12545 7510 12550 7530
rect 12570 7510 12590 7530
rect 12610 7510 12615 7530
rect 12860 7605 12930 7615
rect 12860 7585 12865 7605
rect 12885 7585 12905 7605
rect 12925 7585 12930 7605
rect 12860 7555 12930 7585
rect 12860 7535 12865 7555
rect 12885 7535 12905 7555
rect 12925 7535 12930 7555
rect 12860 7525 12930 7535
rect 12955 7605 12985 7615
rect 12955 7585 12960 7605
rect 12980 7585 12985 7605
rect 12955 7555 12985 7585
rect 12955 7535 12960 7555
rect 12980 7535 12985 7555
rect 12955 7525 12985 7535
rect 13010 7605 13040 7615
rect 13010 7585 13015 7605
rect 13035 7585 13040 7605
rect 13010 7555 13040 7585
rect 13010 7535 13015 7555
rect 13035 7535 13040 7555
rect 13010 7525 13040 7535
rect 13065 7605 13095 7615
rect 13065 7585 13070 7605
rect 13090 7585 13095 7605
rect 13065 7555 13095 7585
rect 13065 7535 13070 7555
rect 13090 7535 13095 7555
rect 13065 7525 13095 7535
rect 13120 7605 13150 7615
rect 13120 7585 13125 7605
rect 13145 7585 13150 7605
rect 13120 7555 13150 7585
rect 13120 7535 13125 7555
rect 13145 7535 13150 7555
rect 13120 7525 13150 7535
rect 13175 7605 13205 7615
rect 13175 7585 13180 7605
rect 13200 7585 13205 7605
rect 13175 7555 13205 7585
rect 13175 7535 13180 7555
rect 13200 7535 13205 7555
rect 13175 7525 13205 7535
rect 13230 7605 13260 7615
rect 13230 7585 13235 7605
rect 13255 7585 13260 7605
rect 13230 7555 13260 7585
rect 13230 7535 13235 7555
rect 13255 7535 13260 7555
rect 13230 7525 13260 7535
rect 13285 7605 13315 7615
rect 13285 7585 13290 7605
rect 13310 7585 13315 7605
rect 13285 7555 13315 7585
rect 13285 7535 13290 7555
rect 13310 7535 13315 7555
rect 13285 7525 13315 7535
rect 13340 7605 13370 7615
rect 13340 7585 13345 7605
rect 13365 7585 13370 7605
rect 13340 7555 13370 7585
rect 13340 7535 13345 7555
rect 13365 7535 13370 7555
rect 13340 7525 13370 7535
rect 13395 7605 13425 7615
rect 13395 7585 13400 7605
rect 13420 7585 13425 7605
rect 13395 7555 13425 7585
rect 13395 7535 13400 7555
rect 13420 7535 13425 7555
rect 13395 7525 13425 7535
rect 13450 7605 13480 7615
rect 13450 7585 13455 7605
rect 13475 7585 13480 7605
rect 13450 7555 13480 7585
rect 13450 7535 13455 7555
rect 13475 7535 13480 7555
rect 13450 7525 13480 7535
rect 13505 7605 13535 7615
rect 13505 7585 13510 7605
rect 13530 7585 13535 7605
rect 13505 7555 13535 7585
rect 13505 7535 13510 7555
rect 13530 7535 13535 7555
rect 13505 7525 13535 7535
rect 13560 7605 13590 7615
rect 13560 7585 13565 7605
rect 13585 7585 13590 7605
rect 13560 7555 13590 7585
rect 13560 7535 13565 7555
rect 13585 7535 13590 7555
rect 13560 7525 13590 7535
rect 13615 7605 13645 7615
rect 13615 7585 13620 7605
rect 13640 7585 13645 7605
rect 13615 7555 13645 7585
rect 13615 7535 13620 7555
rect 13640 7535 13645 7555
rect 13615 7525 13645 7535
rect 13670 7605 13700 7615
rect 13670 7585 13675 7605
rect 13695 7585 13700 7605
rect 13670 7555 13700 7585
rect 13670 7535 13675 7555
rect 13695 7535 13700 7555
rect 13670 7525 13700 7535
rect 13725 7605 13755 7615
rect 13725 7585 13730 7605
rect 13750 7585 13755 7605
rect 13725 7555 13755 7585
rect 13725 7535 13730 7555
rect 13750 7535 13755 7555
rect 13725 7525 13755 7535
rect 13780 7605 13810 7615
rect 13780 7585 13785 7605
rect 13805 7585 13810 7605
rect 13780 7555 13810 7585
rect 13780 7535 13785 7555
rect 13805 7535 13810 7555
rect 13780 7525 13810 7535
rect 13835 7605 13865 7615
rect 13835 7585 13840 7605
rect 13860 7585 13865 7605
rect 13835 7555 13865 7585
rect 13835 7535 13840 7555
rect 13860 7535 13865 7555
rect 13835 7525 13865 7535
rect 13890 7605 13920 7615
rect 13890 7585 13895 7605
rect 13915 7585 13920 7605
rect 13890 7555 13920 7585
rect 13890 7535 13895 7555
rect 13915 7535 13920 7555
rect 13890 7525 13920 7535
rect 13945 7605 13975 7615
rect 13945 7585 13950 7605
rect 13970 7585 13975 7605
rect 13945 7555 13975 7585
rect 13945 7535 13950 7555
rect 13970 7535 13975 7555
rect 13945 7525 13975 7535
rect 14000 7605 14030 7615
rect 14000 7585 14005 7605
rect 14025 7585 14030 7605
rect 14000 7555 14030 7585
rect 14000 7535 14005 7555
rect 14025 7535 14030 7555
rect 14000 7525 14030 7535
rect 14055 7605 14085 7615
rect 14055 7585 14060 7605
rect 14080 7585 14085 7605
rect 14055 7555 14085 7585
rect 14055 7535 14060 7555
rect 14080 7535 14085 7555
rect 14055 7525 14085 7535
rect 14110 7605 14180 7615
rect 14110 7585 14115 7605
rect 14135 7585 14155 7605
rect 14175 7585 14180 7605
rect 14110 7555 14180 7585
rect 14110 7535 14115 7555
rect 14135 7535 14155 7555
rect 14175 7535 14180 7555
rect 14110 7525 14180 7535
rect 17145 7605 17215 7615
rect 17145 7585 17150 7605
rect 17170 7585 17190 7605
rect 17210 7585 17215 7605
rect 17145 7555 17215 7585
rect 17145 7535 17150 7555
rect 17170 7535 17190 7555
rect 17210 7535 17215 7555
rect 17145 7525 17215 7535
rect 17240 7605 17270 7615
rect 17240 7585 17245 7605
rect 17265 7585 17270 7605
rect 17240 7555 17270 7585
rect 17240 7535 17245 7555
rect 17265 7535 17270 7555
rect 17240 7525 17270 7535
rect 17295 7605 17325 7615
rect 17295 7585 17300 7605
rect 17320 7585 17325 7605
rect 17295 7555 17325 7585
rect 17295 7535 17300 7555
rect 17320 7535 17325 7555
rect 17295 7525 17325 7535
rect 17350 7605 17380 7615
rect 17350 7585 17355 7605
rect 17375 7585 17380 7605
rect 17350 7555 17380 7585
rect 17350 7535 17355 7555
rect 17375 7535 17380 7555
rect 17350 7525 17380 7535
rect 17405 7605 17435 7615
rect 17405 7585 17410 7605
rect 17430 7585 17435 7605
rect 17405 7555 17435 7585
rect 17405 7535 17410 7555
rect 17430 7535 17435 7555
rect 17405 7525 17435 7535
rect 17460 7605 17490 7615
rect 17460 7585 17465 7605
rect 17485 7585 17490 7605
rect 17460 7555 17490 7585
rect 17460 7535 17465 7555
rect 17485 7535 17490 7555
rect 17460 7525 17490 7535
rect 17515 7605 17545 7615
rect 17515 7585 17520 7605
rect 17540 7585 17545 7605
rect 17515 7555 17545 7585
rect 17515 7535 17520 7555
rect 17540 7535 17545 7555
rect 17515 7525 17545 7535
rect 17570 7605 17600 7615
rect 17570 7585 17575 7605
rect 17595 7585 17600 7605
rect 17570 7555 17600 7585
rect 17570 7535 17575 7555
rect 17595 7535 17600 7555
rect 17570 7525 17600 7535
rect 17625 7605 17655 7615
rect 17625 7585 17630 7605
rect 17650 7585 17655 7605
rect 17625 7555 17655 7585
rect 17625 7535 17630 7555
rect 17650 7535 17655 7555
rect 17625 7525 17655 7535
rect 17680 7605 17710 7615
rect 17680 7585 17685 7605
rect 17705 7585 17710 7605
rect 17680 7555 17710 7585
rect 17680 7535 17685 7555
rect 17705 7535 17710 7555
rect 17680 7525 17710 7535
rect 17735 7605 17765 7615
rect 17735 7585 17740 7605
rect 17760 7585 17765 7605
rect 17735 7555 17765 7585
rect 17735 7535 17740 7555
rect 17760 7535 17765 7555
rect 17735 7525 17765 7535
rect 17790 7605 17820 7615
rect 17790 7585 17795 7605
rect 17815 7585 17820 7605
rect 17790 7555 17820 7585
rect 17790 7535 17795 7555
rect 17815 7535 17820 7555
rect 17790 7525 17820 7535
rect 17845 7605 17875 7615
rect 17845 7585 17850 7605
rect 17870 7585 17875 7605
rect 17845 7555 17875 7585
rect 17845 7535 17850 7555
rect 17870 7535 17875 7555
rect 17845 7525 17875 7535
rect 17900 7605 17930 7615
rect 17900 7585 17905 7605
rect 17925 7585 17930 7605
rect 17900 7555 17930 7585
rect 17900 7535 17905 7555
rect 17925 7535 17930 7555
rect 17900 7525 17930 7535
rect 17955 7605 17985 7615
rect 17955 7585 17960 7605
rect 17980 7585 17985 7605
rect 17955 7555 17985 7585
rect 17955 7535 17960 7555
rect 17980 7535 17985 7555
rect 17955 7525 17985 7535
rect 18010 7605 18040 7615
rect 18010 7585 18015 7605
rect 18035 7585 18040 7605
rect 18010 7555 18040 7585
rect 18010 7535 18015 7555
rect 18035 7535 18040 7555
rect 18010 7525 18040 7535
rect 18065 7605 18095 7615
rect 18065 7585 18070 7605
rect 18090 7585 18095 7605
rect 18065 7555 18095 7585
rect 18065 7535 18070 7555
rect 18090 7535 18095 7555
rect 18065 7525 18095 7535
rect 18120 7605 18150 7615
rect 18120 7585 18125 7605
rect 18145 7585 18150 7605
rect 18120 7555 18150 7585
rect 18120 7535 18125 7555
rect 18145 7535 18150 7555
rect 18120 7525 18150 7535
rect 18175 7605 18205 7615
rect 18175 7585 18180 7605
rect 18200 7585 18205 7605
rect 18175 7555 18205 7585
rect 18175 7535 18180 7555
rect 18200 7535 18205 7555
rect 18175 7525 18205 7535
rect 18230 7605 18260 7615
rect 18230 7585 18235 7605
rect 18255 7585 18260 7605
rect 18230 7555 18260 7585
rect 18230 7535 18235 7555
rect 18255 7535 18260 7555
rect 18230 7525 18260 7535
rect 18285 7605 18315 7615
rect 18285 7585 18290 7605
rect 18310 7585 18315 7605
rect 18285 7555 18315 7585
rect 18285 7535 18290 7555
rect 18310 7535 18315 7555
rect 18285 7525 18315 7535
rect 18340 7605 18370 7615
rect 18340 7585 18345 7605
rect 18365 7585 18370 7605
rect 18340 7555 18370 7585
rect 18340 7535 18345 7555
rect 18365 7535 18370 7555
rect 18340 7525 18370 7535
rect 18395 7605 18465 7615
rect 18395 7585 18400 7605
rect 18420 7585 18440 7605
rect 18460 7585 18465 7605
rect 18395 7555 18465 7585
rect 18395 7535 18400 7555
rect 18420 7535 18440 7555
rect 18460 7535 18465 7555
rect 18395 7525 18465 7535
rect 18685 7610 18690 7630
rect 18710 7610 18730 7630
rect 18750 7610 18755 7630
rect 18685 7580 18755 7610
rect 18685 7560 18690 7580
rect 18710 7560 18730 7580
rect 18750 7560 18755 7580
rect 18685 7530 18755 7560
rect 12545 7500 12615 7510
rect 12865 7505 12885 7525
rect 13015 7505 13035 7525
rect 13125 7505 13145 7525
rect 13235 7505 13255 7525
rect 13345 7505 13365 7525
rect 13455 7505 13475 7525
rect 13565 7505 13585 7525
rect 13675 7505 13695 7525
rect 13785 7505 13805 7525
rect 13895 7505 13915 7525
rect 14005 7505 14025 7525
rect 14155 7505 14175 7525
rect 17150 7505 17170 7525
rect 17300 7505 17320 7525
rect 17410 7505 17430 7525
rect 17520 7505 17540 7525
rect 17630 7505 17650 7525
rect 17740 7505 17760 7525
rect 17850 7505 17870 7525
rect 17960 7505 17980 7525
rect 18070 7505 18090 7525
rect 18180 7505 18200 7525
rect 18290 7505 18310 7525
rect 18440 7505 18460 7525
rect 18685 7510 18690 7530
rect 18710 7510 18730 7530
rect 18750 7510 18755 7530
rect 10930 7475 10940 7495
rect 10960 7475 10970 7495
rect 11290 7480 11310 7500
rect 11410 7480 11430 7500
rect 11530 7480 11550 7500
rect 11650 7480 11670 7500
rect 11770 7480 11790 7500
rect 11890 7480 11910 7500
rect 12010 7480 12030 7500
rect 12130 7480 12150 7500
rect 12250 7480 12270 7500
rect 12370 7480 12390 7500
rect 12490 7480 12510 7500
rect 12855 7495 12895 7505
rect 10930 7465 10970 7475
rect 11280 7470 11320 7480
rect 11280 7450 11290 7470
rect 11310 7450 11320 7470
rect 10813 7435 10847 7445
rect 11280 7440 11320 7450
rect 11400 7470 11440 7480
rect 11400 7450 11410 7470
rect 11430 7450 11440 7470
rect 11400 7440 11440 7450
rect 11520 7470 11560 7480
rect 11520 7450 11530 7470
rect 11550 7450 11560 7470
rect 11520 7440 11560 7450
rect 11640 7470 11680 7480
rect 11640 7450 11650 7470
rect 11670 7450 11680 7470
rect 11640 7440 11680 7450
rect 11760 7470 11800 7480
rect 11760 7450 11770 7470
rect 11790 7450 11800 7470
rect 11760 7440 11800 7450
rect 11823 7470 11857 7480
rect 11823 7450 11831 7470
rect 11849 7450 11857 7470
rect 11823 7440 11857 7450
rect 11880 7470 11920 7480
rect 11880 7450 11890 7470
rect 11910 7450 11920 7470
rect 11880 7440 11920 7450
rect 12000 7470 12040 7480
rect 12000 7450 12010 7470
rect 12030 7450 12040 7470
rect 12000 7440 12040 7450
rect 12120 7470 12160 7480
rect 12120 7450 12130 7470
rect 12150 7450 12160 7470
rect 12120 7440 12160 7450
rect 12240 7470 12280 7480
rect 12240 7450 12250 7470
rect 12270 7450 12280 7470
rect 12240 7440 12280 7450
rect 12360 7470 12400 7480
rect 12360 7450 12370 7470
rect 12390 7450 12400 7470
rect 12360 7440 12400 7450
rect 12480 7470 12520 7480
rect 12480 7450 12490 7470
rect 12510 7450 12520 7470
rect 12855 7475 12865 7495
rect 12885 7475 12895 7495
rect 12855 7465 12895 7475
rect 13005 7495 13045 7505
rect 13005 7475 13015 7495
rect 13035 7475 13045 7495
rect 13005 7465 13045 7475
rect 13115 7495 13155 7505
rect 13115 7475 13125 7495
rect 13145 7475 13155 7495
rect 13115 7465 13155 7475
rect 13225 7495 13265 7505
rect 13225 7475 13235 7495
rect 13255 7475 13265 7495
rect 13225 7465 13265 7475
rect 13335 7495 13375 7505
rect 13335 7475 13345 7495
rect 13365 7475 13375 7495
rect 13335 7465 13375 7475
rect 13445 7495 13485 7505
rect 13445 7475 13455 7495
rect 13475 7475 13485 7495
rect 13445 7465 13485 7475
rect 13555 7495 13595 7505
rect 13555 7475 13565 7495
rect 13585 7475 13595 7495
rect 13555 7465 13595 7475
rect 13665 7495 13705 7505
rect 13665 7475 13675 7495
rect 13695 7475 13705 7495
rect 13665 7465 13705 7475
rect 13775 7495 13815 7505
rect 13775 7475 13785 7495
rect 13805 7475 13815 7495
rect 13775 7465 13815 7475
rect 13885 7495 13925 7505
rect 13885 7475 13895 7495
rect 13915 7475 13925 7495
rect 13885 7465 13925 7475
rect 13995 7495 14035 7505
rect 13995 7475 14005 7495
rect 14025 7475 14035 7495
rect 13995 7465 14035 7475
rect 14145 7495 14185 7505
rect 14145 7475 14155 7495
rect 14175 7475 14185 7495
rect 14145 7465 14185 7475
rect 17140 7495 17180 7505
rect 17140 7475 17150 7495
rect 17170 7475 17180 7495
rect 17140 7465 17180 7475
rect 17290 7495 17330 7505
rect 17290 7475 17300 7495
rect 17320 7475 17330 7495
rect 17290 7465 17330 7475
rect 17400 7495 17440 7505
rect 17400 7475 17410 7495
rect 17430 7475 17440 7495
rect 17400 7465 17440 7475
rect 17510 7495 17550 7505
rect 17510 7475 17520 7495
rect 17540 7475 17550 7495
rect 17510 7465 17550 7475
rect 17620 7495 17660 7505
rect 17620 7475 17630 7495
rect 17650 7475 17660 7495
rect 17620 7465 17660 7475
rect 17730 7495 17770 7505
rect 17730 7475 17740 7495
rect 17760 7475 17770 7495
rect 17730 7465 17770 7475
rect 17840 7495 17880 7505
rect 17840 7475 17850 7495
rect 17870 7475 17880 7495
rect 17840 7465 17880 7475
rect 17950 7495 17990 7505
rect 17950 7475 17960 7495
rect 17980 7475 17990 7495
rect 17950 7465 17990 7475
rect 18060 7495 18100 7505
rect 18060 7475 18070 7495
rect 18090 7475 18100 7495
rect 18060 7465 18100 7475
rect 18170 7495 18210 7505
rect 18170 7475 18180 7495
rect 18200 7475 18210 7495
rect 18170 7465 18210 7475
rect 18280 7495 18320 7505
rect 18280 7475 18290 7495
rect 18310 7475 18320 7495
rect 18280 7465 18320 7475
rect 18430 7495 18470 7505
rect 18685 7500 18755 7510
rect 18785 7880 18815 7890
rect 18785 7860 18790 7880
rect 18810 7860 18815 7880
rect 18785 7830 18815 7860
rect 18785 7810 18790 7830
rect 18810 7810 18815 7830
rect 18785 7780 18815 7810
rect 18785 7760 18790 7780
rect 18810 7760 18815 7780
rect 18785 7730 18815 7760
rect 18785 7710 18790 7730
rect 18810 7710 18815 7730
rect 18785 7680 18815 7710
rect 18785 7660 18790 7680
rect 18810 7660 18815 7680
rect 18785 7630 18815 7660
rect 18785 7610 18790 7630
rect 18810 7610 18815 7630
rect 18785 7580 18815 7610
rect 18785 7560 18790 7580
rect 18810 7560 18815 7580
rect 18785 7530 18815 7560
rect 18785 7510 18790 7530
rect 18810 7510 18815 7530
rect 18785 7500 18815 7510
rect 18845 7880 18875 7890
rect 18845 7860 18850 7880
rect 18870 7860 18875 7880
rect 18845 7830 18875 7860
rect 18845 7810 18850 7830
rect 18870 7810 18875 7830
rect 18845 7780 18875 7810
rect 18845 7760 18850 7780
rect 18870 7760 18875 7780
rect 18845 7730 18875 7760
rect 18845 7710 18850 7730
rect 18870 7710 18875 7730
rect 18845 7680 18875 7710
rect 18845 7660 18850 7680
rect 18870 7660 18875 7680
rect 18845 7630 18875 7660
rect 18845 7610 18850 7630
rect 18870 7610 18875 7630
rect 18845 7580 18875 7610
rect 18845 7560 18850 7580
rect 18870 7560 18875 7580
rect 18845 7530 18875 7560
rect 18845 7510 18850 7530
rect 18870 7510 18875 7530
rect 18845 7500 18875 7510
rect 18905 7880 18935 7890
rect 18905 7860 18910 7880
rect 18930 7860 18935 7880
rect 18905 7830 18935 7860
rect 18905 7810 18910 7830
rect 18930 7810 18935 7830
rect 18905 7780 18935 7810
rect 18905 7760 18910 7780
rect 18930 7760 18935 7780
rect 18905 7730 18935 7760
rect 18905 7710 18910 7730
rect 18930 7710 18935 7730
rect 18905 7680 18935 7710
rect 18905 7660 18910 7680
rect 18930 7660 18935 7680
rect 18905 7630 18935 7660
rect 18905 7610 18910 7630
rect 18930 7610 18935 7630
rect 18905 7580 18935 7610
rect 18905 7560 18910 7580
rect 18930 7560 18935 7580
rect 18905 7530 18935 7560
rect 18905 7510 18910 7530
rect 18930 7510 18935 7530
rect 18905 7500 18935 7510
rect 18965 7880 18995 7890
rect 18965 7860 18970 7880
rect 18990 7860 18995 7880
rect 18965 7830 18995 7860
rect 18965 7810 18970 7830
rect 18990 7810 18995 7830
rect 18965 7780 18995 7810
rect 18965 7760 18970 7780
rect 18990 7760 18995 7780
rect 18965 7730 18995 7760
rect 18965 7710 18970 7730
rect 18990 7710 18995 7730
rect 18965 7680 18995 7710
rect 18965 7660 18970 7680
rect 18990 7660 18995 7680
rect 18965 7630 18995 7660
rect 18965 7610 18970 7630
rect 18990 7610 18995 7630
rect 18965 7580 18995 7610
rect 18965 7560 18970 7580
rect 18990 7560 18995 7580
rect 18965 7530 18995 7560
rect 18965 7510 18970 7530
rect 18990 7510 18995 7530
rect 18965 7500 18995 7510
rect 19025 7880 19055 7890
rect 19025 7860 19030 7880
rect 19050 7860 19055 7880
rect 19025 7830 19055 7860
rect 19025 7810 19030 7830
rect 19050 7810 19055 7830
rect 19025 7780 19055 7810
rect 19025 7760 19030 7780
rect 19050 7760 19055 7780
rect 19025 7730 19055 7760
rect 19025 7710 19030 7730
rect 19050 7710 19055 7730
rect 19025 7680 19055 7710
rect 19025 7660 19030 7680
rect 19050 7660 19055 7680
rect 19025 7630 19055 7660
rect 19025 7610 19030 7630
rect 19050 7610 19055 7630
rect 19025 7580 19055 7610
rect 19025 7560 19030 7580
rect 19050 7560 19055 7580
rect 19025 7530 19055 7560
rect 19025 7510 19030 7530
rect 19050 7510 19055 7530
rect 19025 7500 19055 7510
rect 19085 7880 19115 7890
rect 19085 7860 19090 7880
rect 19110 7860 19115 7880
rect 19085 7830 19115 7860
rect 19085 7810 19090 7830
rect 19110 7810 19115 7830
rect 19085 7780 19115 7810
rect 19085 7760 19090 7780
rect 19110 7760 19115 7780
rect 19085 7730 19115 7760
rect 19085 7710 19090 7730
rect 19110 7710 19115 7730
rect 19085 7680 19115 7710
rect 19085 7660 19090 7680
rect 19110 7660 19115 7680
rect 19085 7630 19115 7660
rect 19085 7610 19090 7630
rect 19110 7610 19115 7630
rect 19085 7580 19115 7610
rect 19085 7560 19090 7580
rect 19110 7560 19115 7580
rect 19085 7530 19115 7560
rect 19085 7510 19090 7530
rect 19110 7510 19115 7530
rect 19085 7500 19115 7510
rect 19145 7880 19175 7890
rect 19145 7860 19150 7880
rect 19170 7860 19175 7880
rect 19145 7830 19175 7860
rect 19145 7810 19150 7830
rect 19170 7810 19175 7830
rect 19145 7780 19175 7810
rect 19145 7760 19150 7780
rect 19170 7760 19175 7780
rect 19145 7730 19175 7760
rect 19145 7710 19150 7730
rect 19170 7710 19175 7730
rect 19145 7680 19175 7710
rect 19145 7660 19150 7680
rect 19170 7660 19175 7680
rect 19145 7630 19175 7660
rect 19145 7610 19150 7630
rect 19170 7610 19175 7630
rect 19145 7580 19175 7610
rect 19145 7560 19150 7580
rect 19170 7560 19175 7580
rect 19145 7530 19175 7560
rect 19145 7510 19150 7530
rect 19170 7510 19175 7530
rect 19145 7500 19175 7510
rect 19205 7880 19235 7890
rect 19205 7860 19210 7880
rect 19230 7860 19235 7880
rect 19205 7830 19235 7860
rect 19205 7810 19210 7830
rect 19230 7810 19235 7830
rect 19205 7780 19235 7810
rect 19205 7760 19210 7780
rect 19230 7760 19235 7780
rect 19205 7730 19235 7760
rect 19205 7710 19210 7730
rect 19230 7710 19235 7730
rect 19205 7680 19235 7710
rect 19205 7660 19210 7680
rect 19230 7660 19235 7680
rect 19205 7630 19235 7660
rect 19205 7610 19210 7630
rect 19230 7610 19235 7630
rect 19205 7580 19235 7610
rect 19205 7560 19210 7580
rect 19230 7560 19235 7580
rect 19205 7530 19235 7560
rect 19205 7510 19210 7530
rect 19230 7510 19235 7530
rect 19205 7500 19235 7510
rect 19265 7880 19295 7890
rect 19265 7860 19270 7880
rect 19290 7860 19295 7880
rect 19265 7830 19295 7860
rect 19265 7810 19270 7830
rect 19290 7810 19295 7830
rect 19265 7780 19295 7810
rect 19265 7760 19270 7780
rect 19290 7760 19295 7780
rect 19265 7730 19295 7760
rect 19265 7710 19270 7730
rect 19290 7710 19295 7730
rect 19265 7680 19295 7710
rect 19265 7660 19270 7680
rect 19290 7660 19295 7680
rect 19265 7630 19295 7660
rect 19265 7610 19270 7630
rect 19290 7610 19295 7630
rect 19265 7580 19295 7610
rect 19265 7560 19270 7580
rect 19290 7560 19295 7580
rect 19265 7530 19295 7560
rect 19265 7510 19270 7530
rect 19290 7510 19295 7530
rect 19265 7500 19295 7510
rect 19325 7880 19355 7890
rect 19325 7860 19330 7880
rect 19350 7860 19355 7880
rect 19325 7830 19355 7860
rect 19325 7810 19330 7830
rect 19350 7810 19355 7830
rect 19325 7780 19355 7810
rect 19325 7760 19330 7780
rect 19350 7760 19355 7780
rect 19325 7730 19355 7760
rect 19325 7710 19330 7730
rect 19350 7710 19355 7730
rect 19325 7680 19355 7710
rect 19325 7660 19330 7680
rect 19350 7660 19355 7680
rect 19325 7630 19355 7660
rect 19325 7610 19330 7630
rect 19350 7610 19355 7630
rect 19325 7580 19355 7610
rect 19325 7560 19330 7580
rect 19350 7560 19355 7580
rect 19325 7530 19355 7560
rect 19325 7510 19330 7530
rect 19350 7510 19355 7530
rect 19325 7500 19355 7510
rect 19385 7880 19415 7890
rect 19385 7860 19390 7880
rect 19410 7860 19415 7880
rect 19385 7830 19415 7860
rect 19385 7810 19390 7830
rect 19410 7810 19415 7830
rect 19385 7780 19415 7810
rect 19385 7760 19390 7780
rect 19410 7760 19415 7780
rect 19385 7730 19415 7760
rect 19385 7710 19390 7730
rect 19410 7710 19415 7730
rect 19385 7680 19415 7710
rect 19385 7660 19390 7680
rect 19410 7660 19415 7680
rect 19385 7630 19415 7660
rect 19385 7610 19390 7630
rect 19410 7610 19415 7630
rect 19385 7580 19415 7610
rect 19385 7560 19390 7580
rect 19410 7560 19415 7580
rect 19385 7530 19415 7560
rect 19385 7510 19390 7530
rect 19410 7510 19415 7530
rect 19385 7500 19415 7510
rect 19445 7880 19475 7890
rect 19445 7860 19450 7880
rect 19470 7860 19475 7880
rect 19445 7830 19475 7860
rect 19445 7810 19450 7830
rect 19470 7810 19475 7830
rect 19445 7780 19475 7810
rect 19445 7760 19450 7780
rect 19470 7760 19475 7780
rect 19445 7730 19475 7760
rect 19445 7710 19450 7730
rect 19470 7710 19475 7730
rect 19445 7680 19475 7710
rect 19445 7660 19450 7680
rect 19470 7660 19475 7680
rect 19445 7630 19475 7660
rect 19445 7610 19450 7630
rect 19470 7610 19475 7630
rect 19445 7580 19475 7610
rect 19445 7560 19450 7580
rect 19470 7560 19475 7580
rect 19445 7530 19475 7560
rect 19445 7510 19450 7530
rect 19470 7510 19475 7530
rect 19445 7500 19475 7510
rect 19505 7880 19535 7890
rect 19505 7860 19510 7880
rect 19530 7860 19535 7880
rect 19505 7830 19535 7860
rect 19505 7810 19510 7830
rect 19530 7810 19535 7830
rect 19505 7780 19535 7810
rect 19505 7760 19510 7780
rect 19530 7760 19535 7780
rect 19505 7730 19535 7760
rect 19505 7710 19510 7730
rect 19530 7710 19535 7730
rect 19505 7680 19535 7710
rect 19505 7660 19510 7680
rect 19530 7660 19535 7680
rect 19505 7630 19535 7660
rect 19505 7610 19510 7630
rect 19530 7610 19535 7630
rect 19505 7580 19535 7610
rect 19505 7560 19510 7580
rect 19530 7560 19535 7580
rect 19505 7530 19535 7560
rect 19505 7510 19510 7530
rect 19530 7510 19535 7530
rect 19505 7500 19535 7510
rect 19565 7880 19595 7890
rect 19565 7860 19570 7880
rect 19590 7860 19595 7880
rect 19565 7830 19595 7860
rect 19565 7810 19570 7830
rect 19590 7810 19595 7830
rect 19565 7780 19595 7810
rect 19565 7760 19570 7780
rect 19590 7760 19595 7780
rect 19565 7730 19595 7760
rect 19565 7710 19570 7730
rect 19590 7710 19595 7730
rect 19565 7680 19595 7710
rect 19565 7660 19570 7680
rect 19590 7660 19595 7680
rect 19565 7630 19595 7660
rect 19565 7610 19570 7630
rect 19590 7610 19595 7630
rect 19565 7580 19595 7610
rect 19565 7560 19570 7580
rect 19590 7560 19595 7580
rect 19565 7530 19595 7560
rect 19565 7510 19570 7530
rect 19590 7510 19595 7530
rect 19565 7500 19595 7510
rect 19625 7880 19655 7890
rect 19625 7860 19630 7880
rect 19650 7860 19655 7880
rect 19625 7830 19655 7860
rect 19625 7810 19630 7830
rect 19650 7810 19655 7830
rect 19625 7780 19655 7810
rect 19625 7760 19630 7780
rect 19650 7760 19655 7780
rect 19625 7730 19655 7760
rect 19625 7710 19630 7730
rect 19650 7710 19655 7730
rect 19625 7680 19655 7710
rect 19625 7660 19630 7680
rect 19650 7660 19655 7680
rect 19625 7630 19655 7660
rect 19625 7610 19630 7630
rect 19650 7610 19655 7630
rect 19625 7580 19655 7610
rect 19625 7560 19630 7580
rect 19650 7560 19655 7580
rect 19625 7530 19655 7560
rect 19625 7510 19630 7530
rect 19650 7510 19655 7530
rect 19625 7500 19655 7510
rect 19685 7880 19715 7890
rect 19685 7860 19690 7880
rect 19710 7860 19715 7880
rect 19685 7830 19715 7860
rect 19685 7810 19690 7830
rect 19710 7810 19715 7830
rect 19685 7780 19715 7810
rect 19685 7760 19690 7780
rect 19710 7760 19715 7780
rect 19685 7730 19715 7760
rect 19685 7710 19690 7730
rect 19710 7710 19715 7730
rect 19685 7680 19715 7710
rect 19685 7660 19690 7680
rect 19710 7660 19715 7680
rect 19685 7630 19715 7660
rect 19685 7610 19690 7630
rect 19710 7610 19715 7630
rect 19685 7580 19715 7610
rect 19685 7560 19690 7580
rect 19710 7560 19715 7580
rect 19685 7530 19715 7560
rect 19685 7510 19690 7530
rect 19710 7510 19715 7530
rect 19685 7500 19715 7510
rect 19745 7880 19775 7890
rect 19745 7860 19750 7880
rect 19770 7860 19775 7880
rect 19745 7830 19775 7860
rect 19745 7810 19750 7830
rect 19770 7810 19775 7830
rect 19745 7780 19775 7810
rect 19745 7760 19750 7780
rect 19770 7760 19775 7780
rect 19745 7730 19775 7760
rect 19745 7710 19750 7730
rect 19770 7710 19775 7730
rect 19745 7680 19775 7710
rect 19745 7660 19750 7680
rect 19770 7660 19775 7680
rect 19745 7630 19775 7660
rect 19745 7610 19750 7630
rect 19770 7610 19775 7630
rect 19745 7580 19775 7610
rect 19745 7560 19750 7580
rect 19770 7560 19775 7580
rect 19745 7530 19775 7560
rect 19745 7510 19750 7530
rect 19770 7510 19775 7530
rect 19745 7500 19775 7510
rect 19805 7880 19835 7890
rect 19805 7860 19810 7880
rect 19830 7860 19835 7880
rect 19805 7830 19835 7860
rect 19805 7810 19810 7830
rect 19830 7810 19835 7830
rect 19805 7780 19835 7810
rect 19805 7760 19810 7780
rect 19830 7760 19835 7780
rect 19805 7730 19835 7760
rect 19805 7710 19810 7730
rect 19830 7710 19835 7730
rect 19805 7680 19835 7710
rect 19805 7660 19810 7680
rect 19830 7660 19835 7680
rect 19805 7630 19835 7660
rect 19805 7610 19810 7630
rect 19830 7610 19835 7630
rect 19805 7580 19835 7610
rect 19805 7560 19810 7580
rect 19830 7560 19835 7580
rect 19805 7530 19835 7560
rect 19805 7510 19810 7530
rect 19830 7510 19835 7530
rect 19805 7500 19835 7510
rect 19865 7880 19895 7890
rect 19865 7860 19870 7880
rect 19890 7860 19895 7880
rect 19865 7830 19895 7860
rect 19865 7810 19870 7830
rect 19890 7810 19895 7830
rect 19865 7780 19895 7810
rect 19865 7760 19870 7780
rect 19890 7760 19895 7780
rect 19865 7730 19895 7760
rect 19865 7710 19870 7730
rect 19890 7710 19895 7730
rect 19865 7680 19895 7710
rect 19865 7660 19870 7680
rect 19890 7660 19895 7680
rect 19865 7630 19895 7660
rect 19865 7610 19870 7630
rect 19890 7610 19895 7630
rect 19865 7580 19895 7610
rect 19865 7560 19870 7580
rect 19890 7560 19895 7580
rect 19865 7530 19895 7560
rect 19865 7510 19870 7530
rect 19890 7510 19895 7530
rect 19865 7500 19895 7510
rect 19925 7880 19955 7890
rect 19925 7860 19930 7880
rect 19950 7860 19955 7880
rect 19925 7830 19955 7860
rect 19925 7810 19930 7830
rect 19950 7810 19955 7830
rect 19925 7780 19955 7810
rect 19925 7760 19930 7780
rect 19950 7760 19955 7780
rect 19925 7730 19955 7760
rect 19925 7710 19930 7730
rect 19950 7710 19955 7730
rect 19925 7680 19955 7710
rect 19925 7660 19930 7680
rect 19950 7660 19955 7680
rect 19925 7630 19955 7660
rect 19925 7610 19930 7630
rect 19950 7610 19955 7630
rect 19925 7580 19955 7610
rect 19925 7560 19930 7580
rect 19950 7560 19955 7580
rect 19925 7530 19955 7560
rect 19925 7510 19930 7530
rect 19950 7510 19955 7530
rect 19925 7500 19955 7510
rect 19985 7880 20015 7890
rect 19985 7860 19990 7880
rect 20010 7860 20015 7880
rect 19985 7830 20015 7860
rect 19985 7810 19990 7830
rect 20010 7810 20015 7830
rect 19985 7780 20015 7810
rect 19985 7760 19990 7780
rect 20010 7760 20015 7780
rect 19985 7730 20015 7760
rect 19985 7710 19990 7730
rect 20010 7710 20015 7730
rect 19985 7680 20015 7710
rect 19985 7660 19990 7680
rect 20010 7660 20015 7680
rect 19985 7630 20015 7660
rect 19985 7610 19990 7630
rect 20010 7610 20015 7630
rect 19985 7580 20015 7610
rect 19985 7560 19990 7580
rect 20010 7560 20015 7580
rect 19985 7530 20015 7560
rect 19985 7510 19990 7530
rect 20010 7510 20015 7530
rect 19985 7500 20015 7510
rect 20045 7880 20115 7890
rect 20350 7885 20390 7895
rect 20500 7915 20540 7925
rect 20500 7895 20510 7915
rect 20530 7895 20540 7915
rect 20500 7885 20540 7895
rect 20558 7915 20592 7925
rect 20558 7895 20566 7915
rect 20584 7895 20592 7915
rect 20558 7885 20592 7895
rect 20610 7915 20650 7925
rect 20610 7895 20620 7915
rect 20640 7895 20650 7915
rect 20610 7885 20650 7895
rect 20720 7915 20760 7925
rect 20720 7895 20730 7915
rect 20750 7895 20760 7915
rect 20720 7885 20760 7895
rect 20830 7915 20870 7925
rect 20830 7895 20840 7915
rect 20860 7895 20870 7915
rect 20830 7885 20870 7895
rect 20940 7915 20980 7925
rect 20940 7895 20950 7915
rect 20970 7895 20980 7915
rect 20940 7885 20980 7895
rect 21050 7915 21090 7925
rect 21050 7895 21060 7915
rect 21080 7895 21090 7915
rect 21050 7885 21090 7895
rect 21160 7915 21200 7925
rect 21160 7895 21170 7915
rect 21190 7895 21200 7915
rect 21160 7885 21200 7895
rect 21270 7915 21310 7925
rect 21270 7895 21280 7915
rect 21300 7895 21310 7915
rect 21270 7885 21310 7895
rect 21380 7915 21420 7925
rect 21380 7895 21390 7915
rect 21410 7895 21420 7915
rect 21380 7885 21420 7895
rect 21490 7915 21530 7925
rect 21490 7895 21500 7915
rect 21520 7895 21530 7915
rect 21490 7885 21530 7895
rect 21640 7915 21680 7925
rect 21640 7895 21650 7915
rect 21670 7895 21680 7915
rect 21640 7885 21680 7895
rect 20045 7860 20050 7880
rect 20070 7860 20090 7880
rect 20110 7860 20115 7880
rect 20045 7830 20115 7860
rect 20045 7810 20050 7830
rect 20070 7810 20090 7830
rect 20110 7810 20115 7830
rect 20045 7780 20115 7810
rect 20045 7760 20050 7780
rect 20070 7760 20090 7780
rect 20110 7760 20115 7780
rect 20045 7730 20115 7760
rect 20045 7710 20050 7730
rect 20070 7710 20090 7730
rect 20110 7710 20115 7730
rect 20045 7680 20115 7710
rect 20555 7695 20595 7836
rect 20045 7660 20050 7680
rect 20070 7660 20090 7680
rect 20110 7660 20115 7680
rect 20045 7630 20115 7660
rect 20445 7665 20485 7675
rect 20445 7645 20455 7665
rect 20475 7645 20485 7665
rect 20445 7635 20485 7645
rect 20555 7665 20595 7675
rect 20555 7645 20565 7665
rect 20585 7645 20595 7665
rect 20555 7635 20595 7645
rect 20665 7665 20705 7675
rect 20665 7645 20675 7665
rect 20695 7645 20705 7665
rect 20665 7635 20705 7645
rect 20775 7665 20815 7675
rect 20775 7645 20785 7665
rect 20805 7645 20815 7665
rect 20775 7635 20815 7645
rect 20885 7665 20925 7675
rect 20885 7645 20895 7665
rect 20915 7645 20925 7665
rect 20885 7635 20925 7645
rect 20995 7665 21035 7675
rect 20995 7645 21005 7665
rect 21025 7645 21035 7665
rect 20995 7635 21035 7645
rect 21105 7665 21145 7675
rect 21105 7645 21115 7665
rect 21135 7645 21145 7665
rect 21105 7635 21145 7645
rect 21215 7665 21255 7675
rect 21215 7645 21225 7665
rect 21245 7645 21255 7665
rect 21215 7635 21255 7645
rect 21325 7665 21365 7675
rect 21325 7645 21335 7665
rect 21355 7645 21365 7665
rect 21325 7635 21365 7645
rect 21435 7665 21475 7675
rect 21435 7645 21445 7665
rect 21465 7645 21475 7665
rect 21435 7635 21475 7645
rect 21545 7665 21585 7675
rect 21545 7645 21555 7665
rect 21575 7645 21585 7665
rect 21545 7635 21585 7645
rect 20045 7610 20050 7630
rect 20070 7610 20090 7630
rect 20110 7610 20115 7630
rect 20455 7615 20475 7635
rect 20565 7615 20585 7635
rect 20675 7615 20695 7635
rect 20785 7615 20805 7635
rect 20895 7615 20915 7635
rect 21005 7615 21025 7635
rect 21115 7615 21135 7635
rect 21225 7615 21245 7635
rect 21335 7615 21355 7635
rect 21445 7615 21465 7635
rect 21555 7615 21575 7635
rect 20045 7580 20115 7610
rect 20045 7560 20050 7580
rect 20070 7560 20090 7580
rect 20110 7560 20115 7580
rect 20045 7530 20115 7560
rect 20045 7510 20050 7530
rect 20070 7510 20090 7530
rect 20110 7510 20115 7530
rect 20355 7605 20425 7615
rect 20355 7585 20360 7605
rect 20380 7585 20400 7605
rect 20420 7585 20425 7605
rect 20355 7555 20425 7585
rect 20355 7535 20360 7555
rect 20380 7535 20400 7555
rect 20420 7535 20425 7555
rect 20355 7525 20425 7535
rect 20450 7605 20480 7615
rect 20450 7585 20455 7605
rect 20475 7585 20480 7605
rect 20450 7555 20480 7585
rect 20450 7535 20455 7555
rect 20475 7535 20480 7555
rect 20450 7525 20480 7535
rect 20505 7605 20535 7615
rect 20505 7585 20510 7605
rect 20530 7585 20535 7605
rect 20505 7555 20535 7585
rect 20505 7535 20510 7555
rect 20530 7535 20535 7555
rect 20505 7525 20535 7535
rect 20560 7605 20590 7615
rect 20560 7585 20565 7605
rect 20585 7585 20590 7605
rect 20560 7555 20590 7585
rect 20560 7535 20565 7555
rect 20585 7535 20590 7555
rect 20560 7525 20590 7535
rect 20615 7605 20645 7615
rect 20615 7585 20620 7605
rect 20640 7585 20645 7605
rect 20615 7555 20645 7585
rect 20615 7535 20620 7555
rect 20640 7535 20645 7555
rect 20615 7525 20645 7535
rect 20670 7605 20700 7615
rect 20670 7585 20675 7605
rect 20695 7585 20700 7605
rect 20670 7555 20700 7585
rect 20670 7535 20675 7555
rect 20695 7535 20700 7555
rect 20670 7525 20700 7535
rect 20725 7605 20755 7615
rect 20725 7585 20730 7605
rect 20750 7585 20755 7605
rect 20725 7555 20755 7585
rect 20725 7535 20730 7555
rect 20750 7535 20755 7555
rect 20725 7525 20755 7535
rect 20780 7605 20810 7615
rect 20780 7585 20785 7605
rect 20805 7585 20810 7605
rect 20780 7555 20810 7585
rect 20780 7535 20785 7555
rect 20805 7535 20810 7555
rect 20780 7525 20810 7535
rect 20835 7605 20865 7615
rect 20835 7585 20840 7605
rect 20860 7585 20865 7605
rect 20835 7555 20865 7585
rect 20835 7535 20840 7555
rect 20860 7535 20865 7555
rect 20835 7525 20865 7535
rect 20890 7605 20920 7615
rect 20890 7585 20895 7605
rect 20915 7585 20920 7605
rect 20890 7555 20920 7585
rect 20890 7535 20895 7555
rect 20915 7535 20920 7555
rect 20890 7525 20920 7535
rect 20945 7605 20975 7615
rect 20945 7585 20950 7605
rect 20970 7585 20975 7605
rect 20945 7555 20975 7585
rect 20945 7535 20950 7555
rect 20970 7535 20975 7555
rect 20945 7525 20975 7535
rect 21000 7605 21030 7615
rect 21000 7585 21005 7605
rect 21025 7585 21030 7605
rect 21000 7555 21030 7585
rect 21000 7535 21005 7555
rect 21025 7535 21030 7555
rect 21000 7525 21030 7535
rect 21055 7605 21085 7615
rect 21055 7585 21060 7605
rect 21080 7585 21085 7605
rect 21055 7555 21085 7585
rect 21055 7535 21060 7555
rect 21080 7535 21085 7555
rect 21055 7525 21085 7535
rect 21110 7605 21140 7615
rect 21110 7585 21115 7605
rect 21135 7585 21140 7605
rect 21110 7555 21140 7585
rect 21110 7535 21115 7555
rect 21135 7535 21140 7555
rect 21110 7525 21140 7535
rect 21165 7605 21195 7615
rect 21165 7585 21170 7605
rect 21190 7585 21195 7605
rect 21165 7555 21195 7585
rect 21165 7535 21170 7555
rect 21190 7535 21195 7555
rect 21165 7525 21195 7535
rect 21220 7605 21250 7615
rect 21220 7585 21225 7605
rect 21245 7585 21250 7605
rect 21220 7555 21250 7585
rect 21220 7535 21225 7555
rect 21245 7535 21250 7555
rect 21220 7525 21250 7535
rect 21275 7605 21305 7615
rect 21275 7585 21280 7605
rect 21300 7585 21305 7605
rect 21275 7555 21305 7585
rect 21275 7535 21280 7555
rect 21300 7535 21305 7555
rect 21275 7525 21305 7535
rect 21330 7605 21360 7615
rect 21330 7585 21335 7605
rect 21355 7585 21360 7605
rect 21330 7555 21360 7585
rect 21330 7535 21335 7555
rect 21355 7535 21360 7555
rect 21330 7525 21360 7535
rect 21385 7605 21415 7615
rect 21385 7585 21390 7605
rect 21410 7585 21415 7605
rect 21385 7555 21415 7585
rect 21385 7535 21390 7555
rect 21410 7535 21415 7555
rect 21385 7525 21415 7535
rect 21440 7605 21470 7615
rect 21440 7585 21445 7605
rect 21465 7585 21470 7605
rect 21440 7555 21470 7585
rect 21440 7535 21445 7555
rect 21465 7535 21470 7555
rect 21440 7525 21470 7535
rect 21495 7605 21525 7615
rect 21495 7585 21500 7605
rect 21520 7585 21525 7605
rect 21495 7555 21525 7585
rect 21495 7535 21500 7555
rect 21520 7535 21525 7555
rect 21495 7525 21525 7535
rect 21550 7605 21580 7615
rect 21550 7585 21555 7605
rect 21575 7585 21580 7605
rect 21550 7555 21580 7585
rect 21550 7535 21555 7555
rect 21575 7535 21580 7555
rect 21550 7525 21580 7535
rect 21605 7605 21675 7615
rect 21605 7585 21610 7605
rect 21630 7585 21650 7605
rect 21670 7585 21675 7605
rect 21605 7555 21675 7585
rect 21605 7535 21610 7555
rect 21630 7535 21650 7555
rect 21670 7535 21675 7555
rect 21605 7525 21675 7535
rect 20045 7500 20115 7510
rect 20360 7505 20380 7525
rect 20510 7505 20530 7525
rect 20620 7505 20640 7525
rect 20730 7505 20750 7525
rect 20840 7505 20860 7525
rect 20950 7505 20970 7525
rect 21060 7505 21080 7525
rect 21170 7505 21190 7525
rect 21280 7505 21300 7525
rect 21390 7505 21410 7525
rect 21500 7505 21520 7525
rect 21650 7505 21670 7525
rect 18430 7475 18440 7495
rect 18460 7475 18470 7495
rect 18790 7480 18810 7500
rect 18910 7480 18930 7500
rect 19030 7480 19050 7500
rect 19150 7480 19170 7500
rect 19270 7480 19290 7500
rect 19390 7480 19410 7500
rect 19510 7480 19530 7500
rect 19630 7480 19650 7500
rect 19750 7480 19770 7500
rect 19870 7480 19890 7500
rect 19990 7480 20010 7500
rect 20350 7495 20390 7505
rect 18430 7465 18470 7475
rect 18780 7470 18820 7480
rect 12480 7440 12520 7450
rect 18780 7450 18790 7470
rect 18810 7450 18820 7470
rect 10813 7415 10821 7435
rect 10839 7415 10847 7435
rect 10813 7405 10847 7415
rect 12978 7435 13012 7445
rect 12978 7415 12986 7435
rect 13004 7415 13012 7435
rect 12978 7405 13012 7415
rect 18313 7435 18347 7445
rect 18780 7440 18820 7450
rect 18900 7470 18940 7480
rect 18900 7450 18910 7470
rect 18930 7450 18940 7470
rect 18900 7440 18940 7450
rect 19020 7470 19060 7480
rect 19020 7450 19030 7470
rect 19050 7450 19060 7470
rect 19020 7440 19060 7450
rect 19140 7470 19180 7480
rect 19140 7450 19150 7470
rect 19170 7450 19180 7470
rect 19140 7440 19180 7450
rect 19260 7470 19300 7480
rect 19260 7450 19270 7470
rect 19290 7450 19300 7470
rect 19260 7440 19300 7450
rect 19323 7470 19357 7480
rect 19323 7450 19331 7470
rect 19349 7450 19357 7470
rect 19323 7440 19357 7450
rect 19380 7470 19420 7480
rect 19380 7450 19390 7470
rect 19410 7450 19420 7470
rect 19380 7440 19420 7450
rect 19500 7470 19540 7480
rect 19500 7450 19510 7470
rect 19530 7450 19540 7470
rect 19500 7440 19540 7450
rect 19620 7470 19660 7480
rect 19620 7450 19630 7470
rect 19650 7450 19660 7470
rect 19620 7440 19660 7450
rect 19740 7470 19780 7480
rect 19740 7450 19750 7470
rect 19770 7450 19780 7470
rect 19740 7440 19780 7450
rect 19860 7470 19900 7480
rect 19860 7450 19870 7470
rect 19890 7450 19900 7470
rect 19860 7440 19900 7450
rect 19980 7470 20020 7480
rect 19980 7450 19990 7470
rect 20010 7450 20020 7470
rect 20350 7475 20360 7495
rect 20380 7475 20390 7495
rect 20350 7465 20390 7475
rect 20500 7495 20540 7505
rect 20500 7475 20510 7495
rect 20530 7475 20540 7495
rect 20500 7465 20540 7475
rect 20610 7495 20650 7505
rect 20610 7475 20620 7495
rect 20640 7475 20650 7495
rect 20610 7465 20650 7475
rect 20720 7495 20760 7505
rect 20720 7475 20730 7495
rect 20750 7475 20760 7495
rect 20720 7465 20760 7475
rect 20830 7495 20870 7505
rect 20830 7475 20840 7495
rect 20860 7475 20870 7495
rect 20830 7465 20870 7475
rect 20940 7495 20980 7505
rect 20940 7475 20950 7495
rect 20970 7475 20980 7495
rect 20940 7465 20980 7475
rect 21050 7495 21090 7505
rect 21050 7475 21060 7495
rect 21080 7475 21090 7495
rect 21050 7465 21090 7475
rect 21160 7495 21200 7505
rect 21160 7475 21170 7495
rect 21190 7475 21200 7495
rect 21160 7465 21200 7475
rect 21270 7495 21310 7505
rect 21270 7475 21280 7495
rect 21300 7475 21310 7495
rect 21270 7465 21310 7475
rect 21380 7495 21420 7505
rect 21380 7475 21390 7495
rect 21410 7475 21420 7495
rect 21380 7465 21420 7475
rect 21490 7495 21530 7505
rect 21490 7475 21500 7495
rect 21520 7475 21530 7495
rect 21490 7465 21530 7475
rect 21640 7495 21680 7505
rect 21640 7475 21650 7495
rect 21670 7475 21680 7495
rect 21640 7465 21680 7475
rect 19980 7440 20020 7450
rect 18313 7415 18321 7435
rect 18339 7415 18347 7435
rect 18313 7405 18347 7415
rect 20473 7435 20507 7445
rect 20473 7415 20481 7435
rect 20499 7415 20507 7435
rect 20473 7405 20507 7415
rect 9800 7375 9845 7380
rect 9800 7350 9810 7375
rect 9835 7350 9845 7375
rect 9800 7345 9845 7350
rect 10635 7375 10680 7380
rect 10635 7350 10645 7375
rect 10670 7350 10680 7375
rect 10635 7345 10680 7350
rect 13145 7375 13190 7380
rect 13145 7350 13155 7375
rect 13180 7350 13190 7375
rect 13145 7345 13190 7350
rect 13980 7375 14025 7380
rect 13980 7350 13990 7375
rect 14015 7350 14025 7375
rect 13980 7345 14025 7350
rect 17300 7375 17345 7380
rect 17300 7350 17310 7375
rect 17335 7350 17345 7375
rect 17300 7345 17345 7350
rect 18135 7375 18180 7380
rect 18135 7350 18145 7375
rect 18170 7350 18180 7375
rect 18135 7345 18180 7350
rect 20640 7375 20685 7380
rect 20640 7350 20650 7375
rect 20675 7350 20685 7375
rect 20640 7345 20685 7350
rect 21475 7375 21520 7380
rect 21475 7350 21485 7375
rect 21510 7350 21520 7375
rect 21475 7345 21520 7350
rect 9800 7315 9845 7320
rect 9800 7290 9810 7315
rect 9835 7290 9845 7315
rect 9800 7285 9845 7290
rect 10635 7315 10680 7320
rect 10635 7290 10645 7315
rect 10670 7290 10680 7315
rect 10635 7285 10680 7290
rect 13145 7315 13190 7320
rect 13145 7290 13155 7315
rect 13180 7290 13190 7315
rect 13145 7285 13190 7290
rect 13980 7315 14025 7320
rect 13980 7290 13990 7315
rect 14015 7290 14025 7315
rect 13980 7285 14025 7290
rect 17300 7315 17345 7320
rect 17300 7290 17310 7315
rect 17335 7290 17345 7315
rect 17300 7285 17345 7290
rect 18135 7315 18180 7320
rect 18135 7290 18145 7315
rect 18170 7290 18180 7315
rect 18135 7285 18180 7290
rect 20640 7315 20685 7320
rect 20640 7290 20650 7315
rect 20675 7290 20685 7315
rect 20640 7285 20685 7290
rect 21475 7315 21520 7320
rect 21475 7290 21485 7315
rect 21510 7290 21520 7315
rect 21475 7285 21520 7290
rect 10813 7275 10847 7285
rect 10813 7255 10821 7275
rect 10839 7255 10847 7275
rect 10813 7245 10847 7255
rect 12978 7275 13012 7285
rect 12978 7255 12986 7275
rect 13004 7255 13012 7275
rect 12978 7245 13012 7255
rect 18313 7275 18347 7285
rect 18313 7255 18321 7275
rect 18339 7255 18347 7275
rect 18313 7245 18347 7255
rect 20473 7275 20507 7285
rect 20473 7255 20481 7275
rect 20499 7255 20507 7275
rect 20473 7245 20507 7255
rect 9640 7215 9680 7225
rect 9640 7195 9650 7215
rect 9670 7195 9680 7215
rect 9640 7185 9680 7195
rect 9790 7215 9830 7225
rect 9790 7195 9800 7215
rect 9820 7195 9830 7215
rect 9790 7185 9830 7195
rect 9900 7215 9940 7225
rect 9900 7195 9910 7215
rect 9930 7195 9940 7215
rect 9900 7185 9940 7195
rect 10010 7215 10050 7225
rect 10010 7195 10020 7215
rect 10040 7195 10050 7215
rect 10010 7185 10050 7195
rect 10120 7215 10160 7225
rect 10120 7195 10130 7215
rect 10150 7195 10160 7215
rect 10120 7185 10160 7195
rect 10230 7215 10270 7225
rect 10230 7195 10240 7215
rect 10260 7195 10270 7215
rect 10230 7185 10270 7195
rect 10340 7215 10380 7225
rect 10340 7195 10350 7215
rect 10370 7195 10380 7215
rect 10340 7185 10380 7195
rect 10450 7215 10490 7225
rect 10450 7195 10460 7215
rect 10480 7195 10490 7215
rect 10450 7185 10490 7195
rect 10560 7215 10600 7225
rect 10560 7195 10570 7215
rect 10590 7195 10600 7215
rect 10560 7185 10600 7195
rect 10670 7215 10710 7225
rect 10670 7195 10680 7215
rect 10700 7195 10710 7215
rect 10670 7185 10710 7195
rect 10780 7215 10820 7225
rect 10780 7195 10790 7215
rect 10810 7195 10820 7215
rect 10780 7185 10820 7195
rect 10930 7215 10970 7225
rect 10930 7195 10940 7215
rect 10960 7195 10970 7215
rect 10930 7185 10970 7195
rect 12855 7215 12895 7225
rect 12855 7195 12865 7215
rect 12885 7195 12895 7215
rect 12855 7185 12895 7195
rect 13005 7215 13045 7225
rect 13005 7195 13015 7215
rect 13035 7195 13045 7215
rect 13005 7185 13045 7195
rect 13115 7215 13155 7225
rect 13115 7195 13125 7215
rect 13145 7195 13155 7215
rect 13115 7185 13155 7195
rect 13225 7215 13265 7225
rect 13225 7195 13235 7215
rect 13255 7195 13265 7215
rect 13225 7185 13265 7195
rect 13335 7215 13375 7225
rect 13335 7195 13345 7215
rect 13365 7195 13375 7215
rect 13335 7185 13375 7195
rect 13445 7215 13485 7225
rect 13445 7195 13455 7215
rect 13475 7195 13485 7215
rect 13445 7185 13485 7195
rect 13555 7215 13595 7225
rect 13555 7195 13565 7215
rect 13585 7195 13595 7215
rect 13555 7185 13595 7195
rect 13665 7215 13705 7225
rect 13665 7195 13675 7215
rect 13695 7195 13705 7215
rect 13665 7185 13705 7195
rect 13775 7215 13815 7225
rect 13775 7195 13785 7215
rect 13805 7195 13815 7215
rect 13775 7185 13815 7195
rect 13885 7215 13925 7225
rect 13885 7195 13895 7215
rect 13915 7195 13925 7215
rect 13885 7185 13925 7195
rect 13995 7215 14035 7225
rect 13995 7195 14005 7215
rect 14025 7195 14035 7215
rect 13995 7185 14035 7195
rect 14145 7215 14185 7225
rect 14145 7195 14155 7215
rect 14175 7195 14185 7215
rect 14145 7185 14185 7195
rect 17140 7215 17180 7225
rect 17140 7195 17150 7215
rect 17170 7195 17180 7215
rect 17140 7185 17180 7195
rect 17290 7215 17330 7225
rect 17290 7195 17300 7215
rect 17320 7195 17330 7215
rect 17290 7185 17330 7195
rect 17400 7215 17440 7225
rect 17400 7195 17410 7215
rect 17430 7195 17440 7215
rect 17400 7185 17440 7195
rect 17510 7215 17550 7225
rect 17510 7195 17520 7215
rect 17540 7195 17550 7215
rect 17510 7185 17550 7195
rect 17620 7215 17660 7225
rect 17620 7195 17630 7215
rect 17650 7195 17660 7215
rect 17620 7185 17660 7195
rect 17730 7215 17770 7225
rect 17730 7195 17740 7215
rect 17760 7195 17770 7215
rect 17730 7185 17770 7195
rect 17840 7215 17880 7225
rect 17840 7195 17850 7215
rect 17870 7195 17880 7215
rect 17840 7185 17880 7195
rect 17950 7215 17990 7225
rect 17950 7195 17960 7215
rect 17980 7195 17990 7215
rect 17950 7185 17990 7195
rect 18060 7215 18100 7225
rect 18060 7195 18070 7215
rect 18090 7195 18100 7215
rect 18060 7185 18100 7195
rect 18170 7215 18210 7225
rect 18170 7195 18180 7215
rect 18200 7195 18210 7215
rect 18170 7185 18210 7195
rect 18280 7215 18320 7225
rect 18280 7195 18290 7215
rect 18310 7195 18320 7215
rect 18280 7185 18320 7195
rect 18430 7215 18470 7225
rect 18430 7195 18440 7215
rect 18460 7195 18470 7215
rect 18430 7185 18470 7195
rect 20350 7215 20390 7225
rect 20350 7195 20360 7215
rect 20380 7195 20390 7215
rect 20350 7185 20390 7195
rect 20500 7215 20540 7225
rect 20500 7195 20510 7215
rect 20530 7195 20540 7215
rect 20500 7185 20540 7195
rect 20610 7215 20650 7225
rect 20610 7195 20620 7215
rect 20640 7195 20650 7215
rect 20610 7185 20650 7195
rect 20720 7215 20760 7225
rect 20720 7195 20730 7215
rect 20750 7195 20760 7215
rect 20720 7185 20760 7195
rect 20830 7215 20870 7225
rect 20830 7195 20840 7215
rect 20860 7195 20870 7215
rect 20830 7185 20870 7195
rect 20940 7215 20980 7225
rect 20940 7195 20950 7215
rect 20970 7195 20980 7215
rect 20940 7185 20980 7195
rect 21050 7215 21090 7225
rect 21050 7195 21060 7215
rect 21080 7195 21090 7215
rect 21050 7185 21090 7195
rect 21160 7215 21200 7225
rect 21160 7195 21170 7215
rect 21190 7195 21200 7215
rect 21160 7185 21200 7195
rect 21270 7215 21310 7225
rect 21270 7195 21280 7215
rect 21300 7195 21310 7215
rect 21270 7185 21310 7195
rect 21380 7215 21420 7225
rect 21380 7195 21390 7215
rect 21410 7195 21420 7215
rect 21380 7185 21420 7195
rect 21490 7215 21530 7225
rect 21490 7195 21500 7215
rect 21520 7195 21530 7215
rect 21490 7185 21530 7195
rect 21640 7215 21680 7225
rect 21640 7195 21650 7215
rect 21670 7195 21680 7215
rect 21640 7185 21680 7195
rect 9650 7165 9670 7185
rect 9800 7165 9820 7185
rect 9910 7165 9930 7185
rect 10020 7165 10040 7185
rect 10130 7165 10150 7185
rect 10240 7165 10260 7185
rect 10350 7165 10370 7185
rect 10460 7165 10480 7185
rect 10570 7165 10590 7185
rect 10680 7165 10700 7185
rect 10790 7165 10810 7185
rect 10940 7165 10960 7185
rect 11330 7175 11370 7185
rect 9645 7155 9715 7165
rect 9645 7135 9650 7155
rect 9670 7135 9690 7155
rect 9710 7135 9715 7155
rect 9645 7105 9715 7135
rect 9645 7085 9650 7105
rect 9670 7085 9690 7105
rect 9710 7085 9715 7105
rect 9645 7055 9715 7085
rect 9645 7035 9650 7055
rect 9670 7035 9690 7055
rect 9710 7035 9715 7055
rect 9645 7025 9715 7035
rect 9740 7155 9770 7165
rect 9740 7135 9745 7155
rect 9765 7135 9770 7155
rect 9740 7105 9770 7135
rect 9740 7085 9745 7105
rect 9765 7085 9770 7105
rect 9740 7055 9770 7085
rect 9740 7035 9745 7055
rect 9765 7035 9770 7055
rect 9740 7025 9770 7035
rect 9795 7155 9825 7165
rect 9795 7135 9800 7155
rect 9820 7135 9825 7155
rect 9795 7105 9825 7135
rect 9795 7085 9800 7105
rect 9820 7085 9825 7105
rect 9795 7055 9825 7085
rect 9795 7035 9800 7055
rect 9820 7035 9825 7055
rect 9795 7025 9825 7035
rect 9850 7155 9880 7165
rect 9850 7135 9855 7155
rect 9875 7135 9880 7155
rect 9850 7105 9880 7135
rect 9850 7085 9855 7105
rect 9875 7085 9880 7105
rect 9850 7055 9880 7085
rect 9850 7035 9855 7055
rect 9875 7035 9880 7055
rect 9850 7025 9880 7035
rect 9905 7155 9935 7165
rect 9905 7135 9910 7155
rect 9930 7135 9935 7155
rect 9905 7105 9935 7135
rect 9905 7085 9910 7105
rect 9930 7085 9935 7105
rect 9905 7055 9935 7085
rect 9905 7035 9910 7055
rect 9930 7035 9935 7055
rect 9905 7025 9935 7035
rect 9960 7155 9990 7165
rect 9960 7135 9965 7155
rect 9985 7135 9990 7155
rect 9960 7105 9990 7135
rect 9960 7085 9965 7105
rect 9985 7085 9990 7105
rect 9960 7055 9990 7085
rect 9960 7035 9965 7055
rect 9985 7035 9990 7055
rect 9960 7025 9990 7035
rect 10015 7155 10045 7165
rect 10015 7135 10020 7155
rect 10040 7135 10045 7155
rect 10015 7105 10045 7135
rect 10015 7085 10020 7105
rect 10040 7085 10045 7105
rect 10015 7055 10045 7085
rect 10015 7035 10020 7055
rect 10040 7035 10045 7055
rect 10015 7025 10045 7035
rect 10070 7155 10100 7165
rect 10070 7135 10075 7155
rect 10095 7135 10100 7155
rect 10070 7105 10100 7135
rect 10070 7085 10075 7105
rect 10095 7085 10100 7105
rect 10070 7055 10100 7085
rect 10070 7035 10075 7055
rect 10095 7035 10100 7055
rect 10070 7025 10100 7035
rect 10125 7155 10155 7165
rect 10125 7135 10130 7155
rect 10150 7135 10155 7155
rect 10125 7105 10155 7135
rect 10125 7085 10130 7105
rect 10150 7085 10155 7105
rect 10125 7055 10155 7085
rect 10125 7035 10130 7055
rect 10150 7035 10155 7055
rect 10125 7025 10155 7035
rect 10180 7155 10210 7165
rect 10180 7135 10185 7155
rect 10205 7135 10210 7155
rect 10180 7105 10210 7135
rect 10180 7085 10185 7105
rect 10205 7085 10210 7105
rect 10180 7055 10210 7085
rect 10180 7035 10185 7055
rect 10205 7035 10210 7055
rect 10180 7025 10210 7035
rect 10235 7155 10265 7165
rect 10235 7135 10240 7155
rect 10260 7135 10265 7155
rect 10235 7105 10265 7135
rect 10235 7085 10240 7105
rect 10260 7085 10265 7105
rect 10235 7055 10265 7085
rect 10235 7035 10240 7055
rect 10260 7035 10265 7055
rect 10235 7025 10265 7035
rect 10290 7155 10320 7165
rect 10290 7135 10295 7155
rect 10315 7135 10320 7155
rect 10290 7105 10320 7135
rect 10290 7085 10295 7105
rect 10315 7085 10320 7105
rect 10290 7055 10320 7085
rect 10290 7035 10295 7055
rect 10315 7035 10320 7055
rect 10290 7025 10320 7035
rect 10345 7155 10375 7165
rect 10345 7135 10350 7155
rect 10370 7135 10375 7155
rect 10345 7105 10375 7135
rect 10345 7085 10350 7105
rect 10370 7085 10375 7105
rect 10345 7055 10375 7085
rect 10345 7035 10350 7055
rect 10370 7035 10375 7055
rect 10345 7025 10375 7035
rect 10400 7155 10430 7165
rect 10400 7135 10405 7155
rect 10425 7135 10430 7155
rect 10400 7105 10430 7135
rect 10400 7085 10405 7105
rect 10425 7085 10430 7105
rect 10400 7055 10430 7085
rect 10400 7035 10405 7055
rect 10425 7035 10430 7055
rect 10400 7025 10430 7035
rect 10455 7155 10485 7165
rect 10455 7135 10460 7155
rect 10480 7135 10485 7155
rect 10455 7105 10485 7135
rect 10455 7085 10460 7105
rect 10480 7085 10485 7105
rect 10455 7055 10485 7085
rect 10455 7035 10460 7055
rect 10480 7035 10485 7055
rect 10455 7025 10485 7035
rect 10510 7155 10540 7165
rect 10510 7135 10515 7155
rect 10535 7135 10540 7155
rect 10510 7105 10540 7135
rect 10510 7085 10515 7105
rect 10535 7085 10540 7105
rect 10510 7055 10540 7085
rect 10510 7035 10515 7055
rect 10535 7035 10540 7055
rect 10510 7025 10540 7035
rect 10565 7155 10595 7165
rect 10565 7135 10570 7155
rect 10590 7135 10595 7155
rect 10565 7105 10595 7135
rect 10565 7085 10570 7105
rect 10590 7085 10595 7105
rect 10565 7055 10595 7085
rect 10565 7035 10570 7055
rect 10590 7035 10595 7055
rect 10565 7025 10595 7035
rect 10620 7155 10650 7165
rect 10620 7135 10625 7155
rect 10645 7135 10650 7155
rect 10620 7105 10650 7135
rect 10620 7085 10625 7105
rect 10645 7085 10650 7105
rect 10620 7055 10650 7085
rect 10620 7035 10625 7055
rect 10645 7035 10650 7055
rect 10620 7025 10650 7035
rect 10675 7155 10705 7165
rect 10675 7135 10680 7155
rect 10700 7135 10705 7155
rect 10675 7105 10705 7135
rect 10675 7085 10680 7105
rect 10700 7085 10705 7105
rect 10675 7055 10705 7085
rect 10675 7035 10680 7055
rect 10700 7035 10705 7055
rect 10675 7025 10705 7035
rect 10730 7155 10760 7165
rect 10730 7135 10735 7155
rect 10755 7135 10760 7155
rect 10730 7105 10760 7135
rect 10730 7085 10735 7105
rect 10755 7085 10760 7105
rect 10730 7055 10760 7085
rect 10730 7035 10735 7055
rect 10755 7035 10760 7055
rect 10730 7025 10760 7035
rect 10785 7155 10815 7165
rect 10785 7135 10790 7155
rect 10810 7135 10815 7155
rect 10785 7105 10815 7135
rect 10785 7085 10790 7105
rect 10810 7085 10815 7105
rect 10785 7055 10815 7085
rect 10785 7035 10790 7055
rect 10810 7035 10815 7055
rect 10785 7025 10815 7035
rect 10840 7155 10870 7165
rect 10840 7135 10845 7155
rect 10865 7135 10870 7155
rect 10840 7105 10870 7135
rect 10840 7085 10845 7105
rect 10865 7085 10870 7105
rect 10840 7055 10870 7085
rect 10840 7035 10845 7055
rect 10865 7035 10870 7055
rect 10840 7025 10870 7035
rect 10895 7155 10965 7165
rect 10895 7135 10900 7155
rect 10920 7135 10940 7155
rect 10960 7135 10965 7155
rect 11330 7155 11340 7175
rect 11360 7155 11370 7175
rect 11330 7145 11370 7155
rect 11440 7175 11480 7185
rect 11440 7155 11450 7175
rect 11470 7155 11480 7175
rect 11440 7145 11480 7155
rect 11550 7175 11590 7185
rect 11550 7155 11560 7175
rect 11580 7155 11590 7175
rect 11550 7145 11590 7155
rect 11660 7175 11700 7185
rect 11660 7155 11670 7175
rect 11690 7155 11700 7175
rect 11660 7145 11700 7155
rect 11770 7175 11810 7185
rect 11770 7155 11780 7175
rect 11800 7155 11810 7175
rect 11770 7145 11810 7155
rect 11880 7175 11920 7185
rect 11880 7155 11890 7175
rect 11910 7155 11920 7175
rect 11880 7145 11920 7155
rect 11990 7175 12030 7185
rect 11990 7155 12000 7175
rect 12020 7155 12030 7175
rect 11990 7145 12030 7155
rect 12100 7175 12140 7185
rect 12100 7155 12110 7175
rect 12130 7155 12140 7175
rect 12100 7145 12140 7155
rect 12210 7175 12250 7185
rect 12210 7155 12220 7175
rect 12240 7155 12250 7175
rect 12210 7145 12250 7155
rect 12320 7175 12360 7185
rect 12320 7155 12330 7175
rect 12350 7155 12360 7175
rect 12320 7145 12360 7155
rect 12430 7175 12470 7185
rect 12430 7155 12440 7175
rect 12460 7155 12470 7175
rect 12865 7165 12885 7185
rect 13015 7165 13035 7185
rect 13125 7165 13145 7185
rect 13235 7165 13255 7185
rect 13345 7165 13365 7185
rect 13455 7165 13475 7185
rect 13565 7165 13585 7185
rect 13675 7165 13695 7185
rect 13785 7165 13805 7185
rect 13895 7165 13915 7185
rect 14005 7165 14025 7185
rect 14155 7165 14175 7185
rect 17150 7165 17170 7185
rect 17300 7165 17320 7185
rect 17410 7165 17430 7185
rect 17520 7165 17540 7185
rect 17630 7165 17650 7185
rect 17740 7165 17760 7185
rect 17850 7165 17870 7185
rect 17960 7165 17980 7185
rect 18070 7165 18090 7185
rect 18180 7165 18200 7185
rect 18290 7165 18310 7185
rect 18440 7165 18460 7185
rect 18830 7175 18870 7185
rect 12430 7145 12470 7155
rect 12860 7155 12930 7165
rect 10895 7105 10965 7135
rect 11340 7125 11360 7145
rect 11450 7125 11470 7145
rect 11560 7125 11580 7145
rect 11670 7125 11690 7145
rect 11780 7125 11800 7145
rect 11890 7125 11910 7145
rect 12000 7125 12020 7145
rect 12110 7125 12130 7145
rect 12220 7125 12240 7145
rect 12330 7125 12350 7145
rect 12440 7125 12460 7145
rect 12860 7135 12865 7155
rect 12885 7135 12905 7155
rect 12925 7135 12930 7155
rect 10895 7085 10900 7105
rect 10920 7085 10940 7105
rect 10960 7085 10965 7105
rect 10895 7055 10965 7085
rect 10895 7035 10900 7055
rect 10920 7035 10940 7055
rect 10960 7035 10965 7055
rect 10895 7025 10965 7035
rect 11240 7115 11310 7125
rect 11240 7095 11245 7115
rect 11265 7095 11285 7115
rect 11305 7095 11310 7115
rect 11240 7065 11310 7095
rect 11240 7045 11245 7065
rect 11265 7045 11285 7065
rect 11305 7045 11310 7065
rect 9745 7005 9765 7025
rect 9855 7005 9875 7025
rect 9965 7005 9985 7025
rect 10075 7005 10095 7025
rect 10185 7005 10205 7025
rect 10295 7005 10315 7025
rect 10405 7005 10425 7025
rect 10515 7005 10535 7025
rect 10625 7005 10645 7025
rect 10735 7005 10755 7025
rect 10845 7005 10865 7025
rect 11240 7015 11310 7045
rect 9735 6995 9775 7005
rect 9735 6975 9745 6995
rect 9763 6975 9775 6995
rect 9735 6965 9775 6975
rect 9845 6995 9885 7005
rect 9845 6975 9855 6995
rect 9873 6975 9885 6995
rect 9845 6965 9885 6975
rect 9955 6995 9995 7005
rect 9955 6975 9965 6995
rect 9983 6975 9995 6995
rect 9955 6965 9995 6975
rect 10065 6995 10105 7005
rect 10065 6975 10075 6995
rect 10093 6975 10105 6995
rect 10065 6965 10105 6975
rect 10175 6995 10215 7005
rect 10175 6975 10185 6995
rect 10203 6975 10215 6995
rect 10175 6965 10215 6975
rect 10285 6995 10325 7005
rect 10285 6975 10295 6995
rect 10313 6975 10325 6995
rect 10285 6965 10325 6975
rect 10395 6995 10435 7005
rect 10395 6975 10405 6995
rect 10423 6975 10435 6995
rect 10395 6965 10435 6975
rect 10505 6995 10545 7005
rect 10505 6975 10515 6995
rect 10533 6975 10545 6995
rect 10505 6965 10545 6975
rect 10615 6995 10655 7005
rect 10615 6975 10625 6995
rect 10643 6975 10655 6995
rect 10615 6965 10655 6975
rect 10725 6995 10765 7005
rect 10725 6975 10735 6995
rect 10753 6975 10765 6995
rect 10725 6965 10765 6975
rect 10835 6995 10875 7005
rect 10835 6975 10845 6995
rect 10863 6975 10875 6995
rect 11240 6995 11245 7015
rect 11265 6995 11285 7015
rect 11305 6995 11310 7015
rect 11240 6985 11310 6995
rect 11335 7115 11365 7125
rect 11335 7095 11340 7115
rect 11360 7095 11365 7115
rect 11335 7065 11365 7095
rect 11335 7045 11340 7065
rect 11360 7045 11365 7065
rect 11335 7015 11365 7045
rect 11335 6995 11340 7015
rect 11360 6995 11365 7015
rect 11335 6985 11365 6995
rect 11390 7115 11420 7125
rect 11390 7095 11395 7115
rect 11415 7095 11420 7115
rect 11390 7065 11420 7095
rect 11390 7045 11395 7065
rect 11415 7045 11420 7065
rect 11390 7015 11420 7045
rect 11390 6995 11395 7015
rect 11415 6995 11420 7015
rect 11390 6985 11420 6995
rect 11445 7115 11475 7125
rect 11445 7095 11450 7115
rect 11470 7095 11475 7115
rect 11445 7065 11475 7095
rect 11445 7045 11450 7065
rect 11470 7045 11475 7065
rect 11445 7015 11475 7045
rect 11445 6995 11450 7015
rect 11470 6995 11475 7015
rect 11445 6985 11475 6995
rect 11500 7115 11530 7125
rect 11500 7095 11505 7115
rect 11525 7095 11530 7115
rect 11500 7065 11530 7095
rect 11500 7045 11505 7065
rect 11525 7045 11530 7065
rect 11500 7015 11530 7045
rect 11500 6995 11505 7015
rect 11525 6995 11530 7015
rect 11500 6985 11530 6995
rect 11555 7115 11585 7125
rect 11555 7095 11560 7115
rect 11580 7095 11585 7115
rect 11555 7065 11585 7095
rect 11555 7045 11560 7065
rect 11580 7045 11585 7065
rect 11555 7015 11585 7045
rect 11555 6995 11560 7015
rect 11580 6995 11585 7015
rect 11555 6985 11585 6995
rect 11610 7115 11640 7125
rect 11610 7095 11615 7115
rect 11635 7095 11640 7115
rect 11610 7065 11640 7095
rect 11610 7045 11615 7065
rect 11635 7045 11640 7065
rect 11610 7015 11640 7045
rect 11610 6995 11615 7015
rect 11635 6995 11640 7015
rect 11610 6985 11640 6995
rect 11665 7115 11695 7125
rect 11665 7095 11670 7115
rect 11690 7095 11695 7115
rect 11665 7065 11695 7095
rect 11665 7045 11670 7065
rect 11690 7045 11695 7065
rect 11665 7015 11695 7045
rect 11665 6995 11670 7015
rect 11690 6995 11695 7015
rect 11665 6985 11695 6995
rect 11720 7115 11750 7125
rect 11720 7095 11725 7115
rect 11745 7095 11750 7115
rect 11720 7065 11750 7095
rect 11720 7045 11725 7065
rect 11745 7045 11750 7065
rect 11720 7015 11750 7045
rect 11720 6995 11725 7015
rect 11745 6995 11750 7015
rect 11720 6985 11750 6995
rect 11775 7115 11805 7125
rect 11775 7095 11780 7115
rect 11800 7095 11805 7115
rect 11775 7065 11805 7095
rect 11775 7045 11780 7065
rect 11800 7045 11805 7065
rect 11775 7015 11805 7045
rect 11775 6995 11780 7015
rect 11800 6995 11805 7015
rect 11775 6985 11805 6995
rect 11830 7115 11860 7125
rect 11830 7095 11835 7115
rect 11855 7095 11860 7115
rect 11830 7065 11860 7095
rect 11830 7045 11835 7065
rect 11855 7045 11860 7065
rect 11830 7015 11860 7045
rect 11830 6995 11835 7015
rect 11855 6995 11860 7015
rect 11830 6985 11860 6995
rect 11885 7115 11915 7125
rect 11885 7095 11890 7115
rect 11910 7095 11915 7115
rect 11885 7065 11915 7095
rect 11885 7045 11890 7065
rect 11910 7045 11915 7065
rect 11885 7015 11915 7045
rect 11885 6995 11890 7015
rect 11910 6995 11915 7015
rect 11885 6985 11915 6995
rect 11940 7115 11970 7125
rect 11940 7095 11945 7115
rect 11965 7095 11970 7115
rect 11940 7065 11970 7095
rect 11940 7045 11945 7065
rect 11965 7045 11970 7065
rect 11940 7015 11970 7045
rect 11940 6995 11945 7015
rect 11965 6995 11970 7015
rect 11940 6985 11970 6995
rect 11995 7115 12025 7125
rect 11995 7095 12000 7115
rect 12020 7095 12025 7115
rect 11995 7065 12025 7095
rect 11995 7045 12000 7065
rect 12020 7045 12025 7065
rect 11995 7015 12025 7045
rect 11995 6995 12000 7015
rect 12020 6995 12025 7015
rect 11995 6985 12025 6995
rect 12050 7115 12080 7125
rect 12050 7095 12055 7115
rect 12075 7095 12080 7115
rect 12050 7065 12080 7095
rect 12050 7045 12055 7065
rect 12075 7045 12080 7065
rect 12050 7015 12080 7045
rect 12050 6995 12055 7015
rect 12075 6995 12080 7015
rect 12050 6985 12080 6995
rect 12105 7115 12135 7125
rect 12105 7095 12110 7115
rect 12130 7095 12135 7115
rect 12105 7065 12135 7095
rect 12105 7045 12110 7065
rect 12130 7045 12135 7065
rect 12105 7015 12135 7045
rect 12105 6995 12110 7015
rect 12130 6995 12135 7015
rect 12105 6985 12135 6995
rect 12160 7115 12190 7125
rect 12160 7095 12165 7115
rect 12185 7095 12190 7115
rect 12160 7065 12190 7095
rect 12160 7045 12165 7065
rect 12185 7045 12190 7065
rect 12160 7015 12190 7045
rect 12160 6995 12165 7015
rect 12185 6995 12190 7015
rect 12160 6985 12190 6995
rect 12215 7115 12245 7125
rect 12215 7095 12220 7115
rect 12240 7095 12245 7115
rect 12215 7065 12245 7095
rect 12215 7045 12220 7065
rect 12240 7045 12245 7065
rect 12215 7015 12245 7045
rect 12215 6995 12220 7015
rect 12240 6995 12245 7015
rect 12215 6985 12245 6995
rect 12270 7115 12300 7125
rect 12270 7095 12275 7115
rect 12295 7095 12300 7115
rect 12270 7065 12300 7095
rect 12270 7045 12275 7065
rect 12295 7045 12300 7065
rect 12270 7015 12300 7045
rect 12270 6995 12275 7015
rect 12295 6995 12300 7015
rect 12270 6985 12300 6995
rect 12325 7115 12355 7125
rect 12325 7095 12330 7115
rect 12350 7095 12355 7115
rect 12325 7065 12355 7095
rect 12325 7045 12330 7065
rect 12350 7045 12355 7065
rect 12325 7015 12355 7045
rect 12325 6995 12330 7015
rect 12350 6995 12355 7015
rect 12325 6985 12355 6995
rect 12380 7115 12410 7125
rect 12380 7095 12385 7115
rect 12405 7095 12410 7115
rect 12380 7065 12410 7095
rect 12380 7045 12385 7065
rect 12405 7045 12410 7065
rect 12380 7015 12410 7045
rect 12380 6995 12385 7015
rect 12405 6995 12410 7015
rect 12380 6985 12410 6995
rect 12435 7115 12465 7125
rect 12435 7095 12440 7115
rect 12460 7095 12465 7115
rect 12435 7065 12465 7095
rect 12435 7045 12440 7065
rect 12460 7045 12465 7065
rect 12435 7015 12465 7045
rect 12435 6995 12440 7015
rect 12460 6995 12465 7015
rect 12435 6985 12465 6995
rect 12490 7115 12560 7125
rect 12490 7095 12495 7115
rect 12515 7095 12535 7115
rect 12555 7095 12560 7115
rect 12490 7065 12560 7095
rect 12490 7045 12495 7065
rect 12515 7045 12535 7065
rect 12555 7045 12560 7065
rect 12490 7015 12560 7045
rect 12860 7105 12930 7135
rect 12860 7085 12865 7105
rect 12885 7085 12905 7105
rect 12925 7085 12930 7105
rect 12860 7055 12930 7085
rect 12860 7035 12865 7055
rect 12885 7035 12905 7055
rect 12925 7035 12930 7055
rect 12860 7025 12930 7035
rect 12955 7155 12985 7165
rect 12955 7135 12960 7155
rect 12980 7135 12985 7155
rect 12955 7105 12985 7135
rect 12955 7085 12960 7105
rect 12980 7085 12985 7105
rect 12955 7055 12985 7085
rect 12955 7035 12960 7055
rect 12980 7035 12985 7055
rect 12955 7025 12985 7035
rect 13010 7155 13040 7165
rect 13010 7135 13015 7155
rect 13035 7135 13040 7155
rect 13010 7105 13040 7135
rect 13010 7085 13015 7105
rect 13035 7085 13040 7105
rect 13010 7055 13040 7085
rect 13010 7035 13015 7055
rect 13035 7035 13040 7055
rect 13010 7025 13040 7035
rect 13065 7155 13095 7165
rect 13065 7135 13070 7155
rect 13090 7135 13095 7155
rect 13065 7105 13095 7135
rect 13065 7085 13070 7105
rect 13090 7085 13095 7105
rect 13065 7055 13095 7085
rect 13065 7035 13070 7055
rect 13090 7035 13095 7055
rect 13065 7025 13095 7035
rect 13120 7155 13150 7165
rect 13120 7135 13125 7155
rect 13145 7135 13150 7155
rect 13120 7105 13150 7135
rect 13120 7085 13125 7105
rect 13145 7085 13150 7105
rect 13120 7055 13150 7085
rect 13120 7035 13125 7055
rect 13145 7035 13150 7055
rect 13120 7025 13150 7035
rect 13175 7155 13205 7165
rect 13175 7135 13180 7155
rect 13200 7135 13205 7155
rect 13175 7105 13205 7135
rect 13175 7085 13180 7105
rect 13200 7085 13205 7105
rect 13175 7055 13205 7085
rect 13175 7035 13180 7055
rect 13200 7035 13205 7055
rect 13175 7025 13205 7035
rect 13230 7155 13260 7165
rect 13230 7135 13235 7155
rect 13255 7135 13260 7155
rect 13230 7105 13260 7135
rect 13230 7085 13235 7105
rect 13255 7085 13260 7105
rect 13230 7055 13260 7085
rect 13230 7035 13235 7055
rect 13255 7035 13260 7055
rect 13230 7025 13260 7035
rect 13285 7155 13315 7165
rect 13285 7135 13290 7155
rect 13310 7135 13315 7155
rect 13285 7105 13315 7135
rect 13285 7085 13290 7105
rect 13310 7085 13315 7105
rect 13285 7055 13315 7085
rect 13285 7035 13290 7055
rect 13310 7035 13315 7055
rect 13285 7025 13315 7035
rect 13340 7155 13370 7165
rect 13340 7135 13345 7155
rect 13365 7135 13370 7155
rect 13340 7105 13370 7135
rect 13340 7085 13345 7105
rect 13365 7085 13370 7105
rect 13340 7055 13370 7085
rect 13340 7035 13345 7055
rect 13365 7035 13370 7055
rect 13340 7025 13370 7035
rect 13395 7155 13425 7165
rect 13395 7135 13400 7155
rect 13420 7135 13425 7155
rect 13395 7105 13425 7135
rect 13395 7085 13400 7105
rect 13420 7085 13425 7105
rect 13395 7055 13425 7085
rect 13395 7035 13400 7055
rect 13420 7035 13425 7055
rect 13395 7025 13425 7035
rect 13450 7155 13480 7165
rect 13450 7135 13455 7155
rect 13475 7135 13480 7155
rect 13450 7105 13480 7135
rect 13450 7085 13455 7105
rect 13475 7085 13480 7105
rect 13450 7055 13480 7085
rect 13450 7035 13455 7055
rect 13475 7035 13480 7055
rect 13450 7025 13480 7035
rect 13505 7155 13535 7165
rect 13505 7135 13510 7155
rect 13530 7135 13535 7155
rect 13505 7105 13535 7135
rect 13505 7085 13510 7105
rect 13530 7085 13535 7105
rect 13505 7055 13535 7085
rect 13505 7035 13510 7055
rect 13530 7035 13535 7055
rect 13505 7025 13535 7035
rect 13560 7155 13590 7165
rect 13560 7135 13565 7155
rect 13585 7135 13590 7155
rect 13560 7105 13590 7135
rect 13560 7085 13565 7105
rect 13585 7085 13590 7105
rect 13560 7055 13590 7085
rect 13560 7035 13565 7055
rect 13585 7035 13590 7055
rect 13560 7025 13590 7035
rect 13615 7155 13645 7165
rect 13615 7135 13620 7155
rect 13640 7135 13645 7155
rect 13615 7105 13645 7135
rect 13615 7085 13620 7105
rect 13640 7085 13645 7105
rect 13615 7055 13645 7085
rect 13615 7035 13620 7055
rect 13640 7035 13645 7055
rect 13615 7025 13645 7035
rect 13670 7155 13700 7165
rect 13670 7135 13675 7155
rect 13695 7135 13700 7155
rect 13670 7105 13700 7135
rect 13670 7085 13675 7105
rect 13695 7085 13700 7105
rect 13670 7055 13700 7085
rect 13670 7035 13675 7055
rect 13695 7035 13700 7055
rect 13670 7025 13700 7035
rect 13725 7155 13755 7165
rect 13725 7135 13730 7155
rect 13750 7135 13755 7155
rect 13725 7105 13755 7135
rect 13725 7085 13730 7105
rect 13750 7085 13755 7105
rect 13725 7055 13755 7085
rect 13725 7035 13730 7055
rect 13750 7035 13755 7055
rect 13725 7025 13755 7035
rect 13780 7155 13810 7165
rect 13780 7135 13785 7155
rect 13805 7135 13810 7155
rect 13780 7105 13810 7135
rect 13780 7085 13785 7105
rect 13805 7085 13810 7105
rect 13780 7055 13810 7085
rect 13780 7035 13785 7055
rect 13805 7035 13810 7055
rect 13780 7025 13810 7035
rect 13835 7155 13865 7165
rect 13835 7135 13840 7155
rect 13860 7135 13865 7155
rect 13835 7105 13865 7135
rect 13835 7085 13840 7105
rect 13860 7085 13865 7105
rect 13835 7055 13865 7085
rect 13835 7035 13840 7055
rect 13860 7035 13865 7055
rect 13835 7025 13865 7035
rect 13890 7155 13920 7165
rect 13890 7135 13895 7155
rect 13915 7135 13920 7155
rect 13890 7105 13920 7135
rect 13890 7085 13895 7105
rect 13915 7085 13920 7105
rect 13890 7055 13920 7085
rect 13890 7035 13895 7055
rect 13915 7035 13920 7055
rect 13890 7025 13920 7035
rect 13945 7155 13975 7165
rect 13945 7135 13950 7155
rect 13970 7135 13975 7155
rect 13945 7105 13975 7135
rect 13945 7085 13950 7105
rect 13970 7085 13975 7105
rect 13945 7055 13975 7085
rect 13945 7035 13950 7055
rect 13970 7035 13975 7055
rect 13945 7025 13975 7035
rect 14000 7155 14030 7165
rect 14000 7135 14005 7155
rect 14025 7135 14030 7155
rect 14000 7105 14030 7135
rect 14000 7085 14005 7105
rect 14025 7085 14030 7105
rect 14000 7055 14030 7085
rect 14000 7035 14005 7055
rect 14025 7035 14030 7055
rect 14000 7025 14030 7035
rect 14055 7155 14085 7165
rect 14055 7135 14060 7155
rect 14080 7135 14085 7155
rect 14055 7105 14085 7135
rect 14055 7085 14060 7105
rect 14080 7085 14085 7105
rect 14055 7055 14085 7085
rect 14055 7035 14060 7055
rect 14080 7035 14085 7055
rect 14055 7025 14085 7035
rect 14110 7155 14180 7165
rect 14110 7135 14115 7155
rect 14135 7135 14155 7155
rect 14175 7135 14180 7155
rect 14110 7105 14180 7135
rect 14110 7085 14115 7105
rect 14135 7085 14155 7105
rect 14175 7085 14180 7105
rect 14110 7055 14180 7085
rect 14110 7035 14115 7055
rect 14135 7035 14155 7055
rect 14175 7035 14180 7055
rect 14110 7025 14180 7035
rect 17145 7155 17215 7165
rect 17145 7135 17150 7155
rect 17170 7135 17190 7155
rect 17210 7135 17215 7155
rect 17145 7105 17215 7135
rect 17145 7085 17150 7105
rect 17170 7085 17190 7105
rect 17210 7085 17215 7105
rect 17145 7055 17215 7085
rect 17145 7035 17150 7055
rect 17170 7035 17190 7055
rect 17210 7035 17215 7055
rect 17145 7025 17215 7035
rect 17240 7155 17270 7165
rect 17240 7135 17245 7155
rect 17265 7135 17270 7155
rect 17240 7105 17270 7135
rect 17240 7085 17245 7105
rect 17265 7085 17270 7105
rect 17240 7055 17270 7085
rect 17240 7035 17245 7055
rect 17265 7035 17270 7055
rect 17240 7025 17270 7035
rect 17295 7155 17325 7165
rect 17295 7135 17300 7155
rect 17320 7135 17325 7155
rect 17295 7105 17325 7135
rect 17295 7085 17300 7105
rect 17320 7085 17325 7105
rect 17295 7055 17325 7085
rect 17295 7035 17300 7055
rect 17320 7035 17325 7055
rect 17295 7025 17325 7035
rect 17350 7155 17380 7165
rect 17350 7135 17355 7155
rect 17375 7135 17380 7155
rect 17350 7105 17380 7135
rect 17350 7085 17355 7105
rect 17375 7085 17380 7105
rect 17350 7055 17380 7085
rect 17350 7035 17355 7055
rect 17375 7035 17380 7055
rect 17350 7025 17380 7035
rect 17405 7155 17435 7165
rect 17405 7135 17410 7155
rect 17430 7135 17435 7155
rect 17405 7105 17435 7135
rect 17405 7085 17410 7105
rect 17430 7085 17435 7105
rect 17405 7055 17435 7085
rect 17405 7035 17410 7055
rect 17430 7035 17435 7055
rect 17405 7025 17435 7035
rect 17460 7155 17490 7165
rect 17460 7135 17465 7155
rect 17485 7135 17490 7155
rect 17460 7105 17490 7135
rect 17460 7085 17465 7105
rect 17485 7085 17490 7105
rect 17460 7055 17490 7085
rect 17460 7035 17465 7055
rect 17485 7035 17490 7055
rect 17460 7025 17490 7035
rect 17515 7155 17545 7165
rect 17515 7135 17520 7155
rect 17540 7135 17545 7155
rect 17515 7105 17545 7135
rect 17515 7085 17520 7105
rect 17540 7085 17545 7105
rect 17515 7055 17545 7085
rect 17515 7035 17520 7055
rect 17540 7035 17545 7055
rect 17515 7025 17545 7035
rect 17570 7155 17600 7165
rect 17570 7135 17575 7155
rect 17595 7135 17600 7155
rect 17570 7105 17600 7135
rect 17570 7085 17575 7105
rect 17595 7085 17600 7105
rect 17570 7055 17600 7085
rect 17570 7035 17575 7055
rect 17595 7035 17600 7055
rect 17570 7025 17600 7035
rect 17625 7155 17655 7165
rect 17625 7135 17630 7155
rect 17650 7135 17655 7155
rect 17625 7105 17655 7135
rect 17625 7085 17630 7105
rect 17650 7085 17655 7105
rect 17625 7055 17655 7085
rect 17625 7035 17630 7055
rect 17650 7035 17655 7055
rect 17625 7025 17655 7035
rect 17680 7155 17710 7165
rect 17680 7135 17685 7155
rect 17705 7135 17710 7155
rect 17680 7105 17710 7135
rect 17680 7085 17685 7105
rect 17705 7085 17710 7105
rect 17680 7055 17710 7085
rect 17680 7035 17685 7055
rect 17705 7035 17710 7055
rect 17680 7025 17710 7035
rect 17735 7155 17765 7165
rect 17735 7135 17740 7155
rect 17760 7135 17765 7155
rect 17735 7105 17765 7135
rect 17735 7085 17740 7105
rect 17760 7085 17765 7105
rect 17735 7055 17765 7085
rect 17735 7035 17740 7055
rect 17760 7035 17765 7055
rect 17735 7025 17765 7035
rect 17790 7155 17820 7165
rect 17790 7135 17795 7155
rect 17815 7135 17820 7155
rect 17790 7105 17820 7135
rect 17790 7085 17795 7105
rect 17815 7085 17820 7105
rect 17790 7055 17820 7085
rect 17790 7035 17795 7055
rect 17815 7035 17820 7055
rect 17790 7025 17820 7035
rect 17845 7155 17875 7165
rect 17845 7135 17850 7155
rect 17870 7135 17875 7155
rect 17845 7105 17875 7135
rect 17845 7085 17850 7105
rect 17870 7085 17875 7105
rect 17845 7055 17875 7085
rect 17845 7035 17850 7055
rect 17870 7035 17875 7055
rect 17845 7025 17875 7035
rect 17900 7155 17930 7165
rect 17900 7135 17905 7155
rect 17925 7135 17930 7155
rect 17900 7105 17930 7135
rect 17900 7085 17905 7105
rect 17925 7085 17930 7105
rect 17900 7055 17930 7085
rect 17900 7035 17905 7055
rect 17925 7035 17930 7055
rect 17900 7025 17930 7035
rect 17955 7155 17985 7165
rect 17955 7135 17960 7155
rect 17980 7135 17985 7155
rect 17955 7105 17985 7135
rect 17955 7085 17960 7105
rect 17980 7085 17985 7105
rect 17955 7055 17985 7085
rect 17955 7035 17960 7055
rect 17980 7035 17985 7055
rect 17955 7025 17985 7035
rect 18010 7155 18040 7165
rect 18010 7135 18015 7155
rect 18035 7135 18040 7155
rect 18010 7105 18040 7135
rect 18010 7085 18015 7105
rect 18035 7085 18040 7105
rect 18010 7055 18040 7085
rect 18010 7035 18015 7055
rect 18035 7035 18040 7055
rect 18010 7025 18040 7035
rect 18065 7155 18095 7165
rect 18065 7135 18070 7155
rect 18090 7135 18095 7155
rect 18065 7105 18095 7135
rect 18065 7085 18070 7105
rect 18090 7085 18095 7105
rect 18065 7055 18095 7085
rect 18065 7035 18070 7055
rect 18090 7035 18095 7055
rect 18065 7025 18095 7035
rect 18120 7155 18150 7165
rect 18120 7135 18125 7155
rect 18145 7135 18150 7155
rect 18120 7105 18150 7135
rect 18120 7085 18125 7105
rect 18145 7085 18150 7105
rect 18120 7055 18150 7085
rect 18120 7035 18125 7055
rect 18145 7035 18150 7055
rect 18120 7025 18150 7035
rect 18175 7155 18205 7165
rect 18175 7135 18180 7155
rect 18200 7135 18205 7155
rect 18175 7105 18205 7135
rect 18175 7085 18180 7105
rect 18200 7085 18205 7105
rect 18175 7055 18205 7085
rect 18175 7035 18180 7055
rect 18200 7035 18205 7055
rect 18175 7025 18205 7035
rect 18230 7155 18260 7165
rect 18230 7135 18235 7155
rect 18255 7135 18260 7155
rect 18230 7105 18260 7135
rect 18230 7085 18235 7105
rect 18255 7085 18260 7105
rect 18230 7055 18260 7085
rect 18230 7035 18235 7055
rect 18255 7035 18260 7055
rect 18230 7025 18260 7035
rect 18285 7155 18315 7165
rect 18285 7135 18290 7155
rect 18310 7135 18315 7155
rect 18285 7105 18315 7135
rect 18285 7085 18290 7105
rect 18310 7085 18315 7105
rect 18285 7055 18315 7085
rect 18285 7035 18290 7055
rect 18310 7035 18315 7055
rect 18285 7025 18315 7035
rect 18340 7155 18370 7165
rect 18340 7135 18345 7155
rect 18365 7135 18370 7155
rect 18340 7105 18370 7135
rect 18340 7085 18345 7105
rect 18365 7085 18370 7105
rect 18340 7055 18370 7085
rect 18340 7035 18345 7055
rect 18365 7035 18370 7055
rect 18340 7025 18370 7035
rect 18395 7155 18465 7165
rect 18395 7135 18400 7155
rect 18420 7135 18440 7155
rect 18460 7135 18465 7155
rect 18830 7155 18840 7175
rect 18860 7155 18870 7175
rect 18830 7145 18870 7155
rect 18940 7175 18980 7185
rect 18940 7155 18950 7175
rect 18970 7155 18980 7175
rect 18940 7145 18980 7155
rect 19050 7175 19090 7185
rect 19050 7155 19060 7175
rect 19080 7155 19090 7175
rect 19050 7145 19090 7155
rect 19160 7175 19200 7185
rect 19160 7155 19170 7175
rect 19190 7155 19200 7175
rect 19160 7145 19200 7155
rect 19270 7175 19310 7185
rect 19270 7155 19280 7175
rect 19300 7155 19310 7175
rect 19270 7145 19310 7155
rect 19380 7175 19420 7185
rect 19380 7155 19390 7175
rect 19410 7155 19420 7175
rect 19380 7145 19420 7155
rect 19490 7175 19530 7185
rect 19490 7155 19500 7175
rect 19520 7155 19530 7175
rect 19490 7145 19530 7155
rect 19600 7175 19640 7185
rect 19600 7155 19610 7175
rect 19630 7155 19640 7175
rect 19600 7145 19640 7155
rect 19710 7175 19750 7185
rect 19710 7155 19720 7175
rect 19740 7155 19750 7175
rect 19710 7145 19750 7155
rect 19820 7175 19860 7185
rect 19820 7155 19830 7175
rect 19850 7155 19860 7175
rect 19820 7145 19860 7155
rect 19930 7175 19970 7185
rect 19930 7155 19940 7175
rect 19960 7155 19970 7175
rect 20360 7165 20380 7185
rect 20510 7165 20530 7185
rect 20620 7165 20640 7185
rect 20730 7165 20750 7185
rect 20840 7165 20860 7185
rect 20950 7165 20970 7185
rect 21060 7165 21080 7185
rect 21170 7165 21190 7185
rect 21280 7165 21300 7185
rect 21390 7165 21410 7185
rect 21500 7165 21520 7185
rect 21650 7165 21670 7185
rect 19930 7145 19970 7155
rect 20355 7155 20425 7165
rect 18395 7105 18465 7135
rect 18840 7125 18860 7145
rect 18950 7125 18970 7145
rect 19060 7125 19080 7145
rect 19170 7125 19190 7145
rect 19280 7125 19300 7145
rect 19390 7125 19410 7145
rect 19500 7125 19520 7145
rect 19610 7125 19630 7145
rect 19720 7125 19740 7145
rect 19830 7125 19850 7145
rect 19940 7125 19960 7145
rect 20355 7135 20360 7155
rect 20380 7135 20400 7155
rect 20420 7135 20425 7155
rect 18395 7085 18400 7105
rect 18420 7085 18440 7105
rect 18460 7085 18465 7105
rect 18395 7055 18465 7085
rect 18395 7035 18400 7055
rect 18420 7035 18440 7055
rect 18460 7035 18465 7055
rect 18395 7025 18465 7035
rect 18740 7115 18810 7125
rect 18740 7095 18745 7115
rect 18765 7095 18785 7115
rect 18805 7095 18810 7115
rect 18740 7065 18810 7095
rect 18740 7045 18745 7065
rect 18765 7045 18785 7065
rect 18805 7045 18810 7065
rect 12490 6995 12495 7015
rect 12515 6995 12535 7015
rect 12555 6995 12560 7015
rect 12960 7005 12980 7025
rect 13070 7005 13090 7025
rect 13180 7005 13200 7025
rect 13290 7005 13310 7025
rect 13400 7005 13420 7025
rect 13510 7005 13530 7025
rect 13620 7005 13640 7025
rect 13730 7005 13750 7025
rect 13840 7005 13860 7025
rect 13950 7005 13970 7025
rect 14060 7005 14080 7025
rect 17245 7005 17265 7025
rect 17355 7005 17375 7025
rect 17465 7005 17485 7025
rect 17575 7005 17595 7025
rect 17685 7005 17705 7025
rect 17795 7005 17815 7025
rect 17905 7005 17925 7025
rect 18015 7005 18035 7025
rect 18125 7005 18145 7025
rect 18235 7005 18255 7025
rect 18345 7005 18365 7025
rect 18740 7015 18810 7045
rect 12490 6985 12560 6995
rect 12950 6995 12990 7005
rect 10835 6965 10875 6975
rect 11245 6965 11265 6985
rect 11395 6965 11415 6985
rect 11505 6965 11525 6985
rect 11615 6965 11635 6985
rect 11725 6965 11745 6985
rect 11835 6965 11855 6985
rect 11945 6965 11965 6985
rect 12055 6965 12075 6985
rect 12165 6965 12185 6985
rect 12275 6965 12295 6985
rect 12385 6965 12405 6985
rect 12535 6965 12555 6985
rect 12950 6975 12962 6995
rect 12980 6975 12990 6995
rect 12950 6965 12990 6975
rect 13060 6995 13100 7005
rect 13060 6975 13072 6995
rect 13090 6975 13100 6995
rect 13060 6965 13100 6975
rect 13170 6995 13210 7005
rect 13170 6975 13182 6995
rect 13200 6975 13210 6995
rect 13170 6965 13210 6975
rect 13280 6995 13320 7005
rect 13280 6975 13292 6995
rect 13310 6975 13320 6995
rect 13280 6965 13320 6975
rect 13390 6995 13430 7005
rect 13390 6975 13402 6995
rect 13420 6975 13430 6995
rect 13390 6965 13430 6975
rect 13500 6995 13540 7005
rect 13500 6975 13512 6995
rect 13530 6975 13540 6995
rect 13500 6965 13540 6975
rect 13610 6995 13650 7005
rect 13610 6975 13622 6995
rect 13640 6975 13650 6995
rect 13610 6965 13650 6975
rect 13720 6995 13760 7005
rect 13720 6975 13732 6995
rect 13750 6975 13760 6995
rect 13720 6965 13760 6975
rect 13830 6995 13870 7005
rect 13830 6975 13842 6995
rect 13860 6975 13870 6995
rect 13830 6965 13870 6975
rect 13940 6995 13980 7005
rect 13940 6975 13952 6995
rect 13970 6975 13980 6995
rect 13940 6965 13980 6975
rect 14050 6995 14090 7005
rect 14050 6975 14062 6995
rect 14080 6975 14090 6995
rect 14050 6965 14090 6975
rect 17235 6995 17275 7005
rect 17235 6975 17245 6995
rect 17263 6975 17275 6995
rect 17235 6965 17275 6975
rect 17345 6995 17385 7005
rect 17345 6975 17355 6995
rect 17373 6975 17385 6995
rect 17345 6965 17385 6975
rect 17455 6995 17495 7005
rect 17455 6975 17465 6995
rect 17483 6975 17495 6995
rect 17455 6965 17495 6975
rect 17565 6995 17605 7005
rect 17565 6975 17575 6995
rect 17593 6975 17605 6995
rect 17565 6965 17605 6975
rect 17675 6995 17715 7005
rect 17675 6975 17685 6995
rect 17703 6975 17715 6995
rect 17675 6965 17715 6975
rect 17785 6995 17825 7005
rect 17785 6975 17795 6995
rect 17813 6975 17825 6995
rect 17785 6965 17825 6975
rect 17895 6995 17935 7005
rect 17895 6975 17905 6995
rect 17923 6975 17935 6995
rect 17895 6965 17935 6975
rect 18005 6995 18045 7005
rect 18005 6975 18015 6995
rect 18033 6975 18045 6995
rect 18005 6965 18045 6975
rect 18115 6995 18155 7005
rect 18115 6975 18125 6995
rect 18143 6975 18155 6995
rect 18115 6965 18155 6975
rect 18225 6995 18265 7005
rect 18225 6975 18235 6995
rect 18253 6975 18265 6995
rect 18225 6965 18265 6975
rect 18335 6995 18375 7005
rect 18335 6975 18345 6995
rect 18363 6975 18375 6995
rect 18740 6995 18745 7015
rect 18765 6995 18785 7015
rect 18805 6995 18810 7015
rect 18740 6985 18810 6995
rect 18835 7115 18865 7125
rect 18835 7095 18840 7115
rect 18860 7095 18865 7115
rect 18835 7065 18865 7095
rect 18835 7045 18840 7065
rect 18860 7045 18865 7065
rect 18835 7015 18865 7045
rect 18835 6995 18840 7015
rect 18860 6995 18865 7015
rect 18835 6985 18865 6995
rect 18890 7115 18920 7125
rect 18890 7095 18895 7115
rect 18915 7095 18920 7115
rect 18890 7065 18920 7095
rect 18890 7045 18895 7065
rect 18915 7045 18920 7065
rect 18890 7015 18920 7045
rect 18890 6995 18895 7015
rect 18915 6995 18920 7015
rect 18890 6985 18920 6995
rect 18945 7115 18975 7125
rect 18945 7095 18950 7115
rect 18970 7095 18975 7115
rect 18945 7065 18975 7095
rect 18945 7045 18950 7065
rect 18970 7045 18975 7065
rect 18945 7015 18975 7045
rect 18945 6995 18950 7015
rect 18970 6995 18975 7015
rect 18945 6985 18975 6995
rect 19000 7115 19030 7125
rect 19000 7095 19005 7115
rect 19025 7095 19030 7115
rect 19000 7065 19030 7095
rect 19000 7045 19005 7065
rect 19025 7045 19030 7065
rect 19000 7015 19030 7045
rect 19000 6995 19005 7015
rect 19025 6995 19030 7015
rect 19000 6985 19030 6995
rect 19055 7115 19085 7125
rect 19055 7095 19060 7115
rect 19080 7095 19085 7115
rect 19055 7065 19085 7095
rect 19055 7045 19060 7065
rect 19080 7045 19085 7065
rect 19055 7015 19085 7045
rect 19055 6995 19060 7015
rect 19080 6995 19085 7015
rect 19055 6985 19085 6995
rect 19110 7115 19140 7125
rect 19110 7095 19115 7115
rect 19135 7095 19140 7115
rect 19110 7065 19140 7095
rect 19110 7045 19115 7065
rect 19135 7045 19140 7065
rect 19110 7015 19140 7045
rect 19110 6995 19115 7015
rect 19135 6995 19140 7015
rect 19110 6985 19140 6995
rect 19165 7115 19195 7125
rect 19165 7095 19170 7115
rect 19190 7095 19195 7115
rect 19165 7065 19195 7095
rect 19165 7045 19170 7065
rect 19190 7045 19195 7065
rect 19165 7015 19195 7045
rect 19165 6995 19170 7015
rect 19190 6995 19195 7015
rect 19165 6985 19195 6995
rect 19220 7115 19250 7125
rect 19220 7095 19225 7115
rect 19245 7095 19250 7115
rect 19220 7065 19250 7095
rect 19220 7045 19225 7065
rect 19245 7045 19250 7065
rect 19220 7015 19250 7045
rect 19220 6995 19225 7015
rect 19245 6995 19250 7015
rect 19220 6985 19250 6995
rect 19275 7115 19305 7125
rect 19275 7095 19280 7115
rect 19300 7095 19305 7115
rect 19275 7065 19305 7095
rect 19275 7045 19280 7065
rect 19300 7045 19305 7065
rect 19275 7015 19305 7045
rect 19275 6995 19280 7015
rect 19300 6995 19305 7015
rect 19275 6985 19305 6995
rect 19330 7115 19360 7125
rect 19330 7095 19335 7115
rect 19355 7095 19360 7115
rect 19330 7065 19360 7095
rect 19330 7045 19335 7065
rect 19355 7045 19360 7065
rect 19330 7015 19360 7045
rect 19330 6995 19335 7015
rect 19355 6995 19360 7015
rect 19330 6985 19360 6995
rect 19385 7115 19415 7125
rect 19385 7095 19390 7115
rect 19410 7095 19415 7115
rect 19385 7065 19415 7095
rect 19385 7045 19390 7065
rect 19410 7045 19415 7065
rect 19385 7015 19415 7045
rect 19385 6995 19390 7015
rect 19410 6995 19415 7015
rect 19385 6985 19415 6995
rect 19440 7115 19470 7125
rect 19440 7095 19445 7115
rect 19465 7095 19470 7115
rect 19440 7065 19470 7095
rect 19440 7045 19445 7065
rect 19465 7045 19470 7065
rect 19440 7015 19470 7045
rect 19440 6995 19445 7015
rect 19465 6995 19470 7015
rect 19440 6985 19470 6995
rect 19495 7115 19525 7125
rect 19495 7095 19500 7115
rect 19520 7095 19525 7115
rect 19495 7065 19525 7095
rect 19495 7045 19500 7065
rect 19520 7045 19525 7065
rect 19495 7015 19525 7045
rect 19495 6995 19500 7015
rect 19520 6995 19525 7015
rect 19495 6985 19525 6995
rect 19550 7115 19580 7125
rect 19550 7095 19555 7115
rect 19575 7095 19580 7115
rect 19550 7065 19580 7095
rect 19550 7045 19555 7065
rect 19575 7045 19580 7065
rect 19550 7015 19580 7045
rect 19550 6995 19555 7015
rect 19575 6995 19580 7015
rect 19550 6985 19580 6995
rect 19605 7115 19635 7125
rect 19605 7095 19610 7115
rect 19630 7095 19635 7115
rect 19605 7065 19635 7095
rect 19605 7045 19610 7065
rect 19630 7045 19635 7065
rect 19605 7015 19635 7045
rect 19605 6995 19610 7015
rect 19630 6995 19635 7015
rect 19605 6985 19635 6995
rect 19660 7115 19690 7125
rect 19660 7095 19665 7115
rect 19685 7095 19690 7115
rect 19660 7065 19690 7095
rect 19660 7045 19665 7065
rect 19685 7045 19690 7065
rect 19660 7015 19690 7045
rect 19660 6995 19665 7015
rect 19685 6995 19690 7015
rect 19660 6985 19690 6995
rect 19715 7115 19745 7125
rect 19715 7095 19720 7115
rect 19740 7095 19745 7115
rect 19715 7065 19745 7095
rect 19715 7045 19720 7065
rect 19740 7045 19745 7065
rect 19715 7015 19745 7045
rect 19715 6995 19720 7015
rect 19740 6995 19745 7015
rect 19715 6985 19745 6995
rect 19770 7115 19800 7125
rect 19770 7095 19775 7115
rect 19795 7095 19800 7115
rect 19770 7065 19800 7095
rect 19770 7045 19775 7065
rect 19795 7045 19800 7065
rect 19770 7015 19800 7045
rect 19770 6995 19775 7015
rect 19795 6995 19800 7015
rect 19770 6985 19800 6995
rect 19825 7115 19855 7125
rect 19825 7095 19830 7115
rect 19850 7095 19855 7115
rect 19825 7065 19855 7095
rect 19825 7045 19830 7065
rect 19850 7045 19855 7065
rect 19825 7015 19855 7045
rect 19825 6995 19830 7015
rect 19850 6995 19855 7015
rect 19825 6985 19855 6995
rect 19880 7115 19910 7125
rect 19880 7095 19885 7115
rect 19905 7095 19910 7115
rect 19880 7065 19910 7095
rect 19880 7045 19885 7065
rect 19905 7045 19910 7065
rect 19880 7015 19910 7045
rect 19880 6995 19885 7015
rect 19905 6995 19910 7015
rect 19880 6985 19910 6995
rect 19935 7115 19965 7125
rect 19935 7095 19940 7115
rect 19960 7095 19965 7115
rect 19935 7065 19965 7095
rect 19935 7045 19940 7065
rect 19960 7045 19965 7065
rect 19935 7015 19965 7045
rect 19935 6995 19940 7015
rect 19960 6995 19965 7015
rect 19935 6985 19965 6995
rect 19990 7115 20060 7125
rect 19990 7095 19995 7115
rect 20015 7095 20035 7115
rect 20055 7095 20060 7115
rect 19990 7065 20060 7095
rect 19990 7045 19995 7065
rect 20015 7045 20035 7065
rect 20055 7045 20060 7065
rect 19990 7015 20060 7045
rect 20355 7105 20425 7135
rect 20355 7085 20360 7105
rect 20380 7085 20400 7105
rect 20420 7085 20425 7105
rect 20355 7055 20425 7085
rect 20355 7035 20360 7055
rect 20380 7035 20400 7055
rect 20420 7035 20425 7055
rect 20355 7025 20425 7035
rect 20450 7155 20480 7165
rect 20450 7135 20455 7155
rect 20475 7135 20480 7155
rect 20450 7105 20480 7135
rect 20450 7085 20455 7105
rect 20475 7085 20480 7105
rect 20450 7055 20480 7085
rect 20450 7035 20455 7055
rect 20475 7035 20480 7055
rect 20450 7025 20480 7035
rect 20505 7155 20535 7165
rect 20505 7135 20510 7155
rect 20530 7135 20535 7155
rect 20505 7105 20535 7135
rect 20505 7085 20510 7105
rect 20530 7085 20535 7105
rect 20505 7055 20535 7085
rect 20505 7035 20510 7055
rect 20530 7035 20535 7055
rect 20505 7025 20535 7035
rect 20560 7155 20590 7165
rect 20560 7135 20565 7155
rect 20585 7135 20590 7155
rect 20560 7105 20590 7135
rect 20560 7085 20565 7105
rect 20585 7085 20590 7105
rect 20560 7055 20590 7085
rect 20560 7035 20565 7055
rect 20585 7035 20590 7055
rect 20560 7025 20590 7035
rect 20615 7155 20645 7165
rect 20615 7135 20620 7155
rect 20640 7135 20645 7155
rect 20615 7105 20645 7135
rect 20615 7085 20620 7105
rect 20640 7085 20645 7105
rect 20615 7055 20645 7085
rect 20615 7035 20620 7055
rect 20640 7035 20645 7055
rect 20615 7025 20645 7035
rect 20670 7155 20700 7165
rect 20670 7135 20675 7155
rect 20695 7135 20700 7155
rect 20670 7105 20700 7135
rect 20670 7085 20675 7105
rect 20695 7085 20700 7105
rect 20670 7055 20700 7085
rect 20670 7035 20675 7055
rect 20695 7035 20700 7055
rect 20670 7025 20700 7035
rect 20725 7155 20755 7165
rect 20725 7135 20730 7155
rect 20750 7135 20755 7155
rect 20725 7105 20755 7135
rect 20725 7085 20730 7105
rect 20750 7085 20755 7105
rect 20725 7055 20755 7085
rect 20725 7035 20730 7055
rect 20750 7035 20755 7055
rect 20725 7025 20755 7035
rect 20780 7155 20810 7165
rect 20780 7135 20785 7155
rect 20805 7135 20810 7155
rect 20780 7105 20810 7135
rect 20780 7085 20785 7105
rect 20805 7085 20810 7105
rect 20780 7055 20810 7085
rect 20780 7035 20785 7055
rect 20805 7035 20810 7055
rect 20780 7025 20810 7035
rect 20835 7155 20865 7165
rect 20835 7135 20840 7155
rect 20860 7135 20865 7155
rect 20835 7105 20865 7135
rect 20835 7085 20840 7105
rect 20860 7085 20865 7105
rect 20835 7055 20865 7085
rect 20835 7035 20840 7055
rect 20860 7035 20865 7055
rect 20835 7025 20865 7035
rect 20890 7155 20920 7165
rect 20890 7135 20895 7155
rect 20915 7135 20920 7155
rect 20890 7105 20920 7135
rect 20890 7085 20895 7105
rect 20915 7085 20920 7105
rect 20890 7055 20920 7085
rect 20890 7035 20895 7055
rect 20915 7035 20920 7055
rect 20890 7025 20920 7035
rect 20945 7155 20975 7165
rect 20945 7135 20950 7155
rect 20970 7135 20975 7155
rect 20945 7105 20975 7135
rect 20945 7085 20950 7105
rect 20970 7085 20975 7105
rect 20945 7055 20975 7085
rect 20945 7035 20950 7055
rect 20970 7035 20975 7055
rect 20945 7025 20975 7035
rect 21000 7155 21030 7165
rect 21000 7135 21005 7155
rect 21025 7135 21030 7155
rect 21000 7105 21030 7135
rect 21000 7085 21005 7105
rect 21025 7085 21030 7105
rect 21000 7055 21030 7085
rect 21000 7035 21005 7055
rect 21025 7035 21030 7055
rect 21000 7025 21030 7035
rect 21055 7155 21085 7165
rect 21055 7135 21060 7155
rect 21080 7135 21085 7155
rect 21055 7105 21085 7135
rect 21055 7085 21060 7105
rect 21080 7085 21085 7105
rect 21055 7055 21085 7085
rect 21055 7035 21060 7055
rect 21080 7035 21085 7055
rect 21055 7025 21085 7035
rect 21110 7155 21140 7165
rect 21110 7135 21115 7155
rect 21135 7135 21140 7155
rect 21110 7105 21140 7135
rect 21110 7085 21115 7105
rect 21135 7085 21140 7105
rect 21110 7055 21140 7085
rect 21110 7035 21115 7055
rect 21135 7035 21140 7055
rect 21110 7025 21140 7035
rect 21165 7155 21195 7165
rect 21165 7135 21170 7155
rect 21190 7135 21195 7155
rect 21165 7105 21195 7135
rect 21165 7085 21170 7105
rect 21190 7085 21195 7105
rect 21165 7055 21195 7085
rect 21165 7035 21170 7055
rect 21190 7035 21195 7055
rect 21165 7025 21195 7035
rect 21220 7155 21250 7165
rect 21220 7135 21225 7155
rect 21245 7135 21250 7155
rect 21220 7105 21250 7135
rect 21220 7085 21225 7105
rect 21245 7085 21250 7105
rect 21220 7055 21250 7085
rect 21220 7035 21225 7055
rect 21245 7035 21250 7055
rect 21220 7025 21250 7035
rect 21275 7155 21305 7165
rect 21275 7135 21280 7155
rect 21300 7135 21305 7155
rect 21275 7105 21305 7135
rect 21275 7085 21280 7105
rect 21300 7085 21305 7105
rect 21275 7055 21305 7085
rect 21275 7035 21280 7055
rect 21300 7035 21305 7055
rect 21275 7025 21305 7035
rect 21330 7155 21360 7165
rect 21330 7135 21335 7155
rect 21355 7135 21360 7155
rect 21330 7105 21360 7135
rect 21330 7085 21335 7105
rect 21355 7085 21360 7105
rect 21330 7055 21360 7085
rect 21330 7035 21335 7055
rect 21355 7035 21360 7055
rect 21330 7025 21360 7035
rect 21385 7155 21415 7165
rect 21385 7135 21390 7155
rect 21410 7135 21415 7155
rect 21385 7105 21415 7135
rect 21385 7085 21390 7105
rect 21410 7085 21415 7105
rect 21385 7055 21415 7085
rect 21385 7035 21390 7055
rect 21410 7035 21415 7055
rect 21385 7025 21415 7035
rect 21440 7155 21470 7165
rect 21440 7135 21445 7155
rect 21465 7135 21470 7155
rect 21440 7105 21470 7135
rect 21440 7085 21445 7105
rect 21465 7085 21470 7105
rect 21440 7055 21470 7085
rect 21440 7035 21445 7055
rect 21465 7035 21470 7055
rect 21440 7025 21470 7035
rect 21495 7155 21525 7165
rect 21495 7135 21500 7155
rect 21520 7135 21525 7155
rect 21495 7105 21525 7135
rect 21495 7085 21500 7105
rect 21520 7085 21525 7105
rect 21495 7055 21525 7085
rect 21495 7035 21500 7055
rect 21520 7035 21525 7055
rect 21495 7025 21525 7035
rect 21550 7155 21580 7165
rect 21550 7135 21555 7155
rect 21575 7135 21580 7155
rect 21550 7105 21580 7135
rect 21550 7085 21555 7105
rect 21575 7085 21580 7105
rect 21550 7055 21580 7085
rect 21550 7035 21555 7055
rect 21575 7035 21580 7055
rect 21550 7025 21580 7035
rect 21605 7155 21675 7165
rect 21605 7135 21610 7155
rect 21630 7135 21650 7155
rect 21670 7135 21675 7155
rect 21605 7105 21675 7135
rect 21605 7085 21610 7105
rect 21630 7085 21650 7105
rect 21670 7085 21675 7105
rect 21605 7055 21675 7085
rect 21605 7035 21610 7055
rect 21630 7035 21650 7055
rect 21670 7035 21675 7055
rect 21605 7025 21675 7035
rect 19990 6995 19995 7015
rect 20015 6995 20035 7015
rect 20055 6995 20060 7015
rect 20455 7005 20475 7025
rect 20565 7005 20585 7025
rect 20675 7005 20695 7025
rect 20785 7005 20805 7025
rect 20895 7005 20915 7025
rect 21005 7005 21025 7025
rect 21115 7005 21135 7025
rect 21225 7005 21245 7025
rect 21335 7005 21355 7025
rect 21445 7005 21465 7025
rect 21555 7005 21575 7025
rect 19990 6985 20060 6995
rect 20445 6995 20485 7005
rect 18335 6965 18375 6975
rect 18745 6965 18765 6985
rect 18895 6965 18915 6985
rect 19005 6965 19025 6985
rect 19115 6965 19135 6985
rect 19225 6965 19245 6985
rect 19335 6965 19355 6985
rect 19445 6965 19465 6985
rect 19555 6965 19575 6985
rect 19665 6965 19685 6985
rect 19775 6965 19795 6985
rect 19885 6965 19905 6985
rect 20035 6965 20055 6985
rect 20445 6975 20457 6995
rect 20475 6975 20485 6995
rect 20445 6965 20485 6975
rect 20555 6995 20595 7005
rect 20555 6975 20567 6995
rect 20585 6975 20595 6995
rect 20555 6965 20595 6975
rect 20665 6995 20705 7005
rect 20665 6975 20677 6995
rect 20695 6975 20705 6995
rect 20665 6965 20705 6975
rect 20775 6995 20815 7005
rect 20775 6975 20787 6995
rect 20805 6975 20815 6995
rect 20775 6965 20815 6975
rect 20885 6995 20925 7005
rect 20885 6975 20897 6995
rect 20915 6975 20925 6995
rect 20885 6965 20925 6975
rect 20995 6995 21035 7005
rect 20995 6975 21007 6995
rect 21025 6975 21035 6995
rect 20995 6965 21035 6975
rect 21105 6995 21145 7005
rect 21105 6975 21117 6995
rect 21135 6975 21145 6995
rect 21105 6965 21145 6975
rect 21215 6995 21255 7005
rect 21215 6975 21227 6995
rect 21245 6975 21255 6995
rect 21215 6965 21255 6975
rect 21325 6995 21365 7005
rect 21325 6975 21337 6995
rect 21355 6975 21365 6995
rect 21325 6965 21365 6975
rect 21435 6995 21475 7005
rect 21435 6975 21447 6995
rect 21465 6975 21475 6995
rect 21435 6965 21475 6975
rect 21545 6995 21585 7005
rect 21545 6975 21557 6995
rect 21575 6975 21585 6995
rect 21545 6965 21585 6975
rect 11235 6955 11275 6965
rect 11235 6935 11245 6955
rect 11265 6935 11275 6955
rect 11235 6925 11275 6935
rect 11385 6955 11425 6965
rect 11385 6935 11395 6955
rect 11415 6935 11425 6955
rect 11385 6925 11425 6935
rect 11495 6955 11535 6965
rect 11495 6935 11505 6955
rect 11525 6935 11535 6955
rect 11495 6925 11535 6935
rect 11605 6955 11645 6965
rect 11605 6935 11615 6955
rect 11635 6935 11645 6955
rect 11605 6925 11645 6935
rect 11715 6955 11755 6965
rect 11715 6935 11725 6955
rect 11745 6935 11755 6955
rect 11715 6925 11755 6935
rect 11825 6955 11865 6965
rect 11825 6935 11835 6955
rect 11855 6935 11865 6955
rect 11825 6925 11865 6935
rect 11935 6955 11975 6965
rect 11935 6935 11945 6955
rect 11965 6935 11975 6955
rect 11935 6925 11975 6935
rect 12045 6955 12085 6965
rect 12045 6935 12055 6955
rect 12075 6935 12085 6955
rect 12045 6925 12085 6935
rect 12155 6955 12195 6965
rect 12155 6935 12165 6955
rect 12185 6935 12195 6955
rect 12155 6925 12195 6935
rect 12265 6955 12305 6965
rect 12265 6935 12275 6955
rect 12295 6935 12305 6955
rect 12265 6925 12305 6935
rect 12375 6955 12415 6965
rect 12375 6935 12385 6955
rect 12405 6935 12415 6955
rect 12375 6925 12415 6935
rect 12525 6955 12565 6965
rect 12525 6935 12535 6955
rect 12555 6935 12565 6955
rect 12525 6925 12565 6935
rect 18735 6955 18775 6965
rect 18735 6935 18745 6955
rect 18765 6935 18775 6955
rect 18735 6925 18775 6935
rect 18885 6955 18925 6965
rect 18885 6935 18895 6955
rect 18915 6935 18925 6955
rect 18885 6925 18925 6935
rect 18995 6955 19035 6965
rect 18995 6935 19005 6955
rect 19025 6935 19035 6955
rect 18995 6925 19035 6935
rect 19105 6955 19145 6965
rect 19105 6935 19115 6955
rect 19135 6935 19145 6955
rect 19105 6925 19145 6935
rect 19215 6955 19255 6965
rect 19215 6935 19225 6955
rect 19245 6935 19255 6955
rect 19215 6925 19255 6935
rect 19325 6955 19365 6965
rect 19325 6935 19335 6955
rect 19355 6935 19365 6955
rect 19325 6925 19365 6935
rect 19435 6955 19475 6965
rect 19435 6935 19445 6955
rect 19465 6935 19475 6955
rect 19435 6925 19475 6935
rect 19545 6955 19585 6965
rect 19545 6935 19555 6955
rect 19575 6935 19585 6955
rect 19545 6925 19585 6935
rect 19655 6955 19695 6965
rect 19655 6935 19665 6955
rect 19685 6935 19695 6955
rect 19655 6925 19695 6935
rect 19765 6955 19805 6965
rect 19765 6935 19775 6955
rect 19795 6935 19805 6955
rect 19765 6925 19805 6935
rect 19875 6955 19915 6965
rect 19875 6935 19885 6955
rect 19905 6935 19915 6955
rect 19875 6925 19915 6935
rect 20025 6955 20065 6965
rect 20025 6935 20035 6955
rect 20055 6935 20065 6955
rect 20025 6925 20065 6935
rect 20450 6900 20490 6910
rect 20450 6880 20460 6900
rect 20480 6880 20490 6900
rect 20450 6870 20490 6880
rect 20545 6900 20585 6910
rect 20545 6880 20555 6900
rect 20575 6880 20585 6900
rect 20545 6870 20585 6880
rect 20655 6900 20695 6910
rect 20655 6880 20665 6900
rect 20685 6880 20695 6900
rect 20655 6870 20695 6880
rect 20765 6900 20805 6910
rect 20765 6880 20775 6900
rect 20795 6880 20805 6900
rect 20765 6870 20805 6880
rect 20860 6900 20900 6910
rect 20860 6880 20870 6900
rect 20890 6880 20900 6900
rect 20860 6870 20900 6880
rect 20460 6850 20480 6870
rect 20555 6850 20575 6870
rect 20665 6850 20685 6870
rect 20775 6850 20795 6870
rect 20870 6850 20890 6870
rect 20455 6840 20525 6850
rect 20455 6820 20460 6840
rect 20480 6820 20500 6840
rect 20520 6820 20525 6840
rect 20455 6790 20525 6820
rect 11190 6770 11230 6780
rect 11085 6755 11125 6765
rect 11085 6735 11095 6755
rect 11115 6735 11125 6755
rect 11190 6750 11200 6770
rect 11220 6750 11230 6770
rect 11410 6770 11450 6780
rect 11190 6740 11230 6750
rect 11305 6755 11345 6765
rect 11085 6725 11125 6735
rect 11095 6660 11115 6725
rect 11200 6660 11220 6740
rect 11305 6735 11315 6755
rect 11335 6735 11345 6755
rect 11410 6750 11420 6770
rect 11440 6750 11450 6770
rect 11640 6770 11680 6780
rect 11410 6740 11450 6750
rect 11525 6755 11565 6765
rect 11305 6725 11345 6735
rect 11237 6710 11269 6720
rect 11237 6690 11243 6710
rect 11260 6690 11269 6710
rect 11237 6680 11269 6690
rect 11315 6660 11335 6725
rect 11420 6660 11440 6740
rect 11525 6735 11535 6755
rect 11555 6735 11565 6755
rect 11640 6750 11650 6770
rect 11670 6750 11680 6770
rect 12230 6770 12270 6780
rect 11640 6740 11680 6750
rect 12125 6755 12165 6765
rect 11525 6725 11565 6735
rect 11457 6710 11489 6720
rect 11457 6690 11463 6710
rect 11480 6690 11489 6710
rect 11457 6680 11489 6690
rect 11535 6660 11555 6725
rect 11601 6710 11633 6720
rect 11601 6690 11610 6710
rect 11627 6690 11633 6710
rect 11601 6680 11633 6690
rect 11650 6660 11670 6740
rect 12125 6735 12135 6755
rect 12155 6735 12165 6755
rect 12230 6750 12240 6770
rect 12260 6750 12270 6770
rect 12450 6770 12490 6780
rect 12230 6740 12270 6750
rect 12345 6755 12385 6765
rect 12125 6725 12165 6735
rect 11820 6710 11850 6720
rect 11820 6690 11825 6710
rect 11845 6690 11850 6710
rect 11820 6680 11850 6690
rect 11867 6710 11899 6720
rect 11867 6690 11876 6710
rect 11893 6690 11899 6710
rect 11867 6680 11899 6690
rect 11950 6710 11980 6720
rect 11950 6690 11955 6710
rect 11975 6690 11980 6710
rect 11950 6680 11980 6690
rect 11830 6660 11850 6680
rect 11950 6660 11970 6680
rect 12135 6660 12155 6725
rect 12240 6660 12260 6740
rect 12345 6735 12355 6755
rect 12375 6735 12385 6755
rect 12450 6750 12460 6770
rect 12480 6750 12490 6770
rect 12680 6770 12720 6780
rect 12450 6740 12490 6750
rect 12565 6755 12605 6765
rect 12345 6725 12385 6735
rect 12277 6710 12309 6720
rect 12277 6690 12283 6710
rect 12300 6690 12309 6710
rect 12277 6680 12309 6690
rect 12355 6660 12375 6725
rect 12460 6660 12480 6740
rect 12565 6735 12575 6755
rect 12595 6735 12605 6755
rect 12680 6750 12690 6770
rect 12710 6750 12720 6770
rect 18690 6770 18730 6780
rect 12680 6740 12720 6750
rect 18585 6755 18625 6765
rect 12565 6725 12605 6735
rect 12497 6710 12529 6720
rect 12497 6690 12503 6710
rect 12520 6690 12529 6710
rect 12497 6680 12529 6690
rect 12575 6660 12595 6725
rect 12641 6710 12673 6720
rect 12641 6690 12650 6710
rect 12667 6690 12673 6710
rect 12641 6680 12673 6690
rect 12690 6660 12710 6740
rect 18585 6735 18595 6755
rect 18615 6735 18625 6755
rect 18690 6750 18700 6770
rect 18720 6750 18730 6770
rect 18910 6770 18950 6780
rect 18690 6740 18730 6750
rect 18805 6755 18845 6765
rect 18585 6725 18625 6735
rect 18595 6660 18615 6725
rect 18700 6660 18720 6740
rect 18805 6735 18815 6755
rect 18835 6735 18845 6755
rect 18910 6750 18920 6770
rect 18940 6750 18950 6770
rect 19140 6770 19180 6780
rect 18910 6740 18950 6750
rect 19025 6755 19065 6765
rect 18805 6725 18845 6735
rect 18737 6710 18769 6720
rect 18737 6690 18743 6710
rect 18760 6690 18769 6710
rect 18737 6680 18769 6690
rect 18815 6660 18835 6725
rect 18920 6660 18940 6740
rect 19025 6735 19035 6755
rect 19055 6735 19065 6755
rect 19140 6750 19150 6770
rect 19170 6750 19180 6770
rect 19730 6770 19770 6780
rect 19140 6740 19180 6750
rect 19625 6755 19665 6765
rect 19025 6725 19065 6735
rect 18957 6710 18989 6720
rect 18957 6690 18963 6710
rect 18980 6690 18989 6710
rect 18957 6680 18989 6690
rect 19035 6660 19055 6725
rect 19101 6710 19133 6720
rect 19101 6690 19110 6710
rect 19127 6690 19133 6710
rect 19101 6680 19133 6690
rect 19150 6660 19170 6740
rect 19625 6735 19635 6755
rect 19655 6735 19665 6755
rect 19730 6750 19740 6770
rect 19760 6750 19770 6770
rect 19950 6770 19990 6780
rect 19730 6740 19770 6750
rect 19845 6755 19885 6765
rect 19625 6725 19665 6735
rect 19320 6710 19350 6720
rect 19320 6690 19325 6710
rect 19345 6690 19350 6710
rect 19320 6680 19350 6690
rect 19367 6710 19399 6720
rect 19367 6690 19376 6710
rect 19393 6690 19399 6710
rect 19367 6680 19399 6690
rect 19450 6710 19480 6720
rect 19450 6690 19455 6710
rect 19475 6690 19480 6710
rect 19450 6680 19480 6690
rect 19330 6660 19350 6680
rect 19450 6660 19470 6680
rect 19635 6660 19655 6725
rect 19740 6660 19760 6740
rect 19845 6735 19855 6755
rect 19875 6735 19885 6755
rect 19950 6750 19960 6770
rect 19980 6750 19990 6770
rect 20180 6770 20220 6780
rect 19950 6740 19990 6750
rect 20065 6755 20105 6765
rect 19845 6725 19885 6735
rect 19777 6710 19809 6720
rect 19777 6690 19783 6710
rect 19800 6690 19809 6710
rect 19777 6680 19809 6690
rect 19855 6660 19875 6725
rect 19960 6660 19980 6740
rect 20065 6735 20075 6755
rect 20095 6735 20105 6755
rect 20180 6750 20190 6770
rect 20210 6750 20220 6770
rect 20180 6740 20220 6750
rect 20455 6770 20460 6790
rect 20480 6770 20500 6790
rect 20520 6770 20525 6790
rect 20455 6740 20525 6770
rect 20065 6725 20105 6735
rect 19997 6710 20029 6720
rect 19997 6690 20003 6710
rect 20020 6690 20029 6710
rect 19997 6680 20029 6690
rect 20075 6660 20095 6725
rect 20141 6710 20173 6720
rect 20141 6690 20150 6710
rect 20167 6690 20173 6710
rect 20141 6680 20173 6690
rect 20190 6660 20210 6740
rect 20455 6720 20460 6740
rect 20480 6720 20500 6740
rect 20520 6720 20525 6740
rect 20455 6710 20525 6720
rect 20550 6840 20580 6850
rect 20550 6820 20555 6840
rect 20575 6820 20580 6840
rect 20550 6790 20580 6820
rect 20550 6770 20555 6790
rect 20575 6770 20580 6790
rect 20550 6740 20580 6770
rect 20550 6720 20555 6740
rect 20575 6720 20580 6740
rect 20550 6710 20580 6720
rect 20605 6840 20635 6850
rect 20605 6820 20610 6840
rect 20630 6820 20635 6840
rect 20605 6790 20635 6820
rect 20605 6770 20610 6790
rect 20630 6770 20635 6790
rect 20605 6740 20635 6770
rect 20605 6720 20610 6740
rect 20630 6720 20635 6740
rect 20605 6710 20635 6720
rect 20660 6840 20690 6850
rect 20660 6820 20665 6840
rect 20685 6820 20690 6840
rect 20660 6790 20690 6820
rect 20660 6770 20665 6790
rect 20685 6770 20690 6790
rect 20660 6740 20690 6770
rect 20660 6720 20665 6740
rect 20685 6720 20690 6740
rect 20660 6710 20690 6720
rect 20715 6840 20745 6850
rect 20715 6820 20720 6840
rect 20740 6820 20745 6840
rect 20715 6790 20745 6820
rect 20715 6770 20720 6790
rect 20740 6770 20745 6790
rect 20715 6740 20745 6770
rect 20715 6720 20720 6740
rect 20740 6720 20745 6740
rect 20715 6710 20745 6720
rect 20770 6840 20800 6850
rect 20770 6820 20775 6840
rect 20795 6820 20800 6840
rect 20770 6790 20800 6820
rect 20770 6770 20775 6790
rect 20795 6770 20800 6790
rect 20770 6740 20800 6770
rect 20770 6720 20775 6740
rect 20795 6720 20800 6740
rect 20770 6710 20800 6720
rect 20825 6840 20895 6850
rect 20825 6820 20830 6840
rect 20850 6820 20870 6840
rect 20890 6820 20895 6840
rect 20825 6790 20895 6820
rect 20825 6770 20830 6790
rect 20850 6770 20870 6790
rect 20890 6770 20895 6790
rect 20825 6740 20895 6770
rect 20825 6720 20830 6740
rect 20850 6720 20870 6740
rect 20890 6720 20895 6740
rect 20825 6710 20895 6720
rect 20615 6690 20635 6710
rect 20720 6690 20740 6710
rect 20566 6675 20598 6685
rect 10990 6650 11065 6660
rect 10990 6630 11000 6650
rect 11020 6630 11040 6650
rect 11060 6630 11065 6650
rect 10990 6600 11065 6630
rect 10990 6580 11000 6600
rect 11020 6580 11040 6600
rect 11060 6580 11065 6600
rect 10990 6550 11065 6580
rect 10990 6530 11000 6550
rect 11020 6530 11040 6550
rect 11060 6530 11065 6550
rect 10990 6520 11065 6530
rect 11090 6650 11120 6660
rect 11090 6630 11095 6650
rect 11115 6630 11120 6650
rect 11090 6600 11120 6630
rect 11090 6580 11095 6600
rect 11115 6580 11120 6600
rect 11090 6550 11120 6580
rect 11090 6530 11095 6550
rect 11115 6530 11120 6550
rect 11090 6520 11120 6530
rect 11145 6650 11175 6660
rect 11145 6630 11150 6650
rect 11170 6630 11175 6650
rect 11145 6600 11175 6630
rect 11145 6580 11150 6600
rect 11170 6580 11175 6600
rect 11145 6550 11175 6580
rect 11145 6530 11150 6550
rect 11170 6530 11175 6550
rect 11145 6520 11175 6530
rect 11200 6650 11230 6660
rect 11200 6630 11205 6650
rect 11225 6630 11230 6650
rect 11200 6600 11230 6630
rect 11200 6580 11205 6600
rect 11225 6580 11230 6600
rect 11200 6550 11230 6580
rect 11200 6530 11205 6550
rect 11225 6530 11230 6550
rect 11200 6520 11230 6530
rect 11255 6650 11285 6660
rect 11255 6630 11260 6650
rect 11280 6630 11285 6650
rect 11255 6600 11285 6630
rect 11255 6580 11260 6600
rect 11280 6580 11285 6600
rect 11255 6550 11285 6580
rect 11255 6530 11260 6550
rect 11280 6530 11285 6550
rect 11255 6520 11285 6530
rect 11310 6650 11340 6660
rect 11310 6630 11315 6650
rect 11335 6630 11340 6650
rect 11310 6600 11340 6630
rect 11310 6580 11315 6600
rect 11335 6580 11340 6600
rect 11310 6550 11340 6580
rect 11310 6530 11315 6550
rect 11335 6530 11340 6550
rect 11310 6520 11340 6530
rect 11365 6650 11395 6660
rect 11365 6630 11370 6650
rect 11390 6630 11395 6650
rect 11365 6600 11395 6630
rect 11365 6580 11370 6600
rect 11390 6580 11395 6600
rect 11365 6550 11395 6580
rect 11365 6530 11370 6550
rect 11390 6530 11395 6550
rect 11365 6520 11395 6530
rect 11420 6650 11450 6660
rect 11420 6630 11425 6650
rect 11445 6630 11450 6650
rect 11420 6600 11450 6630
rect 11420 6580 11425 6600
rect 11445 6580 11450 6600
rect 11420 6550 11450 6580
rect 11420 6530 11425 6550
rect 11445 6530 11450 6550
rect 11420 6520 11450 6530
rect 11475 6650 11505 6660
rect 11475 6630 11480 6650
rect 11500 6630 11505 6650
rect 11475 6600 11505 6630
rect 11475 6580 11480 6600
rect 11500 6580 11505 6600
rect 11475 6550 11505 6580
rect 11475 6530 11480 6550
rect 11500 6530 11505 6550
rect 11475 6520 11505 6530
rect 11530 6650 11560 6660
rect 11530 6630 11535 6650
rect 11555 6630 11560 6650
rect 11530 6600 11560 6630
rect 11530 6580 11535 6600
rect 11555 6580 11560 6600
rect 11530 6550 11560 6580
rect 11530 6530 11535 6550
rect 11555 6530 11560 6550
rect 11530 6520 11560 6530
rect 11585 6650 11615 6660
rect 11585 6630 11590 6650
rect 11610 6630 11615 6650
rect 11585 6600 11615 6630
rect 11585 6580 11590 6600
rect 11610 6580 11615 6600
rect 11585 6550 11615 6580
rect 11585 6530 11590 6550
rect 11610 6530 11615 6550
rect 11585 6520 11615 6530
rect 11640 6650 11670 6660
rect 11640 6630 11645 6650
rect 11665 6630 11670 6650
rect 11640 6600 11670 6630
rect 11640 6580 11645 6600
rect 11665 6580 11670 6600
rect 11640 6550 11670 6580
rect 11640 6530 11645 6550
rect 11665 6530 11670 6550
rect 11640 6520 11670 6530
rect 11695 6650 11805 6660
rect 11695 6630 11700 6650
rect 11720 6630 11740 6650
rect 11760 6630 11780 6650
rect 11800 6630 11805 6650
rect 11695 6600 11805 6630
rect 11695 6580 11700 6600
rect 11720 6580 11740 6600
rect 11760 6580 11780 6600
rect 11800 6580 11805 6600
rect 11695 6550 11805 6580
rect 11695 6530 11700 6550
rect 11720 6530 11740 6550
rect 11760 6530 11780 6550
rect 11800 6530 11805 6550
rect 11695 6520 11805 6530
rect 11830 6650 11860 6660
rect 11830 6630 11835 6650
rect 11855 6630 11860 6650
rect 11830 6600 11860 6630
rect 11830 6580 11835 6600
rect 11855 6580 11860 6600
rect 11830 6550 11860 6580
rect 11830 6530 11835 6550
rect 11855 6530 11860 6550
rect 11830 6520 11860 6530
rect 11885 6650 11915 6660
rect 11885 6630 11890 6650
rect 11910 6630 11915 6650
rect 11885 6600 11915 6630
rect 11885 6580 11890 6600
rect 11910 6580 11915 6600
rect 11885 6550 11915 6580
rect 11885 6530 11890 6550
rect 11910 6530 11915 6550
rect 11885 6520 11915 6530
rect 11940 6650 11970 6660
rect 11940 6630 11945 6650
rect 11965 6630 11970 6650
rect 11940 6600 11970 6630
rect 11940 6580 11945 6600
rect 11965 6580 11970 6600
rect 11940 6550 11970 6580
rect 11940 6530 11945 6550
rect 11965 6530 11970 6550
rect 11940 6520 11970 6530
rect 11995 6650 12105 6660
rect 11995 6630 12000 6650
rect 12020 6630 12040 6650
rect 12060 6630 12080 6650
rect 12100 6630 12105 6650
rect 11995 6600 12105 6630
rect 11995 6580 12000 6600
rect 12020 6580 12040 6600
rect 12060 6580 12080 6600
rect 12100 6580 12105 6600
rect 11995 6550 12105 6580
rect 11995 6530 12000 6550
rect 12020 6530 12040 6550
rect 12060 6530 12080 6550
rect 12100 6530 12105 6550
rect 11995 6520 12105 6530
rect 12130 6650 12160 6660
rect 12130 6630 12135 6650
rect 12155 6630 12160 6650
rect 12130 6600 12160 6630
rect 12130 6580 12135 6600
rect 12155 6580 12160 6600
rect 12130 6550 12160 6580
rect 12130 6530 12135 6550
rect 12155 6530 12160 6550
rect 12130 6520 12160 6530
rect 12185 6650 12215 6660
rect 12185 6630 12190 6650
rect 12210 6630 12215 6650
rect 12185 6600 12215 6630
rect 12185 6580 12190 6600
rect 12210 6580 12215 6600
rect 12185 6550 12215 6580
rect 12185 6530 12190 6550
rect 12210 6530 12215 6550
rect 12185 6520 12215 6530
rect 12240 6650 12270 6660
rect 12240 6630 12245 6650
rect 12265 6630 12270 6650
rect 12240 6600 12270 6630
rect 12240 6580 12245 6600
rect 12265 6580 12270 6600
rect 12240 6550 12270 6580
rect 12240 6530 12245 6550
rect 12265 6530 12270 6550
rect 12240 6520 12270 6530
rect 12295 6650 12325 6660
rect 12295 6630 12300 6650
rect 12320 6630 12325 6650
rect 12295 6600 12325 6630
rect 12295 6580 12300 6600
rect 12320 6580 12325 6600
rect 12295 6550 12325 6580
rect 12295 6530 12300 6550
rect 12320 6530 12325 6550
rect 12295 6520 12325 6530
rect 12350 6650 12380 6660
rect 12350 6630 12355 6650
rect 12375 6630 12380 6650
rect 12350 6600 12380 6630
rect 12350 6580 12355 6600
rect 12375 6580 12380 6600
rect 12350 6550 12380 6580
rect 12350 6530 12355 6550
rect 12375 6530 12380 6550
rect 12350 6520 12380 6530
rect 12405 6650 12435 6660
rect 12405 6630 12410 6650
rect 12430 6630 12435 6650
rect 12405 6600 12435 6630
rect 12405 6580 12410 6600
rect 12430 6580 12435 6600
rect 12405 6550 12435 6580
rect 12405 6530 12410 6550
rect 12430 6530 12435 6550
rect 12405 6520 12435 6530
rect 12460 6650 12490 6660
rect 12460 6630 12465 6650
rect 12485 6630 12490 6650
rect 12460 6600 12490 6630
rect 12460 6580 12465 6600
rect 12485 6580 12490 6600
rect 12460 6550 12490 6580
rect 12460 6530 12465 6550
rect 12485 6530 12490 6550
rect 12460 6520 12490 6530
rect 12515 6650 12545 6660
rect 12515 6630 12520 6650
rect 12540 6630 12545 6650
rect 12515 6600 12545 6630
rect 12515 6580 12520 6600
rect 12540 6580 12545 6600
rect 12515 6550 12545 6580
rect 12515 6530 12520 6550
rect 12540 6530 12545 6550
rect 12515 6520 12545 6530
rect 12570 6650 12600 6660
rect 12570 6630 12575 6650
rect 12595 6630 12600 6650
rect 12570 6600 12600 6630
rect 12570 6580 12575 6600
rect 12595 6580 12600 6600
rect 12570 6550 12600 6580
rect 12570 6530 12575 6550
rect 12595 6530 12600 6550
rect 12570 6520 12600 6530
rect 12625 6650 12655 6660
rect 12625 6630 12630 6650
rect 12650 6630 12655 6650
rect 12625 6600 12655 6630
rect 12625 6580 12630 6600
rect 12650 6580 12655 6600
rect 12625 6550 12655 6580
rect 12625 6530 12630 6550
rect 12650 6530 12655 6550
rect 12625 6520 12655 6530
rect 12680 6650 12710 6660
rect 12680 6630 12685 6650
rect 12705 6630 12710 6650
rect 12680 6600 12710 6630
rect 12680 6580 12685 6600
rect 12705 6580 12710 6600
rect 12680 6550 12710 6580
rect 12680 6530 12685 6550
rect 12705 6530 12710 6550
rect 12680 6520 12710 6530
rect 12735 6650 12810 6660
rect 12735 6630 12740 6650
rect 12760 6630 12780 6650
rect 12800 6630 12810 6650
rect 12735 6600 12810 6630
rect 12735 6580 12740 6600
rect 12760 6580 12780 6600
rect 12800 6580 12810 6600
rect 12735 6550 12810 6580
rect 12735 6530 12740 6550
rect 12760 6530 12780 6550
rect 12800 6530 12810 6550
rect 12735 6520 12810 6530
rect 18490 6650 18565 6660
rect 18490 6630 18500 6650
rect 18520 6630 18540 6650
rect 18560 6630 18565 6650
rect 18490 6600 18565 6630
rect 18490 6580 18500 6600
rect 18520 6580 18540 6600
rect 18560 6580 18565 6600
rect 18490 6550 18565 6580
rect 18490 6530 18500 6550
rect 18520 6530 18540 6550
rect 18560 6530 18565 6550
rect 18490 6520 18565 6530
rect 18590 6650 18620 6660
rect 18590 6630 18595 6650
rect 18615 6630 18620 6650
rect 18590 6600 18620 6630
rect 18590 6580 18595 6600
rect 18615 6580 18620 6600
rect 18590 6550 18620 6580
rect 18590 6530 18595 6550
rect 18615 6530 18620 6550
rect 18590 6520 18620 6530
rect 18645 6650 18675 6660
rect 18645 6630 18650 6650
rect 18670 6630 18675 6650
rect 18645 6600 18675 6630
rect 18645 6580 18650 6600
rect 18670 6580 18675 6600
rect 18645 6550 18675 6580
rect 18645 6530 18650 6550
rect 18670 6530 18675 6550
rect 18645 6520 18675 6530
rect 18700 6650 18730 6660
rect 18700 6630 18705 6650
rect 18725 6630 18730 6650
rect 18700 6600 18730 6630
rect 18700 6580 18705 6600
rect 18725 6580 18730 6600
rect 18700 6550 18730 6580
rect 18700 6530 18705 6550
rect 18725 6530 18730 6550
rect 18700 6520 18730 6530
rect 18755 6650 18785 6660
rect 18755 6630 18760 6650
rect 18780 6630 18785 6650
rect 18755 6600 18785 6630
rect 18755 6580 18760 6600
rect 18780 6580 18785 6600
rect 18755 6550 18785 6580
rect 18755 6530 18760 6550
rect 18780 6530 18785 6550
rect 18755 6520 18785 6530
rect 18810 6650 18840 6660
rect 18810 6630 18815 6650
rect 18835 6630 18840 6650
rect 18810 6600 18840 6630
rect 18810 6580 18815 6600
rect 18835 6580 18840 6600
rect 18810 6550 18840 6580
rect 18810 6530 18815 6550
rect 18835 6530 18840 6550
rect 18810 6520 18840 6530
rect 18865 6650 18895 6660
rect 18865 6630 18870 6650
rect 18890 6630 18895 6650
rect 18865 6600 18895 6630
rect 18865 6580 18870 6600
rect 18890 6580 18895 6600
rect 18865 6550 18895 6580
rect 18865 6530 18870 6550
rect 18890 6530 18895 6550
rect 18865 6520 18895 6530
rect 18920 6650 18950 6660
rect 18920 6630 18925 6650
rect 18945 6630 18950 6650
rect 18920 6600 18950 6630
rect 18920 6580 18925 6600
rect 18945 6580 18950 6600
rect 18920 6550 18950 6580
rect 18920 6530 18925 6550
rect 18945 6530 18950 6550
rect 18920 6520 18950 6530
rect 18975 6650 19005 6660
rect 18975 6630 18980 6650
rect 19000 6630 19005 6650
rect 18975 6600 19005 6630
rect 18975 6580 18980 6600
rect 19000 6580 19005 6600
rect 18975 6550 19005 6580
rect 18975 6530 18980 6550
rect 19000 6530 19005 6550
rect 18975 6520 19005 6530
rect 19030 6650 19060 6660
rect 19030 6630 19035 6650
rect 19055 6630 19060 6650
rect 19030 6600 19060 6630
rect 19030 6580 19035 6600
rect 19055 6580 19060 6600
rect 19030 6550 19060 6580
rect 19030 6530 19035 6550
rect 19055 6530 19060 6550
rect 19030 6520 19060 6530
rect 19085 6650 19115 6660
rect 19085 6630 19090 6650
rect 19110 6630 19115 6650
rect 19085 6600 19115 6630
rect 19085 6580 19090 6600
rect 19110 6580 19115 6600
rect 19085 6550 19115 6580
rect 19085 6530 19090 6550
rect 19110 6530 19115 6550
rect 19085 6520 19115 6530
rect 19140 6650 19170 6660
rect 19140 6630 19145 6650
rect 19165 6630 19170 6650
rect 19140 6600 19170 6630
rect 19140 6580 19145 6600
rect 19165 6580 19170 6600
rect 19140 6550 19170 6580
rect 19140 6530 19145 6550
rect 19165 6530 19170 6550
rect 19140 6520 19170 6530
rect 19195 6650 19305 6660
rect 19195 6630 19200 6650
rect 19220 6630 19240 6650
rect 19260 6630 19280 6650
rect 19300 6630 19305 6650
rect 19195 6600 19305 6630
rect 19195 6580 19200 6600
rect 19220 6580 19240 6600
rect 19260 6580 19280 6600
rect 19300 6580 19305 6600
rect 19195 6550 19305 6580
rect 19195 6530 19200 6550
rect 19220 6530 19240 6550
rect 19260 6530 19280 6550
rect 19300 6530 19305 6550
rect 19195 6520 19305 6530
rect 19330 6650 19360 6660
rect 19330 6630 19335 6650
rect 19355 6630 19360 6650
rect 19330 6600 19360 6630
rect 19330 6580 19335 6600
rect 19355 6580 19360 6600
rect 19330 6550 19360 6580
rect 19330 6530 19335 6550
rect 19355 6530 19360 6550
rect 19330 6520 19360 6530
rect 19385 6650 19415 6660
rect 19385 6630 19390 6650
rect 19410 6630 19415 6650
rect 19385 6600 19415 6630
rect 19385 6580 19390 6600
rect 19410 6580 19415 6600
rect 19385 6550 19415 6580
rect 19385 6530 19390 6550
rect 19410 6530 19415 6550
rect 19385 6520 19415 6530
rect 19440 6650 19470 6660
rect 19440 6630 19445 6650
rect 19465 6630 19470 6650
rect 19440 6600 19470 6630
rect 19440 6580 19445 6600
rect 19465 6580 19470 6600
rect 19440 6550 19470 6580
rect 19440 6530 19445 6550
rect 19465 6530 19470 6550
rect 19440 6520 19470 6530
rect 19495 6650 19605 6660
rect 19495 6630 19500 6650
rect 19520 6630 19540 6650
rect 19560 6630 19580 6650
rect 19600 6630 19605 6650
rect 19495 6600 19605 6630
rect 19495 6580 19500 6600
rect 19520 6580 19540 6600
rect 19560 6580 19580 6600
rect 19600 6580 19605 6600
rect 19495 6550 19605 6580
rect 19495 6530 19500 6550
rect 19520 6530 19540 6550
rect 19560 6530 19580 6550
rect 19600 6530 19605 6550
rect 19495 6520 19605 6530
rect 19630 6650 19660 6660
rect 19630 6630 19635 6650
rect 19655 6630 19660 6650
rect 19630 6600 19660 6630
rect 19630 6580 19635 6600
rect 19655 6580 19660 6600
rect 19630 6550 19660 6580
rect 19630 6530 19635 6550
rect 19655 6530 19660 6550
rect 19630 6520 19660 6530
rect 19685 6650 19715 6660
rect 19685 6630 19690 6650
rect 19710 6630 19715 6650
rect 19685 6600 19715 6630
rect 19685 6580 19690 6600
rect 19710 6580 19715 6600
rect 19685 6550 19715 6580
rect 19685 6530 19690 6550
rect 19710 6530 19715 6550
rect 19685 6520 19715 6530
rect 19740 6650 19770 6660
rect 19740 6630 19745 6650
rect 19765 6630 19770 6650
rect 19740 6600 19770 6630
rect 19740 6580 19745 6600
rect 19765 6580 19770 6600
rect 19740 6550 19770 6580
rect 19740 6530 19745 6550
rect 19765 6530 19770 6550
rect 19740 6520 19770 6530
rect 19795 6650 19825 6660
rect 19795 6630 19800 6650
rect 19820 6630 19825 6650
rect 19795 6600 19825 6630
rect 19795 6580 19800 6600
rect 19820 6580 19825 6600
rect 19795 6550 19825 6580
rect 19795 6530 19800 6550
rect 19820 6530 19825 6550
rect 19795 6520 19825 6530
rect 19850 6650 19880 6660
rect 19850 6630 19855 6650
rect 19875 6630 19880 6650
rect 19850 6600 19880 6630
rect 19850 6580 19855 6600
rect 19875 6580 19880 6600
rect 19850 6550 19880 6580
rect 19850 6530 19855 6550
rect 19875 6530 19880 6550
rect 19850 6520 19880 6530
rect 19905 6650 19935 6660
rect 19905 6630 19910 6650
rect 19930 6630 19935 6650
rect 19905 6600 19935 6630
rect 19905 6580 19910 6600
rect 19930 6580 19935 6600
rect 19905 6550 19935 6580
rect 19905 6530 19910 6550
rect 19930 6530 19935 6550
rect 19905 6520 19935 6530
rect 19960 6650 19990 6660
rect 19960 6630 19965 6650
rect 19985 6630 19990 6650
rect 19960 6600 19990 6630
rect 19960 6580 19965 6600
rect 19985 6580 19990 6600
rect 19960 6550 19990 6580
rect 19960 6530 19965 6550
rect 19985 6530 19990 6550
rect 19960 6520 19990 6530
rect 20015 6650 20045 6660
rect 20015 6630 20020 6650
rect 20040 6630 20045 6650
rect 20015 6600 20045 6630
rect 20015 6580 20020 6600
rect 20040 6580 20045 6600
rect 20015 6550 20045 6580
rect 20015 6530 20020 6550
rect 20040 6530 20045 6550
rect 20015 6520 20045 6530
rect 20070 6650 20100 6660
rect 20070 6630 20075 6650
rect 20095 6630 20100 6650
rect 20070 6600 20100 6630
rect 20070 6580 20075 6600
rect 20095 6580 20100 6600
rect 20070 6550 20100 6580
rect 20070 6530 20075 6550
rect 20095 6530 20100 6550
rect 20070 6520 20100 6530
rect 20125 6650 20155 6660
rect 20125 6630 20130 6650
rect 20150 6630 20155 6650
rect 20125 6600 20155 6630
rect 20125 6580 20130 6600
rect 20150 6580 20155 6600
rect 20125 6550 20155 6580
rect 20125 6530 20130 6550
rect 20150 6530 20155 6550
rect 20125 6520 20155 6530
rect 20180 6650 20210 6660
rect 20180 6630 20185 6650
rect 20205 6630 20210 6650
rect 20180 6600 20210 6630
rect 20180 6580 20185 6600
rect 20205 6580 20210 6600
rect 20180 6550 20210 6580
rect 20180 6530 20185 6550
rect 20205 6530 20210 6550
rect 20180 6520 20210 6530
rect 20235 6650 20310 6660
rect 20235 6630 20240 6650
rect 20260 6630 20280 6650
rect 20300 6630 20310 6650
rect 20566 6655 20571 6675
rect 20591 6655 20598 6675
rect 20566 6645 20598 6655
rect 20615 6680 20655 6690
rect 20615 6660 20625 6680
rect 20645 6660 20655 6680
rect 20615 6650 20655 6660
rect 20710 6680 20750 6690
rect 20710 6660 20720 6680
rect 20740 6660 20750 6680
rect 20710 6650 20750 6660
rect 20235 6600 20310 6630
rect 20235 6580 20240 6600
rect 20260 6580 20280 6600
rect 20300 6580 20310 6600
rect 20510 6625 20550 6635
rect 20510 6605 20520 6625
rect 20540 6605 20550 6625
rect 20510 6595 20550 6605
rect 20800 6625 20840 6635
rect 20800 6605 20810 6625
rect 20830 6605 20840 6625
rect 20800 6595 20840 6605
rect 20235 6550 20310 6580
rect 20235 6530 20240 6550
rect 20260 6530 20280 6550
rect 20300 6530 20310 6550
rect 20471 6565 20503 6575
rect 20471 6545 20476 6565
rect 20496 6545 20503 6565
rect 20471 6535 20503 6545
rect 20235 6520 20310 6530
rect 11000 6500 11020 6520
rect 10990 6490 11030 6500
rect 10990 6470 11000 6490
rect 11020 6470 11030 6490
rect 10990 6460 11030 6470
rect 11106 6490 11138 6500
rect 11106 6470 11112 6490
rect 11129 6470 11138 6490
rect 11106 6460 11138 6470
rect 9760 6440 9805 6445
rect 9760 6415 9770 6440
rect 9795 6415 9805 6440
rect 9760 6410 9805 6415
rect 10770 6440 10815 6445
rect 11155 6440 11175 6520
rect 11260 6440 11280 6520
rect 11305 6490 11345 6500
rect 11305 6470 11315 6490
rect 11335 6470 11345 6490
rect 11305 6460 11345 6470
rect 11370 6440 11390 6520
rect 11480 6440 11500 6520
rect 11525 6490 11565 6500
rect 11525 6470 11535 6490
rect 11555 6470 11565 6490
rect 11525 6460 11565 6470
rect 11590 6440 11610 6520
rect 11740 6500 11760 6520
rect 11830 6500 11850 6520
rect 11885 6500 11905 6520
rect 12040 6500 12060 6520
rect 11730 6490 11770 6500
rect 11730 6470 11740 6490
rect 11760 6470 11770 6490
rect 11730 6460 11770 6470
rect 11825 6490 11855 6500
rect 11825 6470 11830 6490
rect 11850 6470 11855 6490
rect 11825 6460 11855 6470
rect 11875 6490 11905 6500
rect 11875 6470 11880 6490
rect 11900 6470 11905 6490
rect 11875 6460 11905 6470
rect 11922 6490 11954 6500
rect 11922 6470 11928 6490
rect 11945 6470 11954 6490
rect 11922 6460 11954 6470
rect 12030 6490 12070 6500
rect 12030 6470 12040 6490
rect 12060 6470 12070 6490
rect 12030 6460 12070 6470
rect 12146 6490 12178 6500
rect 12146 6470 12152 6490
rect 12169 6470 12178 6490
rect 12146 6460 12178 6470
rect 12195 6440 12215 6520
rect 12300 6440 12320 6520
rect 12345 6490 12385 6500
rect 12345 6470 12355 6490
rect 12375 6470 12385 6490
rect 12345 6460 12385 6470
rect 12410 6440 12430 6520
rect 12520 6440 12540 6520
rect 12565 6490 12605 6500
rect 12565 6470 12575 6490
rect 12595 6470 12605 6490
rect 12565 6460 12605 6470
rect 12630 6440 12650 6520
rect 12780 6500 12800 6520
rect 18500 6500 18520 6520
rect 12770 6490 12810 6500
rect 12770 6470 12780 6490
rect 12800 6470 12810 6490
rect 12770 6460 12810 6470
rect 18490 6490 18530 6500
rect 18490 6470 18500 6490
rect 18520 6470 18530 6490
rect 18490 6460 18530 6470
rect 18606 6490 18638 6500
rect 18606 6470 18612 6490
rect 18629 6470 18638 6490
rect 18606 6460 18638 6470
rect 12985 6440 13030 6445
rect 10770 6415 10780 6440
rect 10805 6415 10815 6440
rect 10770 6410 10815 6415
rect 11145 6430 11185 6440
rect 11145 6410 11155 6430
rect 11175 6410 11185 6430
rect 11145 6400 11185 6410
rect 11250 6430 11290 6440
rect 11250 6410 11260 6430
rect 11280 6410 11290 6430
rect 11250 6400 11290 6410
rect 11360 6430 11400 6440
rect 11360 6410 11370 6430
rect 11390 6410 11400 6430
rect 11360 6400 11400 6410
rect 11470 6430 11510 6440
rect 11470 6410 11480 6430
rect 11500 6410 11510 6430
rect 11470 6400 11510 6410
rect 11580 6430 11620 6440
rect 11580 6410 11590 6430
rect 11610 6410 11620 6430
rect 11580 6400 11620 6410
rect 12185 6430 12225 6440
rect 12185 6410 12195 6430
rect 12215 6410 12225 6430
rect 12185 6400 12225 6410
rect 12290 6430 12330 6440
rect 12290 6410 12300 6430
rect 12320 6410 12330 6430
rect 12290 6400 12330 6410
rect 12400 6430 12440 6440
rect 12400 6410 12410 6430
rect 12430 6410 12440 6430
rect 12400 6400 12440 6410
rect 12510 6430 12550 6440
rect 12510 6410 12520 6430
rect 12540 6410 12550 6430
rect 12510 6400 12550 6410
rect 12620 6430 12660 6440
rect 12620 6410 12630 6430
rect 12650 6410 12660 6430
rect 12985 6415 12995 6440
rect 13020 6415 13030 6440
rect 12985 6410 13030 6415
rect 13995 6440 14040 6445
rect 18655 6440 18675 6520
rect 18760 6440 18780 6520
rect 18805 6490 18845 6500
rect 18805 6470 18815 6490
rect 18835 6470 18845 6490
rect 18805 6460 18845 6470
rect 18870 6440 18890 6520
rect 18980 6440 19000 6520
rect 19025 6490 19065 6500
rect 19025 6470 19035 6490
rect 19055 6470 19065 6490
rect 19025 6460 19065 6470
rect 19090 6440 19110 6520
rect 19240 6500 19260 6520
rect 19330 6500 19350 6520
rect 19385 6500 19405 6520
rect 19540 6500 19560 6520
rect 19230 6490 19270 6500
rect 19230 6470 19240 6490
rect 19260 6470 19270 6490
rect 19230 6460 19270 6470
rect 19325 6490 19355 6500
rect 19325 6470 19330 6490
rect 19350 6470 19355 6490
rect 19325 6460 19355 6470
rect 19375 6490 19405 6500
rect 19375 6470 19380 6490
rect 19400 6470 19405 6490
rect 19375 6460 19405 6470
rect 19422 6490 19454 6500
rect 19422 6470 19428 6490
rect 19445 6470 19454 6490
rect 19422 6460 19454 6470
rect 19530 6490 19570 6500
rect 19530 6470 19540 6490
rect 19560 6470 19570 6490
rect 19530 6460 19570 6470
rect 19646 6490 19678 6500
rect 19646 6470 19652 6490
rect 19669 6470 19678 6490
rect 19646 6460 19678 6470
rect 19695 6440 19715 6520
rect 19800 6440 19820 6520
rect 19845 6490 19885 6500
rect 19845 6470 19855 6490
rect 19875 6470 19885 6490
rect 19845 6460 19885 6470
rect 19910 6440 19930 6520
rect 20020 6440 20040 6520
rect 20065 6490 20105 6500
rect 20065 6470 20075 6490
rect 20095 6470 20105 6490
rect 20065 6460 20105 6470
rect 20130 6440 20150 6520
rect 20280 6500 20300 6520
rect 20520 6515 20540 6595
rect 20560 6565 20600 6575
rect 20560 6545 20570 6565
rect 20590 6545 20600 6565
rect 20560 6535 20600 6545
rect 20570 6515 20590 6535
rect 20810 6515 20830 6595
rect 20847 6565 20879 6575
rect 20847 6545 20854 6565
rect 20874 6545 20879 6565
rect 20847 6535 20879 6545
rect 20355 6505 20430 6515
rect 20270 6490 20310 6500
rect 20270 6470 20280 6490
rect 20300 6470 20310 6490
rect 20270 6460 20310 6470
rect 20355 6485 20365 6505
rect 20385 6485 20405 6505
rect 20425 6485 20430 6505
rect 20355 6455 20430 6485
rect 13995 6415 14005 6440
rect 14030 6415 14040 6440
rect 13995 6410 14040 6415
rect 18645 6430 18685 6440
rect 18645 6410 18655 6430
rect 18675 6410 18685 6430
rect 12620 6400 12660 6410
rect 18645 6400 18685 6410
rect 18750 6430 18790 6440
rect 18750 6410 18760 6430
rect 18780 6410 18790 6430
rect 18750 6400 18790 6410
rect 18860 6430 18900 6440
rect 18860 6410 18870 6430
rect 18890 6410 18900 6430
rect 18860 6400 18900 6410
rect 18970 6430 19010 6440
rect 18970 6410 18980 6430
rect 19000 6410 19010 6430
rect 18970 6400 19010 6410
rect 19080 6430 19120 6440
rect 19080 6410 19090 6430
rect 19110 6410 19120 6430
rect 19080 6400 19120 6410
rect 19685 6430 19725 6440
rect 19685 6410 19695 6430
rect 19715 6410 19725 6430
rect 19685 6400 19725 6410
rect 19790 6430 19830 6440
rect 19790 6410 19800 6430
rect 19820 6410 19830 6430
rect 19790 6400 19830 6410
rect 19900 6430 19940 6440
rect 19900 6410 19910 6430
rect 19930 6410 19940 6430
rect 19900 6400 19940 6410
rect 20010 6430 20050 6440
rect 20010 6410 20020 6430
rect 20040 6410 20050 6430
rect 20010 6400 20050 6410
rect 20120 6430 20160 6440
rect 20120 6410 20130 6430
rect 20150 6410 20160 6430
rect 20120 6400 20160 6410
rect 20355 6435 20365 6455
rect 20385 6435 20405 6455
rect 20425 6435 20430 6455
rect 20355 6405 20430 6435
rect 19310 6350 19350 6390
rect 20355 6385 20365 6405
rect 20385 6385 20405 6405
rect 20425 6385 20430 6405
rect 20355 6375 20430 6385
rect 20455 6505 20485 6515
rect 20455 6485 20460 6505
rect 20480 6485 20485 6505
rect 20455 6455 20485 6485
rect 20455 6435 20460 6455
rect 20480 6435 20485 6455
rect 20455 6405 20485 6435
rect 20455 6385 20460 6405
rect 20480 6385 20485 6405
rect 20455 6375 20485 6385
rect 20510 6505 20540 6515
rect 20510 6485 20515 6505
rect 20535 6485 20540 6505
rect 20510 6455 20540 6485
rect 20510 6435 20515 6455
rect 20535 6435 20540 6455
rect 20510 6405 20540 6435
rect 20510 6385 20515 6405
rect 20535 6385 20540 6405
rect 20510 6375 20540 6385
rect 20565 6505 20595 6515
rect 20565 6485 20570 6505
rect 20590 6485 20595 6505
rect 20565 6455 20595 6485
rect 20565 6435 20570 6455
rect 20590 6435 20595 6455
rect 20565 6405 20595 6435
rect 20565 6385 20570 6405
rect 20590 6385 20595 6405
rect 20565 6375 20595 6385
rect 20620 6505 20730 6515
rect 20620 6485 20625 6505
rect 20645 6485 20665 6505
rect 20685 6485 20705 6505
rect 20725 6485 20730 6505
rect 20620 6455 20730 6485
rect 20620 6435 20625 6455
rect 20645 6435 20665 6455
rect 20685 6435 20705 6455
rect 20725 6435 20730 6455
rect 20620 6405 20730 6435
rect 20620 6385 20625 6405
rect 20645 6385 20665 6405
rect 20685 6385 20705 6405
rect 20725 6385 20730 6405
rect 20620 6375 20730 6385
rect 20755 6505 20785 6515
rect 20755 6485 20760 6505
rect 20780 6485 20785 6505
rect 20755 6455 20785 6485
rect 20755 6435 20760 6455
rect 20780 6435 20785 6455
rect 20755 6405 20785 6435
rect 20755 6385 20760 6405
rect 20780 6385 20785 6405
rect 20755 6375 20785 6385
rect 20810 6505 20840 6515
rect 20810 6485 20815 6505
rect 20835 6485 20840 6505
rect 20810 6455 20840 6485
rect 20810 6435 20815 6455
rect 20835 6435 20840 6455
rect 20810 6405 20840 6435
rect 20810 6385 20815 6405
rect 20835 6385 20840 6405
rect 20810 6375 20840 6385
rect 20865 6505 20895 6515
rect 20865 6485 20870 6505
rect 20890 6485 20895 6505
rect 20865 6455 20895 6485
rect 20865 6435 20870 6455
rect 20890 6435 20895 6455
rect 20865 6405 20895 6435
rect 20865 6385 20870 6405
rect 20890 6385 20895 6405
rect 20865 6375 20895 6385
rect 20920 6505 20995 6515
rect 20920 6485 20925 6505
rect 20945 6485 20965 6505
rect 20985 6485 20995 6505
rect 20920 6455 20995 6485
rect 20920 6435 20925 6455
rect 20945 6435 20965 6455
rect 20985 6435 20995 6455
rect 20920 6405 20995 6435
rect 20920 6385 20925 6405
rect 20945 6385 20965 6405
rect 20985 6385 20995 6405
rect 20920 6375 20995 6385
rect 20365 6355 20385 6375
rect 9765 6330 9805 6340
rect 9765 6310 9775 6330
rect 9795 6310 9805 6330
rect 9765 6300 9805 6310
rect 9965 6330 10005 6340
rect 9965 6310 9975 6330
rect 9995 6310 10005 6330
rect 9965 6300 10005 6310
rect 10165 6330 10205 6340
rect 10165 6310 10175 6330
rect 10195 6310 10205 6330
rect 10165 6300 10205 6310
rect 10365 6330 10405 6340
rect 10365 6310 10375 6330
rect 10395 6310 10405 6330
rect 10365 6300 10405 6310
rect 10565 6330 10605 6340
rect 10565 6310 10575 6330
rect 10595 6310 10605 6330
rect 10565 6300 10605 6310
rect 10668 6330 10702 6340
rect 10668 6310 10676 6330
rect 10694 6310 10702 6330
rect 10668 6300 10702 6310
rect 10765 6330 10805 6340
rect 10765 6310 10775 6330
rect 10795 6310 10805 6330
rect 11810 6310 11850 6350
rect 20355 6345 20395 6355
rect 12995 6330 13035 6340
rect 12995 6310 13005 6330
rect 13025 6310 13035 6330
rect 10765 6300 10805 6310
rect 12995 6300 13035 6310
rect 13098 6330 13132 6340
rect 13098 6310 13106 6330
rect 13124 6310 13132 6330
rect 13098 6300 13132 6310
rect 13195 6330 13235 6340
rect 13195 6310 13205 6330
rect 13225 6310 13235 6330
rect 13195 6300 13235 6310
rect 13395 6330 13435 6340
rect 13395 6310 13405 6330
rect 13425 6310 13435 6330
rect 13395 6300 13435 6310
rect 13595 6330 13635 6340
rect 13595 6310 13605 6330
rect 13625 6310 13635 6330
rect 13595 6300 13635 6310
rect 13795 6330 13835 6340
rect 13795 6310 13805 6330
rect 13825 6310 13835 6330
rect 13795 6300 13835 6310
rect 13995 6330 14035 6340
rect 13995 6310 14005 6330
rect 14025 6310 14035 6330
rect 13995 6300 14035 6310
rect 18815 6300 18855 6340
rect 19380 6300 19420 6340
rect 20355 6325 20365 6345
rect 20385 6325 20395 6345
rect 20355 6315 20395 6325
rect 9775 6280 9795 6300
rect 9975 6280 9995 6300
rect 10175 6280 10195 6300
rect 10375 6280 10395 6300
rect 10575 6280 10595 6300
rect 10775 6280 10795 6300
rect 9630 6270 9700 6280
rect 9630 6250 9635 6270
rect 9655 6250 9675 6270
rect 9695 6250 9700 6270
rect 9630 6225 9700 6250
rect 9630 6205 9635 6225
rect 9655 6205 9675 6225
rect 9695 6205 9700 6225
rect 9630 6180 9700 6205
rect 9630 6160 9635 6180
rect 9655 6160 9675 6180
rect 9695 6160 9700 6180
rect 9630 6130 9700 6160
rect 9630 6110 9635 6130
rect 9655 6110 9675 6130
rect 9695 6110 9700 6130
rect 9630 6085 9700 6110
rect 9630 6065 9635 6085
rect 9655 6065 9675 6085
rect 9695 6065 9700 6085
rect 9630 6040 9700 6065
rect 9630 6020 9635 6040
rect 9655 6020 9675 6040
rect 9695 6020 9700 6040
rect 9630 6010 9700 6020
rect 9770 6270 9800 6280
rect 9770 6250 9775 6270
rect 9795 6250 9800 6270
rect 9770 6225 9800 6250
rect 9770 6205 9775 6225
rect 9795 6205 9800 6225
rect 9770 6180 9800 6205
rect 9770 6160 9775 6180
rect 9795 6160 9800 6180
rect 9770 6130 9800 6160
rect 9770 6110 9775 6130
rect 9795 6110 9800 6130
rect 9770 6085 9800 6110
rect 9770 6065 9775 6085
rect 9795 6065 9800 6085
rect 9770 6040 9800 6065
rect 9770 6020 9775 6040
rect 9795 6020 9800 6040
rect 9770 6010 9800 6020
rect 9870 6270 9900 6280
rect 9870 6250 9875 6270
rect 9895 6250 9900 6270
rect 9870 6225 9900 6250
rect 9870 6205 9875 6225
rect 9895 6205 9900 6225
rect 9870 6180 9900 6205
rect 9870 6160 9875 6180
rect 9895 6160 9900 6180
rect 9870 6130 9900 6160
rect 9870 6110 9875 6130
rect 9895 6110 9900 6130
rect 9870 6085 9900 6110
rect 9870 6065 9875 6085
rect 9895 6065 9900 6085
rect 9870 6040 9900 6065
rect 9870 6020 9875 6040
rect 9895 6020 9900 6040
rect 9870 6010 9900 6020
rect 9970 6270 10000 6280
rect 9970 6250 9975 6270
rect 9995 6250 10000 6270
rect 9970 6225 10000 6250
rect 9970 6205 9975 6225
rect 9995 6205 10000 6225
rect 9970 6180 10000 6205
rect 9970 6160 9975 6180
rect 9995 6160 10000 6180
rect 9970 6130 10000 6160
rect 9970 6110 9975 6130
rect 9995 6110 10000 6130
rect 9970 6085 10000 6110
rect 9970 6065 9975 6085
rect 9995 6065 10000 6085
rect 9970 6040 10000 6065
rect 9970 6020 9975 6040
rect 9995 6020 10000 6040
rect 9970 6010 10000 6020
rect 10070 6270 10100 6280
rect 10070 6250 10075 6270
rect 10095 6250 10100 6270
rect 10070 6225 10100 6250
rect 10070 6205 10075 6225
rect 10095 6205 10100 6225
rect 10070 6180 10100 6205
rect 10070 6160 10075 6180
rect 10095 6160 10100 6180
rect 10070 6130 10100 6160
rect 10070 6110 10075 6130
rect 10095 6110 10100 6130
rect 10070 6085 10100 6110
rect 10070 6065 10075 6085
rect 10095 6065 10100 6085
rect 10070 6040 10100 6065
rect 10070 6020 10075 6040
rect 10095 6020 10100 6040
rect 10070 6010 10100 6020
rect 10170 6270 10200 6280
rect 10170 6250 10175 6270
rect 10195 6250 10200 6270
rect 10170 6225 10200 6250
rect 10170 6205 10175 6225
rect 10195 6205 10200 6225
rect 10170 6180 10200 6205
rect 10170 6160 10175 6180
rect 10195 6160 10200 6180
rect 10170 6130 10200 6160
rect 10170 6110 10175 6130
rect 10195 6110 10200 6130
rect 10170 6085 10200 6110
rect 10170 6065 10175 6085
rect 10195 6065 10200 6085
rect 10170 6040 10200 6065
rect 10170 6020 10175 6040
rect 10195 6020 10200 6040
rect 10170 6010 10200 6020
rect 10270 6270 10300 6280
rect 10270 6250 10275 6270
rect 10295 6250 10300 6270
rect 10270 6225 10300 6250
rect 10270 6205 10275 6225
rect 10295 6205 10300 6225
rect 10270 6180 10300 6205
rect 10270 6160 10275 6180
rect 10295 6160 10300 6180
rect 10270 6130 10300 6160
rect 10270 6110 10275 6130
rect 10295 6110 10300 6130
rect 10270 6085 10300 6110
rect 10270 6065 10275 6085
rect 10295 6065 10300 6085
rect 10270 6040 10300 6065
rect 10270 6020 10275 6040
rect 10295 6020 10300 6040
rect 10270 6010 10300 6020
rect 10370 6270 10400 6280
rect 10370 6250 10375 6270
rect 10395 6250 10400 6270
rect 10370 6225 10400 6250
rect 10370 6205 10375 6225
rect 10395 6205 10400 6225
rect 10370 6180 10400 6205
rect 10370 6160 10375 6180
rect 10395 6160 10400 6180
rect 10370 6130 10400 6160
rect 10370 6110 10375 6130
rect 10395 6110 10400 6130
rect 10370 6085 10400 6110
rect 10370 6065 10375 6085
rect 10395 6065 10400 6085
rect 10370 6040 10400 6065
rect 10370 6020 10375 6040
rect 10395 6020 10400 6040
rect 10370 6010 10400 6020
rect 10470 6270 10500 6280
rect 10470 6250 10475 6270
rect 10495 6250 10500 6270
rect 10470 6225 10500 6250
rect 10470 6205 10475 6225
rect 10495 6205 10500 6225
rect 10470 6180 10500 6205
rect 10470 6160 10475 6180
rect 10495 6160 10500 6180
rect 10470 6130 10500 6160
rect 10470 6110 10475 6130
rect 10495 6110 10500 6130
rect 10470 6085 10500 6110
rect 10470 6065 10475 6085
rect 10495 6065 10500 6085
rect 10470 6040 10500 6065
rect 10470 6020 10475 6040
rect 10495 6020 10500 6040
rect 10470 6010 10500 6020
rect 10570 6270 10600 6280
rect 10570 6250 10575 6270
rect 10595 6250 10600 6270
rect 10570 6225 10600 6250
rect 10570 6205 10575 6225
rect 10595 6205 10600 6225
rect 10570 6180 10600 6205
rect 10570 6160 10575 6180
rect 10595 6160 10600 6180
rect 10570 6130 10600 6160
rect 10570 6110 10575 6130
rect 10595 6110 10600 6130
rect 10570 6085 10600 6110
rect 10570 6065 10575 6085
rect 10595 6065 10600 6085
rect 10570 6040 10600 6065
rect 10570 6020 10575 6040
rect 10595 6020 10600 6040
rect 10570 6010 10600 6020
rect 10670 6270 10700 6280
rect 10670 6250 10675 6270
rect 10695 6250 10700 6270
rect 10670 6225 10700 6250
rect 10670 6205 10675 6225
rect 10695 6205 10700 6225
rect 10670 6180 10700 6205
rect 10670 6160 10675 6180
rect 10695 6160 10700 6180
rect 10670 6130 10700 6160
rect 10670 6110 10675 6130
rect 10695 6110 10700 6130
rect 10670 6085 10700 6110
rect 10670 6065 10675 6085
rect 10695 6065 10700 6085
rect 10670 6040 10700 6065
rect 10670 6020 10675 6040
rect 10695 6020 10700 6040
rect 10670 6010 10700 6020
rect 10770 6270 10800 6280
rect 10770 6250 10775 6270
rect 10795 6250 10800 6270
rect 10770 6225 10800 6250
rect 10770 6205 10775 6225
rect 10795 6205 10800 6225
rect 10770 6180 10800 6205
rect 10770 6160 10775 6180
rect 10795 6160 10800 6180
rect 10770 6130 10800 6160
rect 10770 6110 10775 6130
rect 10795 6110 10800 6130
rect 10770 6085 10800 6110
rect 10770 6065 10775 6085
rect 10795 6065 10800 6085
rect 10770 6040 10800 6065
rect 10770 6020 10775 6040
rect 10795 6020 10800 6040
rect 10770 6010 10800 6020
rect 10870 6270 10940 6280
rect 10870 6250 10875 6270
rect 10895 6250 10915 6270
rect 10935 6250 10940 6270
rect 11315 6260 11355 6300
rect 11880 6260 11920 6300
rect 13005 6280 13025 6300
rect 13205 6280 13225 6300
rect 13405 6280 13425 6300
rect 13605 6280 13625 6300
rect 13805 6280 13825 6300
rect 14005 6280 14025 6300
rect 20455 6295 20475 6375
rect 20526 6345 20558 6355
rect 20526 6325 20533 6345
rect 20553 6325 20558 6345
rect 20526 6315 20558 6325
rect 20575 6295 20595 6375
rect 20665 6355 20685 6375
rect 20655 6345 20695 6355
rect 20655 6325 20665 6345
rect 20685 6325 20695 6345
rect 20655 6315 20695 6325
rect 20755 6295 20775 6375
rect 20792 6345 20824 6355
rect 20792 6325 20797 6345
rect 20817 6325 20824 6345
rect 20792 6315 20824 6325
rect 20875 6295 20895 6375
rect 20965 6355 20985 6375
rect 20955 6345 20995 6355
rect 20955 6325 20965 6345
rect 20985 6325 20995 6345
rect 20955 6315 20995 6325
rect 20095 6285 20135 6295
rect 12860 6270 12930 6280
rect 10870 6225 10940 6250
rect 12595 6245 12635 6255
rect 10870 6205 10875 6225
rect 10895 6205 10915 6225
rect 10935 6205 10940 6225
rect 10870 6180 10940 6205
rect 11315 6230 11355 6240
rect 11315 6210 11325 6230
rect 11345 6210 11355 6230
rect 11315 6200 11355 6210
rect 11425 6230 11465 6240
rect 11425 6210 11435 6230
rect 11455 6210 11465 6230
rect 11425 6200 11465 6210
rect 11535 6230 11575 6240
rect 11535 6210 11545 6230
rect 11565 6210 11575 6230
rect 11535 6200 11575 6210
rect 11645 6230 11685 6240
rect 11645 6210 11655 6230
rect 11675 6210 11685 6230
rect 11645 6200 11685 6210
rect 11755 6230 11795 6240
rect 11755 6210 11765 6230
rect 11785 6210 11795 6230
rect 11755 6200 11795 6210
rect 11815 6230 11845 6240
rect 11815 6210 11820 6230
rect 11840 6210 11845 6230
rect 11815 6200 11845 6210
rect 11865 6230 11905 6240
rect 11865 6210 11875 6230
rect 11895 6210 11905 6230
rect 11865 6200 11905 6210
rect 11975 6230 12015 6240
rect 11975 6210 11985 6230
rect 12005 6210 12015 6230
rect 11975 6200 12015 6210
rect 12085 6230 12125 6240
rect 12085 6210 12095 6230
rect 12115 6210 12125 6230
rect 12085 6200 12125 6210
rect 12195 6230 12235 6240
rect 12195 6210 12205 6230
rect 12225 6210 12235 6230
rect 12195 6200 12235 6210
rect 12305 6230 12345 6240
rect 12305 6210 12315 6230
rect 12335 6210 12345 6230
rect 12305 6200 12345 6210
rect 12415 6230 12455 6240
rect 12415 6210 12425 6230
rect 12445 6210 12455 6230
rect 12415 6200 12455 6210
rect 12525 6230 12565 6240
rect 12525 6210 12535 6230
rect 12555 6210 12565 6230
rect 12595 6225 12605 6245
rect 12625 6225 12635 6245
rect 12595 6215 12635 6225
rect 12860 6250 12865 6270
rect 12885 6250 12905 6270
rect 12925 6250 12930 6270
rect 12860 6225 12930 6250
rect 12525 6200 12565 6210
rect 12860 6205 12865 6225
rect 12885 6205 12905 6225
rect 12925 6205 12930 6225
rect 11325 6180 11345 6200
rect 11435 6180 11455 6200
rect 11545 6180 11565 6200
rect 11655 6180 11675 6200
rect 11765 6180 11785 6200
rect 11875 6180 11895 6200
rect 11985 6180 12005 6200
rect 12095 6180 12115 6200
rect 12205 6180 12225 6200
rect 12315 6180 12335 6200
rect 12425 6180 12445 6200
rect 12535 6180 12555 6200
rect 12860 6180 12930 6205
rect 10870 6160 10875 6180
rect 10895 6160 10915 6180
rect 10935 6160 10940 6180
rect 10870 6130 10940 6160
rect 10870 6110 10875 6130
rect 10895 6110 10915 6130
rect 10935 6110 10940 6130
rect 10870 6085 10940 6110
rect 10870 6065 10875 6085
rect 10895 6065 10915 6085
rect 10935 6065 10940 6085
rect 10870 6040 10940 6065
rect 10870 6020 10875 6040
rect 10895 6020 10915 6040
rect 10935 6020 10940 6040
rect 10870 6010 10940 6020
rect 11170 6170 11240 6180
rect 11170 6150 11175 6170
rect 11195 6150 11215 6170
rect 11235 6150 11240 6170
rect 11170 6120 11240 6150
rect 11170 6100 11175 6120
rect 11195 6100 11215 6120
rect 11235 6100 11240 6120
rect 11170 6070 11240 6100
rect 11170 6050 11175 6070
rect 11195 6050 11215 6070
rect 11235 6050 11240 6070
rect 11170 6020 11240 6050
rect 9635 5990 9655 6010
rect 9875 5990 9895 6010
rect 10075 5990 10095 6010
rect 10275 5990 10295 6010
rect 10475 5990 10495 6010
rect 10675 5990 10695 6010
rect 10915 5990 10935 6010
rect 11170 6000 11175 6020
rect 11195 6000 11215 6020
rect 11235 6000 11240 6020
rect 9625 5980 9665 5990
rect 9625 5960 9635 5980
rect 9655 5960 9665 5980
rect 9625 5950 9665 5960
rect 9865 5980 9905 5990
rect 9865 5960 9875 5980
rect 9895 5960 9905 5980
rect 9865 5950 9905 5960
rect 10065 5980 10105 5990
rect 10065 5960 10075 5980
rect 10095 5960 10105 5980
rect 10065 5950 10105 5960
rect 10265 5980 10305 5990
rect 10265 5960 10275 5980
rect 10295 5960 10305 5980
rect 10265 5950 10305 5960
rect 10465 5980 10505 5990
rect 10465 5960 10475 5980
rect 10495 5960 10505 5980
rect 10465 5950 10505 5960
rect 10665 5980 10705 5990
rect 10665 5960 10675 5980
rect 10695 5960 10705 5980
rect 10665 5950 10705 5960
rect 10905 5980 10945 5990
rect 10905 5960 10915 5980
rect 10935 5960 10945 5980
rect 10905 5950 10945 5960
rect 11170 5970 11240 6000
rect 11170 5950 11175 5970
rect 11195 5950 11215 5970
rect 11235 5950 11240 5970
rect 11170 5940 11240 5950
rect 11265 6170 11295 6180
rect 11265 6150 11270 6170
rect 11290 6150 11295 6170
rect 11265 6120 11295 6150
rect 11265 6100 11270 6120
rect 11290 6100 11295 6120
rect 11265 6070 11295 6100
rect 11265 6050 11270 6070
rect 11290 6050 11295 6070
rect 11265 6020 11295 6050
rect 11265 6000 11270 6020
rect 11290 6000 11295 6020
rect 11265 5970 11295 6000
rect 11265 5950 11270 5970
rect 11290 5950 11295 5970
rect 11265 5940 11295 5950
rect 11320 6170 11350 6180
rect 11320 6150 11325 6170
rect 11345 6150 11350 6170
rect 11320 6120 11350 6150
rect 11320 6100 11325 6120
rect 11345 6100 11350 6120
rect 11320 6070 11350 6100
rect 11320 6050 11325 6070
rect 11345 6050 11350 6070
rect 11320 6020 11350 6050
rect 11320 6000 11325 6020
rect 11345 6000 11350 6020
rect 11320 5970 11350 6000
rect 11320 5950 11325 5970
rect 11345 5950 11350 5970
rect 11320 5940 11350 5950
rect 11375 6170 11405 6180
rect 11375 6150 11380 6170
rect 11400 6150 11405 6170
rect 11375 6120 11405 6150
rect 11375 6100 11380 6120
rect 11400 6100 11405 6120
rect 11375 6070 11405 6100
rect 11375 6050 11380 6070
rect 11400 6050 11405 6070
rect 11375 6020 11405 6050
rect 11375 6000 11380 6020
rect 11400 6000 11405 6020
rect 11375 5970 11405 6000
rect 11375 5950 11380 5970
rect 11400 5950 11405 5970
rect 11375 5940 11405 5950
rect 11430 6170 11460 6180
rect 11430 6150 11435 6170
rect 11455 6150 11460 6170
rect 11430 6120 11460 6150
rect 11430 6100 11435 6120
rect 11455 6100 11460 6120
rect 11430 6070 11460 6100
rect 11430 6050 11435 6070
rect 11455 6050 11460 6070
rect 11430 6020 11460 6050
rect 11430 6000 11435 6020
rect 11455 6000 11460 6020
rect 11430 5970 11460 6000
rect 11430 5950 11435 5970
rect 11455 5950 11460 5970
rect 11430 5940 11460 5950
rect 11485 6170 11515 6180
rect 11485 6150 11490 6170
rect 11510 6150 11515 6170
rect 11485 6120 11515 6150
rect 11485 6100 11490 6120
rect 11510 6100 11515 6120
rect 11485 6070 11515 6100
rect 11485 6050 11490 6070
rect 11510 6050 11515 6070
rect 11485 6020 11515 6050
rect 11485 6000 11490 6020
rect 11510 6000 11515 6020
rect 11485 5970 11515 6000
rect 11485 5950 11490 5970
rect 11510 5950 11515 5970
rect 11485 5940 11515 5950
rect 11540 6170 11570 6180
rect 11540 6150 11545 6170
rect 11565 6150 11570 6170
rect 11540 6120 11570 6150
rect 11540 6100 11545 6120
rect 11565 6100 11570 6120
rect 11540 6070 11570 6100
rect 11540 6050 11545 6070
rect 11565 6050 11570 6070
rect 11540 6020 11570 6050
rect 11540 6000 11545 6020
rect 11565 6000 11570 6020
rect 11540 5970 11570 6000
rect 11540 5950 11545 5970
rect 11565 5950 11570 5970
rect 11540 5940 11570 5950
rect 11595 6170 11625 6180
rect 11595 6150 11600 6170
rect 11620 6150 11625 6170
rect 11595 6120 11625 6150
rect 11595 6100 11600 6120
rect 11620 6100 11625 6120
rect 11595 6070 11625 6100
rect 11595 6050 11600 6070
rect 11620 6050 11625 6070
rect 11595 6020 11625 6050
rect 11595 6000 11600 6020
rect 11620 6000 11625 6020
rect 11595 5970 11625 6000
rect 11595 5950 11600 5970
rect 11620 5950 11625 5970
rect 11595 5940 11625 5950
rect 11650 6170 11680 6180
rect 11650 6150 11655 6170
rect 11675 6150 11680 6170
rect 11650 6120 11680 6150
rect 11650 6100 11655 6120
rect 11675 6100 11680 6120
rect 11650 6070 11680 6100
rect 11650 6050 11655 6070
rect 11675 6050 11680 6070
rect 11650 6020 11680 6050
rect 11650 6000 11655 6020
rect 11675 6000 11680 6020
rect 11650 5970 11680 6000
rect 11650 5950 11655 5970
rect 11675 5950 11680 5970
rect 11650 5940 11680 5950
rect 11705 6170 11735 6180
rect 11705 6150 11710 6170
rect 11730 6150 11735 6170
rect 11705 6120 11735 6150
rect 11705 6100 11710 6120
rect 11730 6100 11735 6120
rect 11705 6070 11735 6100
rect 11705 6050 11710 6070
rect 11730 6050 11735 6070
rect 11705 6020 11735 6050
rect 11705 6000 11710 6020
rect 11730 6000 11735 6020
rect 11705 5970 11735 6000
rect 11705 5950 11710 5970
rect 11730 5950 11735 5970
rect 11705 5940 11735 5950
rect 11760 6170 11790 6180
rect 11760 6150 11765 6170
rect 11785 6150 11790 6170
rect 11760 6120 11790 6150
rect 11760 6100 11765 6120
rect 11785 6100 11790 6120
rect 11760 6070 11790 6100
rect 11760 6050 11765 6070
rect 11785 6050 11790 6070
rect 11760 6020 11790 6050
rect 11760 6000 11765 6020
rect 11785 6000 11790 6020
rect 11760 5970 11790 6000
rect 11760 5950 11765 5970
rect 11785 5950 11790 5970
rect 11760 5940 11790 5950
rect 11815 6170 11845 6180
rect 11815 6150 11820 6170
rect 11840 6150 11845 6170
rect 11815 6120 11845 6150
rect 11815 6100 11820 6120
rect 11840 6100 11845 6120
rect 11815 6070 11845 6100
rect 11815 6050 11820 6070
rect 11840 6050 11845 6070
rect 11815 6020 11845 6050
rect 11815 6000 11820 6020
rect 11840 6000 11845 6020
rect 11815 5970 11845 6000
rect 11815 5950 11820 5970
rect 11840 5950 11845 5970
rect 11815 5940 11845 5950
rect 11870 6170 11900 6180
rect 11870 6150 11875 6170
rect 11895 6150 11900 6170
rect 11870 6120 11900 6150
rect 11870 6100 11875 6120
rect 11895 6100 11900 6120
rect 11870 6070 11900 6100
rect 11870 6050 11875 6070
rect 11895 6050 11900 6070
rect 11870 6020 11900 6050
rect 11870 6000 11875 6020
rect 11895 6000 11900 6020
rect 11870 5970 11900 6000
rect 11870 5950 11875 5970
rect 11895 5950 11900 5970
rect 11870 5940 11900 5950
rect 11925 6170 11955 6180
rect 11925 6150 11930 6170
rect 11950 6150 11955 6170
rect 11925 6120 11955 6150
rect 11925 6100 11930 6120
rect 11950 6100 11955 6120
rect 11925 6070 11955 6100
rect 11925 6050 11930 6070
rect 11950 6050 11955 6070
rect 11925 6020 11955 6050
rect 11925 6000 11930 6020
rect 11950 6000 11955 6020
rect 11925 5970 11955 6000
rect 11925 5950 11930 5970
rect 11950 5950 11955 5970
rect 11925 5940 11955 5950
rect 11980 6170 12010 6180
rect 11980 6150 11985 6170
rect 12005 6150 12010 6170
rect 11980 6120 12010 6150
rect 11980 6100 11985 6120
rect 12005 6100 12010 6120
rect 11980 6070 12010 6100
rect 11980 6050 11985 6070
rect 12005 6050 12010 6070
rect 11980 6020 12010 6050
rect 11980 6000 11985 6020
rect 12005 6000 12010 6020
rect 11980 5970 12010 6000
rect 11980 5950 11985 5970
rect 12005 5950 12010 5970
rect 11980 5940 12010 5950
rect 12035 6170 12065 6180
rect 12035 6150 12040 6170
rect 12060 6150 12065 6170
rect 12035 6120 12065 6150
rect 12035 6100 12040 6120
rect 12060 6100 12065 6120
rect 12035 6070 12065 6100
rect 12035 6050 12040 6070
rect 12060 6050 12065 6070
rect 12035 6020 12065 6050
rect 12035 6000 12040 6020
rect 12060 6000 12065 6020
rect 12035 5970 12065 6000
rect 12035 5950 12040 5970
rect 12060 5950 12065 5970
rect 12035 5940 12065 5950
rect 12090 6170 12120 6180
rect 12090 6150 12095 6170
rect 12115 6150 12120 6170
rect 12090 6120 12120 6150
rect 12090 6100 12095 6120
rect 12115 6100 12120 6120
rect 12090 6070 12120 6100
rect 12090 6050 12095 6070
rect 12115 6050 12120 6070
rect 12090 6020 12120 6050
rect 12090 6000 12095 6020
rect 12115 6000 12120 6020
rect 12090 5970 12120 6000
rect 12090 5950 12095 5970
rect 12115 5950 12120 5970
rect 12090 5940 12120 5950
rect 12145 6170 12175 6180
rect 12145 6150 12150 6170
rect 12170 6150 12175 6170
rect 12145 6120 12175 6150
rect 12145 6100 12150 6120
rect 12170 6100 12175 6120
rect 12145 6070 12175 6100
rect 12145 6050 12150 6070
rect 12170 6050 12175 6070
rect 12145 6020 12175 6050
rect 12145 6000 12150 6020
rect 12170 6000 12175 6020
rect 12145 5970 12175 6000
rect 12145 5950 12150 5970
rect 12170 5950 12175 5970
rect 12145 5940 12175 5950
rect 12200 6170 12230 6180
rect 12200 6150 12205 6170
rect 12225 6150 12230 6170
rect 12200 6120 12230 6150
rect 12200 6100 12205 6120
rect 12225 6100 12230 6120
rect 12200 6070 12230 6100
rect 12200 6050 12205 6070
rect 12225 6050 12230 6070
rect 12200 6020 12230 6050
rect 12200 6000 12205 6020
rect 12225 6000 12230 6020
rect 12200 5970 12230 6000
rect 12200 5950 12205 5970
rect 12225 5950 12230 5970
rect 12200 5940 12230 5950
rect 12255 6170 12285 6180
rect 12255 6150 12260 6170
rect 12280 6150 12285 6170
rect 12255 6120 12285 6150
rect 12255 6100 12260 6120
rect 12280 6100 12285 6120
rect 12255 6070 12285 6100
rect 12255 6050 12260 6070
rect 12280 6050 12285 6070
rect 12255 6020 12285 6050
rect 12255 6000 12260 6020
rect 12280 6000 12285 6020
rect 12255 5970 12285 6000
rect 12255 5950 12260 5970
rect 12280 5950 12285 5970
rect 12255 5940 12285 5950
rect 12310 6170 12340 6180
rect 12310 6150 12315 6170
rect 12335 6150 12340 6170
rect 12310 6120 12340 6150
rect 12310 6100 12315 6120
rect 12335 6100 12340 6120
rect 12310 6070 12340 6100
rect 12310 6050 12315 6070
rect 12335 6050 12340 6070
rect 12310 6020 12340 6050
rect 12310 6000 12315 6020
rect 12335 6000 12340 6020
rect 12310 5970 12340 6000
rect 12310 5950 12315 5970
rect 12335 5950 12340 5970
rect 12310 5940 12340 5950
rect 12365 6170 12395 6180
rect 12365 6150 12370 6170
rect 12390 6150 12395 6170
rect 12365 6120 12395 6150
rect 12365 6100 12370 6120
rect 12390 6100 12395 6120
rect 12365 6070 12395 6100
rect 12365 6050 12370 6070
rect 12390 6050 12395 6070
rect 12365 6020 12395 6050
rect 12365 6000 12370 6020
rect 12390 6000 12395 6020
rect 12365 5970 12395 6000
rect 12365 5950 12370 5970
rect 12390 5950 12395 5970
rect 12365 5940 12395 5950
rect 12420 6170 12450 6180
rect 12420 6150 12425 6170
rect 12445 6150 12450 6170
rect 12420 6120 12450 6150
rect 12420 6100 12425 6120
rect 12445 6100 12450 6120
rect 12420 6070 12450 6100
rect 12420 6050 12425 6070
rect 12445 6050 12450 6070
rect 12420 6020 12450 6050
rect 12420 6000 12425 6020
rect 12445 6000 12450 6020
rect 12420 5970 12450 6000
rect 12420 5950 12425 5970
rect 12445 5950 12450 5970
rect 12420 5940 12450 5950
rect 12475 6170 12505 6180
rect 12475 6150 12480 6170
rect 12500 6150 12505 6170
rect 12475 6120 12505 6150
rect 12475 6100 12480 6120
rect 12500 6100 12505 6120
rect 12475 6070 12505 6100
rect 12475 6050 12480 6070
rect 12500 6050 12505 6070
rect 12475 6020 12505 6050
rect 12475 6000 12480 6020
rect 12500 6000 12505 6020
rect 12475 5970 12505 6000
rect 12475 5950 12480 5970
rect 12500 5950 12505 5970
rect 12475 5940 12505 5950
rect 12530 6170 12560 6180
rect 12530 6150 12535 6170
rect 12555 6150 12560 6170
rect 12530 6120 12560 6150
rect 12530 6100 12535 6120
rect 12555 6100 12560 6120
rect 12530 6070 12560 6100
rect 12530 6050 12535 6070
rect 12555 6050 12560 6070
rect 12530 6020 12560 6050
rect 12530 6000 12535 6020
rect 12555 6000 12560 6020
rect 12530 5970 12560 6000
rect 12530 5950 12535 5970
rect 12555 5950 12560 5970
rect 12530 5940 12560 5950
rect 12585 6170 12655 6180
rect 12585 6150 12590 6170
rect 12610 6150 12630 6170
rect 12650 6150 12655 6170
rect 12585 6120 12655 6150
rect 12585 6100 12590 6120
rect 12610 6100 12630 6120
rect 12650 6100 12655 6120
rect 12585 6070 12655 6100
rect 12585 6050 12590 6070
rect 12610 6050 12630 6070
rect 12650 6050 12655 6070
rect 12585 6020 12655 6050
rect 12585 6000 12590 6020
rect 12610 6000 12630 6020
rect 12650 6000 12655 6020
rect 12860 6160 12865 6180
rect 12885 6160 12905 6180
rect 12925 6160 12930 6180
rect 12860 6130 12930 6160
rect 12860 6110 12865 6130
rect 12885 6110 12905 6130
rect 12925 6110 12930 6130
rect 12860 6085 12930 6110
rect 12860 6065 12865 6085
rect 12885 6065 12905 6085
rect 12925 6065 12930 6085
rect 12860 6040 12930 6065
rect 12860 6020 12865 6040
rect 12885 6020 12905 6040
rect 12925 6020 12930 6040
rect 12860 6010 12930 6020
rect 13000 6270 13030 6280
rect 13000 6250 13005 6270
rect 13025 6250 13030 6270
rect 13000 6225 13030 6250
rect 13000 6205 13005 6225
rect 13025 6205 13030 6225
rect 13000 6180 13030 6205
rect 13000 6160 13005 6180
rect 13025 6160 13030 6180
rect 13000 6130 13030 6160
rect 13000 6110 13005 6130
rect 13025 6110 13030 6130
rect 13000 6085 13030 6110
rect 13000 6065 13005 6085
rect 13025 6065 13030 6085
rect 13000 6040 13030 6065
rect 13000 6020 13005 6040
rect 13025 6020 13030 6040
rect 13000 6010 13030 6020
rect 13100 6270 13130 6280
rect 13100 6250 13105 6270
rect 13125 6250 13130 6270
rect 13100 6225 13130 6250
rect 13100 6205 13105 6225
rect 13125 6205 13130 6225
rect 13100 6180 13130 6205
rect 13100 6160 13105 6180
rect 13125 6160 13130 6180
rect 13100 6130 13130 6160
rect 13100 6110 13105 6130
rect 13125 6110 13130 6130
rect 13100 6085 13130 6110
rect 13100 6065 13105 6085
rect 13125 6065 13130 6085
rect 13100 6040 13130 6065
rect 13100 6020 13105 6040
rect 13125 6020 13130 6040
rect 13100 6010 13130 6020
rect 13200 6270 13230 6280
rect 13200 6250 13205 6270
rect 13225 6250 13230 6270
rect 13200 6225 13230 6250
rect 13200 6205 13205 6225
rect 13225 6205 13230 6225
rect 13200 6180 13230 6205
rect 13200 6160 13205 6180
rect 13225 6160 13230 6180
rect 13200 6130 13230 6160
rect 13200 6110 13205 6130
rect 13225 6110 13230 6130
rect 13200 6085 13230 6110
rect 13200 6065 13205 6085
rect 13225 6065 13230 6085
rect 13200 6040 13230 6065
rect 13200 6020 13205 6040
rect 13225 6020 13230 6040
rect 13200 6010 13230 6020
rect 13300 6270 13330 6280
rect 13300 6250 13305 6270
rect 13325 6250 13330 6270
rect 13300 6225 13330 6250
rect 13300 6205 13305 6225
rect 13325 6205 13330 6225
rect 13300 6180 13330 6205
rect 13300 6160 13305 6180
rect 13325 6160 13330 6180
rect 13300 6130 13330 6160
rect 13300 6110 13305 6130
rect 13325 6110 13330 6130
rect 13300 6085 13330 6110
rect 13300 6065 13305 6085
rect 13325 6065 13330 6085
rect 13300 6040 13330 6065
rect 13300 6020 13305 6040
rect 13325 6020 13330 6040
rect 13300 6010 13330 6020
rect 13400 6270 13430 6280
rect 13400 6250 13405 6270
rect 13425 6250 13430 6270
rect 13400 6225 13430 6250
rect 13400 6205 13405 6225
rect 13425 6205 13430 6225
rect 13400 6180 13430 6205
rect 13400 6160 13405 6180
rect 13425 6160 13430 6180
rect 13400 6130 13430 6160
rect 13400 6110 13405 6130
rect 13425 6110 13430 6130
rect 13400 6085 13430 6110
rect 13400 6065 13405 6085
rect 13425 6065 13430 6085
rect 13400 6040 13430 6065
rect 13400 6020 13405 6040
rect 13425 6020 13430 6040
rect 13400 6010 13430 6020
rect 13500 6270 13530 6280
rect 13500 6250 13505 6270
rect 13525 6250 13530 6270
rect 13500 6225 13530 6250
rect 13500 6205 13505 6225
rect 13525 6205 13530 6225
rect 13500 6180 13530 6205
rect 13500 6160 13505 6180
rect 13525 6160 13530 6180
rect 13500 6130 13530 6160
rect 13500 6110 13505 6130
rect 13525 6110 13530 6130
rect 13500 6085 13530 6110
rect 13500 6065 13505 6085
rect 13525 6065 13530 6085
rect 13500 6040 13530 6065
rect 13500 6020 13505 6040
rect 13525 6020 13530 6040
rect 13500 6010 13530 6020
rect 13600 6270 13630 6280
rect 13600 6250 13605 6270
rect 13625 6250 13630 6270
rect 13600 6225 13630 6250
rect 13600 6205 13605 6225
rect 13625 6205 13630 6225
rect 13600 6180 13630 6205
rect 13600 6160 13605 6180
rect 13625 6160 13630 6180
rect 13600 6130 13630 6160
rect 13600 6110 13605 6130
rect 13625 6110 13630 6130
rect 13600 6085 13630 6110
rect 13600 6065 13605 6085
rect 13625 6065 13630 6085
rect 13600 6040 13630 6065
rect 13600 6020 13605 6040
rect 13625 6020 13630 6040
rect 13600 6010 13630 6020
rect 13700 6270 13730 6280
rect 13700 6250 13705 6270
rect 13725 6250 13730 6270
rect 13700 6225 13730 6250
rect 13700 6205 13705 6225
rect 13725 6205 13730 6225
rect 13700 6180 13730 6205
rect 13700 6160 13705 6180
rect 13725 6160 13730 6180
rect 13700 6130 13730 6160
rect 13700 6110 13705 6130
rect 13725 6110 13730 6130
rect 13700 6085 13730 6110
rect 13700 6065 13705 6085
rect 13725 6065 13730 6085
rect 13700 6040 13730 6065
rect 13700 6020 13705 6040
rect 13725 6020 13730 6040
rect 13700 6010 13730 6020
rect 13800 6270 13830 6280
rect 13800 6250 13805 6270
rect 13825 6250 13830 6270
rect 13800 6225 13830 6250
rect 13800 6205 13805 6225
rect 13825 6205 13830 6225
rect 13800 6180 13830 6205
rect 13800 6160 13805 6180
rect 13825 6160 13830 6180
rect 13800 6130 13830 6160
rect 13800 6110 13805 6130
rect 13825 6110 13830 6130
rect 13800 6085 13830 6110
rect 13800 6065 13805 6085
rect 13825 6065 13830 6085
rect 13800 6040 13830 6065
rect 13800 6020 13805 6040
rect 13825 6020 13830 6040
rect 13800 6010 13830 6020
rect 13900 6270 13930 6280
rect 13900 6250 13905 6270
rect 13925 6250 13930 6270
rect 13900 6225 13930 6250
rect 13900 6205 13905 6225
rect 13925 6205 13930 6225
rect 13900 6180 13930 6205
rect 13900 6160 13905 6180
rect 13925 6160 13930 6180
rect 13900 6130 13930 6160
rect 13900 6110 13905 6130
rect 13925 6110 13930 6130
rect 13900 6085 13930 6110
rect 13900 6065 13905 6085
rect 13925 6065 13930 6085
rect 13900 6040 13930 6065
rect 13900 6020 13905 6040
rect 13925 6020 13930 6040
rect 13900 6010 13930 6020
rect 14000 6270 14030 6280
rect 14000 6250 14005 6270
rect 14025 6250 14030 6270
rect 14000 6225 14030 6250
rect 14000 6205 14005 6225
rect 14025 6205 14030 6225
rect 14000 6180 14030 6205
rect 14000 6160 14005 6180
rect 14025 6160 14030 6180
rect 14000 6130 14030 6160
rect 14000 6110 14005 6130
rect 14025 6110 14030 6130
rect 14000 6085 14030 6110
rect 14000 6065 14005 6085
rect 14025 6065 14030 6085
rect 14000 6040 14030 6065
rect 14000 6020 14005 6040
rect 14025 6020 14030 6040
rect 14000 6010 14030 6020
rect 14100 6270 14170 6280
rect 14100 6250 14105 6270
rect 14125 6250 14145 6270
rect 14165 6250 14170 6270
rect 14100 6225 14170 6250
rect 18815 6270 18855 6280
rect 18815 6250 18825 6270
rect 18845 6250 18855 6270
rect 18815 6240 18855 6250
rect 18925 6270 18965 6280
rect 18925 6250 18935 6270
rect 18955 6250 18965 6270
rect 18925 6240 18965 6250
rect 19035 6270 19075 6280
rect 19035 6250 19045 6270
rect 19065 6250 19075 6270
rect 19035 6240 19075 6250
rect 19145 6270 19185 6280
rect 19145 6250 19155 6270
rect 19175 6250 19185 6270
rect 19145 6240 19185 6250
rect 19255 6270 19295 6280
rect 19255 6250 19265 6270
rect 19285 6250 19295 6270
rect 19255 6240 19295 6250
rect 19315 6270 19345 6280
rect 19315 6250 19320 6270
rect 19340 6250 19345 6270
rect 19315 6240 19345 6250
rect 19365 6270 19405 6280
rect 19365 6250 19375 6270
rect 19395 6250 19405 6270
rect 19365 6240 19405 6250
rect 19475 6270 19515 6280
rect 19475 6250 19485 6270
rect 19505 6250 19515 6270
rect 19475 6240 19515 6250
rect 19585 6270 19625 6280
rect 19585 6250 19595 6270
rect 19615 6250 19625 6270
rect 19585 6240 19625 6250
rect 19695 6270 19735 6280
rect 19695 6250 19705 6270
rect 19725 6250 19735 6270
rect 19695 6240 19735 6250
rect 19805 6270 19845 6280
rect 19805 6250 19815 6270
rect 19835 6250 19845 6270
rect 19805 6240 19845 6250
rect 19915 6270 19955 6280
rect 19915 6250 19925 6270
rect 19945 6250 19955 6270
rect 19915 6240 19955 6250
rect 20025 6270 20065 6280
rect 20025 6250 20035 6270
rect 20055 6250 20065 6270
rect 20095 6265 20105 6285
rect 20125 6265 20135 6285
rect 20095 6255 20135 6265
rect 20445 6285 20485 6295
rect 20445 6265 20455 6285
rect 20475 6265 20485 6285
rect 20445 6255 20485 6265
rect 20560 6285 20600 6295
rect 20560 6265 20570 6285
rect 20590 6265 20600 6285
rect 20560 6255 20600 6265
rect 20750 6285 20790 6295
rect 20750 6265 20760 6285
rect 20780 6265 20790 6285
rect 20750 6255 20790 6265
rect 20865 6285 20905 6295
rect 20865 6265 20875 6285
rect 20895 6265 20905 6285
rect 20865 6255 20905 6265
rect 20025 6240 20065 6250
rect 14100 6205 14105 6225
rect 14125 6205 14145 6225
rect 14165 6205 14170 6225
rect 18825 6220 18845 6240
rect 18935 6220 18955 6240
rect 19045 6220 19065 6240
rect 19155 6220 19175 6240
rect 19265 6220 19285 6240
rect 19375 6220 19395 6240
rect 19485 6220 19505 6240
rect 19595 6220 19615 6240
rect 19705 6220 19725 6240
rect 19815 6220 19835 6240
rect 19925 6220 19945 6240
rect 20035 6220 20055 6240
rect 20600 6225 20640 6235
rect 14100 6180 14170 6205
rect 14100 6160 14105 6180
rect 14125 6160 14145 6180
rect 14165 6160 14170 6180
rect 14100 6130 14170 6160
rect 14100 6110 14105 6130
rect 14125 6110 14145 6130
rect 14165 6110 14170 6130
rect 14100 6085 14170 6110
rect 14100 6065 14105 6085
rect 14125 6065 14145 6085
rect 14165 6065 14170 6085
rect 14100 6040 14170 6065
rect 14100 6020 14105 6040
rect 14125 6020 14145 6040
rect 14165 6020 14170 6040
rect 14100 6010 14170 6020
rect 18670 6210 18740 6220
rect 18670 6190 18675 6210
rect 18695 6190 18715 6210
rect 18735 6190 18740 6210
rect 18670 6160 18740 6190
rect 18670 6140 18675 6160
rect 18695 6140 18715 6160
rect 18735 6140 18740 6160
rect 18670 6110 18740 6140
rect 18670 6090 18675 6110
rect 18695 6090 18715 6110
rect 18735 6090 18740 6110
rect 18670 6060 18740 6090
rect 18670 6040 18675 6060
rect 18695 6040 18715 6060
rect 18735 6040 18740 6060
rect 18670 6010 18740 6040
rect 12585 5970 12655 6000
rect 12865 5990 12885 6010
rect 13105 5990 13125 6010
rect 13305 5990 13325 6010
rect 13505 5990 13525 6010
rect 13705 5990 13725 6010
rect 13905 5990 13925 6010
rect 14145 5990 14165 6010
rect 18670 5990 18675 6010
rect 18695 5990 18715 6010
rect 18735 5990 18740 6010
rect 12585 5950 12590 5970
rect 12610 5950 12630 5970
rect 12650 5950 12655 5970
rect 12855 5980 12895 5990
rect 12855 5960 12865 5980
rect 12885 5960 12895 5980
rect 12855 5950 12895 5960
rect 13095 5980 13135 5990
rect 13095 5960 13105 5980
rect 13125 5960 13135 5980
rect 13095 5950 13135 5960
rect 13295 5980 13335 5990
rect 13295 5960 13305 5980
rect 13325 5960 13335 5980
rect 13295 5950 13335 5960
rect 13495 5980 13535 5990
rect 13495 5960 13505 5980
rect 13525 5960 13535 5980
rect 13495 5950 13535 5960
rect 13695 5980 13735 5990
rect 13695 5960 13705 5980
rect 13725 5960 13735 5980
rect 13695 5950 13735 5960
rect 13895 5980 13935 5990
rect 13895 5960 13905 5980
rect 13925 5960 13935 5980
rect 13895 5950 13935 5960
rect 14135 5980 14175 5990
rect 18670 5980 18740 5990
rect 18765 6210 18795 6220
rect 18765 6190 18770 6210
rect 18790 6190 18795 6210
rect 18765 6160 18795 6190
rect 18765 6140 18770 6160
rect 18790 6140 18795 6160
rect 18765 6110 18795 6140
rect 18765 6090 18770 6110
rect 18790 6090 18795 6110
rect 18765 6060 18795 6090
rect 18765 6040 18770 6060
rect 18790 6040 18795 6060
rect 18765 6010 18795 6040
rect 18765 5990 18770 6010
rect 18790 5990 18795 6010
rect 18765 5980 18795 5990
rect 18820 6210 18850 6220
rect 18820 6190 18825 6210
rect 18845 6190 18850 6210
rect 18820 6160 18850 6190
rect 18820 6140 18825 6160
rect 18845 6140 18850 6160
rect 18820 6110 18850 6140
rect 18820 6090 18825 6110
rect 18845 6090 18850 6110
rect 18820 6060 18850 6090
rect 18820 6040 18825 6060
rect 18845 6040 18850 6060
rect 18820 6010 18850 6040
rect 18820 5990 18825 6010
rect 18845 5990 18850 6010
rect 18820 5980 18850 5990
rect 18875 6210 18905 6220
rect 18875 6190 18880 6210
rect 18900 6190 18905 6210
rect 18875 6160 18905 6190
rect 18875 6140 18880 6160
rect 18900 6140 18905 6160
rect 18875 6110 18905 6140
rect 18875 6090 18880 6110
rect 18900 6090 18905 6110
rect 18875 6060 18905 6090
rect 18875 6040 18880 6060
rect 18900 6040 18905 6060
rect 18875 6010 18905 6040
rect 18875 5990 18880 6010
rect 18900 5990 18905 6010
rect 18875 5980 18905 5990
rect 18930 6210 18960 6220
rect 18930 6190 18935 6210
rect 18955 6190 18960 6210
rect 18930 6160 18960 6190
rect 18930 6140 18935 6160
rect 18955 6140 18960 6160
rect 18930 6110 18960 6140
rect 18930 6090 18935 6110
rect 18955 6090 18960 6110
rect 18930 6060 18960 6090
rect 18930 6040 18935 6060
rect 18955 6040 18960 6060
rect 18930 6010 18960 6040
rect 18930 5990 18935 6010
rect 18955 5990 18960 6010
rect 18930 5980 18960 5990
rect 18985 6210 19015 6220
rect 18985 6190 18990 6210
rect 19010 6190 19015 6210
rect 18985 6160 19015 6190
rect 18985 6140 18990 6160
rect 19010 6140 19015 6160
rect 18985 6110 19015 6140
rect 18985 6090 18990 6110
rect 19010 6090 19015 6110
rect 18985 6060 19015 6090
rect 18985 6040 18990 6060
rect 19010 6040 19015 6060
rect 18985 6010 19015 6040
rect 18985 5990 18990 6010
rect 19010 5990 19015 6010
rect 18985 5980 19015 5990
rect 19040 6210 19070 6220
rect 19040 6190 19045 6210
rect 19065 6190 19070 6210
rect 19040 6160 19070 6190
rect 19040 6140 19045 6160
rect 19065 6140 19070 6160
rect 19040 6110 19070 6140
rect 19040 6090 19045 6110
rect 19065 6090 19070 6110
rect 19040 6060 19070 6090
rect 19040 6040 19045 6060
rect 19065 6040 19070 6060
rect 19040 6010 19070 6040
rect 19040 5990 19045 6010
rect 19065 5990 19070 6010
rect 19040 5980 19070 5990
rect 19095 6210 19125 6220
rect 19095 6190 19100 6210
rect 19120 6190 19125 6210
rect 19095 6160 19125 6190
rect 19095 6140 19100 6160
rect 19120 6140 19125 6160
rect 19095 6110 19125 6140
rect 19095 6090 19100 6110
rect 19120 6090 19125 6110
rect 19095 6060 19125 6090
rect 19095 6040 19100 6060
rect 19120 6040 19125 6060
rect 19095 6010 19125 6040
rect 19095 5990 19100 6010
rect 19120 5990 19125 6010
rect 19095 5980 19125 5990
rect 19150 6210 19180 6220
rect 19150 6190 19155 6210
rect 19175 6190 19180 6210
rect 19150 6160 19180 6190
rect 19150 6140 19155 6160
rect 19175 6140 19180 6160
rect 19150 6110 19180 6140
rect 19150 6090 19155 6110
rect 19175 6090 19180 6110
rect 19150 6060 19180 6090
rect 19150 6040 19155 6060
rect 19175 6040 19180 6060
rect 19150 6010 19180 6040
rect 19150 5990 19155 6010
rect 19175 5990 19180 6010
rect 19150 5980 19180 5990
rect 19205 6210 19235 6220
rect 19205 6190 19210 6210
rect 19230 6190 19235 6210
rect 19205 6160 19235 6190
rect 19205 6140 19210 6160
rect 19230 6140 19235 6160
rect 19205 6110 19235 6140
rect 19205 6090 19210 6110
rect 19230 6090 19235 6110
rect 19205 6060 19235 6090
rect 19205 6040 19210 6060
rect 19230 6040 19235 6060
rect 19205 6010 19235 6040
rect 19205 5990 19210 6010
rect 19230 5990 19235 6010
rect 19205 5980 19235 5990
rect 19260 6210 19290 6220
rect 19260 6190 19265 6210
rect 19285 6190 19290 6210
rect 19260 6160 19290 6190
rect 19260 6140 19265 6160
rect 19285 6140 19290 6160
rect 19260 6110 19290 6140
rect 19260 6090 19265 6110
rect 19285 6090 19290 6110
rect 19260 6060 19290 6090
rect 19260 6040 19265 6060
rect 19285 6040 19290 6060
rect 19260 6010 19290 6040
rect 19260 5990 19265 6010
rect 19285 5990 19290 6010
rect 19260 5980 19290 5990
rect 19315 6210 19345 6220
rect 19315 6190 19320 6210
rect 19340 6190 19345 6210
rect 19315 6160 19345 6190
rect 19315 6140 19320 6160
rect 19340 6140 19345 6160
rect 19315 6110 19345 6140
rect 19315 6090 19320 6110
rect 19340 6090 19345 6110
rect 19315 6060 19345 6090
rect 19315 6040 19320 6060
rect 19340 6040 19345 6060
rect 19315 6010 19345 6040
rect 19315 5990 19320 6010
rect 19340 5990 19345 6010
rect 19315 5980 19345 5990
rect 19370 6210 19400 6220
rect 19370 6190 19375 6210
rect 19395 6190 19400 6210
rect 19370 6160 19400 6190
rect 19370 6140 19375 6160
rect 19395 6140 19400 6160
rect 19370 6110 19400 6140
rect 19370 6090 19375 6110
rect 19395 6090 19400 6110
rect 19370 6060 19400 6090
rect 19370 6040 19375 6060
rect 19395 6040 19400 6060
rect 19370 6010 19400 6040
rect 19370 5990 19375 6010
rect 19395 5990 19400 6010
rect 19370 5980 19400 5990
rect 19425 6210 19455 6220
rect 19425 6190 19430 6210
rect 19450 6190 19455 6210
rect 19425 6160 19455 6190
rect 19425 6140 19430 6160
rect 19450 6140 19455 6160
rect 19425 6110 19455 6140
rect 19425 6090 19430 6110
rect 19450 6090 19455 6110
rect 19425 6060 19455 6090
rect 19425 6040 19430 6060
rect 19450 6040 19455 6060
rect 19425 6010 19455 6040
rect 19425 5990 19430 6010
rect 19450 5990 19455 6010
rect 19425 5980 19455 5990
rect 19480 6210 19510 6220
rect 19480 6190 19485 6210
rect 19505 6190 19510 6210
rect 19480 6160 19510 6190
rect 19480 6140 19485 6160
rect 19505 6140 19510 6160
rect 19480 6110 19510 6140
rect 19480 6090 19485 6110
rect 19505 6090 19510 6110
rect 19480 6060 19510 6090
rect 19480 6040 19485 6060
rect 19505 6040 19510 6060
rect 19480 6010 19510 6040
rect 19480 5990 19485 6010
rect 19505 5990 19510 6010
rect 19480 5980 19510 5990
rect 19535 6210 19565 6220
rect 19535 6190 19540 6210
rect 19560 6190 19565 6210
rect 19535 6160 19565 6190
rect 19535 6140 19540 6160
rect 19560 6140 19565 6160
rect 19535 6110 19565 6140
rect 19535 6090 19540 6110
rect 19560 6090 19565 6110
rect 19535 6060 19565 6090
rect 19535 6040 19540 6060
rect 19560 6040 19565 6060
rect 19535 6010 19565 6040
rect 19535 5990 19540 6010
rect 19560 5990 19565 6010
rect 19535 5980 19565 5990
rect 19590 6210 19620 6220
rect 19590 6190 19595 6210
rect 19615 6190 19620 6210
rect 19590 6160 19620 6190
rect 19590 6140 19595 6160
rect 19615 6140 19620 6160
rect 19590 6110 19620 6140
rect 19590 6090 19595 6110
rect 19615 6090 19620 6110
rect 19590 6060 19620 6090
rect 19590 6040 19595 6060
rect 19615 6040 19620 6060
rect 19590 6010 19620 6040
rect 19590 5990 19595 6010
rect 19615 5990 19620 6010
rect 19590 5980 19620 5990
rect 19645 6210 19675 6220
rect 19645 6190 19650 6210
rect 19670 6190 19675 6210
rect 19645 6160 19675 6190
rect 19645 6140 19650 6160
rect 19670 6140 19675 6160
rect 19645 6110 19675 6140
rect 19645 6090 19650 6110
rect 19670 6090 19675 6110
rect 19645 6060 19675 6090
rect 19645 6040 19650 6060
rect 19670 6040 19675 6060
rect 19645 6010 19675 6040
rect 19645 5990 19650 6010
rect 19670 5990 19675 6010
rect 19645 5980 19675 5990
rect 19700 6210 19730 6220
rect 19700 6190 19705 6210
rect 19725 6190 19730 6210
rect 19700 6160 19730 6190
rect 19700 6140 19705 6160
rect 19725 6140 19730 6160
rect 19700 6110 19730 6140
rect 19700 6090 19705 6110
rect 19725 6090 19730 6110
rect 19700 6060 19730 6090
rect 19700 6040 19705 6060
rect 19725 6040 19730 6060
rect 19700 6010 19730 6040
rect 19700 5990 19705 6010
rect 19725 5990 19730 6010
rect 19700 5980 19730 5990
rect 19755 6210 19785 6220
rect 19755 6190 19760 6210
rect 19780 6190 19785 6210
rect 19755 6160 19785 6190
rect 19755 6140 19760 6160
rect 19780 6140 19785 6160
rect 19755 6110 19785 6140
rect 19755 6090 19760 6110
rect 19780 6090 19785 6110
rect 19755 6060 19785 6090
rect 19755 6040 19760 6060
rect 19780 6040 19785 6060
rect 19755 6010 19785 6040
rect 19755 5990 19760 6010
rect 19780 5990 19785 6010
rect 19755 5980 19785 5990
rect 19810 6210 19840 6220
rect 19810 6190 19815 6210
rect 19835 6190 19840 6210
rect 19810 6160 19840 6190
rect 19810 6140 19815 6160
rect 19835 6140 19840 6160
rect 19810 6110 19840 6140
rect 19810 6090 19815 6110
rect 19835 6090 19840 6110
rect 19810 6060 19840 6090
rect 19810 6040 19815 6060
rect 19835 6040 19840 6060
rect 19810 6010 19840 6040
rect 19810 5990 19815 6010
rect 19835 5990 19840 6010
rect 19810 5980 19840 5990
rect 19865 6210 19895 6220
rect 19865 6190 19870 6210
rect 19890 6190 19895 6210
rect 19865 6160 19895 6190
rect 19865 6140 19870 6160
rect 19890 6140 19895 6160
rect 19865 6110 19895 6140
rect 19865 6090 19870 6110
rect 19890 6090 19895 6110
rect 19865 6060 19895 6090
rect 19865 6040 19870 6060
rect 19890 6040 19895 6060
rect 19865 6010 19895 6040
rect 19865 5990 19870 6010
rect 19890 5990 19895 6010
rect 19865 5980 19895 5990
rect 19920 6210 19950 6220
rect 19920 6190 19925 6210
rect 19945 6190 19950 6210
rect 19920 6160 19950 6190
rect 19920 6140 19925 6160
rect 19945 6140 19950 6160
rect 19920 6110 19950 6140
rect 19920 6090 19925 6110
rect 19945 6090 19950 6110
rect 19920 6060 19950 6090
rect 19920 6040 19925 6060
rect 19945 6040 19950 6060
rect 19920 6010 19950 6040
rect 19920 5990 19925 6010
rect 19945 5990 19950 6010
rect 19920 5980 19950 5990
rect 19975 6210 20005 6220
rect 19975 6190 19980 6210
rect 20000 6190 20005 6210
rect 19975 6160 20005 6190
rect 19975 6140 19980 6160
rect 20000 6140 20005 6160
rect 19975 6110 20005 6140
rect 19975 6090 19980 6110
rect 20000 6090 20005 6110
rect 19975 6060 20005 6090
rect 19975 6040 19980 6060
rect 20000 6040 20005 6060
rect 19975 6010 20005 6040
rect 19975 5990 19980 6010
rect 20000 5990 20005 6010
rect 19975 5980 20005 5990
rect 20030 6210 20060 6220
rect 20030 6190 20035 6210
rect 20055 6190 20060 6210
rect 20030 6160 20060 6190
rect 20030 6140 20035 6160
rect 20055 6140 20060 6160
rect 20030 6110 20060 6140
rect 20030 6090 20035 6110
rect 20055 6090 20060 6110
rect 20030 6060 20060 6090
rect 20030 6040 20035 6060
rect 20055 6040 20060 6060
rect 20030 6010 20060 6040
rect 20030 5990 20035 6010
rect 20055 5990 20060 6010
rect 20030 5980 20060 5990
rect 20085 6210 20155 6220
rect 20085 6190 20090 6210
rect 20110 6190 20130 6210
rect 20150 6190 20155 6210
rect 20600 6205 20610 6225
rect 20630 6205 20640 6225
rect 20600 6195 20640 6205
rect 20660 6225 20690 6235
rect 20660 6205 20665 6225
rect 20685 6205 20690 6225
rect 20660 6195 20690 6205
rect 20710 6225 20750 6235
rect 20710 6205 20720 6225
rect 20740 6205 20750 6225
rect 20710 6195 20750 6205
rect 20085 6160 20155 6190
rect 20610 6175 20630 6195
rect 20720 6175 20740 6195
rect 20085 6140 20090 6160
rect 20110 6140 20130 6160
rect 20150 6140 20155 6160
rect 20085 6110 20155 6140
rect 20085 6090 20090 6110
rect 20110 6090 20130 6110
rect 20150 6090 20155 6110
rect 20085 6060 20155 6090
rect 20085 6040 20090 6060
rect 20110 6040 20130 6060
rect 20150 6040 20155 6060
rect 20085 6010 20155 6040
rect 20510 6165 20580 6175
rect 20510 6145 20515 6165
rect 20535 6145 20555 6165
rect 20575 6145 20580 6165
rect 20510 6115 20580 6145
rect 20510 6095 20515 6115
rect 20535 6095 20555 6115
rect 20575 6095 20580 6115
rect 20510 6065 20580 6095
rect 20510 6045 20515 6065
rect 20535 6045 20555 6065
rect 20575 6045 20580 6065
rect 20510 6035 20580 6045
rect 20605 6165 20635 6175
rect 20605 6145 20610 6165
rect 20630 6145 20635 6165
rect 20605 6115 20635 6145
rect 20605 6095 20610 6115
rect 20630 6095 20635 6115
rect 20605 6065 20635 6095
rect 20605 6045 20610 6065
rect 20630 6045 20635 6065
rect 20605 6035 20635 6045
rect 20660 6165 20690 6175
rect 20660 6145 20665 6165
rect 20685 6145 20690 6165
rect 20660 6115 20690 6145
rect 20660 6095 20665 6115
rect 20685 6095 20690 6115
rect 20660 6065 20690 6095
rect 20660 6045 20665 6065
rect 20685 6045 20690 6065
rect 20660 6035 20690 6045
rect 20715 6165 20745 6175
rect 20715 6145 20720 6165
rect 20740 6145 20745 6165
rect 20715 6115 20745 6145
rect 20715 6095 20720 6115
rect 20740 6095 20745 6115
rect 20715 6065 20745 6095
rect 20715 6045 20720 6065
rect 20740 6045 20745 6065
rect 20715 6035 20745 6045
rect 20770 6165 20840 6175
rect 20770 6145 20775 6165
rect 20795 6145 20815 6165
rect 20835 6145 20840 6165
rect 20770 6115 20840 6145
rect 20770 6095 20775 6115
rect 20795 6095 20815 6115
rect 20835 6095 20840 6115
rect 20770 6065 20840 6095
rect 20770 6045 20775 6065
rect 20795 6045 20815 6065
rect 20835 6045 20840 6065
rect 20770 6035 20840 6045
rect 20515 6015 20535 6035
rect 20720 6015 20740 6035
rect 20815 6015 20835 6035
rect 20085 5990 20090 6010
rect 20110 5990 20130 6010
rect 20150 5990 20155 6010
rect 20085 5980 20155 5990
rect 20505 6005 20545 6015
rect 20505 5985 20515 6005
rect 20535 5985 20545 6005
rect 14135 5960 14145 5980
rect 14165 5960 14175 5980
rect 18675 5960 18695 5980
rect 18770 5960 18790 5980
rect 18880 5960 18900 5980
rect 18990 5960 19010 5980
rect 19100 5960 19120 5980
rect 19210 5960 19230 5980
rect 19320 5960 19340 5980
rect 19430 5960 19450 5980
rect 19540 5960 19560 5980
rect 19650 5960 19670 5980
rect 19760 5960 19780 5980
rect 19870 5960 19890 5980
rect 19980 5960 20000 5980
rect 20130 5960 20150 5980
rect 20505 5975 20545 5985
rect 20685 6005 20740 6015
rect 20685 5985 20695 6005
rect 20715 5995 20740 6005
rect 20805 6005 20845 6015
rect 20715 5985 20725 5995
rect 20685 5975 20725 5985
rect 20805 5985 20815 6005
rect 20835 5985 20845 6005
rect 20805 5975 20845 5985
rect 14135 5950 14175 5960
rect 18665 5950 18705 5960
rect 12585 5940 12655 5950
rect 11175 5920 11195 5940
rect 11270 5920 11290 5940
rect 11380 5920 11400 5940
rect 11490 5920 11510 5940
rect 11600 5920 11620 5940
rect 11710 5920 11730 5940
rect 11820 5920 11840 5940
rect 11930 5920 11950 5940
rect 12040 5920 12060 5940
rect 12150 5920 12170 5940
rect 12260 5920 12280 5940
rect 12370 5920 12390 5940
rect 12480 5920 12500 5940
rect 12630 5920 12650 5940
rect 18665 5930 18675 5950
rect 18695 5930 18705 5950
rect 18665 5920 18705 5930
rect 18760 5950 18800 5960
rect 18760 5930 18770 5950
rect 18790 5930 18800 5950
rect 18760 5920 18800 5930
rect 18870 5950 18910 5960
rect 18870 5930 18880 5950
rect 18900 5930 18910 5950
rect 18870 5920 18910 5930
rect 18980 5950 19020 5960
rect 18980 5930 18990 5950
rect 19010 5930 19020 5950
rect 18980 5920 19020 5930
rect 19090 5950 19130 5960
rect 19090 5930 19100 5950
rect 19120 5930 19130 5950
rect 19090 5920 19130 5930
rect 19200 5950 19240 5960
rect 19200 5930 19210 5950
rect 19230 5930 19240 5950
rect 19200 5920 19240 5930
rect 19310 5950 19350 5960
rect 19310 5930 19320 5950
rect 19340 5930 19350 5950
rect 19310 5920 19350 5930
rect 19420 5950 19460 5960
rect 19420 5930 19430 5950
rect 19450 5930 19460 5950
rect 19420 5920 19460 5930
rect 19530 5950 19570 5960
rect 19530 5930 19540 5950
rect 19560 5930 19570 5950
rect 19530 5920 19570 5930
rect 19640 5950 19680 5960
rect 19640 5930 19650 5950
rect 19670 5930 19680 5950
rect 19640 5920 19680 5930
rect 19750 5950 19790 5960
rect 19750 5930 19760 5950
rect 19780 5930 19790 5950
rect 19750 5920 19790 5930
rect 19860 5950 19900 5960
rect 19860 5930 19870 5950
rect 19890 5930 19900 5950
rect 19860 5920 19900 5930
rect 19970 5950 20010 5960
rect 19970 5930 19980 5950
rect 20000 5930 20010 5950
rect 19970 5920 20010 5930
rect 20120 5950 20160 5960
rect 20120 5930 20130 5950
rect 20150 5930 20160 5950
rect 20120 5920 20160 5930
rect 11165 5910 11205 5920
rect 11165 5890 11175 5910
rect 11195 5890 11205 5910
rect 11165 5880 11205 5890
rect 11260 5910 11300 5920
rect 11260 5890 11270 5910
rect 11290 5890 11300 5910
rect 11260 5880 11300 5890
rect 11370 5910 11410 5920
rect 11370 5890 11380 5910
rect 11400 5890 11410 5910
rect 11370 5880 11410 5890
rect 11480 5910 11520 5920
rect 11480 5890 11490 5910
rect 11510 5890 11520 5910
rect 11480 5880 11520 5890
rect 11590 5910 11630 5920
rect 11590 5890 11600 5910
rect 11620 5890 11630 5910
rect 11590 5880 11630 5890
rect 11700 5910 11740 5920
rect 11700 5890 11710 5910
rect 11730 5890 11740 5910
rect 11700 5880 11740 5890
rect 11810 5910 11850 5920
rect 11810 5890 11820 5910
rect 11840 5890 11850 5910
rect 11810 5880 11850 5890
rect 11920 5910 11960 5920
rect 11920 5890 11930 5910
rect 11950 5890 11960 5910
rect 11920 5880 11960 5890
rect 12030 5910 12070 5920
rect 12030 5890 12040 5910
rect 12060 5890 12070 5910
rect 12030 5880 12070 5890
rect 12140 5910 12180 5920
rect 12140 5890 12150 5910
rect 12170 5890 12180 5910
rect 12140 5880 12180 5890
rect 12250 5910 12290 5920
rect 12250 5890 12260 5910
rect 12280 5890 12290 5910
rect 12250 5880 12290 5890
rect 12360 5910 12400 5920
rect 12360 5890 12370 5910
rect 12390 5890 12400 5910
rect 12360 5880 12400 5890
rect 12470 5910 12510 5920
rect 12470 5890 12480 5910
rect 12500 5890 12510 5910
rect 12470 5880 12510 5890
rect 12620 5910 12660 5920
rect 12620 5890 12630 5910
rect 12650 5890 12660 5910
rect 12620 5880 12660 5890
rect 11632 4510 11668 4520
rect 11632 4490 11640 4510
rect 11660 4490 11668 4510
rect 11632 4480 11668 4490
rect 11752 4510 11788 4520
rect 11752 4490 11760 4510
rect 11780 4490 11788 4510
rect 11752 4480 11788 4490
rect 11872 4510 11908 4520
rect 11872 4490 11880 4510
rect 11900 4490 11908 4510
rect 11872 4480 11908 4490
rect 11570 4465 11610 4475
rect 11200 4450 11240 4460
rect 11200 4430 11210 4450
rect 11230 4430 11240 4450
rect 11200 4420 11240 4430
rect 11460 4450 11500 4460
rect 11460 4430 11470 4450
rect 11490 4430 11500 4450
rect 11570 4445 11580 4465
rect 11600 4445 11610 4465
rect 11570 4435 11610 4445
rect 11460 4420 11500 4430
rect 11210 4398 11230 4420
rect 11470 4398 11490 4420
rect 11580 4415 11600 4435
rect 11640 4415 11660 4480
rect 11690 4465 11730 4475
rect 11690 4445 11700 4465
rect 11720 4445 11730 4465
rect 11690 4435 11730 4445
rect 11700 4415 11720 4435
rect 11760 4415 11780 4480
rect 11810 4465 11850 4475
rect 11810 4445 11820 4465
rect 11840 4445 11850 4465
rect 11810 4435 11850 4445
rect 11820 4415 11840 4435
rect 11880 4415 11900 4480
rect 11930 4465 11970 4475
rect 11930 4445 11940 4465
rect 11960 4445 11970 4465
rect 11930 4435 11970 4445
rect 12080 4440 12120 4450
rect 11940 4415 11960 4435
rect 12080 4420 12090 4440
rect 12110 4420 12120 4440
rect 11205 4375 11275 4398
rect 11205 4355 11210 4375
rect 11230 4355 11250 4375
rect 11270 4355 11275 4375
rect 11205 4345 11275 4355
rect 11305 4380 11335 4398
rect 11305 4360 11310 4380
rect 11330 4360 11335 4380
rect 11305 4345 11335 4360
rect 11365 4380 11395 4398
rect 11365 4360 11370 4380
rect 11390 4360 11395 4380
rect 11365 4345 11395 4360
rect 11425 4375 11495 4398
rect 11425 4355 11430 4375
rect 11450 4355 11470 4375
rect 11490 4355 11495 4375
rect 11425 4345 11495 4355
rect 11535 4390 11605 4415
rect 11535 4370 11540 4390
rect 11560 4370 11580 4390
rect 11600 4370 11605 4390
rect 11535 4345 11605 4370
rect 11635 4390 11665 4415
rect 11635 4370 11640 4390
rect 11660 4370 11665 4390
rect 11635 4345 11665 4370
rect 11695 4390 11725 4415
rect 11695 4370 11700 4390
rect 11720 4370 11725 4390
rect 11695 4345 11725 4370
rect 11755 4390 11785 4415
rect 11755 4370 11760 4390
rect 11780 4370 11785 4390
rect 11755 4345 11785 4370
rect 11815 4390 11845 4415
rect 11815 4370 11820 4390
rect 11840 4370 11845 4390
rect 11815 4345 11845 4370
rect 11875 4390 11905 4415
rect 11875 4370 11880 4390
rect 11900 4370 11905 4390
rect 11875 4345 11905 4370
rect 11935 4390 12005 4415
rect 12080 4410 12120 4420
rect 12200 4440 12240 4450
rect 12200 4420 12210 4440
rect 12230 4420 12240 4440
rect 12200 4410 12240 4420
rect 12320 4440 12360 4450
rect 12320 4420 12330 4440
rect 12350 4420 12360 4440
rect 12320 4410 12360 4420
rect 12440 4440 12480 4450
rect 12440 4420 12450 4440
rect 12470 4420 12480 4440
rect 12440 4410 12480 4420
rect 12560 4440 12600 4450
rect 12560 4420 12570 4440
rect 12590 4420 12600 4440
rect 12560 4410 12600 4420
rect 12090 4390 12110 4410
rect 12210 4390 12230 4410
rect 12330 4390 12350 4410
rect 12450 4390 12470 4410
rect 12570 4390 12590 4410
rect 11935 4370 11940 4390
rect 11960 4370 11980 4390
rect 12000 4370 12005 4390
rect 11935 4345 12005 4370
rect 12045 4375 12115 4390
rect 12045 4355 12050 4375
rect 12070 4355 12090 4375
rect 12110 4355 12115 4375
rect 11370 4325 11390 4345
rect 12045 4340 12115 4355
rect 12145 4375 12175 4390
rect 12145 4355 12150 4375
rect 12170 4355 12175 4375
rect 12145 4340 12175 4355
rect 12205 4375 12235 4390
rect 12205 4355 12210 4375
rect 12230 4355 12235 4375
rect 12205 4340 12235 4355
rect 12265 4375 12295 4390
rect 12265 4355 12270 4375
rect 12290 4355 12295 4375
rect 12265 4340 12295 4355
rect 12325 4375 12355 4390
rect 12325 4355 12330 4375
rect 12350 4355 12355 4375
rect 12325 4340 12355 4355
rect 12385 4375 12415 4390
rect 12385 4355 12390 4375
rect 12410 4355 12415 4375
rect 12385 4340 12415 4355
rect 12445 4375 12475 4390
rect 12445 4355 12450 4375
rect 12470 4355 12475 4375
rect 12445 4340 12475 4355
rect 12505 4375 12535 4390
rect 12505 4355 12510 4375
rect 12530 4355 12535 4375
rect 12505 4340 12535 4355
rect 12565 4375 12635 4390
rect 12565 4355 12570 4375
rect 12590 4355 12610 4375
rect 12630 4355 12635 4375
rect 12565 4340 12635 4355
rect 11330 4320 11390 4325
rect 12150 4320 12170 4340
rect 12270 4320 12290 4340
rect 12390 4320 12410 4340
rect 12510 4320 12530 4340
rect 11330 4295 11340 4320
rect 11360 4305 11390 4320
rect 11750 4310 11790 4320
rect 11360 4295 11370 4305
rect 11330 4285 11370 4295
rect 11750 4290 11760 4310
rect 11780 4290 11790 4310
rect 11750 4280 11790 4290
rect 12140 4310 12180 4320
rect 12140 4290 12150 4310
rect 12170 4290 12180 4310
rect 12140 4280 12180 4290
rect 12203 4310 12237 4320
rect 12203 4290 12211 4310
rect 12229 4290 12237 4310
rect 12203 4280 12237 4290
rect 12260 4310 12300 4320
rect 12260 4290 12270 4310
rect 12290 4290 12300 4310
rect 12260 4280 12300 4290
rect 12380 4310 12420 4320
rect 12380 4290 12390 4310
rect 12410 4290 12420 4310
rect 12380 4280 12420 4290
rect 12500 4310 12540 4320
rect 12500 4290 12510 4310
rect 12530 4290 12540 4310
rect 12500 4280 12540 4290
rect 11210 4200 11250 4210
rect 11210 4180 11220 4200
rect 11240 4180 11250 4200
rect 11210 4170 11250 4180
rect 11360 4200 11400 4210
rect 11360 4180 11370 4200
rect 11390 4180 11400 4200
rect 11360 4170 11400 4180
rect 11470 4200 11510 4210
rect 11470 4180 11480 4200
rect 11500 4180 11510 4200
rect 11470 4170 11510 4180
rect 11580 4200 11620 4210
rect 11580 4180 11590 4200
rect 11610 4180 11620 4200
rect 11580 4170 11620 4180
rect 11690 4200 11730 4210
rect 11690 4180 11700 4200
rect 11720 4180 11730 4200
rect 11690 4170 11730 4180
rect 11800 4200 11840 4210
rect 11800 4180 11810 4200
rect 11830 4180 11840 4200
rect 11800 4170 11840 4180
rect 11910 4200 11950 4210
rect 11910 4180 11920 4200
rect 11940 4180 11950 4200
rect 11910 4170 11950 4180
rect 12020 4200 12060 4210
rect 12020 4180 12030 4200
rect 12050 4180 12060 4200
rect 12020 4170 12060 4180
rect 12130 4200 12170 4210
rect 12130 4180 12140 4200
rect 12160 4180 12170 4200
rect 12130 4170 12170 4180
rect 12240 4200 12280 4210
rect 12240 4180 12250 4200
rect 12270 4180 12280 4200
rect 12240 4170 12280 4180
rect 12350 4200 12390 4210
rect 12350 4180 12360 4200
rect 12380 4180 12390 4200
rect 12350 4170 12390 4180
rect 12500 4200 12540 4210
rect 12500 4180 12510 4200
rect 12530 4180 12540 4200
rect 12500 4170 12540 4180
rect 11220 4150 11240 4170
rect 11370 4150 11390 4170
rect 11480 4150 11500 4170
rect 11590 4150 11610 4170
rect 11700 4150 11720 4170
rect 11810 4150 11830 4170
rect 11920 4150 11940 4170
rect 12030 4150 12050 4170
rect 12140 4150 12160 4170
rect 12250 4150 12270 4170
rect 12360 4150 12380 4170
rect 12510 4150 12530 4170
rect 11215 4140 11285 4150
rect 11215 4120 11220 4140
rect 11240 4120 11260 4140
rect 11280 4120 11285 4140
rect 11215 4110 11285 4120
rect 11310 4140 11340 4150
rect 11310 4120 11315 4140
rect 11335 4120 11340 4140
rect 11310 4110 11340 4120
rect 11365 4140 11395 4150
rect 11365 4120 11370 4140
rect 11390 4120 11395 4140
rect 11365 4110 11395 4120
rect 11420 4140 11450 4150
rect 11420 4120 11425 4140
rect 11445 4120 11450 4140
rect 11420 4110 11450 4120
rect 11475 4140 11505 4150
rect 11475 4120 11480 4140
rect 11500 4120 11505 4140
rect 11475 4110 11505 4120
rect 11530 4140 11560 4150
rect 11530 4120 11535 4140
rect 11555 4120 11560 4140
rect 11530 4110 11560 4120
rect 11585 4140 11615 4150
rect 11585 4120 11590 4140
rect 11610 4120 11615 4140
rect 11585 4110 11615 4120
rect 11640 4140 11670 4150
rect 11640 4120 11645 4140
rect 11665 4120 11670 4140
rect 11640 4110 11670 4120
rect 11695 4140 11725 4150
rect 11695 4120 11700 4140
rect 11720 4120 11725 4140
rect 11695 4110 11725 4120
rect 11750 4140 11780 4150
rect 11750 4120 11755 4140
rect 11775 4120 11780 4140
rect 11750 4110 11780 4120
rect 11805 4140 11835 4150
rect 11805 4120 11810 4140
rect 11830 4120 11835 4140
rect 11805 4110 11835 4120
rect 11860 4140 11890 4150
rect 11860 4120 11865 4140
rect 11885 4120 11890 4140
rect 11860 4110 11890 4120
rect 11915 4140 11945 4150
rect 11915 4120 11920 4140
rect 11940 4120 11945 4140
rect 11915 4110 11945 4120
rect 11970 4140 12000 4150
rect 11970 4120 11975 4140
rect 11995 4120 12000 4140
rect 11970 4110 12000 4120
rect 12025 4140 12055 4150
rect 12025 4120 12030 4140
rect 12050 4120 12055 4140
rect 12025 4110 12055 4120
rect 12080 4140 12110 4150
rect 12080 4120 12085 4140
rect 12105 4120 12110 4140
rect 12080 4110 12110 4120
rect 12135 4140 12165 4150
rect 12135 4120 12140 4140
rect 12160 4120 12165 4140
rect 12135 4110 12165 4120
rect 12190 4140 12220 4150
rect 12190 4120 12195 4140
rect 12215 4120 12220 4140
rect 12190 4110 12220 4120
rect 12245 4140 12275 4150
rect 12245 4120 12250 4140
rect 12270 4120 12275 4140
rect 12245 4110 12275 4120
rect 12300 4140 12330 4150
rect 12300 4120 12305 4140
rect 12325 4120 12330 4140
rect 12300 4110 12330 4120
rect 12355 4140 12385 4150
rect 12355 4120 12360 4140
rect 12380 4120 12385 4140
rect 12355 4110 12385 4120
rect 12410 4140 12440 4150
rect 12410 4120 12415 4140
rect 12435 4120 12440 4140
rect 12410 4110 12440 4120
rect 12465 4140 12535 4150
rect 12465 4120 12470 4140
rect 12490 4120 12510 4140
rect 12530 4120 12535 4140
rect 12465 4110 12535 4120
rect 11315 4090 11335 4110
rect 11425 4090 11445 4110
rect 11535 4090 11555 4110
rect 11645 4090 11665 4110
rect 11755 4090 11775 4110
rect 11865 4090 11885 4110
rect 11975 4090 11995 4110
rect 12085 4090 12105 4110
rect 12195 4090 12215 4110
rect 12305 4090 12325 4110
rect 12415 4090 12435 4110
rect 11305 4080 11345 4090
rect 11305 4060 11315 4080
rect 11335 4060 11345 4080
rect 11305 4050 11345 4060
rect 11362 4080 11398 4090
rect 11362 4060 11370 4080
rect 11390 4060 11398 4080
rect 11362 4050 11398 4060
rect 11415 4080 11455 4090
rect 11415 4060 11425 4080
rect 11445 4060 11455 4080
rect 11415 4050 11455 4060
rect 11525 4080 11565 4090
rect 11525 4060 11535 4080
rect 11555 4060 11565 4080
rect 11525 4050 11565 4060
rect 11635 4080 11675 4090
rect 11635 4060 11645 4080
rect 11665 4060 11675 4080
rect 11635 4050 11675 4060
rect 11745 4080 11785 4090
rect 11745 4060 11755 4080
rect 11775 4060 11785 4080
rect 11745 4050 11785 4060
rect 11855 4080 11895 4090
rect 11855 4060 11865 4080
rect 11885 4060 11895 4080
rect 11855 4050 11895 4060
rect 11965 4080 12005 4090
rect 11965 4060 11975 4080
rect 11995 4060 12005 4080
rect 11965 4050 12005 4060
rect 12075 4080 12115 4090
rect 12075 4060 12085 4080
rect 12105 4060 12115 4080
rect 12075 4050 12115 4060
rect 12185 4080 12225 4090
rect 12185 4060 12195 4080
rect 12215 4060 12225 4080
rect 12185 4050 12225 4060
rect 12295 4080 12335 4090
rect 12295 4060 12305 4080
rect 12325 4060 12335 4080
rect 12295 4050 12335 4060
rect 12405 4080 12445 4090
rect 12405 4060 12415 4080
rect 12435 4060 12445 4080
rect 12405 4050 12445 4060
rect 11415 3990 11455 4030
rect 11635 3990 11675 4030
rect 11855 3990 11895 4030
rect 12075 3990 12115 4030
rect 12295 3990 12335 4030
rect 11310 3955 11350 3965
rect 11310 3935 11320 3955
rect 11340 3935 11350 3955
rect 11310 3925 11350 3935
rect 11415 3955 11455 3965
rect 11415 3935 11425 3955
rect 11445 3935 11455 3955
rect 11415 3925 11455 3935
rect 11525 3955 11565 3965
rect 11525 3935 11535 3955
rect 11555 3935 11565 3955
rect 11525 3925 11565 3935
rect 11635 3955 11675 3965
rect 11635 3935 11645 3955
rect 11665 3935 11675 3955
rect 11635 3925 11675 3935
rect 11745 3955 11785 3965
rect 11745 3935 11755 3955
rect 11775 3935 11785 3955
rect 11745 3925 11785 3935
rect 12050 3955 12090 3965
rect 12050 3935 12060 3955
rect 12080 3935 12090 3955
rect 12050 3925 12090 3935
rect 12155 3955 12195 3965
rect 12155 3935 12165 3955
rect 12185 3935 12195 3955
rect 12155 3925 12195 3935
rect 12265 3955 12305 3965
rect 12265 3935 12275 3955
rect 12295 3935 12305 3955
rect 12265 3925 12305 3935
rect 12375 3955 12415 3965
rect 12375 3935 12385 3955
rect 12405 3935 12415 3955
rect 12375 3925 12415 3935
rect 12485 3955 12525 3965
rect 12485 3935 12495 3955
rect 12515 3935 12525 3955
rect 12485 3925 12525 3935
rect 11155 3895 11195 3905
rect 11155 3875 11165 3895
rect 11185 3875 11195 3895
rect 11155 3865 11195 3875
rect 11271 3895 11303 3905
rect 11271 3875 11277 3895
rect 11294 3875 11303 3895
rect 11271 3865 11303 3875
rect 11165 3845 11185 3865
rect 11320 3845 11340 3925
rect 11360 3895 11400 3905
rect 11360 3875 11370 3895
rect 11390 3875 11400 3895
rect 11360 3865 11400 3875
rect 11370 3845 11390 3865
rect 11425 3845 11445 3925
rect 11470 3895 11510 3905
rect 11470 3875 11480 3895
rect 11500 3875 11510 3895
rect 11470 3865 11510 3875
rect 11535 3845 11555 3925
rect 11645 3845 11665 3925
rect 11690 3895 11730 3905
rect 11690 3875 11700 3895
rect 11720 3875 11730 3895
rect 11690 3865 11730 3875
rect 11755 3845 11775 3925
rect 11800 3895 11840 3905
rect 11800 3875 11810 3895
rect 11830 3875 11840 3895
rect 11800 3865 11840 3875
rect 11895 3895 11935 3905
rect 11895 3875 11905 3895
rect 11925 3875 11935 3895
rect 11895 3865 11935 3875
rect 12011 3895 12043 3905
rect 12011 3875 12017 3895
rect 12034 3875 12043 3895
rect 12011 3865 12043 3875
rect 11810 3845 11830 3865
rect 11905 3845 11925 3865
rect 12060 3845 12080 3925
rect 12165 3845 12185 3925
rect 12210 3895 12250 3905
rect 12210 3875 12220 3895
rect 12240 3875 12250 3895
rect 12210 3865 12250 3875
rect 12275 3845 12295 3925
rect 12385 3845 12405 3925
rect 12430 3895 12470 3905
rect 12430 3875 12440 3895
rect 12460 3875 12470 3895
rect 12430 3865 12470 3875
rect 12495 3845 12515 3925
rect 12635 3895 12675 3905
rect 12635 3875 12645 3895
rect 12665 3875 12675 3895
rect 12635 3865 12675 3875
rect 12765 3870 12795 3900
rect 12645 3845 12665 3865
rect 11155 3835 11230 3845
rect 11155 3815 11165 3835
rect 11185 3815 11205 3835
rect 11225 3815 11230 3835
rect 11155 3805 11230 3815
rect 11255 3835 11285 3845
rect 11255 3815 11260 3835
rect 11280 3815 11285 3835
rect 11255 3805 11285 3815
rect 11310 3835 11340 3845
rect 11310 3815 11315 3835
rect 11335 3815 11340 3835
rect 11310 3805 11340 3815
rect 11365 3835 11395 3845
rect 11365 3815 11370 3835
rect 11390 3815 11395 3835
rect 11365 3805 11395 3815
rect 11420 3835 11450 3845
rect 11420 3815 11425 3835
rect 11445 3815 11450 3835
rect 11420 3805 11450 3815
rect 11475 3835 11505 3845
rect 11475 3815 11480 3835
rect 11500 3815 11505 3835
rect 11475 3805 11505 3815
rect 11530 3835 11560 3845
rect 11530 3815 11535 3835
rect 11555 3815 11560 3835
rect 11530 3805 11560 3815
rect 11585 3835 11615 3845
rect 11585 3815 11590 3835
rect 11610 3815 11615 3835
rect 11585 3805 11615 3815
rect 11640 3835 11670 3845
rect 11640 3815 11645 3835
rect 11665 3815 11670 3835
rect 11640 3805 11670 3815
rect 11695 3835 11725 3845
rect 11695 3815 11700 3835
rect 11720 3815 11725 3835
rect 11695 3805 11725 3815
rect 11750 3835 11780 3845
rect 11750 3815 11755 3835
rect 11775 3815 11780 3835
rect 11750 3805 11780 3815
rect 11805 3835 11835 3845
rect 11805 3815 11810 3835
rect 11830 3815 11835 3835
rect 11805 3805 11835 3815
rect 11860 3835 11970 3845
rect 11860 3815 11865 3835
rect 11885 3815 11905 3835
rect 11925 3815 11945 3835
rect 11965 3815 11970 3835
rect 11860 3805 11970 3815
rect 11995 3835 12025 3845
rect 11995 3815 12000 3835
rect 12020 3815 12025 3835
rect 11995 3805 12025 3815
rect 12050 3835 12080 3845
rect 12050 3815 12055 3835
rect 12075 3815 12080 3835
rect 12050 3805 12080 3815
rect 12105 3835 12135 3845
rect 12105 3815 12110 3835
rect 12130 3815 12135 3835
rect 12105 3805 12135 3815
rect 12160 3835 12190 3845
rect 12160 3815 12165 3835
rect 12185 3815 12190 3835
rect 12160 3805 12190 3815
rect 12215 3835 12245 3845
rect 12215 3815 12220 3835
rect 12240 3815 12245 3835
rect 12215 3805 12245 3815
rect 12270 3835 12300 3845
rect 12270 3815 12275 3835
rect 12295 3815 12300 3835
rect 12270 3805 12300 3815
rect 12325 3835 12355 3845
rect 12325 3815 12330 3835
rect 12350 3815 12355 3835
rect 12325 3805 12355 3815
rect 12380 3835 12410 3845
rect 12380 3815 12385 3835
rect 12405 3815 12410 3835
rect 12380 3805 12410 3815
rect 12435 3835 12465 3845
rect 12435 3815 12440 3835
rect 12460 3815 12465 3835
rect 12435 3805 12465 3815
rect 12490 3835 12520 3845
rect 12490 3815 12495 3835
rect 12515 3815 12520 3835
rect 12490 3805 12520 3815
rect 12545 3835 12575 3845
rect 12545 3815 12550 3835
rect 12570 3815 12575 3835
rect 12545 3805 12575 3815
rect 12600 3835 12675 3845
rect 12600 3815 12605 3835
rect 12625 3815 12645 3835
rect 12665 3815 12675 3835
rect 12600 3805 12675 3815
rect 11260 3725 11280 3805
rect 11365 3725 11385 3805
rect 11402 3775 11434 3785
rect 11402 3755 11408 3775
rect 11425 3755 11434 3775
rect 11402 3745 11434 3755
rect 11480 3725 11500 3805
rect 11585 3725 11605 3805
rect 11622 3775 11654 3785
rect 11622 3755 11628 3775
rect 11645 3755 11654 3775
rect 11622 3745 11654 3755
rect 11700 3725 11720 3805
rect 11766 3775 11798 3785
rect 11766 3755 11775 3775
rect 11792 3755 11798 3775
rect 11766 3745 11798 3755
rect 11815 3725 11835 3805
rect 12000 3735 12020 3805
rect 11990 3725 12030 3735
rect 11250 3715 11290 3725
rect 11250 3695 11260 3715
rect 11280 3695 11290 3715
rect 11250 3685 11290 3695
rect 11355 3715 11395 3725
rect 11355 3695 11365 3715
rect 11385 3695 11395 3715
rect 11355 3685 11395 3695
rect 11470 3715 11510 3725
rect 11470 3695 11480 3715
rect 11500 3695 11510 3715
rect 11470 3685 11510 3695
rect 11575 3715 11615 3725
rect 11575 3695 11585 3715
rect 11605 3695 11615 3715
rect 11575 3685 11615 3695
rect 11690 3715 11730 3725
rect 11690 3695 11700 3715
rect 11720 3695 11730 3715
rect 11690 3685 11730 3695
rect 11805 3715 11845 3725
rect 11805 3695 11815 3715
rect 11835 3695 11845 3715
rect 11990 3705 12000 3725
rect 12020 3705 12030 3725
rect 11990 3695 12030 3705
rect 11805 3685 11845 3695
rect 12105 3690 12125 3805
rect 12142 3775 12174 3785
rect 12142 3755 12148 3775
rect 12165 3755 12174 3775
rect 12142 3745 12174 3755
rect 12220 3735 12240 3805
rect 12210 3725 12250 3735
rect 12210 3705 12220 3725
rect 12240 3705 12250 3725
rect 12210 3695 12250 3705
rect 12325 3690 12345 3805
rect 12362 3775 12394 3785
rect 12362 3755 12368 3775
rect 12385 3755 12394 3775
rect 12362 3745 12394 3755
rect 12440 3735 12460 3805
rect 12506 3775 12538 3785
rect 12506 3755 12515 3775
rect 12532 3755 12538 3775
rect 12506 3745 12538 3755
rect 12430 3725 12470 3735
rect 12430 3705 12440 3725
rect 12460 3705 12470 3725
rect 12430 3695 12470 3705
rect 12555 3690 12575 3805
rect 12865 3700 12895 3730
rect 12095 3650 12135 3690
rect 12315 3650 12355 3690
rect 12545 3650 12585 3690
rect 12810 3655 12840 3685
rect 10210 3630 10250 3640
rect 10210 3610 10220 3630
rect 10240 3610 10250 3630
rect 10210 3600 10250 3610
rect 10320 3630 10360 3640
rect 10320 3610 10330 3630
rect 10350 3610 10360 3630
rect 10320 3600 10360 3610
rect 10430 3630 10470 3640
rect 10430 3610 10440 3630
rect 10460 3610 10470 3630
rect 10430 3600 10470 3610
rect 10540 3630 10580 3640
rect 10540 3610 10550 3630
rect 10570 3610 10580 3630
rect 10540 3600 10580 3610
rect 10650 3630 10690 3640
rect 10650 3610 10660 3630
rect 10680 3610 10690 3630
rect 10650 3600 10690 3610
rect 10760 3630 10800 3640
rect 13000 3630 13040 3640
rect 10760 3610 10770 3630
rect 10790 3610 10800 3630
rect 10760 3600 10800 3610
rect 11180 3620 11220 3630
rect 11180 3600 11190 3620
rect 11210 3600 11220 3620
rect 10220 3580 10240 3600
rect 10330 3580 10350 3600
rect 10440 3580 10460 3600
rect 10550 3580 10570 3600
rect 10660 3580 10680 3600
rect 10770 3580 10790 3600
rect 11180 3590 11220 3600
rect 11340 3620 11380 3630
rect 11340 3600 11350 3620
rect 11370 3600 11380 3620
rect 11340 3590 11380 3600
rect 11460 3620 11500 3630
rect 11460 3600 11470 3620
rect 11490 3600 11500 3620
rect 11460 3590 11500 3600
rect 11580 3620 11620 3630
rect 11580 3600 11590 3620
rect 11610 3600 11620 3620
rect 11580 3590 11620 3600
rect 11700 3620 11740 3630
rect 11700 3600 11710 3620
rect 11730 3600 11740 3620
rect 11700 3590 11740 3600
rect 11820 3620 11860 3630
rect 11820 3600 11830 3620
rect 11850 3600 11860 3620
rect 11820 3590 11860 3600
rect 11940 3620 11980 3630
rect 11940 3600 11950 3620
rect 11970 3600 11980 3620
rect 11940 3590 11980 3600
rect 12060 3620 12100 3630
rect 12060 3600 12070 3620
rect 12090 3600 12100 3620
rect 12060 3590 12100 3600
rect 12180 3620 12220 3630
rect 12180 3600 12190 3620
rect 12210 3600 12220 3620
rect 12180 3590 12220 3600
rect 12300 3620 12340 3630
rect 12300 3600 12310 3620
rect 12330 3600 12340 3620
rect 12300 3590 12340 3600
rect 12420 3620 12460 3630
rect 12420 3600 12430 3620
rect 12450 3600 12460 3620
rect 12420 3590 12460 3600
rect 12580 3620 12620 3630
rect 12580 3600 12590 3620
rect 12610 3600 12620 3620
rect 13000 3610 13010 3630
rect 13030 3610 13040 3630
rect 13000 3600 13040 3610
rect 13110 3630 13150 3640
rect 13110 3610 13120 3630
rect 13140 3610 13150 3630
rect 13110 3600 13150 3610
rect 13220 3630 13260 3640
rect 13220 3610 13230 3630
rect 13250 3610 13260 3630
rect 13220 3600 13260 3610
rect 13330 3630 13370 3640
rect 13330 3610 13340 3630
rect 13360 3610 13370 3630
rect 13330 3600 13370 3610
rect 13440 3630 13480 3640
rect 13440 3610 13450 3630
rect 13470 3610 13480 3630
rect 13440 3600 13480 3610
rect 13550 3630 13590 3640
rect 13550 3610 13560 3630
rect 13580 3610 13590 3630
rect 26180 3620 26220 3630
rect 13550 3600 13590 3610
rect 25905 3605 26030 3615
rect 12580 3590 12620 3600
rect 10120 3570 10190 3580
rect 1266 3495 1296 3525
rect 9899 3520 10040 3560
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 5145 3415 5175 3445
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 1210 3310 1240 3340
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 5365 3305 5395 3335
rect 10120 3550 10125 3570
rect 10145 3550 10165 3570
rect 10185 3550 10190 3570
rect 10120 3520 10190 3550
rect 10120 3500 10125 3520
rect 10145 3500 10165 3520
rect 10185 3500 10190 3520
rect 10120 3470 10190 3500
rect 10120 3450 10125 3470
rect 10145 3450 10165 3470
rect 10185 3450 10190 3470
rect 10120 3420 10190 3450
rect 10120 3400 10125 3420
rect 10145 3400 10165 3420
rect 10185 3400 10190 3420
rect 10120 3370 10190 3400
rect 10120 3350 10125 3370
rect 10145 3350 10165 3370
rect 10185 3350 10190 3370
rect 10120 3320 10190 3350
rect 10120 3300 10125 3320
rect 10145 3300 10165 3320
rect 10185 3300 10190 3320
rect 1165 3255 1195 3285
rect 4890 3255 4920 3285
rect 5415 3255 5445 3285
rect 10120 3270 10190 3300
rect 10120 3250 10125 3270
rect 10145 3250 10165 3270
rect 10185 3250 10190 3270
rect 2740 3210 2770 3240
rect 10120 3220 10190 3250
rect 46 3200 91 3205
rect 46 3175 56 3200
rect 81 3175 91 3200
rect 46 3170 91 3175
rect 10120 3200 10125 3220
rect 10145 3200 10165 3220
rect 10185 3200 10190 3220
rect 1110 3145 1145 3170
rect 1261 3195 1306 3200
rect 1261 3170 1271 3195
rect 1296 3170 1306 3195
rect 1261 3165 1306 3170
rect 2330 3165 2370 3200
rect 46 3140 91 3145
rect 46 3115 56 3140
rect 81 3115 91 3140
rect 46 3110 91 3115
rect 1261 3135 1306 3140
rect 1261 3110 1271 3135
rect 1296 3110 1306 3135
rect 1261 3105 1306 3110
rect 1165 3070 1195 3100
rect 2295 3080 2330 3105
rect 46 3060 91 3065
rect 46 3035 56 3060
rect 81 3035 91 3060
rect 46 3030 91 3035
rect 1080 3005 1115 3030
rect 46 3000 91 3005
rect 46 2975 56 3000
rect 81 2975 91 3000
rect 46 2970 91 2975
rect 1266 3045 1306 3080
rect 910 2910 1120 2915
rect 910 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1120 2910
rect 910 2875 1120 2880
rect 1266 2900 1286 3045
rect 2350 3020 2370 3165
rect 2625 3155 2655 3185
rect 4445 3155 4475 3185
rect 10120 3170 10190 3200
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 5320 3110 5350 3140
rect 3990 3050 4020 3080
rect 2330 2985 2370 3020
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 1306 2960 1341 2985
rect 2330 2955 2375 2960
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2520 2945 2560 2985
rect 3080 2975 3120 2985
rect 3080 2955 3090 2975
rect 3110 2955 3120 2975
rect 3080 2945 3120 2955
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2975 3305 2985
rect 3265 2955 3275 2975
rect 3295 2955 3305 2975
rect 3265 2945 3305 2955
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2975 3665 2985
rect 3625 2955 3635 2975
rect 3655 2955 3665 2975
rect 3625 2945 3665 2955
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2975 4205 2985
rect 4165 2955 4175 2975
rect 4195 2955 4205 2975
rect 4165 2945 4205 2955
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2975 4565 2985
rect 4525 2955 4535 2975
rect 4555 2955 4565 2975
rect 4525 2945 4565 2955
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 3095 2925 3115 2945
rect 3275 2925 3295 2945
rect 3455 2925 3475 2945
rect 3635 2925 3655 2945
rect 3815 2925 3835 2945
rect 3995 2925 4015 2945
rect 4175 2925 4195 2945
rect 4355 2925 4375 2945
rect 4535 2925 4555 2945
rect 4715 2925 4735 2945
rect 4895 2925 4915 2945
rect 10120 3150 10125 3170
rect 10145 3150 10165 3170
rect 10185 3150 10190 3170
rect 10120 3120 10190 3150
rect 10120 3100 10125 3120
rect 10145 3100 10165 3120
rect 10185 3100 10190 3120
rect 10120 3070 10190 3100
rect 10120 3050 10125 3070
rect 10145 3050 10165 3070
rect 10185 3050 10190 3070
rect 10120 3020 10190 3050
rect 10120 3000 10125 3020
rect 10145 3000 10165 3020
rect 10185 3000 10190 3020
rect 10120 2990 10190 3000
rect 10215 3570 10245 3580
rect 10215 3550 10220 3570
rect 10240 3550 10245 3570
rect 10215 3520 10245 3550
rect 10215 3500 10220 3520
rect 10240 3500 10245 3520
rect 10215 3470 10245 3500
rect 10215 3450 10220 3470
rect 10240 3450 10245 3470
rect 10215 3420 10245 3450
rect 10215 3400 10220 3420
rect 10240 3400 10245 3420
rect 10215 3370 10245 3400
rect 10215 3350 10220 3370
rect 10240 3350 10245 3370
rect 10215 3320 10245 3350
rect 10215 3300 10220 3320
rect 10240 3300 10245 3320
rect 10215 3270 10245 3300
rect 10215 3250 10220 3270
rect 10240 3250 10245 3270
rect 10215 3220 10245 3250
rect 10215 3200 10220 3220
rect 10240 3200 10245 3220
rect 10215 3170 10245 3200
rect 10215 3150 10220 3170
rect 10240 3150 10245 3170
rect 10215 3120 10245 3150
rect 10215 3100 10220 3120
rect 10240 3100 10245 3120
rect 10215 3070 10245 3100
rect 10215 3050 10220 3070
rect 10240 3050 10245 3070
rect 10215 3020 10245 3050
rect 10215 3000 10220 3020
rect 10240 3000 10245 3020
rect 10215 2990 10245 3000
rect 10270 3570 10300 3580
rect 10270 3550 10275 3570
rect 10295 3550 10300 3570
rect 10270 3520 10300 3550
rect 10270 3500 10275 3520
rect 10295 3500 10300 3520
rect 10270 3470 10300 3500
rect 10270 3450 10275 3470
rect 10295 3450 10300 3470
rect 10270 3420 10300 3450
rect 10270 3400 10275 3420
rect 10295 3400 10300 3420
rect 10270 3370 10300 3400
rect 10270 3350 10275 3370
rect 10295 3350 10300 3370
rect 10270 3320 10300 3350
rect 10270 3300 10275 3320
rect 10295 3300 10300 3320
rect 10270 3270 10300 3300
rect 10270 3250 10275 3270
rect 10295 3250 10300 3270
rect 10270 3220 10300 3250
rect 10270 3200 10275 3220
rect 10295 3200 10300 3220
rect 10270 3170 10300 3200
rect 10270 3150 10275 3170
rect 10295 3150 10300 3170
rect 10270 3120 10300 3150
rect 10270 3100 10275 3120
rect 10295 3100 10300 3120
rect 10270 3070 10300 3100
rect 10270 3050 10275 3070
rect 10295 3050 10300 3070
rect 10270 3020 10300 3050
rect 10270 3000 10275 3020
rect 10295 3000 10300 3020
rect 10270 2990 10300 3000
rect 10325 3570 10355 3580
rect 10325 3550 10330 3570
rect 10350 3550 10355 3570
rect 10325 3520 10355 3550
rect 10325 3500 10330 3520
rect 10350 3500 10355 3520
rect 10325 3470 10355 3500
rect 10325 3450 10330 3470
rect 10350 3450 10355 3470
rect 10325 3420 10355 3450
rect 10325 3400 10330 3420
rect 10350 3400 10355 3420
rect 10325 3370 10355 3400
rect 10325 3350 10330 3370
rect 10350 3350 10355 3370
rect 10325 3320 10355 3350
rect 10325 3300 10330 3320
rect 10350 3300 10355 3320
rect 10325 3270 10355 3300
rect 10325 3250 10330 3270
rect 10350 3250 10355 3270
rect 10325 3220 10355 3250
rect 10325 3200 10330 3220
rect 10350 3200 10355 3220
rect 10325 3170 10355 3200
rect 10325 3150 10330 3170
rect 10350 3150 10355 3170
rect 10325 3120 10355 3150
rect 10325 3100 10330 3120
rect 10350 3100 10355 3120
rect 10325 3070 10355 3100
rect 10325 3050 10330 3070
rect 10350 3050 10355 3070
rect 10325 3020 10355 3050
rect 10325 3000 10330 3020
rect 10350 3000 10355 3020
rect 10325 2990 10355 3000
rect 10380 3570 10410 3580
rect 10380 3550 10385 3570
rect 10405 3550 10410 3570
rect 10380 3520 10410 3550
rect 10380 3500 10385 3520
rect 10405 3500 10410 3520
rect 10380 3470 10410 3500
rect 10380 3450 10385 3470
rect 10405 3450 10410 3470
rect 10380 3420 10410 3450
rect 10380 3400 10385 3420
rect 10405 3400 10410 3420
rect 10380 3370 10410 3400
rect 10380 3350 10385 3370
rect 10405 3350 10410 3370
rect 10380 3320 10410 3350
rect 10380 3300 10385 3320
rect 10405 3300 10410 3320
rect 10380 3270 10410 3300
rect 10380 3250 10385 3270
rect 10405 3250 10410 3270
rect 10380 3220 10410 3250
rect 10380 3200 10385 3220
rect 10405 3200 10410 3220
rect 10380 3170 10410 3200
rect 10380 3150 10385 3170
rect 10405 3150 10410 3170
rect 10380 3120 10410 3150
rect 10380 3100 10385 3120
rect 10405 3100 10410 3120
rect 10380 3070 10410 3100
rect 10380 3050 10385 3070
rect 10405 3050 10410 3070
rect 10380 3020 10410 3050
rect 10380 3000 10385 3020
rect 10405 3000 10410 3020
rect 10380 2990 10410 3000
rect 10435 3570 10465 3580
rect 10435 3550 10440 3570
rect 10460 3550 10465 3570
rect 10435 3520 10465 3550
rect 10435 3500 10440 3520
rect 10460 3500 10465 3520
rect 10435 3470 10465 3500
rect 10435 3450 10440 3470
rect 10460 3450 10465 3470
rect 10435 3420 10465 3450
rect 10435 3400 10440 3420
rect 10460 3400 10465 3420
rect 10435 3370 10465 3400
rect 10435 3350 10440 3370
rect 10460 3350 10465 3370
rect 10435 3320 10465 3350
rect 10435 3300 10440 3320
rect 10460 3300 10465 3320
rect 10435 3270 10465 3300
rect 10435 3250 10440 3270
rect 10460 3250 10465 3270
rect 10435 3220 10465 3250
rect 10435 3200 10440 3220
rect 10460 3200 10465 3220
rect 10435 3170 10465 3200
rect 10435 3150 10440 3170
rect 10460 3150 10465 3170
rect 10435 3120 10465 3150
rect 10435 3100 10440 3120
rect 10460 3100 10465 3120
rect 10435 3070 10465 3100
rect 10435 3050 10440 3070
rect 10460 3050 10465 3070
rect 10435 3020 10465 3050
rect 10435 3000 10440 3020
rect 10460 3000 10465 3020
rect 10435 2990 10465 3000
rect 10490 3570 10520 3580
rect 10490 3550 10495 3570
rect 10515 3550 10520 3570
rect 10490 3520 10520 3550
rect 10490 3500 10495 3520
rect 10515 3500 10520 3520
rect 10490 3470 10520 3500
rect 10490 3450 10495 3470
rect 10515 3450 10520 3470
rect 10490 3420 10520 3450
rect 10490 3400 10495 3420
rect 10515 3400 10520 3420
rect 10490 3370 10520 3400
rect 10490 3350 10495 3370
rect 10515 3350 10520 3370
rect 10490 3320 10520 3350
rect 10490 3300 10495 3320
rect 10515 3300 10520 3320
rect 10490 3270 10520 3300
rect 10490 3250 10495 3270
rect 10515 3250 10520 3270
rect 10490 3220 10520 3250
rect 10490 3200 10495 3220
rect 10515 3200 10520 3220
rect 10490 3170 10520 3200
rect 10490 3150 10495 3170
rect 10515 3150 10520 3170
rect 10490 3120 10520 3150
rect 10490 3100 10495 3120
rect 10515 3100 10520 3120
rect 10490 3070 10520 3100
rect 10490 3050 10495 3070
rect 10515 3050 10520 3070
rect 10490 3020 10520 3050
rect 10490 3000 10495 3020
rect 10515 3000 10520 3020
rect 10490 2990 10520 3000
rect 10545 3570 10575 3580
rect 10545 3550 10550 3570
rect 10570 3550 10575 3570
rect 10545 3520 10575 3550
rect 10545 3500 10550 3520
rect 10570 3500 10575 3520
rect 10545 3470 10575 3500
rect 10545 3450 10550 3470
rect 10570 3450 10575 3470
rect 10545 3420 10575 3450
rect 10545 3400 10550 3420
rect 10570 3400 10575 3420
rect 10545 3370 10575 3400
rect 10545 3350 10550 3370
rect 10570 3350 10575 3370
rect 10545 3320 10575 3350
rect 10545 3300 10550 3320
rect 10570 3300 10575 3320
rect 10545 3270 10575 3300
rect 10545 3250 10550 3270
rect 10570 3250 10575 3270
rect 10545 3220 10575 3250
rect 10545 3200 10550 3220
rect 10570 3200 10575 3220
rect 10545 3170 10575 3200
rect 10545 3150 10550 3170
rect 10570 3150 10575 3170
rect 10545 3120 10575 3150
rect 10545 3100 10550 3120
rect 10570 3100 10575 3120
rect 10545 3070 10575 3100
rect 10545 3050 10550 3070
rect 10570 3050 10575 3070
rect 10545 3020 10575 3050
rect 10545 3000 10550 3020
rect 10570 3000 10575 3020
rect 10545 2990 10575 3000
rect 10600 3570 10630 3580
rect 10600 3550 10605 3570
rect 10625 3550 10630 3570
rect 10600 3520 10630 3550
rect 10600 3500 10605 3520
rect 10625 3500 10630 3520
rect 10600 3470 10630 3500
rect 10600 3450 10605 3470
rect 10625 3450 10630 3470
rect 10600 3420 10630 3450
rect 10600 3400 10605 3420
rect 10625 3400 10630 3420
rect 10600 3370 10630 3400
rect 10600 3350 10605 3370
rect 10625 3350 10630 3370
rect 10600 3320 10630 3350
rect 10600 3300 10605 3320
rect 10625 3300 10630 3320
rect 10600 3270 10630 3300
rect 10600 3250 10605 3270
rect 10625 3250 10630 3270
rect 10600 3220 10630 3250
rect 10600 3200 10605 3220
rect 10625 3200 10630 3220
rect 10600 3170 10630 3200
rect 10600 3150 10605 3170
rect 10625 3150 10630 3170
rect 10600 3120 10630 3150
rect 10600 3100 10605 3120
rect 10625 3100 10630 3120
rect 10600 3070 10630 3100
rect 10600 3050 10605 3070
rect 10625 3050 10630 3070
rect 10600 3020 10630 3050
rect 10600 3000 10605 3020
rect 10625 3000 10630 3020
rect 10600 2990 10630 3000
rect 10655 3570 10685 3580
rect 10655 3550 10660 3570
rect 10680 3550 10685 3570
rect 10655 3520 10685 3550
rect 10655 3500 10660 3520
rect 10680 3500 10685 3520
rect 10655 3470 10685 3500
rect 10655 3450 10660 3470
rect 10680 3450 10685 3470
rect 10655 3420 10685 3450
rect 10655 3400 10660 3420
rect 10680 3400 10685 3420
rect 10655 3370 10685 3400
rect 10655 3350 10660 3370
rect 10680 3350 10685 3370
rect 10655 3320 10685 3350
rect 10655 3300 10660 3320
rect 10680 3300 10685 3320
rect 10655 3270 10685 3300
rect 10655 3250 10660 3270
rect 10680 3250 10685 3270
rect 10655 3220 10685 3250
rect 10655 3200 10660 3220
rect 10680 3200 10685 3220
rect 10655 3170 10685 3200
rect 10655 3150 10660 3170
rect 10680 3150 10685 3170
rect 10655 3120 10685 3150
rect 10655 3100 10660 3120
rect 10680 3100 10685 3120
rect 10655 3070 10685 3100
rect 10655 3050 10660 3070
rect 10680 3050 10685 3070
rect 10655 3020 10685 3050
rect 10655 3000 10660 3020
rect 10680 3000 10685 3020
rect 10655 2990 10685 3000
rect 10710 3570 10740 3580
rect 10710 3550 10715 3570
rect 10735 3550 10740 3570
rect 10710 3520 10740 3550
rect 10710 3500 10715 3520
rect 10735 3500 10740 3520
rect 10710 3470 10740 3500
rect 10710 3450 10715 3470
rect 10735 3450 10740 3470
rect 10710 3420 10740 3450
rect 10710 3400 10715 3420
rect 10735 3400 10740 3420
rect 10710 3370 10740 3400
rect 10710 3350 10715 3370
rect 10735 3350 10740 3370
rect 10710 3320 10740 3350
rect 10710 3300 10715 3320
rect 10735 3300 10740 3320
rect 10710 3270 10740 3300
rect 10710 3250 10715 3270
rect 10735 3250 10740 3270
rect 10710 3220 10740 3250
rect 10710 3200 10715 3220
rect 10735 3200 10740 3220
rect 10710 3170 10740 3200
rect 10710 3150 10715 3170
rect 10735 3150 10740 3170
rect 10710 3120 10740 3150
rect 10710 3100 10715 3120
rect 10735 3100 10740 3120
rect 10710 3070 10740 3100
rect 10710 3050 10715 3070
rect 10735 3050 10740 3070
rect 10710 3020 10740 3050
rect 10710 3000 10715 3020
rect 10735 3000 10740 3020
rect 10710 2990 10740 3000
rect 10765 3570 10795 3580
rect 10765 3550 10770 3570
rect 10790 3550 10795 3570
rect 10765 3520 10795 3550
rect 10765 3500 10770 3520
rect 10790 3500 10795 3520
rect 10765 3470 10795 3500
rect 10765 3450 10770 3470
rect 10790 3450 10795 3470
rect 10765 3420 10795 3450
rect 10765 3400 10770 3420
rect 10790 3400 10795 3420
rect 10765 3370 10795 3400
rect 10765 3350 10770 3370
rect 10790 3350 10795 3370
rect 10765 3320 10795 3350
rect 10765 3300 10770 3320
rect 10790 3300 10795 3320
rect 10765 3270 10795 3300
rect 10765 3250 10770 3270
rect 10790 3250 10795 3270
rect 10765 3220 10795 3250
rect 10765 3200 10770 3220
rect 10790 3200 10795 3220
rect 10765 3170 10795 3200
rect 10765 3150 10770 3170
rect 10790 3150 10795 3170
rect 10765 3120 10795 3150
rect 10765 3100 10770 3120
rect 10790 3100 10795 3120
rect 10765 3070 10795 3100
rect 10765 3050 10770 3070
rect 10790 3050 10795 3070
rect 10765 3020 10795 3050
rect 10765 3000 10770 3020
rect 10790 3000 10795 3020
rect 10765 2990 10795 3000
rect 10820 3570 10890 3580
rect 11190 3570 11210 3590
rect 11350 3570 11370 3590
rect 11470 3570 11490 3590
rect 11590 3570 11610 3590
rect 11710 3570 11730 3590
rect 11830 3570 11850 3590
rect 11950 3570 11970 3590
rect 12070 3570 12090 3590
rect 12190 3570 12210 3590
rect 12310 3570 12330 3590
rect 12430 3570 12450 3590
rect 12590 3570 12610 3590
rect 13010 3580 13030 3600
rect 13120 3580 13140 3600
rect 13230 3580 13250 3600
rect 13340 3580 13360 3600
rect 13450 3580 13470 3600
rect 13560 3580 13580 3600
rect 25905 3585 25915 3605
rect 25935 3595 26030 3605
rect 25935 3585 25945 3595
rect 12910 3570 12980 3580
rect 10820 3550 10825 3570
rect 10845 3550 10865 3570
rect 10885 3550 10890 3570
rect 10820 3520 10890 3550
rect 10820 3500 10825 3520
rect 10845 3500 10865 3520
rect 10885 3500 10890 3520
rect 10820 3470 10890 3500
rect 10820 3450 10825 3470
rect 10845 3450 10865 3470
rect 10885 3450 10890 3470
rect 10820 3420 10890 3450
rect 10820 3400 10825 3420
rect 10845 3400 10865 3420
rect 10885 3400 10890 3420
rect 10820 3370 10890 3400
rect 10820 3350 10825 3370
rect 10845 3350 10865 3370
rect 10885 3350 10890 3370
rect 10820 3320 10890 3350
rect 10820 3300 10825 3320
rect 10845 3300 10865 3320
rect 10885 3300 10890 3320
rect 10820 3270 10890 3300
rect 10820 3250 10825 3270
rect 10845 3250 10865 3270
rect 10885 3250 10890 3270
rect 10820 3220 10890 3250
rect 10820 3200 10825 3220
rect 10845 3200 10865 3220
rect 10885 3200 10890 3220
rect 10820 3170 10890 3200
rect 11185 3560 11255 3570
rect 11185 3540 11190 3560
rect 11210 3540 11230 3560
rect 11250 3540 11255 3560
rect 11185 3510 11255 3540
rect 11185 3490 11190 3510
rect 11210 3490 11230 3510
rect 11250 3490 11255 3510
rect 11185 3460 11255 3490
rect 11185 3440 11190 3460
rect 11210 3440 11230 3460
rect 11250 3440 11255 3460
rect 11185 3410 11255 3440
rect 11185 3390 11190 3410
rect 11210 3390 11230 3410
rect 11250 3390 11255 3410
rect 11185 3360 11255 3390
rect 11185 3340 11190 3360
rect 11210 3340 11230 3360
rect 11250 3340 11255 3360
rect 11185 3310 11255 3340
rect 11185 3290 11190 3310
rect 11210 3290 11230 3310
rect 11250 3290 11255 3310
rect 11185 3260 11255 3290
rect 11185 3240 11190 3260
rect 11210 3240 11230 3260
rect 11250 3240 11255 3260
rect 11185 3210 11255 3240
rect 11185 3190 11190 3210
rect 11210 3190 11230 3210
rect 11250 3190 11255 3210
rect 11185 3180 11255 3190
rect 11285 3560 11315 3570
rect 11285 3540 11290 3560
rect 11310 3540 11315 3560
rect 11285 3510 11315 3540
rect 11285 3490 11290 3510
rect 11310 3490 11315 3510
rect 11285 3460 11315 3490
rect 11285 3440 11290 3460
rect 11310 3440 11315 3460
rect 11285 3410 11315 3440
rect 11285 3390 11290 3410
rect 11310 3390 11315 3410
rect 11285 3360 11315 3390
rect 11285 3340 11290 3360
rect 11310 3340 11315 3360
rect 11285 3310 11315 3340
rect 11285 3290 11290 3310
rect 11310 3290 11315 3310
rect 11285 3260 11315 3290
rect 11285 3240 11290 3260
rect 11310 3240 11315 3260
rect 11285 3210 11315 3240
rect 11285 3190 11290 3210
rect 11310 3190 11315 3210
rect 11285 3180 11315 3190
rect 11345 3560 11375 3570
rect 11345 3540 11350 3560
rect 11370 3540 11375 3560
rect 11345 3510 11375 3540
rect 11345 3490 11350 3510
rect 11370 3490 11375 3510
rect 11345 3460 11375 3490
rect 11345 3440 11350 3460
rect 11370 3440 11375 3460
rect 11345 3410 11375 3440
rect 11345 3390 11350 3410
rect 11370 3390 11375 3410
rect 11345 3360 11375 3390
rect 11345 3340 11350 3360
rect 11370 3340 11375 3360
rect 11345 3310 11375 3340
rect 11345 3290 11350 3310
rect 11370 3290 11375 3310
rect 11345 3260 11375 3290
rect 11345 3240 11350 3260
rect 11370 3240 11375 3260
rect 11345 3210 11375 3240
rect 11345 3190 11350 3210
rect 11370 3190 11375 3210
rect 11345 3180 11375 3190
rect 11405 3560 11435 3570
rect 11405 3540 11410 3560
rect 11430 3540 11435 3560
rect 11405 3510 11435 3540
rect 11405 3490 11410 3510
rect 11430 3490 11435 3510
rect 11405 3460 11435 3490
rect 11405 3440 11410 3460
rect 11430 3440 11435 3460
rect 11405 3410 11435 3440
rect 11405 3390 11410 3410
rect 11430 3390 11435 3410
rect 11405 3360 11435 3390
rect 11405 3340 11410 3360
rect 11430 3340 11435 3360
rect 11405 3310 11435 3340
rect 11405 3290 11410 3310
rect 11430 3290 11435 3310
rect 11405 3260 11435 3290
rect 11405 3240 11410 3260
rect 11430 3240 11435 3260
rect 11405 3210 11435 3240
rect 11405 3190 11410 3210
rect 11430 3190 11435 3210
rect 11405 3180 11435 3190
rect 11465 3560 11495 3570
rect 11465 3540 11470 3560
rect 11490 3540 11495 3560
rect 11465 3510 11495 3540
rect 11465 3490 11470 3510
rect 11490 3490 11495 3510
rect 11465 3460 11495 3490
rect 11465 3440 11470 3460
rect 11490 3440 11495 3460
rect 11465 3410 11495 3440
rect 11465 3390 11470 3410
rect 11490 3390 11495 3410
rect 11465 3360 11495 3390
rect 11465 3340 11470 3360
rect 11490 3340 11495 3360
rect 11465 3310 11495 3340
rect 11465 3290 11470 3310
rect 11490 3290 11495 3310
rect 11465 3260 11495 3290
rect 11465 3240 11470 3260
rect 11490 3240 11495 3260
rect 11465 3210 11495 3240
rect 11465 3190 11470 3210
rect 11490 3190 11495 3210
rect 11465 3180 11495 3190
rect 11525 3560 11555 3570
rect 11525 3540 11530 3560
rect 11550 3540 11555 3560
rect 11525 3510 11555 3540
rect 11525 3490 11530 3510
rect 11550 3490 11555 3510
rect 11525 3460 11555 3490
rect 11525 3440 11530 3460
rect 11550 3440 11555 3460
rect 11525 3410 11555 3440
rect 11525 3390 11530 3410
rect 11550 3390 11555 3410
rect 11525 3360 11555 3390
rect 11525 3340 11530 3360
rect 11550 3340 11555 3360
rect 11525 3310 11555 3340
rect 11525 3290 11530 3310
rect 11550 3290 11555 3310
rect 11525 3260 11555 3290
rect 11525 3240 11530 3260
rect 11550 3240 11555 3260
rect 11525 3210 11555 3240
rect 11525 3190 11530 3210
rect 11550 3190 11555 3210
rect 11525 3180 11555 3190
rect 11585 3560 11615 3570
rect 11585 3540 11590 3560
rect 11610 3540 11615 3560
rect 11585 3510 11615 3540
rect 11585 3490 11590 3510
rect 11610 3490 11615 3510
rect 11585 3460 11615 3490
rect 11585 3440 11590 3460
rect 11610 3440 11615 3460
rect 11585 3410 11615 3440
rect 11585 3390 11590 3410
rect 11610 3390 11615 3410
rect 11585 3360 11615 3390
rect 11585 3340 11590 3360
rect 11610 3340 11615 3360
rect 11585 3310 11615 3340
rect 11585 3290 11590 3310
rect 11610 3290 11615 3310
rect 11585 3260 11615 3290
rect 11585 3240 11590 3260
rect 11610 3240 11615 3260
rect 11585 3210 11615 3240
rect 11585 3190 11590 3210
rect 11610 3190 11615 3210
rect 11585 3180 11615 3190
rect 11645 3560 11675 3570
rect 11645 3540 11650 3560
rect 11670 3540 11675 3560
rect 11645 3510 11675 3540
rect 11645 3490 11650 3510
rect 11670 3490 11675 3510
rect 11645 3460 11675 3490
rect 11645 3440 11650 3460
rect 11670 3440 11675 3460
rect 11645 3410 11675 3440
rect 11645 3390 11650 3410
rect 11670 3390 11675 3410
rect 11645 3360 11675 3390
rect 11645 3340 11650 3360
rect 11670 3340 11675 3360
rect 11645 3310 11675 3340
rect 11645 3290 11650 3310
rect 11670 3290 11675 3310
rect 11645 3260 11675 3290
rect 11645 3240 11650 3260
rect 11670 3240 11675 3260
rect 11645 3210 11675 3240
rect 11645 3190 11650 3210
rect 11670 3190 11675 3210
rect 11645 3180 11675 3190
rect 11705 3560 11735 3570
rect 11705 3540 11710 3560
rect 11730 3540 11735 3560
rect 11705 3510 11735 3540
rect 11705 3490 11710 3510
rect 11730 3490 11735 3510
rect 11705 3460 11735 3490
rect 11705 3440 11710 3460
rect 11730 3440 11735 3460
rect 11705 3410 11735 3440
rect 11705 3390 11710 3410
rect 11730 3390 11735 3410
rect 11705 3360 11735 3390
rect 11705 3340 11710 3360
rect 11730 3340 11735 3360
rect 11705 3310 11735 3340
rect 11705 3290 11710 3310
rect 11730 3290 11735 3310
rect 11705 3260 11735 3290
rect 11705 3240 11710 3260
rect 11730 3240 11735 3260
rect 11705 3210 11735 3240
rect 11705 3190 11710 3210
rect 11730 3190 11735 3210
rect 11705 3180 11735 3190
rect 11765 3560 11795 3570
rect 11765 3540 11770 3560
rect 11790 3540 11795 3560
rect 11765 3510 11795 3540
rect 11765 3490 11770 3510
rect 11790 3490 11795 3510
rect 11765 3460 11795 3490
rect 11765 3440 11770 3460
rect 11790 3440 11795 3460
rect 11765 3410 11795 3440
rect 11765 3390 11770 3410
rect 11790 3390 11795 3410
rect 11765 3360 11795 3390
rect 11765 3340 11770 3360
rect 11790 3340 11795 3360
rect 11765 3310 11795 3340
rect 11765 3290 11770 3310
rect 11790 3290 11795 3310
rect 11765 3260 11795 3290
rect 11765 3240 11770 3260
rect 11790 3240 11795 3260
rect 11765 3210 11795 3240
rect 11765 3190 11770 3210
rect 11790 3190 11795 3210
rect 11765 3180 11795 3190
rect 11825 3560 11855 3570
rect 11825 3540 11830 3560
rect 11850 3540 11855 3560
rect 11825 3510 11855 3540
rect 11825 3490 11830 3510
rect 11850 3490 11855 3510
rect 11825 3460 11855 3490
rect 11825 3440 11830 3460
rect 11850 3440 11855 3460
rect 11825 3410 11855 3440
rect 11825 3390 11830 3410
rect 11850 3390 11855 3410
rect 11825 3360 11855 3390
rect 11825 3340 11830 3360
rect 11850 3340 11855 3360
rect 11825 3310 11855 3340
rect 11825 3290 11830 3310
rect 11850 3290 11855 3310
rect 11825 3260 11855 3290
rect 11825 3240 11830 3260
rect 11850 3240 11855 3260
rect 11825 3210 11855 3240
rect 11825 3190 11830 3210
rect 11850 3190 11855 3210
rect 11825 3180 11855 3190
rect 11885 3560 11915 3570
rect 11885 3540 11890 3560
rect 11910 3540 11915 3560
rect 11885 3510 11915 3540
rect 11885 3490 11890 3510
rect 11910 3490 11915 3510
rect 11885 3460 11915 3490
rect 11885 3440 11890 3460
rect 11910 3440 11915 3460
rect 11885 3410 11915 3440
rect 11885 3390 11890 3410
rect 11910 3390 11915 3410
rect 11885 3360 11915 3390
rect 11885 3340 11890 3360
rect 11910 3340 11915 3360
rect 11885 3310 11915 3340
rect 11885 3290 11890 3310
rect 11910 3290 11915 3310
rect 11885 3260 11915 3290
rect 11885 3240 11890 3260
rect 11910 3240 11915 3260
rect 11885 3210 11915 3240
rect 11885 3190 11890 3210
rect 11910 3190 11915 3210
rect 11885 3180 11915 3190
rect 11945 3560 11975 3570
rect 11945 3540 11950 3560
rect 11970 3540 11975 3560
rect 11945 3510 11975 3540
rect 11945 3490 11950 3510
rect 11970 3490 11975 3510
rect 11945 3460 11975 3490
rect 11945 3440 11950 3460
rect 11970 3440 11975 3460
rect 11945 3410 11975 3440
rect 11945 3390 11950 3410
rect 11970 3390 11975 3410
rect 11945 3360 11975 3390
rect 11945 3340 11950 3360
rect 11970 3340 11975 3360
rect 11945 3310 11975 3340
rect 11945 3290 11950 3310
rect 11970 3290 11975 3310
rect 11945 3260 11975 3290
rect 11945 3240 11950 3260
rect 11970 3240 11975 3260
rect 11945 3210 11975 3240
rect 11945 3190 11950 3210
rect 11970 3190 11975 3210
rect 11945 3180 11975 3190
rect 12005 3560 12035 3570
rect 12005 3540 12010 3560
rect 12030 3540 12035 3560
rect 12005 3510 12035 3540
rect 12005 3490 12010 3510
rect 12030 3490 12035 3510
rect 12005 3460 12035 3490
rect 12005 3440 12010 3460
rect 12030 3440 12035 3460
rect 12005 3410 12035 3440
rect 12005 3390 12010 3410
rect 12030 3390 12035 3410
rect 12005 3360 12035 3390
rect 12005 3340 12010 3360
rect 12030 3340 12035 3360
rect 12005 3310 12035 3340
rect 12005 3290 12010 3310
rect 12030 3290 12035 3310
rect 12005 3260 12035 3290
rect 12005 3240 12010 3260
rect 12030 3240 12035 3260
rect 12005 3210 12035 3240
rect 12005 3190 12010 3210
rect 12030 3190 12035 3210
rect 12005 3180 12035 3190
rect 12065 3560 12095 3570
rect 12065 3540 12070 3560
rect 12090 3540 12095 3560
rect 12065 3510 12095 3540
rect 12065 3490 12070 3510
rect 12090 3490 12095 3510
rect 12065 3460 12095 3490
rect 12065 3440 12070 3460
rect 12090 3440 12095 3460
rect 12065 3410 12095 3440
rect 12065 3390 12070 3410
rect 12090 3390 12095 3410
rect 12065 3360 12095 3390
rect 12065 3340 12070 3360
rect 12090 3340 12095 3360
rect 12065 3310 12095 3340
rect 12065 3290 12070 3310
rect 12090 3290 12095 3310
rect 12065 3260 12095 3290
rect 12065 3240 12070 3260
rect 12090 3240 12095 3260
rect 12065 3210 12095 3240
rect 12065 3190 12070 3210
rect 12090 3190 12095 3210
rect 12065 3180 12095 3190
rect 12125 3560 12155 3570
rect 12125 3540 12130 3560
rect 12150 3540 12155 3560
rect 12125 3510 12155 3540
rect 12125 3490 12130 3510
rect 12150 3490 12155 3510
rect 12125 3460 12155 3490
rect 12125 3440 12130 3460
rect 12150 3440 12155 3460
rect 12125 3410 12155 3440
rect 12125 3390 12130 3410
rect 12150 3390 12155 3410
rect 12125 3360 12155 3390
rect 12125 3340 12130 3360
rect 12150 3340 12155 3360
rect 12125 3310 12155 3340
rect 12125 3290 12130 3310
rect 12150 3290 12155 3310
rect 12125 3260 12155 3290
rect 12125 3240 12130 3260
rect 12150 3240 12155 3260
rect 12125 3210 12155 3240
rect 12125 3190 12130 3210
rect 12150 3190 12155 3210
rect 12125 3180 12155 3190
rect 12185 3560 12215 3570
rect 12185 3540 12190 3560
rect 12210 3540 12215 3560
rect 12185 3510 12215 3540
rect 12185 3490 12190 3510
rect 12210 3490 12215 3510
rect 12185 3460 12215 3490
rect 12185 3440 12190 3460
rect 12210 3440 12215 3460
rect 12185 3410 12215 3440
rect 12185 3390 12190 3410
rect 12210 3390 12215 3410
rect 12185 3360 12215 3390
rect 12185 3340 12190 3360
rect 12210 3340 12215 3360
rect 12185 3310 12215 3340
rect 12185 3290 12190 3310
rect 12210 3290 12215 3310
rect 12185 3260 12215 3290
rect 12185 3240 12190 3260
rect 12210 3240 12215 3260
rect 12185 3210 12215 3240
rect 12185 3190 12190 3210
rect 12210 3190 12215 3210
rect 12185 3180 12215 3190
rect 12245 3560 12275 3570
rect 12245 3540 12250 3560
rect 12270 3540 12275 3560
rect 12245 3510 12275 3540
rect 12245 3490 12250 3510
rect 12270 3490 12275 3510
rect 12245 3460 12275 3490
rect 12245 3440 12250 3460
rect 12270 3440 12275 3460
rect 12245 3410 12275 3440
rect 12245 3390 12250 3410
rect 12270 3390 12275 3410
rect 12245 3360 12275 3390
rect 12245 3340 12250 3360
rect 12270 3340 12275 3360
rect 12245 3310 12275 3340
rect 12245 3290 12250 3310
rect 12270 3290 12275 3310
rect 12245 3260 12275 3290
rect 12245 3240 12250 3260
rect 12270 3240 12275 3260
rect 12245 3210 12275 3240
rect 12245 3190 12250 3210
rect 12270 3190 12275 3210
rect 12245 3180 12275 3190
rect 12305 3560 12335 3570
rect 12305 3540 12310 3560
rect 12330 3540 12335 3560
rect 12305 3510 12335 3540
rect 12305 3490 12310 3510
rect 12330 3490 12335 3510
rect 12305 3460 12335 3490
rect 12305 3440 12310 3460
rect 12330 3440 12335 3460
rect 12305 3410 12335 3440
rect 12305 3390 12310 3410
rect 12330 3390 12335 3410
rect 12305 3360 12335 3390
rect 12305 3340 12310 3360
rect 12330 3340 12335 3360
rect 12305 3310 12335 3340
rect 12305 3290 12310 3310
rect 12330 3290 12335 3310
rect 12305 3260 12335 3290
rect 12305 3240 12310 3260
rect 12330 3240 12335 3260
rect 12305 3210 12335 3240
rect 12305 3190 12310 3210
rect 12330 3190 12335 3210
rect 12305 3180 12335 3190
rect 12365 3560 12395 3570
rect 12365 3540 12370 3560
rect 12390 3540 12395 3560
rect 12365 3510 12395 3540
rect 12365 3490 12370 3510
rect 12390 3490 12395 3510
rect 12365 3460 12395 3490
rect 12365 3440 12370 3460
rect 12390 3440 12395 3460
rect 12365 3410 12395 3440
rect 12365 3390 12370 3410
rect 12390 3390 12395 3410
rect 12365 3360 12395 3390
rect 12365 3340 12370 3360
rect 12390 3340 12395 3360
rect 12365 3310 12395 3340
rect 12365 3290 12370 3310
rect 12390 3290 12395 3310
rect 12365 3260 12395 3290
rect 12365 3240 12370 3260
rect 12390 3240 12395 3260
rect 12365 3210 12395 3240
rect 12365 3190 12370 3210
rect 12390 3190 12395 3210
rect 12365 3180 12395 3190
rect 12425 3560 12455 3570
rect 12425 3540 12430 3560
rect 12450 3540 12455 3560
rect 12425 3510 12455 3540
rect 12425 3490 12430 3510
rect 12450 3490 12455 3510
rect 12425 3460 12455 3490
rect 12425 3440 12430 3460
rect 12450 3440 12455 3460
rect 12425 3410 12455 3440
rect 12425 3390 12430 3410
rect 12450 3390 12455 3410
rect 12425 3360 12455 3390
rect 12425 3340 12430 3360
rect 12450 3340 12455 3360
rect 12425 3310 12455 3340
rect 12425 3290 12430 3310
rect 12450 3290 12455 3310
rect 12425 3260 12455 3290
rect 12425 3240 12430 3260
rect 12450 3240 12455 3260
rect 12425 3210 12455 3240
rect 12425 3190 12430 3210
rect 12450 3190 12455 3210
rect 12425 3180 12455 3190
rect 12485 3560 12515 3570
rect 12485 3540 12490 3560
rect 12510 3540 12515 3560
rect 12485 3510 12515 3540
rect 12485 3490 12490 3510
rect 12510 3490 12515 3510
rect 12485 3460 12515 3490
rect 12485 3440 12490 3460
rect 12510 3440 12515 3460
rect 12485 3410 12515 3440
rect 12485 3390 12490 3410
rect 12510 3390 12515 3410
rect 12485 3360 12515 3390
rect 12485 3340 12490 3360
rect 12510 3340 12515 3360
rect 12485 3310 12515 3340
rect 12485 3290 12490 3310
rect 12510 3290 12515 3310
rect 12485 3260 12515 3290
rect 12485 3240 12490 3260
rect 12510 3240 12515 3260
rect 12485 3210 12515 3240
rect 12485 3190 12490 3210
rect 12510 3190 12515 3210
rect 12485 3180 12515 3190
rect 12545 3560 12615 3570
rect 12545 3540 12550 3560
rect 12570 3540 12590 3560
rect 12610 3540 12615 3560
rect 12545 3510 12615 3540
rect 12545 3490 12550 3510
rect 12570 3490 12590 3510
rect 12610 3490 12615 3510
rect 12545 3460 12615 3490
rect 12545 3440 12550 3460
rect 12570 3440 12590 3460
rect 12610 3440 12615 3460
rect 12545 3410 12615 3440
rect 12545 3390 12550 3410
rect 12570 3390 12590 3410
rect 12610 3390 12615 3410
rect 12545 3360 12615 3390
rect 12545 3340 12550 3360
rect 12570 3340 12590 3360
rect 12610 3340 12615 3360
rect 12545 3310 12615 3340
rect 12545 3290 12550 3310
rect 12570 3290 12590 3310
rect 12610 3290 12615 3310
rect 12545 3260 12615 3290
rect 12545 3240 12550 3260
rect 12570 3240 12590 3260
rect 12610 3240 12615 3260
rect 12545 3210 12615 3240
rect 12545 3190 12550 3210
rect 12570 3190 12590 3210
rect 12610 3190 12615 3210
rect 12545 3180 12615 3190
rect 12910 3550 12915 3570
rect 12935 3550 12955 3570
rect 12975 3550 12980 3570
rect 12910 3520 12980 3550
rect 12910 3500 12915 3520
rect 12935 3500 12955 3520
rect 12975 3500 12980 3520
rect 12910 3470 12980 3500
rect 12910 3450 12915 3470
rect 12935 3450 12955 3470
rect 12975 3450 12980 3470
rect 12910 3420 12980 3450
rect 12910 3400 12915 3420
rect 12935 3400 12955 3420
rect 12975 3400 12980 3420
rect 12910 3370 12980 3400
rect 12910 3350 12915 3370
rect 12935 3350 12955 3370
rect 12975 3350 12980 3370
rect 12910 3320 12980 3350
rect 12910 3300 12915 3320
rect 12935 3300 12955 3320
rect 12975 3300 12980 3320
rect 12910 3270 12980 3300
rect 12910 3250 12915 3270
rect 12935 3250 12955 3270
rect 12975 3250 12980 3270
rect 12910 3220 12980 3250
rect 12910 3200 12915 3220
rect 12935 3200 12955 3220
rect 12975 3200 12980 3220
rect 10820 3150 10825 3170
rect 10845 3150 10865 3170
rect 10885 3150 10890 3170
rect 11290 3160 11310 3180
rect 11410 3160 11430 3180
rect 11530 3160 11550 3180
rect 11650 3160 11670 3180
rect 11770 3160 11790 3180
rect 11890 3160 11910 3180
rect 12010 3160 12030 3180
rect 12130 3160 12150 3180
rect 12250 3160 12270 3180
rect 12370 3160 12390 3180
rect 12490 3160 12510 3180
rect 12910 3170 12980 3200
rect 10820 3120 10890 3150
rect 11280 3150 11320 3160
rect 11280 3130 11290 3150
rect 11310 3130 11320 3150
rect 11280 3120 11320 3130
rect 11400 3150 11440 3160
rect 11400 3130 11410 3150
rect 11430 3130 11440 3150
rect 11400 3120 11440 3130
rect 11520 3150 11560 3160
rect 11520 3130 11530 3150
rect 11550 3130 11560 3150
rect 11520 3120 11560 3130
rect 11640 3150 11680 3160
rect 11640 3130 11650 3150
rect 11670 3130 11680 3150
rect 11640 3120 11680 3130
rect 11760 3150 11800 3160
rect 11760 3130 11770 3150
rect 11790 3130 11800 3150
rect 11760 3120 11800 3130
rect 11823 3150 11857 3160
rect 11823 3130 11831 3150
rect 11849 3130 11857 3150
rect 11823 3120 11857 3130
rect 11880 3150 11920 3160
rect 11880 3130 11890 3150
rect 11910 3130 11920 3150
rect 11880 3120 11920 3130
rect 12000 3150 12040 3160
rect 12000 3130 12010 3150
rect 12030 3130 12040 3150
rect 12000 3120 12040 3130
rect 12120 3150 12160 3160
rect 12120 3130 12130 3150
rect 12150 3130 12160 3150
rect 12120 3120 12160 3130
rect 12240 3150 12280 3160
rect 12240 3130 12250 3150
rect 12270 3130 12280 3150
rect 12240 3120 12280 3130
rect 12360 3150 12400 3160
rect 12360 3130 12370 3150
rect 12390 3130 12400 3150
rect 12360 3120 12400 3130
rect 12480 3150 12520 3160
rect 12480 3130 12490 3150
rect 12510 3130 12520 3150
rect 12480 3120 12520 3130
rect 12910 3150 12915 3170
rect 12935 3150 12955 3170
rect 12975 3150 12980 3170
rect 12910 3120 12980 3150
rect 10820 3100 10825 3120
rect 10845 3100 10865 3120
rect 10885 3100 10890 3120
rect 10820 3070 10890 3100
rect 10820 3050 10825 3070
rect 10845 3050 10865 3070
rect 10885 3050 10890 3070
rect 10820 3020 10890 3050
rect 10820 3000 10825 3020
rect 10845 3000 10865 3020
rect 10885 3000 10890 3020
rect 10820 2990 10890 3000
rect 12910 3100 12915 3120
rect 12935 3100 12955 3120
rect 12975 3100 12980 3120
rect 12910 3070 12980 3100
rect 12910 3050 12915 3070
rect 12935 3050 12955 3070
rect 12975 3050 12980 3070
rect 12910 3020 12980 3050
rect 12910 3000 12915 3020
rect 12935 3000 12955 3020
rect 12975 3000 12980 3020
rect 12910 2990 12980 3000
rect 13005 3570 13035 3580
rect 13005 3550 13010 3570
rect 13030 3550 13035 3570
rect 13005 3520 13035 3550
rect 13005 3500 13010 3520
rect 13030 3500 13035 3520
rect 13005 3470 13035 3500
rect 13005 3450 13010 3470
rect 13030 3450 13035 3470
rect 13005 3420 13035 3450
rect 13005 3400 13010 3420
rect 13030 3400 13035 3420
rect 13005 3370 13035 3400
rect 13005 3350 13010 3370
rect 13030 3350 13035 3370
rect 13005 3320 13035 3350
rect 13005 3300 13010 3320
rect 13030 3300 13035 3320
rect 13005 3270 13035 3300
rect 13005 3250 13010 3270
rect 13030 3250 13035 3270
rect 13005 3220 13035 3250
rect 13005 3200 13010 3220
rect 13030 3200 13035 3220
rect 13005 3170 13035 3200
rect 13005 3150 13010 3170
rect 13030 3150 13035 3170
rect 13005 3120 13035 3150
rect 13005 3100 13010 3120
rect 13030 3100 13035 3120
rect 13005 3070 13035 3100
rect 13005 3050 13010 3070
rect 13030 3050 13035 3070
rect 13005 3020 13035 3050
rect 13005 3000 13010 3020
rect 13030 3000 13035 3020
rect 13005 2990 13035 3000
rect 13060 3570 13090 3580
rect 13060 3550 13065 3570
rect 13085 3550 13090 3570
rect 13060 3520 13090 3550
rect 13060 3500 13065 3520
rect 13085 3500 13090 3520
rect 13060 3470 13090 3500
rect 13060 3450 13065 3470
rect 13085 3450 13090 3470
rect 13060 3420 13090 3450
rect 13060 3400 13065 3420
rect 13085 3400 13090 3420
rect 13060 3370 13090 3400
rect 13060 3350 13065 3370
rect 13085 3350 13090 3370
rect 13060 3320 13090 3350
rect 13060 3300 13065 3320
rect 13085 3300 13090 3320
rect 13060 3270 13090 3300
rect 13060 3250 13065 3270
rect 13085 3250 13090 3270
rect 13060 3220 13090 3250
rect 13060 3200 13065 3220
rect 13085 3200 13090 3220
rect 13060 3170 13090 3200
rect 13060 3150 13065 3170
rect 13085 3150 13090 3170
rect 13060 3120 13090 3150
rect 13060 3100 13065 3120
rect 13085 3100 13090 3120
rect 13060 3070 13090 3100
rect 13060 3050 13065 3070
rect 13085 3050 13090 3070
rect 13060 3020 13090 3050
rect 13060 3000 13065 3020
rect 13085 3000 13090 3020
rect 13060 2990 13090 3000
rect 13115 3570 13145 3580
rect 13115 3550 13120 3570
rect 13140 3550 13145 3570
rect 13115 3520 13145 3550
rect 13115 3500 13120 3520
rect 13140 3500 13145 3520
rect 13115 3470 13145 3500
rect 13115 3450 13120 3470
rect 13140 3450 13145 3470
rect 13115 3420 13145 3450
rect 13115 3400 13120 3420
rect 13140 3400 13145 3420
rect 13115 3370 13145 3400
rect 13115 3350 13120 3370
rect 13140 3350 13145 3370
rect 13115 3320 13145 3350
rect 13115 3300 13120 3320
rect 13140 3300 13145 3320
rect 13115 3270 13145 3300
rect 13115 3250 13120 3270
rect 13140 3250 13145 3270
rect 13115 3220 13145 3250
rect 13115 3200 13120 3220
rect 13140 3200 13145 3220
rect 13115 3170 13145 3200
rect 13115 3150 13120 3170
rect 13140 3150 13145 3170
rect 13115 3120 13145 3150
rect 13115 3100 13120 3120
rect 13140 3100 13145 3120
rect 13115 3070 13145 3100
rect 13115 3050 13120 3070
rect 13140 3050 13145 3070
rect 13115 3020 13145 3050
rect 13115 3000 13120 3020
rect 13140 3000 13145 3020
rect 13115 2990 13145 3000
rect 13170 3570 13200 3580
rect 13170 3550 13175 3570
rect 13195 3550 13200 3570
rect 13170 3520 13200 3550
rect 13170 3500 13175 3520
rect 13195 3500 13200 3520
rect 13170 3470 13200 3500
rect 13170 3450 13175 3470
rect 13195 3450 13200 3470
rect 13170 3420 13200 3450
rect 13170 3400 13175 3420
rect 13195 3400 13200 3420
rect 13170 3370 13200 3400
rect 13170 3350 13175 3370
rect 13195 3350 13200 3370
rect 13170 3320 13200 3350
rect 13170 3300 13175 3320
rect 13195 3300 13200 3320
rect 13170 3270 13200 3300
rect 13170 3250 13175 3270
rect 13195 3250 13200 3270
rect 13170 3220 13200 3250
rect 13170 3200 13175 3220
rect 13195 3200 13200 3220
rect 13170 3170 13200 3200
rect 13170 3150 13175 3170
rect 13195 3150 13200 3170
rect 13170 3120 13200 3150
rect 13170 3100 13175 3120
rect 13195 3100 13200 3120
rect 13170 3070 13200 3100
rect 13170 3050 13175 3070
rect 13195 3050 13200 3070
rect 13170 3020 13200 3050
rect 13170 3000 13175 3020
rect 13195 3000 13200 3020
rect 13170 2990 13200 3000
rect 13225 3570 13255 3580
rect 13225 3550 13230 3570
rect 13250 3550 13255 3570
rect 13225 3520 13255 3550
rect 13225 3500 13230 3520
rect 13250 3500 13255 3520
rect 13225 3470 13255 3500
rect 13225 3450 13230 3470
rect 13250 3450 13255 3470
rect 13225 3420 13255 3450
rect 13225 3400 13230 3420
rect 13250 3400 13255 3420
rect 13225 3370 13255 3400
rect 13225 3350 13230 3370
rect 13250 3350 13255 3370
rect 13225 3320 13255 3350
rect 13225 3300 13230 3320
rect 13250 3300 13255 3320
rect 13225 3270 13255 3300
rect 13225 3250 13230 3270
rect 13250 3250 13255 3270
rect 13225 3220 13255 3250
rect 13225 3200 13230 3220
rect 13250 3200 13255 3220
rect 13225 3170 13255 3200
rect 13225 3150 13230 3170
rect 13250 3150 13255 3170
rect 13225 3120 13255 3150
rect 13225 3100 13230 3120
rect 13250 3100 13255 3120
rect 13225 3070 13255 3100
rect 13225 3050 13230 3070
rect 13250 3050 13255 3070
rect 13225 3020 13255 3050
rect 13225 3000 13230 3020
rect 13250 3000 13255 3020
rect 13225 2990 13255 3000
rect 13280 3570 13310 3580
rect 13280 3550 13285 3570
rect 13305 3550 13310 3570
rect 13280 3520 13310 3550
rect 13280 3500 13285 3520
rect 13305 3500 13310 3520
rect 13280 3470 13310 3500
rect 13280 3450 13285 3470
rect 13305 3450 13310 3470
rect 13280 3420 13310 3450
rect 13280 3400 13285 3420
rect 13305 3400 13310 3420
rect 13280 3370 13310 3400
rect 13280 3350 13285 3370
rect 13305 3350 13310 3370
rect 13280 3320 13310 3350
rect 13280 3300 13285 3320
rect 13305 3300 13310 3320
rect 13280 3270 13310 3300
rect 13280 3250 13285 3270
rect 13305 3250 13310 3270
rect 13280 3220 13310 3250
rect 13280 3200 13285 3220
rect 13305 3200 13310 3220
rect 13280 3170 13310 3200
rect 13280 3150 13285 3170
rect 13305 3150 13310 3170
rect 13280 3120 13310 3150
rect 13280 3100 13285 3120
rect 13305 3100 13310 3120
rect 13280 3070 13310 3100
rect 13280 3050 13285 3070
rect 13305 3050 13310 3070
rect 13280 3020 13310 3050
rect 13280 3000 13285 3020
rect 13305 3000 13310 3020
rect 13280 2990 13310 3000
rect 13335 3570 13365 3580
rect 13335 3550 13340 3570
rect 13360 3550 13365 3570
rect 13335 3520 13365 3550
rect 13335 3500 13340 3520
rect 13360 3500 13365 3520
rect 13335 3470 13365 3500
rect 13335 3450 13340 3470
rect 13360 3450 13365 3470
rect 13335 3420 13365 3450
rect 13335 3400 13340 3420
rect 13360 3400 13365 3420
rect 13335 3370 13365 3400
rect 13335 3350 13340 3370
rect 13360 3350 13365 3370
rect 13335 3320 13365 3350
rect 13335 3300 13340 3320
rect 13360 3300 13365 3320
rect 13335 3270 13365 3300
rect 13335 3250 13340 3270
rect 13360 3250 13365 3270
rect 13335 3220 13365 3250
rect 13335 3200 13340 3220
rect 13360 3200 13365 3220
rect 13335 3170 13365 3200
rect 13335 3150 13340 3170
rect 13360 3150 13365 3170
rect 13335 3120 13365 3150
rect 13335 3100 13340 3120
rect 13360 3100 13365 3120
rect 13335 3070 13365 3100
rect 13335 3050 13340 3070
rect 13360 3050 13365 3070
rect 13335 3020 13365 3050
rect 13335 3000 13340 3020
rect 13360 3000 13365 3020
rect 13335 2990 13365 3000
rect 13390 3570 13420 3580
rect 13390 3550 13395 3570
rect 13415 3550 13420 3570
rect 13390 3520 13420 3550
rect 13390 3500 13395 3520
rect 13415 3500 13420 3520
rect 13390 3470 13420 3500
rect 13390 3450 13395 3470
rect 13415 3450 13420 3470
rect 13390 3420 13420 3450
rect 13390 3400 13395 3420
rect 13415 3400 13420 3420
rect 13390 3370 13420 3400
rect 13390 3350 13395 3370
rect 13415 3350 13420 3370
rect 13390 3320 13420 3350
rect 13390 3300 13395 3320
rect 13415 3300 13420 3320
rect 13390 3270 13420 3300
rect 13390 3250 13395 3270
rect 13415 3250 13420 3270
rect 13390 3220 13420 3250
rect 13390 3200 13395 3220
rect 13415 3200 13420 3220
rect 13390 3170 13420 3200
rect 13390 3150 13395 3170
rect 13415 3150 13420 3170
rect 13390 3120 13420 3150
rect 13390 3100 13395 3120
rect 13415 3100 13420 3120
rect 13390 3070 13420 3100
rect 13390 3050 13395 3070
rect 13415 3050 13420 3070
rect 13390 3020 13420 3050
rect 13390 3000 13395 3020
rect 13415 3000 13420 3020
rect 13390 2990 13420 3000
rect 13445 3570 13475 3580
rect 13445 3550 13450 3570
rect 13470 3550 13475 3570
rect 13445 3520 13475 3550
rect 13445 3500 13450 3520
rect 13470 3500 13475 3520
rect 13445 3470 13475 3500
rect 13445 3450 13450 3470
rect 13470 3450 13475 3470
rect 13445 3420 13475 3450
rect 13445 3400 13450 3420
rect 13470 3400 13475 3420
rect 13445 3370 13475 3400
rect 13445 3350 13450 3370
rect 13470 3350 13475 3370
rect 13445 3320 13475 3350
rect 13445 3300 13450 3320
rect 13470 3300 13475 3320
rect 13445 3270 13475 3300
rect 13445 3250 13450 3270
rect 13470 3250 13475 3270
rect 13445 3220 13475 3250
rect 13445 3200 13450 3220
rect 13470 3200 13475 3220
rect 13445 3170 13475 3200
rect 13445 3150 13450 3170
rect 13470 3150 13475 3170
rect 13445 3120 13475 3150
rect 13445 3100 13450 3120
rect 13470 3100 13475 3120
rect 13445 3070 13475 3100
rect 13445 3050 13450 3070
rect 13470 3050 13475 3070
rect 13445 3020 13475 3050
rect 13445 3000 13450 3020
rect 13470 3000 13475 3020
rect 13445 2990 13475 3000
rect 13500 3570 13530 3580
rect 13500 3550 13505 3570
rect 13525 3550 13530 3570
rect 13500 3520 13530 3550
rect 13500 3500 13505 3520
rect 13525 3500 13530 3520
rect 13500 3470 13530 3500
rect 13500 3450 13505 3470
rect 13525 3450 13530 3470
rect 13500 3420 13530 3450
rect 13500 3400 13505 3420
rect 13525 3400 13530 3420
rect 13500 3370 13530 3400
rect 13500 3350 13505 3370
rect 13525 3350 13530 3370
rect 13500 3320 13530 3350
rect 13500 3300 13505 3320
rect 13525 3300 13530 3320
rect 13500 3270 13530 3300
rect 13500 3250 13505 3270
rect 13525 3250 13530 3270
rect 13500 3220 13530 3250
rect 13500 3200 13505 3220
rect 13525 3200 13530 3220
rect 13500 3170 13530 3200
rect 13500 3150 13505 3170
rect 13525 3150 13530 3170
rect 13500 3120 13530 3150
rect 13500 3100 13505 3120
rect 13525 3100 13530 3120
rect 13500 3070 13530 3100
rect 13500 3050 13505 3070
rect 13525 3050 13530 3070
rect 13500 3020 13530 3050
rect 13500 3000 13505 3020
rect 13525 3000 13530 3020
rect 13500 2990 13530 3000
rect 13555 3570 13585 3580
rect 13555 3550 13560 3570
rect 13580 3550 13585 3570
rect 13555 3520 13585 3550
rect 13555 3500 13560 3520
rect 13580 3500 13585 3520
rect 13555 3470 13585 3500
rect 13555 3450 13560 3470
rect 13580 3450 13585 3470
rect 13555 3420 13585 3450
rect 13555 3400 13560 3420
rect 13580 3400 13585 3420
rect 13555 3370 13585 3400
rect 13555 3350 13560 3370
rect 13580 3350 13585 3370
rect 13555 3320 13585 3350
rect 13555 3300 13560 3320
rect 13580 3300 13585 3320
rect 13555 3270 13585 3300
rect 13555 3250 13560 3270
rect 13580 3250 13585 3270
rect 13555 3220 13585 3250
rect 13555 3200 13560 3220
rect 13580 3200 13585 3220
rect 13555 3170 13585 3200
rect 13555 3150 13560 3170
rect 13580 3150 13585 3170
rect 13555 3120 13585 3150
rect 13555 3100 13560 3120
rect 13580 3100 13585 3120
rect 13555 3070 13585 3100
rect 13555 3050 13560 3070
rect 13580 3050 13585 3070
rect 13555 3020 13585 3050
rect 13555 3000 13560 3020
rect 13580 3000 13585 3020
rect 13555 2990 13585 3000
rect 13610 3570 13680 3580
rect 25905 3575 25945 3585
rect 26010 3575 26030 3595
rect 26180 3600 26190 3620
rect 26210 3600 26220 3620
rect 26180 3590 26220 3600
rect 26340 3620 26380 3630
rect 26340 3600 26350 3620
rect 26370 3600 26380 3620
rect 26340 3590 26380 3600
rect 26460 3620 26500 3630
rect 26460 3600 26470 3620
rect 26490 3600 26500 3620
rect 26460 3590 26500 3600
rect 26580 3620 26620 3630
rect 26580 3600 26590 3620
rect 26610 3600 26620 3620
rect 26580 3590 26620 3600
rect 26700 3620 26740 3630
rect 26700 3600 26710 3620
rect 26730 3600 26740 3620
rect 26700 3590 26740 3600
rect 26820 3620 26860 3630
rect 26820 3600 26830 3620
rect 26850 3600 26860 3620
rect 26820 3590 26860 3600
rect 26940 3620 26980 3630
rect 26940 3600 26950 3620
rect 26970 3600 26980 3620
rect 26940 3590 26980 3600
rect 27060 3620 27100 3630
rect 27060 3600 27070 3620
rect 27090 3600 27100 3620
rect 27060 3590 27100 3600
rect 27180 3620 27220 3630
rect 27180 3600 27190 3620
rect 27210 3600 27220 3620
rect 27180 3590 27220 3600
rect 27300 3620 27340 3630
rect 27300 3600 27310 3620
rect 27330 3600 27340 3620
rect 27300 3590 27340 3600
rect 27420 3620 27460 3630
rect 27420 3600 27430 3620
rect 27450 3600 27460 3620
rect 27420 3590 27460 3600
rect 27580 3620 27620 3630
rect 27580 3600 27590 3620
rect 27610 3600 27620 3620
rect 27580 3590 27620 3600
rect 13610 3550 13615 3570
rect 13635 3550 13655 3570
rect 13675 3550 13680 3570
rect 26005 3565 26035 3575
rect 13610 3520 13680 3550
rect 13610 3500 13615 3520
rect 13635 3500 13655 3520
rect 13675 3500 13680 3520
rect 13610 3470 13680 3500
rect 13610 3450 13615 3470
rect 13635 3450 13655 3470
rect 13675 3450 13680 3470
rect 13610 3420 13680 3450
rect 13610 3400 13615 3420
rect 13635 3400 13655 3420
rect 13675 3400 13680 3420
rect 13610 3370 13680 3400
rect 13610 3350 13615 3370
rect 13635 3350 13655 3370
rect 13675 3350 13680 3370
rect 13610 3320 13680 3350
rect 13610 3300 13615 3320
rect 13635 3300 13655 3320
rect 13675 3300 13680 3320
rect 13760 3520 13901 3560
rect 26005 3545 26010 3565
rect 26030 3545 26035 3565
rect 25785 3515 25855 3545
rect 25785 3495 25790 3515
rect 25810 3495 25830 3515
rect 25850 3495 25855 3515
rect 25785 3465 25855 3495
rect 25785 3445 25790 3465
rect 25810 3445 25830 3465
rect 25850 3445 25855 3465
rect 25785 3415 25855 3445
rect 25785 3395 25790 3415
rect 25810 3395 25830 3415
rect 25850 3395 25855 3415
rect 25785 3365 25855 3395
rect 25450 3340 25490 3350
rect 25450 3320 25460 3340
rect 25480 3320 25490 3340
rect 25450 3310 25490 3320
rect 25710 3340 25750 3350
rect 25710 3320 25720 3340
rect 25740 3320 25750 3340
rect 25710 3310 25750 3320
rect 25785 3345 25790 3365
rect 25810 3345 25830 3365
rect 25850 3345 25855 3365
rect 25785 3315 25855 3345
rect 13610 3270 13680 3300
rect 25460 3288 25480 3310
rect 25720 3288 25740 3310
rect 25785 3295 25790 3315
rect 25810 3295 25830 3315
rect 25850 3295 25855 3315
rect 13610 3250 13615 3270
rect 13635 3250 13655 3270
rect 13675 3250 13680 3270
rect 13610 3220 13680 3250
rect 25455 3265 25525 3288
rect 25455 3245 25460 3265
rect 25480 3245 25500 3265
rect 25520 3245 25525 3265
rect 25455 3235 25525 3245
rect 25555 3270 25585 3288
rect 25555 3250 25560 3270
rect 25580 3250 25585 3270
rect 25555 3235 25585 3250
rect 25615 3270 25645 3288
rect 25615 3250 25620 3270
rect 25640 3250 25645 3270
rect 25615 3235 25645 3250
rect 25675 3265 25745 3288
rect 25675 3245 25680 3265
rect 25700 3245 25720 3265
rect 25740 3245 25745 3265
rect 25675 3235 25745 3245
rect 25785 3265 25855 3295
rect 25785 3245 25790 3265
rect 25810 3245 25830 3265
rect 25850 3245 25855 3265
rect 25785 3235 25855 3245
rect 25885 3515 25915 3545
rect 25885 3495 25890 3515
rect 25910 3495 25915 3515
rect 25885 3465 25915 3495
rect 25885 3445 25890 3465
rect 25910 3445 25915 3465
rect 25885 3415 25915 3445
rect 25885 3395 25890 3415
rect 25910 3395 25915 3415
rect 25885 3365 25915 3395
rect 25885 3345 25890 3365
rect 25910 3345 25915 3365
rect 25885 3315 25915 3345
rect 25885 3295 25890 3315
rect 25910 3295 25915 3315
rect 25885 3265 25915 3295
rect 25885 3245 25890 3265
rect 25910 3245 25915 3265
rect 25885 3235 25915 3245
rect 25945 3515 25975 3545
rect 25945 3495 25950 3515
rect 25970 3495 25975 3515
rect 25945 3465 25975 3495
rect 25945 3445 25950 3465
rect 25970 3445 25975 3465
rect 25945 3415 25975 3445
rect 25945 3395 25950 3415
rect 25970 3395 25975 3415
rect 25945 3365 25975 3395
rect 25945 3345 25950 3365
rect 25970 3345 25975 3365
rect 25945 3315 25975 3345
rect 25945 3295 25950 3315
rect 25970 3295 25975 3315
rect 25945 3265 25975 3295
rect 25945 3245 25950 3265
rect 25970 3245 25975 3265
rect 25945 3235 25975 3245
rect 26005 3515 26035 3545
rect 26005 3495 26010 3515
rect 26030 3495 26035 3515
rect 26005 3465 26035 3495
rect 26005 3445 26010 3465
rect 26030 3445 26035 3465
rect 26005 3415 26035 3445
rect 26005 3395 26010 3415
rect 26030 3395 26035 3415
rect 26005 3365 26035 3395
rect 26005 3345 26010 3365
rect 26030 3345 26035 3365
rect 26005 3315 26035 3345
rect 26005 3295 26010 3315
rect 26030 3295 26035 3315
rect 26005 3265 26035 3295
rect 26005 3245 26010 3265
rect 26030 3245 26035 3265
rect 26005 3235 26035 3245
rect 26065 3565 26135 3575
rect 26190 3570 26210 3590
rect 26350 3570 26370 3590
rect 26470 3570 26490 3590
rect 26590 3570 26610 3590
rect 26710 3570 26730 3590
rect 26830 3570 26850 3590
rect 26950 3570 26970 3590
rect 27070 3570 27090 3590
rect 27190 3570 27210 3590
rect 27310 3570 27330 3590
rect 27430 3570 27450 3590
rect 27590 3570 27610 3590
rect 26065 3545 26070 3565
rect 26090 3545 26110 3565
rect 26130 3545 26135 3565
rect 26065 3515 26135 3545
rect 26065 3495 26070 3515
rect 26090 3495 26110 3515
rect 26130 3495 26135 3515
rect 26065 3465 26135 3495
rect 26065 3445 26070 3465
rect 26090 3445 26110 3465
rect 26130 3445 26135 3465
rect 26065 3415 26135 3445
rect 26065 3395 26070 3415
rect 26090 3395 26110 3415
rect 26130 3395 26135 3415
rect 26065 3365 26135 3395
rect 26065 3345 26070 3365
rect 26090 3345 26110 3365
rect 26130 3345 26135 3365
rect 26065 3315 26135 3345
rect 26065 3295 26070 3315
rect 26090 3295 26110 3315
rect 26130 3295 26135 3315
rect 26065 3265 26135 3295
rect 26065 3245 26070 3265
rect 26090 3245 26110 3265
rect 26130 3245 26135 3265
rect 26065 3235 26135 3245
rect 26185 3560 26255 3570
rect 26185 3540 26190 3560
rect 26210 3540 26230 3560
rect 26250 3540 26255 3560
rect 26185 3510 26255 3540
rect 26185 3490 26190 3510
rect 26210 3490 26230 3510
rect 26250 3490 26255 3510
rect 26185 3460 26255 3490
rect 26185 3440 26190 3460
rect 26210 3440 26230 3460
rect 26250 3440 26255 3460
rect 26185 3410 26255 3440
rect 26185 3390 26190 3410
rect 26210 3390 26230 3410
rect 26250 3390 26255 3410
rect 26185 3360 26255 3390
rect 26185 3340 26190 3360
rect 26210 3340 26230 3360
rect 26250 3340 26255 3360
rect 26185 3310 26255 3340
rect 26185 3290 26190 3310
rect 26210 3290 26230 3310
rect 26250 3290 26255 3310
rect 26185 3260 26255 3290
rect 26185 3240 26190 3260
rect 26210 3240 26230 3260
rect 26250 3240 26255 3260
rect 13610 3200 13615 3220
rect 13635 3200 13655 3220
rect 13675 3200 13680 3220
rect 25620 3215 25640 3235
rect 25790 3215 25810 3235
rect 26110 3215 26130 3235
rect 13610 3170 13680 3200
rect 25580 3205 25640 3215
rect 25580 3185 25590 3205
rect 25610 3195 25640 3205
rect 25780 3205 25820 3215
rect 25610 3185 25620 3195
rect 25580 3175 25620 3185
rect 25780 3185 25790 3205
rect 25810 3185 25820 3205
rect 25780 3175 25820 3185
rect 25905 3205 25940 3215
rect 25905 3185 25910 3205
rect 25930 3185 25940 3205
rect 25905 3175 25940 3185
rect 25980 3205 26015 3215
rect 25980 3185 25990 3205
rect 26010 3185 26015 3205
rect 25980 3175 26015 3185
rect 26100 3205 26140 3215
rect 26100 3185 26110 3205
rect 26130 3185 26140 3205
rect 26100 3175 26140 3185
rect 26185 3210 26255 3240
rect 26185 3190 26190 3210
rect 26210 3190 26230 3210
rect 26250 3190 26255 3210
rect 26185 3180 26255 3190
rect 26285 3560 26315 3570
rect 26285 3540 26290 3560
rect 26310 3540 26315 3560
rect 26285 3510 26315 3540
rect 26285 3490 26290 3510
rect 26310 3490 26315 3510
rect 26285 3460 26315 3490
rect 26285 3440 26290 3460
rect 26310 3440 26315 3460
rect 26285 3410 26315 3440
rect 26285 3390 26290 3410
rect 26310 3390 26315 3410
rect 26285 3360 26315 3390
rect 26285 3340 26290 3360
rect 26310 3340 26315 3360
rect 26285 3310 26315 3340
rect 26285 3290 26290 3310
rect 26310 3290 26315 3310
rect 26285 3260 26315 3290
rect 26285 3240 26290 3260
rect 26310 3240 26315 3260
rect 26285 3210 26315 3240
rect 26285 3190 26290 3210
rect 26310 3190 26315 3210
rect 26285 3180 26315 3190
rect 26345 3560 26375 3570
rect 26345 3540 26350 3560
rect 26370 3540 26375 3560
rect 26345 3510 26375 3540
rect 26345 3490 26350 3510
rect 26370 3490 26375 3510
rect 26345 3460 26375 3490
rect 26345 3440 26350 3460
rect 26370 3440 26375 3460
rect 26345 3410 26375 3440
rect 26345 3390 26350 3410
rect 26370 3390 26375 3410
rect 26345 3360 26375 3390
rect 26345 3340 26350 3360
rect 26370 3340 26375 3360
rect 26345 3310 26375 3340
rect 26345 3290 26350 3310
rect 26370 3290 26375 3310
rect 26345 3260 26375 3290
rect 26345 3240 26350 3260
rect 26370 3240 26375 3260
rect 26345 3210 26375 3240
rect 26345 3190 26350 3210
rect 26370 3190 26375 3210
rect 26345 3180 26375 3190
rect 26405 3560 26435 3570
rect 26405 3540 26410 3560
rect 26430 3540 26435 3560
rect 26405 3510 26435 3540
rect 26405 3490 26410 3510
rect 26430 3490 26435 3510
rect 26405 3460 26435 3490
rect 26405 3440 26410 3460
rect 26430 3440 26435 3460
rect 26405 3410 26435 3440
rect 26405 3390 26410 3410
rect 26430 3390 26435 3410
rect 26405 3360 26435 3390
rect 26405 3340 26410 3360
rect 26430 3340 26435 3360
rect 26405 3310 26435 3340
rect 26405 3290 26410 3310
rect 26430 3290 26435 3310
rect 26405 3260 26435 3290
rect 26405 3240 26410 3260
rect 26430 3240 26435 3260
rect 26405 3210 26435 3240
rect 26405 3190 26410 3210
rect 26430 3190 26435 3210
rect 26405 3180 26435 3190
rect 26465 3560 26495 3570
rect 26465 3540 26470 3560
rect 26490 3540 26495 3560
rect 26465 3510 26495 3540
rect 26465 3490 26470 3510
rect 26490 3490 26495 3510
rect 26465 3460 26495 3490
rect 26465 3440 26470 3460
rect 26490 3440 26495 3460
rect 26465 3410 26495 3440
rect 26465 3390 26470 3410
rect 26490 3390 26495 3410
rect 26465 3360 26495 3390
rect 26465 3340 26470 3360
rect 26490 3340 26495 3360
rect 26465 3310 26495 3340
rect 26465 3290 26470 3310
rect 26490 3290 26495 3310
rect 26465 3260 26495 3290
rect 26465 3240 26470 3260
rect 26490 3240 26495 3260
rect 26465 3210 26495 3240
rect 26465 3190 26470 3210
rect 26490 3190 26495 3210
rect 26465 3180 26495 3190
rect 26525 3560 26555 3570
rect 26525 3540 26530 3560
rect 26550 3540 26555 3560
rect 26525 3510 26555 3540
rect 26525 3490 26530 3510
rect 26550 3490 26555 3510
rect 26525 3460 26555 3490
rect 26525 3440 26530 3460
rect 26550 3440 26555 3460
rect 26525 3410 26555 3440
rect 26525 3390 26530 3410
rect 26550 3390 26555 3410
rect 26525 3360 26555 3390
rect 26525 3340 26530 3360
rect 26550 3340 26555 3360
rect 26525 3310 26555 3340
rect 26525 3290 26530 3310
rect 26550 3290 26555 3310
rect 26525 3260 26555 3290
rect 26525 3240 26530 3260
rect 26550 3240 26555 3260
rect 26525 3210 26555 3240
rect 26525 3190 26530 3210
rect 26550 3190 26555 3210
rect 26525 3180 26555 3190
rect 26585 3560 26615 3570
rect 26585 3540 26590 3560
rect 26610 3540 26615 3560
rect 26585 3510 26615 3540
rect 26585 3490 26590 3510
rect 26610 3490 26615 3510
rect 26585 3460 26615 3490
rect 26585 3440 26590 3460
rect 26610 3440 26615 3460
rect 26585 3410 26615 3440
rect 26585 3390 26590 3410
rect 26610 3390 26615 3410
rect 26585 3360 26615 3390
rect 26585 3340 26590 3360
rect 26610 3340 26615 3360
rect 26585 3310 26615 3340
rect 26585 3290 26590 3310
rect 26610 3290 26615 3310
rect 26585 3260 26615 3290
rect 26585 3240 26590 3260
rect 26610 3240 26615 3260
rect 26585 3210 26615 3240
rect 26585 3190 26590 3210
rect 26610 3190 26615 3210
rect 26585 3180 26615 3190
rect 26645 3560 26675 3570
rect 26645 3540 26650 3560
rect 26670 3540 26675 3560
rect 26645 3510 26675 3540
rect 26645 3490 26650 3510
rect 26670 3490 26675 3510
rect 26645 3460 26675 3490
rect 26645 3440 26650 3460
rect 26670 3440 26675 3460
rect 26645 3410 26675 3440
rect 26645 3390 26650 3410
rect 26670 3390 26675 3410
rect 26645 3360 26675 3390
rect 26645 3340 26650 3360
rect 26670 3340 26675 3360
rect 26645 3310 26675 3340
rect 26645 3290 26650 3310
rect 26670 3290 26675 3310
rect 26645 3260 26675 3290
rect 26645 3240 26650 3260
rect 26670 3240 26675 3260
rect 26645 3210 26675 3240
rect 26645 3190 26650 3210
rect 26670 3190 26675 3210
rect 26645 3180 26675 3190
rect 26705 3560 26735 3570
rect 26705 3540 26710 3560
rect 26730 3540 26735 3560
rect 26705 3510 26735 3540
rect 26705 3490 26710 3510
rect 26730 3490 26735 3510
rect 26705 3460 26735 3490
rect 26705 3440 26710 3460
rect 26730 3440 26735 3460
rect 26705 3410 26735 3440
rect 26705 3390 26710 3410
rect 26730 3390 26735 3410
rect 26705 3360 26735 3390
rect 26705 3340 26710 3360
rect 26730 3340 26735 3360
rect 26705 3310 26735 3340
rect 26705 3290 26710 3310
rect 26730 3290 26735 3310
rect 26705 3260 26735 3290
rect 26705 3240 26710 3260
rect 26730 3240 26735 3260
rect 26705 3210 26735 3240
rect 26705 3190 26710 3210
rect 26730 3190 26735 3210
rect 26705 3180 26735 3190
rect 26765 3560 26795 3570
rect 26765 3540 26770 3560
rect 26790 3540 26795 3560
rect 26765 3510 26795 3540
rect 26765 3490 26770 3510
rect 26790 3490 26795 3510
rect 26765 3460 26795 3490
rect 26765 3440 26770 3460
rect 26790 3440 26795 3460
rect 26765 3410 26795 3440
rect 26765 3390 26770 3410
rect 26790 3390 26795 3410
rect 26765 3360 26795 3390
rect 26765 3340 26770 3360
rect 26790 3340 26795 3360
rect 26765 3310 26795 3340
rect 26765 3290 26770 3310
rect 26790 3290 26795 3310
rect 26765 3260 26795 3290
rect 26765 3240 26770 3260
rect 26790 3240 26795 3260
rect 26765 3210 26795 3240
rect 26765 3190 26770 3210
rect 26790 3190 26795 3210
rect 26765 3180 26795 3190
rect 26825 3560 26855 3570
rect 26825 3540 26830 3560
rect 26850 3540 26855 3560
rect 26825 3510 26855 3540
rect 26825 3490 26830 3510
rect 26850 3490 26855 3510
rect 26825 3460 26855 3490
rect 26825 3440 26830 3460
rect 26850 3440 26855 3460
rect 26825 3410 26855 3440
rect 26825 3390 26830 3410
rect 26850 3390 26855 3410
rect 26825 3360 26855 3390
rect 26825 3340 26830 3360
rect 26850 3340 26855 3360
rect 26825 3310 26855 3340
rect 26825 3290 26830 3310
rect 26850 3290 26855 3310
rect 26825 3260 26855 3290
rect 26825 3240 26830 3260
rect 26850 3240 26855 3260
rect 26825 3210 26855 3240
rect 26825 3190 26830 3210
rect 26850 3190 26855 3210
rect 26825 3180 26855 3190
rect 26885 3560 26915 3570
rect 26885 3540 26890 3560
rect 26910 3540 26915 3560
rect 26885 3510 26915 3540
rect 26885 3490 26890 3510
rect 26910 3490 26915 3510
rect 26885 3460 26915 3490
rect 26885 3440 26890 3460
rect 26910 3440 26915 3460
rect 26885 3410 26915 3440
rect 26885 3390 26890 3410
rect 26910 3390 26915 3410
rect 26885 3360 26915 3390
rect 26885 3340 26890 3360
rect 26910 3340 26915 3360
rect 26885 3310 26915 3340
rect 26885 3290 26890 3310
rect 26910 3290 26915 3310
rect 26885 3260 26915 3290
rect 26885 3240 26890 3260
rect 26910 3240 26915 3260
rect 26885 3210 26915 3240
rect 26885 3190 26890 3210
rect 26910 3190 26915 3210
rect 26885 3180 26915 3190
rect 26945 3560 26975 3570
rect 26945 3540 26950 3560
rect 26970 3540 26975 3560
rect 26945 3510 26975 3540
rect 26945 3490 26950 3510
rect 26970 3490 26975 3510
rect 26945 3460 26975 3490
rect 26945 3440 26950 3460
rect 26970 3440 26975 3460
rect 26945 3410 26975 3440
rect 26945 3390 26950 3410
rect 26970 3390 26975 3410
rect 26945 3360 26975 3390
rect 26945 3340 26950 3360
rect 26970 3340 26975 3360
rect 26945 3310 26975 3340
rect 26945 3290 26950 3310
rect 26970 3290 26975 3310
rect 26945 3260 26975 3290
rect 26945 3240 26950 3260
rect 26970 3240 26975 3260
rect 26945 3210 26975 3240
rect 26945 3190 26950 3210
rect 26970 3190 26975 3210
rect 26945 3180 26975 3190
rect 27005 3560 27035 3570
rect 27005 3540 27010 3560
rect 27030 3540 27035 3560
rect 27005 3510 27035 3540
rect 27005 3490 27010 3510
rect 27030 3490 27035 3510
rect 27005 3460 27035 3490
rect 27005 3440 27010 3460
rect 27030 3440 27035 3460
rect 27005 3410 27035 3440
rect 27005 3390 27010 3410
rect 27030 3390 27035 3410
rect 27005 3360 27035 3390
rect 27005 3340 27010 3360
rect 27030 3340 27035 3360
rect 27005 3310 27035 3340
rect 27005 3290 27010 3310
rect 27030 3290 27035 3310
rect 27005 3260 27035 3290
rect 27005 3240 27010 3260
rect 27030 3240 27035 3260
rect 27005 3210 27035 3240
rect 27005 3190 27010 3210
rect 27030 3190 27035 3210
rect 27005 3180 27035 3190
rect 27065 3560 27095 3570
rect 27065 3540 27070 3560
rect 27090 3540 27095 3560
rect 27065 3510 27095 3540
rect 27065 3490 27070 3510
rect 27090 3490 27095 3510
rect 27065 3460 27095 3490
rect 27065 3440 27070 3460
rect 27090 3440 27095 3460
rect 27065 3410 27095 3440
rect 27065 3390 27070 3410
rect 27090 3390 27095 3410
rect 27065 3360 27095 3390
rect 27065 3340 27070 3360
rect 27090 3340 27095 3360
rect 27065 3310 27095 3340
rect 27065 3290 27070 3310
rect 27090 3290 27095 3310
rect 27065 3260 27095 3290
rect 27065 3240 27070 3260
rect 27090 3240 27095 3260
rect 27065 3210 27095 3240
rect 27065 3190 27070 3210
rect 27090 3190 27095 3210
rect 27065 3180 27095 3190
rect 27125 3560 27155 3570
rect 27125 3540 27130 3560
rect 27150 3540 27155 3560
rect 27125 3510 27155 3540
rect 27125 3490 27130 3510
rect 27150 3490 27155 3510
rect 27125 3460 27155 3490
rect 27125 3440 27130 3460
rect 27150 3440 27155 3460
rect 27125 3410 27155 3440
rect 27125 3390 27130 3410
rect 27150 3390 27155 3410
rect 27125 3360 27155 3390
rect 27125 3340 27130 3360
rect 27150 3340 27155 3360
rect 27125 3310 27155 3340
rect 27125 3290 27130 3310
rect 27150 3290 27155 3310
rect 27125 3260 27155 3290
rect 27125 3240 27130 3260
rect 27150 3240 27155 3260
rect 27125 3210 27155 3240
rect 27125 3190 27130 3210
rect 27150 3190 27155 3210
rect 27125 3180 27155 3190
rect 27185 3560 27215 3570
rect 27185 3540 27190 3560
rect 27210 3540 27215 3560
rect 27185 3510 27215 3540
rect 27185 3490 27190 3510
rect 27210 3490 27215 3510
rect 27185 3460 27215 3490
rect 27185 3440 27190 3460
rect 27210 3440 27215 3460
rect 27185 3410 27215 3440
rect 27185 3390 27190 3410
rect 27210 3390 27215 3410
rect 27185 3360 27215 3390
rect 27185 3340 27190 3360
rect 27210 3340 27215 3360
rect 27185 3310 27215 3340
rect 27185 3290 27190 3310
rect 27210 3290 27215 3310
rect 27185 3260 27215 3290
rect 27185 3240 27190 3260
rect 27210 3240 27215 3260
rect 27185 3210 27215 3240
rect 27185 3190 27190 3210
rect 27210 3190 27215 3210
rect 27185 3180 27215 3190
rect 27245 3560 27275 3570
rect 27245 3540 27250 3560
rect 27270 3540 27275 3560
rect 27245 3510 27275 3540
rect 27245 3490 27250 3510
rect 27270 3490 27275 3510
rect 27245 3460 27275 3490
rect 27245 3440 27250 3460
rect 27270 3440 27275 3460
rect 27245 3410 27275 3440
rect 27245 3390 27250 3410
rect 27270 3390 27275 3410
rect 27245 3360 27275 3390
rect 27245 3340 27250 3360
rect 27270 3340 27275 3360
rect 27245 3310 27275 3340
rect 27245 3290 27250 3310
rect 27270 3290 27275 3310
rect 27245 3260 27275 3290
rect 27245 3240 27250 3260
rect 27270 3240 27275 3260
rect 27245 3210 27275 3240
rect 27245 3190 27250 3210
rect 27270 3190 27275 3210
rect 27245 3180 27275 3190
rect 27305 3560 27335 3570
rect 27305 3540 27310 3560
rect 27330 3540 27335 3560
rect 27305 3510 27335 3540
rect 27305 3490 27310 3510
rect 27330 3490 27335 3510
rect 27305 3460 27335 3490
rect 27305 3440 27310 3460
rect 27330 3440 27335 3460
rect 27305 3410 27335 3440
rect 27305 3390 27310 3410
rect 27330 3390 27335 3410
rect 27305 3360 27335 3390
rect 27305 3340 27310 3360
rect 27330 3340 27335 3360
rect 27305 3310 27335 3340
rect 27305 3290 27310 3310
rect 27330 3290 27335 3310
rect 27305 3260 27335 3290
rect 27305 3240 27310 3260
rect 27330 3240 27335 3260
rect 27305 3210 27335 3240
rect 27305 3190 27310 3210
rect 27330 3190 27335 3210
rect 27305 3180 27335 3190
rect 27365 3560 27395 3570
rect 27365 3540 27370 3560
rect 27390 3540 27395 3560
rect 27365 3510 27395 3540
rect 27365 3490 27370 3510
rect 27390 3490 27395 3510
rect 27365 3460 27395 3490
rect 27365 3440 27370 3460
rect 27390 3440 27395 3460
rect 27365 3410 27395 3440
rect 27365 3390 27370 3410
rect 27390 3390 27395 3410
rect 27365 3360 27395 3390
rect 27365 3340 27370 3360
rect 27390 3340 27395 3360
rect 27365 3310 27395 3340
rect 27365 3290 27370 3310
rect 27390 3290 27395 3310
rect 27365 3260 27395 3290
rect 27365 3240 27370 3260
rect 27390 3240 27395 3260
rect 27365 3210 27395 3240
rect 27365 3190 27370 3210
rect 27390 3190 27395 3210
rect 27365 3180 27395 3190
rect 27425 3560 27455 3570
rect 27425 3540 27430 3560
rect 27450 3540 27455 3560
rect 27425 3510 27455 3540
rect 27425 3490 27430 3510
rect 27450 3490 27455 3510
rect 27425 3460 27455 3490
rect 27425 3440 27430 3460
rect 27450 3440 27455 3460
rect 27425 3410 27455 3440
rect 27425 3390 27430 3410
rect 27450 3390 27455 3410
rect 27425 3360 27455 3390
rect 27425 3340 27430 3360
rect 27450 3340 27455 3360
rect 27425 3310 27455 3340
rect 27425 3290 27430 3310
rect 27450 3290 27455 3310
rect 27425 3260 27455 3290
rect 27425 3240 27430 3260
rect 27450 3240 27455 3260
rect 27425 3210 27455 3240
rect 27425 3190 27430 3210
rect 27450 3190 27455 3210
rect 27425 3180 27455 3190
rect 27485 3560 27515 3570
rect 27485 3540 27490 3560
rect 27510 3540 27515 3560
rect 27485 3510 27515 3540
rect 27485 3490 27490 3510
rect 27510 3490 27515 3510
rect 27485 3460 27515 3490
rect 27485 3440 27490 3460
rect 27510 3440 27515 3460
rect 27485 3410 27515 3440
rect 27485 3390 27490 3410
rect 27510 3390 27515 3410
rect 27485 3360 27515 3390
rect 27485 3340 27490 3360
rect 27510 3340 27515 3360
rect 27485 3310 27515 3340
rect 27485 3290 27490 3310
rect 27510 3290 27515 3310
rect 27485 3260 27515 3290
rect 27485 3240 27490 3260
rect 27510 3240 27515 3260
rect 27485 3210 27515 3240
rect 27485 3190 27490 3210
rect 27510 3190 27515 3210
rect 27485 3180 27515 3190
rect 27545 3560 27615 3570
rect 27545 3540 27550 3560
rect 27570 3540 27590 3560
rect 27610 3540 27615 3560
rect 27545 3510 27615 3540
rect 27545 3490 27550 3510
rect 27570 3490 27590 3510
rect 27610 3490 27615 3510
rect 27545 3460 27615 3490
rect 27545 3440 27550 3460
rect 27570 3440 27590 3460
rect 27610 3440 27615 3460
rect 27545 3410 27615 3440
rect 27545 3390 27550 3410
rect 27570 3390 27590 3410
rect 27610 3390 27615 3410
rect 27545 3360 27615 3390
rect 27545 3340 27550 3360
rect 27570 3340 27590 3360
rect 27610 3340 27615 3360
rect 27545 3310 27615 3340
rect 27545 3290 27550 3310
rect 27570 3290 27590 3310
rect 27610 3290 27615 3310
rect 27545 3260 27615 3290
rect 27545 3240 27550 3260
rect 27570 3240 27590 3260
rect 27610 3240 27615 3260
rect 27945 3285 27985 3295
rect 27945 3265 27955 3285
rect 27975 3265 27985 3285
rect 27945 3255 27985 3265
rect 28055 3285 28095 3295
rect 28055 3265 28065 3285
rect 28085 3265 28095 3285
rect 28055 3255 28095 3265
rect 28165 3285 28205 3295
rect 28165 3265 28175 3285
rect 28195 3265 28205 3285
rect 28165 3255 28205 3265
rect 28275 3285 28315 3295
rect 28275 3265 28285 3285
rect 28305 3265 28315 3285
rect 28275 3255 28315 3265
rect 28385 3285 28425 3295
rect 28385 3265 28395 3285
rect 28415 3265 28425 3285
rect 28385 3255 28425 3265
rect 28495 3285 28535 3295
rect 28495 3265 28505 3285
rect 28525 3265 28535 3285
rect 28495 3255 28535 3265
rect 28605 3285 28645 3295
rect 28605 3265 28615 3285
rect 28635 3265 28645 3285
rect 28605 3255 28645 3265
rect 28715 3285 28755 3295
rect 28715 3265 28725 3285
rect 28745 3265 28755 3285
rect 28715 3255 28755 3265
rect 28825 3285 28865 3295
rect 28825 3265 28835 3285
rect 28855 3265 28865 3285
rect 28825 3255 28865 3265
rect 28935 3285 28975 3295
rect 28935 3265 28945 3285
rect 28965 3265 28975 3285
rect 28935 3255 28975 3265
rect 29045 3285 29085 3295
rect 29045 3265 29055 3285
rect 29075 3265 29085 3285
rect 29045 3255 29085 3265
rect 27545 3210 27615 3240
rect 27955 3235 27975 3255
rect 28065 3235 28085 3255
rect 28175 3235 28195 3255
rect 28285 3235 28305 3255
rect 28395 3235 28415 3255
rect 28505 3235 28525 3255
rect 28615 3235 28635 3255
rect 28725 3235 28745 3255
rect 28835 3235 28855 3255
rect 28945 3235 28965 3255
rect 29055 3235 29075 3255
rect 27545 3190 27550 3210
rect 27570 3190 27590 3210
rect 27610 3190 27615 3210
rect 27545 3180 27615 3190
rect 27855 3225 27925 3235
rect 27855 3205 27860 3225
rect 27880 3205 27900 3225
rect 27920 3205 27925 3225
rect 13610 3150 13615 3170
rect 13635 3150 13655 3170
rect 13675 3150 13680 3170
rect 26290 3160 26310 3180
rect 26410 3160 26430 3180
rect 26530 3160 26550 3180
rect 26650 3160 26670 3180
rect 26770 3160 26790 3180
rect 26890 3160 26910 3180
rect 27010 3160 27030 3180
rect 27130 3160 27150 3180
rect 27250 3160 27270 3180
rect 27370 3160 27390 3180
rect 27490 3160 27510 3180
rect 27855 3175 27925 3205
rect 13610 3120 13680 3150
rect 13610 3100 13615 3120
rect 13635 3100 13655 3120
rect 13675 3100 13680 3120
rect 13610 3070 13680 3100
rect 13610 3050 13615 3070
rect 13635 3050 13655 3070
rect 13675 3050 13680 3070
rect 13610 3020 13680 3050
rect 13610 3000 13615 3020
rect 13635 3000 13655 3020
rect 13675 3000 13680 3020
rect 13610 2990 13680 3000
rect 10125 2970 10145 2990
rect 10275 2970 10295 2990
rect 10385 2970 10405 2990
rect 10495 2970 10515 2990
rect 10605 2970 10625 2990
rect 10715 2970 10735 2990
rect 10865 2970 10885 2990
rect 12915 2970 12935 2990
rect 13065 2970 13085 2990
rect 13175 2970 13195 2990
rect 13285 2970 13305 2990
rect 13395 2970 13415 2990
rect 13505 2970 13525 2990
rect 13655 2970 13675 2990
rect 2960 2915 3030 2925
rect 1266 2865 1306 2900
rect 2330 2895 2375 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect 2960 2895 2965 2915
rect 2985 2895 3005 2915
rect 3025 2895 3030 2915
rect 2960 2865 3030 2895
rect -55 2825 -25 2855
rect 51 2850 96 2855
rect 51 2825 61 2850
rect 86 2825 96 2850
rect 51 2820 96 2825
rect 724 2850 769 2855
rect 724 2825 734 2850
rect 759 2825 769 2850
rect 724 2820 769 2825
rect 1210 2820 1240 2850
rect 2960 2845 2965 2865
rect 2985 2845 3005 2865
rect 3025 2845 3030 2865
rect 1261 2835 1306 2840
rect 1261 2810 1271 2835
rect 1296 2810 1306 2835
rect 1261 2805 1306 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2960 2835 3030 2845
rect 3090 2915 3120 2925
rect 3090 2895 3095 2915
rect 3115 2895 3120 2915
rect 3090 2865 3120 2895
rect 3090 2845 3095 2865
rect 3115 2845 3120 2865
rect 3090 2835 3120 2845
rect 3180 2915 3210 2925
rect 3180 2895 3185 2915
rect 3205 2895 3210 2915
rect 3180 2865 3210 2895
rect 3180 2845 3185 2865
rect 3205 2845 3210 2865
rect 3180 2835 3210 2845
rect 3270 2915 3300 2925
rect 3270 2895 3275 2915
rect 3295 2895 3300 2915
rect 3270 2865 3300 2895
rect 3270 2845 3275 2865
rect 3295 2845 3300 2865
rect 3270 2835 3300 2845
rect 3360 2915 3390 2925
rect 3360 2895 3365 2915
rect 3385 2895 3390 2915
rect 3360 2865 3390 2895
rect 3360 2845 3365 2865
rect 3385 2845 3390 2865
rect 3360 2835 3390 2845
rect 3450 2915 3480 2925
rect 3450 2895 3455 2915
rect 3475 2895 3480 2915
rect 3450 2865 3480 2895
rect 3450 2845 3455 2865
rect 3475 2845 3480 2865
rect 3450 2835 3480 2845
rect 3540 2915 3570 2925
rect 3540 2895 3545 2915
rect 3565 2895 3570 2915
rect 3540 2865 3570 2895
rect 3540 2845 3545 2865
rect 3565 2845 3570 2865
rect 3540 2835 3570 2845
rect 3630 2915 3660 2925
rect 3630 2895 3635 2915
rect 3655 2895 3660 2915
rect 3630 2865 3660 2895
rect 3630 2845 3635 2865
rect 3655 2845 3660 2865
rect 3630 2835 3660 2845
rect 3720 2915 3750 2925
rect 3720 2895 3725 2915
rect 3745 2895 3750 2915
rect 3720 2865 3750 2895
rect 3720 2845 3725 2865
rect 3745 2845 3750 2865
rect 3720 2835 3750 2845
rect 3810 2915 3840 2925
rect 3810 2895 3815 2915
rect 3835 2895 3840 2915
rect 3810 2865 3840 2895
rect 3810 2845 3815 2865
rect 3835 2845 3840 2865
rect 3810 2835 3840 2845
rect 3900 2915 3930 2925
rect 3900 2895 3905 2915
rect 3925 2895 3930 2915
rect 3900 2865 3930 2895
rect 3900 2845 3905 2865
rect 3925 2845 3930 2865
rect 3900 2835 3930 2845
rect 3990 2915 4020 2925
rect 3990 2895 3995 2915
rect 4015 2895 4020 2915
rect 3990 2865 4020 2895
rect 3990 2845 3995 2865
rect 4015 2845 4020 2865
rect 3990 2835 4020 2845
rect 4080 2915 4110 2925
rect 4080 2895 4085 2915
rect 4105 2895 4110 2915
rect 4080 2865 4110 2895
rect 4080 2845 4085 2865
rect 4105 2845 4110 2865
rect 4080 2835 4110 2845
rect 4170 2915 4200 2925
rect 4170 2895 4175 2915
rect 4195 2895 4200 2915
rect 4170 2865 4200 2895
rect 4170 2845 4175 2865
rect 4195 2845 4200 2865
rect 4170 2835 4200 2845
rect 4260 2915 4290 2925
rect 4260 2895 4265 2915
rect 4285 2895 4290 2915
rect 4260 2865 4290 2895
rect 4260 2845 4265 2865
rect 4285 2845 4290 2865
rect 4260 2835 4290 2845
rect 4350 2915 4380 2925
rect 4350 2895 4355 2915
rect 4375 2895 4380 2915
rect 4350 2865 4380 2895
rect 4350 2845 4355 2865
rect 4375 2845 4380 2865
rect 4350 2835 4380 2845
rect 4440 2915 4470 2925
rect 4440 2895 4445 2915
rect 4465 2895 4470 2915
rect 4440 2865 4470 2895
rect 4440 2845 4445 2865
rect 4465 2845 4470 2865
rect 4440 2835 4470 2845
rect 4530 2915 4560 2925
rect 4530 2895 4535 2915
rect 4555 2895 4560 2915
rect 4530 2865 4560 2895
rect 4530 2845 4535 2865
rect 4555 2845 4560 2865
rect 4530 2835 4560 2845
rect 4620 2915 4650 2925
rect 4620 2895 4625 2915
rect 4645 2895 4650 2915
rect 4620 2865 4650 2895
rect 4620 2845 4625 2865
rect 4645 2845 4650 2865
rect 4620 2835 4650 2845
rect 4710 2915 4740 2925
rect 4710 2895 4715 2915
rect 4735 2895 4740 2915
rect 4710 2865 4740 2895
rect 4710 2845 4715 2865
rect 4735 2845 4740 2865
rect 4710 2835 4740 2845
rect 4800 2915 4830 2925
rect 4800 2895 4805 2915
rect 4825 2895 4830 2915
rect 4800 2865 4830 2895
rect 4800 2845 4805 2865
rect 4825 2845 4830 2865
rect 4800 2835 4830 2845
rect 4890 2915 4920 2925
rect 4890 2895 4895 2915
rect 4915 2895 4920 2915
rect 4890 2865 4920 2895
rect 4890 2845 4895 2865
rect 4915 2845 4920 2865
rect 4890 2835 4920 2845
rect 4980 2915 5050 2925
rect 4980 2895 4985 2915
rect 5005 2895 5025 2915
rect 5045 2895 5050 2915
rect 9899 2900 10040 2940
rect 10115 2960 10155 2970
rect 10115 2940 10125 2960
rect 10145 2940 10155 2960
rect 10115 2930 10155 2940
rect 10265 2960 10305 2970
rect 10265 2940 10275 2960
rect 10295 2940 10305 2960
rect 10265 2930 10305 2940
rect 10375 2960 10415 2970
rect 10375 2940 10385 2960
rect 10405 2940 10415 2960
rect 10375 2930 10415 2940
rect 10485 2960 10525 2970
rect 10485 2940 10495 2960
rect 10515 2940 10525 2960
rect 10485 2930 10525 2940
rect 10595 2960 10635 2970
rect 10595 2940 10605 2960
rect 10625 2940 10635 2960
rect 10595 2930 10635 2940
rect 10653 2960 10687 2970
rect 10653 2940 10661 2960
rect 10679 2940 10687 2960
rect 10653 2930 10687 2940
rect 10705 2960 10745 2970
rect 10705 2940 10715 2960
rect 10735 2940 10745 2960
rect 10705 2930 10745 2940
rect 10855 2960 10895 2970
rect 10855 2940 10865 2960
rect 10885 2940 10895 2960
rect 12905 2960 12945 2970
rect 10855 2930 10895 2940
rect 11180 2940 11220 2950
rect 11180 2920 11190 2940
rect 11210 2920 11220 2940
rect 11180 2910 11220 2920
rect 11340 2940 11380 2950
rect 11340 2920 11350 2940
rect 11370 2920 11380 2940
rect 11340 2910 11380 2920
rect 11460 2940 11500 2950
rect 11460 2920 11470 2940
rect 11490 2920 11500 2940
rect 11460 2910 11500 2920
rect 11580 2940 11620 2950
rect 11580 2920 11590 2940
rect 11610 2920 11620 2940
rect 11580 2910 11620 2920
rect 11700 2940 11740 2950
rect 11700 2920 11710 2940
rect 11730 2920 11740 2940
rect 11700 2910 11740 2920
rect 11820 2940 11860 2950
rect 11820 2920 11830 2940
rect 11850 2920 11860 2940
rect 11820 2910 11860 2920
rect 11940 2940 11980 2950
rect 11940 2920 11950 2940
rect 11970 2920 11980 2940
rect 11940 2910 11980 2920
rect 12060 2940 12100 2950
rect 12060 2920 12070 2940
rect 12090 2920 12100 2940
rect 12060 2910 12100 2920
rect 12180 2940 12220 2950
rect 12180 2920 12190 2940
rect 12210 2920 12220 2940
rect 12180 2910 12220 2920
rect 12300 2940 12340 2950
rect 12300 2920 12310 2940
rect 12330 2920 12340 2940
rect 12300 2910 12340 2920
rect 12420 2940 12460 2950
rect 12420 2920 12430 2940
rect 12450 2920 12460 2940
rect 12420 2910 12460 2920
rect 12480 2910 12520 2950
rect 12580 2940 12620 2950
rect 12580 2920 12590 2940
rect 12610 2920 12620 2940
rect 12905 2940 12915 2960
rect 12935 2940 12945 2960
rect 12905 2930 12945 2940
rect 13055 2960 13095 2970
rect 13055 2940 13065 2960
rect 13085 2940 13095 2960
rect 13055 2930 13095 2940
rect 13113 2960 13147 2970
rect 13113 2940 13121 2960
rect 13139 2940 13147 2960
rect 13113 2930 13147 2940
rect 13165 2960 13205 2970
rect 13165 2940 13175 2960
rect 13195 2940 13205 2960
rect 13165 2930 13205 2940
rect 13275 2960 13315 2970
rect 13275 2940 13285 2960
rect 13305 2940 13315 2960
rect 13275 2930 13315 2940
rect 13385 2960 13425 2970
rect 13385 2940 13395 2960
rect 13415 2940 13425 2960
rect 13385 2930 13425 2940
rect 13495 2960 13535 2970
rect 13495 2940 13505 2960
rect 13525 2940 13535 2960
rect 13495 2930 13535 2940
rect 13645 2960 13685 2970
rect 13645 2940 13655 2960
rect 13675 2940 13685 2960
rect 13645 2930 13685 2940
rect 26280 3150 26320 3160
rect 26280 3130 26290 3150
rect 26310 3130 26320 3150
rect 26280 3120 26320 3130
rect 26400 3150 26440 3160
rect 26400 3130 26410 3150
rect 26430 3130 26440 3150
rect 26400 3120 26440 3130
rect 26520 3150 26560 3160
rect 26520 3130 26530 3150
rect 26550 3130 26560 3150
rect 26520 3120 26560 3130
rect 26640 3150 26680 3160
rect 26640 3130 26650 3150
rect 26670 3130 26680 3150
rect 26640 3120 26680 3130
rect 26760 3150 26800 3160
rect 26760 3130 26770 3150
rect 26790 3130 26800 3150
rect 26760 3120 26800 3130
rect 26823 3150 26857 3160
rect 26823 3130 26831 3150
rect 26849 3130 26857 3150
rect 26823 3120 26857 3130
rect 26880 3150 26920 3160
rect 26880 3130 26890 3150
rect 26910 3130 26920 3150
rect 26880 3120 26920 3130
rect 27000 3150 27040 3160
rect 27000 3130 27010 3150
rect 27030 3130 27040 3150
rect 27000 3120 27040 3130
rect 27120 3150 27160 3160
rect 27120 3130 27130 3150
rect 27150 3130 27160 3150
rect 27120 3120 27160 3130
rect 27240 3150 27280 3160
rect 27240 3130 27250 3150
rect 27270 3130 27280 3150
rect 27240 3120 27280 3130
rect 27360 3150 27400 3160
rect 27360 3130 27370 3150
rect 27390 3130 27400 3150
rect 27360 3120 27400 3130
rect 27480 3150 27520 3160
rect 27480 3130 27490 3150
rect 27510 3130 27520 3150
rect 27480 3120 27520 3130
rect 27855 3155 27860 3175
rect 27880 3155 27900 3175
rect 27920 3155 27925 3175
rect 27855 3125 27925 3155
rect 27855 3105 27860 3125
rect 27880 3105 27900 3125
rect 27920 3105 27925 3125
rect 27855 3075 27925 3105
rect 27855 3055 27860 3075
rect 27880 3055 27900 3075
rect 27920 3055 27925 3075
rect 27855 3025 27925 3055
rect 27855 3005 27860 3025
rect 27880 3005 27900 3025
rect 27920 3005 27925 3025
rect 27855 2975 27925 3005
rect 27855 2955 27860 2975
rect 27880 2955 27900 2975
rect 27920 2955 27925 2975
rect 12580 2910 12620 2920
rect 4980 2865 5050 2895
rect 11190 2890 11210 2910
rect 11350 2890 11370 2910
rect 11470 2890 11490 2910
rect 11590 2890 11610 2910
rect 11710 2890 11730 2910
rect 11830 2890 11850 2910
rect 11950 2890 11970 2910
rect 12070 2890 12090 2910
rect 12190 2890 12210 2910
rect 12310 2890 12330 2910
rect 12430 2890 12450 2910
rect 12590 2890 12610 2910
rect 13760 2900 13901 2940
rect 26180 2940 26220 2950
rect 26180 2920 26190 2940
rect 26210 2920 26220 2940
rect 26180 2910 26220 2920
rect 26340 2940 26380 2950
rect 26340 2920 26350 2940
rect 26370 2920 26380 2940
rect 26340 2910 26380 2920
rect 26460 2940 26500 2950
rect 26460 2920 26470 2940
rect 26490 2920 26500 2940
rect 26460 2910 26500 2920
rect 26580 2940 26620 2950
rect 26580 2920 26590 2940
rect 26610 2920 26620 2940
rect 26580 2910 26620 2920
rect 26700 2940 26740 2950
rect 26700 2920 26710 2940
rect 26730 2920 26740 2940
rect 26700 2910 26740 2920
rect 26820 2940 26860 2950
rect 26820 2920 26830 2940
rect 26850 2920 26860 2940
rect 26820 2910 26860 2920
rect 26940 2940 26980 2950
rect 26940 2920 26950 2940
rect 26970 2920 26980 2940
rect 26940 2910 26980 2920
rect 27060 2940 27100 2950
rect 27060 2920 27070 2940
rect 27090 2920 27100 2940
rect 27060 2910 27100 2920
rect 27180 2940 27220 2950
rect 27180 2920 27190 2940
rect 27210 2920 27220 2940
rect 27180 2910 27220 2920
rect 27300 2940 27340 2950
rect 27300 2920 27310 2940
rect 27330 2920 27340 2940
rect 27300 2910 27340 2920
rect 27420 2940 27460 2950
rect 27420 2920 27430 2940
rect 27450 2920 27460 2940
rect 27420 2910 27460 2920
rect 27480 2910 27520 2950
rect 27580 2940 27620 2950
rect 27855 2945 27925 2955
rect 27950 3225 27980 3235
rect 27950 3205 27955 3225
rect 27975 3205 27980 3225
rect 27950 3175 27980 3205
rect 27950 3155 27955 3175
rect 27975 3155 27980 3175
rect 27950 3125 27980 3155
rect 27950 3105 27955 3125
rect 27975 3105 27980 3125
rect 27950 3075 27980 3105
rect 27950 3055 27955 3075
rect 27975 3055 27980 3075
rect 27950 3025 27980 3055
rect 27950 3005 27955 3025
rect 27975 3005 27980 3025
rect 27950 2975 27980 3005
rect 27950 2955 27955 2975
rect 27975 2955 27980 2975
rect 27950 2945 27980 2955
rect 28005 3225 28035 3235
rect 28005 3205 28010 3225
rect 28030 3205 28035 3225
rect 28005 3175 28035 3205
rect 28005 3155 28010 3175
rect 28030 3155 28035 3175
rect 28005 3125 28035 3155
rect 28005 3105 28010 3125
rect 28030 3105 28035 3125
rect 28005 3075 28035 3105
rect 28005 3055 28010 3075
rect 28030 3055 28035 3075
rect 28005 3025 28035 3055
rect 28005 3005 28010 3025
rect 28030 3005 28035 3025
rect 28005 2975 28035 3005
rect 28005 2955 28010 2975
rect 28030 2955 28035 2975
rect 28005 2945 28035 2955
rect 28060 3225 28090 3235
rect 28060 3205 28065 3225
rect 28085 3205 28090 3225
rect 28060 3175 28090 3205
rect 28060 3155 28065 3175
rect 28085 3155 28090 3175
rect 28060 3125 28090 3155
rect 28060 3105 28065 3125
rect 28085 3105 28090 3125
rect 28060 3075 28090 3105
rect 28060 3055 28065 3075
rect 28085 3055 28090 3075
rect 28060 3025 28090 3055
rect 28060 3005 28065 3025
rect 28085 3005 28090 3025
rect 28060 2975 28090 3005
rect 28060 2955 28065 2975
rect 28085 2955 28090 2975
rect 28060 2945 28090 2955
rect 28115 3225 28145 3235
rect 28115 3205 28120 3225
rect 28140 3205 28145 3225
rect 28115 3175 28145 3205
rect 28115 3155 28120 3175
rect 28140 3155 28145 3175
rect 28115 3125 28145 3155
rect 28115 3105 28120 3125
rect 28140 3105 28145 3125
rect 28115 3075 28145 3105
rect 28115 3055 28120 3075
rect 28140 3055 28145 3075
rect 28115 3025 28145 3055
rect 28115 3005 28120 3025
rect 28140 3005 28145 3025
rect 28115 2975 28145 3005
rect 28115 2955 28120 2975
rect 28140 2955 28145 2975
rect 28115 2945 28145 2955
rect 28170 3225 28200 3235
rect 28170 3205 28175 3225
rect 28195 3205 28200 3225
rect 28170 3175 28200 3205
rect 28170 3155 28175 3175
rect 28195 3155 28200 3175
rect 28170 3125 28200 3155
rect 28170 3105 28175 3125
rect 28195 3105 28200 3125
rect 28170 3075 28200 3105
rect 28170 3055 28175 3075
rect 28195 3055 28200 3075
rect 28170 3025 28200 3055
rect 28170 3005 28175 3025
rect 28195 3005 28200 3025
rect 28170 2975 28200 3005
rect 28170 2955 28175 2975
rect 28195 2955 28200 2975
rect 28170 2945 28200 2955
rect 28225 3225 28255 3235
rect 28225 3205 28230 3225
rect 28250 3205 28255 3225
rect 28225 3175 28255 3205
rect 28225 3155 28230 3175
rect 28250 3155 28255 3175
rect 28225 3125 28255 3155
rect 28225 3105 28230 3125
rect 28250 3105 28255 3125
rect 28225 3075 28255 3105
rect 28225 3055 28230 3075
rect 28250 3055 28255 3075
rect 28225 3025 28255 3055
rect 28225 3005 28230 3025
rect 28250 3005 28255 3025
rect 28225 2975 28255 3005
rect 28225 2955 28230 2975
rect 28250 2955 28255 2975
rect 28225 2945 28255 2955
rect 28280 3225 28310 3235
rect 28280 3205 28285 3225
rect 28305 3205 28310 3225
rect 28280 3175 28310 3205
rect 28280 3155 28285 3175
rect 28305 3155 28310 3175
rect 28280 3125 28310 3155
rect 28280 3105 28285 3125
rect 28305 3105 28310 3125
rect 28280 3075 28310 3105
rect 28280 3055 28285 3075
rect 28305 3055 28310 3075
rect 28280 3025 28310 3055
rect 28280 3005 28285 3025
rect 28305 3005 28310 3025
rect 28280 2975 28310 3005
rect 28280 2955 28285 2975
rect 28305 2955 28310 2975
rect 28280 2945 28310 2955
rect 28335 3225 28365 3235
rect 28335 3205 28340 3225
rect 28360 3205 28365 3225
rect 28335 3175 28365 3205
rect 28335 3155 28340 3175
rect 28360 3155 28365 3175
rect 28335 3125 28365 3155
rect 28335 3105 28340 3125
rect 28360 3105 28365 3125
rect 28335 3075 28365 3105
rect 28335 3055 28340 3075
rect 28360 3055 28365 3075
rect 28335 3025 28365 3055
rect 28335 3005 28340 3025
rect 28360 3005 28365 3025
rect 28335 2975 28365 3005
rect 28335 2955 28340 2975
rect 28360 2955 28365 2975
rect 28335 2945 28365 2955
rect 28390 3225 28420 3235
rect 28390 3205 28395 3225
rect 28415 3205 28420 3225
rect 28390 3175 28420 3205
rect 28390 3155 28395 3175
rect 28415 3155 28420 3175
rect 28390 3125 28420 3155
rect 28390 3105 28395 3125
rect 28415 3105 28420 3125
rect 28390 3075 28420 3105
rect 28390 3055 28395 3075
rect 28415 3055 28420 3075
rect 28390 3025 28420 3055
rect 28390 3005 28395 3025
rect 28415 3005 28420 3025
rect 28390 2975 28420 3005
rect 28390 2955 28395 2975
rect 28415 2955 28420 2975
rect 28390 2945 28420 2955
rect 28445 3225 28475 3235
rect 28445 3205 28450 3225
rect 28470 3205 28475 3225
rect 28445 3175 28475 3205
rect 28445 3155 28450 3175
rect 28470 3155 28475 3175
rect 28445 3125 28475 3155
rect 28445 3105 28450 3125
rect 28470 3105 28475 3125
rect 28445 3075 28475 3105
rect 28445 3055 28450 3075
rect 28470 3055 28475 3075
rect 28445 3025 28475 3055
rect 28445 3005 28450 3025
rect 28470 3005 28475 3025
rect 28445 2975 28475 3005
rect 28445 2955 28450 2975
rect 28470 2955 28475 2975
rect 28445 2945 28475 2955
rect 28500 3225 28530 3235
rect 28500 3205 28505 3225
rect 28525 3205 28530 3225
rect 28500 3175 28530 3205
rect 28500 3155 28505 3175
rect 28525 3155 28530 3175
rect 28500 3125 28530 3155
rect 28500 3105 28505 3125
rect 28525 3105 28530 3125
rect 28500 3075 28530 3105
rect 28500 3055 28505 3075
rect 28525 3055 28530 3075
rect 28500 3025 28530 3055
rect 28500 3005 28505 3025
rect 28525 3005 28530 3025
rect 28500 2975 28530 3005
rect 28500 2955 28505 2975
rect 28525 2955 28530 2975
rect 28500 2945 28530 2955
rect 28555 3225 28585 3235
rect 28555 3205 28560 3225
rect 28580 3205 28585 3225
rect 28555 3175 28585 3205
rect 28555 3155 28560 3175
rect 28580 3155 28585 3175
rect 28555 3125 28585 3155
rect 28555 3105 28560 3125
rect 28580 3105 28585 3125
rect 28555 3075 28585 3105
rect 28555 3055 28560 3075
rect 28580 3055 28585 3075
rect 28555 3025 28585 3055
rect 28555 3005 28560 3025
rect 28580 3005 28585 3025
rect 28555 2975 28585 3005
rect 28555 2955 28560 2975
rect 28580 2955 28585 2975
rect 28555 2945 28585 2955
rect 28610 3225 28640 3235
rect 28610 3205 28615 3225
rect 28635 3205 28640 3225
rect 28610 3175 28640 3205
rect 28610 3155 28615 3175
rect 28635 3155 28640 3175
rect 28610 3125 28640 3155
rect 28610 3105 28615 3125
rect 28635 3105 28640 3125
rect 28610 3075 28640 3105
rect 28610 3055 28615 3075
rect 28635 3055 28640 3075
rect 28610 3025 28640 3055
rect 28610 3005 28615 3025
rect 28635 3005 28640 3025
rect 28610 2975 28640 3005
rect 28610 2955 28615 2975
rect 28635 2955 28640 2975
rect 28610 2945 28640 2955
rect 28665 3225 28695 3235
rect 28665 3205 28670 3225
rect 28690 3205 28695 3225
rect 28665 3175 28695 3205
rect 28665 3155 28670 3175
rect 28690 3155 28695 3175
rect 28665 3125 28695 3155
rect 28665 3105 28670 3125
rect 28690 3105 28695 3125
rect 28665 3075 28695 3105
rect 28665 3055 28670 3075
rect 28690 3055 28695 3075
rect 28665 3025 28695 3055
rect 28665 3005 28670 3025
rect 28690 3005 28695 3025
rect 28665 2975 28695 3005
rect 28665 2955 28670 2975
rect 28690 2955 28695 2975
rect 28665 2945 28695 2955
rect 28720 3225 28750 3235
rect 28720 3205 28725 3225
rect 28745 3205 28750 3225
rect 28720 3175 28750 3205
rect 28720 3155 28725 3175
rect 28745 3155 28750 3175
rect 28720 3125 28750 3155
rect 28720 3105 28725 3125
rect 28745 3105 28750 3125
rect 28720 3075 28750 3105
rect 28720 3055 28725 3075
rect 28745 3055 28750 3075
rect 28720 3025 28750 3055
rect 28720 3005 28725 3025
rect 28745 3005 28750 3025
rect 28720 2975 28750 3005
rect 28720 2955 28725 2975
rect 28745 2955 28750 2975
rect 28720 2945 28750 2955
rect 28775 3225 28805 3235
rect 28775 3205 28780 3225
rect 28800 3205 28805 3225
rect 28775 3175 28805 3205
rect 28775 3155 28780 3175
rect 28800 3155 28805 3175
rect 28775 3125 28805 3155
rect 28775 3105 28780 3125
rect 28800 3105 28805 3125
rect 28775 3075 28805 3105
rect 28775 3055 28780 3075
rect 28800 3055 28805 3075
rect 28775 3025 28805 3055
rect 28775 3005 28780 3025
rect 28800 3005 28805 3025
rect 28775 2975 28805 3005
rect 28775 2955 28780 2975
rect 28800 2955 28805 2975
rect 28775 2945 28805 2955
rect 28830 3225 28860 3235
rect 28830 3205 28835 3225
rect 28855 3205 28860 3225
rect 28830 3175 28860 3205
rect 28830 3155 28835 3175
rect 28855 3155 28860 3175
rect 28830 3125 28860 3155
rect 28830 3105 28835 3125
rect 28855 3105 28860 3125
rect 28830 3075 28860 3105
rect 28830 3055 28835 3075
rect 28855 3055 28860 3075
rect 28830 3025 28860 3055
rect 28830 3005 28835 3025
rect 28855 3005 28860 3025
rect 28830 2975 28860 3005
rect 28830 2955 28835 2975
rect 28855 2955 28860 2975
rect 28830 2945 28860 2955
rect 28885 3225 28915 3235
rect 28885 3205 28890 3225
rect 28910 3205 28915 3225
rect 28885 3175 28915 3205
rect 28885 3155 28890 3175
rect 28910 3155 28915 3175
rect 28885 3125 28915 3155
rect 28885 3105 28890 3125
rect 28910 3105 28915 3125
rect 28885 3075 28915 3105
rect 28885 3055 28890 3075
rect 28910 3055 28915 3075
rect 28885 3025 28915 3055
rect 28885 3005 28890 3025
rect 28910 3005 28915 3025
rect 28885 2975 28915 3005
rect 28885 2955 28890 2975
rect 28910 2955 28915 2975
rect 28885 2945 28915 2955
rect 28940 3225 28970 3235
rect 28940 3205 28945 3225
rect 28965 3205 28970 3225
rect 28940 3175 28970 3205
rect 28940 3155 28945 3175
rect 28965 3155 28970 3175
rect 28940 3125 28970 3155
rect 28940 3105 28945 3125
rect 28965 3105 28970 3125
rect 28940 3075 28970 3105
rect 28940 3055 28945 3075
rect 28965 3055 28970 3075
rect 28940 3025 28970 3055
rect 28940 3005 28945 3025
rect 28965 3005 28970 3025
rect 28940 2975 28970 3005
rect 28940 2955 28945 2975
rect 28965 2955 28970 2975
rect 28940 2945 28970 2955
rect 28995 3225 29025 3235
rect 28995 3205 29000 3225
rect 29020 3205 29025 3225
rect 28995 3175 29025 3205
rect 28995 3155 29000 3175
rect 29020 3155 29025 3175
rect 28995 3125 29025 3155
rect 28995 3105 29000 3125
rect 29020 3105 29025 3125
rect 28995 3075 29025 3105
rect 28995 3055 29000 3075
rect 29020 3055 29025 3075
rect 28995 3025 29025 3055
rect 28995 3005 29000 3025
rect 29020 3005 29025 3025
rect 28995 2975 29025 3005
rect 28995 2955 29000 2975
rect 29020 2955 29025 2975
rect 28995 2945 29025 2955
rect 29050 3225 29080 3235
rect 29050 3205 29055 3225
rect 29075 3205 29080 3225
rect 29050 3175 29080 3205
rect 29050 3155 29055 3175
rect 29075 3155 29080 3175
rect 29050 3125 29080 3155
rect 29050 3105 29055 3125
rect 29075 3105 29080 3125
rect 29050 3075 29080 3105
rect 29050 3055 29055 3075
rect 29075 3055 29080 3075
rect 29050 3025 29080 3055
rect 29050 3005 29055 3025
rect 29075 3005 29080 3025
rect 29050 2975 29080 3005
rect 29050 2955 29055 2975
rect 29075 2955 29080 2975
rect 29050 2945 29080 2955
rect 29105 3225 29175 3235
rect 29105 3205 29110 3225
rect 29130 3205 29150 3225
rect 29170 3205 29175 3225
rect 29105 3175 29175 3205
rect 29105 3155 29110 3175
rect 29130 3155 29150 3175
rect 29170 3155 29175 3175
rect 29105 3125 29175 3155
rect 29105 3105 29110 3125
rect 29130 3105 29150 3125
rect 29170 3105 29175 3125
rect 29105 3075 29175 3105
rect 29105 3055 29110 3075
rect 29130 3055 29150 3075
rect 29170 3055 29175 3075
rect 29105 3025 29175 3055
rect 29105 3005 29110 3025
rect 29130 3005 29150 3025
rect 29170 3005 29175 3025
rect 29105 2975 29175 3005
rect 29105 2955 29110 2975
rect 29130 2955 29150 2975
rect 29170 2955 29175 2975
rect 29105 2945 29175 2955
rect 27580 2920 27590 2940
rect 27610 2920 27620 2940
rect 27860 2925 27880 2945
rect 28010 2925 28030 2945
rect 28120 2925 28140 2945
rect 28230 2925 28250 2945
rect 28340 2925 28360 2945
rect 28450 2925 28470 2945
rect 28560 2925 28580 2945
rect 28670 2925 28690 2945
rect 28780 2925 28800 2945
rect 28890 2925 28910 2945
rect 29000 2925 29020 2945
rect 29150 2925 29170 2945
rect 27580 2910 27620 2920
rect 27850 2915 27890 2925
rect 26190 2890 26210 2910
rect 26350 2890 26370 2910
rect 26470 2890 26490 2910
rect 26590 2890 26610 2910
rect 26710 2890 26730 2910
rect 26830 2890 26850 2910
rect 26950 2890 26970 2910
rect 27070 2890 27090 2910
rect 27190 2890 27210 2910
rect 27310 2890 27330 2910
rect 27430 2890 27450 2910
rect 27590 2890 27610 2910
rect 27850 2895 27860 2915
rect 27880 2895 27890 2915
rect 4980 2845 4985 2865
rect 5005 2845 5025 2865
rect 5045 2845 5050 2865
rect 4980 2835 5050 2845
rect 11185 2880 11255 2890
rect 11185 2860 11190 2880
rect 11210 2860 11230 2880
rect 11250 2860 11255 2880
rect 3005 2815 3025 2835
rect 3185 2815 3205 2835
rect 3365 2815 3385 2835
rect 3545 2815 3565 2835
rect 3725 2815 3745 2835
rect 3905 2815 3925 2835
rect 4085 2815 4105 2835
rect 4265 2815 4285 2835
rect 4445 2815 4465 2835
rect 4625 2815 4645 2835
rect 4805 2815 4825 2835
rect 4985 2815 5005 2835
rect 11185 2830 11255 2860
rect 2995 2805 3035 2815
rect -10 2765 20 2795
rect 51 2790 96 2795
rect 51 2765 61 2790
rect 86 2765 96 2790
rect 51 2760 96 2765
rect 724 2790 769 2795
rect 724 2765 734 2790
rect 759 2765 769 2790
rect 724 2760 769 2765
rect 2620 2755 2660 2795
rect 2995 2785 3005 2805
rect 3025 2785 3035 2805
rect 2995 2775 3035 2785
rect 3175 2805 3215 2815
rect 3175 2785 3185 2805
rect 3205 2785 3215 2805
rect 3175 2775 3215 2785
rect 3355 2805 3395 2815
rect 3355 2785 3365 2805
rect 3385 2785 3395 2805
rect 3355 2775 3395 2785
rect 3535 2805 3575 2815
rect 3535 2785 3545 2805
rect 3565 2785 3575 2805
rect 3535 2775 3575 2785
rect 3715 2805 3755 2815
rect 3715 2785 3725 2805
rect 3745 2785 3755 2805
rect 3715 2775 3755 2785
rect 3895 2805 3935 2815
rect 3895 2785 3905 2805
rect 3925 2785 3935 2805
rect 3895 2775 3935 2785
rect 4075 2805 4115 2815
rect 4075 2785 4085 2805
rect 4105 2785 4115 2805
rect 4075 2775 4115 2785
rect 4255 2805 4295 2815
rect 4255 2785 4265 2805
rect 4285 2785 4295 2805
rect 4255 2775 4295 2785
rect 4435 2805 4475 2815
rect 4435 2785 4445 2805
rect 4465 2785 4475 2805
rect 4435 2775 4475 2785
rect 4615 2805 4655 2815
rect 4615 2785 4625 2805
rect 4645 2785 4655 2805
rect 4615 2775 4655 2785
rect 4795 2805 4835 2815
rect 4795 2785 4805 2805
rect 4825 2785 4835 2805
rect 4795 2775 4835 2785
rect 4975 2805 5015 2815
rect 4975 2785 4985 2805
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 11185 2810 11190 2830
rect 11210 2810 11230 2830
rect 11250 2810 11255 2830
rect 11185 2780 11255 2810
rect 11185 2760 11190 2780
rect 11210 2760 11230 2780
rect 11250 2760 11255 2780
rect 1266 2715 1296 2745
rect 2150 2710 2190 2750
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2725 3215 2745
rect 3175 2715 3215 2725
rect 3355 2745 3395 2755
rect 3355 2725 3365 2745
rect 3385 2725 3395 2745
rect 3355 2715 3395 2725
rect 3535 2745 3575 2755
rect 3535 2725 3545 2745
rect 3565 2725 3575 2745
rect 3535 2715 3575 2725
rect 3715 2745 3755 2755
rect 3715 2725 3725 2745
rect 3745 2725 3755 2745
rect 3715 2715 3755 2725
rect 3895 2745 3935 2755
rect 3895 2725 3905 2745
rect 3925 2725 3935 2745
rect 3895 2715 3935 2725
rect 4075 2745 4115 2755
rect 4075 2725 4085 2745
rect 4105 2725 4115 2745
rect 4075 2715 4115 2725
rect 4255 2745 4295 2755
rect 4255 2725 4265 2745
rect 4285 2725 4295 2745
rect 4255 2715 4295 2725
rect 4435 2745 4475 2755
rect 4435 2725 4445 2745
rect 4465 2725 4475 2745
rect 4435 2715 4475 2725
rect 4615 2745 4655 2755
rect 4615 2725 4625 2745
rect 4645 2725 4655 2745
rect 4615 2715 4655 2725
rect 4795 2745 4835 2755
rect 4795 2725 4805 2745
rect 4825 2725 4835 2745
rect 4795 2715 4835 2725
rect 11185 2730 11255 2760
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3185 2695 3205 2715
rect 3365 2695 3385 2715
rect 3545 2695 3565 2715
rect 3725 2695 3745 2715
rect 3905 2695 3925 2715
rect 4085 2695 4105 2715
rect 4265 2695 4285 2715
rect 4445 2695 4465 2715
rect 4625 2695 4645 2715
rect 4805 2695 4825 2715
rect 11185 2710 11190 2730
rect 11210 2710 11230 2730
rect 11250 2710 11255 2730
rect 10210 2700 10250 2710
rect 3140 2685 3210 2695
rect 3140 2665 3145 2685
rect 3165 2665 3185 2685
rect 3205 2665 3210 2685
rect 3140 2635 3210 2665
rect 3140 2615 3145 2635
rect 3165 2615 3185 2635
rect 3205 2615 3210 2635
rect 3140 2585 3210 2615
rect 3140 2565 3145 2585
rect 3165 2565 3185 2585
rect 3205 2565 3210 2585
rect 3140 2535 3210 2565
rect 3140 2515 3145 2535
rect 3165 2515 3185 2535
rect 3205 2515 3210 2535
rect 3140 2485 3210 2515
rect 3140 2465 3145 2485
rect 3165 2465 3185 2485
rect 3205 2465 3210 2485
rect 3140 2435 3210 2465
rect 3140 2415 3145 2435
rect 3165 2415 3185 2435
rect 3205 2415 3210 2435
rect 3140 2405 3210 2415
rect 3270 2685 3300 2695
rect 3270 2665 3275 2685
rect 3295 2665 3300 2685
rect 3270 2635 3300 2665
rect 3270 2615 3275 2635
rect 3295 2615 3300 2635
rect 3270 2585 3300 2615
rect 3270 2565 3275 2585
rect 3295 2565 3300 2585
rect 3270 2535 3300 2565
rect 3270 2515 3275 2535
rect 3295 2515 3300 2535
rect 3270 2485 3300 2515
rect 3270 2465 3275 2485
rect 3295 2465 3300 2485
rect 3270 2435 3300 2465
rect 3270 2415 3275 2435
rect 3295 2415 3300 2435
rect 3270 2405 3300 2415
rect 3360 2685 3390 2695
rect 3360 2665 3365 2685
rect 3385 2665 3390 2685
rect 3360 2635 3390 2665
rect 3360 2615 3365 2635
rect 3385 2615 3390 2635
rect 3360 2585 3390 2615
rect 3360 2565 3365 2585
rect 3385 2565 3390 2585
rect 3360 2535 3390 2565
rect 3360 2515 3365 2535
rect 3385 2515 3390 2535
rect 3360 2485 3390 2515
rect 3360 2465 3365 2485
rect 3385 2465 3390 2485
rect 3360 2435 3390 2465
rect 3360 2415 3365 2435
rect 3385 2415 3390 2435
rect 3360 2405 3390 2415
rect 3450 2685 3480 2695
rect 3450 2665 3455 2685
rect 3475 2665 3480 2685
rect 3450 2635 3480 2665
rect 3450 2615 3455 2635
rect 3475 2615 3480 2635
rect 3450 2585 3480 2615
rect 3450 2565 3455 2585
rect 3475 2565 3480 2585
rect 3450 2535 3480 2565
rect 3450 2515 3455 2535
rect 3475 2515 3480 2535
rect 3450 2485 3480 2515
rect 3450 2465 3455 2485
rect 3475 2465 3480 2485
rect 3450 2435 3480 2465
rect 3450 2415 3455 2435
rect 3475 2415 3480 2435
rect 3450 2405 3480 2415
rect 3540 2685 3570 2695
rect 3540 2665 3545 2685
rect 3565 2665 3570 2685
rect 3540 2635 3570 2665
rect 3540 2615 3545 2635
rect 3565 2615 3570 2635
rect 3540 2585 3570 2615
rect 3540 2565 3545 2585
rect 3565 2565 3570 2585
rect 3540 2535 3570 2565
rect 3540 2515 3545 2535
rect 3565 2515 3570 2535
rect 3540 2485 3570 2515
rect 3540 2465 3545 2485
rect 3565 2465 3570 2485
rect 3540 2435 3570 2465
rect 3540 2415 3545 2435
rect 3565 2415 3570 2435
rect 3540 2405 3570 2415
rect 3630 2685 3660 2695
rect 3630 2665 3635 2685
rect 3655 2665 3660 2685
rect 3630 2635 3660 2665
rect 3630 2615 3635 2635
rect 3655 2615 3660 2635
rect 3630 2585 3660 2615
rect 3630 2565 3635 2585
rect 3655 2565 3660 2585
rect 3630 2535 3660 2565
rect 3630 2515 3635 2535
rect 3655 2515 3660 2535
rect 3630 2485 3660 2515
rect 3630 2465 3635 2485
rect 3655 2465 3660 2485
rect 3630 2435 3660 2465
rect 3630 2415 3635 2435
rect 3655 2415 3660 2435
rect 3630 2405 3660 2415
rect 3720 2685 3750 2695
rect 3720 2665 3725 2685
rect 3745 2665 3750 2685
rect 3720 2635 3750 2665
rect 3720 2615 3725 2635
rect 3745 2615 3750 2635
rect 3720 2585 3750 2615
rect 3720 2565 3725 2585
rect 3745 2565 3750 2585
rect 3720 2535 3750 2565
rect 3720 2515 3725 2535
rect 3745 2515 3750 2535
rect 3720 2485 3750 2515
rect 3720 2465 3725 2485
rect 3745 2465 3750 2485
rect 3720 2435 3750 2465
rect 3720 2415 3725 2435
rect 3745 2415 3750 2435
rect 3720 2405 3750 2415
rect 3810 2685 3840 2695
rect 3810 2665 3815 2685
rect 3835 2665 3840 2685
rect 3810 2635 3840 2665
rect 3810 2615 3815 2635
rect 3835 2615 3840 2635
rect 3810 2585 3840 2615
rect 3810 2565 3815 2585
rect 3835 2565 3840 2585
rect 3810 2535 3840 2565
rect 3810 2515 3815 2535
rect 3835 2515 3840 2535
rect 3810 2485 3840 2515
rect 3810 2465 3815 2485
rect 3835 2465 3840 2485
rect 3810 2435 3840 2465
rect 3810 2415 3815 2435
rect 3835 2415 3840 2435
rect 3810 2405 3840 2415
rect 3900 2685 3930 2695
rect 3900 2665 3905 2685
rect 3925 2665 3930 2685
rect 3900 2635 3930 2665
rect 3900 2615 3905 2635
rect 3925 2615 3930 2635
rect 3900 2585 3930 2615
rect 3900 2565 3905 2585
rect 3925 2565 3930 2585
rect 3900 2535 3930 2565
rect 3900 2515 3905 2535
rect 3925 2515 3930 2535
rect 3900 2485 3930 2515
rect 3900 2465 3905 2485
rect 3925 2465 3930 2485
rect 3900 2435 3930 2465
rect 3900 2415 3905 2435
rect 3925 2415 3930 2435
rect 3900 2405 3930 2415
rect 3990 2685 4020 2695
rect 3990 2665 3995 2685
rect 4015 2665 4020 2685
rect 3990 2635 4020 2665
rect 3990 2615 3995 2635
rect 4015 2615 4020 2635
rect 3990 2585 4020 2615
rect 3990 2565 3995 2585
rect 4015 2565 4020 2585
rect 3990 2535 4020 2565
rect 3990 2515 3995 2535
rect 4015 2515 4020 2535
rect 3990 2485 4020 2515
rect 3990 2465 3995 2485
rect 4015 2465 4020 2485
rect 3990 2435 4020 2465
rect 3990 2415 3995 2435
rect 4015 2415 4020 2435
rect 3990 2405 4020 2415
rect 4080 2685 4110 2695
rect 4080 2665 4085 2685
rect 4105 2665 4110 2685
rect 4080 2635 4110 2665
rect 4080 2615 4085 2635
rect 4105 2615 4110 2635
rect 4080 2585 4110 2615
rect 4080 2565 4085 2585
rect 4105 2565 4110 2585
rect 4080 2535 4110 2565
rect 4080 2515 4085 2535
rect 4105 2515 4110 2535
rect 4080 2485 4110 2515
rect 4080 2465 4085 2485
rect 4105 2465 4110 2485
rect 4080 2435 4110 2465
rect 4080 2415 4085 2435
rect 4105 2415 4110 2435
rect 4080 2405 4110 2415
rect 4170 2685 4200 2695
rect 4170 2665 4175 2685
rect 4195 2665 4200 2685
rect 4170 2635 4200 2665
rect 4170 2615 4175 2635
rect 4195 2615 4200 2635
rect 4170 2585 4200 2615
rect 4170 2565 4175 2585
rect 4195 2565 4200 2585
rect 4170 2535 4200 2565
rect 4170 2515 4175 2535
rect 4195 2515 4200 2535
rect 4170 2485 4200 2515
rect 4170 2465 4175 2485
rect 4195 2465 4200 2485
rect 4170 2435 4200 2465
rect 4170 2415 4175 2435
rect 4195 2415 4200 2435
rect 4170 2405 4200 2415
rect 4260 2685 4290 2695
rect 4260 2665 4265 2685
rect 4285 2665 4290 2685
rect 4260 2635 4290 2665
rect 4260 2615 4265 2635
rect 4285 2615 4290 2635
rect 4260 2585 4290 2615
rect 4260 2565 4265 2585
rect 4285 2565 4290 2585
rect 4260 2535 4290 2565
rect 4260 2515 4265 2535
rect 4285 2515 4290 2535
rect 4260 2485 4290 2515
rect 4260 2465 4265 2485
rect 4285 2465 4290 2485
rect 4260 2435 4290 2465
rect 4260 2415 4265 2435
rect 4285 2415 4290 2435
rect 4260 2405 4290 2415
rect 4350 2685 4380 2695
rect 4350 2665 4355 2685
rect 4375 2665 4380 2685
rect 4350 2635 4380 2665
rect 4350 2615 4355 2635
rect 4375 2615 4380 2635
rect 4350 2585 4380 2615
rect 4350 2565 4355 2585
rect 4375 2565 4380 2585
rect 4350 2535 4380 2565
rect 4350 2515 4355 2535
rect 4375 2515 4380 2535
rect 4350 2485 4380 2515
rect 4350 2465 4355 2485
rect 4375 2465 4380 2485
rect 4350 2435 4380 2465
rect 4350 2415 4355 2435
rect 4375 2415 4380 2435
rect 4350 2405 4380 2415
rect 4440 2685 4470 2695
rect 4440 2665 4445 2685
rect 4465 2665 4470 2685
rect 4440 2635 4470 2665
rect 4440 2615 4445 2635
rect 4465 2615 4470 2635
rect 4440 2585 4470 2615
rect 4440 2565 4445 2585
rect 4465 2565 4470 2585
rect 4440 2535 4470 2565
rect 4440 2515 4445 2535
rect 4465 2515 4470 2535
rect 4440 2485 4470 2515
rect 4440 2465 4445 2485
rect 4465 2465 4470 2485
rect 4440 2435 4470 2465
rect 4440 2415 4445 2435
rect 4465 2415 4470 2435
rect 4440 2405 4470 2415
rect 4530 2685 4560 2695
rect 4530 2665 4535 2685
rect 4555 2665 4560 2685
rect 4530 2635 4560 2665
rect 4530 2615 4535 2635
rect 4555 2615 4560 2635
rect 4530 2585 4560 2615
rect 4530 2565 4535 2585
rect 4555 2565 4560 2585
rect 4530 2535 4560 2565
rect 4530 2515 4535 2535
rect 4555 2515 4560 2535
rect 4530 2485 4560 2515
rect 4530 2465 4535 2485
rect 4555 2465 4560 2485
rect 4530 2435 4560 2465
rect 4530 2415 4535 2435
rect 4555 2415 4560 2435
rect 4530 2405 4560 2415
rect 4620 2685 4650 2695
rect 4620 2665 4625 2685
rect 4645 2665 4650 2685
rect 4620 2635 4650 2665
rect 4620 2615 4625 2635
rect 4645 2615 4650 2635
rect 4620 2585 4650 2615
rect 4620 2565 4625 2585
rect 4645 2565 4650 2585
rect 4620 2535 4650 2565
rect 4620 2515 4625 2535
rect 4645 2515 4650 2535
rect 4620 2485 4650 2515
rect 4620 2465 4625 2485
rect 4645 2465 4650 2485
rect 4620 2435 4650 2465
rect 4620 2415 4625 2435
rect 4645 2415 4650 2435
rect 4620 2405 4650 2415
rect 4710 2685 4740 2695
rect 4710 2665 4715 2685
rect 4735 2665 4740 2685
rect 4710 2635 4740 2665
rect 4710 2615 4715 2635
rect 4735 2615 4740 2635
rect 4710 2585 4740 2615
rect 4710 2565 4715 2585
rect 4735 2565 4740 2585
rect 4710 2535 4740 2565
rect 4710 2515 4715 2535
rect 4735 2515 4740 2535
rect 4710 2485 4740 2515
rect 4710 2465 4715 2485
rect 4735 2465 4740 2485
rect 4710 2435 4740 2465
rect 4710 2415 4715 2435
rect 4735 2415 4740 2435
rect 4710 2405 4740 2415
rect 4800 2685 4870 2695
rect 4800 2665 4805 2685
rect 4825 2665 4845 2685
rect 4865 2665 4870 2685
rect 10210 2680 10220 2700
rect 10240 2680 10250 2700
rect 10210 2670 10250 2680
rect 10320 2700 10360 2710
rect 10320 2680 10330 2700
rect 10350 2680 10360 2700
rect 10320 2670 10360 2680
rect 10430 2700 10470 2710
rect 10430 2680 10440 2700
rect 10460 2680 10470 2700
rect 10430 2670 10470 2680
rect 10540 2700 10580 2710
rect 10540 2680 10550 2700
rect 10570 2680 10580 2700
rect 10540 2670 10580 2680
rect 10650 2700 10690 2710
rect 10650 2680 10660 2700
rect 10680 2680 10690 2700
rect 10650 2670 10690 2680
rect 10760 2700 10800 2710
rect 10760 2680 10770 2700
rect 10790 2680 10800 2700
rect 10760 2670 10800 2680
rect 11185 2680 11255 2710
rect 4800 2635 4870 2665
rect 4800 2615 4805 2635
rect 4825 2615 4845 2635
rect 4865 2615 4870 2635
rect 4800 2585 4870 2615
rect 4800 2565 4805 2585
rect 4825 2565 4845 2585
rect 4865 2565 4870 2585
rect 4800 2535 4870 2565
rect 4800 2515 4805 2535
rect 4825 2515 4845 2535
rect 4865 2515 4870 2535
rect 4800 2485 4870 2515
rect 4800 2465 4805 2485
rect 4825 2465 4845 2485
rect 4865 2465 4870 2485
rect 4800 2435 4870 2465
rect 4800 2415 4805 2435
rect 4825 2415 4845 2435
rect 4865 2415 4870 2435
rect 4800 2405 4870 2415
rect 9790 2645 10005 2665
rect 10220 2650 10240 2670
rect 10330 2650 10350 2670
rect 10440 2650 10460 2670
rect 10550 2650 10570 2670
rect 10660 2650 10680 2670
rect 10770 2650 10790 2670
rect 11185 2660 11190 2680
rect 11210 2660 11230 2680
rect 11250 2660 11255 2680
rect 9790 2625 9825 2645
rect 9970 2625 10005 2645
rect 9885 2575 9910 2625
rect 10120 2640 10190 2650
rect 10120 2620 10125 2640
rect 10145 2620 10165 2640
rect 10185 2620 10190 2640
rect 10120 2590 10190 2620
rect 10120 2570 10125 2590
rect 10145 2570 10165 2590
rect 10185 2570 10190 2590
rect 10120 2540 10190 2570
rect 10120 2520 10125 2540
rect 10145 2520 10165 2540
rect 10185 2520 10190 2540
rect 10120 2490 10190 2520
rect 10120 2470 10125 2490
rect 10145 2470 10165 2490
rect 10185 2470 10190 2490
rect 10120 2460 10190 2470
rect 10215 2640 10245 2650
rect 10215 2620 10220 2640
rect 10240 2620 10245 2640
rect 10215 2590 10245 2620
rect 10215 2570 10220 2590
rect 10240 2570 10245 2590
rect 10215 2540 10245 2570
rect 10215 2520 10220 2540
rect 10240 2520 10245 2540
rect 10215 2490 10245 2520
rect 10215 2470 10220 2490
rect 10240 2470 10245 2490
rect 10215 2460 10245 2470
rect 10270 2640 10300 2650
rect 10270 2620 10275 2640
rect 10295 2620 10300 2640
rect 10270 2590 10300 2620
rect 10270 2570 10275 2590
rect 10295 2570 10300 2590
rect 10270 2540 10300 2570
rect 10270 2520 10275 2540
rect 10295 2520 10300 2540
rect 10270 2490 10300 2520
rect 10270 2470 10275 2490
rect 10295 2470 10300 2490
rect 10270 2460 10300 2470
rect 10325 2640 10355 2650
rect 10325 2620 10330 2640
rect 10350 2620 10355 2640
rect 10325 2590 10355 2620
rect 10325 2570 10330 2590
rect 10350 2570 10355 2590
rect 10325 2540 10355 2570
rect 10325 2520 10330 2540
rect 10350 2520 10355 2540
rect 10325 2490 10355 2520
rect 10325 2470 10330 2490
rect 10350 2470 10355 2490
rect 10325 2460 10355 2470
rect 10380 2640 10410 2650
rect 10380 2620 10385 2640
rect 10405 2620 10410 2640
rect 10380 2590 10410 2620
rect 10380 2570 10385 2590
rect 10405 2570 10410 2590
rect 10380 2540 10410 2570
rect 10380 2520 10385 2540
rect 10405 2520 10410 2540
rect 10380 2490 10410 2520
rect 10380 2470 10385 2490
rect 10405 2470 10410 2490
rect 10380 2460 10410 2470
rect 10435 2640 10465 2650
rect 10435 2620 10440 2640
rect 10460 2620 10465 2640
rect 10435 2590 10465 2620
rect 10435 2570 10440 2590
rect 10460 2570 10465 2590
rect 10435 2540 10465 2570
rect 10435 2520 10440 2540
rect 10460 2520 10465 2540
rect 10435 2490 10465 2520
rect 10435 2470 10440 2490
rect 10460 2470 10465 2490
rect 10435 2460 10465 2470
rect 10490 2640 10520 2650
rect 10490 2620 10495 2640
rect 10515 2620 10520 2640
rect 10490 2590 10520 2620
rect 10490 2570 10495 2590
rect 10515 2570 10520 2590
rect 10490 2540 10520 2570
rect 10490 2520 10495 2540
rect 10515 2520 10520 2540
rect 10490 2490 10520 2520
rect 10490 2470 10495 2490
rect 10515 2470 10520 2490
rect 10490 2460 10520 2470
rect 10545 2640 10575 2650
rect 10545 2620 10550 2640
rect 10570 2620 10575 2640
rect 10545 2590 10575 2620
rect 10545 2570 10550 2590
rect 10570 2570 10575 2590
rect 10545 2540 10575 2570
rect 10545 2520 10550 2540
rect 10570 2520 10575 2540
rect 10545 2490 10575 2520
rect 10545 2470 10550 2490
rect 10570 2470 10575 2490
rect 10545 2460 10575 2470
rect 10600 2640 10630 2650
rect 10600 2620 10605 2640
rect 10625 2620 10630 2640
rect 10600 2590 10630 2620
rect 10600 2570 10605 2590
rect 10625 2570 10630 2590
rect 10600 2540 10630 2570
rect 10600 2520 10605 2540
rect 10625 2520 10630 2540
rect 10600 2490 10630 2520
rect 10600 2470 10605 2490
rect 10625 2470 10630 2490
rect 10600 2460 10630 2470
rect 10655 2640 10685 2650
rect 10655 2620 10660 2640
rect 10680 2620 10685 2640
rect 10655 2590 10685 2620
rect 10655 2570 10660 2590
rect 10680 2570 10685 2590
rect 10655 2540 10685 2570
rect 10655 2520 10660 2540
rect 10680 2520 10685 2540
rect 10655 2490 10685 2520
rect 10655 2470 10660 2490
rect 10680 2470 10685 2490
rect 10655 2460 10685 2470
rect 10710 2640 10740 2650
rect 10710 2620 10715 2640
rect 10735 2620 10740 2640
rect 10710 2590 10740 2620
rect 10710 2570 10715 2590
rect 10735 2570 10740 2590
rect 10710 2540 10740 2570
rect 10710 2520 10715 2540
rect 10735 2520 10740 2540
rect 10710 2490 10740 2520
rect 10710 2470 10715 2490
rect 10735 2470 10740 2490
rect 10710 2460 10740 2470
rect 10765 2640 10795 2650
rect 10765 2620 10770 2640
rect 10790 2620 10795 2640
rect 10765 2590 10795 2620
rect 10765 2570 10770 2590
rect 10790 2570 10795 2590
rect 10765 2540 10795 2570
rect 10765 2520 10770 2540
rect 10790 2520 10795 2540
rect 10765 2490 10795 2520
rect 10765 2470 10770 2490
rect 10790 2470 10795 2490
rect 10765 2460 10795 2470
rect 10820 2640 10890 2650
rect 10820 2620 10825 2640
rect 10845 2620 10865 2640
rect 10885 2620 10890 2640
rect 10820 2590 10890 2620
rect 10820 2570 10825 2590
rect 10845 2570 10865 2590
rect 10885 2570 10890 2590
rect 10820 2540 10890 2570
rect 10820 2520 10825 2540
rect 10845 2520 10865 2540
rect 10885 2520 10890 2540
rect 10820 2490 10890 2520
rect 11185 2630 11255 2660
rect 11185 2610 11190 2630
rect 11210 2610 11230 2630
rect 11250 2610 11255 2630
rect 11185 2580 11255 2610
rect 11185 2560 11190 2580
rect 11210 2560 11230 2580
rect 11250 2560 11255 2580
rect 11185 2530 11255 2560
rect 11185 2510 11190 2530
rect 11210 2510 11230 2530
rect 11250 2510 11255 2530
rect 11185 2500 11255 2510
rect 11285 2880 11315 2890
rect 11285 2860 11290 2880
rect 11310 2860 11315 2880
rect 11285 2830 11315 2860
rect 11285 2810 11290 2830
rect 11310 2810 11315 2830
rect 11285 2780 11315 2810
rect 11285 2760 11290 2780
rect 11310 2760 11315 2780
rect 11285 2730 11315 2760
rect 11285 2710 11290 2730
rect 11310 2710 11315 2730
rect 11285 2680 11315 2710
rect 11285 2660 11290 2680
rect 11310 2660 11315 2680
rect 11285 2630 11315 2660
rect 11285 2610 11290 2630
rect 11310 2610 11315 2630
rect 11285 2580 11315 2610
rect 11285 2560 11290 2580
rect 11310 2560 11315 2580
rect 11285 2530 11315 2560
rect 11285 2510 11290 2530
rect 11310 2510 11315 2530
rect 11285 2500 11315 2510
rect 11345 2880 11375 2890
rect 11345 2860 11350 2880
rect 11370 2860 11375 2880
rect 11345 2830 11375 2860
rect 11345 2810 11350 2830
rect 11370 2810 11375 2830
rect 11345 2780 11375 2810
rect 11345 2760 11350 2780
rect 11370 2760 11375 2780
rect 11345 2730 11375 2760
rect 11345 2710 11350 2730
rect 11370 2710 11375 2730
rect 11345 2680 11375 2710
rect 11345 2660 11350 2680
rect 11370 2660 11375 2680
rect 11345 2630 11375 2660
rect 11345 2610 11350 2630
rect 11370 2610 11375 2630
rect 11345 2580 11375 2610
rect 11345 2560 11350 2580
rect 11370 2560 11375 2580
rect 11345 2530 11375 2560
rect 11345 2510 11350 2530
rect 11370 2510 11375 2530
rect 11345 2500 11375 2510
rect 11405 2880 11435 2890
rect 11405 2860 11410 2880
rect 11430 2860 11435 2880
rect 11405 2830 11435 2860
rect 11405 2810 11410 2830
rect 11430 2810 11435 2830
rect 11405 2780 11435 2810
rect 11405 2760 11410 2780
rect 11430 2760 11435 2780
rect 11405 2730 11435 2760
rect 11405 2710 11410 2730
rect 11430 2710 11435 2730
rect 11405 2680 11435 2710
rect 11405 2660 11410 2680
rect 11430 2660 11435 2680
rect 11405 2630 11435 2660
rect 11405 2610 11410 2630
rect 11430 2610 11435 2630
rect 11405 2580 11435 2610
rect 11405 2560 11410 2580
rect 11430 2560 11435 2580
rect 11405 2530 11435 2560
rect 11405 2510 11410 2530
rect 11430 2510 11435 2530
rect 11405 2500 11435 2510
rect 11465 2880 11495 2890
rect 11465 2860 11470 2880
rect 11490 2860 11495 2880
rect 11465 2830 11495 2860
rect 11465 2810 11470 2830
rect 11490 2810 11495 2830
rect 11465 2780 11495 2810
rect 11465 2760 11470 2780
rect 11490 2760 11495 2780
rect 11465 2730 11495 2760
rect 11465 2710 11470 2730
rect 11490 2710 11495 2730
rect 11465 2680 11495 2710
rect 11465 2660 11470 2680
rect 11490 2660 11495 2680
rect 11465 2630 11495 2660
rect 11465 2610 11470 2630
rect 11490 2610 11495 2630
rect 11465 2580 11495 2610
rect 11465 2560 11470 2580
rect 11490 2560 11495 2580
rect 11465 2530 11495 2560
rect 11465 2510 11470 2530
rect 11490 2510 11495 2530
rect 11465 2500 11495 2510
rect 11525 2880 11555 2890
rect 11525 2860 11530 2880
rect 11550 2860 11555 2880
rect 11525 2830 11555 2860
rect 11525 2810 11530 2830
rect 11550 2810 11555 2830
rect 11525 2780 11555 2810
rect 11525 2760 11530 2780
rect 11550 2760 11555 2780
rect 11525 2730 11555 2760
rect 11525 2710 11530 2730
rect 11550 2710 11555 2730
rect 11525 2680 11555 2710
rect 11525 2660 11530 2680
rect 11550 2660 11555 2680
rect 11525 2630 11555 2660
rect 11525 2610 11530 2630
rect 11550 2610 11555 2630
rect 11525 2580 11555 2610
rect 11525 2560 11530 2580
rect 11550 2560 11555 2580
rect 11525 2530 11555 2560
rect 11525 2510 11530 2530
rect 11550 2510 11555 2530
rect 11525 2500 11555 2510
rect 11585 2880 11615 2890
rect 11585 2860 11590 2880
rect 11610 2860 11615 2880
rect 11585 2830 11615 2860
rect 11585 2810 11590 2830
rect 11610 2810 11615 2830
rect 11585 2780 11615 2810
rect 11585 2760 11590 2780
rect 11610 2760 11615 2780
rect 11585 2730 11615 2760
rect 11585 2710 11590 2730
rect 11610 2710 11615 2730
rect 11585 2680 11615 2710
rect 11585 2660 11590 2680
rect 11610 2660 11615 2680
rect 11585 2630 11615 2660
rect 11585 2610 11590 2630
rect 11610 2610 11615 2630
rect 11585 2580 11615 2610
rect 11585 2560 11590 2580
rect 11610 2560 11615 2580
rect 11585 2530 11615 2560
rect 11585 2510 11590 2530
rect 11610 2510 11615 2530
rect 11585 2500 11615 2510
rect 11645 2880 11675 2890
rect 11645 2860 11650 2880
rect 11670 2860 11675 2880
rect 11645 2830 11675 2860
rect 11645 2810 11650 2830
rect 11670 2810 11675 2830
rect 11645 2780 11675 2810
rect 11645 2760 11650 2780
rect 11670 2760 11675 2780
rect 11645 2730 11675 2760
rect 11645 2710 11650 2730
rect 11670 2710 11675 2730
rect 11645 2680 11675 2710
rect 11645 2660 11650 2680
rect 11670 2660 11675 2680
rect 11645 2630 11675 2660
rect 11645 2610 11650 2630
rect 11670 2610 11675 2630
rect 11645 2580 11675 2610
rect 11645 2560 11650 2580
rect 11670 2560 11675 2580
rect 11645 2530 11675 2560
rect 11645 2510 11650 2530
rect 11670 2510 11675 2530
rect 11645 2500 11675 2510
rect 11705 2880 11735 2890
rect 11705 2860 11710 2880
rect 11730 2860 11735 2880
rect 11705 2830 11735 2860
rect 11705 2810 11710 2830
rect 11730 2810 11735 2830
rect 11705 2780 11735 2810
rect 11705 2760 11710 2780
rect 11730 2760 11735 2780
rect 11705 2730 11735 2760
rect 11705 2710 11710 2730
rect 11730 2710 11735 2730
rect 11705 2680 11735 2710
rect 11705 2660 11710 2680
rect 11730 2660 11735 2680
rect 11705 2630 11735 2660
rect 11705 2610 11710 2630
rect 11730 2610 11735 2630
rect 11705 2580 11735 2610
rect 11705 2560 11710 2580
rect 11730 2560 11735 2580
rect 11705 2530 11735 2560
rect 11705 2510 11710 2530
rect 11730 2510 11735 2530
rect 11705 2500 11735 2510
rect 11765 2880 11795 2890
rect 11765 2860 11770 2880
rect 11790 2860 11795 2880
rect 11765 2830 11795 2860
rect 11765 2810 11770 2830
rect 11790 2810 11795 2830
rect 11765 2780 11795 2810
rect 11765 2760 11770 2780
rect 11790 2760 11795 2780
rect 11765 2730 11795 2760
rect 11765 2710 11770 2730
rect 11790 2710 11795 2730
rect 11765 2680 11795 2710
rect 11765 2660 11770 2680
rect 11790 2660 11795 2680
rect 11765 2630 11795 2660
rect 11765 2610 11770 2630
rect 11790 2610 11795 2630
rect 11765 2580 11795 2610
rect 11765 2560 11770 2580
rect 11790 2560 11795 2580
rect 11765 2530 11795 2560
rect 11765 2510 11770 2530
rect 11790 2510 11795 2530
rect 11765 2500 11795 2510
rect 11825 2880 11855 2890
rect 11825 2860 11830 2880
rect 11850 2860 11855 2880
rect 11825 2830 11855 2860
rect 11825 2810 11830 2830
rect 11850 2810 11855 2830
rect 11825 2780 11855 2810
rect 11825 2760 11830 2780
rect 11850 2760 11855 2780
rect 11825 2730 11855 2760
rect 11825 2710 11830 2730
rect 11850 2710 11855 2730
rect 11825 2680 11855 2710
rect 11825 2660 11830 2680
rect 11850 2660 11855 2680
rect 11825 2630 11855 2660
rect 11825 2610 11830 2630
rect 11850 2610 11855 2630
rect 11825 2580 11855 2610
rect 11825 2560 11830 2580
rect 11850 2560 11855 2580
rect 11825 2530 11855 2560
rect 11825 2510 11830 2530
rect 11850 2510 11855 2530
rect 11825 2500 11855 2510
rect 11885 2880 11915 2890
rect 11885 2860 11890 2880
rect 11910 2860 11915 2880
rect 11885 2830 11915 2860
rect 11885 2810 11890 2830
rect 11910 2810 11915 2830
rect 11885 2780 11915 2810
rect 11885 2760 11890 2780
rect 11910 2760 11915 2780
rect 11885 2730 11915 2760
rect 11885 2710 11890 2730
rect 11910 2710 11915 2730
rect 11885 2680 11915 2710
rect 11885 2660 11890 2680
rect 11910 2660 11915 2680
rect 11885 2630 11915 2660
rect 11885 2610 11890 2630
rect 11910 2610 11915 2630
rect 11885 2580 11915 2610
rect 11885 2560 11890 2580
rect 11910 2560 11915 2580
rect 11885 2530 11915 2560
rect 11885 2510 11890 2530
rect 11910 2510 11915 2530
rect 11885 2500 11915 2510
rect 11945 2880 11975 2890
rect 11945 2860 11950 2880
rect 11970 2860 11975 2880
rect 11945 2830 11975 2860
rect 11945 2810 11950 2830
rect 11970 2810 11975 2830
rect 11945 2780 11975 2810
rect 11945 2760 11950 2780
rect 11970 2760 11975 2780
rect 11945 2730 11975 2760
rect 11945 2710 11950 2730
rect 11970 2710 11975 2730
rect 11945 2680 11975 2710
rect 11945 2660 11950 2680
rect 11970 2660 11975 2680
rect 11945 2630 11975 2660
rect 11945 2610 11950 2630
rect 11970 2610 11975 2630
rect 11945 2580 11975 2610
rect 11945 2560 11950 2580
rect 11970 2560 11975 2580
rect 11945 2530 11975 2560
rect 11945 2510 11950 2530
rect 11970 2510 11975 2530
rect 11945 2500 11975 2510
rect 12005 2880 12035 2890
rect 12005 2860 12010 2880
rect 12030 2860 12035 2880
rect 12005 2830 12035 2860
rect 12005 2810 12010 2830
rect 12030 2810 12035 2830
rect 12005 2780 12035 2810
rect 12005 2760 12010 2780
rect 12030 2760 12035 2780
rect 12005 2730 12035 2760
rect 12005 2710 12010 2730
rect 12030 2710 12035 2730
rect 12005 2680 12035 2710
rect 12005 2660 12010 2680
rect 12030 2660 12035 2680
rect 12005 2630 12035 2660
rect 12005 2610 12010 2630
rect 12030 2610 12035 2630
rect 12005 2580 12035 2610
rect 12005 2560 12010 2580
rect 12030 2560 12035 2580
rect 12005 2530 12035 2560
rect 12005 2510 12010 2530
rect 12030 2510 12035 2530
rect 12005 2500 12035 2510
rect 12065 2880 12095 2890
rect 12065 2860 12070 2880
rect 12090 2860 12095 2880
rect 12065 2830 12095 2860
rect 12065 2810 12070 2830
rect 12090 2810 12095 2830
rect 12065 2780 12095 2810
rect 12065 2760 12070 2780
rect 12090 2760 12095 2780
rect 12065 2730 12095 2760
rect 12065 2710 12070 2730
rect 12090 2710 12095 2730
rect 12065 2680 12095 2710
rect 12065 2660 12070 2680
rect 12090 2660 12095 2680
rect 12065 2630 12095 2660
rect 12065 2610 12070 2630
rect 12090 2610 12095 2630
rect 12065 2580 12095 2610
rect 12065 2560 12070 2580
rect 12090 2560 12095 2580
rect 12065 2530 12095 2560
rect 12065 2510 12070 2530
rect 12090 2510 12095 2530
rect 12065 2500 12095 2510
rect 12125 2880 12155 2890
rect 12125 2860 12130 2880
rect 12150 2860 12155 2880
rect 12125 2830 12155 2860
rect 12125 2810 12130 2830
rect 12150 2810 12155 2830
rect 12125 2780 12155 2810
rect 12125 2760 12130 2780
rect 12150 2760 12155 2780
rect 12125 2730 12155 2760
rect 12125 2710 12130 2730
rect 12150 2710 12155 2730
rect 12125 2680 12155 2710
rect 12125 2660 12130 2680
rect 12150 2660 12155 2680
rect 12125 2630 12155 2660
rect 12125 2610 12130 2630
rect 12150 2610 12155 2630
rect 12125 2580 12155 2610
rect 12125 2560 12130 2580
rect 12150 2560 12155 2580
rect 12125 2530 12155 2560
rect 12125 2510 12130 2530
rect 12150 2510 12155 2530
rect 12125 2500 12155 2510
rect 12185 2880 12215 2890
rect 12185 2860 12190 2880
rect 12210 2860 12215 2880
rect 12185 2830 12215 2860
rect 12185 2810 12190 2830
rect 12210 2810 12215 2830
rect 12185 2780 12215 2810
rect 12185 2760 12190 2780
rect 12210 2760 12215 2780
rect 12185 2730 12215 2760
rect 12185 2710 12190 2730
rect 12210 2710 12215 2730
rect 12185 2680 12215 2710
rect 12185 2660 12190 2680
rect 12210 2660 12215 2680
rect 12185 2630 12215 2660
rect 12185 2610 12190 2630
rect 12210 2610 12215 2630
rect 12185 2580 12215 2610
rect 12185 2560 12190 2580
rect 12210 2560 12215 2580
rect 12185 2530 12215 2560
rect 12185 2510 12190 2530
rect 12210 2510 12215 2530
rect 12185 2500 12215 2510
rect 12245 2880 12275 2890
rect 12245 2860 12250 2880
rect 12270 2860 12275 2880
rect 12245 2830 12275 2860
rect 12245 2810 12250 2830
rect 12270 2810 12275 2830
rect 12245 2780 12275 2810
rect 12245 2760 12250 2780
rect 12270 2760 12275 2780
rect 12245 2730 12275 2760
rect 12245 2710 12250 2730
rect 12270 2710 12275 2730
rect 12245 2680 12275 2710
rect 12245 2660 12250 2680
rect 12270 2660 12275 2680
rect 12245 2630 12275 2660
rect 12245 2610 12250 2630
rect 12270 2610 12275 2630
rect 12245 2580 12275 2610
rect 12245 2560 12250 2580
rect 12270 2560 12275 2580
rect 12245 2530 12275 2560
rect 12245 2510 12250 2530
rect 12270 2510 12275 2530
rect 12245 2500 12275 2510
rect 12305 2880 12335 2890
rect 12305 2860 12310 2880
rect 12330 2860 12335 2880
rect 12305 2830 12335 2860
rect 12305 2810 12310 2830
rect 12330 2810 12335 2830
rect 12305 2780 12335 2810
rect 12305 2760 12310 2780
rect 12330 2760 12335 2780
rect 12305 2730 12335 2760
rect 12305 2710 12310 2730
rect 12330 2710 12335 2730
rect 12305 2680 12335 2710
rect 12305 2660 12310 2680
rect 12330 2660 12335 2680
rect 12305 2630 12335 2660
rect 12305 2610 12310 2630
rect 12330 2610 12335 2630
rect 12305 2580 12335 2610
rect 12305 2560 12310 2580
rect 12330 2560 12335 2580
rect 12305 2530 12335 2560
rect 12305 2510 12310 2530
rect 12330 2510 12335 2530
rect 12305 2500 12335 2510
rect 12365 2880 12395 2890
rect 12365 2860 12370 2880
rect 12390 2860 12395 2880
rect 12365 2830 12395 2860
rect 12365 2810 12370 2830
rect 12390 2810 12395 2830
rect 12365 2780 12395 2810
rect 12365 2760 12370 2780
rect 12390 2760 12395 2780
rect 12365 2730 12395 2760
rect 12365 2710 12370 2730
rect 12390 2710 12395 2730
rect 12365 2680 12395 2710
rect 12365 2660 12370 2680
rect 12390 2660 12395 2680
rect 12365 2630 12395 2660
rect 12365 2610 12370 2630
rect 12390 2610 12395 2630
rect 12365 2580 12395 2610
rect 12365 2560 12370 2580
rect 12390 2560 12395 2580
rect 12365 2530 12395 2560
rect 12365 2510 12370 2530
rect 12390 2510 12395 2530
rect 12365 2500 12395 2510
rect 12425 2880 12455 2890
rect 12425 2860 12430 2880
rect 12450 2860 12455 2880
rect 12425 2830 12455 2860
rect 12425 2810 12430 2830
rect 12450 2810 12455 2830
rect 12425 2780 12455 2810
rect 12425 2760 12430 2780
rect 12450 2760 12455 2780
rect 12425 2730 12455 2760
rect 12425 2710 12430 2730
rect 12450 2710 12455 2730
rect 12425 2680 12455 2710
rect 12425 2660 12430 2680
rect 12450 2660 12455 2680
rect 12425 2630 12455 2660
rect 12425 2610 12430 2630
rect 12450 2610 12455 2630
rect 12425 2580 12455 2610
rect 12425 2560 12430 2580
rect 12450 2560 12455 2580
rect 12425 2530 12455 2560
rect 12425 2510 12430 2530
rect 12450 2510 12455 2530
rect 12425 2500 12455 2510
rect 12485 2880 12515 2890
rect 12485 2860 12490 2880
rect 12510 2860 12515 2880
rect 12485 2830 12515 2860
rect 12485 2810 12490 2830
rect 12510 2810 12515 2830
rect 12485 2780 12515 2810
rect 12485 2760 12490 2780
rect 12510 2760 12515 2780
rect 12485 2730 12515 2760
rect 12485 2710 12490 2730
rect 12510 2710 12515 2730
rect 12485 2680 12515 2710
rect 12485 2660 12490 2680
rect 12510 2660 12515 2680
rect 12485 2630 12515 2660
rect 12485 2610 12490 2630
rect 12510 2610 12515 2630
rect 12485 2580 12515 2610
rect 12485 2560 12490 2580
rect 12510 2560 12515 2580
rect 12485 2530 12515 2560
rect 12485 2510 12490 2530
rect 12510 2510 12515 2530
rect 12485 2500 12515 2510
rect 12545 2880 12615 2890
rect 12545 2860 12550 2880
rect 12570 2860 12590 2880
rect 12610 2860 12615 2880
rect 12545 2830 12615 2860
rect 12545 2810 12550 2830
rect 12570 2810 12590 2830
rect 12610 2810 12615 2830
rect 12545 2780 12615 2810
rect 12545 2760 12550 2780
rect 12570 2760 12590 2780
rect 12610 2760 12615 2780
rect 12545 2730 12615 2760
rect 12545 2710 12550 2730
rect 12570 2710 12590 2730
rect 12610 2710 12615 2730
rect 26185 2880 26255 2890
rect 26185 2860 26190 2880
rect 26210 2860 26230 2880
rect 26250 2860 26255 2880
rect 26185 2830 26255 2860
rect 26185 2810 26190 2830
rect 26210 2810 26230 2830
rect 26250 2810 26255 2830
rect 26185 2780 26255 2810
rect 26185 2760 26190 2780
rect 26210 2760 26230 2780
rect 26250 2760 26255 2780
rect 26185 2730 26255 2760
rect 26185 2710 26190 2730
rect 26210 2710 26230 2730
rect 26250 2710 26255 2730
rect 12545 2680 12615 2710
rect 12545 2660 12550 2680
rect 12570 2660 12590 2680
rect 12610 2660 12615 2680
rect 13000 2700 13040 2710
rect 13000 2680 13010 2700
rect 13030 2680 13040 2700
rect 13000 2670 13040 2680
rect 13110 2700 13150 2710
rect 13110 2680 13120 2700
rect 13140 2680 13150 2700
rect 13110 2670 13150 2680
rect 13220 2700 13260 2710
rect 13220 2680 13230 2700
rect 13250 2680 13260 2700
rect 13220 2670 13260 2680
rect 13330 2700 13370 2710
rect 13330 2680 13340 2700
rect 13360 2680 13370 2700
rect 13330 2670 13370 2680
rect 13440 2700 13480 2710
rect 13440 2680 13450 2700
rect 13470 2680 13480 2700
rect 13440 2670 13480 2680
rect 13550 2700 13590 2710
rect 13550 2680 13560 2700
rect 13580 2680 13590 2700
rect 13550 2670 13590 2680
rect 26185 2680 26255 2710
rect 12545 2630 12615 2660
rect 13010 2650 13030 2670
rect 13120 2650 13140 2670
rect 13230 2650 13250 2670
rect 13340 2650 13360 2670
rect 13450 2650 13470 2670
rect 13560 2650 13580 2670
rect 24735 2665 24775 2675
rect 12545 2610 12550 2630
rect 12570 2610 12590 2630
rect 12610 2610 12615 2630
rect 12545 2580 12615 2610
rect 12545 2560 12550 2580
rect 12570 2560 12590 2580
rect 12610 2560 12615 2580
rect 12545 2530 12615 2560
rect 12545 2510 12550 2530
rect 12570 2510 12590 2530
rect 12610 2510 12615 2530
rect 12545 2500 12615 2510
rect 12910 2640 12980 2650
rect 12910 2620 12915 2640
rect 12935 2620 12955 2640
rect 12975 2620 12980 2640
rect 12910 2590 12980 2620
rect 12910 2570 12915 2590
rect 12935 2570 12955 2590
rect 12975 2570 12980 2590
rect 12910 2540 12980 2570
rect 12910 2520 12915 2540
rect 12935 2520 12955 2540
rect 12975 2520 12980 2540
rect 10820 2470 10825 2490
rect 10845 2470 10865 2490
rect 10885 2470 10890 2490
rect 11290 2480 11310 2500
rect 11410 2480 11430 2500
rect 11530 2480 11550 2500
rect 11650 2480 11670 2500
rect 11770 2480 11790 2500
rect 11890 2480 11910 2500
rect 12010 2480 12030 2500
rect 12130 2480 12150 2500
rect 12250 2480 12270 2500
rect 12370 2480 12390 2500
rect 12490 2480 12510 2500
rect 12910 2490 12980 2520
rect 10820 2460 10890 2470
rect 11280 2470 11320 2480
rect 10125 2440 10145 2460
rect 10275 2440 10295 2460
rect 10385 2440 10405 2460
rect 10495 2440 10515 2460
rect 10605 2440 10625 2460
rect 10715 2440 10735 2460
rect 10865 2440 10885 2460
rect 11280 2450 11290 2470
rect 11310 2450 11320 2470
rect 11280 2440 11320 2450
rect 11400 2470 11440 2480
rect 11400 2450 11410 2470
rect 11430 2450 11440 2470
rect 11400 2440 11440 2450
rect 11520 2470 11560 2480
rect 11520 2450 11530 2470
rect 11550 2450 11560 2470
rect 11520 2440 11560 2450
rect 11640 2470 11680 2480
rect 11640 2450 11650 2470
rect 11670 2450 11680 2470
rect 11640 2440 11680 2450
rect 11760 2470 11800 2480
rect 11760 2450 11770 2470
rect 11790 2450 11800 2470
rect 11760 2440 11800 2450
rect 11823 2470 11857 2480
rect 11823 2450 11831 2470
rect 11849 2450 11857 2470
rect 11823 2440 11857 2450
rect 11880 2470 11920 2480
rect 11880 2450 11890 2470
rect 11910 2450 11920 2470
rect 11880 2440 11920 2450
rect 12000 2470 12040 2480
rect 12000 2450 12010 2470
rect 12030 2450 12040 2470
rect 12000 2440 12040 2450
rect 12120 2470 12160 2480
rect 12120 2450 12130 2470
rect 12150 2450 12160 2470
rect 12120 2440 12160 2450
rect 12240 2470 12280 2480
rect 12240 2450 12250 2470
rect 12270 2450 12280 2470
rect 12240 2440 12280 2450
rect 12360 2470 12400 2480
rect 12360 2450 12370 2470
rect 12390 2450 12400 2470
rect 12360 2440 12400 2450
rect 12480 2470 12520 2480
rect 12480 2450 12490 2470
rect 12510 2450 12520 2470
rect 12910 2470 12915 2490
rect 12935 2470 12955 2490
rect 12975 2470 12980 2490
rect 12910 2460 12980 2470
rect 13005 2640 13035 2650
rect 13005 2620 13010 2640
rect 13030 2620 13035 2640
rect 13005 2590 13035 2620
rect 13005 2570 13010 2590
rect 13030 2570 13035 2590
rect 13005 2540 13035 2570
rect 13005 2520 13010 2540
rect 13030 2520 13035 2540
rect 13005 2490 13035 2520
rect 13005 2470 13010 2490
rect 13030 2470 13035 2490
rect 13005 2460 13035 2470
rect 13060 2640 13090 2650
rect 13060 2620 13065 2640
rect 13085 2620 13090 2640
rect 13060 2590 13090 2620
rect 13060 2570 13065 2590
rect 13085 2570 13090 2590
rect 13060 2540 13090 2570
rect 13060 2520 13065 2540
rect 13085 2520 13090 2540
rect 13060 2490 13090 2520
rect 13060 2470 13065 2490
rect 13085 2470 13090 2490
rect 13060 2460 13090 2470
rect 13115 2640 13145 2650
rect 13115 2620 13120 2640
rect 13140 2620 13145 2640
rect 13115 2590 13145 2620
rect 13115 2570 13120 2590
rect 13140 2570 13145 2590
rect 13115 2540 13145 2570
rect 13115 2520 13120 2540
rect 13140 2520 13145 2540
rect 13115 2490 13145 2520
rect 13115 2470 13120 2490
rect 13140 2470 13145 2490
rect 13115 2460 13145 2470
rect 13170 2640 13200 2650
rect 13170 2620 13175 2640
rect 13195 2620 13200 2640
rect 13170 2590 13200 2620
rect 13170 2570 13175 2590
rect 13195 2570 13200 2590
rect 13170 2540 13200 2570
rect 13170 2520 13175 2540
rect 13195 2520 13200 2540
rect 13170 2490 13200 2520
rect 13170 2470 13175 2490
rect 13195 2470 13200 2490
rect 13170 2460 13200 2470
rect 13225 2640 13255 2650
rect 13225 2620 13230 2640
rect 13250 2620 13255 2640
rect 13225 2590 13255 2620
rect 13225 2570 13230 2590
rect 13250 2570 13255 2590
rect 13225 2540 13255 2570
rect 13225 2520 13230 2540
rect 13250 2520 13255 2540
rect 13225 2490 13255 2520
rect 13225 2470 13230 2490
rect 13250 2470 13255 2490
rect 13225 2460 13255 2470
rect 13280 2640 13310 2650
rect 13280 2620 13285 2640
rect 13305 2620 13310 2640
rect 13280 2590 13310 2620
rect 13280 2570 13285 2590
rect 13305 2570 13310 2590
rect 13280 2540 13310 2570
rect 13280 2520 13285 2540
rect 13305 2520 13310 2540
rect 13280 2490 13310 2520
rect 13280 2470 13285 2490
rect 13305 2470 13310 2490
rect 13280 2460 13310 2470
rect 13335 2640 13365 2650
rect 13335 2620 13340 2640
rect 13360 2620 13365 2640
rect 13335 2590 13365 2620
rect 13335 2570 13340 2590
rect 13360 2570 13365 2590
rect 13335 2540 13365 2570
rect 13335 2520 13340 2540
rect 13360 2520 13365 2540
rect 13335 2490 13365 2520
rect 13335 2470 13340 2490
rect 13360 2470 13365 2490
rect 13335 2460 13365 2470
rect 13390 2640 13420 2650
rect 13390 2620 13395 2640
rect 13415 2620 13420 2640
rect 13390 2590 13420 2620
rect 13390 2570 13395 2590
rect 13415 2570 13420 2590
rect 13390 2540 13420 2570
rect 13390 2520 13395 2540
rect 13415 2520 13420 2540
rect 13390 2490 13420 2520
rect 13390 2470 13395 2490
rect 13415 2470 13420 2490
rect 13390 2460 13420 2470
rect 13445 2640 13475 2650
rect 13445 2620 13450 2640
rect 13470 2620 13475 2640
rect 13445 2590 13475 2620
rect 13445 2570 13450 2590
rect 13470 2570 13475 2590
rect 13445 2540 13475 2570
rect 13445 2520 13450 2540
rect 13470 2520 13475 2540
rect 13445 2490 13475 2520
rect 13445 2470 13450 2490
rect 13470 2470 13475 2490
rect 13445 2460 13475 2470
rect 13500 2640 13530 2650
rect 13500 2620 13505 2640
rect 13525 2620 13530 2640
rect 13500 2590 13530 2620
rect 13500 2570 13505 2590
rect 13525 2570 13530 2590
rect 13500 2540 13530 2570
rect 13500 2520 13505 2540
rect 13525 2520 13530 2540
rect 13500 2490 13530 2520
rect 13500 2470 13505 2490
rect 13525 2470 13530 2490
rect 13500 2460 13530 2470
rect 13555 2640 13585 2650
rect 13555 2620 13560 2640
rect 13580 2620 13585 2640
rect 13555 2590 13585 2620
rect 13555 2570 13560 2590
rect 13580 2570 13585 2590
rect 13555 2540 13585 2570
rect 13555 2520 13560 2540
rect 13580 2520 13585 2540
rect 13555 2490 13585 2520
rect 13555 2470 13560 2490
rect 13580 2470 13585 2490
rect 13555 2460 13585 2470
rect 13610 2640 13680 2650
rect 13610 2620 13615 2640
rect 13635 2620 13655 2640
rect 13675 2620 13680 2640
rect 13610 2590 13680 2620
rect 13610 2570 13615 2590
rect 13635 2570 13655 2590
rect 13675 2570 13680 2590
rect 13610 2540 13680 2570
rect 13610 2520 13615 2540
rect 13635 2520 13655 2540
rect 13675 2520 13680 2540
rect 13610 2490 13680 2520
rect 13610 2470 13615 2490
rect 13635 2470 13655 2490
rect 13675 2470 13680 2490
rect 13610 2460 13680 2470
rect 13795 2645 14010 2665
rect 13795 2625 13830 2645
rect 13975 2625 14010 2645
rect 24735 2645 24745 2665
rect 24765 2645 24775 2665
rect 24735 2635 24775 2645
rect 24845 2665 24885 2675
rect 24845 2645 24855 2665
rect 24875 2645 24885 2665
rect 24845 2635 24885 2645
rect 24955 2665 24995 2675
rect 24955 2645 24965 2665
rect 24985 2645 24995 2665
rect 24955 2635 24995 2645
rect 25065 2665 25105 2675
rect 25065 2645 25075 2665
rect 25095 2645 25105 2665
rect 25065 2635 25105 2645
rect 25175 2665 25215 2675
rect 25175 2645 25185 2665
rect 25205 2645 25215 2665
rect 25175 2635 25215 2645
rect 25285 2665 25325 2675
rect 25285 2645 25295 2665
rect 25315 2645 25325 2665
rect 25285 2635 25325 2645
rect 25395 2665 25435 2675
rect 25395 2645 25405 2665
rect 25425 2645 25435 2665
rect 25395 2635 25435 2645
rect 25505 2665 25545 2675
rect 25505 2645 25515 2665
rect 25535 2645 25545 2665
rect 25505 2635 25545 2645
rect 25615 2665 25655 2675
rect 25615 2645 25625 2665
rect 25645 2645 25655 2665
rect 25615 2635 25655 2645
rect 25725 2665 25765 2675
rect 25725 2645 25735 2665
rect 25755 2645 25765 2665
rect 25725 2635 25765 2645
rect 25835 2665 25875 2675
rect 25835 2645 25845 2665
rect 25865 2645 25875 2665
rect 25835 2635 25875 2645
rect 26185 2660 26190 2680
rect 26210 2660 26230 2680
rect 26250 2660 26255 2680
rect 12480 2440 12520 2450
rect 12915 2440 12935 2460
rect 13065 2440 13085 2460
rect 13175 2440 13195 2460
rect 13285 2440 13305 2460
rect 13395 2440 13415 2460
rect 13505 2440 13525 2460
rect 13655 2440 13675 2460
rect 10115 2430 10155 2440
rect 10115 2410 10125 2430
rect 10145 2410 10155 2430
rect 3275 2385 3295 2405
rect 3455 2385 3475 2405
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2370 3395 2380
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 2625 2315 2655 2345
rect 3355 2340 3395 2350
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3635 2340 3655 2405
rect 3815 2385 3835 2405
rect 3995 2385 4015 2405
rect 4175 2385 4195 2405
rect 3805 2375 3845 2385
rect 3805 2355 3815 2375
rect 3835 2355 3845 2375
rect 3805 2345 3845 2355
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2375 4205 2385
rect 4165 2355 4175 2375
rect 4195 2355 4205 2375
rect 4165 2345 4205 2355
rect 4355 2340 4375 2405
rect 4535 2385 4555 2405
rect 4715 2385 4735 2405
rect 10115 2400 10155 2410
rect 10265 2430 10305 2440
rect 10265 2410 10275 2430
rect 10295 2410 10305 2430
rect 10265 2400 10305 2410
rect 10375 2430 10415 2440
rect 10375 2410 10385 2430
rect 10405 2410 10415 2430
rect 10375 2400 10415 2410
rect 10485 2430 10525 2440
rect 10485 2410 10495 2430
rect 10515 2410 10525 2430
rect 10485 2400 10525 2410
rect 10595 2430 10635 2440
rect 10595 2410 10605 2430
rect 10625 2410 10635 2430
rect 10595 2400 10635 2410
rect 10705 2430 10745 2440
rect 10705 2410 10715 2430
rect 10735 2410 10745 2430
rect 10705 2400 10745 2410
rect 10855 2430 10895 2440
rect 10855 2410 10865 2430
rect 10885 2410 10895 2430
rect 10855 2400 10895 2410
rect 12905 2430 12945 2440
rect 12905 2410 12915 2430
rect 12935 2410 12945 2430
rect 12905 2400 12945 2410
rect 13055 2430 13095 2440
rect 13055 2410 13065 2430
rect 13085 2410 13095 2430
rect 13055 2400 13095 2410
rect 13165 2430 13205 2440
rect 13165 2410 13175 2430
rect 13195 2410 13205 2430
rect 13165 2400 13205 2410
rect 13275 2430 13315 2440
rect 13275 2410 13285 2430
rect 13305 2410 13315 2430
rect 13275 2400 13315 2410
rect 13385 2430 13425 2440
rect 13385 2410 13395 2430
rect 13415 2410 13425 2430
rect 13385 2400 13425 2410
rect 13495 2430 13535 2440
rect 13495 2410 13505 2430
rect 13525 2410 13535 2430
rect 13495 2400 13535 2410
rect 13645 2430 13685 2440
rect 13645 2410 13655 2430
rect 13675 2410 13685 2430
rect 13645 2400 13685 2410
rect 13890 2575 13915 2625
rect 24745 2615 24765 2635
rect 24855 2615 24875 2635
rect 24965 2615 24985 2635
rect 25075 2615 25095 2635
rect 25185 2615 25205 2635
rect 25295 2615 25315 2635
rect 25405 2615 25425 2635
rect 25515 2615 25535 2635
rect 25625 2615 25645 2635
rect 25735 2615 25755 2635
rect 25845 2615 25865 2635
rect 26185 2630 26255 2660
rect 24645 2605 24715 2615
rect 24645 2585 24650 2605
rect 24670 2585 24690 2605
rect 24710 2585 24715 2605
rect 24645 2555 24715 2585
rect 24645 2535 24650 2555
rect 24670 2535 24690 2555
rect 24710 2535 24715 2555
rect 24645 2525 24715 2535
rect 24740 2605 24770 2615
rect 24740 2585 24745 2605
rect 24765 2585 24770 2605
rect 24740 2555 24770 2585
rect 24740 2535 24745 2555
rect 24765 2535 24770 2555
rect 24740 2525 24770 2535
rect 24795 2605 24825 2615
rect 24795 2585 24800 2605
rect 24820 2585 24825 2605
rect 24795 2555 24825 2585
rect 24795 2535 24800 2555
rect 24820 2535 24825 2555
rect 24795 2525 24825 2535
rect 24850 2605 24880 2615
rect 24850 2585 24855 2605
rect 24875 2585 24880 2605
rect 24850 2555 24880 2585
rect 24850 2535 24855 2555
rect 24875 2535 24880 2555
rect 24850 2525 24880 2535
rect 24905 2605 24935 2615
rect 24905 2585 24910 2605
rect 24930 2585 24935 2605
rect 24905 2555 24935 2585
rect 24905 2535 24910 2555
rect 24930 2535 24935 2555
rect 24905 2525 24935 2535
rect 24960 2605 24990 2615
rect 24960 2585 24965 2605
rect 24985 2585 24990 2605
rect 24960 2555 24990 2585
rect 24960 2535 24965 2555
rect 24985 2535 24990 2555
rect 24960 2525 24990 2535
rect 25015 2605 25045 2615
rect 25015 2585 25020 2605
rect 25040 2585 25045 2605
rect 25015 2555 25045 2585
rect 25015 2535 25020 2555
rect 25040 2535 25045 2555
rect 25015 2525 25045 2535
rect 25070 2605 25100 2615
rect 25070 2585 25075 2605
rect 25095 2585 25100 2605
rect 25070 2555 25100 2585
rect 25070 2535 25075 2555
rect 25095 2535 25100 2555
rect 25070 2525 25100 2535
rect 25125 2605 25155 2615
rect 25125 2585 25130 2605
rect 25150 2585 25155 2605
rect 25125 2555 25155 2585
rect 25125 2535 25130 2555
rect 25150 2535 25155 2555
rect 25125 2525 25155 2535
rect 25180 2605 25210 2615
rect 25180 2585 25185 2605
rect 25205 2585 25210 2605
rect 25180 2555 25210 2585
rect 25180 2535 25185 2555
rect 25205 2535 25210 2555
rect 25180 2525 25210 2535
rect 25235 2605 25265 2615
rect 25235 2585 25240 2605
rect 25260 2585 25265 2605
rect 25235 2555 25265 2585
rect 25235 2535 25240 2555
rect 25260 2535 25265 2555
rect 25235 2525 25265 2535
rect 25290 2605 25320 2615
rect 25290 2585 25295 2605
rect 25315 2585 25320 2605
rect 25290 2555 25320 2585
rect 25290 2535 25295 2555
rect 25315 2535 25320 2555
rect 25290 2525 25320 2535
rect 25345 2605 25375 2615
rect 25345 2585 25350 2605
rect 25370 2585 25375 2605
rect 25345 2555 25375 2585
rect 25345 2535 25350 2555
rect 25370 2535 25375 2555
rect 25345 2525 25375 2535
rect 25400 2605 25430 2615
rect 25400 2585 25405 2605
rect 25425 2585 25430 2605
rect 25400 2555 25430 2585
rect 25400 2535 25405 2555
rect 25425 2535 25430 2555
rect 25400 2525 25430 2535
rect 25455 2605 25485 2615
rect 25455 2585 25460 2605
rect 25480 2585 25485 2605
rect 25455 2555 25485 2585
rect 25455 2535 25460 2555
rect 25480 2535 25485 2555
rect 25455 2525 25485 2535
rect 25510 2605 25540 2615
rect 25510 2585 25515 2605
rect 25535 2585 25540 2605
rect 25510 2555 25540 2585
rect 25510 2535 25515 2555
rect 25535 2535 25540 2555
rect 25510 2525 25540 2535
rect 25565 2605 25595 2615
rect 25565 2585 25570 2605
rect 25590 2585 25595 2605
rect 25565 2555 25595 2585
rect 25565 2535 25570 2555
rect 25590 2535 25595 2555
rect 25565 2525 25595 2535
rect 25620 2605 25650 2615
rect 25620 2585 25625 2605
rect 25645 2585 25650 2605
rect 25620 2555 25650 2585
rect 25620 2535 25625 2555
rect 25645 2535 25650 2555
rect 25620 2525 25650 2535
rect 25675 2605 25705 2615
rect 25675 2585 25680 2605
rect 25700 2585 25705 2605
rect 25675 2555 25705 2585
rect 25675 2535 25680 2555
rect 25700 2535 25705 2555
rect 25675 2525 25705 2535
rect 25730 2605 25760 2615
rect 25730 2585 25735 2605
rect 25755 2585 25760 2605
rect 25730 2555 25760 2585
rect 25730 2535 25735 2555
rect 25755 2535 25760 2555
rect 25730 2525 25760 2535
rect 25785 2605 25815 2615
rect 25785 2585 25790 2605
rect 25810 2585 25815 2605
rect 25785 2555 25815 2585
rect 25785 2535 25790 2555
rect 25810 2535 25815 2555
rect 25785 2525 25815 2535
rect 25840 2605 25870 2615
rect 25840 2585 25845 2605
rect 25865 2585 25870 2605
rect 25840 2555 25870 2585
rect 25840 2535 25845 2555
rect 25865 2535 25870 2555
rect 25840 2525 25870 2535
rect 25895 2605 25965 2615
rect 25895 2585 25900 2605
rect 25920 2585 25940 2605
rect 25960 2585 25965 2605
rect 25895 2555 25965 2585
rect 25895 2535 25900 2555
rect 25920 2535 25940 2555
rect 25960 2535 25965 2555
rect 25895 2525 25965 2535
rect 26185 2610 26190 2630
rect 26210 2610 26230 2630
rect 26250 2610 26255 2630
rect 26185 2580 26255 2610
rect 26185 2560 26190 2580
rect 26210 2560 26230 2580
rect 26250 2560 26255 2580
rect 26185 2530 26255 2560
rect 24650 2505 24670 2525
rect 24800 2505 24820 2525
rect 24910 2505 24930 2525
rect 25020 2505 25040 2525
rect 25130 2505 25150 2525
rect 25240 2505 25260 2525
rect 25350 2505 25370 2525
rect 25460 2505 25480 2525
rect 25570 2505 25590 2525
rect 25680 2505 25700 2525
rect 25790 2505 25810 2525
rect 25940 2505 25960 2525
rect 26185 2510 26190 2530
rect 26210 2510 26230 2530
rect 26250 2510 26255 2530
rect 24640 2495 24680 2505
rect 24640 2475 24650 2495
rect 24670 2475 24680 2495
rect 24640 2465 24680 2475
rect 24790 2495 24830 2505
rect 24790 2475 24800 2495
rect 24820 2475 24830 2495
rect 24790 2465 24830 2475
rect 24900 2495 24940 2505
rect 24900 2475 24910 2495
rect 24930 2475 24940 2495
rect 24900 2465 24940 2475
rect 25010 2495 25050 2505
rect 25010 2475 25020 2495
rect 25040 2475 25050 2495
rect 25010 2465 25050 2475
rect 25120 2495 25160 2505
rect 25120 2475 25130 2495
rect 25150 2475 25160 2495
rect 25120 2465 25160 2475
rect 25230 2495 25270 2505
rect 25230 2475 25240 2495
rect 25260 2475 25270 2495
rect 25230 2465 25270 2475
rect 25340 2495 25380 2505
rect 25340 2475 25350 2495
rect 25370 2475 25380 2495
rect 25340 2465 25380 2475
rect 25450 2495 25490 2505
rect 25450 2475 25460 2495
rect 25480 2475 25490 2495
rect 25450 2465 25490 2475
rect 25560 2495 25600 2505
rect 25560 2475 25570 2495
rect 25590 2475 25600 2495
rect 25560 2465 25600 2475
rect 25670 2495 25710 2505
rect 25670 2475 25680 2495
rect 25700 2475 25710 2495
rect 25670 2465 25710 2475
rect 25780 2495 25820 2505
rect 25780 2475 25790 2495
rect 25810 2475 25820 2495
rect 25780 2465 25820 2475
rect 25930 2495 25970 2505
rect 26185 2500 26255 2510
rect 26285 2880 26315 2890
rect 26285 2860 26290 2880
rect 26310 2860 26315 2880
rect 26285 2830 26315 2860
rect 26285 2810 26290 2830
rect 26310 2810 26315 2830
rect 26285 2780 26315 2810
rect 26285 2760 26290 2780
rect 26310 2760 26315 2780
rect 26285 2730 26315 2760
rect 26285 2710 26290 2730
rect 26310 2710 26315 2730
rect 26285 2680 26315 2710
rect 26285 2660 26290 2680
rect 26310 2660 26315 2680
rect 26285 2630 26315 2660
rect 26285 2610 26290 2630
rect 26310 2610 26315 2630
rect 26285 2580 26315 2610
rect 26285 2560 26290 2580
rect 26310 2560 26315 2580
rect 26285 2530 26315 2560
rect 26285 2510 26290 2530
rect 26310 2510 26315 2530
rect 26285 2500 26315 2510
rect 26345 2880 26375 2890
rect 26345 2860 26350 2880
rect 26370 2860 26375 2880
rect 26345 2830 26375 2860
rect 26345 2810 26350 2830
rect 26370 2810 26375 2830
rect 26345 2780 26375 2810
rect 26345 2760 26350 2780
rect 26370 2760 26375 2780
rect 26345 2730 26375 2760
rect 26345 2710 26350 2730
rect 26370 2710 26375 2730
rect 26345 2680 26375 2710
rect 26345 2660 26350 2680
rect 26370 2660 26375 2680
rect 26345 2630 26375 2660
rect 26345 2610 26350 2630
rect 26370 2610 26375 2630
rect 26345 2580 26375 2610
rect 26345 2560 26350 2580
rect 26370 2560 26375 2580
rect 26345 2530 26375 2560
rect 26345 2510 26350 2530
rect 26370 2510 26375 2530
rect 26345 2500 26375 2510
rect 26405 2880 26435 2890
rect 26405 2860 26410 2880
rect 26430 2860 26435 2880
rect 26405 2830 26435 2860
rect 26405 2810 26410 2830
rect 26430 2810 26435 2830
rect 26405 2780 26435 2810
rect 26405 2760 26410 2780
rect 26430 2760 26435 2780
rect 26405 2730 26435 2760
rect 26405 2710 26410 2730
rect 26430 2710 26435 2730
rect 26405 2680 26435 2710
rect 26405 2660 26410 2680
rect 26430 2660 26435 2680
rect 26405 2630 26435 2660
rect 26405 2610 26410 2630
rect 26430 2610 26435 2630
rect 26405 2580 26435 2610
rect 26405 2560 26410 2580
rect 26430 2560 26435 2580
rect 26405 2530 26435 2560
rect 26405 2510 26410 2530
rect 26430 2510 26435 2530
rect 26405 2500 26435 2510
rect 26465 2880 26495 2890
rect 26465 2860 26470 2880
rect 26490 2860 26495 2880
rect 26465 2830 26495 2860
rect 26465 2810 26470 2830
rect 26490 2810 26495 2830
rect 26465 2780 26495 2810
rect 26465 2760 26470 2780
rect 26490 2760 26495 2780
rect 26465 2730 26495 2760
rect 26465 2710 26470 2730
rect 26490 2710 26495 2730
rect 26465 2680 26495 2710
rect 26465 2660 26470 2680
rect 26490 2660 26495 2680
rect 26465 2630 26495 2660
rect 26465 2610 26470 2630
rect 26490 2610 26495 2630
rect 26465 2580 26495 2610
rect 26465 2560 26470 2580
rect 26490 2560 26495 2580
rect 26465 2530 26495 2560
rect 26465 2510 26470 2530
rect 26490 2510 26495 2530
rect 26465 2500 26495 2510
rect 26525 2880 26555 2890
rect 26525 2860 26530 2880
rect 26550 2860 26555 2880
rect 26525 2830 26555 2860
rect 26525 2810 26530 2830
rect 26550 2810 26555 2830
rect 26525 2780 26555 2810
rect 26525 2760 26530 2780
rect 26550 2760 26555 2780
rect 26525 2730 26555 2760
rect 26525 2710 26530 2730
rect 26550 2710 26555 2730
rect 26525 2680 26555 2710
rect 26525 2660 26530 2680
rect 26550 2660 26555 2680
rect 26525 2630 26555 2660
rect 26525 2610 26530 2630
rect 26550 2610 26555 2630
rect 26525 2580 26555 2610
rect 26525 2560 26530 2580
rect 26550 2560 26555 2580
rect 26525 2530 26555 2560
rect 26525 2510 26530 2530
rect 26550 2510 26555 2530
rect 26525 2500 26555 2510
rect 26585 2880 26615 2890
rect 26585 2860 26590 2880
rect 26610 2860 26615 2880
rect 26585 2830 26615 2860
rect 26585 2810 26590 2830
rect 26610 2810 26615 2830
rect 26585 2780 26615 2810
rect 26585 2760 26590 2780
rect 26610 2760 26615 2780
rect 26585 2730 26615 2760
rect 26585 2710 26590 2730
rect 26610 2710 26615 2730
rect 26585 2680 26615 2710
rect 26585 2660 26590 2680
rect 26610 2660 26615 2680
rect 26585 2630 26615 2660
rect 26585 2610 26590 2630
rect 26610 2610 26615 2630
rect 26585 2580 26615 2610
rect 26585 2560 26590 2580
rect 26610 2560 26615 2580
rect 26585 2530 26615 2560
rect 26585 2510 26590 2530
rect 26610 2510 26615 2530
rect 26585 2500 26615 2510
rect 26645 2880 26675 2890
rect 26645 2860 26650 2880
rect 26670 2860 26675 2880
rect 26645 2830 26675 2860
rect 26645 2810 26650 2830
rect 26670 2810 26675 2830
rect 26645 2780 26675 2810
rect 26645 2760 26650 2780
rect 26670 2760 26675 2780
rect 26645 2730 26675 2760
rect 26645 2710 26650 2730
rect 26670 2710 26675 2730
rect 26645 2680 26675 2710
rect 26645 2660 26650 2680
rect 26670 2660 26675 2680
rect 26645 2630 26675 2660
rect 26645 2610 26650 2630
rect 26670 2610 26675 2630
rect 26645 2580 26675 2610
rect 26645 2560 26650 2580
rect 26670 2560 26675 2580
rect 26645 2530 26675 2560
rect 26645 2510 26650 2530
rect 26670 2510 26675 2530
rect 26645 2500 26675 2510
rect 26705 2880 26735 2890
rect 26705 2860 26710 2880
rect 26730 2860 26735 2880
rect 26705 2830 26735 2860
rect 26705 2810 26710 2830
rect 26730 2810 26735 2830
rect 26705 2780 26735 2810
rect 26705 2760 26710 2780
rect 26730 2760 26735 2780
rect 26705 2730 26735 2760
rect 26705 2710 26710 2730
rect 26730 2710 26735 2730
rect 26705 2680 26735 2710
rect 26705 2660 26710 2680
rect 26730 2660 26735 2680
rect 26705 2630 26735 2660
rect 26705 2610 26710 2630
rect 26730 2610 26735 2630
rect 26705 2580 26735 2610
rect 26705 2560 26710 2580
rect 26730 2560 26735 2580
rect 26705 2530 26735 2560
rect 26705 2510 26710 2530
rect 26730 2510 26735 2530
rect 26705 2500 26735 2510
rect 26765 2880 26795 2890
rect 26765 2860 26770 2880
rect 26790 2860 26795 2880
rect 26765 2830 26795 2860
rect 26765 2810 26770 2830
rect 26790 2810 26795 2830
rect 26765 2780 26795 2810
rect 26765 2760 26770 2780
rect 26790 2760 26795 2780
rect 26765 2730 26795 2760
rect 26765 2710 26770 2730
rect 26790 2710 26795 2730
rect 26765 2680 26795 2710
rect 26765 2660 26770 2680
rect 26790 2660 26795 2680
rect 26765 2630 26795 2660
rect 26765 2610 26770 2630
rect 26790 2610 26795 2630
rect 26765 2580 26795 2610
rect 26765 2560 26770 2580
rect 26790 2560 26795 2580
rect 26765 2530 26795 2560
rect 26765 2510 26770 2530
rect 26790 2510 26795 2530
rect 26765 2500 26795 2510
rect 26825 2880 26855 2890
rect 26825 2860 26830 2880
rect 26850 2860 26855 2880
rect 26825 2830 26855 2860
rect 26825 2810 26830 2830
rect 26850 2810 26855 2830
rect 26825 2780 26855 2810
rect 26825 2760 26830 2780
rect 26850 2760 26855 2780
rect 26825 2730 26855 2760
rect 26825 2710 26830 2730
rect 26850 2710 26855 2730
rect 26825 2680 26855 2710
rect 26825 2660 26830 2680
rect 26850 2660 26855 2680
rect 26825 2630 26855 2660
rect 26825 2610 26830 2630
rect 26850 2610 26855 2630
rect 26825 2580 26855 2610
rect 26825 2560 26830 2580
rect 26850 2560 26855 2580
rect 26825 2530 26855 2560
rect 26825 2510 26830 2530
rect 26850 2510 26855 2530
rect 26825 2500 26855 2510
rect 26885 2880 26915 2890
rect 26885 2860 26890 2880
rect 26910 2860 26915 2880
rect 26885 2830 26915 2860
rect 26885 2810 26890 2830
rect 26910 2810 26915 2830
rect 26885 2780 26915 2810
rect 26885 2760 26890 2780
rect 26910 2760 26915 2780
rect 26885 2730 26915 2760
rect 26885 2710 26890 2730
rect 26910 2710 26915 2730
rect 26885 2680 26915 2710
rect 26885 2660 26890 2680
rect 26910 2660 26915 2680
rect 26885 2630 26915 2660
rect 26885 2610 26890 2630
rect 26910 2610 26915 2630
rect 26885 2580 26915 2610
rect 26885 2560 26890 2580
rect 26910 2560 26915 2580
rect 26885 2530 26915 2560
rect 26885 2510 26890 2530
rect 26910 2510 26915 2530
rect 26885 2500 26915 2510
rect 26945 2880 26975 2890
rect 26945 2860 26950 2880
rect 26970 2860 26975 2880
rect 26945 2830 26975 2860
rect 26945 2810 26950 2830
rect 26970 2810 26975 2830
rect 26945 2780 26975 2810
rect 26945 2760 26950 2780
rect 26970 2760 26975 2780
rect 26945 2730 26975 2760
rect 26945 2710 26950 2730
rect 26970 2710 26975 2730
rect 26945 2680 26975 2710
rect 26945 2660 26950 2680
rect 26970 2660 26975 2680
rect 26945 2630 26975 2660
rect 26945 2610 26950 2630
rect 26970 2610 26975 2630
rect 26945 2580 26975 2610
rect 26945 2560 26950 2580
rect 26970 2560 26975 2580
rect 26945 2530 26975 2560
rect 26945 2510 26950 2530
rect 26970 2510 26975 2530
rect 26945 2500 26975 2510
rect 27005 2880 27035 2890
rect 27005 2860 27010 2880
rect 27030 2860 27035 2880
rect 27005 2830 27035 2860
rect 27005 2810 27010 2830
rect 27030 2810 27035 2830
rect 27005 2780 27035 2810
rect 27005 2760 27010 2780
rect 27030 2760 27035 2780
rect 27005 2730 27035 2760
rect 27005 2710 27010 2730
rect 27030 2710 27035 2730
rect 27005 2680 27035 2710
rect 27005 2660 27010 2680
rect 27030 2660 27035 2680
rect 27005 2630 27035 2660
rect 27005 2610 27010 2630
rect 27030 2610 27035 2630
rect 27005 2580 27035 2610
rect 27005 2560 27010 2580
rect 27030 2560 27035 2580
rect 27005 2530 27035 2560
rect 27005 2510 27010 2530
rect 27030 2510 27035 2530
rect 27005 2500 27035 2510
rect 27065 2880 27095 2890
rect 27065 2860 27070 2880
rect 27090 2860 27095 2880
rect 27065 2830 27095 2860
rect 27065 2810 27070 2830
rect 27090 2810 27095 2830
rect 27065 2780 27095 2810
rect 27065 2760 27070 2780
rect 27090 2760 27095 2780
rect 27065 2730 27095 2760
rect 27065 2710 27070 2730
rect 27090 2710 27095 2730
rect 27065 2680 27095 2710
rect 27065 2660 27070 2680
rect 27090 2660 27095 2680
rect 27065 2630 27095 2660
rect 27065 2610 27070 2630
rect 27090 2610 27095 2630
rect 27065 2580 27095 2610
rect 27065 2560 27070 2580
rect 27090 2560 27095 2580
rect 27065 2530 27095 2560
rect 27065 2510 27070 2530
rect 27090 2510 27095 2530
rect 27065 2500 27095 2510
rect 27125 2880 27155 2890
rect 27125 2860 27130 2880
rect 27150 2860 27155 2880
rect 27125 2830 27155 2860
rect 27125 2810 27130 2830
rect 27150 2810 27155 2830
rect 27125 2780 27155 2810
rect 27125 2760 27130 2780
rect 27150 2760 27155 2780
rect 27125 2730 27155 2760
rect 27125 2710 27130 2730
rect 27150 2710 27155 2730
rect 27125 2680 27155 2710
rect 27125 2660 27130 2680
rect 27150 2660 27155 2680
rect 27125 2630 27155 2660
rect 27125 2610 27130 2630
rect 27150 2610 27155 2630
rect 27125 2580 27155 2610
rect 27125 2560 27130 2580
rect 27150 2560 27155 2580
rect 27125 2530 27155 2560
rect 27125 2510 27130 2530
rect 27150 2510 27155 2530
rect 27125 2500 27155 2510
rect 27185 2880 27215 2890
rect 27185 2860 27190 2880
rect 27210 2860 27215 2880
rect 27185 2830 27215 2860
rect 27185 2810 27190 2830
rect 27210 2810 27215 2830
rect 27185 2780 27215 2810
rect 27185 2760 27190 2780
rect 27210 2760 27215 2780
rect 27185 2730 27215 2760
rect 27185 2710 27190 2730
rect 27210 2710 27215 2730
rect 27185 2680 27215 2710
rect 27185 2660 27190 2680
rect 27210 2660 27215 2680
rect 27185 2630 27215 2660
rect 27185 2610 27190 2630
rect 27210 2610 27215 2630
rect 27185 2580 27215 2610
rect 27185 2560 27190 2580
rect 27210 2560 27215 2580
rect 27185 2530 27215 2560
rect 27185 2510 27190 2530
rect 27210 2510 27215 2530
rect 27185 2500 27215 2510
rect 27245 2880 27275 2890
rect 27245 2860 27250 2880
rect 27270 2860 27275 2880
rect 27245 2830 27275 2860
rect 27245 2810 27250 2830
rect 27270 2810 27275 2830
rect 27245 2780 27275 2810
rect 27245 2760 27250 2780
rect 27270 2760 27275 2780
rect 27245 2730 27275 2760
rect 27245 2710 27250 2730
rect 27270 2710 27275 2730
rect 27245 2680 27275 2710
rect 27245 2660 27250 2680
rect 27270 2660 27275 2680
rect 27245 2630 27275 2660
rect 27245 2610 27250 2630
rect 27270 2610 27275 2630
rect 27245 2580 27275 2610
rect 27245 2560 27250 2580
rect 27270 2560 27275 2580
rect 27245 2530 27275 2560
rect 27245 2510 27250 2530
rect 27270 2510 27275 2530
rect 27245 2500 27275 2510
rect 27305 2880 27335 2890
rect 27305 2860 27310 2880
rect 27330 2860 27335 2880
rect 27305 2830 27335 2860
rect 27305 2810 27310 2830
rect 27330 2810 27335 2830
rect 27305 2780 27335 2810
rect 27305 2760 27310 2780
rect 27330 2760 27335 2780
rect 27305 2730 27335 2760
rect 27305 2710 27310 2730
rect 27330 2710 27335 2730
rect 27305 2680 27335 2710
rect 27305 2660 27310 2680
rect 27330 2660 27335 2680
rect 27305 2630 27335 2660
rect 27305 2610 27310 2630
rect 27330 2610 27335 2630
rect 27305 2580 27335 2610
rect 27305 2560 27310 2580
rect 27330 2560 27335 2580
rect 27305 2530 27335 2560
rect 27305 2510 27310 2530
rect 27330 2510 27335 2530
rect 27305 2500 27335 2510
rect 27365 2880 27395 2890
rect 27365 2860 27370 2880
rect 27390 2860 27395 2880
rect 27365 2830 27395 2860
rect 27365 2810 27370 2830
rect 27390 2810 27395 2830
rect 27365 2780 27395 2810
rect 27365 2760 27370 2780
rect 27390 2760 27395 2780
rect 27365 2730 27395 2760
rect 27365 2710 27370 2730
rect 27390 2710 27395 2730
rect 27365 2680 27395 2710
rect 27365 2660 27370 2680
rect 27390 2660 27395 2680
rect 27365 2630 27395 2660
rect 27365 2610 27370 2630
rect 27390 2610 27395 2630
rect 27365 2580 27395 2610
rect 27365 2560 27370 2580
rect 27390 2560 27395 2580
rect 27365 2530 27395 2560
rect 27365 2510 27370 2530
rect 27390 2510 27395 2530
rect 27365 2500 27395 2510
rect 27425 2880 27455 2890
rect 27425 2860 27430 2880
rect 27450 2860 27455 2880
rect 27425 2830 27455 2860
rect 27425 2810 27430 2830
rect 27450 2810 27455 2830
rect 27425 2780 27455 2810
rect 27425 2760 27430 2780
rect 27450 2760 27455 2780
rect 27425 2730 27455 2760
rect 27425 2710 27430 2730
rect 27450 2710 27455 2730
rect 27425 2680 27455 2710
rect 27425 2660 27430 2680
rect 27450 2660 27455 2680
rect 27425 2630 27455 2660
rect 27425 2610 27430 2630
rect 27450 2610 27455 2630
rect 27425 2580 27455 2610
rect 27425 2560 27430 2580
rect 27450 2560 27455 2580
rect 27425 2530 27455 2560
rect 27425 2510 27430 2530
rect 27450 2510 27455 2530
rect 27425 2500 27455 2510
rect 27485 2880 27515 2890
rect 27485 2860 27490 2880
rect 27510 2860 27515 2880
rect 27485 2830 27515 2860
rect 27485 2810 27490 2830
rect 27510 2810 27515 2830
rect 27485 2780 27515 2810
rect 27485 2760 27490 2780
rect 27510 2760 27515 2780
rect 27485 2730 27515 2760
rect 27485 2710 27490 2730
rect 27510 2710 27515 2730
rect 27485 2680 27515 2710
rect 27485 2660 27490 2680
rect 27510 2660 27515 2680
rect 27485 2630 27515 2660
rect 27485 2610 27490 2630
rect 27510 2610 27515 2630
rect 27485 2580 27515 2610
rect 27485 2560 27490 2580
rect 27510 2560 27515 2580
rect 27485 2530 27515 2560
rect 27485 2510 27490 2530
rect 27510 2510 27515 2530
rect 27485 2500 27515 2510
rect 27545 2880 27615 2890
rect 27850 2885 27890 2895
rect 28000 2915 28040 2925
rect 28000 2895 28010 2915
rect 28030 2895 28040 2915
rect 28000 2885 28040 2895
rect 28058 2915 28092 2925
rect 28058 2895 28066 2915
rect 28084 2895 28092 2915
rect 28058 2885 28092 2895
rect 28110 2915 28150 2925
rect 28110 2895 28120 2915
rect 28140 2895 28150 2915
rect 28110 2885 28150 2895
rect 28220 2915 28260 2925
rect 28220 2895 28230 2915
rect 28250 2895 28260 2915
rect 28220 2885 28260 2895
rect 28330 2915 28370 2925
rect 28330 2895 28340 2915
rect 28360 2895 28370 2915
rect 28330 2885 28370 2895
rect 28440 2915 28480 2925
rect 28440 2895 28450 2915
rect 28470 2895 28480 2915
rect 28440 2885 28480 2895
rect 28550 2915 28590 2925
rect 28550 2895 28560 2915
rect 28580 2895 28590 2915
rect 28550 2885 28590 2895
rect 28660 2915 28700 2925
rect 28660 2895 28670 2915
rect 28690 2895 28700 2915
rect 28660 2885 28700 2895
rect 28770 2915 28810 2925
rect 28770 2895 28780 2915
rect 28800 2895 28810 2915
rect 28770 2885 28810 2895
rect 28880 2915 28920 2925
rect 28880 2895 28890 2915
rect 28910 2895 28920 2915
rect 28880 2885 28920 2895
rect 28990 2915 29030 2925
rect 28990 2895 29000 2915
rect 29020 2895 29030 2915
rect 28990 2885 29030 2895
rect 29140 2915 29180 2925
rect 29140 2895 29150 2915
rect 29170 2895 29180 2915
rect 29140 2885 29180 2895
rect 27545 2860 27550 2880
rect 27570 2860 27590 2880
rect 27610 2860 27615 2880
rect 27545 2830 27615 2860
rect 27545 2810 27550 2830
rect 27570 2810 27590 2830
rect 27610 2810 27615 2830
rect 27545 2780 27615 2810
rect 27545 2760 27550 2780
rect 27570 2760 27590 2780
rect 27610 2760 27615 2780
rect 27545 2730 27615 2760
rect 27545 2710 27550 2730
rect 27570 2710 27590 2730
rect 27610 2710 27615 2730
rect 27545 2680 27615 2710
rect 28055 2695 28095 2836
rect 27545 2660 27550 2680
rect 27570 2660 27590 2680
rect 27610 2660 27615 2680
rect 27545 2630 27615 2660
rect 27945 2665 27985 2675
rect 27945 2645 27955 2665
rect 27975 2645 27985 2665
rect 27945 2635 27985 2645
rect 28055 2665 28095 2675
rect 28055 2645 28065 2665
rect 28085 2645 28095 2665
rect 28055 2635 28095 2645
rect 28165 2665 28205 2675
rect 28165 2645 28175 2665
rect 28195 2645 28205 2665
rect 28165 2635 28205 2645
rect 28275 2665 28315 2675
rect 28275 2645 28285 2665
rect 28305 2645 28315 2665
rect 28275 2635 28315 2645
rect 28385 2665 28425 2675
rect 28385 2645 28395 2665
rect 28415 2645 28425 2665
rect 28385 2635 28425 2645
rect 28495 2665 28535 2675
rect 28495 2645 28505 2665
rect 28525 2645 28535 2665
rect 28495 2635 28535 2645
rect 28605 2665 28645 2675
rect 28605 2645 28615 2665
rect 28635 2645 28645 2665
rect 28605 2635 28645 2645
rect 28715 2665 28755 2675
rect 28715 2645 28725 2665
rect 28745 2645 28755 2665
rect 28715 2635 28755 2645
rect 28825 2665 28865 2675
rect 28825 2645 28835 2665
rect 28855 2645 28865 2665
rect 28825 2635 28865 2645
rect 28935 2665 28975 2675
rect 28935 2645 28945 2665
rect 28965 2645 28975 2665
rect 28935 2635 28975 2645
rect 29045 2665 29085 2675
rect 29045 2645 29055 2665
rect 29075 2645 29085 2665
rect 29045 2635 29085 2645
rect 27545 2610 27550 2630
rect 27570 2610 27590 2630
rect 27610 2610 27615 2630
rect 27955 2615 27975 2635
rect 28065 2615 28085 2635
rect 28175 2615 28195 2635
rect 28285 2615 28305 2635
rect 28395 2615 28415 2635
rect 28505 2615 28525 2635
rect 28615 2615 28635 2635
rect 28725 2615 28745 2635
rect 28835 2615 28855 2635
rect 28945 2615 28965 2635
rect 29055 2615 29075 2635
rect 27545 2580 27615 2610
rect 27545 2560 27550 2580
rect 27570 2560 27590 2580
rect 27610 2560 27615 2580
rect 27545 2530 27615 2560
rect 27545 2510 27550 2530
rect 27570 2510 27590 2530
rect 27610 2510 27615 2530
rect 27855 2605 27925 2615
rect 27855 2585 27860 2605
rect 27880 2585 27900 2605
rect 27920 2585 27925 2605
rect 27855 2555 27925 2585
rect 27855 2535 27860 2555
rect 27880 2535 27900 2555
rect 27920 2535 27925 2555
rect 27855 2525 27925 2535
rect 27950 2605 27980 2615
rect 27950 2585 27955 2605
rect 27975 2585 27980 2605
rect 27950 2555 27980 2585
rect 27950 2535 27955 2555
rect 27975 2535 27980 2555
rect 27950 2525 27980 2535
rect 28005 2605 28035 2615
rect 28005 2585 28010 2605
rect 28030 2585 28035 2605
rect 28005 2555 28035 2585
rect 28005 2535 28010 2555
rect 28030 2535 28035 2555
rect 28005 2525 28035 2535
rect 28060 2605 28090 2615
rect 28060 2585 28065 2605
rect 28085 2585 28090 2605
rect 28060 2555 28090 2585
rect 28060 2535 28065 2555
rect 28085 2535 28090 2555
rect 28060 2525 28090 2535
rect 28115 2605 28145 2615
rect 28115 2585 28120 2605
rect 28140 2585 28145 2605
rect 28115 2555 28145 2585
rect 28115 2535 28120 2555
rect 28140 2535 28145 2555
rect 28115 2525 28145 2535
rect 28170 2605 28200 2615
rect 28170 2585 28175 2605
rect 28195 2585 28200 2605
rect 28170 2555 28200 2585
rect 28170 2535 28175 2555
rect 28195 2535 28200 2555
rect 28170 2525 28200 2535
rect 28225 2605 28255 2615
rect 28225 2585 28230 2605
rect 28250 2585 28255 2605
rect 28225 2555 28255 2585
rect 28225 2535 28230 2555
rect 28250 2535 28255 2555
rect 28225 2525 28255 2535
rect 28280 2605 28310 2615
rect 28280 2585 28285 2605
rect 28305 2585 28310 2605
rect 28280 2555 28310 2585
rect 28280 2535 28285 2555
rect 28305 2535 28310 2555
rect 28280 2525 28310 2535
rect 28335 2605 28365 2615
rect 28335 2585 28340 2605
rect 28360 2585 28365 2605
rect 28335 2555 28365 2585
rect 28335 2535 28340 2555
rect 28360 2535 28365 2555
rect 28335 2525 28365 2535
rect 28390 2605 28420 2615
rect 28390 2585 28395 2605
rect 28415 2585 28420 2605
rect 28390 2555 28420 2585
rect 28390 2535 28395 2555
rect 28415 2535 28420 2555
rect 28390 2525 28420 2535
rect 28445 2605 28475 2615
rect 28445 2585 28450 2605
rect 28470 2585 28475 2605
rect 28445 2555 28475 2585
rect 28445 2535 28450 2555
rect 28470 2535 28475 2555
rect 28445 2525 28475 2535
rect 28500 2605 28530 2615
rect 28500 2585 28505 2605
rect 28525 2585 28530 2605
rect 28500 2555 28530 2585
rect 28500 2535 28505 2555
rect 28525 2535 28530 2555
rect 28500 2525 28530 2535
rect 28555 2605 28585 2615
rect 28555 2585 28560 2605
rect 28580 2585 28585 2605
rect 28555 2555 28585 2585
rect 28555 2535 28560 2555
rect 28580 2535 28585 2555
rect 28555 2525 28585 2535
rect 28610 2605 28640 2615
rect 28610 2585 28615 2605
rect 28635 2585 28640 2605
rect 28610 2555 28640 2585
rect 28610 2535 28615 2555
rect 28635 2535 28640 2555
rect 28610 2525 28640 2535
rect 28665 2605 28695 2615
rect 28665 2585 28670 2605
rect 28690 2585 28695 2605
rect 28665 2555 28695 2585
rect 28665 2535 28670 2555
rect 28690 2535 28695 2555
rect 28665 2525 28695 2535
rect 28720 2605 28750 2615
rect 28720 2585 28725 2605
rect 28745 2585 28750 2605
rect 28720 2555 28750 2585
rect 28720 2535 28725 2555
rect 28745 2535 28750 2555
rect 28720 2525 28750 2535
rect 28775 2605 28805 2615
rect 28775 2585 28780 2605
rect 28800 2585 28805 2605
rect 28775 2555 28805 2585
rect 28775 2535 28780 2555
rect 28800 2535 28805 2555
rect 28775 2525 28805 2535
rect 28830 2605 28860 2615
rect 28830 2585 28835 2605
rect 28855 2585 28860 2605
rect 28830 2555 28860 2585
rect 28830 2535 28835 2555
rect 28855 2535 28860 2555
rect 28830 2525 28860 2535
rect 28885 2605 28915 2615
rect 28885 2585 28890 2605
rect 28910 2585 28915 2605
rect 28885 2555 28915 2585
rect 28885 2535 28890 2555
rect 28910 2535 28915 2555
rect 28885 2525 28915 2535
rect 28940 2605 28970 2615
rect 28940 2585 28945 2605
rect 28965 2585 28970 2605
rect 28940 2555 28970 2585
rect 28940 2535 28945 2555
rect 28965 2535 28970 2555
rect 28940 2525 28970 2535
rect 28995 2605 29025 2615
rect 28995 2585 29000 2605
rect 29020 2585 29025 2605
rect 28995 2555 29025 2585
rect 28995 2535 29000 2555
rect 29020 2535 29025 2555
rect 28995 2525 29025 2535
rect 29050 2605 29080 2615
rect 29050 2585 29055 2605
rect 29075 2585 29080 2605
rect 29050 2555 29080 2585
rect 29050 2535 29055 2555
rect 29075 2535 29080 2555
rect 29050 2525 29080 2535
rect 29105 2605 29175 2615
rect 29105 2585 29110 2605
rect 29130 2585 29150 2605
rect 29170 2585 29175 2605
rect 29105 2555 29175 2585
rect 29105 2535 29110 2555
rect 29130 2535 29150 2555
rect 29170 2535 29175 2555
rect 29105 2525 29175 2535
rect 27545 2500 27615 2510
rect 27860 2505 27880 2525
rect 28010 2505 28030 2525
rect 28120 2505 28140 2525
rect 28230 2505 28250 2525
rect 28340 2505 28360 2525
rect 28450 2505 28470 2525
rect 28560 2505 28580 2525
rect 28670 2505 28690 2525
rect 28780 2505 28800 2525
rect 28890 2505 28910 2525
rect 29000 2505 29020 2525
rect 29150 2505 29170 2525
rect 25930 2475 25940 2495
rect 25960 2475 25970 2495
rect 26290 2480 26310 2500
rect 26410 2480 26430 2500
rect 26530 2480 26550 2500
rect 26650 2480 26670 2500
rect 26770 2480 26790 2500
rect 26890 2480 26910 2500
rect 27010 2480 27030 2500
rect 27130 2480 27150 2500
rect 27250 2480 27270 2500
rect 27370 2480 27390 2500
rect 27490 2480 27510 2500
rect 27850 2495 27890 2505
rect 25930 2465 25970 2475
rect 26280 2470 26320 2480
rect 26280 2450 26290 2470
rect 26310 2450 26320 2470
rect 25813 2435 25847 2445
rect 26280 2440 26320 2450
rect 26400 2470 26440 2480
rect 26400 2450 26410 2470
rect 26430 2450 26440 2470
rect 26400 2440 26440 2450
rect 26520 2470 26560 2480
rect 26520 2450 26530 2470
rect 26550 2450 26560 2470
rect 26520 2440 26560 2450
rect 26640 2470 26680 2480
rect 26640 2450 26650 2470
rect 26670 2450 26680 2470
rect 26640 2440 26680 2450
rect 26760 2470 26800 2480
rect 26760 2450 26770 2470
rect 26790 2450 26800 2470
rect 26760 2440 26800 2450
rect 26823 2470 26857 2480
rect 26823 2450 26831 2470
rect 26849 2450 26857 2470
rect 26823 2440 26857 2450
rect 26880 2470 26920 2480
rect 26880 2450 26890 2470
rect 26910 2450 26920 2470
rect 26880 2440 26920 2450
rect 27000 2470 27040 2480
rect 27000 2450 27010 2470
rect 27030 2450 27040 2470
rect 27000 2440 27040 2450
rect 27120 2470 27160 2480
rect 27120 2450 27130 2470
rect 27150 2450 27160 2470
rect 27120 2440 27160 2450
rect 27240 2470 27280 2480
rect 27240 2450 27250 2470
rect 27270 2450 27280 2470
rect 27240 2440 27280 2450
rect 27360 2470 27400 2480
rect 27360 2450 27370 2470
rect 27390 2450 27400 2470
rect 27360 2440 27400 2450
rect 27480 2470 27520 2480
rect 27480 2450 27490 2470
rect 27510 2450 27520 2470
rect 27850 2475 27860 2495
rect 27880 2475 27890 2495
rect 27850 2465 27890 2475
rect 28000 2495 28040 2505
rect 28000 2475 28010 2495
rect 28030 2475 28040 2495
rect 28000 2465 28040 2475
rect 28110 2495 28150 2505
rect 28110 2475 28120 2495
rect 28140 2475 28150 2495
rect 28110 2465 28150 2475
rect 28220 2495 28260 2505
rect 28220 2475 28230 2495
rect 28250 2475 28260 2495
rect 28220 2465 28260 2475
rect 28330 2495 28370 2505
rect 28330 2475 28340 2495
rect 28360 2475 28370 2495
rect 28330 2465 28370 2475
rect 28440 2495 28480 2505
rect 28440 2475 28450 2495
rect 28470 2475 28480 2495
rect 28440 2465 28480 2475
rect 28550 2495 28590 2505
rect 28550 2475 28560 2495
rect 28580 2475 28590 2495
rect 28550 2465 28590 2475
rect 28660 2495 28700 2505
rect 28660 2475 28670 2495
rect 28690 2475 28700 2495
rect 28660 2465 28700 2475
rect 28770 2495 28810 2505
rect 28770 2475 28780 2495
rect 28800 2475 28810 2495
rect 28770 2465 28810 2475
rect 28880 2495 28920 2505
rect 28880 2475 28890 2495
rect 28910 2475 28920 2495
rect 28880 2465 28920 2475
rect 28990 2495 29030 2505
rect 28990 2475 29000 2495
rect 29020 2475 29030 2495
rect 28990 2465 29030 2475
rect 29140 2495 29180 2505
rect 29140 2475 29150 2495
rect 29170 2475 29180 2495
rect 29140 2465 29180 2475
rect 27480 2440 27520 2450
rect 25813 2415 25821 2435
rect 25839 2415 25847 2435
rect 25813 2405 25847 2415
rect 27973 2435 28007 2445
rect 27973 2415 27981 2435
rect 27999 2415 28007 2435
rect 27973 2405 28007 2415
rect 10765 2385 10805 2395
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 10765 2365 10775 2385
rect 10795 2365 10805 2385
rect 10765 2355 10805 2365
rect 13025 2370 13065 2380
rect 4705 2345 4745 2355
rect 13025 2350 13035 2370
rect 13055 2350 13065 2370
rect 13025 2340 13065 2350
rect 24800 2375 24845 2380
rect 24800 2350 24810 2375
rect 24835 2350 24845 2375
rect 24800 2345 24845 2350
rect 25635 2375 25680 2380
rect 25635 2350 25645 2375
rect 25670 2350 25680 2375
rect 25635 2345 25680 2350
rect 28140 2375 28185 2380
rect 28140 2350 28150 2375
rect 28175 2350 28185 2375
rect 28140 2345 28185 2350
rect 28975 2375 29020 2380
rect 28975 2350 28985 2375
rect 29010 2350 29020 2375
rect 28975 2345 29020 2350
rect 3625 2330 3665 2340
rect 3625 2310 3635 2330
rect 3655 2310 3665 2330
rect 3625 2300 3665 2310
rect 4345 2330 4385 2340
rect 4345 2310 4355 2330
rect 4375 2310 4385 2330
rect 4345 2300 4385 2310
rect 10115 2310 10155 2320
rect 2740 2260 2770 2290
rect 3445 2285 3485 2295
rect 3445 2265 3455 2285
rect 3475 2265 3485 2285
rect 3445 2255 3485 2265
rect 4525 2285 4565 2295
rect 10115 2290 10125 2310
rect 10145 2290 10155 2310
rect 4525 2265 4535 2285
rect 4555 2265 4565 2285
rect 4525 2255 4565 2265
rect 5275 2260 5305 2290
rect 10115 2280 10155 2290
rect 10265 2310 10305 2320
rect 10265 2290 10275 2310
rect 10295 2290 10305 2310
rect 10265 2280 10305 2290
rect 10375 2310 10415 2320
rect 10375 2290 10385 2310
rect 10405 2290 10415 2310
rect 10375 2280 10415 2290
rect 10485 2310 10525 2320
rect 10485 2290 10495 2310
rect 10515 2290 10525 2310
rect 10485 2280 10525 2290
rect 10595 2310 10635 2320
rect 10595 2290 10605 2310
rect 10625 2290 10635 2310
rect 10595 2280 10635 2290
rect 10705 2310 10745 2320
rect 10705 2290 10715 2310
rect 10735 2290 10745 2310
rect 10705 2280 10745 2290
rect 10855 2310 10895 2320
rect 10855 2290 10865 2310
rect 10885 2290 10895 2310
rect 10855 2280 10895 2290
rect 12905 2310 12945 2320
rect 12905 2290 12915 2310
rect 12935 2290 12945 2310
rect 12905 2280 12945 2290
rect 13055 2310 13095 2320
rect 13055 2290 13065 2310
rect 13085 2290 13095 2310
rect 13055 2280 13095 2290
rect 13165 2310 13205 2320
rect 13165 2290 13175 2310
rect 13195 2290 13205 2310
rect 13165 2280 13205 2290
rect 13275 2310 13315 2320
rect 13275 2290 13285 2310
rect 13305 2290 13315 2310
rect 13275 2280 13315 2290
rect 13385 2310 13425 2320
rect 13385 2290 13395 2310
rect 13415 2290 13425 2310
rect 13385 2280 13425 2290
rect 13495 2310 13535 2320
rect 13495 2290 13505 2310
rect 13525 2290 13535 2310
rect 13495 2280 13535 2290
rect 13645 2310 13685 2320
rect 13645 2290 13655 2310
rect 13675 2290 13685 2310
rect 13645 2280 13685 2290
rect 24800 2315 24845 2320
rect 24800 2290 24810 2315
rect 24835 2290 24845 2315
rect 24800 2285 24845 2290
rect 25635 2315 25680 2320
rect 25635 2290 25645 2315
rect 25670 2290 25680 2315
rect 25635 2285 25680 2290
rect 28140 2315 28185 2320
rect 28140 2290 28150 2315
rect 28175 2290 28185 2315
rect 28140 2285 28185 2290
rect 28975 2315 29020 2320
rect 28975 2290 28985 2315
rect 29010 2290 29020 2315
rect 28975 2285 29020 2290
rect 10125 2260 10145 2280
rect 10275 2260 10295 2280
rect 10385 2260 10405 2280
rect 10495 2260 10515 2280
rect 10605 2260 10625 2280
rect 10715 2260 10735 2280
rect 10865 2260 10885 2280
rect 12915 2260 12935 2280
rect 13065 2260 13085 2280
rect 13175 2260 13195 2280
rect 13285 2260 13305 2280
rect 13395 2260 13415 2280
rect 13505 2260 13525 2280
rect 13655 2260 13675 2280
rect 25813 2275 25847 2285
rect 10120 2250 10190 2260
rect 2430 2215 2460 2245
rect 3810 2215 3840 2245
rect 10120 2230 10125 2250
rect 10145 2230 10165 2250
rect 10185 2230 10190 2250
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 3630 2120 3660 2150
rect 4090 2115 4120 2145
rect 5320 2115 5350 2145
rect 2745 2090 2785 2100
rect 2745 2070 2755 2090
rect 2775 2070 2785 2090
rect 2745 2060 2785 2070
rect 2865 2090 2905 2100
rect 2865 2070 2875 2090
rect 2895 2070 2905 2090
rect 2865 2060 2905 2070
rect 2985 2090 3025 2100
rect 2985 2070 2995 2090
rect 3015 2070 3025 2090
rect 2985 2060 3025 2070
rect 3105 2090 3145 2100
rect 3105 2070 3115 2090
rect 3135 2070 3145 2090
rect 3105 2060 3145 2070
rect 3225 2090 3265 2100
rect 3225 2070 3235 2090
rect 3255 2070 3265 2090
rect 3225 2060 3265 2070
rect 3345 2090 3385 2100
rect 3345 2070 3355 2090
rect 3375 2070 3385 2090
rect 3345 2060 3385 2070
rect 3465 2090 3505 2100
rect 3465 2070 3475 2090
rect 3495 2070 3505 2090
rect 3465 2060 3505 2070
rect 3585 2090 3625 2100
rect 3585 2070 3595 2090
rect 3615 2070 3625 2090
rect 3585 2060 3625 2070
rect 3705 2090 3745 2100
rect 3705 2070 3715 2090
rect 3735 2070 3745 2090
rect 3705 2060 3745 2070
rect 3825 2090 3865 2100
rect 3825 2070 3835 2090
rect 3855 2070 3865 2090
rect 3825 2060 3865 2070
rect 3985 2090 4025 2100
rect 3985 2070 3995 2090
rect 4015 2070 4025 2090
rect 3985 2060 4025 2070
rect 4145 2090 4185 2100
rect 4145 2070 4155 2090
rect 4175 2070 4185 2090
rect 4145 2060 4185 2070
rect 4265 2090 4305 2100
rect 4265 2070 4275 2090
rect 4295 2070 4305 2090
rect 4265 2060 4305 2070
rect 4385 2090 4425 2100
rect 4385 2070 4395 2090
rect 4415 2070 4425 2090
rect 4385 2060 4425 2070
rect 4505 2090 4545 2100
rect 4505 2070 4515 2090
rect 4535 2070 4545 2090
rect 4505 2060 4545 2070
rect 4625 2090 4665 2100
rect 4625 2070 4635 2090
rect 4655 2070 4665 2090
rect 4625 2060 4665 2070
rect 4745 2090 4785 2100
rect 4745 2070 4755 2090
rect 4775 2070 4785 2090
rect 4745 2060 4785 2070
rect 4865 2090 4905 2100
rect 4865 2070 4875 2090
rect 4895 2070 4905 2090
rect 4865 2060 4905 2070
rect 4985 2090 5025 2100
rect 4985 2070 4995 2090
rect 5015 2070 5025 2090
rect 4985 2060 5025 2070
rect 5105 2090 5145 2100
rect 5105 2070 5115 2090
rect 5135 2070 5145 2090
rect 5105 2060 5145 2070
rect 5225 2090 5265 2100
rect 5225 2070 5235 2090
rect 5255 2070 5265 2090
rect 5225 2060 5265 2070
rect 125 2015 2135 2055
rect 2620 2045 2660 2055
rect 2620 2025 2630 2045
rect 2650 2025 2660 2045
rect 2620 2015 2660 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2010 1375 2135 2015
rect 2630 1995 2650 2015
rect 2755 1995 2775 2060
rect 2805 2045 2845 2055
rect 2805 2025 2815 2045
rect 2835 2025 2845 2045
rect 2805 2015 2845 2025
rect 2815 1995 2835 2015
rect 2875 1995 2895 2060
rect 2995 1995 3015 2060
rect 3115 1995 3135 2060
rect 3165 2045 3205 2055
rect 3165 2025 3175 2045
rect 3195 2025 3205 2045
rect 3165 2015 3205 2025
rect 3175 1995 3195 2015
rect 3235 1995 3255 2060
rect 3355 1995 3375 2060
rect 3475 1995 3495 2060
rect 3525 2045 3565 2055
rect 3525 2025 3535 2045
rect 3555 2025 3565 2045
rect 3525 2015 3565 2025
rect 3535 1995 3555 2015
rect 3595 1995 3615 2060
rect 3715 1995 3735 2060
rect 3835 1995 3855 2060
rect 3885 2045 3925 2055
rect 3885 2025 3895 2045
rect 3915 2025 3925 2045
rect 3885 2015 3925 2025
rect 3895 1995 3915 2015
rect 3995 1995 4015 2060
rect 4085 2045 4125 2055
rect 4085 2025 4095 2045
rect 4115 2025 4125 2045
rect 4085 2015 4125 2025
rect 4095 1995 4115 2015
rect 4155 1995 4175 2060
rect 4275 1995 4295 2060
rect 4395 1995 4415 2060
rect 4445 2045 4485 2055
rect 4445 2025 4455 2045
rect 4475 2025 4485 2045
rect 4445 2015 4485 2025
rect 4455 1995 4475 2015
rect 4515 1995 4535 2060
rect 4635 1995 4655 2060
rect 4755 1995 4775 2060
rect 4805 2045 4845 2055
rect 4805 2025 4815 2045
rect 4835 2025 4845 2045
rect 4805 2015 4845 2025
rect 4815 1995 4835 2015
rect 4875 1995 4895 2060
rect 4995 1995 5015 2060
rect 5115 1995 5135 2060
rect 5165 2045 5205 2055
rect 5165 2025 5175 2045
rect 5195 2025 5205 2045
rect 5165 2015 5205 2025
rect 5175 1995 5195 2015
rect 5235 1995 5255 2060
rect 9790 2000 9825 2010
rect 2570 1985 2600 1995
rect 2570 1965 2575 1985
rect 2595 1965 2600 1985
rect 2570 1935 2600 1965
rect 2570 1915 2575 1935
rect 2595 1915 2600 1935
rect 2570 1905 2600 1915
rect 2625 1985 2655 1995
rect 2625 1965 2630 1985
rect 2650 1965 2655 1985
rect 2625 1935 2655 1965
rect 2625 1915 2630 1935
rect 2650 1915 2655 1935
rect 2625 1905 2655 1915
rect 2680 1985 2710 1995
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1905 2710 1915
rect 2750 1985 2780 1995
rect 2750 1965 2755 1985
rect 2775 1965 2780 1985
rect 2750 1935 2780 1965
rect 2750 1915 2755 1935
rect 2775 1915 2780 1935
rect 2750 1905 2780 1915
rect 2810 1985 2840 1995
rect 2810 1965 2815 1985
rect 2835 1965 2840 1985
rect 2810 1935 2840 1965
rect 2810 1915 2815 1935
rect 2835 1915 2840 1935
rect 2810 1905 2840 1915
rect 2870 1985 2900 1995
rect 2870 1965 2875 1985
rect 2895 1965 2900 1985
rect 2870 1935 2900 1965
rect 2870 1915 2875 1935
rect 2895 1915 2900 1935
rect 2870 1905 2900 1915
rect 2930 1985 2960 1995
rect 2930 1965 2935 1985
rect 2955 1965 2960 1985
rect 2930 1935 2960 1965
rect 2930 1915 2935 1935
rect 2955 1915 2960 1935
rect 2930 1905 2960 1915
rect 2990 1985 3020 1995
rect 2990 1965 2995 1985
rect 3015 1965 3020 1985
rect 2990 1935 3020 1965
rect 2990 1915 2995 1935
rect 3015 1915 3020 1935
rect 2990 1905 3020 1915
rect 3050 1985 3080 1995
rect 3050 1965 3055 1985
rect 3075 1965 3080 1985
rect 3050 1935 3080 1965
rect 3050 1915 3055 1935
rect 3075 1915 3080 1935
rect 3050 1905 3080 1915
rect 3110 1985 3140 1995
rect 3110 1965 3115 1985
rect 3135 1965 3140 1985
rect 3110 1935 3140 1965
rect 3110 1915 3115 1935
rect 3135 1915 3140 1935
rect 3110 1905 3140 1915
rect 3170 1985 3200 1995
rect 3170 1965 3175 1985
rect 3195 1965 3200 1985
rect 3170 1935 3200 1965
rect 3170 1915 3175 1935
rect 3195 1915 3200 1935
rect 3170 1905 3200 1915
rect 3230 1985 3260 1995
rect 3230 1965 3235 1985
rect 3255 1965 3260 1985
rect 3230 1935 3260 1965
rect 3230 1915 3235 1935
rect 3255 1915 3260 1935
rect 3230 1905 3260 1915
rect 3290 1985 3320 1995
rect 3290 1965 3295 1985
rect 3315 1965 3320 1985
rect 3290 1935 3320 1965
rect 3290 1915 3295 1935
rect 3315 1915 3320 1935
rect 3290 1905 3320 1915
rect 3350 1985 3380 1995
rect 3350 1965 3355 1985
rect 3375 1965 3380 1985
rect 3350 1935 3380 1965
rect 3350 1915 3355 1935
rect 3375 1915 3380 1935
rect 3350 1905 3380 1915
rect 3410 1985 3440 1995
rect 3410 1965 3415 1985
rect 3435 1965 3440 1985
rect 3410 1935 3440 1965
rect 3410 1915 3415 1935
rect 3435 1915 3440 1935
rect 3410 1905 3440 1915
rect 3470 1985 3500 1995
rect 3470 1965 3475 1985
rect 3495 1965 3500 1985
rect 3470 1935 3500 1965
rect 3470 1915 3475 1935
rect 3495 1915 3500 1935
rect 3470 1905 3500 1915
rect 3530 1985 3560 1995
rect 3530 1965 3535 1985
rect 3555 1965 3560 1985
rect 3530 1935 3560 1965
rect 3530 1915 3535 1935
rect 3555 1915 3560 1935
rect 3530 1905 3560 1915
rect 3590 1985 3620 1995
rect 3590 1965 3595 1985
rect 3615 1965 3620 1985
rect 3590 1935 3620 1965
rect 3590 1915 3595 1935
rect 3615 1915 3620 1935
rect 3590 1905 3620 1915
rect 3650 1985 3680 1995
rect 3650 1965 3655 1985
rect 3675 1965 3680 1985
rect 3650 1935 3680 1965
rect 3650 1915 3655 1935
rect 3675 1915 3680 1935
rect 3650 1905 3680 1915
rect 3710 1985 3740 1995
rect 3710 1965 3715 1985
rect 3735 1965 3740 1985
rect 3710 1935 3740 1965
rect 3710 1915 3715 1935
rect 3735 1915 3740 1935
rect 3710 1905 3740 1915
rect 3770 1985 3800 1995
rect 3770 1965 3775 1985
rect 3795 1965 3800 1985
rect 3770 1935 3800 1965
rect 3770 1915 3775 1935
rect 3795 1915 3800 1935
rect 3770 1905 3800 1915
rect 3830 1985 3860 1995
rect 3830 1965 3835 1985
rect 3855 1965 3860 1985
rect 3830 1935 3860 1965
rect 3830 1915 3835 1935
rect 3855 1915 3860 1935
rect 3830 1905 3860 1915
rect 3890 1985 3920 1995
rect 3890 1965 3895 1985
rect 3915 1965 3920 1985
rect 3890 1935 3920 1965
rect 3890 1915 3895 1935
rect 3915 1915 3920 1935
rect 3890 1905 3920 1915
rect 3950 1985 4060 1995
rect 3950 1965 3955 1985
rect 3975 1965 3995 1985
rect 4015 1965 4035 1985
rect 4055 1965 4060 1985
rect 3950 1935 4060 1965
rect 3950 1915 3955 1935
rect 3975 1915 3995 1935
rect 4015 1915 4035 1935
rect 4055 1915 4060 1935
rect 3950 1905 4060 1915
rect 4090 1985 4120 1995
rect 4090 1965 4095 1985
rect 4115 1965 4120 1985
rect 4090 1935 4120 1965
rect 4090 1915 4095 1935
rect 4115 1915 4120 1935
rect 4090 1905 4120 1915
rect 4150 1985 4180 1995
rect 4150 1965 4155 1985
rect 4175 1965 4180 1985
rect 4150 1935 4180 1965
rect 4150 1915 4155 1935
rect 4175 1915 4180 1935
rect 4150 1905 4180 1915
rect 4210 1985 4240 1995
rect 4210 1965 4215 1985
rect 4235 1965 4240 1985
rect 4210 1935 4240 1965
rect 4210 1915 4215 1935
rect 4235 1915 4240 1935
rect 4210 1905 4240 1915
rect 4270 1985 4300 1995
rect 4270 1965 4275 1985
rect 4295 1965 4300 1985
rect 4270 1935 4300 1965
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1905 4300 1915
rect 4330 1985 4360 1995
rect 4330 1965 4335 1985
rect 4355 1965 4360 1985
rect 4330 1935 4360 1965
rect 4330 1915 4335 1935
rect 4355 1915 4360 1935
rect 4330 1905 4360 1915
rect 4390 1985 4420 1995
rect 4390 1965 4395 1985
rect 4415 1965 4420 1985
rect 4390 1935 4420 1965
rect 4390 1915 4395 1935
rect 4415 1915 4420 1935
rect 4390 1905 4420 1915
rect 4450 1985 4480 1995
rect 4450 1965 4455 1985
rect 4475 1965 4480 1985
rect 4450 1935 4480 1965
rect 4450 1915 4455 1935
rect 4475 1915 4480 1935
rect 4450 1905 4480 1915
rect 4510 1985 4540 1995
rect 4510 1965 4515 1985
rect 4535 1965 4540 1985
rect 4510 1935 4540 1965
rect 4510 1915 4515 1935
rect 4535 1915 4540 1935
rect 4510 1905 4540 1915
rect 4570 1985 4600 1995
rect 4570 1965 4575 1985
rect 4595 1965 4600 1985
rect 4570 1935 4600 1965
rect 4570 1915 4575 1935
rect 4595 1915 4600 1935
rect 4570 1905 4600 1915
rect 4630 1985 4660 1995
rect 4630 1965 4635 1985
rect 4655 1965 4660 1985
rect 4630 1935 4660 1965
rect 4630 1915 4635 1935
rect 4655 1915 4660 1935
rect 4630 1905 4660 1915
rect 4690 1985 4720 1995
rect 4690 1965 4695 1985
rect 4715 1965 4720 1985
rect 4690 1935 4720 1965
rect 4690 1915 4695 1935
rect 4715 1915 4720 1935
rect 4690 1905 4720 1915
rect 4750 1985 4780 1995
rect 4750 1965 4755 1985
rect 4775 1965 4780 1985
rect 4750 1935 4780 1965
rect 4750 1915 4755 1935
rect 4775 1915 4780 1935
rect 4750 1905 4780 1915
rect 4810 1985 4840 1995
rect 4810 1965 4815 1985
rect 4835 1965 4840 1985
rect 4810 1935 4840 1965
rect 4810 1915 4815 1935
rect 4835 1915 4840 1935
rect 4810 1905 4840 1915
rect 4870 1985 4900 1995
rect 4870 1965 4875 1985
rect 4895 1965 4900 1985
rect 4870 1935 4900 1965
rect 4870 1915 4875 1935
rect 4895 1915 4900 1935
rect 4870 1905 4900 1915
rect 4930 1985 4960 1995
rect 4930 1965 4935 1985
rect 4955 1965 4960 1985
rect 4930 1935 4960 1965
rect 4930 1915 4935 1935
rect 4955 1915 4960 1935
rect 4930 1905 4960 1915
rect 4990 1985 5020 1995
rect 4990 1965 4995 1985
rect 5015 1965 5020 1985
rect 4990 1935 5020 1965
rect 4990 1915 4995 1935
rect 5015 1915 5020 1935
rect 4990 1905 5020 1915
rect 5050 1985 5080 1995
rect 5050 1965 5055 1985
rect 5075 1965 5080 1985
rect 5050 1935 5080 1965
rect 5050 1915 5055 1935
rect 5075 1915 5080 1935
rect 5050 1905 5080 1915
rect 5110 1985 5140 1995
rect 5110 1965 5115 1985
rect 5135 1965 5140 1985
rect 5110 1935 5140 1965
rect 5110 1915 5115 1935
rect 5135 1915 5140 1935
rect 5110 1905 5140 1915
rect 5170 1985 5200 1995
rect 5170 1965 5175 1985
rect 5195 1965 5200 1985
rect 5170 1935 5200 1965
rect 5170 1915 5175 1935
rect 5195 1915 5200 1935
rect 5170 1905 5200 1915
rect 5230 1985 5260 1995
rect 5230 1965 5235 1985
rect 5255 1965 5260 1985
rect 9790 1975 9795 2000
rect 9820 1975 9825 2000
rect 9790 1965 9825 1975
rect 9850 2000 9885 2010
rect 9850 1975 9855 2000
rect 9880 1975 9885 2000
rect 9850 1965 9885 1975
rect 9910 2000 9945 2010
rect 9910 1975 9915 2000
rect 9940 1975 9945 2000
rect 9910 1965 9945 1975
rect 9970 2000 10005 2010
rect 9970 1975 9975 2000
rect 10000 1975 10005 2000
rect 9970 1965 10005 1975
rect 10120 2200 10190 2230
rect 10120 2180 10125 2200
rect 10145 2180 10165 2200
rect 10185 2180 10190 2200
rect 10120 2150 10190 2180
rect 10120 2130 10125 2150
rect 10145 2130 10165 2150
rect 10185 2130 10190 2150
rect 10120 2100 10190 2130
rect 10120 2080 10125 2100
rect 10145 2080 10165 2100
rect 10185 2080 10190 2100
rect 10120 2050 10190 2080
rect 10120 2030 10125 2050
rect 10145 2030 10165 2050
rect 10185 2030 10190 2050
rect 10120 2000 10190 2030
rect 10120 1980 10125 2000
rect 10145 1980 10165 2000
rect 10185 1980 10190 2000
rect 10120 1970 10190 1980
rect 10215 2250 10245 2260
rect 10215 2230 10220 2250
rect 10240 2230 10245 2250
rect 10215 2200 10245 2230
rect 10215 2180 10220 2200
rect 10240 2180 10245 2200
rect 10215 2150 10245 2180
rect 10215 2130 10220 2150
rect 10240 2130 10245 2150
rect 10215 2100 10245 2130
rect 10215 2080 10220 2100
rect 10240 2080 10245 2100
rect 10215 2050 10245 2080
rect 10215 2030 10220 2050
rect 10240 2030 10245 2050
rect 10215 2000 10245 2030
rect 10215 1980 10220 2000
rect 10240 1980 10245 2000
rect 10215 1970 10245 1980
rect 10270 2250 10300 2260
rect 10270 2230 10275 2250
rect 10295 2230 10300 2250
rect 10270 2200 10300 2230
rect 10270 2180 10275 2200
rect 10295 2180 10300 2200
rect 10270 2150 10300 2180
rect 10270 2130 10275 2150
rect 10295 2130 10300 2150
rect 10270 2100 10300 2130
rect 10270 2080 10275 2100
rect 10295 2080 10300 2100
rect 10270 2050 10300 2080
rect 10270 2030 10275 2050
rect 10295 2030 10300 2050
rect 10270 2000 10300 2030
rect 10270 1980 10275 2000
rect 10295 1980 10300 2000
rect 10270 1970 10300 1980
rect 10325 2250 10355 2260
rect 10325 2230 10330 2250
rect 10350 2230 10355 2250
rect 10325 2200 10355 2230
rect 10325 2180 10330 2200
rect 10350 2180 10355 2200
rect 10325 2150 10355 2180
rect 10325 2130 10330 2150
rect 10350 2130 10355 2150
rect 10325 2100 10355 2130
rect 10325 2080 10330 2100
rect 10350 2080 10355 2100
rect 10325 2050 10355 2080
rect 10325 2030 10330 2050
rect 10350 2030 10355 2050
rect 10325 2000 10355 2030
rect 10325 1980 10330 2000
rect 10350 1980 10355 2000
rect 10325 1970 10355 1980
rect 10380 2250 10410 2260
rect 10380 2230 10385 2250
rect 10405 2230 10410 2250
rect 10380 2200 10410 2230
rect 10380 2180 10385 2200
rect 10405 2180 10410 2200
rect 10380 2150 10410 2180
rect 10380 2130 10385 2150
rect 10405 2130 10410 2150
rect 10380 2100 10410 2130
rect 10380 2080 10385 2100
rect 10405 2080 10410 2100
rect 10380 2050 10410 2080
rect 10380 2030 10385 2050
rect 10405 2030 10410 2050
rect 10380 2000 10410 2030
rect 10380 1980 10385 2000
rect 10405 1980 10410 2000
rect 10380 1970 10410 1980
rect 10435 2250 10465 2260
rect 10435 2230 10440 2250
rect 10460 2230 10465 2250
rect 10435 2200 10465 2230
rect 10435 2180 10440 2200
rect 10460 2180 10465 2200
rect 10435 2150 10465 2180
rect 10435 2130 10440 2150
rect 10460 2130 10465 2150
rect 10435 2100 10465 2130
rect 10435 2080 10440 2100
rect 10460 2080 10465 2100
rect 10435 2050 10465 2080
rect 10435 2030 10440 2050
rect 10460 2030 10465 2050
rect 10435 2000 10465 2030
rect 10435 1980 10440 2000
rect 10460 1980 10465 2000
rect 10435 1970 10465 1980
rect 10490 2250 10520 2260
rect 10490 2230 10495 2250
rect 10515 2230 10520 2250
rect 10490 2200 10520 2230
rect 10490 2180 10495 2200
rect 10515 2180 10520 2200
rect 10490 2150 10520 2180
rect 10490 2130 10495 2150
rect 10515 2130 10520 2150
rect 10490 2100 10520 2130
rect 10490 2080 10495 2100
rect 10515 2080 10520 2100
rect 10490 2050 10520 2080
rect 10490 2030 10495 2050
rect 10515 2030 10520 2050
rect 10490 2000 10520 2030
rect 10490 1980 10495 2000
rect 10515 1980 10520 2000
rect 10490 1970 10520 1980
rect 10545 2250 10575 2260
rect 10545 2230 10550 2250
rect 10570 2230 10575 2250
rect 10545 2200 10575 2230
rect 10545 2180 10550 2200
rect 10570 2180 10575 2200
rect 10545 2150 10575 2180
rect 10545 2130 10550 2150
rect 10570 2130 10575 2150
rect 10545 2100 10575 2130
rect 10545 2080 10550 2100
rect 10570 2080 10575 2100
rect 10545 2050 10575 2080
rect 10545 2030 10550 2050
rect 10570 2030 10575 2050
rect 10545 2000 10575 2030
rect 10545 1980 10550 2000
rect 10570 1980 10575 2000
rect 10545 1970 10575 1980
rect 10600 2250 10630 2260
rect 10600 2230 10605 2250
rect 10625 2230 10630 2250
rect 10600 2200 10630 2230
rect 10600 2180 10605 2200
rect 10625 2180 10630 2200
rect 10600 2150 10630 2180
rect 10600 2130 10605 2150
rect 10625 2130 10630 2150
rect 10600 2100 10630 2130
rect 10600 2080 10605 2100
rect 10625 2080 10630 2100
rect 10600 2050 10630 2080
rect 10600 2030 10605 2050
rect 10625 2030 10630 2050
rect 10600 2000 10630 2030
rect 10600 1980 10605 2000
rect 10625 1980 10630 2000
rect 10600 1970 10630 1980
rect 10655 2250 10685 2260
rect 10655 2230 10660 2250
rect 10680 2230 10685 2250
rect 10655 2200 10685 2230
rect 10655 2180 10660 2200
rect 10680 2180 10685 2200
rect 10655 2150 10685 2180
rect 10655 2130 10660 2150
rect 10680 2130 10685 2150
rect 10655 2100 10685 2130
rect 10655 2080 10660 2100
rect 10680 2080 10685 2100
rect 10655 2050 10685 2080
rect 10655 2030 10660 2050
rect 10680 2030 10685 2050
rect 10655 2000 10685 2030
rect 10655 1980 10660 2000
rect 10680 1980 10685 2000
rect 10655 1970 10685 1980
rect 10710 2250 10740 2260
rect 10710 2230 10715 2250
rect 10735 2230 10740 2250
rect 10710 2200 10740 2230
rect 10710 2180 10715 2200
rect 10735 2180 10740 2200
rect 10710 2150 10740 2180
rect 10710 2130 10715 2150
rect 10735 2130 10740 2150
rect 10710 2100 10740 2130
rect 10710 2080 10715 2100
rect 10735 2080 10740 2100
rect 10710 2050 10740 2080
rect 10710 2030 10715 2050
rect 10735 2030 10740 2050
rect 10710 2000 10740 2030
rect 10710 1980 10715 2000
rect 10735 1980 10740 2000
rect 10710 1970 10740 1980
rect 10765 2250 10795 2260
rect 10765 2230 10770 2250
rect 10790 2230 10795 2250
rect 10765 2200 10795 2230
rect 10765 2180 10770 2200
rect 10790 2180 10795 2200
rect 10765 2150 10795 2180
rect 10765 2130 10770 2150
rect 10790 2130 10795 2150
rect 10765 2100 10795 2130
rect 10765 2080 10770 2100
rect 10790 2080 10795 2100
rect 10765 2050 10795 2080
rect 10765 2030 10770 2050
rect 10790 2030 10795 2050
rect 10765 2000 10795 2030
rect 10765 1980 10770 2000
rect 10790 1980 10795 2000
rect 10765 1970 10795 1980
rect 10820 2250 10890 2260
rect 10820 2230 10825 2250
rect 10845 2230 10865 2250
rect 10885 2230 10890 2250
rect 10820 2200 10890 2230
rect 10820 2180 10825 2200
rect 10845 2180 10865 2200
rect 10885 2180 10890 2200
rect 12910 2250 12980 2260
rect 12910 2230 12915 2250
rect 12935 2230 12955 2250
rect 12975 2230 12980 2250
rect 12910 2200 12980 2230
rect 10820 2150 10890 2180
rect 10820 2130 10825 2150
rect 10845 2130 10865 2150
rect 10885 2130 10890 2150
rect 11330 2175 11370 2185
rect 11330 2155 11340 2175
rect 11360 2155 11370 2175
rect 11330 2145 11370 2155
rect 11440 2175 11480 2185
rect 11440 2155 11450 2175
rect 11470 2155 11480 2175
rect 11440 2145 11480 2155
rect 11550 2175 11590 2185
rect 11550 2155 11560 2175
rect 11580 2155 11590 2175
rect 11550 2145 11590 2155
rect 11660 2175 11700 2185
rect 11660 2155 11670 2175
rect 11690 2155 11700 2175
rect 11660 2145 11700 2155
rect 11770 2175 11810 2185
rect 11770 2155 11780 2175
rect 11800 2155 11810 2175
rect 11770 2145 11810 2155
rect 11828 2175 11862 2185
rect 11828 2155 11836 2175
rect 11854 2155 11862 2175
rect 11828 2145 11862 2155
rect 11880 2175 11920 2185
rect 11880 2155 11890 2175
rect 11910 2155 11920 2175
rect 11880 2145 11920 2155
rect 11990 2175 12030 2185
rect 11990 2155 12000 2175
rect 12020 2155 12030 2175
rect 11990 2145 12030 2155
rect 12100 2175 12140 2185
rect 12100 2155 12110 2175
rect 12130 2155 12140 2175
rect 12100 2145 12140 2155
rect 12210 2175 12250 2185
rect 12210 2155 12220 2175
rect 12240 2155 12250 2175
rect 12210 2145 12250 2155
rect 12320 2175 12360 2185
rect 12320 2155 12330 2175
rect 12350 2155 12360 2175
rect 12320 2145 12360 2155
rect 12430 2175 12470 2185
rect 12430 2155 12440 2175
rect 12460 2155 12470 2175
rect 12430 2145 12470 2155
rect 12910 2180 12915 2200
rect 12935 2180 12955 2200
rect 12975 2180 12980 2200
rect 12910 2150 12980 2180
rect 10820 2100 10890 2130
rect 11340 2125 11360 2145
rect 11450 2125 11470 2145
rect 11560 2125 11580 2145
rect 11670 2125 11690 2145
rect 11780 2125 11800 2145
rect 11890 2125 11910 2145
rect 12000 2125 12020 2145
rect 12110 2125 12130 2145
rect 12220 2125 12240 2145
rect 12330 2125 12350 2145
rect 12440 2125 12460 2145
rect 12910 2130 12915 2150
rect 12935 2130 12955 2150
rect 12975 2130 12980 2150
rect 10820 2080 10825 2100
rect 10845 2080 10865 2100
rect 10885 2080 10890 2100
rect 10820 2050 10890 2080
rect 10820 2030 10825 2050
rect 10845 2030 10865 2050
rect 10885 2030 10890 2050
rect 10820 2000 10890 2030
rect 10820 1980 10825 2000
rect 10845 1980 10865 2000
rect 10885 1980 10890 2000
rect 11240 2115 11310 2125
rect 11240 2095 11245 2115
rect 11265 2095 11285 2115
rect 11305 2095 11310 2115
rect 11240 2065 11310 2095
rect 11240 2045 11245 2065
rect 11265 2045 11285 2065
rect 11305 2045 11310 2065
rect 11240 2015 11310 2045
rect 11240 1995 11245 2015
rect 11265 1995 11285 2015
rect 11305 1995 11310 2015
rect 11240 1985 11310 1995
rect 11335 2115 11365 2125
rect 11335 2095 11340 2115
rect 11360 2095 11365 2115
rect 11335 2065 11365 2095
rect 11335 2045 11340 2065
rect 11360 2045 11365 2065
rect 11335 2015 11365 2045
rect 11335 1995 11340 2015
rect 11360 1995 11365 2015
rect 11335 1985 11365 1995
rect 11390 2115 11420 2125
rect 11390 2095 11395 2115
rect 11415 2095 11420 2115
rect 11390 2065 11420 2095
rect 11390 2045 11395 2065
rect 11415 2045 11420 2065
rect 11390 2015 11420 2045
rect 11390 1995 11395 2015
rect 11415 1995 11420 2015
rect 11390 1985 11420 1995
rect 11445 2115 11475 2125
rect 11445 2095 11450 2115
rect 11470 2095 11475 2115
rect 11445 2065 11475 2095
rect 11445 2045 11450 2065
rect 11470 2045 11475 2065
rect 11445 2015 11475 2045
rect 11445 1995 11450 2015
rect 11470 1995 11475 2015
rect 11445 1985 11475 1995
rect 11500 2115 11530 2125
rect 11500 2095 11505 2115
rect 11525 2095 11530 2115
rect 11500 2065 11530 2095
rect 11500 2045 11505 2065
rect 11525 2045 11530 2065
rect 11500 2015 11530 2045
rect 11500 1995 11505 2015
rect 11525 1995 11530 2015
rect 11500 1985 11530 1995
rect 11555 2115 11585 2125
rect 11555 2095 11560 2115
rect 11580 2095 11585 2115
rect 11555 2065 11585 2095
rect 11555 2045 11560 2065
rect 11580 2045 11585 2065
rect 11555 2015 11585 2045
rect 11555 1995 11560 2015
rect 11580 1995 11585 2015
rect 11555 1985 11585 1995
rect 11610 2115 11640 2125
rect 11610 2095 11615 2115
rect 11635 2095 11640 2115
rect 11610 2065 11640 2095
rect 11610 2045 11615 2065
rect 11635 2045 11640 2065
rect 11610 2015 11640 2045
rect 11610 1995 11615 2015
rect 11635 1995 11640 2015
rect 11610 1985 11640 1995
rect 11665 2115 11695 2125
rect 11665 2095 11670 2115
rect 11690 2095 11695 2115
rect 11665 2065 11695 2095
rect 11665 2045 11670 2065
rect 11690 2045 11695 2065
rect 11665 2015 11695 2045
rect 11665 1995 11670 2015
rect 11690 1995 11695 2015
rect 11665 1985 11695 1995
rect 11720 2115 11750 2125
rect 11720 2095 11725 2115
rect 11745 2095 11750 2115
rect 11720 2065 11750 2095
rect 11720 2045 11725 2065
rect 11745 2045 11750 2065
rect 11720 2015 11750 2045
rect 11720 1995 11725 2015
rect 11745 1995 11750 2015
rect 11720 1985 11750 1995
rect 11775 2115 11805 2125
rect 11775 2095 11780 2115
rect 11800 2095 11805 2115
rect 11775 2065 11805 2095
rect 11775 2045 11780 2065
rect 11800 2045 11805 2065
rect 11775 2015 11805 2045
rect 11775 1995 11780 2015
rect 11800 1995 11805 2015
rect 11775 1985 11805 1995
rect 11830 2115 11860 2125
rect 11830 2095 11835 2115
rect 11855 2095 11860 2115
rect 11830 2065 11860 2095
rect 11830 2045 11835 2065
rect 11855 2045 11860 2065
rect 11830 2015 11860 2045
rect 11830 1995 11835 2015
rect 11855 1995 11860 2015
rect 11830 1985 11860 1995
rect 11885 2115 11915 2125
rect 11885 2095 11890 2115
rect 11910 2095 11915 2115
rect 11885 2065 11915 2095
rect 11885 2045 11890 2065
rect 11910 2045 11915 2065
rect 11885 2015 11915 2045
rect 11885 1995 11890 2015
rect 11910 1995 11915 2015
rect 11885 1985 11915 1995
rect 11940 2115 11970 2125
rect 11940 2095 11945 2115
rect 11965 2095 11970 2115
rect 11940 2065 11970 2095
rect 11940 2045 11945 2065
rect 11965 2045 11970 2065
rect 11940 2015 11970 2045
rect 11940 1995 11945 2015
rect 11965 1995 11970 2015
rect 11940 1985 11970 1995
rect 11995 2115 12025 2125
rect 11995 2095 12000 2115
rect 12020 2095 12025 2115
rect 11995 2065 12025 2095
rect 11995 2045 12000 2065
rect 12020 2045 12025 2065
rect 11995 2015 12025 2045
rect 11995 1995 12000 2015
rect 12020 1995 12025 2015
rect 11995 1985 12025 1995
rect 12050 2115 12080 2125
rect 12050 2095 12055 2115
rect 12075 2095 12080 2115
rect 12050 2065 12080 2095
rect 12050 2045 12055 2065
rect 12075 2045 12080 2065
rect 12050 2015 12080 2045
rect 12050 1995 12055 2015
rect 12075 1995 12080 2015
rect 12050 1985 12080 1995
rect 12105 2115 12135 2125
rect 12105 2095 12110 2115
rect 12130 2095 12135 2115
rect 12105 2065 12135 2095
rect 12105 2045 12110 2065
rect 12130 2045 12135 2065
rect 12105 2015 12135 2045
rect 12105 1995 12110 2015
rect 12130 1995 12135 2015
rect 12105 1985 12135 1995
rect 12160 2115 12190 2125
rect 12160 2095 12165 2115
rect 12185 2095 12190 2115
rect 12160 2065 12190 2095
rect 12160 2045 12165 2065
rect 12185 2045 12190 2065
rect 12160 2015 12190 2045
rect 12160 1995 12165 2015
rect 12185 1995 12190 2015
rect 12160 1985 12190 1995
rect 12215 2115 12245 2125
rect 12215 2095 12220 2115
rect 12240 2095 12245 2115
rect 12215 2065 12245 2095
rect 12215 2045 12220 2065
rect 12240 2045 12245 2065
rect 12215 2015 12245 2045
rect 12215 1995 12220 2015
rect 12240 1995 12245 2015
rect 12215 1985 12245 1995
rect 12270 2115 12300 2125
rect 12270 2095 12275 2115
rect 12295 2095 12300 2115
rect 12270 2065 12300 2095
rect 12270 2045 12275 2065
rect 12295 2045 12300 2065
rect 12270 2015 12300 2045
rect 12270 1995 12275 2015
rect 12295 1995 12300 2015
rect 12270 1985 12300 1995
rect 12325 2115 12355 2125
rect 12325 2095 12330 2115
rect 12350 2095 12355 2115
rect 12325 2065 12355 2095
rect 12325 2045 12330 2065
rect 12350 2045 12355 2065
rect 12325 2015 12355 2045
rect 12325 1995 12330 2015
rect 12350 1995 12355 2015
rect 12325 1985 12355 1995
rect 12380 2115 12410 2125
rect 12380 2095 12385 2115
rect 12405 2095 12410 2115
rect 12380 2065 12410 2095
rect 12380 2045 12385 2065
rect 12405 2045 12410 2065
rect 12380 2015 12410 2045
rect 12380 1995 12385 2015
rect 12405 1995 12410 2015
rect 12380 1985 12410 1995
rect 12435 2115 12465 2125
rect 12435 2095 12440 2115
rect 12460 2095 12465 2115
rect 12435 2065 12465 2095
rect 12435 2045 12440 2065
rect 12460 2045 12465 2065
rect 12435 2015 12465 2045
rect 12435 1995 12440 2015
rect 12460 1995 12465 2015
rect 12435 1985 12465 1995
rect 12490 2115 12560 2125
rect 12490 2095 12495 2115
rect 12515 2095 12535 2115
rect 12555 2095 12560 2115
rect 12490 2065 12560 2095
rect 12490 2045 12495 2065
rect 12515 2045 12535 2065
rect 12555 2045 12560 2065
rect 12490 2015 12560 2045
rect 12490 1995 12495 2015
rect 12515 1995 12535 2015
rect 12555 1995 12560 2015
rect 12490 1985 12560 1995
rect 12910 2100 12980 2130
rect 12910 2080 12915 2100
rect 12935 2080 12955 2100
rect 12975 2080 12980 2100
rect 12910 2050 12980 2080
rect 12910 2030 12915 2050
rect 12935 2030 12955 2050
rect 12975 2030 12980 2050
rect 12910 2000 12980 2030
rect 10820 1970 10890 1980
rect 5230 1935 5260 1965
rect 10220 1950 10240 1970
rect 10330 1950 10350 1970
rect 10440 1950 10460 1970
rect 10550 1950 10570 1970
rect 10660 1950 10680 1970
rect 10770 1950 10790 1970
rect 11245 1965 11265 1985
rect 11395 1965 11415 1985
rect 11505 1965 11525 1985
rect 11615 1965 11635 1985
rect 11725 1965 11745 1985
rect 11835 1965 11855 1985
rect 11945 1965 11965 1985
rect 12055 1965 12075 1985
rect 12165 1965 12185 1985
rect 12275 1965 12295 1985
rect 12385 1965 12405 1985
rect 12535 1965 12555 1985
rect 12910 1980 12915 2000
rect 12935 1980 12955 2000
rect 12975 1980 12980 2000
rect 12910 1970 12980 1980
rect 13005 2250 13035 2260
rect 13005 2230 13010 2250
rect 13030 2230 13035 2250
rect 13005 2200 13035 2230
rect 13005 2180 13010 2200
rect 13030 2180 13035 2200
rect 13005 2150 13035 2180
rect 13005 2130 13010 2150
rect 13030 2130 13035 2150
rect 13005 2100 13035 2130
rect 13005 2080 13010 2100
rect 13030 2080 13035 2100
rect 13005 2050 13035 2080
rect 13005 2030 13010 2050
rect 13030 2030 13035 2050
rect 13005 2000 13035 2030
rect 13005 1980 13010 2000
rect 13030 1980 13035 2000
rect 13005 1970 13035 1980
rect 13060 2250 13090 2260
rect 13060 2230 13065 2250
rect 13085 2230 13090 2250
rect 13060 2200 13090 2230
rect 13060 2180 13065 2200
rect 13085 2180 13090 2200
rect 13060 2150 13090 2180
rect 13060 2130 13065 2150
rect 13085 2130 13090 2150
rect 13060 2100 13090 2130
rect 13060 2080 13065 2100
rect 13085 2080 13090 2100
rect 13060 2050 13090 2080
rect 13060 2030 13065 2050
rect 13085 2030 13090 2050
rect 13060 2000 13090 2030
rect 13060 1980 13065 2000
rect 13085 1980 13090 2000
rect 13060 1970 13090 1980
rect 13115 2250 13145 2260
rect 13115 2230 13120 2250
rect 13140 2230 13145 2250
rect 13115 2200 13145 2230
rect 13115 2180 13120 2200
rect 13140 2180 13145 2200
rect 13115 2150 13145 2180
rect 13115 2130 13120 2150
rect 13140 2130 13145 2150
rect 13115 2100 13145 2130
rect 13115 2080 13120 2100
rect 13140 2080 13145 2100
rect 13115 2050 13145 2080
rect 13115 2030 13120 2050
rect 13140 2030 13145 2050
rect 13115 2000 13145 2030
rect 13115 1980 13120 2000
rect 13140 1980 13145 2000
rect 13115 1970 13145 1980
rect 13170 2250 13200 2260
rect 13170 2230 13175 2250
rect 13195 2230 13200 2250
rect 13170 2200 13200 2230
rect 13170 2180 13175 2200
rect 13195 2180 13200 2200
rect 13170 2150 13200 2180
rect 13170 2130 13175 2150
rect 13195 2130 13200 2150
rect 13170 2100 13200 2130
rect 13170 2080 13175 2100
rect 13195 2080 13200 2100
rect 13170 2050 13200 2080
rect 13170 2030 13175 2050
rect 13195 2030 13200 2050
rect 13170 2000 13200 2030
rect 13170 1980 13175 2000
rect 13195 1980 13200 2000
rect 13170 1970 13200 1980
rect 13225 2250 13255 2260
rect 13225 2230 13230 2250
rect 13250 2230 13255 2250
rect 13225 2200 13255 2230
rect 13225 2180 13230 2200
rect 13250 2180 13255 2200
rect 13225 2150 13255 2180
rect 13225 2130 13230 2150
rect 13250 2130 13255 2150
rect 13225 2100 13255 2130
rect 13225 2080 13230 2100
rect 13250 2080 13255 2100
rect 13225 2050 13255 2080
rect 13225 2030 13230 2050
rect 13250 2030 13255 2050
rect 13225 2000 13255 2030
rect 13225 1980 13230 2000
rect 13250 1980 13255 2000
rect 13225 1970 13255 1980
rect 13280 2250 13310 2260
rect 13280 2230 13285 2250
rect 13305 2230 13310 2250
rect 13280 2200 13310 2230
rect 13280 2180 13285 2200
rect 13305 2180 13310 2200
rect 13280 2150 13310 2180
rect 13280 2130 13285 2150
rect 13305 2130 13310 2150
rect 13280 2100 13310 2130
rect 13280 2080 13285 2100
rect 13305 2080 13310 2100
rect 13280 2050 13310 2080
rect 13280 2030 13285 2050
rect 13305 2030 13310 2050
rect 13280 2000 13310 2030
rect 13280 1980 13285 2000
rect 13305 1980 13310 2000
rect 13280 1970 13310 1980
rect 13335 2250 13365 2260
rect 13335 2230 13340 2250
rect 13360 2230 13365 2250
rect 13335 2200 13365 2230
rect 13335 2180 13340 2200
rect 13360 2180 13365 2200
rect 13335 2150 13365 2180
rect 13335 2130 13340 2150
rect 13360 2130 13365 2150
rect 13335 2100 13365 2130
rect 13335 2080 13340 2100
rect 13360 2080 13365 2100
rect 13335 2050 13365 2080
rect 13335 2030 13340 2050
rect 13360 2030 13365 2050
rect 13335 2000 13365 2030
rect 13335 1980 13340 2000
rect 13360 1980 13365 2000
rect 13335 1970 13365 1980
rect 13390 2250 13420 2260
rect 13390 2230 13395 2250
rect 13415 2230 13420 2250
rect 13390 2200 13420 2230
rect 13390 2180 13395 2200
rect 13415 2180 13420 2200
rect 13390 2150 13420 2180
rect 13390 2130 13395 2150
rect 13415 2130 13420 2150
rect 13390 2100 13420 2130
rect 13390 2080 13395 2100
rect 13415 2080 13420 2100
rect 13390 2050 13420 2080
rect 13390 2030 13395 2050
rect 13415 2030 13420 2050
rect 13390 2000 13420 2030
rect 13390 1980 13395 2000
rect 13415 1980 13420 2000
rect 13390 1970 13420 1980
rect 13445 2250 13475 2260
rect 13445 2230 13450 2250
rect 13470 2230 13475 2250
rect 13445 2200 13475 2230
rect 13445 2180 13450 2200
rect 13470 2180 13475 2200
rect 13445 2150 13475 2180
rect 13445 2130 13450 2150
rect 13470 2130 13475 2150
rect 13445 2100 13475 2130
rect 13445 2080 13450 2100
rect 13470 2080 13475 2100
rect 13445 2050 13475 2080
rect 13445 2030 13450 2050
rect 13470 2030 13475 2050
rect 13445 2000 13475 2030
rect 13445 1980 13450 2000
rect 13470 1980 13475 2000
rect 13445 1970 13475 1980
rect 13500 2250 13530 2260
rect 13500 2230 13505 2250
rect 13525 2230 13530 2250
rect 13500 2200 13530 2230
rect 13500 2180 13505 2200
rect 13525 2180 13530 2200
rect 13500 2150 13530 2180
rect 13500 2130 13505 2150
rect 13525 2130 13530 2150
rect 13500 2100 13530 2130
rect 13500 2080 13505 2100
rect 13525 2080 13530 2100
rect 13500 2050 13530 2080
rect 13500 2030 13505 2050
rect 13525 2030 13530 2050
rect 13500 2000 13530 2030
rect 13500 1980 13505 2000
rect 13525 1980 13530 2000
rect 13500 1970 13530 1980
rect 13555 2250 13585 2260
rect 13555 2230 13560 2250
rect 13580 2230 13585 2250
rect 13555 2200 13585 2230
rect 13555 2180 13560 2200
rect 13580 2180 13585 2200
rect 13555 2150 13585 2180
rect 13555 2130 13560 2150
rect 13580 2130 13585 2150
rect 13555 2100 13585 2130
rect 13555 2080 13560 2100
rect 13580 2080 13585 2100
rect 13555 2050 13585 2080
rect 13555 2030 13560 2050
rect 13580 2030 13585 2050
rect 13555 2000 13585 2030
rect 13555 1980 13560 2000
rect 13580 1980 13585 2000
rect 13555 1970 13585 1980
rect 13610 2250 13680 2260
rect 13610 2230 13615 2250
rect 13635 2230 13655 2250
rect 13675 2230 13680 2250
rect 25813 2255 25821 2275
rect 25839 2255 25847 2275
rect 25813 2245 25847 2255
rect 27973 2275 28007 2285
rect 27973 2255 27981 2275
rect 27999 2255 28007 2275
rect 27973 2245 28007 2255
rect 13610 2200 13680 2230
rect 13610 2180 13615 2200
rect 13635 2180 13655 2200
rect 13675 2180 13680 2200
rect 13610 2150 13680 2180
rect 13610 2130 13615 2150
rect 13635 2130 13655 2150
rect 13675 2130 13680 2150
rect 13610 2100 13680 2130
rect 13610 2080 13615 2100
rect 13635 2080 13655 2100
rect 13675 2080 13680 2100
rect 13610 2050 13680 2080
rect 13610 2030 13615 2050
rect 13635 2030 13655 2050
rect 13675 2030 13680 2050
rect 13610 2000 13680 2030
rect 13610 1980 13615 2000
rect 13635 1980 13655 2000
rect 13675 1980 13680 2000
rect 13610 1970 13680 1980
rect 13795 2000 13830 2010
rect 13795 1975 13800 2000
rect 13825 1975 13830 2000
rect 11235 1955 11275 1965
rect 5230 1915 5235 1935
rect 5255 1915 5260 1935
rect 5230 1905 5260 1915
rect 10210 1940 10250 1950
rect 10210 1920 10220 1940
rect 10238 1920 10250 1940
rect 10210 1910 10250 1920
rect 10320 1940 10360 1950
rect 10320 1920 10330 1940
rect 10348 1920 10360 1940
rect 10320 1910 10360 1920
rect 10430 1940 10470 1950
rect 10430 1920 10440 1940
rect 10458 1920 10470 1940
rect 10430 1910 10470 1920
rect 10540 1940 10580 1950
rect 10540 1920 10550 1940
rect 10568 1920 10580 1940
rect 10540 1910 10580 1920
rect 10650 1940 10690 1950
rect 10650 1920 10660 1940
rect 10678 1920 10690 1940
rect 10650 1910 10690 1920
rect 10760 1940 10800 1950
rect 10760 1920 10770 1940
rect 10788 1920 10800 1940
rect 11235 1935 11245 1955
rect 11265 1935 11275 1955
rect 11235 1925 11275 1935
rect 11385 1955 11425 1965
rect 11385 1935 11395 1955
rect 11415 1935 11425 1955
rect 11385 1925 11425 1935
rect 11495 1955 11535 1965
rect 11495 1935 11505 1955
rect 11525 1935 11535 1955
rect 11495 1925 11535 1935
rect 11605 1955 11645 1965
rect 11605 1935 11615 1955
rect 11635 1935 11645 1955
rect 11605 1925 11645 1935
rect 11715 1955 11755 1965
rect 11715 1935 11725 1955
rect 11745 1935 11755 1955
rect 11715 1925 11755 1935
rect 11825 1955 11865 1965
rect 11825 1935 11835 1955
rect 11855 1935 11865 1955
rect 11825 1925 11865 1935
rect 11935 1955 11975 1965
rect 11935 1935 11945 1955
rect 11965 1935 11975 1955
rect 11935 1925 11975 1935
rect 12045 1955 12085 1965
rect 12045 1935 12055 1955
rect 12075 1935 12085 1955
rect 12045 1925 12085 1935
rect 12155 1955 12195 1965
rect 12155 1935 12165 1955
rect 12185 1935 12195 1955
rect 12155 1925 12195 1935
rect 12265 1955 12305 1965
rect 12265 1935 12275 1955
rect 12295 1935 12305 1955
rect 12265 1925 12305 1935
rect 12375 1955 12415 1965
rect 12375 1935 12385 1955
rect 12405 1935 12415 1955
rect 12375 1925 12415 1935
rect 12525 1955 12565 1965
rect 12525 1935 12535 1955
rect 12555 1935 12565 1955
rect 13010 1950 13030 1970
rect 13120 1950 13140 1970
rect 13230 1950 13250 1970
rect 13340 1950 13360 1970
rect 13450 1950 13470 1970
rect 13560 1950 13580 1970
rect 13795 1965 13830 1975
rect 13855 2000 13890 2010
rect 13855 1975 13860 2000
rect 13885 1975 13890 2000
rect 13855 1965 13890 1975
rect 13915 2000 13950 2010
rect 13915 1975 13920 2000
rect 13945 1975 13950 2000
rect 13915 1965 13950 1975
rect 24640 2215 24680 2225
rect 24640 2195 24650 2215
rect 24670 2195 24680 2215
rect 24640 2185 24680 2195
rect 24790 2215 24830 2225
rect 24790 2195 24800 2215
rect 24820 2195 24830 2215
rect 24790 2185 24830 2195
rect 24900 2215 24940 2225
rect 24900 2195 24910 2215
rect 24930 2195 24940 2215
rect 24900 2185 24940 2195
rect 25010 2215 25050 2225
rect 25010 2195 25020 2215
rect 25040 2195 25050 2215
rect 25010 2185 25050 2195
rect 25120 2215 25160 2225
rect 25120 2195 25130 2215
rect 25150 2195 25160 2215
rect 25120 2185 25160 2195
rect 25230 2215 25270 2225
rect 25230 2195 25240 2215
rect 25260 2195 25270 2215
rect 25230 2185 25270 2195
rect 25340 2215 25380 2225
rect 25340 2195 25350 2215
rect 25370 2195 25380 2215
rect 25340 2185 25380 2195
rect 25450 2215 25490 2225
rect 25450 2195 25460 2215
rect 25480 2195 25490 2215
rect 25450 2185 25490 2195
rect 25560 2215 25600 2225
rect 25560 2195 25570 2215
rect 25590 2195 25600 2215
rect 25560 2185 25600 2195
rect 25670 2215 25710 2225
rect 25670 2195 25680 2215
rect 25700 2195 25710 2215
rect 25670 2185 25710 2195
rect 25780 2215 25820 2225
rect 25780 2195 25790 2215
rect 25810 2195 25820 2215
rect 25780 2185 25820 2195
rect 25930 2215 25970 2225
rect 25930 2195 25940 2215
rect 25960 2195 25970 2215
rect 25930 2185 25970 2195
rect 27850 2215 27890 2225
rect 27850 2195 27860 2215
rect 27880 2195 27890 2215
rect 27850 2185 27890 2195
rect 28000 2215 28040 2225
rect 28000 2195 28010 2215
rect 28030 2195 28040 2215
rect 28000 2185 28040 2195
rect 28110 2215 28150 2225
rect 28110 2195 28120 2215
rect 28140 2195 28150 2215
rect 28110 2185 28150 2195
rect 28220 2215 28260 2225
rect 28220 2195 28230 2215
rect 28250 2195 28260 2215
rect 28220 2185 28260 2195
rect 28330 2215 28370 2225
rect 28330 2195 28340 2215
rect 28360 2195 28370 2215
rect 28330 2185 28370 2195
rect 28440 2215 28480 2225
rect 28440 2195 28450 2215
rect 28470 2195 28480 2215
rect 28440 2185 28480 2195
rect 28550 2215 28590 2225
rect 28550 2195 28560 2215
rect 28580 2195 28590 2215
rect 28550 2185 28590 2195
rect 28660 2215 28700 2225
rect 28660 2195 28670 2215
rect 28690 2195 28700 2215
rect 28660 2185 28700 2195
rect 28770 2215 28810 2225
rect 28770 2195 28780 2215
rect 28800 2195 28810 2215
rect 28770 2185 28810 2195
rect 28880 2215 28920 2225
rect 28880 2195 28890 2215
rect 28910 2195 28920 2215
rect 28880 2185 28920 2195
rect 28990 2215 29030 2225
rect 28990 2195 29000 2215
rect 29020 2195 29030 2215
rect 28990 2185 29030 2195
rect 29140 2215 29180 2225
rect 29140 2195 29150 2215
rect 29170 2195 29180 2215
rect 29140 2185 29180 2195
rect 24650 2165 24670 2185
rect 24800 2165 24820 2185
rect 24910 2165 24930 2185
rect 25020 2165 25040 2185
rect 25130 2165 25150 2185
rect 25240 2165 25260 2185
rect 25350 2165 25370 2185
rect 25460 2165 25480 2185
rect 25570 2165 25590 2185
rect 25680 2165 25700 2185
rect 25790 2165 25810 2185
rect 25940 2165 25960 2185
rect 26330 2175 26370 2185
rect 24645 2155 24715 2165
rect 24645 2135 24650 2155
rect 24670 2135 24690 2155
rect 24710 2135 24715 2155
rect 24645 2105 24715 2135
rect 24645 2085 24650 2105
rect 24670 2085 24690 2105
rect 24710 2085 24715 2105
rect 24645 2055 24715 2085
rect 24645 2035 24650 2055
rect 24670 2035 24690 2055
rect 24710 2035 24715 2055
rect 24645 2025 24715 2035
rect 24740 2155 24770 2165
rect 24740 2135 24745 2155
rect 24765 2135 24770 2155
rect 24740 2105 24770 2135
rect 24740 2085 24745 2105
rect 24765 2085 24770 2105
rect 24740 2055 24770 2085
rect 24740 2035 24745 2055
rect 24765 2035 24770 2055
rect 24740 2025 24770 2035
rect 24795 2155 24825 2165
rect 24795 2135 24800 2155
rect 24820 2135 24825 2155
rect 24795 2105 24825 2135
rect 24795 2085 24800 2105
rect 24820 2085 24825 2105
rect 24795 2055 24825 2085
rect 24795 2035 24800 2055
rect 24820 2035 24825 2055
rect 24795 2025 24825 2035
rect 24850 2155 24880 2165
rect 24850 2135 24855 2155
rect 24875 2135 24880 2155
rect 24850 2105 24880 2135
rect 24850 2085 24855 2105
rect 24875 2085 24880 2105
rect 24850 2055 24880 2085
rect 24850 2035 24855 2055
rect 24875 2035 24880 2055
rect 24850 2025 24880 2035
rect 24905 2155 24935 2165
rect 24905 2135 24910 2155
rect 24930 2135 24935 2155
rect 24905 2105 24935 2135
rect 24905 2085 24910 2105
rect 24930 2085 24935 2105
rect 24905 2055 24935 2085
rect 24905 2035 24910 2055
rect 24930 2035 24935 2055
rect 24905 2025 24935 2035
rect 24960 2155 24990 2165
rect 24960 2135 24965 2155
rect 24985 2135 24990 2155
rect 24960 2105 24990 2135
rect 24960 2085 24965 2105
rect 24985 2085 24990 2105
rect 24960 2055 24990 2085
rect 24960 2035 24965 2055
rect 24985 2035 24990 2055
rect 24960 2025 24990 2035
rect 25015 2155 25045 2165
rect 25015 2135 25020 2155
rect 25040 2135 25045 2155
rect 25015 2105 25045 2135
rect 25015 2085 25020 2105
rect 25040 2085 25045 2105
rect 25015 2055 25045 2085
rect 25015 2035 25020 2055
rect 25040 2035 25045 2055
rect 25015 2025 25045 2035
rect 25070 2155 25100 2165
rect 25070 2135 25075 2155
rect 25095 2135 25100 2155
rect 25070 2105 25100 2135
rect 25070 2085 25075 2105
rect 25095 2085 25100 2105
rect 25070 2055 25100 2085
rect 25070 2035 25075 2055
rect 25095 2035 25100 2055
rect 25070 2025 25100 2035
rect 25125 2155 25155 2165
rect 25125 2135 25130 2155
rect 25150 2135 25155 2155
rect 25125 2105 25155 2135
rect 25125 2085 25130 2105
rect 25150 2085 25155 2105
rect 25125 2055 25155 2085
rect 25125 2035 25130 2055
rect 25150 2035 25155 2055
rect 25125 2025 25155 2035
rect 25180 2155 25210 2165
rect 25180 2135 25185 2155
rect 25205 2135 25210 2155
rect 25180 2105 25210 2135
rect 25180 2085 25185 2105
rect 25205 2085 25210 2105
rect 25180 2055 25210 2085
rect 25180 2035 25185 2055
rect 25205 2035 25210 2055
rect 25180 2025 25210 2035
rect 25235 2155 25265 2165
rect 25235 2135 25240 2155
rect 25260 2135 25265 2155
rect 25235 2105 25265 2135
rect 25235 2085 25240 2105
rect 25260 2085 25265 2105
rect 25235 2055 25265 2085
rect 25235 2035 25240 2055
rect 25260 2035 25265 2055
rect 25235 2025 25265 2035
rect 25290 2155 25320 2165
rect 25290 2135 25295 2155
rect 25315 2135 25320 2155
rect 25290 2105 25320 2135
rect 25290 2085 25295 2105
rect 25315 2085 25320 2105
rect 25290 2055 25320 2085
rect 25290 2035 25295 2055
rect 25315 2035 25320 2055
rect 25290 2025 25320 2035
rect 25345 2155 25375 2165
rect 25345 2135 25350 2155
rect 25370 2135 25375 2155
rect 25345 2105 25375 2135
rect 25345 2085 25350 2105
rect 25370 2085 25375 2105
rect 25345 2055 25375 2085
rect 25345 2035 25350 2055
rect 25370 2035 25375 2055
rect 25345 2025 25375 2035
rect 25400 2155 25430 2165
rect 25400 2135 25405 2155
rect 25425 2135 25430 2155
rect 25400 2105 25430 2135
rect 25400 2085 25405 2105
rect 25425 2085 25430 2105
rect 25400 2055 25430 2085
rect 25400 2035 25405 2055
rect 25425 2035 25430 2055
rect 25400 2025 25430 2035
rect 25455 2155 25485 2165
rect 25455 2135 25460 2155
rect 25480 2135 25485 2155
rect 25455 2105 25485 2135
rect 25455 2085 25460 2105
rect 25480 2085 25485 2105
rect 25455 2055 25485 2085
rect 25455 2035 25460 2055
rect 25480 2035 25485 2055
rect 25455 2025 25485 2035
rect 25510 2155 25540 2165
rect 25510 2135 25515 2155
rect 25535 2135 25540 2155
rect 25510 2105 25540 2135
rect 25510 2085 25515 2105
rect 25535 2085 25540 2105
rect 25510 2055 25540 2085
rect 25510 2035 25515 2055
rect 25535 2035 25540 2055
rect 25510 2025 25540 2035
rect 25565 2155 25595 2165
rect 25565 2135 25570 2155
rect 25590 2135 25595 2155
rect 25565 2105 25595 2135
rect 25565 2085 25570 2105
rect 25590 2085 25595 2105
rect 25565 2055 25595 2085
rect 25565 2035 25570 2055
rect 25590 2035 25595 2055
rect 25565 2025 25595 2035
rect 25620 2155 25650 2165
rect 25620 2135 25625 2155
rect 25645 2135 25650 2155
rect 25620 2105 25650 2135
rect 25620 2085 25625 2105
rect 25645 2085 25650 2105
rect 25620 2055 25650 2085
rect 25620 2035 25625 2055
rect 25645 2035 25650 2055
rect 25620 2025 25650 2035
rect 25675 2155 25705 2165
rect 25675 2135 25680 2155
rect 25700 2135 25705 2155
rect 25675 2105 25705 2135
rect 25675 2085 25680 2105
rect 25700 2085 25705 2105
rect 25675 2055 25705 2085
rect 25675 2035 25680 2055
rect 25700 2035 25705 2055
rect 25675 2025 25705 2035
rect 25730 2155 25760 2165
rect 25730 2135 25735 2155
rect 25755 2135 25760 2155
rect 25730 2105 25760 2135
rect 25730 2085 25735 2105
rect 25755 2085 25760 2105
rect 25730 2055 25760 2085
rect 25730 2035 25735 2055
rect 25755 2035 25760 2055
rect 25730 2025 25760 2035
rect 25785 2155 25815 2165
rect 25785 2135 25790 2155
rect 25810 2135 25815 2155
rect 25785 2105 25815 2135
rect 25785 2085 25790 2105
rect 25810 2085 25815 2105
rect 25785 2055 25815 2085
rect 25785 2035 25790 2055
rect 25810 2035 25815 2055
rect 25785 2025 25815 2035
rect 25840 2155 25870 2165
rect 25840 2135 25845 2155
rect 25865 2135 25870 2155
rect 25840 2105 25870 2135
rect 25840 2085 25845 2105
rect 25865 2085 25870 2105
rect 25840 2055 25870 2085
rect 25840 2035 25845 2055
rect 25865 2035 25870 2055
rect 25840 2025 25870 2035
rect 25895 2155 25965 2165
rect 25895 2135 25900 2155
rect 25920 2135 25940 2155
rect 25960 2135 25965 2155
rect 26330 2155 26340 2175
rect 26360 2155 26370 2175
rect 26330 2145 26370 2155
rect 26440 2175 26480 2185
rect 26440 2155 26450 2175
rect 26470 2155 26480 2175
rect 26440 2145 26480 2155
rect 26550 2175 26590 2185
rect 26550 2155 26560 2175
rect 26580 2155 26590 2175
rect 26550 2145 26590 2155
rect 26660 2175 26700 2185
rect 26660 2155 26670 2175
rect 26690 2155 26700 2175
rect 26660 2145 26700 2155
rect 26770 2175 26810 2185
rect 26770 2155 26780 2175
rect 26800 2155 26810 2175
rect 26770 2145 26810 2155
rect 26880 2175 26920 2185
rect 26880 2155 26890 2175
rect 26910 2155 26920 2175
rect 26880 2145 26920 2155
rect 26990 2175 27030 2185
rect 26990 2155 27000 2175
rect 27020 2155 27030 2175
rect 26990 2145 27030 2155
rect 27100 2175 27140 2185
rect 27100 2155 27110 2175
rect 27130 2155 27140 2175
rect 27100 2145 27140 2155
rect 27210 2175 27250 2185
rect 27210 2155 27220 2175
rect 27240 2155 27250 2175
rect 27210 2145 27250 2155
rect 27320 2175 27360 2185
rect 27320 2155 27330 2175
rect 27350 2155 27360 2175
rect 27320 2145 27360 2155
rect 27430 2175 27470 2185
rect 27430 2155 27440 2175
rect 27460 2155 27470 2175
rect 27860 2165 27880 2185
rect 28010 2165 28030 2185
rect 28120 2165 28140 2185
rect 28230 2165 28250 2185
rect 28340 2165 28360 2185
rect 28450 2165 28470 2185
rect 28560 2165 28580 2185
rect 28670 2165 28690 2185
rect 28780 2165 28800 2185
rect 28890 2165 28910 2185
rect 29000 2165 29020 2185
rect 29150 2165 29170 2185
rect 27430 2145 27470 2155
rect 27855 2155 27925 2165
rect 25895 2105 25965 2135
rect 26340 2125 26360 2145
rect 26450 2125 26470 2145
rect 26560 2125 26580 2145
rect 26670 2125 26690 2145
rect 26780 2125 26800 2145
rect 26890 2125 26910 2145
rect 27000 2125 27020 2145
rect 27110 2125 27130 2145
rect 27220 2125 27240 2145
rect 27330 2125 27350 2145
rect 27440 2125 27460 2145
rect 27855 2135 27860 2155
rect 27880 2135 27900 2155
rect 27920 2135 27925 2155
rect 25895 2085 25900 2105
rect 25920 2085 25940 2105
rect 25960 2085 25965 2105
rect 25895 2055 25965 2085
rect 25895 2035 25900 2055
rect 25920 2035 25940 2055
rect 25960 2035 25965 2055
rect 25895 2025 25965 2035
rect 26240 2115 26310 2125
rect 26240 2095 26245 2115
rect 26265 2095 26285 2115
rect 26305 2095 26310 2115
rect 26240 2065 26310 2095
rect 26240 2045 26245 2065
rect 26265 2045 26285 2065
rect 26305 2045 26310 2065
rect 13975 2000 14010 2010
rect 24745 2005 24765 2025
rect 24855 2005 24875 2025
rect 24965 2005 24985 2025
rect 25075 2005 25095 2025
rect 25185 2005 25205 2025
rect 25295 2005 25315 2025
rect 25405 2005 25425 2025
rect 25515 2005 25535 2025
rect 25625 2005 25645 2025
rect 25735 2005 25755 2025
rect 25845 2005 25865 2025
rect 26240 2015 26310 2045
rect 13975 1975 13980 2000
rect 14005 1975 14010 2000
rect 13975 1965 14010 1975
rect 24735 1995 24775 2005
rect 24735 1975 24745 1995
rect 24763 1975 24775 1995
rect 24735 1965 24775 1975
rect 24845 1995 24885 2005
rect 24845 1975 24855 1995
rect 24873 1975 24885 1995
rect 24845 1965 24885 1975
rect 24955 1995 24995 2005
rect 24955 1975 24965 1995
rect 24983 1975 24995 1995
rect 24955 1965 24995 1975
rect 25065 1995 25105 2005
rect 25065 1975 25075 1995
rect 25093 1975 25105 1995
rect 25065 1965 25105 1975
rect 25175 1995 25215 2005
rect 25175 1975 25185 1995
rect 25203 1975 25215 1995
rect 25175 1965 25215 1975
rect 25285 1995 25325 2005
rect 25285 1975 25295 1995
rect 25313 1975 25325 1995
rect 25285 1965 25325 1975
rect 25395 1995 25435 2005
rect 25395 1975 25405 1995
rect 25423 1975 25435 1995
rect 25395 1965 25435 1975
rect 25505 1995 25545 2005
rect 25505 1975 25515 1995
rect 25533 1975 25545 1995
rect 25505 1965 25545 1975
rect 25615 1995 25655 2005
rect 25615 1975 25625 1995
rect 25643 1975 25655 1995
rect 25615 1965 25655 1975
rect 25725 1995 25765 2005
rect 25725 1975 25735 1995
rect 25753 1975 25765 1995
rect 25725 1965 25765 1975
rect 25835 1995 25875 2005
rect 25835 1975 25845 1995
rect 25863 1975 25875 1995
rect 26240 1995 26245 2015
rect 26265 1995 26285 2015
rect 26305 1995 26310 2015
rect 26240 1985 26310 1995
rect 26335 2115 26365 2125
rect 26335 2095 26340 2115
rect 26360 2095 26365 2115
rect 26335 2065 26365 2095
rect 26335 2045 26340 2065
rect 26360 2045 26365 2065
rect 26335 2015 26365 2045
rect 26335 1995 26340 2015
rect 26360 1995 26365 2015
rect 26335 1985 26365 1995
rect 26390 2115 26420 2125
rect 26390 2095 26395 2115
rect 26415 2095 26420 2115
rect 26390 2065 26420 2095
rect 26390 2045 26395 2065
rect 26415 2045 26420 2065
rect 26390 2015 26420 2045
rect 26390 1995 26395 2015
rect 26415 1995 26420 2015
rect 26390 1985 26420 1995
rect 26445 2115 26475 2125
rect 26445 2095 26450 2115
rect 26470 2095 26475 2115
rect 26445 2065 26475 2095
rect 26445 2045 26450 2065
rect 26470 2045 26475 2065
rect 26445 2015 26475 2045
rect 26445 1995 26450 2015
rect 26470 1995 26475 2015
rect 26445 1985 26475 1995
rect 26500 2115 26530 2125
rect 26500 2095 26505 2115
rect 26525 2095 26530 2115
rect 26500 2065 26530 2095
rect 26500 2045 26505 2065
rect 26525 2045 26530 2065
rect 26500 2015 26530 2045
rect 26500 1995 26505 2015
rect 26525 1995 26530 2015
rect 26500 1985 26530 1995
rect 26555 2115 26585 2125
rect 26555 2095 26560 2115
rect 26580 2095 26585 2115
rect 26555 2065 26585 2095
rect 26555 2045 26560 2065
rect 26580 2045 26585 2065
rect 26555 2015 26585 2045
rect 26555 1995 26560 2015
rect 26580 1995 26585 2015
rect 26555 1985 26585 1995
rect 26610 2115 26640 2125
rect 26610 2095 26615 2115
rect 26635 2095 26640 2115
rect 26610 2065 26640 2095
rect 26610 2045 26615 2065
rect 26635 2045 26640 2065
rect 26610 2015 26640 2045
rect 26610 1995 26615 2015
rect 26635 1995 26640 2015
rect 26610 1985 26640 1995
rect 26665 2115 26695 2125
rect 26665 2095 26670 2115
rect 26690 2095 26695 2115
rect 26665 2065 26695 2095
rect 26665 2045 26670 2065
rect 26690 2045 26695 2065
rect 26665 2015 26695 2045
rect 26665 1995 26670 2015
rect 26690 1995 26695 2015
rect 26665 1985 26695 1995
rect 26720 2115 26750 2125
rect 26720 2095 26725 2115
rect 26745 2095 26750 2115
rect 26720 2065 26750 2095
rect 26720 2045 26725 2065
rect 26745 2045 26750 2065
rect 26720 2015 26750 2045
rect 26720 1995 26725 2015
rect 26745 1995 26750 2015
rect 26720 1985 26750 1995
rect 26775 2115 26805 2125
rect 26775 2095 26780 2115
rect 26800 2095 26805 2115
rect 26775 2065 26805 2095
rect 26775 2045 26780 2065
rect 26800 2045 26805 2065
rect 26775 2015 26805 2045
rect 26775 1995 26780 2015
rect 26800 1995 26805 2015
rect 26775 1985 26805 1995
rect 26830 2115 26860 2125
rect 26830 2095 26835 2115
rect 26855 2095 26860 2115
rect 26830 2065 26860 2095
rect 26830 2045 26835 2065
rect 26855 2045 26860 2065
rect 26830 2015 26860 2045
rect 26830 1995 26835 2015
rect 26855 1995 26860 2015
rect 26830 1985 26860 1995
rect 26885 2115 26915 2125
rect 26885 2095 26890 2115
rect 26910 2095 26915 2115
rect 26885 2065 26915 2095
rect 26885 2045 26890 2065
rect 26910 2045 26915 2065
rect 26885 2015 26915 2045
rect 26885 1995 26890 2015
rect 26910 1995 26915 2015
rect 26885 1985 26915 1995
rect 26940 2115 26970 2125
rect 26940 2095 26945 2115
rect 26965 2095 26970 2115
rect 26940 2065 26970 2095
rect 26940 2045 26945 2065
rect 26965 2045 26970 2065
rect 26940 2015 26970 2045
rect 26940 1995 26945 2015
rect 26965 1995 26970 2015
rect 26940 1985 26970 1995
rect 26995 2115 27025 2125
rect 26995 2095 27000 2115
rect 27020 2095 27025 2115
rect 26995 2065 27025 2095
rect 26995 2045 27000 2065
rect 27020 2045 27025 2065
rect 26995 2015 27025 2045
rect 26995 1995 27000 2015
rect 27020 1995 27025 2015
rect 26995 1985 27025 1995
rect 27050 2115 27080 2125
rect 27050 2095 27055 2115
rect 27075 2095 27080 2115
rect 27050 2065 27080 2095
rect 27050 2045 27055 2065
rect 27075 2045 27080 2065
rect 27050 2015 27080 2045
rect 27050 1995 27055 2015
rect 27075 1995 27080 2015
rect 27050 1985 27080 1995
rect 27105 2115 27135 2125
rect 27105 2095 27110 2115
rect 27130 2095 27135 2115
rect 27105 2065 27135 2095
rect 27105 2045 27110 2065
rect 27130 2045 27135 2065
rect 27105 2015 27135 2045
rect 27105 1995 27110 2015
rect 27130 1995 27135 2015
rect 27105 1985 27135 1995
rect 27160 2115 27190 2125
rect 27160 2095 27165 2115
rect 27185 2095 27190 2115
rect 27160 2065 27190 2095
rect 27160 2045 27165 2065
rect 27185 2045 27190 2065
rect 27160 2015 27190 2045
rect 27160 1995 27165 2015
rect 27185 1995 27190 2015
rect 27160 1985 27190 1995
rect 27215 2115 27245 2125
rect 27215 2095 27220 2115
rect 27240 2095 27245 2115
rect 27215 2065 27245 2095
rect 27215 2045 27220 2065
rect 27240 2045 27245 2065
rect 27215 2015 27245 2045
rect 27215 1995 27220 2015
rect 27240 1995 27245 2015
rect 27215 1985 27245 1995
rect 27270 2115 27300 2125
rect 27270 2095 27275 2115
rect 27295 2095 27300 2115
rect 27270 2065 27300 2095
rect 27270 2045 27275 2065
rect 27295 2045 27300 2065
rect 27270 2015 27300 2045
rect 27270 1995 27275 2015
rect 27295 1995 27300 2015
rect 27270 1985 27300 1995
rect 27325 2115 27355 2125
rect 27325 2095 27330 2115
rect 27350 2095 27355 2115
rect 27325 2065 27355 2095
rect 27325 2045 27330 2065
rect 27350 2045 27355 2065
rect 27325 2015 27355 2045
rect 27325 1995 27330 2015
rect 27350 1995 27355 2015
rect 27325 1985 27355 1995
rect 27380 2115 27410 2125
rect 27380 2095 27385 2115
rect 27405 2095 27410 2115
rect 27380 2065 27410 2095
rect 27380 2045 27385 2065
rect 27405 2045 27410 2065
rect 27380 2015 27410 2045
rect 27380 1995 27385 2015
rect 27405 1995 27410 2015
rect 27380 1985 27410 1995
rect 27435 2115 27465 2125
rect 27435 2095 27440 2115
rect 27460 2095 27465 2115
rect 27435 2065 27465 2095
rect 27435 2045 27440 2065
rect 27460 2045 27465 2065
rect 27435 2015 27465 2045
rect 27435 1995 27440 2015
rect 27460 1995 27465 2015
rect 27435 1985 27465 1995
rect 27490 2115 27560 2125
rect 27490 2095 27495 2115
rect 27515 2095 27535 2115
rect 27555 2095 27560 2115
rect 27490 2065 27560 2095
rect 27490 2045 27495 2065
rect 27515 2045 27535 2065
rect 27555 2045 27560 2065
rect 27490 2015 27560 2045
rect 27855 2105 27925 2135
rect 27855 2085 27860 2105
rect 27880 2085 27900 2105
rect 27920 2085 27925 2105
rect 27855 2055 27925 2085
rect 27855 2035 27860 2055
rect 27880 2035 27900 2055
rect 27920 2035 27925 2055
rect 27855 2025 27925 2035
rect 27950 2155 27980 2165
rect 27950 2135 27955 2155
rect 27975 2135 27980 2155
rect 27950 2105 27980 2135
rect 27950 2085 27955 2105
rect 27975 2085 27980 2105
rect 27950 2055 27980 2085
rect 27950 2035 27955 2055
rect 27975 2035 27980 2055
rect 27950 2025 27980 2035
rect 28005 2155 28035 2165
rect 28005 2135 28010 2155
rect 28030 2135 28035 2155
rect 28005 2105 28035 2135
rect 28005 2085 28010 2105
rect 28030 2085 28035 2105
rect 28005 2055 28035 2085
rect 28005 2035 28010 2055
rect 28030 2035 28035 2055
rect 28005 2025 28035 2035
rect 28060 2155 28090 2165
rect 28060 2135 28065 2155
rect 28085 2135 28090 2155
rect 28060 2105 28090 2135
rect 28060 2085 28065 2105
rect 28085 2085 28090 2105
rect 28060 2055 28090 2085
rect 28060 2035 28065 2055
rect 28085 2035 28090 2055
rect 28060 2025 28090 2035
rect 28115 2155 28145 2165
rect 28115 2135 28120 2155
rect 28140 2135 28145 2155
rect 28115 2105 28145 2135
rect 28115 2085 28120 2105
rect 28140 2085 28145 2105
rect 28115 2055 28145 2085
rect 28115 2035 28120 2055
rect 28140 2035 28145 2055
rect 28115 2025 28145 2035
rect 28170 2155 28200 2165
rect 28170 2135 28175 2155
rect 28195 2135 28200 2155
rect 28170 2105 28200 2135
rect 28170 2085 28175 2105
rect 28195 2085 28200 2105
rect 28170 2055 28200 2085
rect 28170 2035 28175 2055
rect 28195 2035 28200 2055
rect 28170 2025 28200 2035
rect 28225 2155 28255 2165
rect 28225 2135 28230 2155
rect 28250 2135 28255 2155
rect 28225 2105 28255 2135
rect 28225 2085 28230 2105
rect 28250 2085 28255 2105
rect 28225 2055 28255 2085
rect 28225 2035 28230 2055
rect 28250 2035 28255 2055
rect 28225 2025 28255 2035
rect 28280 2155 28310 2165
rect 28280 2135 28285 2155
rect 28305 2135 28310 2155
rect 28280 2105 28310 2135
rect 28280 2085 28285 2105
rect 28305 2085 28310 2105
rect 28280 2055 28310 2085
rect 28280 2035 28285 2055
rect 28305 2035 28310 2055
rect 28280 2025 28310 2035
rect 28335 2155 28365 2165
rect 28335 2135 28340 2155
rect 28360 2135 28365 2155
rect 28335 2105 28365 2135
rect 28335 2085 28340 2105
rect 28360 2085 28365 2105
rect 28335 2055 28365 2085
rect 28335 2035 28340 2055
rect 28360 2035 28365 2055
rect 28335 2025 28365 2035
rect 28390 2155 28420 2165
rect 28390 2135 28395 2155
rect 28415 2135 28420 2155
rect 28390 2105 28420 2135
rect 28390 2085 28395 2105
rect 28415 2085 28420 2105
rect 28390 2055 28420 2085
rect 28390 2035 28395 2055
rect 28415 2035 28420 2055
rect 28390 2025 28420 2035
rect 28445 2155 28475 2165
rect 28445 2135 28450 2155
rect 28470 2135 28475 2155
rect 28445 2105 28475 2135
rect 28445 2085 28450 2105
rect 28470 2085 28475 2105
rect 28445 2055 28475 2085
rect 28445 2035 28450 2055
rect 28470 2035 28475 2055
rect 28445 2025 28475 2035
rect 28500 2155 28530 2165
rect 28500 2135 28505 2155
rect 28525 2135 28530 2155
rect 28500 2105 28530 2135
rect 28500 2085 28505 2105
rect 28525 2085 28530 2105
rect 28500 2055 28530 2085
rect 28500 2035 28505 2055
rect 28525 2035 28530 2055
rect 28500 2025 28530 2035
rect 28555 2155 28585 2165
rect 28555 2135 28560 2155
rect 28580 2135 28585 2155
rect 28555 2105 28585 2135
rect 28555 2085 28560 2105
rect 28580 2085 28585 2105
rect 28555 2055 28585 2085
rect 28555 2035 28560 2055
rect 28580 2035 28585 2055
rect 28555 2025 28585 2035
rect 28610 2155 28640 2165
rect 28610 2135 28615 2155
rect 28635 2135 28640 2155
rect 28610 2105 28640 2135
rect 28610 2085 28615 2105
rect 28635 2085 28640 2105
rect 28610 2055 28640 2085
rect 28610 2035 28615 2055
rect 28635 2035 28640 2055
rect 28610 2025 28640 2035
rect 28665 2155 28695 2165
rect 28665 2135 28670 2155
rect 28690 2135 28695 2155
rect 28665 2105 28695 2135
rect 28665 2085 28670 2105
rect 28690 2085 28695 2105
rect 28665 2055 28695 2085
rect 28665 2035 28670 2055
rect 28690 2035 28695 2055
rect 28665 2025 28695 2035
rect 28720 2155 28750 2165
rect 28720 2135 28725 2155
rect 28745 2135 28750 2155
rect 28720 2105 28750 2135
rect 28720 2085 28725 2105
rect 28745 2085 28750 2105
rect 28720 2055 28750 2085
rect 28720 2035 28725 2055
rect 28745 2035 28750 2055
rect 28720 2025 28750 2035
rect 28775 2155 28805 2165
rect 28775 2135 28780 2155
rect 28800 2135 28805 2155
rect 28775 2105 28805 2135
rect 28775 2085 28780 2105
rect 28800 2085 28805 2105
rect 28775 2055 28805 2085
rect 28775 2035 28780 2055
rect 28800 2035 28805 2055
rect 28775 2025 28805 2035
rect 28830 2155 28860 2165
rect 28830 2135 28835 2155
rect 28855 2135 28860 2155
rect 28830 2105 28860 2135
rect 28830 2085 28835 2105
rect 28855 2085 28860 2105
rect 28830 2055 28860 2085
rect 28830 2035 28835 2055
rect 28855 2035 28860 2055
rect 28830 2025 28860 2035
rect 28885 2155 28915 2165
rect 28885 2135 28890 2155
rect 28910 2135 28915 2155
rect 28885 2105 28915 2135
rect 28885 2085 28890 2105
rect 28910 2085 28915 2105
rect 28885 2055 28915 2085
rect 28885 2035 28890 2055
rect 28910 2035 28915 2055
rect 28885 2025 28915 2035
rect 28940 2155 28970 2165
rect 28940 2135 28945 2155
rect 28965 2135 28970 2155
rect 28940 2105 28970 2135
rect 28940 2085 28945 2105
rect 28965 2085 28970 2105
rect 28940 2055 28970 2085
rect 28940 2035 28945 2055
rect 28965 2035 28970 2055
rect 28940 2025 28970 2035
rect 28995 2155 29025 2165
rect 28995 2135 29000 2155
rect 29020 2135 29025 2155
rect 28995 2105 29025 2135
rect 28995 2085 29000 2105
rect 29020 2085 29025 2105
rect 28995 2055 29025 2085
rect 28995 2035 29000 2055
rect 29020 2035 29025 2055
rect 28995 2025 29025 2035
rect 29050 2155 29080 2165
rect 29050 2135 29055 2155
rect 29075 2135 29080 2155
rect 29050 2105 29080 2135
rect 29050 2085 29055 2105
rect 29075 2085 29080 2105
rect 29050 2055 29080 2085
rect 29050 2035 29055 2055
rect 29075 2035 29080 2055
rect 29050 2025 29080 2035
rect 29105 2155 29175 2165
rect 29105 2135 29110 2155
rect 29130 2135 29150 2155
rect 29170 2135 29175 2155
rect 29105 2105 29175 2135
rect 29105 2085 29110 2105
rect 29130 2085 29150 2105
rect 29170 2085 29175 2105
rect 29105 2055 29175 2085
rect 29105 2035 29110 2055
rect 29130 2035 29150 2055
rect 29170 2035 29175 2055
rect 29105 2025 29175 2035
rect 27490 1995 27495 2015
rect 27515 1995 27535 2015
rect 27555 1995 27560 2015
rect 27955 2005 27975 2025
rect 28065 2005 28085 2025
rect 28175 2005 28195 2025
rect 28285 2005 28305 2025
rect 28395 2005 28415 2025
rect 28505 2005 28525 2025
rect 28615 2005 28635 2025
rect 28725 2005 28745 2025
rect 28835 2005 28855 2025
rect 28945 2005 28965 2025
rect 29055 2005 29075 2025
rect 27490 1985 27560 1995
rect 27945 1995 27985 2005
rect 25835 1965 25875 1975
rect 26245 1965 26265 1985
rect 26395 1965 26415 1985
rect 26505 1965 26525 1985
rect 26615 1965 26635 1985
rect 26725 1965 26745 1985
rect 26835 1965 26855 1985
rect 26945 1965 26965 1985
rect 27055 1965 27075 1985
rect 27165 1965 27185 1985
rect 27275 1965 27295 1985
rect 27385 1965 27405 1985
rect 27535 1965 27555 1985
rect 27945 1975 27957 1995
rect 27975 1975 27985 1995
rect 27945 1965 27985 1975
rect 28055 1995 28095 2005
rect 28055 1975 28067 1995
rect 28085 1975 28095 1995
rect 28055 1965 28095 1975
rect 28165 1995 28205 2005
rect 28165 1975 28177 1995
rect 28195 1975 28205 1995
rect 28165 1965 28205 1975
rect 28275 1995 28315 2005
rect 28275 1975 28287 1995
rect 28305 1975 28315 1995
rect 28275 1965 28315 1975
rect 28385 1995 28425 2005
rect 28385 1975 28397 1995
rect 28415 1975 28425 1995
rect 28385 1965 28425 1975
rect 28495 1995 28535 2005
rect 28495 1975 28507 1995
rect 28525 1975 28535 1995
rect 28495 1965 28535 1975
rect 28605 1995 28645 2005
rect 28605 1975 28617 1995
rect 28635 1975 28645 1995
rect 28605 1965 28645 1975
rect 28715 1995 28755 2005
rect 28715 1975 28727 1995
rect 28745 1975 28755 1995
rect 28715 1965 28755 1975
rect 28825 1995 28865 2005
rect 28825 1975 28837 1995
rect 28855 1975 28865 1995
rect 28825 1965 28865 1975
rect 28935 1995 28975 2005
rect 28935 1975 28947 1995
rect 28965 1975 28975 1995
rect 28935 1965 28975 1975
rect 29045 1995 29085 2005
rect 29045 1975 29057 1995
rect 29075 1975 29085 1995
rect 29045 1965 29085 1975
rect 26235 1955 26275 1965
rect 12525 1925 12565 1935
rect 13000 1940 13040 1950
rect 10760 1910 10800 1920
rect 13000 1920 13012 1940
rect 13030 1920 13040 1940
rect 13000 1910 13040 1920
rect 13110 1940 13150 1950
rect 13110 1920 13122 1940
rect 13140 1920 13150 1940
rect 13110 1910 13150 1920
rect 13220 1940 13260 1950
rect 13220 1920 13232 1940
rect 13250 1920 13260 1940
rect 13220 1910 13260 1920
rect 13330 1940 13370 1950
rect 13330 1920 13342 1940
rect 13360 1920 13370 1940
rect 13330 1910 13370 1920
rect 13440 1940 13480 1950
rect 13440 1920 13452 1940
rect 13470 1920 13480 1940
rect 13440 1910 13480 1920
rect 13550 1940 13590 1950
rect 13550 1920 13562 1940
rect 13580 1920 13590 1940
rect 26235 1935 26245 1955
rect 26265 1935 26275 1955
rect 26235 1925 26275 1935
rect 26385 1955 26425 1965
rect 26385 1935 26395 1955
rect 26415 1935 26425 1955
rect 26385 1925 26425 1935
rect 26495 1955 26535 1965
rect 26495 1935 26505 1955
rect 26525 1935 26535 1955
rect 26495 1925 26535 1935
rect 26605 1955 26645 1965
rect 26605 1935 26615 1955
rect 26635 1935 26645 1955
rect 26605 1925 26645 1935
rect 26715 1955 26755 1965
rect 26715 1935 26725 1955
rect 26745 1935 26755 1955
rect 26715 1925 26755 1935
rect 26825 1955 26865 1965
rect 26825 1935 26835 1955
rect 26855 1935 26865 1955
rect 26825 1925 26865 1935
rect 26935 1955 26975 1965
rect 26935 1935 26945 1955
rect 26965 1935 26975 1955
rect 26935 1925 26975 1935
rect 27045 1955 27085 1965
rect 27045 1935 27055 1955
rect 27075 1935 27085 1955
rect 27045 1925 27085 1935
rect 27155 1955 27195 1965
rect 27155 1935 27165 1955
rect 27185 1935 27195 1955
rect 27155 1925 27195 1935
rect 27265 1955 27305 1965
rect 27265 1935 27275 1955
rect 27295 1935 27305 1955
rect 27265 1925 27305 1935
rect 27375 1955 27415 1965
rect 27375 1935 27385 1955
rect 27405 1935 27415 1955
rect 27375 1925 27415 1935
rect 27525 1955 27565 1965
rect 27525 1935 27535 1955
rect 27555 1935 27565 1955
rect 27525 1925 27565 1935
rect 13550 1910 13590 1920
rect 2575 1885 2595 1905
rect 2685 1885 2705 1905
rect 2755 1885 2775 1905
rect 2935 1885 2955 1905
rect 3055 1885 3075 1905
rect 3295 1885 3315 1905
rect 3415 1885 3435 1905
rect 3655 1885 3675 1905
rect 3775 1885 3795 1905
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2755 1875 2805 1885
rect 2755 1855 2775 1875
rect 2795 1855 2805 1875
rect 2755 1845 2805 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1875 2965 1885
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1875 3325 1885
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1875 3685 1885
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3995 1880 4015 1905
rect 4215 1885 4235 1905
rect 4335 1885 4355 1905
rect 4575 1885 4595 1905
rect 4695 1885 4715 1905
rect 4935 1885 4955 1905
rect 5055 1885 5075 1905
rect 5235 1885 5255 1905
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1880
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1875 4365 1885
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1875 4725 1885
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1875 5085 1885
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5255 1885
rect 5205 1855 5215 1875
rect 5235 1855 5255 1875
rect 27950 1900 27990 1910
rect 27950 1880 27960 1900
rect 27980 1880 27990 1900
rect 27950 1870 27990 1880
rect 28045 1900 28085 1910
rect 28045 1880 28055 1900
rect 28075 1880 28085 1900
rect 28045 1870 28085 1880
rect 28155 1900 28195 1910
rect 28155 1880 28165 1900
rect 28185 1880 28195 1900
rect 28155 1870 28195 1880
rect 28265 1900 28305 1910
rect 28265 1880 28275 1900
rect 28295 1880 28305 1900
rect 28265 1870 28305 1880
rect 28360 1900 28400 1910
rect 28360 1880 28370 1900
rect 28390 1880 28400 1900
rect 28360 1870 28400 1880
rect 5205 1845 5255 1855
rect 27960 1850 27980 1870
rect 28055 1850 28075 1870
rect 28165 1850 28185 1870
rect 28275 1850 28295 1870
rect 28370 1850 28390 1870
rect 27955 1840 28025 1850
rect 2475 1790 2505 1820
rect 2835 1785 2875 1825
rect 3045 1815 3085 1825
rect 3045 1795 3055 1815
rect 3075 1795 3085 1815
rect 3045 1785 3085 1795
rect 3165 1785 3205 1825
rect 3405 1815 3445 1825
rect 3405 1795 3415 1815
rect 3435 1795 3445 1815
rect 3405 1785 3445 1795
rect 3525 1785 3565 1825
rect 3765 1815 3805 1825
rect 3765 1795 3775 1815
rect 3795 1795 3805 1815
rect 3765 1785 3805 1795
rect 3855 1785 3895 1825
rect 4115 1785 4155 1825
rect 4205 1815 4245 1825
rect 4205 1795 4215 1815
rect 4235 1795 4245 1815
rect 4205 1785 4245 1795
rect 4445 1785 4485 1825
rect 4565 1815 4605 1825
rect 4565 1795 4575 1815
rect 4595 1795 4605 1815
rect 4565 1785 4605 1795
rect 4805 1785 4845 1825
rect 4925 1815 4965 1825
rect 4925 1795 4935 1815
rect 4955 1795 4965 1815
rect 4925 1785 4965 1795
rect 5135 1785 5175 1825
rect 27955 1820 27960 1840
rect 27980 1820 28000 1840
rect 28020 1820 28025 1840
rect 5365 1790 5395 1820
rect 27955 1790 28025 1820
rect 11190 1770 11230 1780
rect 2430 1730 2460 1760
rect 2570 1730 2600 1760
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1725 3265 1735
rect 3285 1755 3325 1765
rect 3285 1735 3295 1755
rect 3315 1735 3325 1755
rect 3285 1725 3325 1735
rect 3525 1755 3565 1765
rect 3525 1735 3535 1755
rect 3555 1735 3565 1755
rect 3525 1725 3565 1735
rect 3765 1755 3805 1765
rect 3765 1735 3775 1755
rect 3795 1735 3805 1755
rect 3765 1725 3805 1735
rect 4205 1755 4245 1765
rect 4205 1735 4215 1755
rect 4235 1735 4245 1755
rect 4205 1725 4245 1735
rect 4445 1755 4485 1765
rect 4445 1735 4455 1755
rect 4475 1735 4485 1755
rect 4445 1725 4485 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1725 4725 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1725 4785 1735
rect 5275 1730 5305 1760
rect 11085 1755 11125 1765
rect 11085 1735 11095 1755
rect 11115 1735 11125 1755
rect 11190 1750 11200 1770
rect 11220 1750 11230 1770
rect 11410 1770 11450 1780
rect 11190 1740 11230 1750
rect 11305 1755 11345 1765
rect 11085 1725 11125 1735
rect 3165 1710 3205 1720
rect 2805 1680 2835 1710
rect 3165 1690 3175 1710
rect 3195 1690 3205 1710
rect 3165 1680 3205 1690
rect 2385 1635 2415 1665
rect 2625 1635 2655 1665
rect 3175 1660 3195 1680
rect 3295 1660 3315 1725
rect 3405 1710 3445 1720
rect 3405 1690 3415 1710
rect 3435 1690 3445 1710
rect 3405 1680 3445 1690
rect 3415 1660 3435 1680
rect 3535 1660 3555 1725
rect 3645 1710 3685 1720
rect 3645 1690 3655 1710
rect 3675 1690 3685 1710
rect 3645 1680 3685 1690
rect 3655 1660 3675 1680
rect 3775 1660 3795 1725
rect 4215 1660 4235 1725
rect 4325 1710 4365 1720
rect 4325 1690 4335 1710
rect 4355 1690 4365 1710
rect 4325 1680 4365 1690
rect 4335 1660 4355 1680
rect 4455 1660 4475 1725
rect 4565 1710 4605 1720
rect 4565 1690 4575 1710
rect 4595 1690 4605 1710
rect 4565 1680 4605 1690
rect 4575 1660 4595 1680
rect 4695 1660 4715 1725
rect 4805 1710 4845 1720
rect 4805 1690 4815 1710
rect 4835 1690 4845 1710
rect 4805 1680 4845 1690
rect 10255 1700 10295 1710
rect 10255 1680 10265 1700
rect 10285 1680 10295 1700
rect 4815 1660 4835 1680
rect 10255 1670 10295 1680
rect 10455 1700 10495 1710
rect 10455 1680 10465 1700
rect 10485 1680 10495 1700
rect 10455 1670 10495 1680
rect 10558 1700 10592 1710
rect 10558 1680 10566 1700
rect 10584 1680 10592 1700
rect 10558 1670 10592 1680
rect 10655 1700 10695 1710
rect 10655 1680 10665 1700
rect 10685 1680 10695 1700
rect 10655 1670 10695 1680
rect 3170 1650 3200 1660
rect 3170 1630 3175 1650
rect 3195 1630 3200 1650
rect 3170 1620 3200 1630
rect 3230 1650 3260 1660
rect 3230 1630 3235 1650
rect 3255 1630 3260 1650
rect 3230 1620 3260 1630
rect 3290 1650 3320 1660
rect 3290 1630 3295 1650
rect 3315 1630 3320 1650
rect 3290 1620 3320 1630
rect 3350 1650 3380 1660
rect 3350 1630 3355 1650
rect 3375 1630 3380 1650
rect 3350 1620 3380 1630
rect 3410 1650 3440 1660
rect 3410 1630 3415 1650
rect 3435 1630 3440 1650
rect 3410 1620 3440 1630
rect 3470 1650 3500 1660
rect 3470 1630 3475 1650
rect 3495 1630 3500 1650
rect 3470 1620 3500 1630
rect 3530 1650 3560 1660
rect 3530 1630 3535 1650
rect 3555 1630 3560 1650
rect 3530 1620 3560 1630
rect 3590 1650 3620 1660
rect 3590 1630 3595 1650
rect 3615 1630 3620 1650
rect 3590 1620 3620 1630
rect 3650 1650 3680 1660
rect 3650 1630 3655 1650
rect 3675 1630 3680 1650
rect 3650 1620 3680 1630
rect 3710 1650 3740 1660
rect 3710 1630 3715 1650
rect 3735 1630 3740 1650
rect 3710 1620 3740 1630
rect 3770 1650 3800 1660
rect 3770 1630 3775 1650
rect 3795 1630 3800 1650
rect 3770 1620 3800 1630
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 4210 1650 4240 1660
rect 4210 1630 4215 1650
rect 4235 1630 4240 1650
rect 4210 1620 4240 1630
rect 4270 1650 4300 1660
rect 4270 1630 4275 1650
rect 4295 1630 4300 1650
rect 4270 1620 4300 1630
rect 4330 1650 4360 1660
rect 4330 1630 4335 1650
rect 4355 1630 4360 1650
rect 4330 1620 4360 1630
rect 4390 1650 4420 1660
rect 4390 1630 4395 1650
rect 4415 1630 4420 1650
rect 4390 1620 4420 1630
rect 4450 1650 4480 1660
rect 4450 1630 4455 1650
rect 4475 1630 4480 1650
rect 4450 1620 4480 1630
rect 4510 1650 4540 1660
rect 4510 1630 4515 1650
rect 4535 1630 4540 1650
rect 4510 1620 4540 1630
rect 4570 1650 4600 1660
rect 4570 1630 4575 1650
rect 4595 1630 4600 1650
rect 4570 1620 4600 1630
rect 4630 1650 4660 1660
rect 4630 1630 4635 1650
rect 4655 1630 4660 1650
rect 4630 1620 4660 1630
rect 4690 1650 4720 1660
rect 4690 1630 4695 1650
rect 4715 1630 4720 1650
rect 4690 1620 4720 1630
rect 4750 1650 4780 1660
rect 4750 1630 4755 1650
rect 4775 1630 4780 1650
rect 4750 1620 4780 1630
rect 4810 1650 4840 1660
rect 10265 1650 10285 1670
rect 10465 1650 10485 1670
rect 10665 1650 10685 1670
rect 11095 1660 11115 1725
rect 11200 1660 11220 1740
rect 11305 1735 11315 1755
rect 11335 1735 11345 1755
rect 11410 1750 11420 1770
rect 11440 1750 11450 1770
rect 11640 1770 11680 1780
rect 11410 1740 11450 1750
rect 11525 1755 11565 1765
rect 11305 1725 11345 1735
rect 11237 1710 11269 1720
rect 11237 1690 11243 1710
rect 11260 1690 11269 1710
rect 11237 1680 11269 1690
rect 11315 1660 11335 1725
rect 11420 1660 11440 1740
rect 11525 1735 11535 1755
rect 11555 1735 11565 1755
rect 11640 1750 11650 1770
rect 11670 1750 11680 1770
rect 12230 1770 12270 1780
rect 11640 1740 11680 1750
rect 12125 1755 12165 1765
rect 11525 1725 11565 1735
rect 11457 1710 11489 1720
rect 11457 1690 11463 1710
rect 11480 1690 11489 1710
rect 11457 1680 11489 1690
rect 11535 1660 11555 1725
rect 11601 1710 11633 1720
rect 11601 1690 11610 1710
rect 11627 1690 11633 1710
rect 11601 1680 11633 1690
rect 11650 1660 11670 1740
rect 12125 1735 12135 1755
rect 12155 1735 12165 1755
rect 12230 1750 12240 1770
rect 12260 1750 12270 1770
rect 12450 1770 12490 1780
rect 12230 1740 12270 1750
rect 12345 1755 12385 1765
rect 12125 1725 12165 1735
rect 11820 1710 11850 1720
rect 11820 1690 11825 1710
rect 11845 1690 11850 1710
rect 11820 1680 11850 1690
rect 11867 1710 11899 1720
rect 11867 1690 11876 1710
rect 11893 1690 11899 1710
rect 11867 1680 11899 1690
rect 11950 1710 11980 1720
rect 11950 1690 11955 1710
rect 11975 1690 11980 1710
rect 11950 1680 11980 1690
rect 11830 1660 11850 1680
rect 11950 1660 11970 1680
rect 12135 1660 12155 1725
rect 12240 1660 12260 1740
rect 12345 1735 12355 1755
rect 12375 1735 12385 1755
rect 12450 1750 12460 1770
rect 12480 1750 12490 1770
rect 12680 1770 12720 1780
rect 12450 1740 12490 1750
rect 12565 1755 12605 1765
rect 12345 1725 12385 1735
rect 12277 1710 12309 1720
rect 12277 1690 12283 1710
rect 12300 1690 12309 1710
rect 12277 1680 12309 1690
rect 12355 1660 12375 1725
rect 12460 1660 12480 1740
rect 12565 1735 12575 1755
rect 12595 1735 12605 1755
rect 12680 1750 12690 1770
rect 12710 1750 12720 1770
rect 26190 1770 26230 1780
rect 12680 1740 12720 1750
rect 26085 1755 26125 1765
rect 12565 1725 12605 1735
rect 12497 1710 12529 1720
rect 12497 1690 12503 1710
rect 12520 1690 12529 1710
rect 12497 1680 12529 1690
rect 12575 1660 12595 1725
rect 12641 1710 12673 1720
rect 12641 1690 12650 1710
rect 12667 1690 12673 1710
rect 12641 1680 12673 1690
rect 12690 1660 12710 1740
rect 26085 1735 26095 1755
rect 26115 1735 26125 1755
rect 26190 1750 26200 1770
rect 26220 1750 26230 1770
rect 26410 1770 26450 1780
rect 26190 1740 26230 1750
rect 26305 1755 26345 1765
rect 26085 1725 26125 1735
rect 13105 1700 13145 1710
rect 13105 1680 13115 1700
rect 13135 1680 13145 1700
rect 13105 1670 13145 1680
rect 13208 1700 13242 1710
rect 13208 1680 13216 1700
rect 13234 1680 13242 1700
rect 13208 1670 13242 1680
rect 13305 1700 13345 1710
rect 13305 1680 13315 1700
rect 13335 1680 13345 1700
rect 13305 1670 13345 1680
rect 13505 1700 13545 1710
rect 13505 1680 13515 1700
rect 13535 1680 13545 1700
rect 13505 1670 13545 1680
rect 10990 1650 11065 1660
rect 4810 1630 4815 1650
rect 4835 1630 4840 1650
rect 4810 1620 4840 1630
rect 9970 1640 10005 1650
rect 2335 1565 2365 1595
rect 3165 1590 3205 1600
rect 3165 1570 3175 1590
rect 3195 1570 3205 1590
rect 3165 1560 3205 1570
rect 3235 1550 3255 1620
rect 3355 1550 3375 1620
rect 3475 1550 3495 1620
rect 3595 1550 3615 1620
rect 3715 1550 3735 1620
rect 4275 1550 4295 1620
rect 4395 1550 4415 1620
rect 4515 1550 4535 1620
rect 4635 1550 4655 1620
rect 4755 1550 4775 1620
rect 9970 1615 9975 1640
rect 10000 1615 10005 1640
rect 9970 1605 10005 1615
rect 4805 1590 4845 1600
rect 4805 1570 4815 1590
rect 4835 1570 4845 1590
rect 4805 1560 4845 1570
rect 5415 1565 5445 1595
rect 3225 1540 3265 1550
rect 3225 1520 3235 1540
rect 3255 1520 3265 1540
rect 3225 1510 3265 1520
rect 3345 1540 3385 1550
rect 3345 1520 3355 1540
rect 3375 1520 3385 1540
rect 3345 1510 3385 1520
rect 3465 1540 3505 1550
rect 3465 1520 3475 1540
rect 3495 1520 3505 1540
rect 3465 1510 3505 1520
rect 3585 1540 3625 1550
rect 3585 1520 3595 1540
rect 3615 1520 3625 1540
rect 3585 1510 3625 1520
rect 3705 1540 3745 1550
rect 3705 1520 3715 1540
rect 3735 1520 3745 1540
rect 3705 1510 3745 1520
rect 4265 1540 4305 1550
rect 4265 1520 4275 1540
rect 4295 1520 4305 1540
rect 4265 1510 4305 1520
rect 4385 1540 4425 1550
rect 4385 1520 4395 1540
rect 4415 1520 4425 1540
rect 4385 1510 4425 1520
rect 4505 1540 4545 1550
rect 4505 1520 4515 1540
rect 4535 1520 4545 1540
rect 4505 1510 4545 1520
rect 4625 1540 4665 1550
rect 4625 1520 4635 1540
rect 4655 1520 4665 1540
rect 4625 1510 4665 1520
rect 4745 1540 4785 1550
rect 4745 1520 4755 1540
rect 4775 1520 4785 1540
rect 4745 1510 4785 1520
rect 2925 1495 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1465 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1465 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1465 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1465 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1465 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1465 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 4205 1495 4245 1505
rect 3765 1465 3805 1475
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1465 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1465 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1465 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1465 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1465 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1465 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1465 5085 1475
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1440 2870 1450
rect 2840 1420 2845 1440
rect 2865 1420 2870 1440
rect 2840 1390 2870 1420
rect 2840 1370 2845 1390
rect 2865 1370 2870 1390
rect 2840 1340 2870 1370
rect 2840 1320 2845 1340
rect 2865 1320 2870 1340
rect 2840 1290 2870 1320
rect 2840 1270 2845 1290
rect 2865 1270 2870 1290
rect 2840 1240 2870 1270
rect 2840 1220 2845 1240
rect 2865 1220 2870 1240
rect 2840 1210 2870 1220
rect 3380 1440 3410 1450
rect 3380 1420 3385 1440
rect 3405 1420 3410 1440
rect 3380 1390 3410 1420
rect 3380 1370 3385 1390
rect 3405 1370 3410 1390
rect 3380 1340 3410 1370
rect 3380 1320 3385 1340
rect 3405 1320 3410 1340
rect 3380 1290 3410 1320
rect 3380 1270 3385 1290
rect 3405 1270 3410 1290
rect 3380 1240 3410 1270
rect 3380 1220 3385 1240
rect 3405 1220 3410 1240
rect 3380 1210 3410 1220
rect 3920 1440 3950 1450
rect 3920 1420 3925 1440
rect 3945 1420 3950 1440
rect 3920 1390 3950 1420
rect 3920 1370 3925 1390
rect 3945 1370 3950 1390
rect 3920 1340 3950 1370
rect 3920 1320 3925 1340
rect 3945 1320 3950 1340
rect 3920 1290 3950 1320
rect 3920 1270 3925 1290
rect 3945 1270 3950 1290
rect 3920 1240 3950 1270
rect 3920 1220 3925 1240
rect 3945 1220 3950 1240
rect 3920 1210 3950 1220
rect 4060 1440 4090 1450
rect 4060 1420 4065 1440
rect 4085 1420 4090 1440
rect 4060 1390 4090 1420
rect 4060 1370 4065 1390
rect 4085 1370 4090 1390
rect 4060 1340 4090 1370
rect 4060 1320 4065 1340
rect 4085 1320 4090 1340
rect 4060 1290 4090 1320
rect 4060 1270 4065 1290
rect 4085 1270 4090 1290
rect 4060 1240 4090 1270
rect 4060 1220 4065 1240
rect 4085 1220 4090 1240
rect 4060 1210 4090 1220
rect 4600 1440 4630 1450
rect 4600 1420 4605 1440
rect 4625 1420 4630 1440
rect 4600 1390 4630 1420
rect 4600 1370 4605 1390
rect 4625 1370 4630 1390
rect 4600 1340 4630 1370
rect 4600 1320 4605 1340
rect 4625 1320 4630 1340
rect 4600 1290 4630 1320
rect 4600 1270 4605 1290
rect 4625 1270 4630 1290
rect 4600 1240 4630 1270
rect 4600 1220 4605 1240
rect 4625 1220 4630 1240
rect 4600 1210 4630 1220
rect 5140 1440 5170 1450
rect 5140 1420 5145 1440
rect 5165 1420 5170 1440
rect 5140 1390 5170 1420
rect 5140 1370 5145 1390
rect 5165 1370 5170 1390
rect 10030 1640 10065 1650
rect 10030 1615 10035 1640
rect 10060 1615 10065 1640
rect 10030 1605 10065 1615
rect 10120 1640 10190 1650
rect 10120 1620 10125 1640
rect 10145 1620 10165 1640
rect 10185 1620 10190 1640
rect 10120 1590 10190 1620
rect 10120 1570 10125 1590
rect 10145 1570 10165 1590
rect 10185 1570 10190 1590
rect 10120 1540 10190 1570
rect 10120 1520 10125 1540
rect 10145 1520 10165 1540
rect 10185 1520 10190 1540
rect 10120 1490 10190 1520
rect 10120 1470 10125 1490
rect 10145 1470 10165 1490
rect 10185 1470 10190 1490
rect 10120 1440 10190 1470
rect 10120 1420 10125 1440
rect 10145 1420 10165 1440
rect 10185 1420 10190 1440
rect 10120 1390 10190 1420
rect 5140 1340 5170 1370
rect 5140 1320 5145 1340
rect 5165 1320 5170 1340
rect 5140 1290 5170 1320
rect 5140 1270 5145 1290
rect 5165 1270 5170 1290
rect 5140 1240 5170 1270
rect 5140 1220 5145 1240
rect 5165 1220 5170 1240
rect 5140 1210 5170 1220
rect 10120 1370 10125 1390
rect 10145 1370 10165 1390
rect 10185 1370 10190 1390
rect 10120 1340 10190 1370
rect 10120 1320 10125 1340
rect 10145 1320 10165 1340
rect 10185 1320 10190 1340
rect 10120 1290 10190 1320
rect 10120 1270 10125 1290
rect 10145 1270 10165 1290
rect 10185 1270 10190 1290
rect 10120 1240 10190 1270
rect 10120 1220 10125 1240
rect 10145 1220 10165 1240
rect 10185 1220 10190 1240
rect 3385 1190 3405 1210
rect 4605 1190 4625 1210
rect 10120 1190 10190 1220
rect 3375 1180 3415 1190
rect 3375 1160 3385 1180
rect 3405 1160 3415 1180
rect 3375 1150 3415 1160
rect 3990 1155 4020 1185
rect 4595 1180 4635 1190
rect 4595 1160 4605 1180
rect 4625 1160 4635 1180
rect 4595 1150 4635 1160
rect 10120 1170 10125 1190
rect 10145 1170 10165 1190
rect 10185 1170 10190 1190
rect 10120 1140 10190 1170
rect 2945 1120 2985 1130
rect 2945 1100 2955 1120
rect 2975 1100 2985 1120
rect 2945 1090 2985 1100
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 3985 1120 4025 1130
rect 3985 1100 3995 1120
rect 4015 1100 4025 1120
rect 3985 1090 4025 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2955 1070 2975 1090
rect 3995 1070 4015 1090
rect 2950 1060 2980 1070
rect 2950 1045 2955 1060
rect 2935 1040 2955 1045
rect 2975 1040 2980 1060
rect 2625 1010 2655 1040
rect 2910 1035 2980 1040
rect 2910 1015 2915 1035
rect 2935 1015 2980 1035
rect 2910 1010 2980 1015
rect 2935 1005 2955 1010
rect 2950 990 2955 1005
rect 2975 990 2980 1010
rect 2950 980 2980 990
rect 3990 1060 4020 1070
rect 3990 1040 3995 1060
rect 4015 1040 4020 1060
rect 3990 1010 4020 1040
rect 3990 990 3995 1010
rect 4015 990 4020 1010
rect 3990 980 4020 990
rect 5030 1060 5100 1070
rect 5030 1040 5035 1060
rect 5055 1040 5075 1060
rect 5095 1045 5100 1060
rect 5095 1040 5150 1045
rect 5030 1035 5150 1040
rect 5030 1015 5120 1035
rect 5140 1015 5150 1035
rect 5030 1010 5150 1015
rect 5030 990 5035 1010
rect 5055 990 5075 1010
rect 5095 1005 5150 1010
rect 5095 990 5100 1005
rect 5030 980 5100 990
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 2995 895 3035 905
rect 3175 925 3215 935
rect 3175 905 3185 925
rect 3205 905 3215 925
rect 3175 895 3215 905
rect 3355 925 3395 935
rect 3355 905 3365 925
rect 3385 905 3395 925
rect 3355 895 3395 905
rect 3535 925 3575 935
rect 3535 905 3545 925
rect 3565 905 3575 925
rect 3535 895 3575 905
rect 3715 925 3755 935
rect 3715 905 3725 925
rect 3745 905 3755 925
rect 3715 895 3755 905
rect 3895 925 3935 935
rect 3895 905 3905 925
rect 3925 905 3935 925
rect 3895 895 3935 905
rect 4075 925 4115 935
rect 4075 905 4085 925
rect 4105 905 4115 925
rect 4075 895 4115 905
rect 4255 925 4295 935
rect 4255 905 4265 925
rect 4285 905 4295 925
rect 4255 895 4295 905
rect 4435 925 4475 935
rect 4435 905 4445 925
rect 4465 905 4475 925
rect 4435 895 4475 905
rect 4615 925 4655 935
rect 4615 905 4625 925
rect 4645 905 4655 925
rect 4615 895 4655 905
rect 4795 925 4835 935
rect 4795 905 4805 925
rect 4825 905 4835 925
rect 4795 895 4835 905
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 10005 910 10030 960
rect 10120 1120 10125 1140
rect 10145 1120 10165 1140
rect 10185 1120 10190 1140
rect 10120 1090 10190 1120
rect 10120 1070 10125 1090
rect 10145 1070 10165 1090
rect 10185 1070 10190 1090
rect 10120 1040 10190 1070
rect 10120 1020 10125 1040
rect 10145 1020 10165 1040
rect 10185 1020 10190 1040
rect 10120 990 10190 1020
rect 10120 970 10125 990
rect 10145 970 10165 990
rect 10185 970 10190 990
rect 10120 960 10190 970
rect 10260 1640 10290 1650
rect 10260 1620 10265 1640
rect 10285 1620 10290 1640
rect 10260 1590 10290 1620
rect 10260 1570 10265 1590
rect 10285 1570 10290 1590
rect 10260 1540 10290 1570
rect 10260 1520 10265 1540
rect 10285 1520 10290 1540
rect 10260 1490 10290 1520
rect 10260 1470 10265 1490
rect 10285 1470 10290 1490
rect 10260 1440 10290 1470
rect 10260 1420 10265 1440
rect 10285 1420 10290 1440
rect 10260 1390 10290 1420
rect 10260 1370 10265 1390
rect 10285 1370 10290 1390
rect 10260 1340 10290 1370
rect 10260 1320 10265 1340
rect 10285 1320 10290 1340
rect 10260 1290 10290 1320
rect 10260 1270 10265 1290
rect 10285 1270 10290 1290
rect 10260 1240 10290 1270
rect 10260 1220 10265 1240
rect 10285 1220 10290 1240
rect 10260 1190 10290 1220
rect 10260 1170 10265 1190
rect 10285 1170 10290 1190
rect 10260 1140 10290 1170
rect 10260 1120 10265 1140
rect 10285 1120 10290 1140
rect 10260 1090 10290 1120
rect 10260 1070 10265 1090
rect 10285 1070 10290 1090
rect 10260 1040 10290 1070
rect 10260 1020 10265 1040
rect 10285 1020 10290 1040
rect 10260 990 10290 1020
rect 10260 970 10265 990
rect 10285 970 10290 990
rect 10260 960 10290 970
rect 10360 1640 10390 1650
rect 10360 1620 10365 1640
rect 10385 1620 10390 1640
rect 10360 1590 10390 1620
rect 10360 1570 10365 1590
rect 10385 1570 10390 1590
rect 10360 1540 10390 1570
rect 10360 1520 10365 1540
rect 10385 1520 10390 1540
rect 10360 1490 10390 1520
rect 10360 1470 10365 1490
rect 10385 1470 10390 1490
rect 10360 1440 10390 1470
rect 10360 1420 10365 1440
rect 10385 1420 10390 1440
rect 10360 1390 10390 1420
rect 10360 1370 10365 1390
rect 10385 1370 10390 1390
rect 10360 1340 10390 1370
rect 10360 1320 10365 1340
rect 10385 1320 10390 1340
rect 10360 1290 10390 1320
rect 10360 1270 10365 1290
rect 10385 1270 10390 1290
rect 10360 1240 10390 1270
rect 10360 1220 10365 1240
rect 10385 1220 10390 1240
rect 10360 1190 10390 1220
rect 10360 1170 10365 1190
rect 10385 1170 10390 1190
rect 10360 1140 10390 1170
rect 10360 1120 10365 1140
rect 10385 1120 10390 1140
rect 10360 1090 10390 1120
rect 10360 1070 10365 1090
rect 10385 1070 10390 1090
rect 10360 1040 10390 1070
rect 10360 1020 10365 1040
rect 10385 1020 10390 1040
rect 10360 990 10390 1020
rect 10360 970 10365 990
rect 10385 970 10390 990
rect 10360 960 10390 970
rect 10460 1640 10490 1650
rect 10460 1620 10465 1640
rect 10485 1620 10490 1640
rect 10460 1590 10490 1620
rect 10460 1570 10465 1590
rect 10485 1570 10490 1590
rect 10460 1540 10490 1570
rect 10460 1520 10465 1540
rect 10485 1520 10490 1540
rect 10460 1490 10490 1520
rect 10460 1470 10465 1490
rect 10485 1470 10490 1490
rect 10460 1440 10490 1470
rect 10460 1420 10465 1440
rect 10485 1420 10490 1440
rect 10460 1390 10490 1420
rect 10460 1370 10465 1390
rect 10485 1370 10490 1390
rect 10460 1340 10490 1370
rect 10460 1320 10465 1340
rect 10485 1320 10490 1340
rect 10460 1290 10490 1320
rect 10460 1270 10465 1290
rect 10485 1270 10490 1290
rect 10460 1240 10490 1270
rect 10460 1220 10465 1240
rect 10485 1220 10490 1240
rect 10460 1190 10490 1220
rect 10460 1170 10465 1190
rect 10485 1170 10490 1190
rect 10460 1140 10490 1170
rect 10460 1120 10465 1140
rect 10485 1120 10490 1140
rect 10460 1090 10490 1120
rect 10460 1070 10465 1090
rect 10485 1070 10490 1090
rect 10460 1040 10490 1070
rect 10460 1020 10465 1040
rect 10485 1020 10490 1040
rect 10460 990 10490 1020
rect 10460 970 10465 990
rect 10485 970 10490 990
rect 10460 960 10490 970
rect 10560 1640 10590 1650
rect 10560 1620 10565 1640
rect 10585 1620 10590 1640
rect 10560 1590 10590 1620
rect 10560 1570 10565 1590
rect 10585 1570 10590 1590
rect 10560 1540 10590 1570
rect 10560 1520 10565 1540
rect 10585 1520 10590 1540
rect 10560 1490 10590 1520
rect 10560 1470 10565 1490
rect 10585 1470 10590 1490
rect 10560 1440 10590 1470
rect 10560 1420 10565 1440
rect 10585 1420 10590 1440
rect 10560 1390 10590 1420
rect 10560 1370 10565 1390
rect 10585 1370 10590 1390
rect 10560 1340 10590 1370
rect 10560 1320 10565 1340
rect 10585 1320 10590 1340
rect 10560 1290 10590 1320
rect 10560 1270 10565 1290
rect 10585 1270 10590 1290
rect 10560 1240 10590 1270
rect 10560 1220 10565 1240
rect 10585 1220 10590 1240
rect 10560 1190 10590 1220
rect 10560 1170 10565 1190
rect 10585 1170 10590 1190
rect 10560 1140 10590 1170
rect 10560 1120 10565 1140
rect 10585 1120 10590 1140
rect 10560 1090 10590 1120
rect 10560 1070 10565 1090
rect 10585 1070 10590 1090
rect 10560 1040 10590 1070
rect 10560 1020 10565 1040
rect 10585 1020 10590 1040
rect 10560 990 10590 1020
rect 10560 970 10565 990
rect 10585 970 10590 990
rect 10560 960 10590 970
rect 10660 1640 10690 1650
rect 10660 1620 10665 1640
rect 10685 1620 10690 1640
rect 10660 1590 10690 1620
rect 10660 1570 10665 1590
rect 10685 1570 10690 1590
rect 10660 1540 10690 1570
rect 10660 1520 10665 1540
rect 10685 1520 10690 1540
rect 10660 1490 10690 1520
rect 10660 1470 10665 1490
rect 10685 1470 10690 1490
rect 10660 1440 10690 1470
rect 10660 1420 10665 1440
rect 10685 1420 10690 1440
rect 10660 1390 10690 1420
rect 10660 1370 10665 1390
rect 10685 1370 10690 1390
rect 10660 1340 10690 1370
rect 10660 1320 10665 1340
rect 10685 1320 10690 1340
rect 10660 1290 10690 1320
rect 10660 1270 10665 1290
rect 10685 1270 10690 1290
rect 10660 1240 10690 1270
rect 10660 1220 10665 1240
rect 10685 1220 10690 1240
rect 10660 1190 10690 1220
rect 10660 1170 10665 1190
rect 10685 1170 10690 1190
rect 10660 1140 10690 1170
rect 10660 1120 10665 1140
rect 10685 1120 10690 1140
rect 10660 1090 10690 1120
rect 10660 1070 10665 1090
rect 10685 1070 10690 1090
rect 10660 1040 10690 1070
rect 10660 1020 10665 1040
rect 10685 1020 10690 1040
rect 10660 990 10690 1020
rect 10660 970 10665 990
rect 10685 970 10690 990
rect 10660 960 10690 970
rect 10760 1640 10830 1650
rect 10760 1620 10765 1640
rect 10785 1620 10805 1640
rect 10825 1620 10830 1640
rect 10760 1590 10830 1620
rect 10760 1570 10765 1590
rect 10785 1570 10805 1590
rect 10825 1570 10830 1590
rect 10760 1540 10830 1570
rect 10760 1520 10765 1540
rect 10785 1520 10805 1540
rect 10825 1520 10830 1540
rect 10990 1630 11000 1650
rect 11020 1630 11040 1650
rect 11060 1630 11065 1650
rect 10990 1600 11065 1630
rect 10990 1580 11000 1600
rect 11020 1580 11040 1600
rect 11060 1580 11065 1600
rect 10990 1550 11065 1580
rect 10990 1530 11000 1550
rect 11020 1530 11040 1550
rect 11060 1530 11065 1550
rect 10990 1520 11065 1530
rect 11090 1650 11120 1660
rect 11090 1630 11095 1650
rect 11115 1630 11120 1650
rect 11090 1600 11120 1630
rect 11090 1580 11095 1600
rect 11115 1580 11120 1600
rect 11090 1550 11120 1580
rect 11090 1530 11095 1550
rect 11115 1530 11120 1550
rect 11090 1520 11120 1530
rect 11145 1650 11175 1660
rect 11145 1630 11150 1650
rect 11170 1630 11175 1650
rect 11145 1600 11175 1630
rect 11145 1580 11150 1600
rect 11170 1580 11175 1600
rect 11145 1550 11175 1580
rect 11145 1530 11150 1550
rect 11170 1530 11175 1550
rect 11145 1520 11175 1530
rect 11200 1650 11230 1660
rect 11200 1630 11205 1650
rect 11225 1630 11230 1650
rect 11200 1600 11230 1630
rect 11200 1580 11205 1600
rect 11225 1580 11230 1600
rect 11200 1550 11230 1580
rect 11200 1530 11205 1550
rect 11225 1530 11230 1550
rect 11200 1520 11230 1530
rect 11255 1650 11285 1660
rect 11255 1630 11260 1650
rect 11280 1630 11285 1650
rect 11255 1600 11285 1630
rect 11255 1580 11260 1600
rect 11280 1580 11285 1600
rect 11255 1550 11285 1580
rect 11255 1530 11260 1550
rect 11280 1530 11285 1550
rect 11255 1520 11285 1530
rect 11310 1650 11340 1660
rect 11310 1630 11315 1650
rect 11335 1630 11340 1650
rect 11310 1600 11340 1630
rect 11310 1580 11315 1600
rect 11335 1580 11340 1600
rect 11310 1550 11340 1580
rect 11310 1530 11315 1550
rect 11335 1530 11340 1550
rect 11310 1520 11340 1530
rect 11365 1650 11395 1660
rect 11365 1630 11370 1650
rect 11390 1630 11395 1650
rect 11365 1600 11395 1630
rect 11365 1580 11370 1600
rect 11390 1580 11395 1600
rect 11365 1550 11395 1580
rect 11365 1530 11370 1550
rect 11390 1530 11395 1550
rect 11365 1520 11395 1530
rect 11420 1650 11450 1660
rect 11420 1630 11425 1650
rect 11445 1630 11450 1650
rect 11420 1600 11450 1630
rect 11420 1580 11425 1600
rect 11445 1580 11450 1600
rect 11420 1550 11450 1580
rect 11420 1530 11425 1550
rect 11445 1530 11450 1550
rect 11420 1520 11450 1530
rect 11475 1650 11505 1660
rect 11475 1630 11480 1650
rect 11500 1630 11505 1650
rect 11475 1600 11505 1630
rect 11475 1580 11480 1600
rect 11500 1580 11505 1600
rect 11475 1550 11505 1580
rect 11475 1530 11480 1550
rect 11500 1530 11505 1550
rect 11475 1520 11505 1530
rect 11530 1650 11560 1660
rect 11530 1630 11535 1650
rect 11555 1630 11560 1650
rect 11530 1600 11560 1630
rect 11530 1580 11535 1600
rect 11555 1580 11560 1600
rect 11530 1550 11560 1580
rect 11530 1530 11535 1550
rect 11555 1530 11560 1550
rect 11530 1520 11560 1530
rect 11585 1650 11615 1660
rect 11585 1630 11590 1650
rect 11610 1630 11615 1650
rect 11585 1600 11615 1630
rect 11585 1580 11590 1600
rect 11610 1580 11615 1600
rect 11585 1550 11615 1580
rect 11585 1530 11590 1550
rect 11610 1530 11615 1550
rect 11585 1520 11615 1530
rect 11640 1650 11670 1660
rect 11640 1630 11645 1650
rect 11665 1630 11670 1650
rect 11640 1600 11670 1630
rect 11640 1580 11645 1600
rect 11665 1580 11670 1600
rect 11640 1550 11670 1580
rect 11640 1530 11645 1550
rect 11665 1530 11670 1550
rect 11640 1520 11670 1530
rect 11695 1650 11805 1660
rect 11695 1630 11700 1650
rect 11720 1630 11740 1650
rect 11760 1630 11780 1650
rect 11800 1630 11805 1650
rect 11695 1600 11805 1630
rect 11695 1580 11700 1600
rect 11720 1580 11740 1600
rect 11760 1580 11780 1600
rect 11800 1580 11805 1600
rect 11695 1550 11805 1580
rect 11695 1530 11700 1550
rect 11720 1530 11740 1550
rect 11760 1530 11780 1550
rect 11800 1530 11805 1550
rect 11695 1520 11805 1530
rect 11830 1650 11860 1660
rect 11830 1630 11835 1650
rect 11855 1630 11860 1650
rect 11830 1600 11860 1630
rect 11830 1580 11835 1600
rect 11855 1580 11860 1600
rect 11830 1550 11860 1580
rect 11830 1530 11835 1550
rect 11855 1530 11860 1550
rect 11830 1520 11860 1530
rect 11885 1650 11915 1660
rect 11885 1630 11890 1650
rect 11910 1630 11915 1650
rect 11885 1600 11915 1630
rect 11885 1580 11890 1600
rect 11910 1580 11915 1600
rect 11885 1550 11915 1580
rect 11885 1530 11890 1550
rect 11910 1530 11915 1550
rect 11885 1520 11915 1530
rect 11940 1650 11970 1660
rect 11940 1630 11945 1650
rect 11965 1630 11970 1650
rect 11940 1600 11970 1630
rect 11940 1580 11945 1600
rect 11965 1580 11970 1600
rect 11940 1550 11970 1580
rect 11940 1530 11945 1550
rect 11965 1530 11970 1550
rect 11940 1520 11970 1530
rect 11995 1650 12105 1660
rect 11995 1630 12000 1650
rect 12020 1630 12040 1650
rect 12060 1630 12080 1650
rect 12100 1630 12105 1650
rect 11995 1600 12105 1630
rect 11995 1580 12000 1600
rect 12020 1580 12040 1600
rect 12060 1580 12080 1600
rect 12100 1580 12105 1600
rect 11995 1550 12105 1580
rect 11995 1530 12000 1550
rect 12020 1530 12040 1550
rect 12060 1530 12080 1550
rect 12100 1530 12105 1550
rect 11995 1520 12105 1530
rect 12130 1650 12160 1660
rect 12130 1630 12135 1650
rect 12155 1630 12160 1650
rect 12130 1600 12160 1630
rect 12130 1580 12135 1600
rect 12155 1580 12160 1600
rect 12130 1550 12160 1580
rect 12130 1530 12135 1550
rect 12155 1530 12160 1550
rect 12130 1520 12160 1530
rect 12185 1650 12215 1660
rect 12185 1630 12190 1650
rect 12210 1630 12215 1650
rect 12185 1600 12215 1630
rect 12185 1580 12190 1600
rect 12210 1580 12215 1600
rect 12185 1550 12215 1580
rect 12185 1530 12190 1550
rect 12210 1530 12215 1550
rect 12185 1520 12215 1530
rect 12240 1650 12270 1660
rect 12240 1630 12245 1650
rect 12265 1630 12270 1650
rect 12240 1600 12270 1630
rect 12240 1580 12245 1600
rect 12265 1580 12270 1600
rect 12240 1550 12270 1580
rect 12240 1530 12245 1550
rect 12265 1530 12270 1550
rect 12240 1520 12270 1530
rect 12295 1650 12325 1660
rect 12295 1630 12300 1650
rect 12320 1630 12325 1650
rect 12295 1600 12325 1630
rect 12295 1580 12300 1600
rect 12320 1580 12325 1600
rect 12295 1550 12325 1580
rect 12295 1530 12300 1550
rect 12320 1530 12325 1550
rect 12295 1520 12325 1530
rect 12350 1650 12380 1660
rect 12350 1630 12355 1650
rect 12375 1630 12380 1650
rect 12350 1600 12380 1630
rect 12350 1580 12355 1600
rect 12375 1580 12380 1600
rect 12350 1550 12380 1580
rect 12350 1530 12355 1550
rect 12375 1530 12380 1550
rect 12350 1520 12380 1530
rect 12405 1650 12435 1660
rect 12405 1630 12410 1650
rect 12430 1630 12435 1650
rect 12405 1600 12435 1630
rect 12405 1580 12410 1600
rect 12430 1580 12435 1600
rect 12405 1550 12435 1580
rect 12405 1530 12410 1550
rect 12430 1530 12435 1550
rect 12405 1520 12435 1530
rect 12460 1650 12490 1660
rect 12460 1630 12465 1650
rect 12485 1630 12490 1650
rect 12460 1600 12490 1630
rect 12460 1580 12465 1600
rect 12485 1580 12490 1600
rect 12460 1550 12490 1580
rect 12460 1530 12465 1550
rect 12485 1530 12490 1550
rect 12460 1520 12490 1530
rect 12515 1650 12545 1660
rect 12515 1630 12520 1650
rect 12540 1630 12545 1650
rect 12515 1600 12545 1630
rect 12515 1580 12520 1600
rect 12540 1580 12545 1600
rect 12515 1550 12545 1580
rect 12515 1530 12520 1550
rect 12540 1530 12545 1550
rect 12515 1520 12545 1530
rect 12570 1650 12600 1660
rect 12570 1630 12575 1650
rect 12595 1630 12600 1650
rect 12570 1600 12600 1630
rect 12570 1580 12575 1600
rect 12595 1580 12600 1600
rect 12570 1550 12600 1580
rect 12570 1530 12575 1550
rect 12595 1530 12600 1550
rect 12570 1520 12600 1530
rect 12625 1650 12655 1660
rect 12625 1630 12630 1650
rect 12650 1630 12655 1650
rect 12625 1600 12655 1630
rect 12625 1580 12630 1600
rect 12650 1580 12655 1600
rect 12625 1550 12655 1580
rect 12625 1530 12630 1550
rect 12650 1530 12655 1550
rect 12625 1520 12655 1530
rect 12680 1650 12710 1660
rect 12680 1630 12685 1650
rect 12705 1630 12710 1650
rect 12680 1600 12710 1630
rect 12680 1580 12685 1600
rect 12705 1580 12710 1600
rect 12680 1550 12710 1580
rect 12680 1530 12685 1550
rect 12705 1530 12710 1550
rect 12680 1520 12710 1530
rect 12735 1650 12810 1660
rect 13115 1650 13135 1670
rect 13315 1650 13335 1670
rect 13515 1650 13535 1670
rect 26095 1660 26115 1725
rect 26200 1660 26220 1740
rect 26305 1735 26315 1755
rect 26335 1735 26345 1755
rect 26410 1750 26420 1770
rect 26440 1750 26450 1770
rect 26640 1770 26680 1780
rect 26410 1740 26450 1750
rect 26525 1755 26565 1765
rect 26305 1725 26345 1735
rect 26237 1710 26269 1720
rect 26237 1690 26243 1710
rect 26260 1690 26269 1710
rect 26237 1680 26269 1690
rect 26315 1660 26335 1725
rect 26420 1660 26440 1740
rect 26525 1735 26535 1755
rect 26555 1735 26565 1755
rect 26640 1750 26650 1770
rect 26670 1750 26680 1770
rect 27230 1770 27270 1780
rect 26640 1740 26680 1750
rect 27125 1755 27165 1765
rect 26525 1725 26565 1735
rect 26457 1710 26489 1720
rect 26457 1690 26463 1710
rect 26480 1690 26489 1710
rect 26457 1680 26489 1690
rect 26535 1660 26555 1725
rect 26601 1710 26633 1720
rect 26601 1690 26610 1710
rect 26627 1690 26633 1710
rect 26601 1680 26633 1690
rect 26650 1660 26670 1740
rect 27125 1735 27135 1755
rect 27155 1735 27165 1755
rect 27230 1750 27240 1770
rect 27260 1750 27270 1770
rect 27450 1770 27490 1780
rect 27230 1740 27270 1750
rect 27345 1755 27385 1765
rect 27125 1725 27165 1735
rect 26820 1710 26850 1720
rect 26820 1690 26825 1710
rect 26845 1690 26850 1710
rect 26820 1680 26850 1690
rect 26867 1710 26899 1720
rect 26867 1690 26876 1710
rect 26893 1690 26899 1710
rect 26867 1680 26899 1690
rect 26950 1710 26980 1720
rect 26950 1690 26955 1710
rect 26975 1690 26980 1710
rect 26950 1680 26980 1690
rect 26830 1660 26850 1680
rect 26950 1660 26970 1680
rect 27135 1660 27155 1725
rect 27240 1660 27260 1740
rect 27345 1735 27355 1755
rect 27375 1735 27385 1755
rect 27450 1750 27460 1770
rect 27480 1750 27490 1770
rect 27680 1770 27720 1780
rect 27450 1740 27490 1750
rect 27565 1755 27605 1765
rect 27345 1725 27385 1735
rect 27277 1710 27309 1720
rect 27277 1690 27283 1710
rect 27300 1690 27309 1710
rect 27277 1680 27309 1690
rect 27355 1660 27375 1725
rect 27460 1660 27480 1740
rect 27565 1735 27575 1755
rect 27595 1735 27605 1755
rect 27680 1750 27690 1770
rect 27710 1750 27720 1770
rect 27680 1740 27720 1750
rect 27955 1770 27960 1790
rect 27980 1770 28000 1790
rect 28020 1770 28025 1790
rect 27955 1740 28025 1770
rect 27565 1725 27605 1735
rect 27497 1710 27529 1720
rect 27497 1690 27503 1710
rect 27520 1690 27529 1710
rect 27497 1680 27529 1690
rect 27575 1660 27595 1725
rect 27641 1710 27673 1720
rect 27641 1690 27650 1710
rect 27667 1690 27673 1710
rect 27641 1680 27673 1690
rect 27690 1660 27710 1740
rect 27955 1720 27960 1740
rect 27980 1720 28000 1740
rect 28020 1720 28025 1740
rect 27955 1710 28025 1720
rect 28050 1840 28080 1850
rect 28050 1820 28055 1840
rect 28075 1820 28080 1840
rect 28050 1790 28080 1820
rect 28050 1770 28055 1790
rect 28075 1770 28080 1790
rect 28050 1740 28080 1770
rect 28050 1720 28055 1740
rect 28075 1720 28080 1740
rect 28050 1710 28080 1720
rect 28105 1840 28135 1850
rect 28105 1820 28110 1840
rect 28130 1820 28135 1840
rect 28105 1790 28135 1820
rect 28105 1770 28110 1790
rect 28130 1770 28135 1790
rect 28105 1740 28135 1770
rect 28105 1720 28110 1740
rect 28130 1720 28135 1740
rect 28105 1710 28135 1720
rect 28160 1840 28190 1850
rect 28160 1820 28165 1840
rect 28185 1820 28190 1840
rect 28160 1790 28190 1820
rect 28160 1770 28165 1790
rect 28185 1770 28190 1790
rect 28160 1740 28190 1770
rect 28160 1720 28165 1740
rect 28185 1720 28190 1740
rect 28160 1710 28190 1720
rect 28215 1840 28245 1850
rect 28215 1820 28220 1840
rect 28240 1820 28245 1840
rect 28215 1790 28245 1820
rect 28215 1770 28220 1790
rect 28240 1770 28245 1790
rect 28215 1740 28245 1770
rect 28215 1720 28220 1740
rect 28240 1720 28245 1740
rect 28215 1710 28245 1720
rect 28270 1840 28300 1850
rect 28270 1820 28275 1840
rect 28295 1820 28300 1840
rect 28270 1790 28300 1820
rect 28270 1770 28275 1790
rect 28295 1770 28300 1790
rect 28270 1740 28300 1770
rect 28270 1720 28275 1740
rect 28295 1720 28300 1740
rect 28270 1710 28300 1720
rect 28325 1840 28395 1850
rect 28325 1820 28330 1840
rect 28350 1820 28370 1840
rect 28390 1820 28395 1840
rect 28325 1790 28395 1820
rect 28325 1770 28330 1790
rect 28350 1770 28370 1790
rect 28390 1770 28395 1790
rect 28325 1740 28395 1770
rect 28325 1720 28330 1740
rect 28350 1720 28370 1740
rect 28390 1720 28395 1740
rect 28325 1710 28395 1720
rect 28115 1690 28135 1710
rect 28220 1690 28240 1710
rect 28066 1675 28098 1685
rect 25990 1650 26065 1660
rect 12735 1630 12740 1650
rect 12760 1630 12780 1650
rect 12800 1630 12810 1650
rect 12735 1600 12810 1630
rect 12735 1580 12740 1600
rect 12760 1580 12780 1600
rect 12800 1580 12810 1600
rect 12735 1550 12810 1580
rect 12735 1530 12740 1550
rect 12760 1530 12780 1550
rect 12800 1530 12810 1550
rect 12735 1520 12810 1530
rect 12970 1640 13040 1650
rect 12970 1620 12975 1640
rect 12995 1620 13015 1640
rect 13035 1620 13040 1640
rect 12970 1590 13040 1620
rect 12970 1570 12975 1590
rect 12995 1570 13015 1590
rect 13035 1570 13040 1590
rect 12970 1540 13040 1570
rect 12970 1520 12975 1540
rect 12995 1520 13015 1540
rect 13035 1520 13040 1540
rect 10760 1490 10830 1520
rect 11000 1500 11020 1520
rect 10760 1470 10765 1490
rect 10785 1470 10805 1490
rect 10825 1470 10830 1490
rect 10760 1440 10830 1470
rect 10990 1490 11030 1500
rect 10990 1470 11000 1490
rect 11020 1470 11030 1490
rect 10990 1460 11030 1470
rect 11106 1490 11138 1500
rect 11106 1470 11112 1490
rect 11129 1470 11138 1490
rect 11106 1460 11138 1470
rect 11155 1440 11175 1520
rect 11260 1440 11280 1520
rect 11305 1490 11345 1500
rect 11305 1470 11315 1490
rect 11335 1470 11345 1490
rect 11305 1460 11345 1470
rect 11370 1440 11390 1520
rect 11480 1440 11500 1520
rect 11525 1490 11565 1500
rect 11525 1470 11535 1490
rect 11555 1470 11565 1490
rect 11525 1460 11565 1470
rect 11590 1440 11610 1520
rect 11740 1500 11760 1520
rect 11830 1500 11850 1520
rect 11885 1500 11905 1520
rect 12040 1500 12060 1520
rect 11730 1490 11770 1500
rect 11730 1470 11740 1490
rect 11760 1470 11770 1490
rect 11730 1460 11770 1470
rect 11825 1490 11855 1500
rect 11825 1470 11830 1490
rect 11850 1470 11855 1490
rect 11825 1460 11855 1470
rect 11875 1490 11905 1500
rect 11875 1470 11880 1490
rect 11900 1470 11905 1490
rect 11875 1460 11905 1470
rect 11922 1490 11954 1500
rect 11922 1470 11928 1490
rect 11945 1470 11954 1490
rect 11922 1460 11954 1470
rect 12030 1490 12070 1500
rect 12030 1470 12040 1490
rect 12060 1470 12070 1490
rect 12030 1460 12070 1470
rect 12146 1490 12178 1500
rect 12146 1470 12152 1490
rect 12169 1470 12178 1490
rect 12146 1460 12178 1470
rect 12195 1440 12215 1520
rect 12300 1440 12320 1520
rect 12345 1490 12385 1500
rect 12345 1470 12355 1490
rect 12375 1470 12385 1490
rect 12345 1460 12385 1470
rect 12410 1440 12430 1520
rect 12520 1440 12540 1520
rect 12565 1490 12605 1500
rect 12565 1470 12575 1490
rect 12595 1470 12605 1490
rect 12565 1460 12605 1470
rect 12630 1440 12650 1520
rect 12780 1500 12800 1520
rect 12770 1490 12810 1500
rect 12770 1470 12780 1490
rect 12800 1470 12810 1490
rect 12770 1460 12810 1470
rect 12970 1490 13040 1520
rect 12970 1470 12975 1490
rect 12995 1470 13015 1490
rect 13035 1470 13040 1490
rect 12970 1440 13040 1470
rect 10760 1420 10765 1440
rect 10785 1420 10805 1440
rect 10825 1420 10830 1440
rect 10760 1390 10830 1420
rect 11145 1430 11185 1440
rect 11145 1410 11155 1430
rect 11175 1410 11185 1430
rect 11145 1400 11185 1410
rect 11250 1430 11290 1440
rect 11250 1410 11260 1430
rect 11280 1410 11290 1430
rect 11250 1400 11290 1410
rect 11360 1430 11400 1440
rect 11360 1410 11370 1430
rect 11390 1410 11400 1430
rect 11360 1400 11400 1410
rect 11470 1430 11510 1440
rect 11470 1410 11480 1430
rect 11500 1410 11510 1430
rect 11470 1400 11510 1410
rect 11580 1430 11620 1440
rect 11580 1410 11590 1430
rect 11610 1410 11620 1430
rect 11580 1400 11620 1410
rect 12185 1430 12225 1440
rect 12185 1410 12195 1430
rect 12215 1410 12225 1430
rect 12185 1400 12225 1410
rect 12290 1430 12330 1440
rect 12290 1410 12300 1430
rect 12320 1410 12330 1430
rect 12290 1400 12330 1410
rect 12400 1430 12440 1440
rect 12400 1410 12410 1430
rect 12430 1410 12440 1430
rect 12400 1400 12440 1410
rect 12510 1430 12550 1440
rect 12510 1410 12520 1430
rect 12540 1410 12550 1430
rect 12510 1400 12550 1410
rect 12620 1430 12660 1440
rect 12620 1410 12630 1430
rect 12650 1410 12660 1430
rect 12620 1400 12660 1410
rect 12970 1420 12975 1440
rect 12995 1420 13015 1440
rect 13035 1420 13040 1440
rect 10760 1370 10765 1390
rect 10785 1370 10805 1390
rect 10825 1370 10830 1390
rect 10760 1340 10830 1370
rect 12970 1390 13040 1420
rect 12970 1370 12975 1390
rect 12995 1370 13015 1390
rect 13035 1370 13040 1390
rect 10760 1320 10765 1340
rect 10785 1320 10805 1340
rect 10825 1320 10830 1340
rect 10760 1290 10830 1320
rect 11810 1310 11850 1350
rect 12970 1340 13040 1370
rect 12970 1320 12975 1340
rect 12995 1320 13015 1340
rect 13035 1320 13040 1340
rect 10760 1270 10765 1290
rect 10785 1270 10805 1290
rect 10825 1270 10830 1290
rect 10760 1240 10830 1270
rect 11315 1260 11355 1300
rect 11880 1260 11920 1300
rect 12970 1290 13040 1320
rect 12970 1270 12975 1290
rect 12995 1270 13015 1290
rect 13035 1270 13040 1290
rect 12595 1245 12635 1255
rect 10760 1220 10765 1240
rect 10785 1220 10805 1240
rect 10825 1220 10830 1240
rect 10760 1190 10830 1220
rect 11315 1230 11355 1240
rect 11315 1210 11325 1230
rect 11345 1210 11355 1230
rect 11315 1200 11355 1210
rect 11425 1230 11465 1240
rect 11425 1210 11435 1230
rect 11455 1210 11465 1230
rect 11425 1200 11465 1210
rect 11535 1230 11575 1240
rect 11535 1210 11545 1230
rect 11565 1210 11575 1230
rect 11535 1200 11575 1210
rect 11645 1230 11685 1240
rect 11645 1210 11655 1230
rect 11675 1210 11685 1230
rect 11645 1200 11685 1210
rect 11755 1230 11795 1240
rect 11755 1210 11765 1230
rect 11785 1210 11795 1230
rect 11755 1200 11795 1210
rect 11815 1230 11845 1240
rect 11815 1210 11820 1230
rect 11840 1210 11845 1230
rect 11815 1200 11845 1210
rect 11865 1230 11905 1240
rect 11865 1210 11875 1230
rect 11895 1210 11905 1230
rect 11865 1200 11905 1210
rect 11975 1230 12015 1240
rect 11975 1210 11985 1230
rect 12005 1210 12015 1230
rect 11975 1200 12015 1210
rect 12085 1230 12125 1240
rect 12085 1210 12095 1230
rect 12115 1210 12125 1230
rect 12085 1200 12125 1210
rect 12195 1230 12235 1240
rect 12195 1210 12205 1230
rect 12225 1210 12235 1230
rect 12195 1200 12235 1210
rect 12305 1230 12345 1240
rect 12305 1210 12315 1230
rect 12335 1210 12345 1230
rect 12305 1200 12345 1210
rect 12415 1230 12455 1240
rect 12415 1210 12425 1230
rect 12445 1210 12455 1230
rect 12415 1200 12455 1210
rect 12525 1230 12565 1240
rect 12525 1210 12535 1230
rect 12555 1210 12565 1230
rect 12595 1225 12605 1245
rect 12625 1225 12635 1245
rect 12595 1215 12635 1225
rect 12970 1240 13040 1270
rect 12970 1220 12975 1240
rect 12995 1220 13015 1240
rect 13035 1220 13040 1240
rect 12525 1200 12565 1210
rect 10760 1170 10765 1190
rect 10785 1170 10805 1190
rect 10825 1170 10830 1190
rect 11325 1180 11345 1200
rect 11435 1180 11455 1200
rect 11545 1180 11565 1200
rect 11655 1180 11675 1200
rect 11765 1180 11785 1200
rect 11875 1180 11895 1200
rect 11985 1180 12005 1200
rect 12095 1180 12115 1200
rect 12205 1180 12225 1200
rect 12315 1180 12335 1200
rect 12425 1180 12445 1200
rect 12535 1180 12555 1200
rect 12970 1190 13040 1220
rect 10760 1140 10830 1170
rect 10760 1120 10765 1140
rect 10785 1120 10805 1140
rect 10825 1120 10830 1140
rect 10760 1090 10830 1120
rect 10760 1070 10765 1090
rect 10785 1070 10805 1090
rect 10825 1070 10830 1090
rect 10760 1040 10830 1070
rect 10760 1020 10765 1040
rect 10785 1020 10805 1040
rect 10825 1020 10830 1040
rect 10760 990 10830 1020
rect 10760 970 10765 990
rect 10785 970 10805 990
rect 10825 970 10830 990
rect 10760 960 10830 970
rect 11170 1170 11240 1180
rect 11170 1150 11175 1170
rect 11195 1150 11215 1170
rect 11235 1150 11240 1170
rect 11170 1120 11240 1150
rect 11170 1100 11175 1120
rect 11195 1100 11215 1120
rect 11235 1100 11240 1120
rect 11170 1070 11240 1100
rect 11170 1050 11175 1070
rect 11195 1050 11215 1070
rect 11235 1050 11240 1070
rect 11170 1020 11240 1050
rect 11170 1000 11175 1020
rect 11195 1000 11215 1020
rect 11235 1000 11240 1020
rect 11170 970 11240 1000
rect 10125 940 10145 960
rect 10365 940 10385 960
rect 10565 940 10585 960
rect 10805 940 10825 960
rect 11170 950 11175 970
rect 11195 950 11215 970
rect 11235 950 11240 970
rect 11170 940 11240 950
rect 11265 1170 11295 1180
rect 11265 1150 11270 1170
rect 11290 1150 11295 1170
rect 11265 1120 11295 1150
rect 11265 1100 11270 1120
rect 11290 1100 11295 1120
rect 11265 1070 11295 1100
rect 11265 1050 11270 1070
rect 11290 1050 11295 1070
rect 11265 1020 11295 1050
rect 11265 1000 11270 1020
rect 11290 1000 11295 1020
rect 11265 970 11295 1000
rect 11265 950 11270 970
rect 11290 950 11295 970
rect 11265 940 11295 950
rect 11320 1170 11350 1180
rect 11320 1150 11325 1170
rect 11345 1150 11350 1170
rect 11320 1120 11350 1150
rect 11320 1100 11325 1120
rect 11345 1100 11350 1120
rect 11320 1070 11350 1100
rect 11320 1050 11325 1070
rect 11345 1050 11350 1070
rect 11320 1020 11350 1050
rect 11320 1000 11325 1020
rect 11345 1000 11350 1020
rect 11320 970 11350 1000
rect 11320 950 11325 970
rect 11345 950 11350 970
rect 11320 940 11350 950
rect 11375 1170 11405 1180
rect 11375 1150 11380 1170
rect 11400 1150 11405 1170
rect 11375 1120 11405 1150
rect 11375 1100 11380 1120
rect 11400 1100 11405 1120
rect 11375 1070 11405 1100
rect 11375 1050 11380 1070
rect 11400 1050 11405 1070
rect 11375 1020 11405 1050
rect 11375 1000 11380 1020
rect 11400 1000 11405 1020
rect 11375 970 11405 1000
rect 11375 950 11380 970
rect 11400 950 11405 970
rect 11375 940 11405 950
rect 11430 1170 11460 1180
rect 11430 1150 11435 1170
rect 11455 1150 11460 1170
rect 11430 1120 11460 1150
rect 11430 1100 11435 1120
rect 11455 1100 11460 1120
rect 11430 1070 11460 1100
rect 11430 1050 11435 1070
rect 11455 1050 11460 1070
rect 11430 1020 11460 1050
rect 11430 1000 11435 1020
rect 11455 1000 11460 1020
rect 11430 970 11460 1000
rect 11430 950 11435 970
rect 11455 950 11460 970
rect 11430 940 11460 950
rect 11485 1170 11515 1180
rect 11485 1150 11490 1170
rect 11510 1150 11515 1170
rect 11485 1120 11515 1150
rect 11485 1100 11490 1120
rect 11510 1100 11515 1120
rect 11485 1070 11515 1100
rect 11485 1050 11490 1070
rect 11510 1050 11515 1070
rect 11485 1020 11515 1050
rect 11485 1000 11490 1020
rect 11510 1000 11515 1020
rect 11485 970 11515 1000
rect 11485 950 11490 970
rect 11510 950 11515 970
rect 11485 940 11515 950
rect 11540 1170 11570 1180
rect 11540 1150 11545 1170
rect 11565 1150 11570 1170
rect 11540 1120 11570 1150
rect 11540 1100 11545 1120
rect 11565 1100 11570 1120
rect 11540 1070 11570 1100
rect 11540 1050 11545 1070
rect 11565 1050 11570 1070
rect 11540 1020 11570 1050
rect 11540 1000 11545 1020
rect 11565 1000 11570 1020
rect 11540 970 11570 1000
rect 11540 950 11545 970
rect 11565 950 11570 970
rect 11540 940 11570 950
rect 11595 1170 11625 1180
rect 11595 1150 11600 1170
rect 11620 1150 11625 1170
rect 11595 1120 11625 1150
rect 11595 1100 11600 1120
rect 11620 1100 11625 1120
rect 11595 1070 11625 1100
rect 11595 1050 11600 1070
rect 11620 1050 11625 1070
rect 11595 1020 11625 1050
rect 11595 1000 11600 1020
rect 11620 1000 11625 1020
rect 11595 970 11625 1000
rect 11595 950 11600 970
rect 11620 950 11625 970
rect 11595 940 11625 950
rect 11650 1170 11680 1180
rect 11650 1150 11655 1170
rect 11675 1150 11680 1170
rect 11650 1120 11680 1150
rect 11650 1100 11655 1120
rect 11675 1100 11680 1120
rect 11650 1070 11680 1100
rect 11650 1050 11655 1070
rect 11675 1050 11680 1070
rect 11650 1020 11680 1050
rect 11650 1000 11655 1020
rect 11675 1000 11680 1020
rect 11650 970 11680 1000
rect 11650 950 11655 970
rect 11675 950 11680 970
rect 11650 940 11680 950
rect 11705 1170 11735 1180
rect 11705 1150 11710 1170
rect 11730 1150 11735 1170
rect 11705 1120 11735 1150
rect 11705 1100 11710 1120
rect 11730 1100 11735 1120
rect 11705 1070 11735 1100
rect 11705 1050 11710 1070
rect 11730 1050 11735 1070
rect 11705 1020 11735 1050
rect 11705 1000 11710 1020
rect 11730 1000 11735 1020
rect 11705 970 11735 1000
rect 11705 950 11710 970
rect 11730 950 11735 970
rect 11705 940 11735 950
rect 11760 1170 11790 1180
rect 11760 1150 11765 1170
rect 11785 1150 11790 1170
rect 11760 1120 11790 1150
rect 11760 1100 11765 1120
rect 11785 1100 11790 1120
rect 11760 1070 11790 1100
rect 11760 1050 11765 1070
rect 11785 1050 11790 1070
rect 11760 1020 11790 1050
rect 11760 1000 11765 1020
rect 11785 1000 11790 1020
rect 11760 970 11790 1000
rect 11760 950 11765 970
rect 11785 950 11790 970
rect 11760 940 11790 950
rect 11815 1170 11845 1180
rect 11815 1150 11820 1170
rect 11840 1150 11845 1170
rect 11815 1120 11845 1150
rect 11815 1100 11820 1120
rect 11840 1100 11845 1120
rect 11815 1070 11845 1100
rect 11815 1050 11820 1070
rect 11840 1050 11845 1070
rect 11815 1020 11845 1050
rect 11815 1000 11820 1020
rect 11840 1000 11845 1020
rect 11815 970 11845 1000
rect 11815 950 11820 970
rect 11840 950 11845 970
rect 11815 940 11845 950
rect 11870 1170 11900 1180
rect 11870 1150 11875 1170
rect 11895 1150 11900 1170
rect 11870 1120 11900 1150
rect 11870 1100 11875 1120
rect 11895 1100 11900 1120
rect 11870 1070 11900 1100
rect 11870 1050 11875 1070
rect 11895 1050 11900 1070
rect 11870 1020 11900 1050
rect 11870 1000 11875 1020
rect 11895 1000 11900 1020
rect 11870 970 11900 1000
rect 11870 950 11875 970
rect 11895 950 11900 970
rect 11870 940 11900 950
rect 11925 1170 11955 1180
rect 11925 1150 11930 1170
rect 11950 1150 11955 1170
rect 11925 1120 11955 1150
rect 11925 1100 11930 1120
rect 11950 1100 11955 1120
rect 11925 1070 11955 1100
rect 11925 1050 11930 1070
rect 11950 1050 11955 1070
rect 11925 1020 11955 1050
rect 11925 1000 11930 1020
rect 11950 1000 11955 1020
rect 11925 970 11955 1000
rect 11925 950 11930 970
rect 11950 950 11955 970
rect 11925 940 11955 950
rect 11980 1170 12010 1180
rect 11980 1150 11985 1170
rect 12005 1150 12010 1170
rect 11980 1120 12010 1150
rect 11980 1100 11985 1120
rect 12005 1100 12010 1120
rect 11980 1070 12010 1100
rect 11980 1050 11985 1070
rect 12005 1050 12010 1070
rect 11980 1020 12010 1050
rect 11980 1000 11985 1020
rect 12005 1000 12010 1020
rect 11980 970 12010 1000
rect 11980 950 11985 970
rect 12005 950 12010 970
rect 11980 940 12010 950
rect 12035 1170 12065 1180
rect 12035 1150 12040 1170
rect 12060 1150 12065 1170
rect 12035 1120 12065 1150
rect 12035 1100 12040 1120
rect 12060 1100 12065 1120
rect 12035 1070 12065 1100
rect 12035 1050 12040 1070
rect 12060 1050 12065 1070
rect 12035 1020 12065 1050
rect 12035 1000 12040 1020
rect 12060 1000 12065 1020
rect 12035 970 12065 1000
rect 12035 950 12040 970
rect 12060 950 12065 970
rect 12035 940 12065 950
rect 12090 1170 12120 1180
rect 12090 1150 12095 1170
rect 12115 1150 12120 1170
rect 12090 1120 12120 1150
rect 12090 1100 12095 1120
rect 12115 1100 12120 1120
rect 12090 1070 12120 1100
rect 12090 1050 12095 1070
rect 12115 1050 12120 1070
rect 12090 1020 12120 1050
rect 12090 1000 12095 1020
rect 12115 1000 12120 1020
rect 12090 970 12120 1000
rect 12090 950 12095 970
rect 12115 950 12120 970
rect 12090 940 12120 950
rect 12145 1170 12175 1180
rect 12145 1150 12150 1170
rect 12170 1150 12175 1170
rect 12145 1120 12175 1150
rect 12145 1100 12150 1120
rect 12170 1100 12175 1120
rect 12145 1070 12175 1100
rect 12145 1050 12150 1070
rect 12170 1050 12175 1070
rect 12145 1020 12175 1050
rect 12145 1000 12150 1020
rect 12170 1000 12175 1020
rect 12145 970 12175 1000
rect 12145 950 12150 970
rect 12170 950 12175 970
rect 12145 940 12175 950
rect 12200 1170 12230 1180
rect 12200 1150 12205 1170
rect 12225 1150 12230 1170
rect 12200 1120 12230 1150
rect 12200 1100 12205 1120
rect 12225 1100 12230 1120
rect 12200 1070 12230 1100
rect 12200 1050 12205 1070
rect 12225 1050 12230 1070
rect 12200 1020 12230 1050
rect 12200 1000 12205 1020
rect 12225 1000 12230 1020
rect 12200 970 12230 1000
rect 12200 950 12205 970
rect 12225 950 12230 970
rect 12200 940 12230 950
rect 12255 1170 12285 1180
rect 12255 1150 12260 1170
rect 12280 1150 12285 1170
rect 12255 1120 12285 1150
rect 12255 1100 12260 1120
rect 12280 1100 12285 1120
rect 12255 1070 12285 1100
rect 12255 1050 12260 1070
rect 12280 1050 12285 1070
rect 12255 1020 12285 1050
rect 12255 1000 12260 1020
rect 12280 1000 12285 1020
rect 12255 970 12285 1000
rect 12255 950 12260 970
rect 12280 950 12285 970
rect 12255 940 12285 950
rect 12310 1170 12340 1180
rect 12310 1150 12315 1170
rect 12335 1150 12340 1170
rect 12310 1120 12340 1150
rect 12310 1100 12315 1120
rect 12335 1100 12340 1120
rect 12310 1070 12340 1100
rect 12310 1050 12315 1070
rect 12335 1050 12340 1070
rect 12310 1020 12340 1050
rect 12310 1000 12315 1020
rect 12335 1000 12340 1020
rect 12310 970 12340 1000
rect 12310 950 12315 970
rect 12335 950 12340 970
rect 12310 940 12340 950
rect 12365 1170 12395 1180
rect 12365 1150 12370 1170
rect 12390 1150 12395 1170
rect 12365 1120 12395 1150
rect 12365 1100 12370 1120
rect 12390 1100 12395 1120
rect 12365 1070 12395 1100
rect 12365 1050 12370 1070
rect 12390 1050 12395 1070
rect 12365 1020 12395 1050
rect 12365 1000 12370 1020
rect 12390 1000 12395 1020
rect 12365 970 12395 1000
rect 12365 950 12370 970
rect 12390 950 12395 970
rect 12365 940 12395 950
rect 12420 1170 12450 1180
rect 12420 1150 12425 1170
rect 12445 1150 12450 1170
rect 12420 1120 12450 1150
rect 12420 1100 12425 1120
rect 12445 1100 12450 1120
rect 12420 1070 12450 1100
rect 12420 1050 12425 1070
rect 12445 1050 12450 1070
rect 12420 1020 12450 1050
rect 12420 1000 12425 1020
rect 12445 1000 12450 1020
rect 12420 970 12450 1000
rect 12420 950 12425 970
rect 12445 950 12450 970
rect 12420 940 12450 950
rect 12475 1170 12505 1180
rect 12475 1150 12480 1170
rect 12500 1150 12505 1170
rect 12475 1120 12505 1150
rect 12475 1100 12480 1120
rect 12500 1100 12505 1120
rect 12475 1070 12505 1100
rect 12475 1050 12480 1070
rect 12500 1050 12505 1070
rect 12475 1020 12505 1050
rect 12475 1000 12480 1020
rect 12500 1000 12505 1020
rect 12475 970 12505 1000
rect 12475 950 12480 970
rect 12500 950 12505 970
rect 12475 940 12505 950
rect 12530 1170 12560 1180
rect 12530 1150 12535 1170
rect 12555 1150 12560 1170
rect 12530 1120 12560 1150
rect 12530 1100 12535 1120
rect 12555 1100 12560 1120
rect 12530 1070 12560 1100
rect 12530 1050 12535 1070
rect 12555 1050 12560 1070
rect 12530 1020 12560 1050
rect 12530 1000 12535 1020
rect 12555 1000 12560 1020
rect 12530 970 12560 1000
rect 12530 950 12535 970
rect 12555 950 12560 970
rect 12530 940 12560 950
rect 12585 1170 12655 1180
rect 12585 1150 12590 1170
rect 12610 1150 12630 1170
rect 12650 1150 12655 1170
rect 12585 1120 12655 1150
rect 12585 1100 12590 1120
rect 12610 1100 12630 1120
rect 12650 1100 12655 1120
rect 12585 1070 12655 1100
rect 12585 1050 12590 1070
rect 12610 1050 12630 1070
rect 12650 1050 12655 1070
rect 12585 1020 12655 1050
rect 12585 1000 12590 1020
rect 12610 1000 12630 1020
rect 12650 1000 12655 1020
rect 12585 970 12655 1000
rect 12585 950 12590 970
rect 12610 950 12630 970
rect 12650 950 12655 970
rect 12970 1170 12975 1190
rect 12995 1170 13015 1190
rect 13035 1170 13040 1190
rect 12970 1140 13040 1170
rect 12970 1120 12975 1140
rect 12995 1120 13015 1140
rect 13035 1120 13040 1140
rect 12970 1090 13040 1120
rect 12970 1070 12975 1090
rect 12995 1070 13015 1090
rect 13035 1070 13040 1090
rect 12970 1040 13040 1070
rect 12970 1020 12975 1040
rect 12995 1020 13015 1040
rect 13035 1020 13040 1040
rect 12970 990 13040 1020
rect 12970 970 12975 990
rect 12995 970 13015 990
rect 13035 970 13040 990
rect 12970 960 13040 970
rect 13110 1640 13140 1650
rect 13110 1620 13115 1640
rect 13135 1620 13140 1640
rect 13110 1590 13140 1620
rect 13110 1570 13115 1590
rect 13135 1570 13140 1590
rect 13110 1540 13140 1570
rect 13110 1520 13115 1540
rect 13135 1520 13140 1540
rect 13110 1490 13140 1520
rect 13110 1470 13115 1490
rect 13135 1470 13140 1490
rect 13110 1440 13140 1470
rect 13110 1420 13115 1440
rect 13135 1420 13140 1440
rect 13110 1390 13140 1420
rect 13110 1370 13115 1390
rect 13135 1370 13140 1390
rect 13110 1340 13140 1370
rect 13110 1320 13115 1340
rect 13135 1320 13140 1340
rect 13110 1290 13140 1320
rect 13110 1270 13115 1290
rect 13135 1270 13140 1290
rect 13110 1240 13140 1270
rect 13110 1220 13115 1240
rect 13135 1220 13140 1240
rect 13110 1190 13140 1220
rect 13110 1170 13115 1190
rect 13135 1170 13140 1190
rect 13110 1140 13140 1170
rect 13110 1120 13115 1140
rect 13135 1120 13140 1140
rect 13110 1090 13140 1120
rect 13110 1070 13115 1090
rect 13135 1070 13140 1090
rect 13110 1040 13140 1070
rect 13110 1020 13115 1040
rect 13135 1020 13140 1040
rect 13110 990 13140 1020
rect 13110 970 13115 990
rect 13135 970 13140 990
rect 13110 960 13140 970
rect 13210 1640 13240 1650
rect 13210 1620 13215 1640
rect 13235 1620 13240 1640
rect 13210 1590 13240 1620
rect 13210 1570 13215 1590
rect 13235 1570 13240 1590
rect 13210 1540 13240 1570
rect 13210 1520 13215 1540
rect 13235 1520 13240 1540
rect 13210 1490 13240 1520
rect 13210 1470 13215 1490
rect 13235 1470 13240 1490
rect 13210 1440 13240 1470
rect 13210 1420 13215 1440
rect 13235 1420 13240 1440
rect 13210 1390 13240 1420
rect 13210 1370 13215 1390
rect 13235 1370 13240 1390
rect 13210 1340 13240 1370
rect 13210 1320 13215 1340
rect 13235 1320 13240 1340
rect 13210 1290 13240 1320
rect 13210 1270 13215 1290
rect 13235 1270 13240 1290
rect 13210 1240 13240 1270
rect 13210 1220 13215 1240
rect 13235 1220 13240 1240
rect 13210 1190 13240 1220
rect 13210 1170 13215 1190
rect 13235 1170 13240 1190
rect 13210 1140 13240 1170
rect 13210 1120 13215 1140
rect 13235 1120 13240 1140
rect 13210 1090 13240 1120
rect 13210 1070 13215 1090
rect 13235 1070 13240 1090
rect 13210 1040 13240 1070
rect 13210 1020 13215 1040
rect 13235 1020 13240 1040
rect 13210 990 13240 1020
rect 13210 970 13215 990
rect 13235 970 13240 990
rect 13210 960 13240 970
rect 13310 1640 13340 1650
rect 13310 1620 13315 1640
rect 13335 1620 13340 1640
rect 13310 1590 13340 1620
rect 13310 1570 13315 1590
rect 13335 1570 13340 1590
rect 13310 1540 13340 1570
rect 13310 1520 13315 1540
rect 13335 1520 13340 1540
rect 13310 1490 13340 1520
rect 13310 1470 13315 1490
rect 13335 1470 13340 1490
rect 13310 1440 13340 1470
rect 13310 1420 13315 1440
rect 13335 1420 13340 1440
rect 13310 1390 13340 1420
rect 13310 1370 13315 1390
rect 13335 1370 13340 1390
rect 13310 1340 13340 1370
rect 13310 1320 13315 1340
rect 13335 1320 13340 1340
rect 13310 1290 13340 1320
rect 13310 1270 13315 1290
rect 13335 1270 13340 1290
rect 13310 1240 13340 1270
rect 13310 1220 13315 1240
rect 13335 1220 13340 1240
rect 13310 1190 13340 1220
rect 13310 1170 13315 1190
rect 13335 1170 13340 1190
rect 13310 1140 13340 1170
rect 13310 1120 13315 1140
rect 13335 1120 13340 1140
rect 13310 1090 13340 1120
rect 13310 1070 13315 1090
rect 13335 1070 13340 1090
rect 13310 1040 13340 1070
rect 13310 1020 13315 1040
rect 13335 1020 13340 1040
rect 13310 990 13340 1020
rect 13310 970 13315 990
rect 13335 970 13340 990
rect 13310 960 13340 970
rect 13410 1640 13440 1650
rect 13410 1620 13415 1640
rect 13435 1620 13440 1640
rect 13410 1590 13440 1620
rect 13410 1570 13415 1590
rect 13435 1570 13440 1590
rect 13410 1540 13440 1570
rect 13410 1520 13415 1540
rect 13435 1520 13440 1540
rect 13410 1490 13440 1520
rect 13410 1470 13415 1490
rect 13435 1470 13440 1490
rect 13410 1440 13440 1470
rect 13410 1420 13415 1440
rect 13435 1420 13440 1440
rect 13410 1390 13440 1420
rect 13410 1370 13415 1390
rect 13435 1370 13440 1390
rect 13410 1340 13440 1370
rect 13410 1320 13415 1340
rect 13435 1320 13440 1340
rect 13410 1290 13440 1320
rect 13410 1270 13415 1290
rect 13435 1270 13440 1290
rect 13410 1240 13440 1270
rect 13410 1220 13415 1240
rect 13435 1220 13440 1240
rect 13410 1190 13440 1220
rect 13410 1170 13415 1190
rect 13435 1170 13440 1190
rect 13410 1140 13440 1170
rect 13410 1120 13415 1140
rect 13435 1120 13440 1140
rect 13410 1090 13440 1120
rect 13410 1070 13415 1090
rect 13435 1070 13440 1090
rect 13410 1040 13440 1070
rect 13410 1020 13415 1040
rect 13435 1020 13440 1040
rect 13410 990 13440 1020
rect 13410 970 13415 990
rect 13435 970 13440 990
rect 13410 960 13440 970
rect 13510 1640 13540 1650
rect 13510 1620 13515 1640
rect 13535 1620 13540 1640
rect 13510 1590 13540 1620
rect 13510 1570 13515 1590
rect 13535 1570 13540 1590
rect 13510 1540 13540 1570
rect 13510 1520 13515 1540
rect 13535 1520 13540 1540
rect 13510 1490 13540 1520
rect 13510 1470 13515 1490
rect 13535 1470 13540 1490
rect 13510 1440 13540 1470
rect 13510 1420 13515 1440
rect 13535 1420 13540 1440
rect 13510 1390 13540 1420
rect 13510 1370 13515 1390
rect 13535 1370 13540 1390
rect 13510 1340 13540 1370
rect 13510 1320 13515 1340
rect 13535 1320 13540 1340
rect 13510 1290 13540 1320
rect 13510 1270 13515 1290
rect 13535 1270 13540 1290
rect 13510 1240 13540 1270
rect 13510 1220 13515 1240
rect 13535 1220 13540 1240
rect 13510 1190 13540 1220
rect 13510 1170 13515 1190
rect 13535 1170 13540 1190
rect 13510 1140 13540 1170
rect 13510 1120 13515 1140
rect 13535 1120 13540 1140
rect 13510 1090 13540 1120
rect 13510 1070 13515 1090
rect 13535 1070 13540 1090
rect 13510 1040 13540 1070
rect 13510 1020 13515 1040
rect 13535 1020 13540 1040
rect 13510 990 13540 1020
rect 13510 970 13515 990
rect 13535 970 13540 990
rect 13510 960 13540 970
rect 13610 1640 13680 1650
rect 13610 1620 13615 1640
rect 13635 1620 13655 1640
rect 13675 1620 13680 1640
rect 13610 1590 13680 1620
rect 13610 1570 13615 1590
rect 13635 1570 13655 1590
rect 13675 1570 13680 1590
rect 13610 1540 13680 1570
rect 13610 1520 13615 1540
rect 13635 1520 13655 1540
rect 13675 1520 13680 1540
rect 13610 1490 13680 1520
rect 13610 1470 13615 1490
rect 13635 1470 13655 1490
rect 13675 1470 13680 1490
rect 13610 1440 13680 1470
rect 13610 1420 13615 1440
rect 13635 1420 13655 1440
rect 13675 1420 13680 1440
rect 13610 1390 13680 1420
rect 13610 1370 13615 1390
rect 13635 1370 13655 1390
rect 13675 1370 13680 1390
rect 13735 1640 13770 1650
rect 13735 1615 13740 1640
rect 13765 1615 13770 1640
rect 13735 1605 13770 1615
rect 13795 1640 13830 1650
rect 13795 1615 13800 1640
rect 13825 1615 13830 1640
rect 13795 1605 13830 1615
rect 25990 1630 26000 1650
rect 26020 1630 26040 1650
rect 26060 1630 26065 1650
rect 25990 1600 26065 1630
rect 25990 1580 26000 1600
rect 26020 1580 26040 1600
rect 26060 1580 26065 1600
rect 25990 1550 26065 1580
rect 25990 1530 26000 1550
rect 26020 1530 26040 1550
rect 26060 1530 26065 1550
rect 25990 1520 26065 1530
rect 26090 1650 26120 1660
rect 26090 1630 26095 1650
rect 26115 1630 26120 1650
rect 26090 1600 26120 1630
rect 26090 1580 26095 1600
rect 26115 1580 26120 1600
rect 26090 1550 26120 1580
rect 26090 1530 26095 1550
rect 26115 1530 26120 1550
rect 26090 1520 26120 1530
rect 26145 1650 26175 1660
rect 26145 1630 26150 1650
rect 26170 1630 26175 1650
rect 26145 1600 26175 1630
rect 26145 1580 26150 1600
rect 26170 1580 26175 1600
rect 26145 1550 26175 1580
rect 26145 1530 26150 1550
rect 26170 1530 26175 1550
rect 26145 1520 26175 1530
rect 26200 1650 26230 1660
rect 26200 1630 26205 1650
rect 26225 1630 26230 1650
rect 26200 1600 26230 1630
rect 26200 1580 26205 1600
rect 26225 1580 26230 1600
rect 26200 1550 26230 1580
rect 26200 1530 26205 1550
rect 26225 1530 26230 1550
rect 26200 1520 26230 1530
rect 26255 1650 26285 1660
rect 26255 1630 26260 1650
rect 26280 1630 26285 1650
rect 26255 1600 26285 1630
rect 26255 1580 26260 1600
rect 26280 1580 26285 1600
rect 26255 1550 26285 1580
rect 26255 1530 26260 1550
rect 26280 1530 26285 1550
rect 26255 1520 26285 1530
rect 26310 1650 26340 1660
rect 26310 1630 26315 1650
rect 26335 1630 26340 1650
rect 26310 1600 26340 1630
rect 26310 1580 26315 1600
rect 26335 1580 26340 1600
rect 26310 1550 26340 1580
rect 26310 1530 26315 1550
rect 26335 1530 26340 1550
rect 26310 1520 26340 1530
rect 26365 1650 26395 1660
rect 26365 1630 26370 1650
rect 26390 1630 26395 1650
rect 26365 1600 26395 1630
rect 26365 1580 26370 1600
rect 26390 1580 26395 1600
rect 26365 1550 26395 1580
rect 26365 1530 26370 1550
rect 26390 1530 26395 1550
rect 26365 1520 26395 1530
rect 26420 1650 26450 1660
rect 26420 1630 26425 1650
rect 26445 1630 26450 1650
rect 26420 1600 26450 1630
rect 26420 1580 26425 1600
rect 26445 1580 26450 1600
rect 26420 1550 26450 1580
rect 26420 1530 26425 1550
rect 26445 1530 26450 1550
rect 26420 1520 26450 1530
rect 26475 1650 26505 1660
rect 26475 1630 26480 1650
rect 26500 1630 26505 1650
rect 26475 1600 26505 1630
rect 26475 1580 26480 1600
rect 26500 1580 26505 1600
rect 26475 1550 26505 1580
rect 26475 1530 26480 1550
rect 26500 1530 26505 1550
rect 26475 1520 26505 1530
rect 26530 1650 26560 1660
rect 26530 1630 26535 1650
rect 26555 1630 26560 1650
rect 26530 1600 26560 1630
rect 26530 1580 26535 1600
rect 26555 1580 26560 1600
rect 26530 1550 26560 1580
rect 26530 1530 26535 1550
rect 26555 1530 26560 1550
rect 26530 1520 26560 1530
rect 26585 1650 26615 1660
rect 26585 1630 26590 1650
rect 26610 1630 26615 1650
rect 26585 1600 26615 1630
rect 26585 1580 26590 1600
rect 26610 1580 26615 1600
rect 26585 1550 26615 1580
rect 26585 1530 26590 1550
rect 26610 1530 26615 1550
rect 26585 1520 26615 1530
rect 26640 1650 26670 1660
rect 26640 1630 26645 1650
rect 26665 1630 26670 1650
rect 26640 1600 26670 1630
rect 26640 1580 26645 1600
rect 26665 1580 26670 1600
rect 26640 1550 26670 1580
rect 26640 1530 26645 1550
rect 26665 1530 26670 1550
rect 26640 1520 26670 1530
rect 26695 1650 26805 1660
rect 26695 1630 26700 1650
rect 26720 1630 26740 1650
rect 26760 1630 26780 1650
rect 26800 1630 26805 1650
rect 26695 1600 26805 1630
rect 26695 1580 26700 1600
rect 26720 1580 26740 1600
rect 26760 1580 26780 1600
rect 26800 1580 26805 1600
rect 26695 1550 26805 1580
rect 26695 1530 26700 1550
rect 26720 1530 26740 1550
rect 26760 1530 26780 1550
rect 26800 1530 26805 1550
rect 26695 1520 26805 1530
rect 26830 1650 26860 1660
rect 26830 1630 26835 1650
rect 26855 1630 26860 1650
rect 26830 1600 26860 1630
rect 26830 1580 26835 1600
rect 26855 1580 26860 1600
rect 26830 1550 26860 1580
rect 26830 1530 26835 1550
rect 26855 1530 26860 1550
rect 26830 1520 26860 1530
rect 26885 1650 26915 1660
rect 26885 1630 26890 1650
rect 26910 1630 26915 1650
rect 26885 1600 26915 1630
rect 26885 1580 26890 1600
rect 26910 1580 26915 1600
rect 26885 1550 26915 1580
rect 26885 1530 26890 1550
rect 26910 1530 26915 1550
rect 26885 1520 26915 1530
rect 26940 1650 26970 1660
rect 26940 1630 26945 1650
rect 26965 1630 26970 1650
rect 26940 1600 26970 1630
rect 26940 1580 26945 1600
rect 26965 1580 26970 1600
rect 26940 1550 26970 1580
rect 26940 1530 26945 1550
rect 26965 1530 26970 1550
rect 26940 1520 26970 1530
rect 26995 1650 27105 1660
rect 26995 1630 27000 1650
rect 27020 1630 27040 1650
rect 27060 1630 27080 1650
rect 27100 1630 27105 1650
rect 26995 1600 27105 1630
rect 26995 1580 27000 1600
rect 27020 1580 27040 1600
rect 27060 1580 27080 1600
rect 27100 1580 27105 1600
rect 26995 1550 27105 1580
rect 26995 1530 27000 1550
rect 27020 1530 27040 1550
rect 27060 1530 27080 1550
rect 27100 1530 27105 1550
rect 26995 1520 27105 1530
rect 27130 1650 27160 1660
rect 27130 1630 27135 1650
rect 27155 1630 27160 1650
rect 27130 1600 27160 1630
rect 27130 1580 27135 1600
rect 27155 1580 27160 1600
rect 27130 1550 27160 1580
rect 27130 1530 27135 1550
rect 27155 1530 27160 1550
rect 27130 1520 27160 1530
rect 27185 1650 27215 1660
rect 27185 1630 27190 1650
rect 27210 1630 27215 1650
rect 27185 1600 27215 1630
rect 27185 1580 27190 1600
rect 27210 1580 27215 1600
rect 27185 1550 27215 1580
rect 27185 1530 27190 1550
rect 27210 1530 27215 1550
rect 27185 1520 27215 1530
rect 27240 1650 27270 1660
rect 27240 1630 27245 1650
rect 27265 1630 27270 1650
rect 27240 1600 27270 1630
rect 27240 1580 27245 1600
rect 27265 1580 27270 1600
rect 27240 1550 27270 1580
rect 27240 1530 27245 1550
rect 27265 1530 27270 1550
rect 27240 1520 27270 1530
rect 27295 1650 27325 1660
rect 27295 1630 27300 1650
rect 27320 1630 27325 1650
rect 27295 1600 27325 1630
rect 27295 1580 27300 1600
rect 27320 1580 27325 1600
rect 27295 1550 27325 1580
rect 27295 1530 27300 1550
rect 27320 1530 27325 1550
rect 27295 1520 27325 1530
rect 27350 1650 27380 1660
rect 27350 1630 27355 1650
rect 27375 1630 27380 1650
rect 27350 1600 27380 1630
rect 27350 1580 27355 1600
rect 27375 1580 27380 1600
rect 27350 1550 27380 1580
rect 27350 1530 27355 1550
rect 27375 1530 27380 1550
rect 27350 1520 27380 1530
rect 27405 1650 27435 1660
rect 27405 1630 27410 1650
rect 27430 1630 27435 1650
rect 27405 1600 27435 1630
rect 27405 1580 27410 1600
rect 27430 1580 27435 1600
rect 27405 1550 27435 1580
rect 27405 1530 27410 1550
rect 27430 1530 27435 1550
rect 27405 1520 27435 1530
rect 27460 1650 27490 1660
rect 27460 1630 27465 1650
rect 27485 1630 27490 1650
rect 27460 1600 27490 1630
rect 27460 1580 27465 1600
rect 27485 1580 27490 1600
rect 27460 1550 27490 1580
rect 27460 1530 27465 1550
rect 27485 1530 27490 1550
rect 27460 1520 27490 1530
rect 27515 1650 27545 1660
rect 27515 1630 27520 1650
rect 27540 1630 27545 1650
rect 27515 1600 27545 1630
rect 27515 1580 27520 1600
rect 27540 1580 27545 1600
rect 27515 1550 27545 1580
rect 27515 1530 27520 1550
rect 27540 1530 27545 1550
rect 27515 1520 27545 1530
rect 27570 1650 27600 1660
rect 27570 1630 27575 1650
rect 27595 1630 27600 1650
rect 27570 1600 27600 1630
rect 27570 1580 27575 1600
rect 27595 1580 27600 1600
rect 27570 1550 27600 1580
rect 27570 1530 27575 1550
rect 27595 1530 27600 1550
rect 27570 1520 27600 1530
rect 27625 1650 27655 1660
rect 27625 1630 27630 1650
rect 27650 1630 27655 1650
rect 27625 1600 27655 1630
rect 27625 1580 27630 1600
rect 27650 1580 27655 1600
rect 27625 1550 27655 1580
rect 27625 1530 27630 1550
rect 27650 1530 27655 1550
rect 27625 1520 27655 1530
rect 27680 1650 27710 1660
rect 27680 1630 27685 1650
rect 27705 1630 27710 1650
rect 27680 1600 27710 1630
rect 27680 1580 27685 1600
rect 27705 1580 27710 1600
rect 27680 1550 27710 1580
rect 27680 1530 27685 1550
rect 27705 1530 27710 1550
rect 27680 1520 27710 1530
rect 27735 1650 27810 1660
rect 27735 1630 27740 1650
rect 27760 1630 27780 1650
rect 27800 1630 27810 1650
rect 28066 1655 28071 1675
rect 28091 1655 28098 1675
rect 28066 1645 28098 1655
rect 28115 1680 28155 1690
rect 28115 1660 28125 1680
rect 28145 1660 28155 1680
rect 28115 1650 28155 1660
rect 28210 1680 28250 1690
rect 28210 1660 28220 1680
rect 28240 1660 28250 1680
rect 28210 1650 28250 1660
rect 27735 1600 27810 1630
rect 27735 1580 27740 1600
rect 27760 1580 27780 1600
rect 27800 1580 27810 1600
rect 28010 1625 28050 1635
rect 28010 1605 28020 1625
rect 28040 1605 28050 1625
rect 28010 1595 28050 1605
rect 28300 1625 28340 1635
rect 28300 1605 28310 1625
rect 28330 1605 28340 1625
rect 28300 1595 28340 1605
rect 27735 1550 27810 1580
rect 27735 1530 27740 1550
rect 27760 1530 27780 1550
rect 27800 1530 27810 1550
rect 27971 1565 28003 1575
rect 27971 1545 27976 1565
rect 27996 1545 28003 1565
rect 27971 1535 28003 1545
rect 27735 1520 27810 1530
rect 26000 1500 26020 1520
rect 25990 1490 26030 1500
rect 25990 1470 26000 1490
rect 26020 1470 26030 1490
rect 25990 1460 26030 1470
rect 26106 1490 26138 1500
rect 26106 1470 26112 1490
rect 26129 1470 26138 1490
rect 26106 1460 26138 1470
rect 26155 1440 26175 1520
rect 26260 1440 26280 1520
rect 26305 1490 26345 1500
rect 26305 1470 26315 1490
rect 26335 1470 26345 1490
rect 26305 1460 26345 1470
rect 26370 1440 26390 1520
rect 26480 1440 26500 1520
rect 26525 1490 26565 1500
rect 26525 1470 26535 1490
rect 26555 1470 26565 1490
rect 26525 1460 26565 1470
rect 26590 1440 26610 1520
rect 26740 1500 26760 1520
rect 26830 1500 26850 1520
rect 26885 1500 26905 1520
rect 27040 1500 27060 1520
rect 26730 1490 26770 1500
rect 26730 1470 26740 1490
rect 26760 1470 26770 1490
rect 26730 1460 26770 1470
rect 26825 1490 26855 1500
rect 26825 1470 26830 1490
rect 26850 1470 26855 1490
rect 26825 1460 26855 1470
rect 26875 1490 26905 1500
rect 26875 1470 26880 1490
rect 26900 1470 26905 1490
rect 26875 1460 26905 1470
rect 26922 1490 26954 1500
rect 26922 1470 26928 1490
rect 26945 1470 26954 1490
rect 26922 1460 26954 1470
rect 27030 1490 27070 1500
rect 27030 1470 27040 1490
rect 27060 1470 27070 1490
rect 27030 1460 27070 1470
rect 27146 1490 27178 1500
rect 27146 1470 27152 1490
rect 27169 1470 27178 1490
rect 27146 1460 27178 1470
rect 27195 1440 27215 1520
rect 27300 1440 27320 1520
rect 27345 1490 27385 1500
rect 27345 1470 27355 1490
rect 27375 1470 27385 1490
rect 27345 1460 27385 1470
rect 27410 1440 27430 1520
rect 27520 1440 27540 1520
rect 27565 1490 27605 1500
rect 27565 1470 27575 1490
rect 27595 1470 27605 1490
rect 27565 1460 27605 1470
rect 27630 1440 27650 1520
rect 27780 1500 27800 1520
rect 28020 1515 28040 1595
rect 28060 1565 28100 1575
rect 28060 1545 28070 1565
rect 28090 1545 28100 1565
rect 28060 1535 28100 1545
rect 28070 1515 28090 1535
rect 28310 1515 28330 1595
rect 28347 1565 28379 1575
rect 28347 1545 28354 1565
rect 28374 1545 28379 1565
rect 28347 1535 28379 1545
rect 27855 1505 27930 1515
rect 27770 1490 27810 1500
rect 27770 1470 27780 1490
rect 27800 1470 27810 1490
rect 27770 1460 27810 1470
rect 27855 1485 27865 1505
rect 27885 1485 27905 1505
rect 27925 1485 27930 1505
rect 27855 1455 27930 1485
rect 26145 1430 26185 1440
rect 26145 1410 26155 1430
rect 26175 1410 26185 1430
rect 26145 1400 26185 1410
rect 26250 1430 26290 1440
rect 26250 1410 26260 1430
rect 26280 1410 26290 1430
rect 26250 1400 26290 1410
rect 26360 1430 26400 1440
rect 26360 1410 26370 1430
rect 26390 1410 26400 1430
rect 26360 1400 26400 1410
rect 26470 1430 26510 1440
rect 26470 1410 26480 1430
rect 26500 1410 26510 1430
rect 26470 1400 26510 1410
rect 26580 1430 26620 1440
rect 26580 1410 26590 1430
rect 26610 1410 26620 1430
rect 26580 1400 26620 1410
rect 27185 1430 27225 1440
rect 27185 1410 27195 1430
rect 27215 1410 27225 1430
rect 27185 1400 27225 1410
rect 27290 1430 27330 1440
rect 27290 1410 27300 1430
rect 27320 1410 27330 1430
rect 27290 1400 27330 1410
rect 27400 1430 27440 1440
rect 27400 1410 27410 1430
rect 27430 1410 27440 1430
rect 27400 1400 27440 1410
rect 27510 1430 27550 1440
rect 27510 1410 27520 1430
rect 27540 1410 27550 1430
rect 27510 1400 27550 1410
rect 27620 1430 27660 1440
rect 27620 1410 27630 1430
rect 27650 1410 27660 1430
rect 27620 1400 27660 1410
rect 27855 1435 27865 1455
rect 27885 1435 27905 1455
rect 27925 1435 27930 1455
rect 27855 1405 27930 1435
rect 13610 1340 13680 1370
rect 26810 1350 26850 1390
rect 27855 1385 27865 1405
rect 27885 1385 27905 1405
rect 27925 1385 27930 1405
rect 27855 1375 27930 1385
rect 27955 1505 27985 1515
rect 27955 1485 27960 1505
rect 27980 1485 27985 1505
rect 27955 1455 27985 1485
rect 27955 1435 27960 1455
rect 27980 1435 27985 1455
rect 27955 1405 27985 1435
rect 27955 1385 27960 1405
rect 27980 1385 27985 1405
rect 27955 1375 27985 1385
rect 28010 1505 28040 1515
rect 28010 1485 28015 1505
rect 28035 1485 28040 1505
rect 28010 1455 28040 1485
rect 28010 1435 28015 1455
rect 28035 1435 28040 1455
rect 28010 1405 28040 1435
rect 28010 1385 28015 1405
rect 28035 1385 28040 1405
rect 28010 1375 28040 1385
rect 28065 1505 28095 1515
rect 28065 1485 28070 1505
rect 28090 1485 28095 1505
rect 28065 1455 28095 1485
rect 28065 1435 28070 1455
rect 28090 1435 28095 1455
rect 28065 1405 28095 1435
rect 28065 1385 28070 1405
rect 28090 1385 28095 1405
rect 28065 1375 28095 1385
rect 28120 1505 28230 1515
rect 28120 1485 28125 1505
rect 28145 1485 28165 1505
rect 28185 1485 28205 1505
rect 28225 1485 28230 1505
rect 28120 1455 28230 1485
rect 28120 1435 28125 1455
rect 28145 1435 28165 1455
rect 28185 1435 28205 1455
rect 28225 1435 28230 1455
rect 28120 1405 28230 1435
rect 28120 1385 28125 1405
rect 28145 1385 28165 1405
rect 28185 1385 28205 1405
rect 28225 1385 28230 1405
rect 28120 1375 28230 1385
rect 28255 1505 28285 1515
rect 28255 1485 28260 1505
rect 28280 1485 28285 1505
rect 28255 1455 28285 1485
rect 28255 1435 28260 1455
rect 28280 1435 28285 1455
rect 28255 1405 28285 1435
rect 28255 1385 28260 1405
rect 28280 1385 28285 1405
rect 28255 1375 28285 1385
rect 28310 1505 28340 1515
rect 28310 1485 28315 1505
rect 28335 1485 28340 1505
rect 28310 1455 28340 1485
rect 28310 1435 28315 1455
rect 28335 1435 28340 1455
rect 28310 1405 28340 1435
rect 28310 1385 28315 1405
rect 28335 1385 28340 1405
rect 28310 1375 28340 1385
rect 28365 1505 28395 1515
rect 28365 1485 28370 1505
rect 28390 1485 28395 1505
rect 28365 1455 28395 1485
rect 28365 1435 28370 1455
rect 28390 1435 28395 1455
rect 28365 1405 28395 1435
rect 28365 1385 28370 1405
rect 28390 1385 28395 1405
rect 28365 1375 28395 1385
rect 28420 1505 28495 1515
rect 28420 1485 28425 1505
rect 28445 1485 28465 1505
rect 28485 1485 28495 1505
rect 28420 1455 28495 1485
rect 28420 1435 28425 1455
rect 28445 1435 28465 1455
rect 28485 1435 28495 1455
rect 28420 1405 28495 1435
rect 28420 1385 28425 1405
rect 28445 1385 28465 1405
rect 28485 1385 28495 1405
rect 28420 1375 28495 1385
rect 27865 1355 27885 1375
rect 27855 1345 27895 1355
rect 13610 1320 13615 1340
rect 13635 1320 13655 1340
rect 13675 1320 13680 1340
rect 13610 1290 13680 1320
rect 26315 1300 26355 1340
rect 26880 1300 26920 1340
rect 27855 1325 27865 1345
rect 27885 1325 27895 1345
rect 27855 1315 27895 1325
rect 27955 1295 27975 1375
rect 28026 1345 28058 1355
rect 28026 1325 28033 1345
rect 28053 1325 28058 1345
rect 28026 1315 28058 1325
rect 28075 1295 28095 1375
rect 28165 1355 28185 1375
rect 28155 1345 28195 1355
rect 28155 1325 28165 1345
rect 28185 1325 28195 1345
rect 28155 1315 28195 1325
rect 28255 1295 28275 1375
rect 28292 1345 28324 1355
rect 28292 1325 28297 1345
rect 28317 1325 28324 1345
rect 28292 1315 28324 1325
rect 28375 1295 28395 1375
rect 28465 1355 28485 1375
rect 28455 1345 28495 1355
rect 28455 1325 28465 1345
rect 28485 1325 28495 1345
rect 28455 1315 28495 1325
rect 13610 1270 13615 1290
rect 13635 1270 13655 1290
rect 13675 1270 13680 1290
rect 27595 1285 27635 1295
rect 13610 1240 13680 1270
rect 26315 1270 26355 1280
rect 26315 1250 26325 1270
rect 26345 1250 26355 1270
rect 26315 1240 26355 1250
rect 26425 1270 26465 1280
rect 26425 1250 26435 1270
rect 26455 1250 26465 1270
rect 26425 1240 26465 1250
rect 26535 1270 26575 1280
rect 26535 1250 26545 1270
rect 26565 1250 26575 1270
rect 26535 1240 26575 1250
rect 26645 1270 26685 1280
rect 26645 1250 26655 1270
rect 26675 1250 26685 1270
rect 26645 1240 26685 1250
rect 26755 1270 26795 1280
rect 26755 1250 26765 1270
rect 26785 1250 26795 1270
rect 26755 1240 26795 1250
rect 26815 1270 26845 1280
rect 26815 1250 26820 1270
rect 26840 1250 26845 1270
rect 26815 1240 26845 1250
rect 26865 1270 26905 1280
rect 26865 1250 26875 1270
rect 26895 1250 26905 1270
rect 26865 1240 26905 1250
rect 26975 1270 27015 1280
rect 26975 1250 26985 1270
rect 27005 1250 27015 1270
rect 26975 1240 27015 1250
rect 27085 1270 27125 1280
rect 27085 1250 27095 1270
rect 27115 1250 27125 1270
rect 27085 1240 27125 1250
rect 27195 1270 27235 1280
rect 27195 1250 27205 1270
rect 27225 1250 27235 1270
rect 27195 1240 27235 1250
rect 27305 1270 27345 1280
rect 27305 1250 27315 1270
rect 27335 1250 27345 1270
rect 27305 1240 27345 1250
rect 27415 1270 27455 1280
rect 27415 1250 27425 1270
rect 27445 1250 27455 1270
rect 27415 1240 27455 1250
rect 27525 1270 27565 1280
rect 27525 1250 27535 1270
rect 27555 1250 27565 1270
rect 27595 1265 27605 1285
rect 27625 1265 27635 1285
rect 27595 1255 27635 1265
rect 27945 1285 27985 1295
rect 27945 1265 27955 1285
rect 27975 1265 27985 1285
rect 27945 1255 27985 1265
rect 28060 1285 28100 1295
rect 28060 1265 28070 1285
rect 28090 1265 28100 1285
rect 28060 1255 28100 1265
rect 28250 1285 28290 1295
rect 28250 1265 28260 1285
rect 28280 1265 28290 1285
rect 28250 1255 28290 1265
rect 28365 1285 28405 1295
rect 28365 1265 28375 1285
rect 28395 1265 28405 1285
rect 28365 1255 28405 1265
rect 27525 1240 27565 1250
rect 13610 1220 13615 1240
rect 13635 1220 13655 1240
rect 13675 1220 13680 1240
rect 26325 1220 26345 1240
rect 26435 1220 26455 1240
rect 26545 1220 26565 1240
rect 26655 1220 26675 1240
rect 26765 1220 26785 1240
rect 26875 1220 26895 1240
rect 26985 1220 27005 1240
rect 27095 1220 27115 1240
rect 27205 1220 27225 1240
rect 27315 1220 27335 1240
rect 27425 1220 27445 1240
rect 27535 1220 27555 1240
rect 28100 1225 28140 1235
rect 13610 1190 13680 1220
rect 13610 1170 13615 1190
rect 13635 1170 13655 1190
rect 13675 1170 13680 1190
rect 13610 1140 13680 1170
rect 13610 1120 13615 1140
rect 13635 1120 13655 1140
rect 13675 1120 13680 1140
rect 26170 1210 26240 1220
rect 26170 1190 26175 1210
rect 26195 1190 26215 1210
rect 26235 1190 26240 1210
rect 26170 1160 26240 1190
rect 26170 1140 26175 1160
rect 26195 1140 26215 1160
rect 26235 1140 26240 1160
rect 13610 1090 13680 1120
rect 13610 1070 13615 1090
rect 13635 1070 13655 1090
rect 13675 1070 13680 1090
rect 13610 1040 13680 1070
rect 13610 1020 13615 1040
rect 13635 1020 13655 1040
rect 13675 1020 13680 1040
rect 13610 990 13680 1020
rect 13610 970 13615 990
rect 13635 970 13655 990
rect 13675 970 13680 990
rect 13610 960 13680 970
rect 12585 940 12655 950
rect 12975 940 12995 960
rect 13215 940 13235 960
rect 13415 940 13435 960
rect 13655 940 13675 960
rect 10115 930 10155 940
rect 10115 910 10125 930
rect 10145 910 10155 930
rect 4975 895 5015 905
rect 10115 900 10155 910
rect 10355 930 10395 940
rect 10355 910 10365 930
rect 10385 910 10395 930
rect 10355 900 10395 910
rect 10555 930 10595 940
rect 10555 910 10565 930
rect 10585 910 10595 930
rect 10555 900 10595 910
rect 10795 930 10835 940
rect 10795 910 10805 930
rect 10825 910 10835 930
rect 11175 920 11195 940
rect 11270 920 11290 940
rect 11380 920 11400 940
rect 11490 920 11510 940
rect 11600 920 11620 940
rect 11710 920 11730 940
rect 11820 920 11840 940
rect 11930 920 11950 940
rect 12040 920 12060 940
rect 12150 920 12170 940
rect 12260 920 12280 940
rect 12370 920 12390 940
rect 12480 920 12500 940
rect 12630 920 12650 940
rect 12965 930 13005 940
rect 10795 900 10835 910
rect 11165 910 11205 920
rect 3005 875 3025 895
rect 3185 875 3205 895
rect 3365 875 3385 895
rect 3545 875 3565 895
rect 3725 875 3745 895
rect 3905 875 3925 895
rect 4085 875 4105 895
rect 4265 875 4285 895
rect 4445 875 4465 895
rect 4625 875 4645 895
rect 4805 875 4825 895
rect 4985 875 5005 895
rect 11165 890 11175 910
rect 11195 890 11205 910
rect 11165 880 11205 890
rect 11260 910 11300 920
rect 11260 890 11270 910
rect 11290 890 11300 910
rect 11260 880 11300 890
rect 11370 910 11410 920
rect 11370 890 11380 910
rect 11400 890 11410 910
rect 11370 880 11410 890
rect 11480 910 11520 920
rect 11480 890 11490 910
rect 11510 890 11520 910
rect 11480 880 11520 890
rect 11590 910 11630 920
rect 11590 890 11600 910
rect 11620 890 11630 910
rect 11590 880 11630 890
rect 11700 910 11740 920
rect 11700 890 11710 910
rect 11730 890 11740 910
rect 11700 880 11740 890
rect 11810 910 11850 920
rect 11810 890 11820 910
rect 11840 890 11850 910
rect 11810 880 11850 890
rect 11920 910 11960 920
rect 11920 890 11930 910
rect 11950 890 11960 910
rect 11920 880 11960 890
rect 12030 910 12070 920
rect 12030 890 12040 910
rect 12060 890 12070 910
rect 12030 880 12070 890
rect 12140 910 12180 920
rect 12140 890 12150 910
rect 12170 890 12180 910
rect 12140 880 12180 890
rect 12250 910 12290 920
rect 12250 890 12260 910
rect 12280 890 12290 910
rect 12250 880 12290 890
rect 12360 910 12400 920
rect 12360 890 12370 910
rect 12390 890 12400 910
rect 12360 880 12400 890
rect 12470 910 12510 920
rect 12470 890 12480 910
rect 12500 890 12510 910
rect 12470 880 12510 890
rect 12620 910 12660 920
rect 12620 890 12630 910
rect 12650 890 12660 910
rect 12965 910 12975 930
rect 12995 910 13005 930
rect 12965 900 13005 910
rect 13205 930 13245 940
rect 13205 910 13215 930
rect 13235 910 13245 930
rect 13205 900 13245 910
rect 13405 930 13445 940
rect 13405 910 13415 930
rect 13435 910 13445 930
rect 13405 900 13445 910
rect 13645 930 13685 940
rect 13645 910 13655 930
rect 13675 910 13685 930
rect 13770 910 13795 960
rect 26170 1110 26240 1140
rect 26170 1090 26175 1110
rect 26195 1090 26215 1110
rect 26235 1090 26240 1110
rect 26170 1060 26240 1090
rect 26170 1040 26175 1060
rect 26195 1040 26215 1060
rect 26235 1040 26240 1060
rect 26170 1010 26240 1040
rect 26170 990 26175 1010
rect 26195 990 26215 1010
rect 26235 990 26240 1010
rect 26170 980 26240 990
rect 26265 1210 26295 1220
rect 26265 1190 26270 1210
rect 26290 1190 26295 1210
rect 26265 1160 26295 1190
rect 26265 1140 26270 1160
rect 26290 1140 26295 1160
rect 26265 1110 26295 1140
rect 26265 1090 26270 1110
rect 26290 1090 26295 1110
rect 26265 1060 26295 1090
rect 26265 1040 26270 1060
rect 26290 1040 26295 1060
rect 26265 1010 26295 1040
rect 26265 990 26270 1010
rect 26290 990 26295 1010
rect 26265 980 26295 990
rect 26320 1210 26350 1220
rect 26320 1190 26325 1210
rect 26345 1190 26350 1210
rect 26320 1160 26350 1190
rect 26320 1140 26325 1160
rect 26345 1140 26350 1160
rect 26320 1110 26350 1140
rect 26320 1090 26325 1110
rect 26345 1090 26350 1110
rect 26320 1060 26350 1090
rect 26320 1040 26325 1060
rect 26345 1040 26350 1060
rect 26320 1010 26350 1040
rect 26320 990 26325 1010
rect 26345 990 26350 1010
rect 26320 980 26350 990
rect 26375 1210 26405 1220
rect 26375 1190 26380 1210
rect 26400 1190 26405 1210
rect 26375 1160 26405 1190
rect 26375 1140 26380 1160
rect 26400 1140 26405 1160
rect 26375 1110 26405 1140
rect 26375 1090 26380 1110
rect 26400 1090 26405 1110
rect 26375 1060 26405 1090
rect 26375 1040 26380 1060
rect 26400 1040 26405 1060
rect 26375 1010 26405 1040
rect 26375 990 26380 1010
rect 26400 990 26405 1010
rect 26375 980 26405 990
rect 26430 1210 26460 1220
rect 26430 1190 26435 1210
rect 26455 1190 26460 1210
rect 26430 1160 26460 1190
rect 26430 1140 26435 1160
rect 26455 1140 26460 1160
rect 26430 1110 26460 1140
rect 26430 1090 26435 1110
rect 26455 1090 26460 1110
rect 26430 1060 26460 1090
rect 26430 1040 26435 1060
rect 26455 1040 26460 1060
rect 26430 1010 26460 1040
rect 26430 990 26435 1010
rect 26455 990 26460 1010
rect 26430 980 26460 990
rect 26485 1210 26515 1220
rect 26485 1190 26490 1210
rect 26510 1190 26515 1210
rect 26485 1160 26515 1190
rect 26485 1140 26490 1160
rect 26510 1140 26515 1160
rect 26485 1110 26515 1140
rect 26485 1090 26490 1110
rect 26510 1090 26515 1110
rect 26485 1060 26515 1090
rect 26485 1040 26490 1060
rect 26510 1040 26515 1060
rect 26485 1010 26515 1040
rect 26485 990 26490 1010
rect 26510 990 26515 1010
rect 26485 980 26515 990
rect 26540 1210 26570 1220
rect 26540 1190 26545 1210
rect 26565 1190 26570 1210
rect 26540 1160 26570 1190
rect 26540 1140 26545 1160
rect 26565 1140 26570 1160
rect 26540 1110 26570 1140
rect 26540 1090 26545 1110
rect 26565 1090 26570 1110
rect 26540 1060 26570 1090
rect 26540 1040 26545 1060
rect 26565 1040 26570 1060
rect 26540 1010 26570 1040
rect 26540 990 26545 1010
rect 26565 990 26570 1010
rect 26540 980 26570 990
rect 26595 1210 26625 1220
rect 26595 1190 26600 1210
rect 26620 1190 26625 1210
rect 26595 1160 26625 1190
rect 26595 1140 26600 1160
rect 26620 1140 26625 1160
rect 26595 1110 26625 1140
rect 26595 1090 26600 1110
rect 26620 1090 26625 1110
rect 26595 1060 26625 1090
rect 26595 1040 26600 1060
rect 26620 1040 26625 1060
rect 26595 1010 26625 1040
rect 26595 990 26600 1010
rect 26620 990 26625 1010
rect 26595 980 26625 990
rect 26650 1210 26680 1220
rect 26650 1190 26655 1210
rect 26675 1190 26680 1210
rect 26650 1160 26680 1190
rect 26650 1140 26655 1160
rect 26675 1140 26680 1160
rect 26650 1110 26680 1140
rect 26650 1090 26655 1110
rect 26675 1090 26680 1110
rect 26650 1060 26680 1090
rect 26650 1040 26655 1060
rect 26675 1040 26680 1060
rect 26650 1010 26680 1040
rect 26650 990 26655 1010
rect 26675 990 26680 1010
rect 26650 980 26680 990
rect 26705 1210 26735 1220
rect 26705 1190 26710 1210
rect 26730 1190 26735 1210
rect 26705 1160 26735 1190
rect 26705 1140 26710 1160
rect 26730 1140 26735 1160
rect 26705 1110 26735 1140
rect 26705 1090 26710 1110
rect 26730 1090 26735 1110
rect 26705 1060 26735 1090
rect 26705 1040 26710 1060
rect 26730 1040 26735 1060
rect 26705 1010 26735 1040
rect 26705 990 26710 1010
rect 26730 990 26735 1010
rect 26705 980 26735 990
rect 26760 1210 26790 1220
rect 26760 1190 26765 1210
rect 26785 1190 26790 1210
rect 26760 1160 26790 1190
rect 26760 1140 26765 1160
rect 26785 1140 26790 1160
rect 26760 1110 26790 1140
rect 26760 1090 26765 1110
rect 26785 1090 26790 1110
rect 26760 1060 26790 1090
rect 26760 1040 26765 1060
rect 26785 1040 26790 1060
rect 26760 1010 26790 1040
rect 26760 990 26765 1010
rect 26785 990 26790 1010
rect 26760 980 26790 990
rect 26815 1210 26845 1220
rect 26815 1190 26820 1210
rect 26840 1190 26845 1210
rect 26815 1160 26845 1190
rect 26815 1140 26820 1160
rect 26840 1140 26845 1160
rect 26815 1110 26845 1140
rect 26815 1090 26820 1110
rect 26840 1090 26845 1110
rect 26815 1060 26845 1090
rect 26815 1040 26820 1060
rect 26840 1040 26845 1060
rect 26815 1010 26845 1040
rect 26815 990 26820 1010
rect 26840 990 26845 1010
rect 26815 980 26845 990
rect 26870 1210 26900 1220
rect 26870 1190 26875 1210
rect 26895 1190 26900 1210
rect 26870 1160 26900 1190
rect 26870 1140 26875 1160
rect 26895 1140 26900 1160
rect 26870 1110 26900 1140
rect 26870 1090 26875 1110
rect 26895 1090 26900 1110
rect 26870 1060 26900 1090
rect 26870 1040 26875 1060
rect 26895 1040 26900 1060
rect 26870 1010 26900 1040
rect 26870 990 26875 1010
rect 26895 990 26900 1010
rect 26870 980 26900 990
rect 26925 1210 26955 1220
rect 26925 1190 26930 1210
rect 26950 1190 26955 1210
rect 26925 1160 26955 1190
rect 26925 1140 26930 1160
rect 26950 1140 26955 1160
rect 26925 1110 26955 1140
rect 26925 1090 26930 1110
rect 26950 1090 26955 1110
rect 26925 1060 26955 1090
rect 26925 1040 26930 1060
rect 26950 1040 26955 1060
rect 26925 1010 26955 1040
rect 26925 990 26930 1010
rect 26950 990 26955 1010
rect 26925 980 26955 990
rect 26980 1210 27010 1220
rect 26980 1190 26985 1210
rect 27005 1190 27010 1210
rect 26980 1160 27010 1190
rect 26980 1140 26985 1160
rect 27005 1140 27010 1160
rect 26980 1110 27010 1140
rect 26980 1090 26985 1110
rect 27005 1090 27010 1110
rect 26980 1060 27010 1090
rect 26980 1040 26985 1060
rect 27005 1040 27010 1060
rect 26980 1010 27010 1040
rect 26980 990 26985 1010
rect 27005 990 27010 1010
rect 26980 980 27010 990
rect 27035 1210 27065 1220
rect 27035 1190 27040 1210
rect 27060 1190 27065 1210
rect 27035 1160 27065 1190
rect 27035 1140 27040 1160
rect 27060 1140 27065 1160
rect 27035 1110 27065 1140
rect 27035 1090 27040 1110
rect 27060 1090 27065 1110
rect 27035 1060 27065 1090
rect 27035 1040 27040 1060
rect 27060 1040 27065 1060
rect 27035 1010 27065 1040
rect 27035 990 27040 1010
rect 27060 990 27065 1010
rect 27035 980 27065 990
rect 27090 1210 27120 1220
rect 27090 1190 27095 1210
rect 27115 1190 27120 1210
rect 27090 1160 27120 1190
rect 27090 1140 27095 1160
rect 27115 1140 27120 1160
rect 27090 1110 27120 1140
rect 27090 1090 27095 1110
rect 27115 1090 27120 1110
rect 27090 1060 27120 1090
rect 27090 1040 27095 1060
rect 27115 1040 27120 1060
rect 27090 1010 27120 1040
rect 27090 990 27095 1010
rect 27115 990 27120 1010
rect 27090 980 27120 990
rect 27145 1210 27175 1220
rect 27145 1190 27150 1210
rect 27170 1190 27175 1210
rect 27145 1160 27175 1190
rect 27145 1140 27150 1160
rect 27170 1140 27175 1160
rect 27145 1110 27175 1140
rect 27145 1090 27150 1110
rect 27170 1090 27175 1110
rect 27145 1060 27175 1090
rect 27145 1040 27150 1060
rect 27170 1040 27175 1060
rect 27145 1010 27175 1040
rect 27145 990 27150 1010
rect 27170 990 27175 1010
rect 27145 980 27175 990
rect 27200 1210 27230 1220
rect 27200 1190 27205 1210
rect 27225 1190 27230 1210
rect 27200 1160 27230 1190
rect 27200 1140 27205 1160
rect 27225 1140 27230 1160
rect 27200 1110 27230 1140
rect 27200 1090 27205 1110
rect 27225 1090 27230 1110
rect 27200 1060 27230 1090
rect 27200 1040 27205 1060
rect 27225 1040 27230 1060
rect 27200 1010 27230 1040
rect 27200 990 27205 1010
rect 27225 990 27230 1010
rect 27200 980 27230 990
rect 27255 1210 27285 1220
rect 27255 1190 27260 1210
rect 27280 1190 27285 1210
rect 27255 1160 27285 1190
rect 27255 1140 27260 1160
rect 27280 1140 27285 1160
rect 27255 1110 27285 1140
rect 27255 1090 27260 1110
rect 27280 1090 27285 1110
rect 27255 1060 27285 1090
rect 27255 1040 27260 1060
rect 27280 1040 27285 1060
rect 27255 1010 27285 1040
rect 27255 990 27260 1010
rect 27280 990 27285 1010
rect 27255 980 27285 990
rect 27310 1210 27340 1220
rect 27310 1190 27315 1210
rect 27335 1190 27340 1210
rect 27310 1160 27340 1190
rect 27310 1140 27315 1160
rect 27335 1140 27340 1160
rect 27310 1110 27340 1140
rect 27310 1090 27315 1110
rect 27335 1090 27340 1110
rect 27310 1060 27340 1090
rect 27310 1040 27315 1060
rect 27335 1040 27340 1060
rect 27310 1010 27340 1040
rect 27310 990 27315 1010
rect 27335 990 27340 1010
rect 27310 980 27340 990
rect 27365 1210 27395 1220
rect 27365 1190 27370 1210
rect 27390 1190 27395 1210
rect 27365 1160 27395 1190
rect 27365 1140 27370 1160
rect 27390 1140 27395 1160
rect 27365 1110 27395 1140
rect 27365 1090 27370 1110
rect 27390 1090 27395 1110
rect 27365 1060 27395 1090
rect 27365 1040 27370 1060
rect 27390 1040 27395 1060
rect 27365 1010 27395 1040
rect 27365 990 27370 1010
rect 27390 990 27395 1010
rect 27365 980 27395 990
rect 27420 1210 27450 1220
rect 27420 1190 27425 1210
rect 27445 1190 27450 1210
rect 27420 1160 27450 1190
rect 27420 1140 27425 1160
rect 27445 1140 27450 1160
rect 27420 1110 27450 1140
rect 27420 1090 27425 1110
rect 27445 1090 27450 1110
rect 27420 1060 27450 1090
rect 27420 1040 27425 1060
rect 27445 1040 27450 1060
rect 27420 1010 27450 1040
rect 27420 990 27425 1010
rect 27445 990 27450 1010
rect 27420 980 27450 990
rect 27475 1210 27505 1220
rect 27475 1190 27480 1210
rect 27500 1190 27505 1210
rect 27475 1160 27505 1190
rect 27475 1140 27480 1160
rect 27500 1140 27505 1160
rect 27475 1110 27505 1140
rect 27475 1090 27480 1110
rect 27500 1090 27505 1110
rect 27475 1060 27505 1090
rect 27475 1040 27480 1060
rect 27500 1040 27505 1060
rect 27475 1010 27505 1040
rect 27475 990 27480 1010
rect 27500 990 27505 1010
rect 27475 980 27505 990
rect 27530 1210 27560 1220
rect 27530 1190 27535 1210
rect 27555 1190 27560 1210
rect 27530 1160 27560 1190
rect 27530 1140 27535 1160
rect 27555 1140 27560 1160
rect 27530 1110 27560 1140
rect 27530 1090 27535 1110
rect 27555 1090 27560 1110
rect 27530 1060 27560 1090
rect 27530 1040 27535 1060
rect 27555 1040 27560 1060
rect 27530 1010 27560 1040
rect 27530 990 27535 1010
rect 27555 990 27560 1010
rect 27530 980 27560 990
rect 27585 1210 27655 1220
rect 27585 1190 27590 1210
rect 27610 1190 27630 1210
rect 27650 1190 27655 1210
rect 28100 1205 28110 1225
rect 28130 1205 28140 1225
rect 28100 1195 28140 1205
rect 28160 1225 28190 1235
rect 28160 1205 28165 1225
rect 28185 1205 28190 1225
rect 28160 1195 28190 1205
rect 28210 1225 28250 1235
rect 28210 1205 28220 1225
rect 28240 1205 28250 1225
rect 28210 1195 28250 1205
rect 27585 1160 27655 1190
rect 28110 1175 28130 1195
rect 28220 1175 28240 1195
rect 27585 1140 27590 1160
rect 27610 1140 27630 1160
rect 27650 1140 27655 1160
rect 27585 1110 27655 1140
rect 27585 1090 27590 1110
rect 27610 1090 27630 1110
rect 27650 1090 27655 1110
rect 27585 1060 27655 1090
rect 27585 1040 27590 1060
rect 27610 1040 27630 1060
rect 27650 1040 27655 1060
rect 27585 1010 27655 1040
rect 28010 1165 28080 1175
rect 28010 1145 28015 1165
rect 28035 1145 28055 1165
rect 28075 1145 28080 1165
rect 28010 1115 28080 1145
rect 28010 1095 28015 1115
rect 28035 1095 28055 1115
rect 28075 1095 28080 1115
rect 28010 1065 28080 1095
rect 28010 1045 28015 1065
rect 28035 1045 28055 1065
rect 28075 1045 28080 1065
rect 28010 1035 28080 1045
rect 28105 1165 28135 1175
rect 28105 1145 28110 1165
rect 28130 1145 28135 1165
rect 28105 1115 28135 1145
rect 28105 1095 28110 1115
rect 28130 1095 28135 1115
rect 28105 1065 28135 1095
rect 28105 1045 28110 1065
rect 28130 1045 28135 1065
rect 28105 1035 28135 1045
rect 28160 1165 28190 1175
rect 28160 1145 28165 1165
rect 28185 1145 28190 1165
rect 28160 1115 28190 1145
rect 28160 1095 28165 1115
rect 28185 1095 28190 1115
rect 28160 1065 28190 1095
rect 28160 1045 28165 1065
rect 28185 1045 28190 1065
rect 28160 1035 28190 1045
rect 28215 1165 28245 1175
rect 28215 1145 28220 1165
rect 28240 1145 28245 1165
rect 28215 1115 28245 1145
rect 28215 1095 28220 1115
rect 28240 1095 28245 1115
rect 28215 1065 28245 1095
rect 28215 1045 28220 1065
rect 28240 1045 28245 1065
rect 28215 1035 28245 1045
rect 28270 1165 28340 1175
rect 28270 1145 28275 1165
rect 28295 1145 28315 1165
rect 28335 1145 28340 1165
rect 28270 1115 28340 1145
rect 28270 1095 28275 1115
rect 28295 1095 28315 1115
rect 28335 1095 28340 1115
rect 28270 1065 28340 1095
rect 28270 1045 28275 1065
rect 28295 1045 28315 1065
rect 28335 1045 28340 1065
rect 28270 1035 28340 1045
rect 28015 1015 28035 1035
rect 28220 1015 28240 1035
rect 28315 1015 28335 1035
rect 27585 990 27590 1010
rect 27610 990 27630 1010
rect 27650 990 27655 1010
rect 27585 980 27655 990
rect 28005 1005 28045 1015
rect 28005 985 28015 1005
rect 28035 985 28045 1005
rect 26175 960 26195 980
rect 26270 960 26290 980
rect 26380 960 26400 980
rect 26490 960 26510 980
rect 26600 960 26620 980
rect 26710 960 26730 980
rect 26820 960 26840 980
rect 26930 960 26950 980
rect 27040 960 27060 980
rect 27150 960 27170 980
rect 27260 960 27280 980
rect 27370 960 27390 980
rect 27480 960 27500 980
rect 27630 960 27650 980
rect 28005 975 28045 985
rect 28185 1005 28240 1015
rect 28185 985 28195 1005
rect 28215 995 28240 1005
rect 28305 1005 28345 1015
rect 28215 985 28225 995
rect 28185 975 28225 985
rect 28305 985 28315 1005
rect 28335 985 28345 1005
rect 28305 975 28345 985
rect 26165 950 26205 960
rect 26165 930 26175 950
rect 26195 930 26205 950
rect 26165 920 26205 930
rect 26260 950 26300 960
rect 26260 930 26270 950
rect 26290 930 26300 950
rect 26260 920 26300 930
rect 26370 950 26410 960
rect 26370 930 26380 950
rect 26400 930 26410 950
rect 26370 920 26410 930
rect 26480 950 26520 960
rect 26480 930 26490 950
rect 26510 930 26520 950
rect 26480 920 26520 930
rect 26590 950 26630 960
rect 26590 930 26600 950
rect 26620 930 26630 950
rect 26590 920 26630 930
rect 26700 950 26740 960
rect 26700 930 26710 950
rect 26730 930 26740 950
rect 26700 920 26740 930
rect 26810 950 26850 960
rect 26810 930 26820 950
rect 26840 930 26850 950
rect 26810 920 26850 930
rect 26920 950 26960 960
rect 26920 930 26930 950
rect 26950 930 26960 950
rect 26920 920 26960 930
rect 27030 950 27070 960
rect 27030 930 27040 950
rect 27060 930 27070 950
rect 27030 920 27070 930
rect 27140 950 27180 960
rect 27140 930 27150 950
rect 27170 930 27180 950
rect 27140 920 27180 930
rect 27250 950 27290 960
rect 27250 930 27260 950
rect 27280 930 27290 950
rect 27250 920 27290 930
rect 27360 950 27400 960
rect 27360 930 27370 950
rect 27390 930 27400 950
rect 27360 920 27400 930
rect 27470 950 27510 960
rect 27470 930 27480 950
rect 27500 930 27510 950
rect 27470 920 27510 930
rect 27620 950 27660 960
rect 27620 930 27630 950
rect 27650 930 27660 950
rect 27620 920 27660 930
rect 13645 900 13685 910
rect 12620 880 12660 890
rect 2960 865 3030 875
rect 2960 845 2965 865
rect 2985 845 3005 865
rect 3025 845 3030 865
rect 2960 815 3030 845
rect 2960 795 2965 815
rect 2985 795 3005 815
rect 3025 795 3030 815
rect 2960 785 3030 795
rect 3090 865 3120 875
rect 3090 845 3095 865
rect 3115 845 3120 865
rect 3090 815 3120 845
rect 3090 795 3095 815
rect 3115 795 3120 815
rect 3090 785 3120 795
rect 3180 865 3210 875
rect 3180 845 3185 865
rect 3205 845 3210 865
rect 3180 815 3210 845
rect 3180 795 3185 815
rect 3205 795 3210 815
rect 3180 785 3210 795
rect 3270 865 3300 875
rect 3270 845 3275 865
rect 3295 845 3300 865
rect 3270 815 3300 845
rect 3270 795 3275 815
rect 3295 795 3300 815
rect 3270 785 3300 795
rect 3360 865 3390 875
rect 3360 845 3365 865
rect 3385 845 3390 865
rect 3360 815 3390 845
rect 3360 795 3365 815
rect 3385 795 3390 815
rect 3360 785 3390 795
rect 3450 865 3480 875
rect 3450 845 3455 865
rect 3475 845 3480 865
rect 3450 815 3480 845
rect 3450 795 3455 815
rect 3475 795 3480 815
rect 3450 785 3480 795
rect 3540 865 3570 875
rect 3540 845 3545 865
rect 3565 845 3570 865
rect 3540 815 3570 845
rect 3540 795 3545 815
rect 3565 795 3570 815
rect 3540 785 3570 795
rect 3630 865 3660 875
rect 3630 845 3635 865
rect 3655 845 3660 865
rect 3630 815 3660 845
rect 3630 795 3635 815
rect 3655 795 3660 815
rect 3630 785 3660 795
rect 3720 865 3750 875
rect 3720 845 3725 865
rect 3745 845 3750 865
rect 3720 815 3750 845
rect 3720 795 3725 815
rect 3745 795 3750 815
rect 3720 785 3750 795
rect 3810 865 3840 875
rect 3810 845 3815 865
rect 3835 845 3840 865
rect 3810 815 3840 845
rect 3810 795 3815 815
rect 3835 795 3840 815
rect 3810 785 3840 795
rect 3900 865 3930 875
rect 3900 845 3905 865
rect 3925 845 3930 865
rect 3900 815 3930 845
rect 3900 795 3905 815
rect 3925 795 3930 815
rect 3900 785 3930 795
rect 3990 865 4020 875
rect 3990 845 3995 865
rect 4015 845 4020 865
rect 3990 815 4020 845
rect 3990 795 3995 815
rect 4015 795 4020 815
rect 3990 785 4020 795
rect 4080 865 4110 875
rect 4080 845 4085 865
rect 4105 845 4110 865
rect 4080 815 4110 845
rect 4080 795 4085 815
rect 4105 795 4110 815
rect 4080 785 4110 795
rect 4170 865 4200 875
rect 4170 845 4175 865
rect 4195 845 4200 865
rect 4170 815 4200 845
rect 4170 795 4175 815
rect 4195 795 4200 815
rect 4170 785 4200 795
rect 4260 865 4290 875
rect 4260 845 4265 865
rect 4285 845 4290 865
rect 4260 815 4290 845
rect 4260 795 4265 815
rect 4285 795 4290 815
rect 4260 785 4290 795
rect 4350 865 4380 875
rect 4350 845 4355 865
rect 4375 845 4380 865
rect 4350 815 4380 845
rect 4350 795 4355 815
rect 4375 795 4380 815
rect 4350 785 4380 795
rect 4440 865 4470 875
rect 4440 845 4445 865
rect 4465 845 4470 865
rect 4440 815 4470 845
rect 4440 795 4445 815
rect 4465 795 4470 815
rect 4440 785 4470 795
rect 4530 865 4560 875
rect 4530 845 4535 865
rect 4555 845 4560 865
rect 4530 815 4560 845
rect 4530 795 4535 815
rect 4555 795 4560 815
rect 4530 785 4560 795
rect 4620 865 4650 875
rect 4620 845 4625 865
rect 4645 845 4650 865
rect 4620 815 4650 845
rect 4620 795 4625 815
rect 4645 795 4650 815
rect 4620 785 4650 795
rect 4710 865 4740 875
rect 4710 845 4715 865
rect 4735 845 4740 865
rect 4710 815 4740 845
rect 4710 795 4715 815
rect 4735 795 4740 815
rect 4710 785 4740 795
rect 4800 865 4830 875
rect 4800 845 4805 865
rect 4825 845 4830 865
rect 4800 815 4830 845
rect 4800 795 4805 815
rect 4825 795 4830 815
rect 4800 785 4830 795
rect 4890 865 4920 875
rect 4890 845 4895 865
rect 4915 845 4920 865
rect 4890 815 4920 845
rect 4890 795 4895 815
rect 4915 795 4920 815
rect 4890 785 4920 795
rect 4980 865 5050 875
rect 4980 845 4985 865
rect 5005 845 5025 865
rect 5045 845 5050 865
rect 4980 815 5050 845
rect 11010 825 11040 855
rect 11495 820 11535 860
rect 11940 830 11970 860
rect 12160 830 12190 860
rect 12380 830 12410 860
rect 12865 830 12895 860
rect 4980 795 4985 815
rect 5005 795 5025 815
rect 5045 795 5050 815
rect 4980 785 5050 795
rect 3095 765 3115 785
rect 3275 765 3295 785
rect 3455 765 3475 785
rect 3635 765 3655 785
rect 3815 765 3835 785
rect 3995 765 4015 785
rect 4175 765 4195 785
rect 4355 765 4375 785
rect 4535 765 4555 785
rect 4715 765 4735 785
rect 4895 765 4915 785
rect 10955 765 10985 795
rect 11305 790 11345 800
rect 11305 780 11315 790
rect 11275 770 11315 780
rect 11335 770 11345 790
rect 2525 730 2555 760
rect 3095 755 3170 765
rect 3095 745 3140 755
rect 3130 735 3140 745
rect 3160 735 3170 755
rect 3130 725 3170 735
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 755 3665 765
rect 3625 735 3635 755
rect 3655 735 3665 755
rect 3625 725 3665 735
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 755 4025 765
rect 3985 735 3995 755
rect 4015 735 4025 755
rect 3985 725 4025 735
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 755 4385 765
rect 4345 735 4355 755
rect 4375 735 4385 755
rect 4345 725 4385 735
rect 4525 755 4565 765
rect 4525 735 4535 755
rect 4555 735 4565 755
rect 4525 725 4565 735
rect 4705 755 4745 765
rect 4705 735 4715 755
rect 4735 735 4745 755
rect 4705 725 4745 735
rect 4885 755 4925 765
rect 4885 735 4895 755
rect 4915 735 4925 755
rect 11275 760 11345 770
rect 11375 790 11415 800
rect 11375 770 11385 790
rect 11405 770 11415 790
rect 11375 760 11415 770
rect 11445 790 11485 800
rect 11445 770 11455 790
rect 11475 770 11485 790
rect 11445 760 11485 770
rect 11275 740 11295 760
rect 11505 740 11525 820
rect 11935 795 11975 805
rect 11935 775 11945 795
rect 11965 775 11975 795
rect 11935 765 11975 775
rect 12045 795 12085 805
rect 12045 775 12055 795
rect 12075 775 12085 795
rect 12045 765 12085 775
rect 12155 795 12195 805
rect 12155 775 12165 795
rect 12185 775 12195 795
rect 12155 765 12195 775
rect 12265 795 12305 805
rect 12265 775 12275 795
rect 12295 775 12305 795
rect 12265 765 12305 775
rect 12375 795 12415 805
rect 12375 775 12385 795
rect 12405 775 12415 795
rect 12375 765 12415 775
rect 12485 795 12525 805
rect 12485 775 12495 795
rect 12515 775 12525 795
rect 12485 765 12525 775
rect 12810 770 12840 800
rect 11945 745 11965 765
rect 12055 745 12075 765
rect 12165 745 12185 765
rect 12275 745 12295 765
rect 12385 745 12405 765
rect 12495 745 12515 765
rect 4885 725 4925 735
rect 11265 730 11295 740
rect 11265 710 11270 730
rect 11290 710 11295 730
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 11265 680 11295 710
rect 11265 660 11270 680
rect 11290 660 11295 680
rect 11265 650 11295 660
rect 11495 730 11525 740
rect 11495 710 11500 730
rect 11520 710 11525 730
rect 11495 680 11525 710
rect 11845 735 11915 745
rect 11845 715 11850 735
rect 11870 715 11890 735
rect 11910 715 11915 735
rect 11845 705 11915 715
rect 11940 735 11970 745
rect 11940 715 11945 735
rect 11965 715 11970 735
rect 11940 705 11970 715
rect 11995 735 12025 745
rect 11995 715 12000 735
rect 12020 715 12025 735
rect 11995 705 12025 715
rect 12050 735 12080 745
rect 12050 715 12055 735
rect 12075 715 12080 735
rect 12050 705 12080 715
rect 12105 735 12135 745
rect 12105 715 12110 735
rect 12130 715 12135 735
rect 12105 705 12135 715
rect 12160 735 12190 745
rect 12160 715 12165 735
rect 12185 715 12190 735
rect 12160 705 12190 715
rect 12215 735 12245 745
rect 12215 715 12220 735
rect 12240 715 12245 735
rect 12215 705 12245 715
rect 12270 735 12300 745
rect 12270 715 12275 735
rect 12295 715 12300 735
rect 12270 705 12300 715
rect 12325 735 12355 745
rect 12325 715 12330 735
rect 12350 715 12355 735
rect 12325 705 12355 715
rect 12380 735 12410 745
rect 12380 715 12385 735
rect 12405 715 12410 735
rect 12380 705 12410 715
rect 12435 735 12465 745
rect 12435 715 12440 735
rect 12460 715 12465 735
rect 12435 705 12465 715
rect 12490 735 12520 745
rect 12490 715 12495 735
rect 12515 715 12520 735
rect 12490 705 12520 715
rect 12545 735 12615 745
rect 12545 715 12550 735
rect 12570 715 12590 735
rect 12610 715 12615 735
rect 12545 705 12615 715
rect 11850 685 11870 705
rect 12000 685 12020 705
rect 12110 685 12130 705
rect 12220 685 12240 705
rect 12330 685 12350 705
rect 12440 685 12460 705
rect 12590 685 12610 705
rect 11495 660 11500 680
rect 11520 660 11525 680
rect 11495 650 11525 660
rect 11840 675 11880 685
rect 11840 655 11850 675
rect 11870 655 11880 675
rect 11840 645 11880 655
rect 11990 675 12030 685
rect 11990 655 12000 675
rect 12020 655 12030 675
rect 11990 645 12030 655
rect 12100 675 12140 685
rect 12100 655 12110 675
rect 12130 655 12140 675
rect 12100 645 12140 655
rect 12210 675 12250 685
rect 12210 655 12220 675
rect 12240 655 12250 675
rect 12210 645 12250 655
rect 12320 675 12360 685
rect 12320 655 12330 675
rect 12350 655 12360 675
rect 12320 645 12360 655
rect 12430 675 12470 685
rect 12430 655 12440 675
rect 12460 655 12470 675
rect 12430 645 12470 655
rect 12580 675 12620 685
rect 12580 655 12590 675
rect 12610 655 12620 675
rect 12580 645 12620 655
rect 11180 -1380 11220 -1370
rect 10905 -1395 11030 -1385
rect 10905 -1415 10915 -1395
rect 10935 -1405 11030 -1395
rect 10935 -1415 10945 -1405
rect 10905 -1425 10945 -1415
rect 11010 -1425 11030 -1405
rect 11180 -1400 11190 -1380
rect 11210 -1400 11220 -1380
rect 11180 -1410 11220 -1400
rect 11340 -1380 11380 -1370
rect 11340 -1400 11350 -1380
rect 11370 -1400 11380 -1380
rect 11340 -1410 11380 -1400
rect 11460 -1380 11500 -1370
rect 11460 -1400 11470 -1380
rect 11490 -1400 11500 -1380
rect 11460 -1410 11500 -1400
rect 11580 -1380 11620 -1370
rect 11580 -1400 11590 -1380
rect 11610 -1400 11620 -1380
rect 11580 -1410 11620 -1400
rect 11700 -1380 11740 -1370
rect 11700 -1400 11710 -1380
rect 11730 -1400 11740 -1380
rect 11700 -1410 11740 -1400
rect 11820 -1380 11860 -1370
rect 11820 -1400 11830 -1380
rect 11850 -1400 11860 -1380
rect 11820 -1410 11860 -1400
rect 11940 -1380 11980 -1370
rect 11940 -1400 11950 -1380
rect 11970 -1400 11980 -1380
rect 11940 -1410 11980 -1400
rect 12060 -1380 12100 -1370
rect 12060 -1400 12070 -1380
rect 12090 -1400 12100 -1380
rect 12060 -1410 12100 -1400
rect 12180 -1380 12220 -1370
rect 12180 -1400 12190 -1380
rect 12210 -1400 12220 -1380
rect 12180 -1410 12220 -1400
rect 12300 -1380 12340 -1370
rect 12300 -1400 12310 -1380
rect 12330 -1400 12340 -1380
rect 12300 -1410 12340 -1400
rect 12420 -1380 12460 -1370
rect 12420 -1400 12430 -1380
rect 12450 -1400 12460 -1380
rect 12420 -1410 12460 -1400
rect 12580 -1380 12620 -1370
rect 12580 -1400 12590 -1380
rect 12610 -1400 12620 -1380
rect 12580 -1410 12620 -1400
rect 11005 -1435 11035 -1425
rect 11005 -1455 11010 -1435
rect 11030 -1455 11035 -1435
rect 10785 -1485 10855 -1455
rect 10785 -1505 10790 -1485
rect 10810 -1505 10830 -1485
rect 10850 -1505 10855 -1485
rect 10785 -1535 10855 -1505
rect 10785 -1555 10790 -1535
rect 10810 -1555 10830 -1535
rect 10850 -1555 10855 -1535
rect 10785 -1585 10855 -1555
rect 10785 -1605 10790 -1585
rect 10810 -1605 10830 -1585
rect 10850 -1605 10855 -1585
rect 10785 -1635 10855 -1605
rect 10450 -1660 10490 -1650
rect 10450 -1680 10460 -1660
rect 10480 -1680 10490 -1660
rect 10450 -1690 10490 -1680
rect 10710 -1660 10750 -1650
rect 10710 -1680 10720 -1660
rect 10740 -1680 10750 -1660
rect 10710 -1690 10750 -1680
rect 10785 -1655 10790 -1635
rect 10810 -1655 10830 -1635
rect 10850 -1655 10855 -1635
rect 10785 -1685 10855 -1655
rect 10460 -1712 10480 -1690
rect 10720 -1712 10740 -1690
rect 10785 -1705 10790 -1685
rect 10810 -1705 10830 -1685
rect 10850 -1705 10855 -1685
rect 10455 -1735 10525 -1712
rect 10455 -1755 10460 -1735
rect 10480 -1755 10500 -1735
rect 10520 -1755 10525 -1735
rect 10455 -1765 10525 -1755
rect 10555 -1730 10585 -1712
rect 10555 -1750 10560 -1730
rect 10580 -1750 10585 -1730
rect 10555 -1765 10585 -1750
rect 10615 -1730 10645 -1712
rect 10615 -1750 10620 -1730
rect 10640 -1750 10645 -1730
rect 10615 -1765 10645 -1750
rect 10675 -1735 10745 -1712
rect 10675 -1755 10680 -1735
rect 10700 -1755 10720 -1735
rect 10740 -1755 10745 -1735
rect 10675 -1765 10745 -1755
rect 10785 -1735 10855 -1705
rect 10785 -1755 10790 -1735
rect 10810 -1755 10830 -1735
rect 10850 -1755 10855 -1735
rect 10785 -1765 10855 -1755
rect 10885 -1485 10915 -1455
rect 10885 -1505 10890 -1485
rect 10910 -1505 10915 -1485
rect 10885 -1535 10915 -1505
rect 10885 -1555 10890 -1535
rect 10910 -1555 10915 -1535
rect 10885 -1585 10915 -1555
rect 10885 -1605 10890 -1585
rect 10910 -1605 10915 -1585
rect 10885 -1635 10915 -1605
rect 10885 -1655 10890 -1635
rect 10910 -1655 10915 -1635
rect 10885 -1685 10915 -1655
rect 10885 -1705 10890 -1685
rect 10910 -1705 10915 -1685
rect 10885 -1735 10915 -1705
rect 10885 -1755 10890 -1735
rect 10910 -1755 10915 -1735
rect 10885 -1765 10915 -1755
rect 10945 -1485 10975 -1455
rect 10945 -1505 10950 -1485
rect 10970 -1505 10975 -1485
rect 10945 -1535 10975 -1505
rect 10945 -1555 10950 -1535
rect 10970 -1555 10975 -1535
rect 10945 -1585 10975 -1555
rect 10945 -1605 10950 -1585
rect 10970 -1605 10975 -1585
rect 10945 -1635 10975 -1605
rect 10945 -1655 10950 -1635
rect 10970 -1655 10975 -1635
rect 10945 -1685 10975 -1655
rect 10945 -1705 10950 -1685
rect 10970 -1705 10975 -1685
rect 10945 -1735 10975 -1705
rect 10945 -1755 10950 -1735
rect 10970 -1755 10975 -1735
rect 10945 -1765 10975 -1755
rect 11005 -1485 11035 -1455
rect 11005 -1505 11010 -1485
rect 11030 -1505 11035 -1485
rect 11005 -1535 11035 -1505
rect 11005 -1555 11010 -1535
rect 11030 -1555 11035 -1535
rect 11005 -1585 11035 -1555
rect 11005 -1605 11010 -1585
rect 11030 -1605 11035 -1585
rect 11005 -1635 11035 -1605
rect 11005 -1655 11010 -1635
rect 11030 -1655 11035 -1635
rect 11005 -1685 11035 -1655
rect 11005 -1705 11010 -1685
rect 11030 -1705 11035 -1685
rect 11005 -1735 11035 -1705
rect 11005 -1755 11010 -1735
rect 11030 -1755 11035 -1735
rect 11005 -1765 11035 -1755
rect 11065 -1435 11135 -1425
rect 11190 -1430 11210 -1410
rect 11350 -1430 11370 -1410
rect 11470 -1430 11490 -1410
rect 11590 -1430 11610 -1410
rect 11710 -1430 11730 -1410
rect 11830 -1430 11850 -1410
rect 11950 -1430 11970 -1410
rect 12070 -1430 12090 -1410
rect 12190 -1430 12210 -1410
rect 12310 -1430 12330 -1410
rect 12430 -1430 12450 -1410
rect 12590 -1430 12610 -1410
rect 11065 -1455 11070 -1435
rect 11090 -1455 11110 -1435
rect 11130 -1455 11135 -1435
rect 11065 -1485 11135 -1455
rect 11065 -1505 11070 -1485
rect 11090 -1505 11110 -1485
rect 11130 -1505 11135 -1485
rect 11065 -1535 11135 -1505
rect 11065 -1555 11070 -1535
rect 11090 -1555 11110 -1535
rect 11130 -1555 11135 -1535
rect 11065 -1585 11135 -1555
rect 11065 -1605 11070 -1585
rect 11090 -1605 11110 -1585
rect 11130 -1605 11135 -1585
rect 11065 -1635 11135 -1605
rect 11065 -1655 11070 -1635
rect 11090 -1655 11110 -1635
rect 11130 -1655 11135 -1635
rect 11065 -1685 11135 -1655
rect 11065 -1705 11070 -1685
rect 11090 -1705 11110 -1685
rect 11130 -1705 11135 -1685
rect 11065 -1735 11135 -1705
rect 11065 -1755 11070 -1735
rect 11090 -1755 11110 -1735
rect 11130 -1755 11135 -1735
rect 11065 -1765 11135 -1755
rect 11185 -1440 11255 -1430
rect 11185 -1460 11190 -1440
rect 11210 -1460 11230 -1440
rect 11250 -1460 11255 -1440
rect 11185 -1490 11255 -1460
rect 11185 -1510 11190 -1490
rect 11210 -1510 11230 -1490
rect 11250 -1510 11255 -1490
rect 11185 -1540 11255 -1510
rect 11185 -1560 11190 -1540
rect 11210 -1560 11230 -1540
rect 11250 -1560 11255 -1540
rect 11185 -1590 11255 -1560
rect 11185 -1610 11190 -1590
rect 11210 -1610 11230 -1590
rect 11250 -1610 11255 -1590
rect 11185 -1640 11255 -1610
rect 11185 -1660 11190 -1640
rect 11210 -1660 11230 -1640
rect 11250 -1660 11255 -1640
rect 11185 -1690 11255 -1660
rect 11185 -1710 11190 -1690
rect 11210 -1710 11230 -1690
rect 11250 -1710 11255 -1690
rect 11185 -1740 11255 -1710
rect 11185 -1760 11190 -1740
rect 11210 -1760 11230 -1740
rect 11250 -1760 11255 -1740
rect 10620 -1785 10640 -1765
rect 10790 -1785 10810 -1765
rect 11110 -1785 11130 -1765
rect 10580 -1795 10640 -1785
rect 10580 -1815 10590 -1795
rect 10610 -1805 10640 -1795
rect 10780 -1795 10820 -1785
rect 10610 -1815 10620 -1805
rect 10580 -1825 10620 -1815
rect 10780 -1815 10790 -1795
rect 10810 -1815 10820 -1795
rect 10780 -1825 10820 -1815
rect 10905 -1795 10940 -1785
rect 10905 -1815 10910 -1795
rect 10930 -1815 10940 -1795
rect 10905 -1825 10940 -1815
rect 10980 -1795 11015 -1785
rect 10980 -1815 10990 -1795
rect 11010 -1815 11015 -1795
rect 10980 -1825 11015 -1815
rect 11100 -1795 11140 -1785
rect 11100 -1815 11110 -1795
rect 11130 -1815 11140 -1795
rect 11100 -1825 11140 -1815
rect 11185 -1790 11255 -1760
rect 11185 -1810 11190 -1790
rect 11210 -1810 11230 -1790
rect 11250 -1810 11255 -1790
rect 11185 -1820 11255 -1810
rect 11285 -1440 11315 -1430
rect 11285 -1460 11290 -1440
rect 11310 -1460 11315 -1440
rect 11285 -1490 11315 -1460
rect 11285 -1510 11290 -1490
rect 11310 -1510 11315 -1490
rect 11285 -1540 11315 -1510
rect 11285 -1560 11290 -1540
rect 11310 -1560 11315 -1540
rect 11285 -1590 11315 -1560
rect 11285 -1610 11290 -1590
rect 11310 -1610 11315 -1590
rect 11285 -1640 11315 -1610
rect 11285 -1660 11290 -1640
rect 11310 -1660 11315 -1640
rect 11285 -1690 11315 -1660
rect 11285 -1710 11290 -1690
rect 11310 -1710 11315 -1690
rect 11285 -1740 11315 -1710
rect 11285 -1760 11290 -1740
rect 11310 -1760 11315 -1740
rect 11285 -1790 11315 -1760
rect 11285 -1810 11290 -1790
rect 11310 -1810 11315 -1790
rect 11285 -1820 11315 -1810
rect 11345 -1440 11375 -1430
rect 11345 -1460 11350 -1440
rect 11370 -1460 11375 -1440
rect 11345 -1490 11375 -1460
rect 11345 -1510 11350 -1490
rect 11370 -1510 11375 -1490
rect 11345 -1540 11375 -1510
rect 11345 -1560 11350 -1540
rect 11370 -1560 11375 -1540
rect 11345 -1590 11375 -1560
rect 11345 -1610 11350 -1590
rect 11370 -1610 11375 -1590
rect 11345 -1640 11375 -1610
rect 11345 -1660 11350 -1640
rect 11370 -1660 11375 -1640
rect 11345 -1690 11375 -1660
rect 11345 -1710 11350 -1690
rect 11370 -1710 11375 -1690
rect 11345 -1740 11375 -1710
rect 11345 -1760 11350 -1740
rect 11370 -1760 11375 -1740
rect 11345 -1790 11375 -1760
rect 11345 -1810 11350 -1790
rect 11370 -1810 11375 -1790
rect 11345 -1820 11375 -1810
rect 11405 -1440 11435 -1430
rect 11405 -1460 11410 -1440
rect 11430 -1460 11435 -1440
rect 11405 -1490 11435 -1460
rect 11405 -1510 11410 -1490
rect 11430 -1510 11435 -1490
rect 11405 -1540 11435 -1510
rect 11405 -1560 11410 -1540
rect 11430 -1560 11435 -1540
rect 11405 -1590 11435 -1560
rect 11405 -1610 11410 -1590
rect 11430 -1610 11435 -1590
rect 11405 -1640 11435 -1610
rect 11405 -1660 11410 -1640
rect 11430 -1660 11435 -1640
rect 11405 -1690 11435 -1660
rect 11405 -1710 11410 -1690
rect 11430 -1710 11435 -1690
rect 11405 -1740 11435 -1710
rect 11405 -1760 11410 -1740
rect 11430 -1760 11435 -1740
rect 11405 -1790 11435 -1760
rect 11405 -1810 11410 -1790
rect 11430 -1810 11435 -1790
rect 11405 -1820 11435 -1810
rect 11465 -1440 11495 -1430
rect 11465 -1460 11470 -1440
rect 11490 -1460 11495 -1440
rect 11465 -1490 11495 -1460
rect 11465 -1510 11470 -1490
rect 11490 -1510 11495 -1490
rect 11465 -1540 11495 -1510
rect 11465 -1560 11470 -1540
rect 11490 -1560 11495 -1540
rect 11465 -1590 11495 -1560
rect 11465 -1610 11470 -1590
rect 11490 -1610 11495 -1590
rect 11465 -1640 11495 -1610
rect 11465 -1660 11470 -1640
rect 11490 -1660 11495 -1640
rect 11465 -1690 11495 -1660
rect 11465 -1710 11470 -1690
rect 11490 -1710 11495 -1690
rect 11465 -1740 11495 -1710
rect 11465 -1760 11470 -1740
rect 11490 -1760 11495 -1740
rect 11465 -1790 11495 -1760
rect 11465 -1810 11470 -1790
rect 11490 -1810 11495 -1790
rect 11465 -1820 11495 -1810
rect 11525 -1440 11555 -1430
rect 11525 -1460 11530 -1440
rect 11550 -1460 11555 -1440
rect 11525 -1490 11555 -1460
rect 11525 -1510 11530 -1490
rect 11550 -1510 11555 -1490
rect 11525 -1540 11555 -1510
rect 11525 -1560 11530 -1540
rect 11550 -1560 11555 -1540
rect 11525 -1590 11555 -1560
rect 11525 -1610 11530 -1590
rect 11550 -1610 11555 -1590
rect 11525 -1640 11555 -1610
rect 11525 -1660 11530 -1640
rect 11550 -1660 11555 -1640
rect 11525 -1690 11555 -1660
rect 11525 -1710 11530 -1690
rect 11550 -1710 11555 -1690
rect 11525 -1740 11555 -1710
rect 11525 -1760 11530 -1740
rect 11550 -1760 11555 -1740
rect 11525 -1790 11555 -1760
rect 11525 -1810 11530 -1790
rect 11550 -1810 11555 -1790
rect 11525 -1820 11555 -1810
rect 11585 -1440 11615 -1430
rect 11585 -1460 11590 -1440
rect 11610 -1460 11615 -1440
rect 11585 -1490 11615 -1460
rect 11585 -1510 11590 -1490
rect 11610 -1510 11615 -1490
rect 11585 -1540 11615 -1510
rect 11585 -1560 11590 -1540
rect 11610 -1560 11615 -1540
rect 11585 -1590 11615 -1560
rect 11585 -1610 11590 -1590
rect 11610 -1610 11615 -1590
rect 11585 -1640 11615 -1610
rect 11585 -1660 11590 -1640
rect 11610 -1660 11615 -1640
rect 11585 -1690 11615 -1660
rect 11585 -1710 11590 -1690
rect 11610 -1710 11615 -1690
rect 11585 -1740 11615 -1710
rect 11585 -1760 11590 -1740
rect 11610 -1760 11615 -1740
rect 11585 -1790 11615 -1760
rect 11585 -1810 11590 -1790
rect 11610 -1810 11615 -1790
rect 11585 -1820 11615 -1810
rect 11645 -1440 11675 -1430
rect 11645 -1460 11650 -1440
rect 11670 -1460 11675 -1440
rect 11645 -1490 11675 -1460
rect 11645 -1510 11650 -1490
rect 11670 -1510 11675 -1490
rect 11645 -1540 11675 -1510
rect 11645 -1560 11650 -1540
rect 11670 -1560 11675 -1540
rect 11645 -1590 11675 -1560
rect 11645 -1610 11650 -1590
rect 11670 -1610 11675 -1590
rect 11645 -1640 11675 -1610
rect 11645 -1660 11650 -1640
rect 11670 -1660 11675 -1640
rect 11645 -1690 11675 -1660
rect 11645 -1710 11650 -1690
rect 11670 -1710 11675 -1690
rect 11645 -1740 11675 -1710
rect 11645 -1760 11650 -1740
rect 11670 -1760 11675 -1740
rect 11645 -1790 11675 -1760
rect 11645 -1810 11650 -1790
rect 11670 -1810 11675 -1790
rect 11645 -1820 11675 -1810
rect 11705 -1440 11735 -1430
rect 11705 -1460 11710 -1440
rect 11730 -1460 11735 -1440
rect 11705 -1490 11735 -1460
rect 11705 -1510 11710 -1490
rect 11730 -1510 11735 -1490
rect 11705 -1540 11735 -1510
rect 11705 -1560 11710 -1540
rect 11730 -1560 11735 -1540
rect 11705 -1590 11735 -1560
rect 11705 -1610 11710 -1590
rect 11730 -1610 11735 -1590
rect 11705 -1640 11735 -1610
rect 11705 -1660 11710 -1640
rect 11730 -1660 11735 -1640
rect 11705 -1690 11735 -1660
rect 11705 -1710 11710 -1690
rect 11730 -1710 11735 -1690
rect 11705 -1740 11735 -1710
rect 11705 -1760 11710 -1740
rect 11730 -1760 11735 -1740
rect 11705 -1790 11735 -1760
rect 11705 -1810 11710 -1790
rect 11730 -1810 11735 -1790
rect 11705 -1820 11735 -1810
rect 11765 -1440 11795 -1430
rect 11765 -1460 11770 -1440
rect 11790 -1460 11795 -1440
rect 11765 -1490 11795 -1460
rect 11765 -1510 11770 -1490
rect 11790 -1510 11795 -1490
rect 11765 -1540 11795 -1510
rect 11765 -1560 11770 -1540
rect 11790 -1560 11795 -1540
rect 11765 -1590 11795 -1560
rect 11765 -1610 11770 -1590
rect 11790 -1610 11795 -1590
rect 11765 -1640 11795 -1610
rect 11765 -1660 11770 -1640
rect 11790 -1660 11795 -1640
rect 11765 -1690 11795 -1660
rect 11765 -1710 11770 -1690
rect 11790 -1710 11795 -1690
rect 11765 -1740 11795 -1710
rect 11765 -1760 11770 -1740
rect 11790 -1760 11795 -1740
rect 11765 -1790 11795 -1760
rect 11765 -1810 11770 -1790
rect 11790 -1810 11795 -1790
rect 11765 -1820 11795 -1810
rect 11825 -1440 11855 -1430
rect 11825 -1460 11830 -1440
rect 11850 -1460 11855 -1440
rect 11825 -1490 11855 -1460
rect 11825 -1510 11830 -1490
rect 11850 -1510 11855 -1490
rect 11825 -1540 11855 -1510
rect 11825 -1560 11830 -1540
rect 11850 -1560 11855 -1540
rect 11825 -1590 11855 -1560
rect 11825 -1610 11830 -1590
rect 11850 -1610 11855 -1590
rect 11825 -1640 11855 -1610
rect 11825 -1660 11830 -1640
rect 11850 -1660 11855 -1640
rect 11825 -1690 11855 -1660
rect 11825 -1710 11830 -1690
rect 11850 -1710 11855 -1690
rect 11825 -1740 11855 -1710
rect 11825 -1760 11830 -1740
rect 11850 -1760 11855 -1740
rect 11825 -1790 11855 -1760
rect 11825 -1810 11830 -1790
rect 11850 -1810 11855 -1790
rect 11825 -1820 11855 -1810
rect 11885 -1440 11915 -1430
rect 11885 -1460 11890 -1440
rect 11910 -1460 11915 -1440
rect 11885 -1490 11915 -1460
rect 11885 -1510 11890 -1490
rect 11910 -1510 11915 -1490
rect 11885 -1540 11915 -1510
rect 11885 -1560 11890 -1540
rect 11910 -1560 11915 -1540
rect 11885 -1590 11915 -1560
rect 11885 -1610 11890 -1590
rect 11910 -1610 11915 -1590
rect 11885 -1640 11915 -1610
rect 11885 -1660 11890 -1640
rect 11910 -1660 11915 -1640
rect 11885 -1690 11915 -1660
rect 11885 -1710 11890 -1690
rect 11910 -1710 11915 -1690
rect 11885 -1740 11915 -1710
rect 11885 -1760 11890 -1740
rect 11910 -1760 11915 -1740
rect 11885 -1790 11915 -1760
rect 11885 -1810 11890 -1790
rect 11910 -1810 11915 -1790
rect 11885 -1820 11915 -1810
rect 11945 -1440 11975 -1430
rect 11945 -1460 11950 -1440
rect 11970 -1460 11975 -1440
rect 11945 -1490 11975 -1460
rect 11945 -1510 11950 -1490
rect 11970 -1510 11975 -1490
rect 11945 -1540 11975 -1510
rect 11945 -1560 11950 -1540
rect 11970 -1560 11975 -1540
rect 11945 -1590 11975 -1560
rect 11945 -1610 11950 -1590
rect 11970 -1610 11975 -1590
rect 11945 -1640 11975 -1610
rect 11945 -1660 11950 -1640
rect 11970 -1660 11975 -1640
rect 11945 -1690 11975 -1660
rect 11945 -1710 11950 -1690
rect 11970 -1710 11975 -1690
rect 11945 -1740 11975 -1710
rect 11945 -1760 11950 -1740
rect 11970 -1760 11975 -1740
rect 11945 -1790 11975 -1760
rect 11945 -1810 11950 -1790
rect 11970 -1810 11975 -1790
rect 11945 -1820 11975 -1810
rect 12005 -1440 12035 -1430
rect 12005 -1460 12010 -1440
rect 12030 -1460 12035 -1440
rect 12005 -1490 12035 -1460
rect 12005 -1510 12010 -1490
rect 12030 -1510 12035 -1490
rect 12005 -1540 12035 -1510
rect 12005 -1560 12010 -1540
rect 12030 -1560 12035 -1540
rect 12005 -1590 12035 -1560
rect 12005 -1610 12010 -1590
rect 12030 -1610 12035 -1590
rect 12005 -1640 12035 -1610
rect 12005 -1660 12010 -1640
rect 12030 -1660 12035 -1640
rect 12005 -1690 12035 -1660
rect 12005 -1710 12010 -1690
rect 12030 -1710 12035 -1690
rect 12005 -1740 12035 -1710
rect 12005 -1760 12010 -1740
rect 12030 -1760 12035 -1740
rect 12005 -1790 12035 -1760
rect 12005 -1810 12010 -1790
rect 12030 -1810 12035 -1790
rect 12005 -1820 12035 -1810
rect 12065 -1440 12095 -1430
rect 12065 -1460 12070 -1440
rect 12090 -1460 12095 -1440
rect 12065 -1490 12095 -1460
rect 12065 -1510 12070 -1490
rect 12090 -1510 12095 -1490
rect 12065 -1540 12095 -1510
rect 12065 -1560 12070 -1540
rect 12090 -1560 12095 -1540
rect 12065 -1590 12095 -1560
rect 12065 -1610 12070 -1590
rect 12090 -1610 12095 -1590
rect 12065 -1640 12095 -1610
rect 12065 -1660 12070 -1640
rect 12090 -1660 12095 -1640
rect 12065 -1690 12095 -1660
rect 12065 -1710 12070 -1690
rect 12090 -1710 12095 -1690
rect 12065 -1740 12095 -1710
rect 12065 -1760 12070 -1740
rect 12090 -1760 12095 -1740
rect 12065 -1790 12095 -1760
rect 12065 -1810 12070 -1790
rect 12090 -1810 12095 -1790
rect 12065 -1820 12095 -1810
rect 12125 -1440 12155 -1430
rect 12125 -1460 12130 -1440
rect 12150 -1460 12155 -1440
rect 12125 -1490 12155 -1460
rect 12125 -1510 12130 -1490
rect 12150 -1510 12155 -1490
rect 12125 -1540 12155 -1510
rect 12125 -1560 12130 -1540
rect 12150 -1560 12155 -1540
rect 12125 -1590 12155 -1560
rect 12125 -1610 12130 -1590
rect 12150 -1610 12155 -1590
rect 12125 -1640 12155 -1610
rect 12125 -1660 12130 -1640
rect 12150 -1660 12155 -1640
rect 12125 -1690 12155 -1660
rect 12125 -1710 12130 -1690
rect 12150 -1710 12155 -1690
rect 12125 -1740 12155 -1710
rect 12125 -1760 12130 -1740
rect 12150 -1760 12155 -1740
rect 12125 -1790 12155 -1760
rect 12125 -1810 12130 -1790
rect 12150 -1810 12155 -1790
rect 12125 -1820 12155 -1810
rect 12185 -1440 12215 -1430
rect 12185 -1460 12190 -1440
rect 12210 -1460 12215 -1440
rect 12185 -1490 12215 -1460
rect 12185 -1510 12190 -1490
rect 12210 -1510 12215 -1490
rect 12185 -1540 12215 -1510
rect 12185 -1560 12190 -1540
rect 12210 -1560 12215 -1540
rect 12185 -1590 12215 -1560
rect 12185 -1610 12190 -1590
rect 12210 -1610 12215 -1590
rect 12185 -1640 12215 -1610
rect 12185 -1660 12190 -1640
rect 12210 -1660 12215 -1640
rect 12185 -1690 12215 -1660
rect 12185 -1710 12190 -1690
rect 12210 -1710 12215 -1690
rect 12185 -1740 12215 -1710
rect 12185 -1760 12190 -1740
rect 12210 -1760 12215 -1740
rect 12185 -1790 12215 -1760
rect 12185 -1810 12190 -1790
rect 12210 -1810 12215 -1790
rect 12185 -1820 12215 -1810
rect 12245 -1440 12275 -1430
rect 12245 -1460 12250 -1440
rect 12270 -1460 12275 -1440
rect 12245 -1490 12275 -1460
rect 12245 -1510 12250 -1490
rect 12270 -1510 12275 -1490
rect 12245 -1540 12275 -1510
rect 12245 -1560 12250 -1540
rect 12270 -1560 12275 -1540
rect 12245 -1590 12275 -1560
rect 12245 -1610 12250 -1590
rect 12270 -1610 12275 -1590
rect 12245 -1640 12275 -1610
rect 12245 -1660 12250 -1640
rect 12270 -1660 12275 -1640
rect 12245 -1690 12275 -1660
rect 12245 -1710 12250 -1690
rect 12270 -1710 12275 -1690
rect 12245 -1740 12275 -1710
rect 12245 -1760 12250 -1740
rect 12270 -1760 12275 -1740
rect 12245 -1790 12275 -1760
rect 12245 -1810 12250 -1790
rect 12270 -1810 12275 -1790
rect 12245 -1820 12275 -1810
rect 12305 -1440 12335 -1430
rect 12305 -1460 12310 -1440
rect 12330 -1460 12335 -1440
rect 12305 -1490 12335 -1460
rect 12305 -1510 12310 -1490
rect 12330 -1510 12335 -1490
rect 12305 -1540 12335 -1510
rect 12305 -1560 12310 -1540
rect 12330 -1560 12335 -1540
rect 12305 -1590 12335 -1560
rect 12305 -1610 12310 -1590
rect 12330 -1610 12335 -1590
rect 12305 -1640 12335 -1610
rect 12305 -1660 12310 -1640
rect 12330 -1660 12335 -1640
rect 12305 -1690 12335 -1660
rect 12305 -1710 12310 -1690
rect 12330 -1710 12335 -1690
rect 12305 -1740 12335 -1710
rect 12305 -1760 12310 -1740
rect 12330 -1760 12335 -1740
rect 12305 -1790 12335 -1760
rect 12305 -1810 12310 -1790
rect 12330 -1810 12335 -1790
rect 12305 -1820 12335 -1810
rect 12365 -1440 12395 -1430
rect 12365 -1460 12370 -1440
rect 12390 -1460 12395 -1440
rect 12365 -1490 12395 -1460
rect 12365 -1510 12370 -1490
rect 12390 -1510 12395 -1490
rect 12365 -1540 12395 -1510
rect 12365 -1560 12370 -1540
rect 12390 -1560 12395 -1540
rect 12365 -1590 12395 -1560
rect 12365 -1610 12370 -1590
rect 12390 -1610 12395 -1590
rect 12365 -1640 12395 -1610
rect 12365 -1660 12370 -1640
rect 12390 -1660 12395 -1640
rect 12365 -1690 12395 -1660
rect 12365 -1710 12370 -1690
rect 12390 -1710 12395 -1690
rect 12365 -1740 12395 -1710
rect 12365 -1760 12370 -1740
rect 12390 -1760 12395 -1740
rect 12365 -1790 12395 -1760
rect 12365 -1810 12370 -1790
rect 12390 -1810 12395 -1790
rect 12365 -1820 12395 -1810
rect 12425 -1440 12455 -1430
rect 12425 -1460 12430 -1440
rect 12450 -1460 12455 -1440
rect 12425 -1490 12455 -1460
rect 12425 -1510 12430 -1490
rect 12450 -1510 12455 -1490
rect 12425 -1540 12455 -1510
rect 12425 -1560 12430 -1540
rect 12450 -1560 12455 -1540
rect 12425 -1590 12455 -1560
rect 12425 -1610 12430 -1590
rect 12450 -1610 12455 -1590
rect 12425 -1640 12455 -1610
rect 12425 -1660 12430 -1640
rect 12450 -1660 12455 -1640
rect 12425 -1690 12455 -1660
rect 12425 -1710 12430 -1690
rect 12450 -1710 12455 -1690
rect 12425 -1740 12455 -1710
rect 12425 -1760 12430 -1740
rect 12450 -1760 12455 -1740
rect 12425 -1790 12455 -1760
rect 12425 -1810 12430 -1790
rect 12450 -1810 12455 -1790
rect 12425 -1820 12455 -1810
rect 12485 -1440 12515 -1430
rect 12485 -1460 12490 -1440
rect 12510 -1460 12515 -1440
rect 12485 -1490 12515 -1460
rect 12485 -1510 12490 -1490
rect 12510 -1510 12515 -1490
rect 12485 -1540 12515 -1510
rect 12485 -1560 12490 -1540
rect 12510 -1560 12515 -1540
rect 12485 -1590 12515 -1560
rect 12485 -1610 12490 -1590
rect 12510 -1610 12515 -1590
rect 12485 -1640 12515 -1610
rect 12485 -1660 12490 -1640
rect 12510 -1660 12515 -1640
rect 12485 -1690 12515 -1660
rect 12485 -1710 12490 -1690
rect 12510 -1710 12515 -1690
rect 12485 -1740 12515 -1710
rect 12485 -1760 12490 -1740
rect 12510 -1760 12515 -1740
rect 12485 -1790 12515 -1760
rect 12485 -1810 12490 -1790
rect 12510 -1810 12515 -1790
rect 12485 -1820 12515 -1810
rect 12545 -1440 12615 -1430
rect 12545 -1460 12550 -1440
rect 12570 -1460 12590 -1440
rect 12610 -1460 12615 -1440
rect 12545 -1490 12615 -1460
rect 12545 -1510 12550 -1490
rect 12570 -1510 12590 -1490
rect 12610 -1510 12615 -1490
rect 12545 -1540 12615 -1510
rect 12545 -1560 12550 -1540
rect 12570 -1560 12590 -1540
rect 12610 -1560 12615 -1540
rect 12545 -1590 12615 -1560
rect 12545 -1610 12550 -1590
rect 12570 -1610 12590 -1590
rect 12610 -1610 12615 -1590
rect 12545 -1640 12615 -1610
rect 12545 -1660 12550 -1640
rect 12570 -1660 12590 -1640
rect 12610 -1660 12615 -1640
rect 12545 -1690 12615 -1660
rect 12545 -1710 12550 -1690
rect 12570 -1710 12590 -1690
rect 12610 -1710 12615 -1690
rect 12545 -1740 12615 -1710
rect 12545 -1760 12550 -1740
rect 12570 -1760 12590 -1740
rect 12610 -1760 12615 -1740
rect 12545 -1790 12615 -1760
rect 12545 -1810 12550 -1790
rect 12570 -1810 12590 -1790
rect 12610 -1810 12615 -1790
rect 12545 -1820 12615 -1810
rect 11290 -1840 11310 -1820
rect 11410 -1840 11430 -1820
rect 11530 -1840 11550 -1820
rect 11650 -1840 11670 -1820
rect 11770 -1840 11790 -1820
rect 11890 -1840 11910 -1820
rect 12010 -1840 12030 -1820
rect 12130 -1840 12150 -1820
rect 12250 -1840 12270 -1820
rect 12370 -1840 12390 -1820
rect 12490 -1840 12510 -1820
rect 11280 -1850 11320 -1840
rect 11280 -1870 11290 -1850
rect 11310 -1870 11320 -1850
rect 11280 -1880 11320 -1870
rect 11400 -1850 11440 -1840
rect 11400 -1870 11410 -1850
rect 11430 -1870 11440 -1850
rect 11400 -1880 11440 -1870
rect 11520 -1850 11560 -1840
rect 11520 -1870 11530 -1850
rect 11550 -1870 11560 -1850
rect 11520 -1880 11560 -1870
rect 11640 -1850 11680 -1840
rect 11640 -1870 11650 -1850
rect 11670 -1870 11680 -1850
rect 11640 -1880 11680 -1870
rect 11760 -1850 11800 -1840
rect 11760 -1870 11770 -1850
rect 11790 -1870 11800 -1850
rect 11760 -1880 11800 -1870
rect 11823 -1850 11857 -1840
rect 11823 -1870 11831 -1850
rect 11849 -1870 11857 -1850
rect 11823 -1880 11857 -1870
rect 11880 -1850 11920 -1840
rect 11880 -1870 11890 -1850
rect 11910 -1870 11920 -1850
rect 11880 -1880 11920 -1870
rect 12000 -1850 12040 -1840
rect 12000 -1870 12010 -1850
rect 12030 -1870 12040 -1850
rect 12000 -1880 12040 -1870
rect 12120 -1850 12160 -1840
rect 12120 -1870 12130 -1850
rect 12150 -1870 12160 -1850
rect 12120 -1880 12160 -1870
rect 12240 -1850 12280 -1840
rect 12240 -1870 12250 -1850
rect 12270 -1870 12280 -1850
rect 12240 -1880 12280 -1870
rect 12360 -1850 12400 -1840
rect 12360 -1870 12370 -1850
rect 12390 -1870 12400 -1850
rect 12360 -1880 12400 -1870
rect 12480 -1850 12520 -1840
rect 12480 -1870 12490 -1850
rect 12510 -1870 12520 -1850
rect 12480 -1880 12520 -1870
rect 12950 -1970 12990 -1960
rect 12950 -1990 12960 -1970
rect 12980 -1990 12990 -1970
rect 12950 -2000 12990 -1990
rect 13060 -1970 13100 -1960
rect 13060 -1990 13070 -1970
rect 13090 -1990 13100 -1970
rect 13060 -2000 13100 -1990
rect 13170 -1970 13210 -1960
rect 13170 -1990 13180 -1970
rect 13200 -1990 13210 -1970
rect 13170 -2000 13210 -1990
rect 13280 -1970 13320 -1960
rect 13280 -1990 13290 -1970
rect 13310 -1990 13320 -1970
rect 13280 -2000 13320 -1990
rect 13390 -1970 13430 -1960
rect 13390 -1990 13400 -1970
rect 13420 -1990 13430 -1970
rect 13390 -2000 13430 -1990
rect 13500 -1970 13540 -1960
rect 13500 -1990 13510 -1970
rect 13530 -1990 13540 -1970
rect 13500 -2000 13540 -1990
rect 13610 -1970 13650 -1960
rect 13610 -1990 13620 -1970
rect 13640 -1990 13650 -1970
rect 13610 -2000 13650 -1990
rect 13720 -1970 13760 -1960
rect 13720 -1990 13730 -1970
rect 13750 -1990 13760 -1970
rect 13720 -2000 13760 -1990
rect 13830 -1970 13870 -1960
rect 13830 -1990 13840 -1970
rect 13860 -1990 13870 -1970
rect 13830 -2000 13870 -1990
rect 13940 -1970 13980 -1960
rect 13940 -1990 13950 -1970
rect 13970 -1990 13980 -1970
rect 13940 -2000 13980 -1990
rect 14050 -1970 14090 -1960
rect 14050 -1990 14060 -1970
rect 14080 -1990 14090 -1970
rect 14050 -2000 14090 -1990
rect 12960 -2020 12980 -2000
rect 13070 -2020 13090 -2000
rect 13180 -2020 13200 -2000
rect 13290 -2020 13310 -2000
rect 13400 -2020 13420 -2000
rect 13510 -2020 13530 -2000
rect 13620 -2020 13640 -2000
rect 13730 -2020 13750 -2000
rect 13840 -2020 13860 -2000
rect 13950 -2020 13970 -2000
rect 14060 -2020 14080 -2000
rect 12860 -2030 12930 -2020
rect 12860 -2050 12865 -2030
rect 12885 -2050 12905 -2030
rect 12925 -2050 12930 -2030
rect 11180 -2060 11220 -2050
rect 11180 -2080 11190 -2060
rect 11210 -2080 11220 -2060
rect 11180 -2090 11220 -2080
rect 11340 -2060 11380 -2050
rect 11340 -2080 11350 -2060
rect 11370 -2080 11380 -2060
rect 11340 -2090 11380 -2080
rect 11460 -2060 11500 -2050
rect 11460 -2080 11470 -2060
rect 11490 -2080 11500 -2060
rect 11460 -2090 11500 -2080
rect 11580 -2060 11620 -2050
rect 11580 -2080 11590 -2060
rect 11610 -2080 11620 -2060
rect 11580 -2090 11620 -2080
rect 11700 -2060 11740 -2050
rect 11700 -2080 11710 -2060
rect 11730 -2080 11740 -2060
rect 11700 -2090 11740 -2080
rect 11820 -2060 11860 -2050
rect 11820 -2080 11830 -2060
rect 11850 -2080 11860 -2060
rect 11820 -2090 11860 -2080
rect 11940 -2060 11980 -2050
rect 11940 -2080 11950 -2060
rect 11970 -2080 11980 -2060
rect 11940 -2090 11980 -2080
rect 12060 -2060 12100 -2050
rect 12060 -2080 12070 -2060
rect 12090 -2080 12100 -2060
rect 12060 -2090 12100 -2080
rect 12180 -2060 12220 -2050
rect 12180 -2080 12190 -2060
rect 12210 -2080 12220 -2060
rect 12180 -2090 12220 -2080
rect 12300 -2060 12340 -2050
rect 12300 -2080 12310 -2060
rect 12330 -2080 12340 -2060
rect 12300 -2090 12340 -2080
rect 12420 -2060 12460 -2050
rect 12420 -2080 12430 -2060
rect 12450 -2080 12460 -2060
rect 12420 -2090 12460 -2080
rect 12480 -2090 12520 -2050
rect 12580 -2060 12620 -2050
rect 12580 -2080 12590 -2060
rect 12610 -2080 12620 -2060
rect 12580 -2090 12620 -2080
rect 12860 -2080 12930 -2050
rect 11190 -2110 11210 -2090
rect 11350 -2110 11370 -2090
rect 11470 -2110 11490 -2090
rect 11590 -2110 11610 -2090
rect 11710 -2110 11730 -2090
rect 11830 -2110 11850 -2090
rect 11950 -2110 11970 -2090
rect 12070 -2110 12090 -2090
rect 12190 -2110 12210 -2090
rect 12310 -2110 12330 -2090
rect 12430 -2110 12450 -2090
rect 12590 -2110 12610 -2090
rect 12860 -2100 12865 -2080
rect 12885 -2100 12905 -2080
rect 12925 -2100 12930 -2080
rect 11185 -2120 11255 -2110
rect 11185 -2140 11190 -2120
rect 11210 -2140 11230 -2120
rect 11250 -2140 11255 -2120
rect 11185 -2170 11255 -2140
rect 11185 -2190 11190 -2170
rect 11210 -2190 11230 -2170
rect 11250 -2190 11255 -2170
rect 11185 -2220 11255 -2190
rect 11185 -2240 11190 -2220
rect 11210 -2240 11230 -2220
rect 11250 -2240 11255 -2220
rect 11185 -2270 11255 -2240
rect 11185 -2290 11190 -2270
rect 11210 -2290 11230 -2270
rect 11250 -2290 11255 -2270
rect 11185 -2320 11255 -2290
rect 11185 -2340 11190 -2320
rect 11210 -2340 11230 -2320
rect 11250 -2340 11255 -2320
rect 11185 -2370 11255 -2340
rect 11185 -2390 11190 -2370
rect 11210 -2390 11230 -2370
rect 11250 -2390 11255 -2370
rect 11185 -2420 11255 -2390
rect 11185 -2440 11190 -2420
rect 11210 -2440 11230 -2420
rect 11250 -2440 11255 -2420
rect 11185 -2470 11255 -2440
rect 11185 -2490 11190 -2470
rect 11210 -2490 11230 -2470
rect 11250 -2490 11255 -2470
rect 11185 -2500 11255 -2490
rect 11285 -2120 11315 -2110
rect 11285 -2140 11290 -2120
rect 11310 -2140 11315 -2120
rect 11285 -2170 11315 -2140
rect 11285 -2190 11290 -2170
rect 11310 -2190 11315 -2170
rect 11285 -2220 11315 -2190
rect 11285 -2240 11290 -2220
rect 11310 -2240 11315 -2220
rect 11285 -2270 11315 -2240
rect 11285 -2290 11290 -2270
rect 11310 -2290 11315 -2270
rect 11285 -2320 11315 -2290
rect 11285 -2340 11290 -2320
rect 11310 -2340 11315 -2320
rect 11285 -2370 11315 -2340
rect 11285 -2390 11290 -2370
rect 11310 -2390 11315 -2370
rect 11285 -2420 11315 -2390
rect 11285 -2440 11290 -2420
rect 11310 -2440 11315 -2420
rect 11285 -2470 11315 -2440
rect 11285 -2490 11290 -2470
rect 11310 -2490 11315 -2470
rect 11285 -2500 11315 -2490
rect 11345 -2120 11375 -2110
rect 11345 -2140 11350 -2120
rect 11370 -2140 11375 -2120
rect 11345 -2170 11375 -2140
rect 11345 -2190 11350 -2170
rect 11370 -2190 11375 -2170
rect 11345 -2220 11375 -2190
rect 11345 -2240 11350 -2220
rect 11370 -2240 11375 -2220
rect 11345 -2270 11375 -2240
rect 11345 -2290 11350 -2270
rect 11370 -2290 11375 -2270
rect 11345 -2320 11375 -2290
rect 11345 -2340 11350 -2320
rect 11370 -2340 11375 -2320
rect 11345 -2370 11375 -2340
rect 11345 -2390 11350 -2370
rect 11370 -2390 11375 -2370
rect 11345 -2420 11375 -2390
rect 11345 -2440 11350 -2420
rect 11370 -2440 11375 -2420
rect 11345 -2470 11375 -2440
rect 11345 -2490 11350 -2470
rect 11370 -2490 11375 -2470
rect 11345 -2500 11375 -2490
rect 11405 -2120 11435 -2110
rect 11405 -2140 11410 -2120
rect 11430 -2140 11435 -2120
rect 11405 -2170 11435 -2140
rect 11405 -2190 11410 -2170
rect 11430 -2190 11435 -2170
rect 11405 -2220 11435 -2190
rect 11405 -2240 11410 -2220
rect 11430 -2240 11435 -2220
rect 11405 -2270 11435 -2240
rect 11405 -2290 11410 -2270
rect 11430 -2290 11435 -2270
rect 11405 -2320 11435 -2290
rect 11405 -2340 11410 -2320
rect 11430 -2340 11435 -2320
rect 11405 -2370 11435 -2340
rect 11405 -2390 11410 -2370
rect 11430 -2390 11435 -2370
rect 11405 -2420 11435 -2390
rect 11405 -2440 11410 -2420
rect 11430 -2440 11435 -2420
rect 11405 -2470 11435 -2440
rect 11405 -2490 11410 -2470
rect 11430 -2490 11435 -2470
rect 11405 -2500 11435 -2490
rect 11465 -2120 11495 -2110
rect 11465 -2140 11470 -2120
rect 11490 -2140 11495 -2120
rect 11465 -2170 11495 -2140
rect 11465 -2190 11470 -2170
rect 11490 -2190 11495 -2170
rect 11465 -2220 11495 -2190
rect 11465 -2240 11470 -2220
rect 11490 -2240 11495 -2220
rect 11465 -2270 11495 -2240
rect 11465 -2290 11470 -2270
rect 11490 -2290 11495 -2270
rect 11465 -2320 11495 -2290
rect 11465 -2340 11470 -2320
rect 11490 -2340 11495 -2320
rect 11465 -2370 11495 -2340
rect 11465 -2390 11470 -2370
rect 11490 -2390 11495 -2370
rect 11465 -2420 11495 -2390
rect 11465 -2440 11470 -2420
rect 11490 -2440 11495 -2420
rect 11465 -2470 11495 -2440
rect 11465 -2490 11470 -2470
rect 11490 -2490 11495 -2470
rect 11465 -2500 11495 -2490
rect 11525 -2120 11555 -2110
rect 11525 -2140 11530 -2120
rect 11550 -2140 11555 -2120
rect 11525 -2170 11555 -2140
rect 11525 -2190 11530 -2170
rect 11550 -2190 11555 -2170
rect 11525 -2220 11555 -2190
rect 11525 -2240 11530 -2220
rect 11550 -2240 11555 -2220
rect 11525 -2270 11555 -2240
rect 11525 -2290 11530 -2270
rect 11550 -2290 11555 -2270
rect 11525 -2320 11555 -2290
rect 11525 -2340 11530 -2320
rect 11550 -2340 11555 -2320
rect 11525 -2370 11555 -2340
rect 11525 -2390 11530 -2370
rect 11550 -2390 11555 -2370
rect 11525 -2420 11555 -2390
rect 11525 -2440 11530 -2420
rect 11550 -2440 11555 -2420
rect 11525 -2470 11555 -2440
rect 11525 -2490 11530 -2470
rect 11550 -2490 11555 -2470
rect 11525 -2500 11555 -2490
rect 11585 -2120 11615 -2110
rect 11585 -2140 11590 -2120
rect 11610 -2140 11615 -2120
rect 11585 -2170 11615 -2140
rect 11585 -2190 11590 -2170
rect 11610 -2190 11615 -2170
rect 11585 -2220 11615 -2190
rect 11585 -2240 11590 -2220
rect 11610 -2240 11615 -2220
rect 11585 -2270 11615 -2240
rect 11585 -2290 11590 -2270
rect 11610 -2290 11615 -2270
rect 11585 -2320 11615 -2290
rect 11585 -2340 11590 -2320
rect 11610 -2340 11615 -2320
rect 11585 -2370 11615 -2340
rect 11585 -2390 11590 -2370
rect 11610 -2390 11615 -2370
rect 11585 -2420 11615 -2390
rect 11585 -2440 11590 -2420
rect 11610 -2440 11615 -2420
rect 11585 -2470 11615 -2440
rect 11585 -2490 11590 -2470
rect 11610 -2490 11615 -2470
rect 11585 -2500 11615 -2490
rect 11645 -2120 11675 -2110
rect 11645 -2140 11650 -2120
rect 11670 -2140 11675 -2120
rect 11645 -2170 11675 -2140
rect 11645 -2190 11650 -2170
rect 11670 -2190 11675 -2170
rect 11645 -2220 11675 -2190
rect 11645 -2240 11650 -2220
rect 11670 -2240 11675 -2220
rect 11645 -2270 11675 -2240
rect 11645 -2290 11650 -2270
rect 11670 -2290 11675 -2270
rect 11645 -2320 11675 -2290
rect 11645 -2340 11650 -2320
rect 11670 -2340 11675 -2320
rect 11645 -2370 11675 -2340
rect 11645 -2390 11650 -2370
rect 11670 -2390 11675 -2370
rect 11645 -2420 11675 -2390
rect 11645 -2440 11650 -2420
rect 11670 -2440 11675 -2420
rect 11645 -2470 11675 -2440
rect 11645 -2490 11650 -2470
rect 11670 -2490 11675 -2470
rect 11645 -2500 11675 -2490
rect 11705 -2120 11735 -2110
rect 11705 -2140 11710 -2120
rect 11730 -2140 11735 -2120
rect 11705 -2170 11735 -2140
rect 11705 -2190 11710 -2170
rect 11730 -2190 11735 -2170
rect 11705 -2220 11735 -2190
rect 11705 -2240 11710 -2220
rect 11730 -2240 11735 -2220
rect 11705 -2270 11735 -2240
rect 11705 -2290 11710 -2270
rect 11730 -2290 11735 -2270
rect 11705 -2320 11735 -2290
rect 11705 -2340 11710 -2320
rect 11730 -2340 11735 -2320
rect 11705 -2370 11735 -2340
rect 11705 -2390 11710 -2370
rect 11730 -2390 11735 -2370
rect 11705 -2420 11735 -2390
rect 11705 -2440 11710 -2420
rect 11730 -2440 11735 -2420
rect 11705 -2470 11735 -2440
rect 11705 -2490 11710 -2470
rect 11730 -2490 11735 -2470
rect 11705 -2500 11735 -2490
rect 11765 -2120 11795 -2110
rect 11765 -2140 11770 -2120
rect 11790 -2140 11795 -2120
rect 11765 -2170 11795 -2140
rect 11765 -2190 11770 -2170
rect 11790 -2190 11795 -2170
rect 11765 -2220 11795 -2190
rect 11765 -2240 11770 -2220
rect 11790 -2240 11795 -2220
rect 11765 -2270 11795 -2240
rect 11765 -2290 11770 -2270
rect 11790 -2290 11795 -2270
rect 11765 -2320 11795 -2290
rect 11765 -2340 11770 -2320
rect 11790 -2340 11795 -2320
rect 11765 -2370 11795 -2340
rect 11765 -2390 11770 -2370
rect 11790 -2390 11795 -2370
rect 11765 -2420 11795 -2390
rect 11765 -2440 11770 -2420
rect 11790 -2440 11795 -2420
rect 11765 -2470 11795 -2440
rect 11765 -2490 11770 -2470
rect 11790 -2490 11795 -2470
rect 11765 -2500 11795 -2490
rect 11825 -2120 11855 -2110
rect 11825 -2140 11830 -2120
rect 11850 -2140 11855 -2120
rect 11825 -2170 11855 -2140
rect 11825 -2190 11830 -2170
rect 11850 -2190 11855 -2170
rect 11825 -2220 11855 -2190
rect 11825 -2240 11830 -2220
rect 11850 -2240 11855 -2220
rect 11825 -2270 11855 -2240
rect 11825 -2290 11830 -2270
rect 11850 -2290 11855 -2270
rect 11825 -2320 11855 -2290
rect 11825 -2340 11830 -2320
rect 11850 -2340 11855 -2320
rect 11825 -2370 11855 -2340
rect 11825 -2390 11830 -2370
rect 11850 -2390 11855 -2370
rect 11825 -2420 11855 -2390
rect 11825 -2440 11830 -2420
rect 11850 -2440 11855 -2420
rect 11825 -2470 11855 -2440
rect 11825 -2490 11830 -2470
rect 11850 -2490 11855 -2470
rect 11825 -2500 11855 -2490
rect 11885 -2120 11915 -2110
rect 11885 -2140 11890 -2120
rect 11910 -2140 11915 -2120
rect 11885 -2170 11915 -2140
rect 11885 -2190 11890 -2170
rect 11910 -2190 11915 -2170
rect 11885 -2220 11915 -2190
rect 11885 -2240 11890 -2220
rect 11910 -2240 11915 -2220
rect 11885 -2270 11915 -2240
rect 11885 -2290 11890 -2270
rect 11910 -2290 11915 -2270
rect 11885 -2320 11915 -2290
rect 11885 -2340 11890 -2320
rect 11910 -2340 11915 -2320
rect 11885 -2370 11915 -2340
rect 11885 -2390 11890 -2370
rect 11910 -2390 11915 -2370
rect 11885 -2420 11915 -2390
rect 11885 -2440 11890 -2420
rect 11910 -2440 11915 -2420
rect 11885 -2470 11915 -2440
rect 11885 -2490 11890 -2470
rect 11910 -2490 11915 -2470
rect 11885 -2500 11915 -2490
rect 11945 -2120 11975 -2110
rect 11945 -2140 11950 -2120
rect 11970 -2140 11975 -2120
rect 11945 -2170 11975 -2140
rect 11945 -2190 11950 -2170
rect 11970 -2190 11975 -2170
rect 11945 -2220 11975 -2190
rect 11945 -2240 11950 -2220
rect 11970 -2240 11975 -2220
rect 11945 -2270 11975 -2240
rect 11945 -2290 11950 -2270
rect 11970 -2290 11975 -2270
rect 11945 -2320 11975 -2290
rect 11945 -2340 11950 -2320
rect 11970 -2340 11975 -2320
rect 11945 -2370 11975 -2340
rect 11945 -2390 11950 -2370
rect 11970 -2390 11975 -2370
rect 11945 -2420 11975 -2390
rect 11945 -2440 11950 -2420
rect 11970 -2440 11975 -2420
rect 11945 -2470 11975 -2440
rect 11945 -2490 11950 -2470
rect 11970 -2490 11975 -2470
rect 11945 -2500 11975 -2490
rect 12005 -2120 12035 -2110
rect 12005 -2140 12010 -2120
rect 12030 -2140 12035 -2120
rect 12005 -2170 12035 -2140
rect 12005 -2190 12010 -2170
rect 12030 -2190 12035 -2170
rect 12005 -2220 12035 -2190
rect 12005 -2240 12010 -2220
rect 12030 -2240 12035 -2220
rect 12005 -2270 12035 -2240
rect 12005 -2290 12010 -2270
rect 12030 -2290 12035 -2270
rect 12005 -2320 12035 -2290
rect 12005 -2340 12010 -2320
rect 12030 -2340 12035 -2320
rect 12005 -2370 12035 -2340
rect 12005 -2390 12010 -2370
rect 12030 -2390 12035 -2370
rect 12005 -2420 12035 -2390
rect 12005 -2440 12010 -2420
rect 12030 -2440 12035 -2420
rect 12005 -2470 12035 -2440
rect 12005 -2490 12010 -2470
rect 12030 -2490 12035 -2470
rect 12005 -2500 12035 -2490
rect 12065 -2120 12095 -2110
rect 12065 -2140 12070 -2120
rect 12090 -2140 12095 -2120
rect 12065 -2170 12095 -2140
rect 12065 -2190 12070 -2170
rect 12090 -2190 12095 -2170
rect 12065 -2220 12095 -2190
rect 12065 -2240 12070 -2220
rect 12090 -2240 12095 -2220
rect 12065 -2270 12095 -2240
rect 12065 -2290 12070 -2270
rect 12090 -2290 12095 -2270
rect 12065 -2320 12095 -2290
rect 12065 -2340 12070 -2320
rect 12090 -2340 12095 -2320
rect 12065 -2370 12095 -2340
rect 12065 -2390 12070 -2370
rect 12090 -2390 12095 -2370
rect 12065 -2420 12095 -2390
rect 12065 -2440 12070 -2420
rect 12090 -2440 12095 -2420
rect 12065 -2470 12095 -2440
rect 12065 -2490 12070 -2470
rect 12090 -2490 12095 -2470
rect 12065 -2500 12095 -2490
rect 12125 -2120 12155 -2110
rect 12125 -2140 12130 -2120
rect 12150 -2140 12155 -2120
rect 12125 -2170 12155 -2140
rect 12125 -2190 12130 -2170
rect 12150 -2190 12155 -2170
rect 12125 -2220 12155 -2190
rect 12125 -2240 12130 -2220
rect 12150 -2240 12155 -2220
rect 12125 -2270 12155 -2240
rect 12125 -2290 12130 -2270
rect 12150 -2290 12155 -2270
rect 12125 -2320 12155 -2290
rect 12125 -2340 12130 -2320
rect 12150 -2340 12155 -2320
rect 12125 -2370 12155 -2340
rect 12125 -2390 12130 -2370
rect 12150 -2390 12155 -2370
rect 12125 -2420 12155 -2390
rect 12125 -2440 12130 -2420
rect 12150 -2440 12155 -2420
rect 12125 -2470 12155 -2440
rect 12125 -2490 12130 -2470
rect 12150 -2490 12155 -2470
rect 12125 -2500 12155 -2490
rect 12185 -2120 12215 -2110
rect 12185 -2140 12190 -2120
rect 12210 -2140 12215 -2120
rect 12185 -2170 12215 -2140
rect 12185 -2190 12190 -2170
rect 12210 -2190 12215 -2170
rect 12185 -2220 12215 -2190
rect 12185 -2240 12190 -2220
rect 12210 -2240 12215 -2220
rect 12185 -2270 12215 -2240
rect 12185 -2290 12190 -2270
rect 12210 -2290 12215 -2270
rect 12185 -2320 12215 -2290
rect 12185 -2340 12190 -2320
rect 12210 -2340 12215 -2320
rect 12185 -2370 12215 -2340
rect 12185 -2390 12190 -2370
rect 12210 -2390 12215 -2370
rect 12185 -2420 12215 -2390
rect 12185 -2440 12190 -2420
rect 12210 -2440 12215 -2420
rect 12185 -2470 12215 -2440
rect 12185 -2490 12190 -2470
rect 12210 -2490 12215 -2470
rect 12185 -2500 12215 -2490
rect 12245 -2120 12275 -2110
rect 12245 -2140 12250 -2120
rect 12270 -2140 12275 -2120
rect 12245 -2170 12275 -2140
rect 12245 -2190 12250 -2170
rect 12270 -2190 12275 -2170
rect 12245 -2220 12275 -2190
rect 12245 -2240 12250 -2220
rect 12270 -2240 12275 -2220
rect 12245 -2270 12275 -2240
rect 12245 -2290 12250 -2270
rect 12270 -2290 12275 -2270
rect 12245 -2320 12275 -2290
rect 12245 -2340 12250 -2320
rect 12270 -2340 12275 -2320
rect 12245 -2370 12275 -2340
rect 12245 -2390 12250 -2370
rect 12270 -2390 12275 -2370
rect 12245 -2420 12275 -2390
rect 12245 -2440 12250 -2420
rect 12270 -2440 12275 -2420
rect 12245 -2470 12275 -2440
rect 12245 -2490 12250 -2470
rect 12270 -2490 12275 -2470
rect 12245 -2500 12275 -2490
rect 12305 -2120 12335 -2110
rect 12305 -2140 12310 -2120
rect 12330 -2140 12335 -2120
rect 12305 -2170 12335 -2140
rect 12305 -2190 12310 -2170
rect 12330 -2190 12335 -2170
rect 12305 -2220 12335 -2190
rect 12305 -2240 12310 -2220
rect 12330 -2240 12335 -2220
rect 12305 -2270 12335 -2240
rect 12305 -2290 12310 -2270
rect 12330 -2290 12335 -2270
rect 12305 -2320 12335 -2290
rect 12305 -2340 12310 -2320
rect 12330 -2340 12335 -2320
rect 12305 -2370 12335 -2340
rect 12305 -2390 12310 -2370
rect 12330 -2390 12335 -2370
rect 12305 -2420 12335 -2390
rect 12305 -2440 12310 -2420
rect 12330 -2440 12335 -2420
rect 12305 -2470 12335 -2440
rect 12305 -2490 12310 -2470
rect 12330 -2490 12335 -2470
rect 12305 -2500 12335 -2490
rect 12365 -2120 12395 -2110
rect 12365 -2140 12370 -2120
rect 12390 -2140 12395 -2120
rect 12365 -2170 12395 -2140
rect 12365 -2190 12370 -2170
rect 12390 -2190 12395 -2170
rect 12365 -2220 12395 -2190
rect 12365 -2240 12370 -2220
rect 12390 -2240 12395 -2220
rect 12365 -2270 12395 -2240
rect 12365 -2290 12370 -2270
rect 12390 -2290 12395 -2270
rect 12365 -2320 12395 -2290
rect 12365 -2340 12370 -2320
rect 12390 -2340 12395 -2320
rect 12365 -2370 12395 -2340
rect 12365 -2390 12370 -2370
rect 12390 -2390 12395 -2370
rect 12365 -2420 12395 -2390
rect 12365 -2440 12370 -2420
rect 12390 -2440 12395 -2420
rect 12365 -2470 12395 -2440
rect 12365 -2490 12370 -2470
rect 12390 -2490 12395 -2470
rect 12365 -2500 12395 -2490
rect 12425 -2120 12455 -2110
rect 12425 -2140 12430 -2120
rect 12450 -2140 12455 -2120
rect 12425 -2170 12455 -2140
rect 12425 -2190 12430 -2170
rect 12450 -2190 12455 -2170
rect 12425 -2220 12455 -2190
rect 12425 -2240 12430 -2220
rect 12450 -2240 12455 -2220
rect 12425 -2270 12455 -2240
rect 12425 -2290 12430 -2270
rect 12450 -2290 12455 -2270
rect 12425 -2320 12455 -2290
rect 12425 -2340 12430 -2320
rect 12450 -2340 12455 -2320
rect 12425 -2370 12455 -2340
rect 12425 -2390 12430 -2370
rect 12450 -2390 12455 -2370
rect 12425 -2420 12455 -2390
rect 12425 -2440 12430 -2420
rect 12450 -2440 12455 -2420
rect 12425 -2470 12455 -2440
rect 12425 -2490 12430 -2470
rect 12450 -2490 12455 -2470
rect 12425 -2500 12455 -2490
rect 12485 -2120 12515 -2110
rect 12485 -2140 12490 -2120
rect 12510 -2140 12515 -2120
rect 12485 -2170 12515 -2140
rect 12485 -2190 12490 -2170
rect 12510 -2190 12515 -2170
rect 12485 -2220 12515 -2190
rect 12485 -2240 12490 -2220
rect 12510 -2240 12515 -2220
rect 12485 -2270 12515 -2240
rect 12485 -2290 12490 -2270
rect 12510 -2290 12515 -2270
rect 12485 -2320 12515 -2290
rect 12485 -2340 12490 -2320
rect 12510 -2340 12515 -2320
rect 12485 -2370 12515 -2340
rect 12485 -2390 12490 -2370
rect 12510 -2390 12515 -2370
rect 12485 -2420 12515 -2390
rect 12485 -2440 12490 -2420
rect 12510 -2440 12515 -2420
rect 12485 -2470 12515 -2440
rect 12485 -2490 12490 -2470
rect 12510 -2490 12515 -2470
rect 12485 -2500 12515 -2490
rect 12545 -2120 12615 -2110
rect 12545 -2140 12550 -2120
rect 12570 -2140 12590 -2120
rect 12610 -2140 12615 -2120
rect 12545 -2170 12615 -2140
rect 12545 -2190 12550 -2170
rect 12570 -2190 12590 -2170
rect 12610 -2190 12615 -2170
rect 12545 -2220 12615 -2190
rect 12545 -2240 12550 -2220
rect 12570 -2240 12590 -2220
rect 12610 -2240 12615 -2220
rect 12545 -2270 12615 -2240
rect 12545 -2290 12550 -2270
rect 12570 -2290 12590 -2270
rect 12610 -2290 12615 -2270
rect 12545 -2320 12615 -2290
rect 12860 -2130 12930 -2100
rect 12860 -2150 12865 -2130
rect 12885 -2150 12905 -2130
rect 12925 -2150 12930 -2130
rect 12860 -2180 12930 -2150
rect 12860 -2200 12865 -2180
rect 12885 -2200 12905 -2180
rect 12925 -2200 12930 -2180
rect 12860 -2230 12930 -2200
rect 12860 -2250 12865 -2230
rect 12885 -2250 12905 -2230
rect 12925 -2250 12930 -2230
rect 12860 -2280 12930 -2250
rect 12860 -2300 12865 -2280
rect 12885 -2300 12905 -2280
rect 12925 -2300 12930 -2280
rect 12860 -2310 12930 -2300
rect 12955 -2030 12985 -2020
rect 12955 -2050 12960 -2030
rect 12980 -2050 12985 -2030
rect 12955 -2080 12985 -2050
rect 12955 -2100 12960 -2080
rect 12980 -2100 12985 -2080
rect 12955 -2130 12985 -2100
rect 12955 -2150 12960 -2130
rect 12980 -2150 12985 -2130
rect 12955 -2180 12985 -2150
rect 12955 -2200 12960 -2180
rect 12980 -2200 12985 -2180
rect 12955 -2230 12985 -2200
rect 12955 -2250 12960 -2230
rect 12980 -2250 12985 -2230
rect 12955 -2280 12985 -2250
rect 12955 -2300 12960 -2280
rect 12980 -2300 12985 -2280
rect 12955 -2310 12985 -2300
rect 13010 -2030 13040 -2020
rect 13010 -2050 13015 -2030
rect 13035 -2050 13040 -2030
rect 13010 -2080 13040 -2050
rect 13010 -2100 13015 -2080
rect 13035 -2100 13040 -2080
rect 13010 -2130 13040 -2100
rect 13010 -2150 13015 -2130
rect 13035 -2150 13040 -2130
rect 13010 -2180 13040 -2150
rect 13010 -2200 13015 -2180
rect 13035 -2200 13040 -2180
rect 13010 -2230 13040 -2200
rect 13010 -2250 13015 -2230
rect 13035 -2250 13040 -2230
rect 13010 -2280 13040 -2250
rect 13010 -2300 13015 -2280
rect 13035 -2300 13040 -2280
rect 13010 -2310 13040 -2300
rect 13065 -2030 13095 -2020
rect 13065 -2050 13070 -2030
rect 13090 -2050 13095 -2030
rect 13065 -2080 13095 -2050
rect 13065 -2100 13070 -2080
rect 13090 -2100 13095 -2080
rect 13065 -2130 13095 -2100
rect 13065 -2150 13070 -2130
rect 13090 -2150 13095 -2130
rect 13065 -2180 13095 -2150
rect 13065 -2200 13070 -2180
rect 13090 -2200 13095 -2180
rect 13065 -2230 13095 -2200
rect 13065 -2250 13070 -2230
rect 13090 -2250 13095 -2230
rect 13065 -2280 13095 -2250
rect 13065 -2300 13070 -2280
rect 13090 -2300 13095 -2280
rect 13065 -2310 13095 -2300
rect 13120 -2030 13150 -2020
rect 13120 -2050 13125 -2030
rect 13145 -2050 13150 -2030
rect 13120 -2080 13150 -2050
rect 13120 -2100 13125 -2080
rect 13145 -2100 13150 -2080
rect 13120 -2130 13150 -2100
rect 13120 -2150 13125 -2130
rect 13145 -2150 13150 -2130
rect 13120 -2180 13150 -2150
rect 13120 -2200 13125 -2180
rect 13145 -2200 13150 -2180
rect 13120 -2230 13150 -2200
rect 13120 -2250 13125 -2230
rect 13145 -2250 13150 -2230
rect 13120 -2280 13150 -2250
rect 13120 -2300 13125 -2280
rect 13145 -2300 13150 -2280
rect 13120 -2310 13150 -2300
rect 13175 -2030 13205 -2020
rect 13175 -2050 13180 -2030
rect 13200 -2050 13205 -2030
rect 13175 -2080 13205 -2050
rect 13175 -2100 13180 -2080
rect 13200 -2100 13205 -2080
rect 13175 -2130 13205 -2100
rect 13175 -2150 13180 -2130
rect 13200 -2150 13205 -2130
rect 13175 -2180 13205 -2150
rect 13175 -2200 13180 -2180
rect 13200 -2200 13205 -2180
rect 13175 -2230 13205 -2200
rect 13175 -2250 13180 -2230
rect 13200 -2250 13205 -2230
rect 13175 -2280 13205 -2250
rect 13175 -2300 13180 -2280
rect 13200 -2300 13205 -2280
rect 13175 -2310 13205 -2300
rect 13230 -2030 13260 -2020
rect 13230 -2050 13235 -2030
rect 13255 -2050 13260 -2030
rect 13230 -2080 13260 -2050
rect 13230 -2100 13235 -2080
rect 13255 -2100 13260 -2080
rect 13230 -2130 13260 -2100
rect 13230 -2150 13235 -2130
rect 13255 -2150 13260 -2130
rect 13230 -2180 13260 -2150
rect 13230 -2200 13235 -2180
rect 13255 -2200 13260 -2180
rect 13230 -2230 13260 -2200
rect 13230 -2250 13235 -2230
rect 13255 -2250 13260 -2230
rect 13230 -2280 13260 -2250
rect 13230 -2300 13235 -2280
rect 13255 -2300 13260 -2280
rect 13230 -2310 13260 -2300
rect 13285 -2030 13315 -2020
rect 13285 -2050 13290 -2030
rect 13310 -2050 13315 -2030
rect 13285 -2080 13315 -2050
rect 13285 -2100 13290 -2080
rect 13310 -2100 13315 -2080
rect 13285 -2130 13315 -2100
rect 13285 -2150 13290 -2130
rect 13310 -2150 13315 -2130
rect 13285 -2180 13315 -2150
rect 13285 -2200 13290 -2180
rect 13310 -2200 13315 -2180
rect 13285 -2230 13315 -2200
rect 13285 -2250 13290 -2230
rect 13310 -2250 13315 -2230
rect 13285 -2280 13315 -2250
rect 13285 -2300 13290 -2280
rect 13310 -2300 13315 -2280
rect 13285 -2310 13315 -2300
rect 13340 -2030 13370 -2020
rect 13340 -2050 13345 -2030
rect 13365 -2050 13370 -2030
rect 13340 -2080 13370 -2050
rect 13340 -2100 13345 -2080
rect 13365 -2100 13370 -2080
rect 13340 -2130 13370 -2100
rect 13340 -2150 13345 -2130
rect 13365 -2150 13370 -2130
rect 13340 -2180 13370 -2150
rect 13340 -2200 13345 -2180
rect 13365 -2200 13370 -2180
rect 13340 -2230 13370 -2200
rect 13340 -2250 13345 -2230
rect 13365 -2250 13370 -2230
rect 13340 -2280 13370 -2250
rect 13340 -2300 13345 -2280
rect 13365 -2300 13370 -2280
rect 13340 -2310 13370 -2300
rect 13395 -2030 13425 -2020
rect 13395 -2050 13400 -2030
rect 13420 -2050 13425 -2030
rect 13395 -2080 13425 -2050
rect 13395 -2100 13400 -2080
rect 13420 -2100 13425 -2080
rect 13395 -2130 13425 -2100
rect 13395 -2150 13400 -2130
rect 13420 -2150 13425 -2130
rect 13395 -2180 13425 -2150
rect 13395 -2200 13400 -2180
rect 13420 -2200 13425 -2180
rect 13395 -2230 13425 -2200
rect 13395 -2250 13400 -2230
rect 13420 -2250 13425 -2230
rect 13395 -2280 13425 -2250
rect 13395 -2300 13400 -2280
rect 13420 -2300 13425 -2280
rect 13395 -2310 13425 -2300
rect 13450 -2030 13480 -2020
rect 13450 -2050 13455 -2030
rect 13475 -2050 13480 -2030
rect 13450 -2080 13480 -2050
rect 13450 -2100 13455 -2080
rect 13475 -2100 13480 -2080
rect 13450 -2130 13480 -2100
rect 13450 -2150 13455 -2130
rect 13475 -2150 13480 -2130
rect 13450 -2180 13480 -2150
rect 13450 -2200 13455 -2180
rect 13475 -2200 13480 -2180
rect 13450 -2230 13480 -2200
rect 13450 -2250 13455 -2230
rect 13475 -2250 13480 -2230
rect 13450 -2280 13480 -2250
rect 13450 -2300 13455 -2280
rect 13475 -2300 13480 -2280
rect 13450 -2310 13480 -2300
rect 13505 -2030 13535 -2020
rect 13505 -2050 13510 -2030
rect 13530 -2050 13535 -2030
rect 13505 -2080 13535 -2050
rect 13505 -2100 13510 -2080
rect 13530 -2100 13535 -2080
rect 13505 -2130 13535 -2100
rect 13505 -2150 13510 -2130
rect 13530 -2150 13535 -2130
rect 13505 -2180 13535 -2150
rect 13505 -2200 13510 -2180
rect 13530 -2200 13535 -2180
rect 13505 -2230 13535 -2200
rect 13505 -2250 13510 -2230
rect 13530 -2250 13535 -2230
rect 13505 -2280 13535 -2250
rect 13505 -2300 13510 -2280
rect 13530 -2300 13535 -2280
rect 13505 -2310 13535 -2300
rect 13560 -2030 13590 -2020
rect 13560 -2050 13565 -2030
rect 13585 -2050 13590 -2030
rect 13560 -2080 13590 -2050
rect 13560 -2100 13565 -2080
rect 13585 -2100 13590 -2080
rect 13560 -2130 13590 -2100
rect 13560 -2150 13565 -2130
rect 13585 -2150 13590 -2130
rect 13560 -2180 13590 -2150
rect 13560 -2200 13565 -2180
rect 13585 -2200 13590 -2180
rect 13560 -2230 13590 -2200
rect 13560 -2250 13565 -2230
rect 13585 -2250 13590 -2230
rect 13560 -2280 13590 -2250
rect 13560 -2300 13565 -2280
rect 13585 -2300 13590 -2280
rect 13560 -2310 13590 -2300
rect 13615 -2030 13645 -2020
rect 13615 -2050 13620 -2030
rect 13640 -2050 13645 -2030
rect 13615 -2080 13645 -2050
rect 13615 -2100 13620 -2080
rect 13640 -2100 13645 -2080
rect 13615 -2130 13645 -2100
rect 13615 -2150 13620 -2130
rect 13640 -2150 13645 -2130
rect 13615 -2180 13645 -2150
rect 13615 -2200 13620 -2180
rect 13640 -2200 13645 -2180
rect 13615 -2230 13645 -2200
rect 13615 -2250 13620 -2230
rect 13640 -2250 13645 -2230
rect 13615 -2280 13645 -2250
rect 13615 -2300 13620 -2280
rect 13640 -2300 13645 -2280
rect 13615 -2310 13645 -2300
rect 13670 -2030 13700 -2020
rect 13670 -2050 13675 -2030
rect 13695 -2050 13700 -2030
rect 13670 -2080 13700 -2050
rect 13670 -2100 13675 -2080
rect 13695 -2100 13700 -2080
rect 13670 -2130 13700 -2100
rect 13670 -2150 13675 -2130
rect 13695 -2150 13700 -2130
rect 13670 -2180 13700 -2150
rect 13670 -2200 13675 -2180
rect 13695 -2200 13700 -2180
rect 13670 -2230 13700 -2200
rect 13670 -2250 13675 -2230
rect 13695 -2250 13700 -2230
rect 13670 -2280 13700 -2250
rect 13670 -2300 13675 -2280
rect 13695 -2300 13700 -2280
rect 13670 -2310 13700 -2300
rect 13725 -2030 13755 -2020
rect 13725 -2050 13730 -2030
rect 13750 -2050 13755 -2030
rect 13725 -2080 13755 -2050
rect 13725 -2100 13730 -2080
rect 13750 -2100 13755 -2080
rect 13725 -2130 13755 -2100
rect 13725 -2150 13730 -2130
rect 13750 -2150 13755 -2130
rect 13725 -2180 13755 -2150
rect 13725 -2200 13730 -2180
rect 13750 -2200 13755 -2180
rect 13725 -2230 13755 -2200
rect 13725 -2250 13730 -2230
rect 13750 -2250 13755 -2230
rect 13725 -2280 13755 -2250
rect 13725 -2300 13730 -2280
rect 13750 -2300 13755 -2280
rect 13725 -2310 13755 -2300
rect 13780 -2030 13810 -2020
rect 13780 -2050 13785 -2030
rect 13805 -2050 13810 -2030
rect 13780 -2080 13810 -2050
rect 13780 -2100 13785 -2080
rect 13805 -2100 13810 -2080
rect 13780 -2130 13810 -2100
rect 13780 -2150 13785 -2130
rect 13805 -2150 13810 -2130
rect 13780 -2180 13810 -2150
rect 13780 -2200 13785 -2180
rect 13805 -2200 13810 -2180
rect 13780 -2230 13810 -2200
rect 13780 -2250 13785 -2230
rect 13805 -2250 13810 -2230
rect 13780 -2280 13810 -2250
rect 13780 -2300 13785 -2280
rect 13805 -2300 13810 -2280
rect 13780 -2310 13810 -2300
rect 13835 -2030 13865 -2020
rect 13835 -2050 13840 -2030
rect 13860 -2050 13865 -2030
rect 13835 -2080 13865 -2050
rect 13835 -2100 13840 -2080
rect 13860 -2100 13865 -2080
rect 13835 -2130 13865 -2100
rect 13835 -2150 13840 -2130
rect 13860 -2150 13865 -2130
rect 13835 -2180 13865 -2150
rect 13835 -2200 13840 -2180
rect 13860 -2200 13865 -2180
rect 13835 -2230 13865 -2200
rect 13835 -2250 13840 -2230
rect 13860 -2250 13865 -2230
rect 13835 -2280 13865 -2250
rect 13835 -2300 13840 -2280
rect 13860 -2300 13865 -2280
rect 13835 -2310 13865 -2300
rect 13890 -2030 13920 -2020
rect 13890 -2050 13895 -2030
rect 13915 -2050 13920 -2030
rect 13890 -2080 13920 -2050
rect 13890 -2100 13895 -2080
rect 13915 -2100 13920 -2080
rect 13890 -2130 13920 -2100
rect 13890 -2150 13895 -2130
rect 13915 -2150 13920 -2130
rect 13890 -2180 13920 -2150
rect 13890 -2200 13895 -2180
rect 13915 -2200 13920 -2180
rect 13890 -2230 13920 -2200
rect 13890 -2250 13895 -2230
rect 13915 -2250 13920 -2230
rect 13890 -2280 13920 -2250
rect 13890 -2300 13895 -2280
rect 13915 -2300 13920 -2280
rect 13890 -2310 13920 -2300
rect 13945 -2030 13975 -2020
rect 13945 -2050 13950 -2030
rect 13970 -2050 13975 -2030
rect 13945 -2080 13975 -2050
rect 13945 -2100 13950 -2080
rect 13970 -2100 13975 -2080
rect 13945 -2130 13975 -2100
rect 13945 -2150 13950 -2130
rect 13970 -2150 13975 -2130
rect 13945 -2180 13975 -2150
rect 13945 -2200 13950 -2180
rect 13970 -2200 13975 -2180
rect 13945 -2230 13975 -2200
rect 13945 -2250 13950 -2230
rect 13970 -2250 13975 -2230
rect 13945 -2280 13975 -2250
rect 13945 -2300 13950 -2280
rect 13970 -2300 13975 -2280
rect 13945 -2310 13975 -2300
rect 14000 -2030 14030 -2020
rect 14000 -2050 14005 -2030
rect 14025 -2050 14030 -2030
rect 14000 -2080 14030 -2050
rect 14000 -2100 14005 -2080
rect 14025 -2100 14030 -2080
rect 14000 -2130 14030 -2100
rect 14000 -2150 14005 -2130
rect 14025 -2150 14030 -2130
rect 14000 -2180 14030 -2150
rect 14000 -2200 14005 -2180
rect 14025 -2200 14030 -2180
rect 14000 -2230 14030 -2200
rect 14000 -2250 14005 -2230
rect 14025 -2250 14030 -2230
rect 14000 -2280 14030 -2250
rect 14000 -2300 14005 -2280
rect 14025 -2300 14030 -2280
rect 14000 -2310 14030 -2300
rect 14055 -2030 14085 -2020
rect 14055 -2050 14060 -2030
rect 14080 -2050 14085 -2030
rect 14055 -2080 14085 -2050
rect 14055 -2100 14060 -2080
rect 14080 -2100 14085 -2080
rect 14055 -2130 14085 -2100
rect 14055 -2150 14060 -2130
rect 14080 -2150 14085 -2130
rect 14055 -2180 14085 -2150
rect 14055 -2200 14060 -2180
rect 14080 -2200 14085 -2180
rect 14055 -2230 14085 -2200
rect 14055 -2250 14060 -2230
rect 14080 -2250 14085 -2230
rect 14055 -2280 14085 -2250
rect 14055 -2300 14060 -2280
rect 14080 -2300 14085 -2280
rect 14055 -2310 14085 -2300
rect 14110 -2030 14180 -2020
rect 14110 -2050 14115 -2030
rect 14135 -2050 14155 -2030
rect 14175 -2050 14180 -2030
rect 14110 -2080 14180 -2050
rect 14110 -2100 14115 -2080
rect 14135 -2100 14155 -2080
rect 14175 -2100 14180 -2080
rect 14110 -2130 14180 -2100
rect 14110 -2150 14115 -2130
rect 14135 -2150 14155 -2130
rect 14175 -2150 14180 -2130
rect 14110 -2180 14180 -2150
rect 14110 -2200 14115 -2180
rect 14135 -2200 14155 -2180
rect 14175 -2200 14180 -2180
rect 14110 -2230 14180 -2200
rect 14110 -2250 14115 -2230
rect 14135 -2250 14155 -2230
rect 14175 -2250 14180 -2230
rect 14110 -2280 14180 -2250
rect 14110 -2300 14115 -2280
rect 14135 -2300 14155 -2280
rect 14175 -2300 14180 -2280
rect 14110 -2310 14180 -2300
rect 12545 -2340 12550 -2320
rect 12570 -2340 12590 -2320
rect 12610 -2340 12615 -2320
rect 12865 -2330 12885 -2310
rect 13015 -2330 13035 -2310
rect 13125 -2330 13145 -2310
rect 13235 -2330 13255 -2310
rect 13345 -2330 13365 -2310
rect 13455 -2330 13475 -2310
rect 13565 -2330 13585 -2310
rect 13675 -2330 13695 -2310
rect 13785 -2330 13805 -2310
rect 13895 -2330 13915 -2310
rect 14005 -2330 14025 -2310
rect 14155 -2330 14175 -2310
rect 12545 -2370 12615 -2340
rect 12855 -2340 12895 -2330
rect 12855 -2360 12865 -2340
rect 12885 -2360 12895 -2340
rect 12855 -2370 12895 -2360
rect 13005 -2340 13045 -2330
rect 13005 -2360 13015 -2340
rect 13035 -2360 13045 -2340
rect 13005 -2370 13045 -2360
rect 13063 -2340 13097 -2330
rect 13063 -2360 13071 -2340
rect 13089 -2360 13097 -2340
rect 13063 -2370 13097 -2360
rect 13115 -2340 13155 -2330
rect 13115 -2360 13125 -2340
rect 13145 -2360 13155 -2340
rect 13115 -2370 13155 -2360
rect 13225 -2340 13265 -2330
rect 13225 -2360 13235 -2340
rect 13255 -2360 13265 -2340
rect 13225 -2370 13265 -2360
rect 13335 -2340 13375 -2330
rect 13335 -2360 13345 -2340
rect 13365 -2360 13375 -2340
rect 13335 -2370 13375 -2360
rect 13445 -2340 13485 -2330
rect 13445 -2360 13455 -2340
rect 13475 -2360 13485 -2340
rect 13445 -2370 13485 -2360
rect 13555 -2340 13595 -2330
rect 13555 -2360 13565 -2340
rect 13585 -2360 13595 -2340
rect 13555 -2370 13595 -2360
rect 13665 -2340 13705 -2330
rect 13665 -2360 13675 -2340
rect 13695 -2360 13705 -2340
rect 13665 -2370 13705 -2360
rect 13775 -2340 13815 -2330
rect 13775 -2360 13785 -2340
rect 13805 -2360 13815 -2340
rect 13775 -2370 13815 -2360
rect 13885 -2340 13925 -2330
rect 13885 -2360 13895 -2340
rect 13915 -2360 13925 -2340
rect 13885 -2370 13925 -2360
rect 13995 -2340 14035 -2330
rect 13995 -2360 14005 -2340
rect 14025 -2360 14035 -2340
rect 13995 -2370 14035 -2360
rect 14145 -2340 14185 -2330
rect 14145 -2360 14155 -2340
rect 14175 -2360 14185 -2340
rect 14145 -2370 14185 -2360
rect 12545 -2390 12550 -2370
rect 12570 -2390 12590 -2370
rect 12610 -2390 12615 -2370
rect 12545 -2420 12615 -2390
rect 12545 -2440 12550 -2420
rect 12570 -2440 12590 -2420
rect 12610 -2440 12615 -2420
rect 12950 -2400 12990 -2390
rect 12950 -2420 12960 -2400
rect 12980 -2420 12990 -2400
rect 12950 -2430 12990 -2420
rect 13060 -2400 13100 -2390
rect 13060 -2420 13070 -2400
rect 13090 -2420 13100 -2400
rect 13060 -2430 13100 -2420
rect 13170 -2400 13210 -2390
rect 13170 -2420 13180 -2400
rect 13200 -2420 13210 -2400
rect 13170 -2430 13210 -2420
rect 13280 -2400 13320 -2390
rect 13280 -2420 13290 -2400
rect 13310 -2420 13320 -2400
rect 13280 -2430 13320 -2420
rect 13390 -2400 13430 -2390
rect 13390 -2420 13400 -2400
rect 13420 -2420 13430 -2400
rect 13390 -2430 13430 -2420
rect 13500 -2400 13540 -2390
rect 13500 -2420 13510 -2400
rect 13530 -2420 13540 -2400
rect 13500 -2430 13540 -2420
rect 13610 -2400 13650 -2390
rect 13610 -2420 13620 -2400
rect 13640 -2420 13650 -2400
rect 13610 -2430 13650 -2420
rect 13720 -2400 13760 -2390
rect 13720 -2420 13730 -2400
rect 13750 -2420 13760 -2400
rect 13720 -2430 13760 -2420
rect 13830 -2400 13870 -2390
rect 13830 -2420 13840 -2400
rect 13860 -2420 13870 -2400
rect 13830 -2430 13870 -2420
rect 13940 -2400 13980 -2390
rect 13940 -2420 13950 -2400
rect 13970 -2420 13980 -2400
rect 13940 -2430 13980 -2420
rect 14050 -2400 14090 -2390
rect 14050 -2420 14060 -2400
rect 14080 -2420 14090 -2400
rect 14050 -2430 14090 -2420
rect 12545 -2470 12615 -2440
rect 12960 -2450 12980 -2430
rect 13070 -2450 13090 -2430
rect 13180 -2450 13200 -2430
rect 13290 -2450 13310 -2430
rect 13400 -2450 13420 -2430
rect 13510 -2450 13530 -2430
rect 13620 -2450 13640 -2430
rect 13730 -2450 13750 -2430
rect 13840 -2450 13860 -2430
rect 13950 -2450 13970 -2430
rect 14060 -2450 14080 -2430
rect 12545 -2490 12550 -2470
rect 12570 -2490 12590 -2470
rect 12610 -2490 12615 -2470
rect 12545 -2500 12615 -2490
rect 12860 -2460 12930 -2450
rect 12860 -2480 12865 -2460
rect 12885 -2480 12905 -2460
rect 12925 -2480 12930 -2460
rect 11290 -2520 11310 -2500
rect 11410 -2520 11430 -2500
rect 11530 -2520 11550 -2500
rect 11650 -2520 11670 -2500
rect 11770 -2520 11790 -2500
rect 11890 -2520 11910 -2500
rect 12010 -2520 12030 -2500
rect 12130 -2520 12150 -2500
rect 12250 -2520 12270 -2500
rect 12370 -2520 12390 -2500
rect 12490 -2520 12510 -2500
rect 12860 -2510 12930 -2480
rect 11280 -2530 11320 -2520
rect 11280 -2550 11290 -2530
rect 11310 -2550 11320 -2530
rect 11280 -2560 11320 -2550
rect 11400 -2530 11440 -2520
rect 11400 -2550 11410 -2530
rect 11430 -2550 11440 -2530
rect 11400 -2560 11440 -2550
rect 11520 -2530 11560 -2520
rect 11520 -2550 11530 -2530
rect 11550 -2550 11560 -2530
rect 11520 -2560 11560 -2550
rect 11640 -2530 11680 -2520
rect 11640 -2550 11650 -2530
rect 11670 -2550 11680 -2530
rect 11640 -2560 11680 -2550
rect 11760 -2530 11800 -2520
rect 11760 -2550 11770 -2530
rect 11790 -2550 11800 -2530
rect 11760 -2560 11800 -2550
rect 11823 -2530 11857 -2520
rect 11823 -2550 11831 -2530
rect 11849 -2550 11857 -2530
rect 11823 -2560 11857 -2550
rect 11880 -2530 11920 -2520
rect 11880 -2550 11890 -2530
rect 11910 -2550 11920 -2530
rect 11880 -2560 11920 -2550
rect 12000 -2530 12040 -2520
rect 12000 -2550 12010 -2530
rect 12030 -2550 12040 -2530
rect 12000 -2560 12040 -2550
rect 12120 -2530 12160 -2520
rect 12120 -2550 12130 -2530
rect 12150 -2550 12160 -2530
rect 12120 -2560 12160 -2550
rect 12240 -2530 12280 -2520
rect 12240 -2550 12250 -2530
rect 12270 -2550 12280 -2530
rect 12240 -2560 12280 -2550
rect 12360 -2530 12400 -2520
rect 12360 -2550 12370 -2530
rect 12390 -2550 12400 -2530
rect 12360 -2560 12400 -2550
rect 12480 -2530 12520 -2520
rect 12480 -2550 12490 -2530
rect 12510 -2550 12520 -2530
rect 12860 -2530 12865 -2510
rect 12885 -2530 12905 -2510
rect 12925 -2530 12930 -2510
rect 12860 -2540 12930 -2530
rect 12955 -2460 12985 -2450
rect 12955 -2480 12960 -2460
rect 12980 -2480 12985 -2460
rect 12955 -2510 12985 -2480
rect 12955 -2530 12960 -2510
rect 12980 -2530 12985 -2510
rect 12955 -2540 12985 -2530
rect 13010 -2460 13040 -2450
rect 13010 -2480 13015 -2460
rect 13035 -2480 13040 -2460
rect 13010 -2510 13040 -2480
rect 13010 -2530 13015 -2510
rect 13035 -2530 13040 -2510
rect 13010 -2540 13040 -2530
rect 13065 -2460 13095 -2450
rect 13065 -2480 13070 -2460
rect 13090 -2480 13095 -2460
rect 13065 -2510 13095 -2480
rect 13065 -2530 13070 -2510
rect 13090 -2530 13095 -2510
rect 13065 -2540 13095 -2530
rect 13120 -2460 13150 -2450
rect 13120 -2480 13125 -2460
rect 13145 -2480 13150 -2460
rect 13120 -2510 13150 -2480
rect 13120 -2530 13125 -2510
rect 13145 -2530 13150 -2510
rect 13120 -2540 13150 -2530
rect 13175 -2460 13205 -2450
rect 13175 -2480 13180 -2460
rect 13200 -2480 13205 -2460
rect 13175 -2510 13205 -2480
rect 13175 -2530 13180 -2510
rect 13200 -2530 13205 -2510
rect 13175 -2540 13205 -2530
rect 13230 -2460 13260 -2450
rect 13230 -2480 13235 -2460
rect 13255 -2480 13260 -2460
rect 13230 -2510 13260 -2480
rect 13230 -2530 13235 -2510
rect 13255 -2530 13260 -2510
rect 13230 -2540 13260 -2530
rect 13285 -2460 13315 -2450
rect 13285 -2480 13290 -2460
rect 13310 -2480 13315 -2460
rect 13285 -2510 13315 -2480
rect 13285 -2530 13290 -2510
rect 13310 -2530 13315 -2510
rect 13285 -2540 13315 -2530
rect 13340 -2460 13370 -2450
rect 13340 -2480 13345 -2460
rect 13365 -2480 13370 -2460
rect 13340 -2510 13370 -2480
rect 13340 -2530 13345 -2510
rect 13365 -2530 13370 -2510
rect 13340 -2540 13370 -2530
rect 13395 -2460 13425 -2450
rect 13395 -2480 13400 -2460
rect 13420 -2480 13425 -2460
rect 13395 -2510 13425 -2480
rect 13395 -2530 13400 -2510
rect 13420 -2530 13425 -2510
rect 13395 -2540 13425 -2530
rect 13450 -2460 13480 -2450
rect 13450 -2480 13455 -2460
rect 13475 -2480 13480 -2460
rect 13450 -2510 13480 -2480
rect 13450 -2530 13455 -2510
rect 13475 -2530 13480 -2510
rect 13450 -2540 13480 -2530
rect 13505 -2460 13535 -2450
rect 13505 -2480 13510 -2460
rect 13530 -2480 13535 -2460
rect 13505 -2510 13535 -2480
rect 13505 -2530 13510 -2510
rect 13530 -2530 13535 -2510
rect 13505 -2540 13535 -2530
rect 13560 -2460 13590 -2450
rect 13560 -2480 13565 -2460
rect 13585 -2480 13590 -2460
rect 13560 -2510 13590 -2480
rect 13560 -2530 13565 -2510
rect 13585 -2530 13590 -2510
rect 13560 -2540 13590 -2530
rect 13615 -2460 13645 -2450
rect 13615 -2480 13620 -2460
rect 13640 -2480 13645 -2460
rect 13615 -2510 13645 -2480
rect 13615 -2530 13620 -2510
rect 13640 -2530 13645 -2510
rect 13615 -2540 13645 -2530
rect 13670 -2460 13700 -2450
rect 13670 -2480 13675 -2460
rect 13695 -2480 13700 -2460
rect 13670 -2510 13700 -2480
rect 13670 -2530 13675 -2510
rect 13695 -2530 13700 -2510
rect 13670 -2540 13700 -2530
rect 13725 -2460 13755 -2450
rect 13725 -2480 13730 -2460
rect 13750 -2480 13755 -2460
rect 13725 -2510 13755 -2480
rect 13725 -2530 13730 -2510
rect 13750 -2530 13755 -2510
rect 13725 -2540 13755 -2530
rect 13780 -2460 13810 -2450
rect 13780 -2480 13785 -2460
rect 13805 -2480 13810 -2460
rect 13780 -2510 13810 -2480
rect 13780 -2530 13785 -2510
rect 13805 -2530 13810 -2510
rect 13780 -2540 13810 -2530
rect 13835 -2460 13865 -2450
rect 13835 -2480 13840 -2460
rect 13860 -2480 13865 -2460
rect 13835 -2510 13865 -2480
rect 13835 -2530 13840 -2510
rect 13860 -2530 13865 -2510
rect 13835 -2540 13865 -2530
rect 13890 -2460 13920 -2450
rect 13890 -2480 13895 -2460
rect 13915 -2480 13920 -2460
rect 13890 -2510 13920 -2480
rect 13890 -2530 13895 -2510
rect 13915 -2530 13920 -2510
rect 13890 -2540 13920 -2530
rect 13945 -2460 13975 -2450
rect 13945 -2480 13950 -2460
rect 13970 -2480 13975 -2460
rect 13945 -2510 13975 -2480
rect 13945 -2530 13950 -2510
rect 13970 -2530 13975 -2510
rect 13945 -2540 13975 -2530
rect 14000 -2460 14030 -2450
rect 14000 -2480 14005 -2460
rect 14025 -2480 14030 -2460
rect 14000 -2510 14030 -2480
rect 14000 -2530 14005 -2510
rect 14025 -2530 14030 -2510
rect 14000 -2540 14030 -2530
rect 14055 -2460 14085 -2450
rect 14055 -2480 14060 -2460
rect 14080 -2480 14085 -2460
rect 14055 -2510 14085 -2480
rect 14055 -2530 14060 -2510
rect 14080 -2530 14085 -2510
rect 14055 -2540 14085 -2530
rect 14110 -2460 14180 -2450
rect 14110 -2480 14115 -2460
rect 14135 -2480 14155 -2460
rect 14175 -2480 14180 -2460
rect 14110 -2510 14180 -2480
rect 14110 -2530 14115 -2510
rect 14135 -2530 14155 -2510
rect 14175 -2530 14180 -2510
rect 14110 -2540 14180 -2530
rect 12480 -2560 12520 -2550
rect 12865 -2560 12885 -2540
rect 13015 -2560 13035 -2540
rect 13125 -2560 13145 -2540
rect 13235 -2560 13255 -2540
rect 13345 -2560 13365 -2540
rect 13455 -2560 13475 -2540
rect 13565 -2560 13585 -2540
rect 13675 -2560 13695 -2540
rect 13785 -2560 13805 -2540
rect 13895 -2560 13915 -2540
rect 14005 -2560 14025 -2540
rect 14155 -2560 14175 -2540
rect 12855 -2570 12895 -2560
rect 12855 -2590 12865 -2570
rect 12885 -2590 12895 -2570
rect 12855 -2600 12895 -2590
rect 13005 -2570 13045 -2560
rect 13005 -2590 13015 -2570
rect 13035 -2590 13045 -2570
rect 13005 -2600 13045 -2590
rect 13115 -2570 13155 -2560
rect 13115 -2590 13125 -2570
rect 13145 -2590 13155 -2570
rect 13115 -2600 13155 -2590
rect 13225 -2570 13265 -2560
rect 13225 -2590 13235 -2570
rect 13255 -2590 13265 -2570
rect 13225 -2600 13265 -2590
rect 13335 -2570 13375 -2560
rect 13335 -2590 13345 -2570
rect 13365 -2590 13375 -2570
rect 13335 -2600 13375 -2590
rect 13445 -2570 13485 -2560
rect 13445 -2590 13455 -2570
rect 13475 -2590 13485 -2570
rect 13445 -2600 13485 -2590
rect 13555 -2570 13595 -2560
rect 13555 -2590 13565 -2570
rect 13585 -2590 13595 -2570
rect 13555 -2600 13595 -2590
rect 13665 -2570 13705 -2560
rect 13665 -2590 13675 -2570
rect 13695 -2590 13705 -2570
rect 13665 -2600 13705 -2590
rect 13775 -2570 13815 -2560
rect 13775 -2590 13785 -2570
rect 13805 -2590 13815 -2570
rect 13775 -2600 13815 -2590
rect 13885 -2570 13925 -2560
rect 13885 -2590 13895 -2570
rect 13915 -2590 13925 -2570
rect 13885 -2600 13925 -2590
rect 13995 -2570 14035 -2560
rect 13995 -2590 14005 -2570
rect 14025 -2590 14035 -2570
rect 13995 -2600 14035 -2590
rect 14145 -2570 14185 -2560
rect 14145 -2590 14155 -2570
rect 14175 -2590 14185 -2570
rect 14145 -2600 14185 -2590
rect 12975 -2630 13015 -2620
rect 12975 -2650 12985 -2630
rect 13005 -2650 13015 -2630
rect 12975 -2660 13015 -2650
rect 12855 -2690 12895 -2680
rect 12855 -2710 12865 -2690
rect 12885 -2710 12895 -2690
rect 12855 -2720 12895 -2710
rect 13005 -2690 13045 -2680
rect 13005 -2710 13015 -2690
rect 13035 -2710 13045 -2690
rect 13005 -2720 13045 -2710
rect 13115 -2690 13155 -2680
rect 13115 -2710 13125 -2690
rect 13145 -2710 13155 -2690
rect 13115 -2720 13155 -2710
rect 13225 -2690 13265 -2680
rect 13225 -2710 13235 -2690
rect 13255 -2710 13265 -2690
rect 13225 -2720 13265 -2710
rect 13335 -2690 13375 -2680
rect 13335 -2710 13345 -2690
rect 13365 -2710 13375 -2690
rect 13335 -2720 13375 -2710
rect 13445 -2690 13485 -2680
rect 13445 -2710 13455 -2690
rect 13475 -2710 13485 -2690
rect 13445 -2720 13485 -2710
rect 13555 -2690 13595 -2680
rect 13555 -2710 13565 -2690
rect 13585 -2710 13595 -2690
rect 13555 -2720 13595 -2710
rect 13665 -2690 13705 -2680
rect 13665 -2710 13675 -2690
rect 13695 -2710 13705 -2690
rect 13665 -2720 13705 -2710
rect 13775 -2690 13815 -2680
rect 13775 -2710 13785 -2690
rect 13805 -2710 13815 -2690
rect 13775 -2720 13815 -2710
rect 13885 -2690 13925 -2680
rect 13885 -2710 13895 -2690
rect 13915 -2710 13925 -2690
rect 13885 -2720 13925 -2710
rect 13995 -2690 14035 -2680
rect 13995 -2710 14005 -2690
rect 14025 -2710 14035 -2690
rect 13995 -2720 14035 -2710
rect 14145 -2690 14185 -2680
rect 14145 -2710 14155 -2690
rect 14175 -2710 14185 -2690
rect 14145 -2720 14185 -2710
rect 12865 -2740 12885 -2720
rect 13015 -2740 13035 -2720
rect 13125 -2740 13145 -2720
rect 13235 -2740 13255 -2720
rect 13345 -2740 13365 -2720
rect 13455 -2740 13475 -2720
rect 13565 -2740 13585 -2720
rect 13675 -2740 13695 -2720
rect 13785 -2740 13805 -2720
rect 13895 -2740 13915 -2720
rect 14005 -2740 14025 -2720
rect 14155 -2740 14175 -2720
rect 12860 -2750 12930 -2740
rect 12860 -2770 12865 -2750
rect 12885 -2770 12905 -2750
rect 12925 -2770 12930 -2750
rect 12860 -2800 12930 -2770
rect 11330 -2825 11370 -2815
rect 11330 -2845 11340 -2825
rect 11360 -2845 11370 -2825
rect 11330 -2855 11370 -2845
rect 11440 -2825 11480 -2815
rect 11440 -2845 11450 -2825
rect 11470 -2845 11480 -2825
rect 11440 -2855 11480 -2845
rect 11550 -2825 11590 -2815
rect 11550 -2845 11560 -2825
rect 11580 -2845 11590 -2825
rect 11550 -2855 11590 -2845
rect 11660 -2825 11700 -2815
rect 11660 -2845 11670 -2825
rect 11690 -2845 11700 -2825
rect 11660 -2855 11700 -2845
rect 11770 -2825 11810 -2815
rect 11770 -2845 11780 -2825
rect 11800 -2845 11810 -2825
rect 11770 -2855 11810 -2845
rect 11880 -2825 11920 -2815
rect 11880 -2845 11890 -2825
rect 11910 -2845 11920 -2825
rect 11880 -2855 11920 -2845
rect 11990 -2825 12030 -2815
rect 11990 -2845 12000 -2825
rect 12020 -2845 12030 -2825
rect 11990 -2855 12030 -2845
rect 12100 -2825 12140 -2815
rect 12100 -2845 12110 -2825
rect 12130 -2845 12140 -2825
rect 12100 -2855 12140 -2845
rect 12210 -2825 12250 -2815
rect 12210 -2845 12220 -2825
rect 12240 -2845 12250 -2825
rect 12210 -2855 12250 -2845
rect 12320 -2825 12360 -2815
rect 12320 -2845 12330 -2825
rect 12350 -2845 12360 -2825
rect 12320 -2855 12360 -2845
rect 12430 -2825 12470 -2815
rect 12430 -2845 12440 -2825
rect 12460 -2845 12470 -2825
rect 12430 -2855 12470 -2845
rect 12860 -2820 12865 -2800
rect 12885 -2820 12905 -2800
rect 12925 -2820 12930 -2800
rect 12860 -2850 12930 -2820
rect 11340 -2875 11360 -2855
rect 11450 -2875 11470 -2855
rect 11560 -2875 11580 -2855
rect 11670 -2875 11690 -2855
rect 11780 -2875 11800 -2855
rect 11890 -2875 11910 -2855
rect 12000 -2875 12020 -2855
rect 12110 -2875 12130 -2855
rect 12220 -2875 12240 -2855
rect 12330 -2875 12350 -2855
rect 12440 -2875 12460 -2855
rect 12860 -2870 12865 -2850
rect 12885 -2870 12905 -2850
rect 12925 -2870 12930 -2850
rect 11240 -2885 11310 -2875
rect 11240 -2905 11245 -2885
rect 11265 -2905 11285 -2885
rect 11305 -2905 11310 -2885
rect 11240 -2935 11310 -2905
rect 11240 -2955 11245 -2935
rect 11265 -2955 11285 -2935
rect 11305 -2955 11310 -2935
rect 11240 -2985 11310 -2955
rect 11240 -3005 11245 -2985
rect 11265 -3005 11285 -2985
rect 11305 -3005 11310 -2985
rect 11240 -3015 11310 -3005
rect 11335 -2885 11365 -2875
rect 11335 -2905 11340 -2885
rect 11360 -2905 11365 -2885
rect 11335 -2935 11365 -2905
rect 11335 -2955 11340 -2935
rect 11360 -2955 11365 -2935
rect 11335 -2985 11365 -2955
rect 11335 -3005 11340 -2985
rect 11360 -3005 11365 -2985
rect 11335 -3015 11365 -3005
rect 11390 -2885 11420 -2875
rect 11390 -2905 11395 -2885
rect 11415 -2905 11420 -2885
rect 11390 -2935 11420 -2905
rect 11390 -2955 11395 -2935
rect 11415 -2955 11420 -2935
rect 11390 -2985 11420 -2955
rect 11390 -3005 11395 -2985
rect 11415 -3005 11420 -2985
rect 11390 -3015 11420 -3005
rect 11445 -2885 11475 -2875
rect 11445 -2905 11450 -2885
rect 11470 -2905 11475 -2885
rect 11445 -2935 11475 -2905
rect 11445 -2955 11450 -2935
rect 11470 -2955 11475 -2935
rect 11445 -2985 11475 -2955
rect 11445 -3005 11450 -2985
rect 11470 -3005 11475 -2985
rect 11445 -3015 11475 -3005
rect 11500 -2885 11530 -2875
rect 11500 -2905 11505 -2885
rect 11525 -2905 11530 -2885
rect 11500 -2935 11530 -2905
rect 11500 -2955 11505 -2935
rect 11525 -2955 11530 -2935
rect 11500 -2985 11530 -2955
rect 11500 -3005 11505 -2985
rect 11525 -3005 11530 -2985
rect 11500 -3015 11530 -3005
rect 11555 -2885 11585 -2875
rect 11555 -2905 11560 -2885
rect 11580 -2905 11585 -2885
rect 11555 -2935 11585 -2905
rect 11555 -2955 11560 -2935
rect 11580 -2955 11585 -2935
rect 11555 -2985 11585 -2955
rect 11555 -3005 11560 -2985
rect 11580 -3005 11585 -2985
rect 11555 -3015 11585 -3005
rect 11610 -2885 11640 -2875
rect 11610 -2905 11615 -2885
rect 11635 -2905 11640 -2885
rect 11610 -2935 11640 -2905
rect 11610 -2955 11615 -2935
rect 11635 -2955 11640 -2935
rect 11610 -2985 11640 -2955
rect 11610 -3005 11615 -2985
rect 11635 -3005 11640 -2985
rect 11610 -3015 11640 -3005
rect 11665 -2885 11695 -2875
rect 11665 -2905 11670 -2885
rect 11690 -2905 11695 -2885
rect 11665 -2935 11695 -2905
rect 11665 -2955 11670 -2935
rect 11690 -2955 11695 -2935
rect 11665 -2985 11695 -2955
rect 11665 -3005 11670 -2985
rect 11690 -3005 11695 -2985
rect 11665 -3015 11695 -3005
rect 11720 -2885 11750 -2875
rect 11720 -2905 11725 -2885
rect 11745 -2905 11750 -2885
rect 11720 -2935 11750 -2905
rect 11720 -2955 11725 -2935
rect 11745 -2955 11750 -2935
rect 11720 -2985 11750 -2955
rect 11720 -3005 11725 -2985
rect 11745 -3005 11750 -2985
rect 11720 -3015 11750 -3005
rect 11775 -2885 11805 -2875
rect 11775 -2905 11780 -2885
rect 11800 -2905 11805 -2885
rect 11775 -2935 11805 -2905
rect 11775 -2955 11780 -2935
rect 11800 -2955 11805 -2935
rect 11775 -2985 11805 -2955
rect 11775 -3005 11780 -2985
rect 11800 -3005 11805 -2985
rect 11775 -3015 11805 -3005
rect 11830 -2885 11860 -2875
rect 11830 -2905 11835 -2885
rect 11855 -2905 11860 -2885
rect 11830 -2935 11860 -2905
rect 11830 -2955 11835 -2935
rect 11855 -2955 11860 -2935
rect 11830 -2985 11860 -2955
rect 11830 -3005 11835 -2985
rect 11855 -3005 11860 -2985
rect 11830 -3015 11860 -3005
rect 11885 -2885 11915 -2875
rect 11885 -2905 11890 -2885
rect 11910 -2905 11915 -2885
rect 11885 -2935 11915 -2905
rect 11885 -2955 11890 -2935
rect 11910 -2955 11915 -2935
rect 11885 -2985 11915 -2955
rect 11885 -3005 11890 -2985
rect 11910 -3005 11915 -2985
rect 11885 -3015 11915 -3005
rect 11940 -2885 11970 -2875
rect 11940 -2905 11945 -2885
rect 11965 -2905 11970 -2885
rect 11940 -2935 11970 -2905
rect 11940 -2955 11945 -2935
rect 11965 -2955 11970 -2935
rect 11940 -2985 11970 -2955
rect 11940 -3005 11945 -2985
rect 11965 -3005 11970 -2985
rect 11940 -3015 11970 -3005
rect 11995 -2885 12025 -2875
rect 11995 -2905 12000 -2885
rect 12020 -2905 12025 -2885
rect 11995 -2935 12025 -2905
rect 11995 -2955 12000 -2935
rect 12020 -2955 12025 -2935
rect 11995 -2985 12025 -2955
rect 11995 -3005 12000 -2985
rect 12020 -3005 12025 -2985
rect 11995 -3015 12025 -3005
rect 12050 -2885 12080 -2875
rect 12050 -2905 12055 -2885
rect 12075 -2905 12080 -2885
rect 12050 -2935 12080 -2905
rect 12050 -2955 12055 -2935
rect 12075 -2955 12080 -2935
rect 12050 -2985 12080 -2955
rect 12050 -3005 12055 -2985
rect 12075 -3005 12080 -2985
rect 12050 -3015 12080 -3005
rect 12105 -2885 12135 -2875
rect 12105 -2905 12110 -2885
rect 12130 -2905 12135 -2885
rect 12105 -2935 12135 -2905
rect 12105 -2955 12110 -2935
rect 12130 -2955 12135 -2935
rect 12105 -2985 12135 -2955
rect 12105 -3005 12110 -2985
rect 12130 -3005 12135 -2985
rect 12105 -3015 12135 -3005
rect 12160 -2885 12190 -2875
rect 12160 -2905 12165 -2885
rect 12185 -2905 12190 -2885
rect 12160 -2935 12190 -2905
rect 12160 -2955 12165 -2935
rect 12185 -2955 12190 -2935
rect 12160 -2985 12190 -2955
rect 12160 -3005 12165 -2985
rect 12185 -3005 12190 -2985
rect 12160 -3015 12190 -3005
rect 12215 -2885 12245 -2875
rect 12215 -2905 12220 -2885
rect 12240 -2905 12245 -2885
rect 12215 -2935 12245 -2905
rect 12215 -2955 12220 -2935
rect 12240 -2955 12245 -2935
rect 12215 -2985 12245 -2955
rect 12215 -3005 12220 -2985
rect 12240 -3005 12245 -2985
rect 12215 -3015 12245 -3005
rect 12270 -2885 12300 -2875
rect 12270 -2905 12275 -2885
rect 12295 -2905 12300 -2885
rect 12270 -2935 12300 -2905
rect 12270 -2955 12275 -2935
rect 12295 -2955 12300 -2935
rect 12270 -2985 12300 -2955
rect 12270 -3005 12275 -2985
rect 12295 -3005 12300 -2985
rect 12270 -3015 12300 -3005
rect 12325 -2885 12355 -2875
rect 12325 -2905 12330 -2885
rect 12350 -2905 12355 -2885
rect 12325 -2935 12355 -2905
rect 12325 -2955 12330 -2935
rect 12350 -2955 12355 -2935
rect 12325 -2985 12355 -2955
rect 12325 -3005 12330 -2985
rect 12350 -3005 12355 -2985
rect 12325 -3015 12355 -3005
rect 12380 -2885 12410 -2875
rect 12380 -2905 12385 -2885
rect 12405 -2905 12410 -2885
rect 12380 -2935 12410 -2905
rect 12380 -2955 12385 -2935
rect 12405 -2955 12410 -2935
rect 12380 -2985 12410 -2955
rect 12380 -3005 12385 -2985
rect 12405 -3005 12410 -2985
rect 12380 -3015 12410 -3005
rect 12435 -2885 12465 -2875
rect 12435 -2905 12440 -2885
rect 12460 -2905 12465 -2885
rect 12435 -2935 12465 -2905
rect 12435 -2955 12440 -2935
rect 12460 -2955 12465 -2935
rect 12435 -2985 12465 -2955
rect 12435 -3005 12440 -2985
rect 12460 -3005 12465 -2985
rect 12435 -3015 12465 -3005
rect 12490 -2885 12560 -2875
rect 12860 -2880 12930 -2870
rect 12955 -2750 12985 -2740
rect 12955 -2770 12960 -2750
rect 12980 -2770 12985 -2750
rect 12955 -2800 12985 -2770
rect 12955 -2820 12960 -2800
rect 12980 -2820 12985 -2800
rect 12955 -2850 12985 -2820
rect 12955 -2870 12960 -2850
rect 12980 -2870 12985 -2850
rect 12955 -2880 12985 -2870
rect 13010 -2750 13040 -2740
rect 13010 -2770 13015 -2750
rect 13035 -2770 13040 -2750
rect 13010 -2800 13040 -2770
rect 13010 -2820 13015 -2800
rect 13035 -2820 13040 -2800
rect 13010 -2850 13040 -2820
rect 13010 -2870 13015 -2850
rect 13035 -2870 13040 -2850
rect 13010 -2880 13040 -2870
rect 13065 -2750 13095 -2740
rect 13065 -2770 13070 -2750
rect 13090 -2770 13095 -2750
rect 13065 -2800 13095 -2770
rect 13065 -2820 13070 -2800
rect 13090 -2820 13095 -2800
rect 13065 -2850 13095 -2820
rect 13065 -2870 13070 -2850
rect 13090 -2870 13095 -2850
rect 13065 -2880 13095 -2870
rect 13120 -2750 13150 -2740
rect 13120 -2770 13125 -2750
rect 13145 -2770 13150 -2750
rect 13120 -2800 13150 -2770
rect 13120 -2820 13125 -2800
rect 13145 -2820 13150 -2800
rect 13120 -2850 13150 -2820
rect 13120 -2870 13125 -2850
rect 13145 -2870 13150 -2850
rect 13120 -2880 13150 -2870
rect 13175 -2750 13205 -2740
rect 13175 -2770 13180 -2750
rect 13200 -2770 13205 -2750
rect 13175 -2800 13205 -2770
rect 13175 -2820 13180 -2800
rect 13200 -2820 13205 -2800
rect 13175 -2850 13205 -2820
rect 13175 -2870 13180 -2850
rect 13200 -2870 13205 -2850
rect 13175 -2880 13205 -2870
rect 13230 -2750 13260 -2740
rect 13230 -2770 13235 -2750
rect 13255 -2770 13260 -2750
rect 13230 -2800 13260 -2770
rect 13230 -2820 13235 -2800
rect 13255 -2820 13260 -2800
rect 13230 -2850 13260 -2820
rect 13230 -2870 13235 -2850
rect 13255 -2870 13260 -2850
rect 13230 -2880 13260 -2870
rect 13285 -2750 13315 -2740
rect 13285 -2770 13290 -2750
rect 13310 -2770 13315 -2750
rect 13285 -2800 13315 -2770
rect 13285 -2820 13290 -2800
rect 13310 -2820 13315 -2800
rect 13285 -2850 13315 -2820
rect 13285 -2870 13290 -2850
rect 13310 -2870 13315 -2850
rect 13285 -2880 13315 -2870
rect 13340 -2750 13370 -2740
rect 13340 -2770 13345 -2750
rect 13365 -2770 13370 -2750
rect 13340 -2800 13370 -2770
rect 13340 -2820 13345 -2800
rect 13365 -2820 13370 -2800
rect 13340 -2850 13370 -2820
rect 13340 -2870 13345 -2850
rect 13365 -2870 13370 -2850
rect 13340 -2880 13370 -2870
rect 13395 -2750 13425 -2740
rect 13395 -2770 13400 -2750
rect 13420 -2770 13425 -2750
rect 13395 -2800 13425 -2770
rect 13395 -2820 13400 -2800
rect 13420 -2820 13425 -2800
rect 13395 -2850 13425 -2820
rect 13395 -2870 13400 -2850
rect 13420 -2870 13425 -2850
rect 13395 -2880 13425 -2870
rect 13450 -2750 13480 -2740
rect 13450 -2770 13455 -2750
rect 13475 -2770 13480 -2750
rect 13450 -2800 13480 -2770
rect 13450 -2820 13455 -2800
rect 13475 -2820 13480 -2800
rect 13450 -2850 13480 -2820
rect 13450 -2870 13455 -2850
rect 13475 -2870 13480 -2850
rect 13450 -2880 13480 -2870
rect 13505 -2750 13535 -2740
rect 13505 -2770 13510 -2750
rect 13530 -2770 13535 -2750
rect 13505 -2800 13535 -2770
rect 13505 -2820 13510 -2800
rect 13530 -2820 13535 -2800
rect 13505 -2850 13535 -2820
rect 13505 -2870 13510 -2850
rect 13530 -2870 13535 -2850
rect 13505 -2880 13535 -2870
rect 13560 -2750 13590 -2740
rect 13560 -2770 13565 -2750
rect 13585 -2770 13590 -2750
rect 13560 -2800 13590 -2770
rect 13560 -2820 13565 -2800
rect 13585 -2820 13590 -2800
rect 13560 -2850 13590 -2820
rect 13560 -2870 13565 -2850
rect 13585 -2870 13590 -2850
rect 13560 -2880 13590 -2870
rect 13615 -2750 13645 -2740
rect 13615 -2770 13620 -2750
rect 13640 -2770 13645 -2750
rect 13615 -2800 13645 -2770
rect 13615 -2820 13620 -2800
rect 13640 -2820 13645 -2800
rect 13615 -2850 13645 -2820
rect 13615 -2870 13620 -2850
rect 13640 -2870 13645 -2850
rect 13615 -2880 13645 -2870
rect 13670 -2750 13700 -2740
rect 13670 -2770 13675 -2750
rect 13695 -2770 13700 -2750
rect 13670 -2800 13700 -2770
rect 13670 -2820 13675 -2800
rect 13695 -2820 13700 -2800
rect 13670 -2850 13700 -2820
rect 13670 -2870 13675 -2850
rect 13695 -2870 13700 -2850
rect 13670 -2880 13700 -2870
rect 13725 -2750 13755 -2740
rect 13725 -2770 13730 -2750
rect 13750 -2770 13755 -2750
rect 13725 -2800 13755 -2770
rect 13725 -2820 13730 -2800
rect 13750 -2820 13755 -2800
rect 13725 -2850 13755 -2820
rect 13725 -2870 13730 -2850
rect 13750 -2870 13755 -2850
rect 13725 -2880 13755 -2870
rect 13780 -2750 13810 -2740
rect 13780 -2770 13785 -2750
rect 13805 -2770 13810 -2750
rect 13780 -2800 13810 -2770
rect 13780 -2820 13785 -2800
rect 13805 -2820 13810 -2800
rect 13780 -2850 13810 -2820
rect 13780 -2870 13785 -2850
rect 13805 -2870 13810 -2850
rect 13780 -2880 13810 -2870
rect 13835 -2750 13865 -2740
rect 13835 -2770 13840 -2750
rect 13860 -2770 13865 -2750
rect 13835 -2800 13865 -2770
rect 13835 -2820 13840 -2800
rect 13860 -2820 13865 -2800
rect 13835 -2850 13865 -2820
rect 13835 -2870 13840 -2850
rect 13860 -2870 13865 -2850
rect 13835 -2880 13865 -2870
rect 13890 -2750 13920 -2740
rect 13890 -2770 13895 -2750
rect 13915 -2770 13920 -2750
rect 13890 -2800 13920 -2770
rect 13890 -2820 13895 -2800
rect 13915 -2820 13920 -2800
rect 13890 -2850 13920 -2820
rect 13890 -2870 13895 -2850
rect 13915 -2870 13920 -2850
rect 13890 -2880 13920 -2870
rect 13945 -2750 13975 -2740
rect 13945 -2770 13950 -2750
rect 13970 -2770 13975 -2750
rect 13945 -2800 13975 -2770
rect 13945 -2820 13950 -2800
rect 13970 -2820 13975 -2800
rect 13945 -2850 13975 -2820
rect 13945 -2870 13950 -2850
rect 13970 -2870 13975 -2850
rect 13945 -2880 13975 -2870
rect 14000 -2750 14030 -2740
rect 14000 -2770 14005 -2750
rect 14025 -2770 14030 -2750
rect 14000 -2800 14030 -2770
rect 14000 -2820 14005 -2800
rect 14025 -2820 14030 -2800
rect 14000 -2850 14030 -2820
rect 14000 -2870 14005 -2850
rect 14025 -2870 14030 -2850
rect 14000 -2880 14030 -2870
rect 14055 -2750 14085 -2740
rect 14055 -2770 14060 -2750
rect 14080 -2770 14085 -2750
rect 14055 -2800 14085 -2770
rect 14055 -2820 14060 -2800
rect 14080 -2820 14085 -2800
rect 14055 -2850 14085 -2820
rect 14055 -2870 14060 -2850
rect 14080 -2870 14085 -2850
rect 14055 -2880 14085 -2870
rect 14110 -2750 14180 -2740
rect 14110 -2770 14115 -2750
rect 14135 -2770 14155 -2750
rect 14175 -2770 14180 -2750
rect 14110 -2800 14180 -2770
rect 14110 -2820 14115 -2800
rect 14135 -2820 14155 -2800
rect 14175 -2820 14180 -2800
rect 14110 -2850 14180 -2820
rect 14110 -2870 14115 -2850
rect 14135 -2870 14155 -2850
rect 14175 -2870 14180 -2850
rect 14110 -2880 14180 -2870
rect 12490 -2905 12495 -2885
rect 12515 -2905 12535 -2885
rect 12555 -2905 12560 -2885
rect 12960 -2900 12980 -2880
rect 13070 -2900 13090 -2880
rect 13180 -2900 13200 -2880
rect 13290 -2900 13310 -2880
rect 13400 -2900 13420 -2880
rect 13510 -2900 13530 -2880
rect 13620 -2900 13640 -2880
rect 13730 -2900 13750 -2880
rect 13840 -2900 13860 -2880
rect 13950 -2900 13970 -2880
rect 14060 -2900 14080 -2880
rect 12490 -2935 12560 -2905
rect 12490 -2955 12495 -2935
rect 12515 -2955 12535 -2935
rect 12555 -2955 12560 -2935
rect 12950 -2910 12990 -2900
rect 12950 -2930 12962 -2910
rect 12980 -2930 12990 -2910
rect 12950 -2940 12990 -2930
rect 13060 -2910 13100 -2900
rect 13060 -2930 13072 -2910
rect 13090 -2930 13100 -2910
rect 13060 -2940 13100 -2930
rect 13170 -2910 13210 -2900
rect 13170 -2930 13182 -2910
rect 13200 -2930 13210 -2910
rect 13170 -2940 13210 -2930
rect 13280 -2910 13320 -2900
rect 13280 -2930 13292 -2910
rect 13310 -2930 13320 -2910
rect 13280 -2940 13320 -2930
rect 13390 -2910 13430 -2900
rect 13390 -2930 13402 -2910
rect 13420 -2930 13430 -2910
rect 13390 -2940 13430 -2930
rect 13500 -2910 13540 -2900
rect 13500 -2930 13512 -2910
rect 13530 -2930 13540 -2910
rect 13500 -2940 13540 -2930
rect 13610 -2910 13650 -2900
rect 13610 -2930 13622 -2910
rect 13640 -2930 13650 -2910
rect 13610 -2940 13650 -2930
rect 13720 -2910 13760 -2900
rect 13720 -2930 13732 -2910
rect 13750 -2930 13760 -2910
rect 13720 -2940 13760 -2930
rect 13830 -2910 13870 -2900
rect 13830 -2930 13842 -2910
rect 13860 -2930 13870 -2910
rect 13830 -2940 13870 -2930
rect 13940 -2910 13980 -2900
rect 13940 -2930 13952 -2910
rect 13970 -2930 13980 -2910
rect 13940 -2940 13980 -2930
rect 14050 -2910 14090 -2900
rect 14050 -2930 14062 -2910
rect 14080 -2930 14090 -2910
rect 14050 -2940 14090 -2930
rect 12490 -2985 12560 -2955
rect 12490 -3005 12495 -2985
rect 12515 -3005 12535 -2985
rect 12555 -3005 12560 -2985
rect 12995 -2970 13035 -2960
rect 12995 -2990 13005 -2970
rect 13025 -2990 13035 -2970
rect 12995 -3000 13035 -2990
rect 13098 -2970 13132 -2960
rect 13098 -2990 13106 -2970
rect 13124 -2990 13132 -2970
rect 13098 -3000 13132 -2990
rect 13195 -2970 13235 -2960
rect 13195 -2990 13205 -2970
rect 13225 -2990 13235 -2970
rect 13195 -3000 13235 -2990
rect 13395 -2970 13435 -2960
rect 13395 -2990 13405 -2970
rect 13425 -2990 13435 -2970
rect 13395 -3000 13435 -2990
rect 13595 -2970 13635 -2960
rect 13595 -2990 13605 -2970
rect 13625 -2990 13635 -2970
rect 13595 -3000 13635 -2990
rect 13795 -2970 13835 -2960
rect 13795 -2990 13805 -2970
rect 13825 -2990 13835 -2970
rect 13795 -3000 13835 -2990
rect 13995 -2970 14035 -2960
rect 13995 -2990 14005 -2970
rect 14025 -2990 14035 -2970
rect 13995 -3000 14035 -2990
rect 12490 -3015 12560 -3005
rect 11245 -3035 11265 -3015
rect 11395 -3035 11415 -3015
rect 11505 -3035 11525 -3015
rect 11615 -3035 11635 -3015
rect 11725 -3035 11745 -3015
rect 11835 -3035 11855 -3015
rect 11945 -3035 11965 -3015
rect 12055 -3035 12075 -3015
rect 12165 -3035 12185 -3015
rect 12275 -3035 12295 -3015
rect 12385 -3035 12405 -3015
rect 12535 -3035 12555 -3015
rect 13005 -3020 13025 -3000
rect 13205 -3020 13225 -3000
rect 13405 -3020 13425 -3000
rect 13605 -3020 13625 -3000
rect 13805 -3020 13825 -3000
rect 14005 -3020 14025 -3000
rect 12860 -3030 12930 -3020
rect 11235 -3045 11275 -3035
rect 11235 -3065 11245 -3045
rect 11265 -3065 11275 -3045
rect 11235 -3075 11275 -3065
rect 11385 -3045 11425 -3035
rect 11385 -3065 11395 -3045
rect 11415 -3065 11425 -3045
rect 11385 -3075 11425 -3065
rect 11495 -3045 11535 -3035
rect 11495 -3065 11505 -3045
rect 11525 -3065 11535 -3045
rect 11495 -3075 11535 -3065
rect 11605 -3045 11645 -3035
rect 11605 -3065 11615 -3045
rect 11635 -3065 11645 -3045
rect 11605 -3075 11645 -3065
rect 11715 -3045 11755 -3035
rect 11715 -3065 11725 -3045
rect 11745 -3065 11755 -3045
rect 11715 -3075 11755 -3065
rect 11825 -3045 11865 -3035
rect 11825 -3065 11835 -3045
rect 11855 -3065 11865 -3045
rect 11825 -3075 11865 -3065
rect 11935 -3045 11975 -3035
rect 11935 -3065 11945 -3045
rect 11965 -3065 11975 -3045
rect 11935 -3075 11975 -3065
rect 12045 -3045 12085 -3035
rect 12045 -3065 12055 -3045
rect 12075 -3065 12085 -3045
rect 12045 -3075 12085 -3065
rect 12155 -3045 12195 -3035
rect 12155 -3065 12165 -3045
rect 12185 -3065 12195 -3045
rect 12155 -3075 12195 -3065
rect 12265 -3045 12305 -3035
rect 12265 -3065 12275 -3045
rect 12295 -3065 12305 -3045
rect 12265 -3075 12305 -3065
rect 12375 -3045 12415 -3035
rect 12375 -3065 12385 -3045
rect 12405 -3065 12415 -3045
rect 12375 -3075 12415 -3065
rect 12525 -3045 12565 -3035
rect 12525 -3065 12535 -3045
rect 12555 -3065 12565 -3045
rect 12525 -3075 12565 -3065
rect 12860 -3050 12865 -3030
rect 12885 -3050 12905 -3030
rect 12925 -3050 12930 -3030
rect 12860 -3075 12930 -3050
rect 12860 -3095 12865 -3075
rect 12885 -3095 12905 -3075
rect 12925 -3095 12930 -3075
rect 12860 -3120 12930 -3095
rect 12860 -3140 12865 -3120
rect 12885 -3140 12905 -3120
rect 12925 -3140 12930 -3120
rect 12860 -3170 12930 -3140
rect 12860 -3190 12865 -3170
rect 12885 -3190 12905 -3170
rect 12925 -3190 12930 -3170
rect 12860 -3215 12930 -3190
rect 11190 -3230 11230 -3220
rect 11085 -3245 11125 -3235
rect 11085 -3265 11095 -3245
rect 11115 -3265 11125 -3245
rect 11190 -3250 11200 -3230
rect 11220 -3250 11230 -3230
rect 11410 -3230 11450 -3220
rect 11190 -3260 11230 -3250
rect 11305 -3245 11345 -3235
rect 11085 -3275 11125 -3265
rect 11095 -3340 11115 -3275
rect 11200 -3340 11220 -3260
rect 11305 -3265 11315 -3245
rect 11335 -3265 11345 -3245
rect 11410 -3250 11420 -3230
rect 11440 -3250 11450 -3230
rect 11640 -3230 11680 -3220
rect 11410 -3260 11450 -3250
rect 11525 -3245 11565 -3235
rect 11305 -3275 11345 -3265
rect 11237 -3290 11269 -3280
rect 11237 -3310 11243 -3290
rect 11260 -3310 11269 -3290
rect 11237 -3320 11269 -3310
rect 11315 -3340 11335 -3275
rect 11420 -3340 11440 -3260
rect 11525 -3265 11535 -3245
rect 11555 -3265 11565 -3245
rect 11640 -3250 11650 -3230
rect 11670 -3250 11680 -3230
rect 12230 -3230 12270 -3220
rect 11640 -3260 11680 -3250
rect 12125 -3245 12165 -3235
rect 11525 -3275 11565 -3265
rect 11457 -3290 11489 -3280
rect 11457 -3310 11463 -3290
rect 11480 -3310 11489 -3290
rect 11457 -3320 11489 -3310
rect 11535 -3340 11555 -3275
rect 11601 -3290 11633 -3280
rect 11601 -3310 11610 -3290
rect 11627 -3310 11633 -3290
rect 11601 -3320 11633 -3310
rect 11650 -3340 11670 -3260
rect 12125 -3265 12135 -3245
rect 12155 -3265 12165 -3245
rect 12230 -3250 12240 -3230
rect 12260 -3250 12270 -3230
rect 12450 -3230 12490 -3220
rect 12230 -3260 12270 -3250
rect 12345 -3245 12385 -3235
rect 12125 -3275 12165 -3265
rect 11820 -3290 11850 -3280
rect 11820 -3310 11825 -3290
rect 11845 -3310 11850 -3290
rect 11820 -3320 11850 -3310
rect 11867 -3290 11899 -3280
rect 11867 -3310 11876 -3290
rect 11893 -3310 11899 -3290
rect 11867 -3320 11899 -3310
rect 11950 -3290 11980 -3280
rect 11950 -3310 11955 -3290
rect 11975 -3310 11980 -3290
rect 11950 -3320 11980 -3310
rect 11830 -3340 11850 -3320
rect 11950 -3340 11970 -3320
rect 12135 -3340 12155 -3275
rect 12240 -3340 12260 -3260
rect 12345 -3265 12355 -3245
rect 12375 -3265 12385 -3245
rect 12450 -3250 12460 -3230
rect 12480 -3250 12490 -3230
rect 12680 -3230 12720 -3220
rect 12450 -3260 12490 -3250
rect 12565 -3245 12605 -3235
rect 12345 -3275 12385 -3265
rect 12277 -3290 12309 -3280
rect 12277 -3310 12283 -3290
rect 12300 -3310 12309 -3290
rect 12277 -3320 12309 -3310
rect 12355 -3340 12375 -3275
rect 12460 -3340 12480 -3260
rect 12565 -3265 12575 -3245
rect 12595 -3265 12605 -3245
rect 12680 -3250 12690 -3230
rect 12710 -3250 12720 -3230
rect 12680 -3260 12720 -3250
rect 12860 -3235 12865 -3215
rect 12885 -3235 12905 -3215
rect 12925 -3235 12930 -3215
rect 12860 -3260 12930 -3235
rect 12565 -3275 12605 -3265
rect 12497 -3290 12529 -3280
rect 12497 -3310 12503 -3290
rect 12520 -3310 12529 -3290
rect 12497 -3320 12529 -3310
rect 12575 -3340 12595 -3275
rect 12641 -3290 12673 -3280
rect 12641 -3310 12650 -3290
rect 12667 -3310 12673 -3290
rect 12641 -3320 12673 -3310
rect 12690 -3340 12710 -3260
rect 12860 -3280 12865 -3260
rect 12885 -3280 12905 -3260
rect 12925 -3280 12930 -3260
rect 12860 -3290 12930 -3280
rect 13000 -3030 13030 -3020
rect 13000 -3050 13005 -3030
rect 13025 -3050 13030 -3030
rect 13000 -3075 13030 -3050
rect 13000 -3095 13005 -3075
rect 13025 -3095 13030 -3075
rect 13000 -3120 13030 -3095
rect 13000 -3140 13005 -3120
rect 13025 -3140 13030 -3120
rect 13000 -3170 13030 -3140
rect 13000 -3190 13005 -3170
rect 13025 -3190 13030 -3170
rect 13000 -3215 13030 -3190
rect 13000 -3235 13005 -3215
rect 13025 -3235 13030 -3215
rect 13000 -3260 13030 -3235
rect 13000 -3280 13005 -3260
rect 13025 -3280 13030 -3260
rect 13000 -3290 13030 -3280
rect 13100 -3030 13130 -3020
rect 13100 -3050 13105 -3030
rect 13125 -3050 13130 -3030
rect 13100 -3075 13130 -3050
rect 13100 -3095 13105 -3075
rect 13125 -3095 13130 -3075
rect 13100 -3120 13130 -3095
rect 13100 -3140 13105 -3120
rect 13125 -3140 13130 -3120
rect 13100 -3170 13130 -3140
rect 13100 -3190 13105 -3170
rect 13125 -3190 13130 -3170
rect 13100 -3215 13130 -3190
rect 13100 -3235 13105 -3215
rect 13125 -3235 13130 -3215
rect 13100 -3260 13130 -3235
rect 13100 -3280 13105 -3260
rect 13125 -3280 13130 -3260
rect 13100 -3290 13130 -3280
rect 13200 -3030 13230 -3020
rect 13200 -3050 13205 -3030
rect 13225 -3050 13230 -3030
rect 13200 -3075 13230 -3050
rect 13200 -3095 13205 -3075
rect 13225 -3095 13230 -3075
rect 13200 -3120 13230 -3095
rect 13200 -3140 13205 -3120
rect 13225 -3140 13230 -3120
rect 13200 -3170 13230 -3140
rect 13200 -3190 13205 -3170
rect 13225 -3190 13230 -3170
rect 13200 -3215 13230 -3190
rect 13200 -3235 13205 -3215
rect 13225 -3235 13230 -3215
rect 13200 -3260 13230 -3235
rect 13200 -3280 13205 -3260
rect 13225 -3280 13230 -3260
rect 13200 -3290 13230 -3280
rect 13300 -3030 13330 -3020
rect 13300 -3050 13305 -3030
rect 13325 -3050 13330 -3030
rect 13300 -3075 13330 -3050
rect 13300 -3095 13305 -3075
rect 13325 -3095 13330 -3075
rect 13300 -3120 13330 -3095
rect 13300 -3140 13305 -3120
rect 13325 -3140 13330 -3120
rect 13300 -3170 13330 -3140
rect 13300 -3190 13305 -3170
rect 13325 -3190 13330 -3170
rect 13300 -3215 13330 -3190
rect 13300 -3235 13305 -3215
rect 13325 -3235 13330 -3215
rect 13300 -3260 13330 -3235
rect 13300 -3280 13305 -3260
rect 13325 -3280 13330 -3260
rect 13300 -3290 13330 -3280
rect 13400 -3030 13430 -3020
rect 13400 -3050 13405 -3030
rect 13425 -3050 13430 -3030
rect 13400 -3075 13430 -3050
rect 13400 -3095 13405 -3075
rect 13425 -3095 13430 -3075
rect 13400 -3120 13430 -3095
rect 13400 -3140 13405 -3120
rect 13425 -3140 13430 -3120
rect 13400 -3170 13430 -3140
rect 13400 -3190 13405 -3170
rect 13425 -3190 13430 -3170
rect 13400 -3215 13430 -3190
rect 13400 -3235 13405 -3215
rect 13425 -3235 13430 -3215
rect 13400 -3260 13430 -3235
rect 13400 -3280 13405 -3260
rect 13425 -3280 13430 -3260
rect 13400 -3290 13430 -3280
rect 13500 -3030 13530 -3020
rect 13500 -3050 13505 -3030
rect 13525 -3050 13530 -3030
rect 13500 -3075 13530 -3050
rect 13500 -3095 13505 -3075
rect 13525 -3095 13530 -3075
rect 13500 -3120 13530 -3095
rect 13500 -3140 13505 -3120
rect 13525 -3140 13530 -3120
rect 13500 -3170 13530 -3140
rect 13500 -3190 13505 -3170
rect 13525 -3190 13530 -3170
rect 13500 -3215 13530 -3190
rect 13500 -3235 13505 -3215
rect 13525 -3235 13530 -3215
rect 13500 -3260 13530 -3235
rect 13500 -3280 13505 -3260
rect 13525 -3280 13530 -3260
rect 13500 -3290 13530 -3280
rect 13600 -3030 13630 -3020
rect 13600 -3050 13605 -3030
rect 13625 -3050 13630 -3030
rect 13600 -3075 13630 -3050
rect 13600 -3095 13605 -3075
rect 13625 -3095 13630 -3075
rect 13600 -3120 13630 -3095
rect 13600 -3140 13605 -3120
rect 13625 -3140 13630 -3120
rect 13600 -3170 13630 -3140
rect 13600 -3190 13605 -3170
rect 13625 -3190 13630 -3170
rect 13600 -3215 13630 -3190
rect 13600 -3235 13605 -3215
rect 13625 -3235 13630 -3215
rect 13600 -3260 13630 -3235
rect 13600 -3280 13605 -3260
rect 13625 -3280 13630 -3260
rect 13600 -3290 13630 -3280
rect 13700 -3030 13730 -3020
rect 13700 -3050 13705 -3030
rect 13725 -3050 13730 -3030
rect 13700 -3075 13730 -3050
rect 13700 -3095 13705 -3075
rect 13725 -3095 13730 -3075
rect 13700 -3120 13730 -3095
rect 13700 -3140 13705 -3120
rect 13725 -3140 13730 -3120
rect 13700 -3170 13730 -3140
rect 13700 -3190 13705 -3170
rect 13725 -3190 13730 -3170
rect 13700 -3215 13730 -3190
rect 13700 -3235 13705 -3215
rect 13725 -3235 13730 -3215
rect 13700 -3260 13730 -3235
rect 13700 -3280 13705 -3260
rect 13725 -3280 13730 -3260
rect 13700 -3290 13730 -3280
rect 13800 -3030 13830 -3020
rect 13800 -3050 13805 -3030
rect 13825 -3050 13830 -3030
rect 13800 -3075 13830 -3050
rect 13800 -3095 13805 -3075
rect 13825 -3095 13830 -3075
rect 13800 -3120 13830 -3095
rect 13800 -3140 13805 -3120
rect 13825 -3140 13830 -3120
rect 13800 -3170 13830 -3140
rect 13800 -3190 13805 -3170
rect 13825 -3190 13830 -3170
rect 13800 -3215 13830 -3190
rect 13800 -3235 13805 -3215
rect 13825 -3235 13830 -3215
rect 13800 -3260 13830 -3235
rect 13800 -3280 13805 -3260
rect 13825 -3280 13830 -3260
rect 13800 -3290 13830 -3280
rect 13900 -3030 13930 -3020
rect 13900 -3050 13905 -3030
rect 13925 -3050 13930 -3030
rect 13900 -3075 13930 -3050
rect 13900 -3095 13905 -3075
rect 13925 -3095 13930 -3075
rect 13900 -3120 13930 -3095
rect 13900 -3140 13905 -3120
rect 13925 -3140 13930 -3120
rect 13900 -3170 13930 -3140
rect 13900 -3190 13905 -3170
rect 13925 -3190 13930 -3170
rect 13900 -3215 13930 -3190
rect 13900 -3235 13905 -3215
rect 13925 -3235 13930 -3215
rect 13900 -3260 13930 -3235
rect 13900 -3280 13905 -3260
rect 13925 -3280 13930 -3260
rect 13900 -3290 13930 -3280
rect 14000 -3030 14030 -3020
rect 14000 -3050 14005 -3030
rect 14025 -3050 14030 -3030
rect 14000 -3075 14030 -3050
rect 14000 -3095 14005 -3075
rect 14025 -3095 14030 -3075
rect 14000 -3120 14030 -3095
rect 14000 -3140 14005 -3120
rect 14025 -3140 14030 -3120
rect 14000 -3170 14030 -3140
rect 14000 -3190 14005 -3170
rect 14025 -3190 14030 -3170
rect 14000 -3215 14030 -3190
rect 14000 -3235 14005 -3215
rect 14025 -3235 14030 -3215
rect 14000 -3260 14030 -3235
rect 14000 -3280 14005 -3260
rect 14025 -3280 14030 -3260
rect 14000 -3290 14030 -3280
rect 14100 -3030 14170 -3020
rect 14100 -3050 14105 -3030
rect 14125 -3050 14145 -3030
rect 14165 -3050 14170 -3030
rect 14100 -3075 14170 -3050
rect 14100 -3095 14105 -3075
rect 14125 -3095 14145 -3075
rect 14165 -3095 14170 -3075
rect 14100 -3120 14170 -3095
rect 14100 -3140 14105 -3120
rect 14125 -3140 14145 -3120
rect 14165 -3140 14170 -3120
rect 14100 -3170 14170 -3140
rect 14100 -3190 14105 -3170
rect 14125 -3190 14145 -3170
rect 14165 -3190 14170 -3170
rect 14100 -3215 14170 -3190
rect 14100 -3235 14105 -3215
rect 14125 -3235 14145 -3215
rect 14165 -3235 14170 -3215
rect 14100 -3260 14170 -3235
rect 14100 -3280 14105 -3260
rect 14125 -3280 14145 -3260
rect 14165 -3280 14170 -3260
rect 14100 -3290 14170 -3280
rect 12865 -3310 12885 -3290
rect 13105 -3310 13125 -3290
rect 13305 -3310 13325 -3290
rect 13505 -3310 13525 -3290
rect 13705 -3310 13725 -3290
rect 13905 -3310 13925 -3290
rect 14145 -3310 14165 -3290
rect 12855 -3320 12895 -3310
rect 12855 -3340 12865 -3320
rect 12885 -3340 12895 -3320
rect 10990 -3350 11065 -3340
rect 10990 -3370 11000 -3350
rect 11020 -3370 11040 -3350
rect 11060 -3370 11065 -3350
rect 10990 -3400 11065 -3370
rect 10990 -3420 11000 -3400
rect 11020 -3420 11040 -3400
rect 11060 -3420 11065 -3400
rect 10990 -3450 11065 -3420
rect 10990 -3470 11000 -3450
rect 11020 -3470 11040 -3450
rect 11060 -3470 11065 -3450
rect 10990 -3480 11065 -3470
rect 11090 -3350 11120 -3340
rect 11090 -3370 11095 -3350
rect 11115 -3370 11120 -3350
rect 11090 -3400 11120 -3370
rect 11090 -3420 11095 -3400
rect 11115 -3420 11120 -3400
rect 11090 -3450 11120 -3420
rect 11090 -3470 11095 -3450
rect 11115 -3470 11120 -3450
rect 11090 -3480 11120 -3470
rect 11145 -3350 11175 -3340
rect 11145 -3370 11150 -3350
rect 11170 -3370 11175 -3350
rect 11145 -3400 11175 -3370
rect 11145 -3420 11150 -3400
rect 11170 -3420 11175 -3400
rect 11145 -3450 11175 -3420
rect 11145 -3470 11150 -3450
rect 11170 -3470 11175 -3450
rect 11145 -3480 11175 -3470
rect 11200 -3350 11230 -3340
rect 11200 -3370 11205 -3350
rect 11225 -3370 11230 -3350
rect 11200 -3400 11230 -3370
rect 11200 -3420 11205 -3400
rect 11225 -3420 11230 -3400
rect 11200 -3450 11230 -3420
rect 11200 -3470 11205 -3450
rect 11225 -3470 11230 -3450
rect 11200 -3480 11230 -3470
rect 11255 -3350 11285 -3340
rect 11255 -3370 11260 -3350
rect 11280 -3370 11285 -3350
rect 11255 -3400 11285 -3370
rect 11255 -3420 11260 -3400
rect 11280 -3420 11285 -3400
rect 11255 -3450 11285 -3420
rect 11255 -3470 11260 -3450
rect 11280 -3470 11285 -3450
rect 11255 -3480 11285 -3470
rect 11310 -3350 11340 -3340
rect 11310 -3370 11315 -3350
rect 11335 -3370 11340 -3350
rect 11310 -3400 11340 -3370
rect 11310 -3420 11315 -3400
rect 11335 -3420 11340 -3400
rect 11310 -3450 11340 -3420
rect 11310 -3470 11315 -3450
rect 11335 -3470 11340 -3450
rect 11310 -3480 11340 -3470
rect 11365 -3350 11395 -3340
rect 11365 -3370 11370 -3350
rect 11390 -3370 11395 -3350
rect 11365 -3400 11395 -3370
rect 11365 -3420 11370 -3400
rect 11390 -3420 11395 -3400
rect 11365 -3450 11395 -3420
rect 11365 -3470 11370 -3450
rect 11390 -3470 11395 -3450
rect 11365 -3480 11395 -3470
rect 11420 -3350 11450 -3340
rect 11420 -3370 11425 -3350
rect 11445 -3370 11450 -3350
rect 11420 -3400 11450 -3370
rect 11420 -3420 11425 -3400
rect 11445 -3420 11450 -3400
rect 11420 -3450 11450 -3420
rect 11420 -3470 11425 -3450
rect 11445 -3470 11450 -3450
rect 11420 -3480 11450 -3470
rect 11475 -3350 11505 -3340
rect 11475 -3370 11480 -3350
rect 11500 -3370 11505 -3350
rect 11475 -3400 11505 -3370
rect 11475 -3420 11480 -3400
rect 11500 -3420 11505 -3400
rect 11475 -3450 11505 -3420
rect 11475 -3470 11480 -3450
rect 11500 -3470 11505 -3450
rect 11475 -3480 11505 -3470
rect 11530 -3350 11560 -3340
rect 11530 -3370 11535 -3350
rect 11555 -3370 11560 -3350
rect 11530 -3400 11560 -3370
rect 11530 -3420 11535 -3400
rect 11555 -3420 11560 -3400
rect 11530 -3450 11560 -3420
rect 11530 -3470 11535 -3450
rect 11555 -3470 11560 -3450
rect 11530 -3480 11560 -3470
rect 11585 -3350 11615 -3340
rect 11585 -3370 11590 -3350
rect 11610 -3370 11615 -3350
rect 11585 -3400 11615 -3370
rect 11585 -3420 11590 -3400
rect 11610 -3420 11615 -3400
rect 11585 -3450 11615 -3420
rect 11585 -3470 11590 -3450
rect 11610 -3470 11615 -3450
rect 11585 -3480 11615 -3470
rect 11640 -3350 11670 -3340
rect 11640 -3370 11645 -3350
rect 11665 -3370 11670 -3350
rect 11640 -3400 11670 -3370
rect 11640 -3420 11645 -3400
rect 11665 -3420 11670 -3400
rect 11640 -3450 11670 -3420
rect 11640 -3470 11645 -3450
rect 11665 -3470 11670 -3450
rect 11640 -3480 11670 -3470
rect 11695 -3350 11805 -3340
rect 11695 -3370 11700 -3350
rect 11720 -3370 11740 -3350
rect 11760 -3370 11780 -3350
rect 11800 -3370 11805 -3350
rect 11695 -3400 11805 -3370
rect 11695 -3420 11700 -3400
rect 11720 -3420 11740 -3400
rect 11760 -3420 11780 -3400
rect 11800 -3420 11805 -3400
rect 11695 -3450 11805 -3420
rect 11695 -3470 11700 -3450
rect 11720 -3470 11740 -3450
rect 11760 -3470 11780 -3450
rect 11800 -3470 11805 -3450
rect 11695 -3480 11805 -3470
rect 11830 -3350 11860 -3340
rect 11830 -3370 11835 -3350
rect 11855 -3370 11860 -3350
rect 11830 -3400 11860 -3370
rect 11830 -3420 11835 -3400
rect 11855 -3420 11860 -3400
rect 11830 -3450 11860 -3420
rect 11830 -3470 11835 -3450
rect 11855 -3470 11860 -3450
rect 11830 -3480 11860 -3470
rect 11885 -3350 11915 -3340
rect 11885 -3370 11890 -3350
rect 11910 -3370 11915 -3350
rect 11885 -3400 11915 -3370
rect 11885 -3420 11890 -3400
rect 11910 -3420 11915 -3400
rect 11885 -3450 11915 -3420
rect 11885 -3470 11890 -3450
rect 11910 -3470 11915 -3450
rect 11885 -3480 11915 -3470
rect 11940 -3350 11970 -3340
rect 11940 -3370 11945 -3350
rect 11965 -3370 11970 -3350
rect 11940 -3400 11970 -3370
rect 11940 -3420 11945 -3400
rect 11965 -3420 11970 -3400
rect 11940 -3450 11970 -3420
rect 11940 -3470 11945 -3450
rect 11965 -3470 11970 -3450
rect 11940 -3480 11970 -3470
rect 11995 -3350 12105 -3340
rect 11995 -3370 12000 -3350
rect 12020 -3370 12040 -3350
rect 12060 -3370 12080 -3350
rect 12100 -3370 12105 -3350
rect 11995 -3400 12105 -3370
rect 11995 -3420 12000 -3400
rect 12020 -3420 12040 -3400
rect 12060 -3420 12080 -3400
rect 12100 -3420 12105 -3400
rect 11995 -3450 12105 -3420
rect 11995 -3470 12000 -3450
rect 12020 -3470 12040 -3450
rect 12060 -3470 12080 -3450
rect 12100 -3470 12105 -3450
rect 11995 -3480 12105 -3470
rect 12130 -3350 12160 -3340
rect 12130 -3370 12135 -3350
rect 12155 -3370 12160 -3350
rect 12130 -3400 12160 -3370
rect 12130 -3420 12135 -3400
rect 12155 -3420 12160 -3400
rect 12130 -3450 12160 -3420
rect 12130 -3470 12135 -3450
rect 12155 -3470 12160 -3450
rect 12130 -3480 12160 -3470
rect 12185 -3350 12215 -3340
rect 12185 -3370 12190 -3350
rect 12210 -3370 12215 -3350
rect 12185 -3400 12215 -3370
rect 12185 -3420 12190 -3400
rect 12210 -3420 12215 -3400
rect 12185 -3450 12215 -3420
rect 12185 -3470 12190 -3450
rect 12210 -3470 12215 -3450
rect 12185 -3480 12215 -3470
rect 12240 -3350 12270 -3340
rect 12240 -3370 12245 -3350
rect 12265 -3370 12270 -3350
rect 12240 -3400 12270 -3370
rect 12240 -3420 12245 -3400
rect 12265 -3420 12270 -3400
rect 12240 -3450 12270 -3420
rect 12240 -3470 12245 -3450
rect 12265 -3470 12270 -3450
rect 12240 -3480 12270 -3470
rect 12295 -3350 12325 -3340
rect 12295 -3370 12300 -3350
rect 12320 -3370 12325 -3350
rect 12295 -3400 12325 -3370
rect 12295 -3420 12300 -3400
rect 12320 -3420 12325 -3400
rect 12295 -3450 12325 -3420
rect 12295 -3470 12300 -3450
rect 12320 -3470 12325 -3450
rect 12295 -3480 12325 -3470
rect 12350 -3350 12380 -3340
rect 12350 -3370 12355 -3350
rect 12375 -3370 12380 -3350
rect 12350 -3400 12380 -3370
rect 12350 -3420 12355 -3400
rect 12375 -3420 12380 -3400
rect 12350 -3450 12380 -3420
rect 12350 -3470 12355 -3450
rect 12375 -3470 12380 -3450
rect 12350 -3480 12380 -3470
rect 12405 -3350 12435 -3340
rect 12405 -3370 12410 -3350
rect 12430 -3370 12435 -3350
rect 12405 -3400 12435 -3370
rect 12405 -3420 12410 -3400
rect 12430 -3420 12435 -3400
rect 12405 -3450 12435 -3420
rect 12405 -3470 12410 -3450
rect 12430 -3470 12435 -3450
rect 12405 -3480 12435 -3470
rect 12460 -3350 12490 -3340
rect 12460 -3370 12465 -3350
rect 12485 -3370 12490 -3350
rect 12460 -3400 12490 -3370
rect 12460 -3420 12465 -3400
rect 12485 -3420 12490 -3400
rect 12460 -3450 12490 -3420
rect 12460 -3470 12465 -3450
rect 12485 -3470 12490 -3450
rect 12460 -3480 12490 -3470
rect 12515 -3350 12545 -3340
rect 12515 -3370 12520 -3350
rect 12540 -3370 12545 -3350
rect 12515 -3400 12545 -3370
rect 12515 -3420 12520 -3400
rect 12540 -3420 12545 -3400
rect 12515 -3450 12545 -3420
rect 12515 -3470 12520 -3450
rect 12540 -3470 12545 -3450
rect 12515 -3480 12545 -3470
rect 12570 -3350 12600 -3340
rect 12570 -3370 12575 -3350
rect 12595 -3370 12600 -3350
rect 12570 -3400 12600 -3370
rect 12570 -3420 12575 -3400
rect 12595 -3420 12600 -3400
rect 12570 -3450 12600 -3420
rect 12570 -3470 12575 -3450
rect 12595 -3470 12600 -3450
rect 12570 -3480 12600 -3470
rect 12625 -3350 12655 -3340
rect 12625 -3370 12630 -3350
rect 12650 -3370 12655 -3350
rect 12625 -3400 12655 -3370
rect 12625 -3420 12630 -3400
rect 12650 -3420 12655 -3400
rect 12625 -3450 12655 -3420
rect 12625 -3470 12630 -3450
rect 12650 -3470 12655 -3450
rect 12625 -3480 12655 -3470
rect 12680 -3350 12710 -3340
rect 12680 -3370 12685 -3350
rect 12705 -3370 12710 -3350
rect 12680 -3400 12710 -3370
rect 12680 -3420 12685 -3400
rect 12705 -3420 12710 -3400
rect 12680 -3450 12710 -3420
rect 12680 -3470 12685 -3450
rect 12705 -3470 12710 -3450
rect 12680 -3480 12710 -3470
rect 12735 -3350 12810 -3340
rect 12855 -3350 12895 -3340
rect 13095 -3320 13135 -3310
rect 13095 -3340 13105 -3320
rect 13125 -3340 13135 -3320
rect 13095 -3350 13135 -3340
rect 13295 -3320 13335 -3310
rect 13295 -3340 13305 -3320
rect 13325 -3340 13335 -3320
rect 13295 -3350 13335 -3340
rect 13495 -3320 13535 -3310
rect 13495 -3340 13505 -3320
rect 13525 -3340 13535 -3320
rect 13495 -3350 13535 -3340
rect 13695 -3320 13735 -3310
rect 13695 -3340 13705 -3320
rect 13725 -3340 13735 -3320
rect 13695 -3350 13735 -3340
rect 13895 -3320 13935 -3310
rect 13895 -3340 13905 -3320
rect 13925 -3340 13935 -3320
rect 13895 -3350 13935 -3340
rect 14135 -3320 14175 -3310
rect 14135 -3340 14145 -3320
rect 14165 -3340 14175 -3320
rect 14135 -3350 14175 -3340
rect 12735 -3370 12740 -3350
rect 12760 -3370 12780 -3350
rect 12800 -3370 12810 -3350
rect 12735 -3400 12810 -3370
rect 12735 -3420 12740 -3400
rect 12760 -3420 12780 -3400
rect 12800 -3420 12810 -3400
rect 12735 -3450 12810 -3420
rect 12735 -3470 12740 -3450
rect 12760 -3470 12780 -3450
rect 12800 -3470 12810 -3450
rect 12735 -3480 12810 -3470
rect 11000 -3500 11020 -3480
rect 10990 -3510 11030 -3500
rect 10990 -3530 11000 -3510
rect 11020 -3530 11030 -3510
rect 10990 -3540 11030 -3530
rect 11106 -3510 11138 -3500
rect 11106 -3530 11112 -3510
rect 11129 -3530 11138 -3510
rect 11106 -3540 11138 -3530
rect 11155 -3560 11175 -3480
rect 11260 -3560 11280 -3480
rect 11305 -3510 11345 -3500
rect 11305 -3530 11315 -3510
rect 11335 -3530 11345 -3510
rect 11305 -3540 11345 -3530
rect 11370 -3560 11390 -3480
rect 11480 -3560 11500 -3480
rect 11525 -3510 11565 -3500
rect 11525 -3530 11535 -3510
rect 11555 -3530 11565 -3510
rect 11525 -3540 11565 -3530
rect 11590 -3560 11610 -3480
rect 11740 -3500 11760 -3480
rect 11830 -3500 11850 -3480
rect 11885 -3500 11905 -3480
rect 12040 -3500 12060 -3480
rect 11730 -3510 11770 -3500
rect 11730 -3530 11740 -3510
rect 11760 -3530 11770 -3510
rect 11730 -3540 11770 -3530
rect 11825 -3510 11855 -3500
rect 11825 -3530 11830 -3510
rect 11850 -3530 11855 -3510
rect 11825 -3540 11855 -3530
rect 11875 -3510 11905 -3500
rect 11875 -3530 11880 -3510
rect 11900 -3530 11905 -3510
rect 11875 -3540 11905 -3530
rect 11922 -3510 11954 -3500
rect 11922 -3530 11928 -3510
rect 11945 -3530 11954 -3510
rect 11922 -3540 11954 -3530
rect 12030 -3510 12070 -3500
rect 12030 -3530 12040 -3510
rect 12060 -3530 12070 -3510
rect 12030 -3540 12070 -3530
rect 12146 -3510 12178 -3500
rect 12146 -3530 12152 -3510
rect 12169 -3530 12178 -3510
rect 12146 -3540 12178 -3530
rect 12195 -3560 12215 -3480
rect 12300 -3560 12320 -3480
rect 12345 -3510 12385 -3500
rect 12345 -3530 12355 -3510
rect 12375 -3530 12385 -3510
rect 12345 -3540 12385 -3530
rect 12410 -3560 12430 -3480
rect 12520 -3560 12540 -3480
rect 12565 -3510 12605 -3500
rect 12565 -3530 12575 -3510
rect 12595 -3530 12605 -3510
rect 12565 -3540 12605 -3530
rect 12630 -3560 12650 -3480
rect 12780 -3500 12800 -3480
rect 12770 -3510 12810 -3500
rect 12770 -3530 12780 -3510
rect 12800 -3530 12810 -3510
rect 12770 -3540 12810 -3530
rect 11145 -3570 11185 -3560
rect 11145 -3590 11155 -3570
rect 11175 -3590 11185 -3570
rect 11145 -3600 11185 -3590
rect 11250 -3570 11290 -3560
rect 11250 -3590 11260 -3570
rect 11280 -3590 11290 -3570
rect 11250 -3600 11290 -3590
rect 11360 -3570 11400 -3560
rect 11360 -3590 11370 -3570
rect 11390 -3590 11400 -3570
rect 11360 -3600 11400 -3590
rect 11470 -3570 11510 -3560
rect 11470 -3590 11480 -3570
rect 11500 -3590 11510 -3570
rect 11470 -3600 11510 -3590
rect 11580 -3570 11620 -3560
rect 11580 -3590 11590 -3570
rect 11610 -3590 11620 -3570
rect 11580 -3600 11620 -3590
rect 12185 -3570 12225 -3560
rect 12185 -3590 12195 -3570
rect 12215 -3590 12225 -3570
rect 12185 -3600 12225 -3590
rect 12290 -3570 12330 -3560
rect 12290 -3590 12300 -3570
rect 12320 -3590 12330 -3570
rect 12290 -3600 12330 -3590
rect 12400 -3570 12440 -3560
rect 12400 -3590 12410 -3570
rect 12430 -3590 12440 -3570
rect 12400 -3600 12440 -3590
rect 12510 -3570 12550 -3560
rect 12510 -3590 12520 -3570
rect 12540 -3590 12550 -3570
rect 12510 -3600 12550 -3590
rect 12620 -3570 12660 -3560
rect 12620 -3590 12630 -3570
rect 12650 -3590 12660 -3570
rect 12620 -3600 12660 -3590
rect 11810 -3690 11850 -3650
rect 11315 -3740 11355 -3700
rect 11880 -3740 11920 -3700
rect 12595 -3755 12635 -3745
rect 11315 -3770 11355 -3760
rect 11315 -3790 11325 -3770
rect 11345 -3790 11355 -3770
rect 11315 -3800 11355 -3790
rect 11425 -3770 11465 -3760
rect 11425 -3790 11435 -3770
rect 11455 -3790 11465 -3770
rect 11425 -3800 11465 -3790
rect 11535 -3770 11575 -3760
rect 11535 -3790 11545 -3770
rect 11565 -3790 11575 -3770
rect 11535 -3800 11575 -3790
rect 11645 -3770 11685 -3760
rect 11645 -3790 11655 -3770
rect 11675 -3790 11685 -3770
rect 11645 -3800 11685 -3790
rect 11755 -3770 11795 -3760
rect 11755 -3790 11765 -3770
rect 11785 -3790 11795 -3770
rect 11755 -3800 11795 -3790
rect 11815 -3770 11845 -3760
rect 11815 -3790 11820 -3770
rect 11840 -3790 11845 -3770
rect 11815 -3800 11845 -3790
rect 11865 -3770 11905 -3760
rect 11865 -3790 11875 -3770
rect 11895 -3790 11905 -3770
rect 11865 -3800 11905 -3790
rect 11975 -3770 12015 -3760
rect 11975 -3790 11985 -3770
rect 12005 -3790 12015 -3770
rect 11975 -3800 12015 -3790
rect 12085 -3770 12125 -3760
rect 12085 -3790 12095 -3770
rect 12115 -3790 12125 -3770
rect 12085 -3800 12125 -3790
rect 12195 -3770 12235 -3760
rect 12195 -3790 12205 -3770
rect 12225 -3790 12235 -3770
rect 12195 -3800 12235 -3790
rect 12305 -3770 12345 -3760
rect 12305 -3790 12315 -3770
rect 12335 -3790 12345 -3770
rect 12305 -3800 12345 -3790
rect 12415 -3770 12455 -3760
rect 12415 -3790 12425 -3770
rect 12445 -3790 12455 -3770
rect 12415 -3800 12455 -3790
rect 12525 -3770 12565 -3760
rect 12525 -3790 12535 -3770
rect 12555 -3790 12565 -3770
rect 12595 -3775 12605 -3755
rect 12625 -3775 12635 -3755
rect 12595 -3785 12635 -3775
rect 12525 -3800 12565 -3790
rect 11325 -3820 11345 -3800
rect 11435 -3820 11455 -3800
rect 11545 -3820 11565 -3800
rect 11655 -3820 11675 -3800
rect 11765 -3820 11785 -3800
rect 11875 -3820 11895 -3800
rect 11985 -3820 12005 -3800
rect 12095 -3820 12115 -3800
rect 12205 -3820 12225 -3800
rect 12315 -3820 12335 -3800
rect 12425 -3820 12445 -3800
rect 12535 -3820 12555 -3800
rect 11170 -3830 11240 -3820
rect 11170 -3850 11175 -3830
rect 11195 -3850 11215 -3830
rect 11235 -3850 11240 -3830
rect 11170 -3880 11240 -3850
rect 11170 -3900 11175 -3880
rect 11195 -3900 11215 -3880
rect 11235 -3900 11240 -3880
rect 11170 -3930 11240 -3900
rect 11170 -3950 11175 -3930
rect 11195 -3950 11215 -3930
rect 11235 -3950 11240 -3930
rect 11170 -3980 11240 -3950
rect 11170 -4000 11175 -3980
rect 11195 -4000 11215 -3980
rect 11235 -4000 11240 -3980
rect 11170 -4030 11240 -4000
rect 11170 -4050 11175 -4030
rect 11195 -4050 11215 -4030
rect 11235 -4050 11240 -4030
rect 11170 -4060 11240 -4050
rect 11265 -3830 11295 -3820
rect 11265 -3850 11270 -3830
rect 11290 -3850 11295 -3830
rect 11265 -3880 11295 -3850
rect 11265 -3900 11270 -3880
rect 11290 -3900 11295 -3880
rect 11265 -3930 11295 -3900
rect 11265 -3950 11270 -3930
rect 11290 -3950 11295 -3930
rect 11265 -3980 11295 -3950
rect 11265 -4000 11270 -3980
rect 11290 -4000 11295 -3980
rect 11265 -4030 11295 -4000
rect 11265 -4050 11270 -4030
rect 11290 -4050 11295 -4030
rect 11265 -4060 11295 -4050
rect 11320 -3830 11350 -3820
rect 11320 -3850 11325 -3830
rect 11345 -3850 11350 -3830
rect 11320 -3880 11350 -3850
rect 11320 -3900 11325 -3880
rect 11345 -3900 11350 -3880
rect 11320 -3930 11350 -3900
rect 11320 -3950 11325 -3930
rect 11345 -3950 11350 -3930
rect 11320 -3980 11350 -3950
rect 11320 -4000 11325 -3980
rect 11345 -4000 11350 -3980
rect 11320 -4030 11350 -4000
rect 11320 -4050 11325 -4030
rect 11345 -4050 11350 -4030
rect 11320 -4060 11350 -4050
rect 11375 -3830 11405 -3820
rect 11375 -3850 11380 -3830
rect 11400 -3850 11405 -3830
rect 11375 -3880 11405 -3850
rect 11375 -3900 11380 -3880
rect 11400 -3900 11405 -3880
rect 11375 -3930 11405 -3900
rect 11375 -3950 11380 -3930
rect 11400 -3950 11405 -3930
rect 11375 -3980 11405 -3950
rect 11375 -4000 11380 -3980
rect 11400 -4000 11405 -3980
rect 11375 -4030 11405 -4000
rect 11375 -4050 11380 -4030
rect 11400 -4050 11405 -4030
rect 11375 -4060 11405 -4050
rect 11430 -3830 11460 -3820
rect 11430 -3850 11435 -3830
rect 11455 -3850 11460 -3830
rect 11430 -3880 11460 -3850
rect 11430 -3900 11435 -3880
rect 11455 -3900 11460 -3880
rect 11430 -3930 11460 -3900
rect 11430 -3950 11435 -3930
rect 11455 -3950 11460 -3930
rect 11430 -3980 11460 -3950
rect 11430 -4000 11435 -3980
rect 11455 -4000 11460 -3980
rect 11430 -4030 11460 -4000
rect 11430 -4050 11435 -4030
rect 11455 -4050 11460 -4030
rect 11430 -4060 11460 -4050
rect 11485 -3830 11515 -3820
rect 11485 -3850 11490 -3830
rect 11510 -3850 11515 -3830
rect 11485 -3880 11515 -3850
rect 11485 -3900 11490 -3880
rect 11510 -3900 11515 -3880
rect 11485 -3930 11515 -3900
rect 11485 -3950 11490 -3930
rect 11510 -3950 11515 -3930
rect 11485 -3980 11515 -3950
rect 11485 -4000 11490 -3980
rect 11510 -4000 11515 -3980
rect 11485 -4030 11515 -4000
rect 11485 -4050 11490 -4030
rect 11510 -4050 11515 -4030
rect 11485 -4060 11515 -4050
rect 11540 -3830 11570 -3820
rect 11540 -3850 11545 -3830
rect 11565 -3850 11570 -3830
rect 11540 -3880 11570 -3850
rect 11540 -3900 11545 -3880
rect 11565 -3900 11570 -3880
rect 11540 -3930 11570 -3900
rect 11540 -3950 11545 -3930
rect 11565 -3950 11570 -3930
rect 11540 -3980 11570 -3950
rect 11540 -4000 11545 -3980
rect 11565 -4000 11570 -3980
rect 11540 -4030 11570 -4000
rect 11540 -4050 11545 -4030
rect 11565 -4050 11570 -4030
rect 11540 -4060 11570 -4050
rect 11595 -3830 11625 -3820
rect 11595 -3850 11600 -3830
rect 11620 -3850 11625 -3830
rect 11595 -3880 11625 -3850
rect 11595 -3900 11600 -3880
rect 11620 -3900 11625 -3880
rect 11595 -3930 11625 -3900
rect 11595 -3950 11600 -3930
rect 11620 -3950 11625 -3930
rect 11595 -3980 11625 -3950
rect 11595 -4000 11600 -3980
rect 11620 -4000 11625 -3980
rect 11595 -4030 11625 -4000
rect 11595 -4050 11600 -4030
rect 11620 -4050 11625 -4030
rect 11595 -4060 11625 -4050
rect 11650 -3830 11680 -3820
rect 11650 -3850 11655 -3830
rect 11675 -3850 11680 -3830
rect 11650 -3880 11680 -3850
rect 11650 -3900 11655 -3880
rect 11675 -3900 11680 -3880
rect 11650 -3930 11680 -3900
rect 11650 -3950 11655 -3930
rect 11675 -3950 11680 -3930
rect 11650 -3980 11680 -3950
rect 11650 -4000 11655 -3980
rect 11675 -4000 11680 -3980
rect 11650 -4030 11680 -4000
rect 11650 -4050 11655 -4030
rect 11675 -4050 11680 -4030
rect 11650 -4060 11680 -4050
rect 11705 -3830 11735 -3820
rect 11705 -3850 11710 -3830
rect 11730 -3850 11735 -3830
rect 11705 -3880 11735 -3850
rect 11705 -3900 11710 -3880
rect 11730 -3900 11735 -3880
rect 11705 -3930 11735 -3900
rect 11705 -3950 11710 -3930
rect 11730 -3950 11735 -3930
rect 11705 -3980 11735 -3950
rect 11705 -4000 11710 -3980
rect 11730 -4000 11735 -3980
rect 11705 -4030 11735 -4000
rect 11705 -4050 11710 -4030
rect 11730 -4050 11735 -4030
rect 11705 -4060 11735 -4050
rect 11760 -3830 11790 -3820
rect 11760 -3850 11765 -3830
rect 11785 -3850 11790 -3830
rect 11760 -3880 11790 -3850
rect 11760 -3900 11765 -3880
rect 11785 -3900 11790 -3880
rect 11760 -3930 11790 -3900
rect 11760 -3950 11765 -3930
rect 11785 -3950 11790 -3930
rect 11760 -3980 11790 -3950
rect 11760 -4000 11765 -3980
rect 11785 -4000 11790 -3980
rect 11760 -4030 11790 -4000
rect 11760 -4050 11765 -4030
rect 11785 -4050 11790 -4030
rect 11760 -4060 11790 -4050
rect 11815 -3830 11845 -3820
rect 11815 -3850 11820 -3830
rect 11840 -3850 11845 -3830
rect 11815 -3880 11845 -3850
rect 11815 -3900 11820 -3880
rect 11840 -3900 11845 -3880
rect 11815 -3930 11845 -3900
rect 11815 -3950 11820 -3930
rect 11840 -3950 11845 -3930
rect 11815 -3980 11845 -3950
rect 11815 -4000 11820 -3980
rect 11840 -4000 11845 -3980
rect 11815 -4030 11845 -4000
rect 11815 -4050 11820 -4030
rect 11840 -4050 11845 -4030
rect 11815 -4060 11845 -4050
rect 11870 -3830 11900 -3820
rect 11870 -3850 11875 -3830
rect 11895 -3850 11900 -3830
rect 11870 -3880 11900 -3850
rect 11870 -3900 11875 -3880
rect 11895 -3900 11900 -3880
rect 11870 -3930 11900 -3900
rect 11870 -3950 11875 -3930
rect 11895 -3950 11900 -3930
rect 11870 -3980 11900 -3950
rect 11870 -4000 11875 -3980
rect 11895 -4000 11900 -3980
rect 11870 -4030 11900 -4000
rect 11870 -4050 11875 -4030
rect 11895 -4050 11900 -4030
rect 11870 -4060 11900 -4050
rect 11925 -3830 11955 -3820
rect 11925 -3850 11930 -3830
rect 11950 -3850 11955 -3830
rect 11925 -3880 11955 -3850
rect 11925 -3900 11930 -3880
rect 11950 -3900 11955 -3880
rect 11925 -3930 11955 -3900
rect 11925 -3950 11930 -3930
rect 11950 -3950 11955 -3930
rect 11925 -3980 11955 -3950
rect 11925 -4000 11930 -3980
rect 11950 -4000 11955 -3980
rect 11925 -4030 11955 -4000
rect 11925 -4050 11930 -4030
rect 11950 -4050 11955 -4030
rect 11925 -4060 11955 -4050
rect 11980 -3830 12010 -3820
rect 11980 -3850 11985 -3830
rect 12005 -3850 12010 -3830
rect 11980 -3880 12010 -3850
rect 11980 -3900 11985 -3880
rect 12005 -3900 12010 -3880
rect 11980 -3930 12010 -3900
rect 11980 -3950 11985 -3930
rect 12005 -3950 12010 -3930
rect 11980 -3980 12010 -3950
rect 11980 -4000 11985 -3980
rect 12005 -4000 12010 -3980
rect 11980 -4030 12010 -4000
rect 11980 -4050 11985 -4030
rect 12005 -4050 12010 -4030
rect 11980 -4060 12010 -4050
rect 12035 -3830 12065 -3820
rect 12035 -3850 12040 -3830
rect 12060 -3850 12065 -3830
rect 12035 -3880 12065 -3850
rect 12035 -3900 12040 -3880
rect 12060 -3900 12065 -3880
rect 12035 -3930 12065 -3900
rect 12035 -3950 12040 -3930
rect 12060 -3950 12065 -3930
rect 12035 -3980 12065 -3950
rect 12035 -4000 12040 -3980
rect 12060 -4000 12065 -3980
rect 12035 -4030 12065 -4000
rect 12035 -4050 12040 -4030
rect 12060 -4050 12065 -4030
rect 12035 -4060 12065 -4050
rect 12090 -3830 12120 -3820
rect 12090 -3850 12095 -3830
rect 12115 -3850 12120 -3830
rect 12090 -3880 12120 -3850
rect 12090 -3900 12095 -3880
rect 12115 -3900 12120 -3880
rect 12090 -3930 12120 -3900
rect 12090 -3950 12095 -3930
rect 12115 -3950 12120 -3930
rect 12090 -3980 12120 -3950
rect 12090 -4000 12095 -3980
rect 12115 -4000 12120 -3980
rect 12090 -4030 12120 -4000
rect 12090 -4050 12095 -4030
rect 12115 -4050 12120 -4030
rect 12090 -4060 12120 -4050
rect 12145 -3830 12175 -3820
rect 12145 -3850 12150 -3830
rect 12170 -3850 12175 -3830
rect 12145 -3880 12175 -3850
rect 12145 -3900 12150 -3880
rect 12170 -3900 12175 -3880
rect 12145 -3930 12175 -3900
rect 12145 -3950 12150 -3930
rect 12170 -3950 12175 -3930
rect 12145 -3980 12175 -3950
rect 12145 -4000 12150 -3980
rect 12170 -4000 12175 -3980
rect 12145 -4030 12175 -4000
rect 12145 -4050 12150 -4030
rect 12170 -4050 12175 -4030
rect 12145 -4060 12175 -4050
rect 12200 -3830 12230 -3820
rect 12200 -3850 12205 -3830
rect 12225 -3850 12230 -3830
rect 12200 -3880 12230 -3850
rect 12200 -3900 12205 -3880
rect 12225 -3900 12230 -3880
rect 12200 -3930 12230 -3900
rect 12200 -3950 12205 -3930
rect 12225 -3950 12230 -3930
rect 12200 -3980 12230 -3950
rect 12200 -4000 12205 -3980
rect 12225 -4000 12230 -3980
rect 12200 -4030 12230 -4000
rect 12200 -4050 12205 -4030
rect 12225 -4050 12230 -4030
rect 12200 -4060 12230 -4050
rect 12255 -3830 12285 -3820
rect 12255 -3850 12260 -3830
rect 12280 -3850 12285 -3830
rect 12255 -3880 12285 -3850
rect 12255 -3900 12260 -3880
rect 12280 -3900 12285 -3880
rect 12255 -3930 12285 -3900
rect 12255 -3950 12260 -3930
rect 12280 -3950 12285 -3930
rect 12255 -3980 12285 -3950
rect 12255 -4000 12260 -3980
rect 12280 -4000 12285 -3980
rect 12255 -4030 12285 -4000
rect 12255 -4050 12260 -4030
rect 12280 -4050 12285 -4030
rect 12255 -4060 12285 -4050
rect 12310 -3830 12340 -3820
rect 12310 -3850 12315 -3830
rect 12335 -3850 12340 -3830
rect 12310 -3880 12340 -3850
rect 12310 -3900 12315 -3880
rect 12335 -3900 12340 -3880
rect 12310 -3930 12340 -3900
rect 12310 -3950 12315 -3930
rect 12335 -3950 12340 -3930
rect 12310 -3980 12340 -3950
rect 12310 -4000 12315 -3980
rect 12335 -4000 12340 -3980
rect 12310 -4030 12340 -4000
rect 12310 -4050 12315 -4030
rect 12335 -4050 12340 -4030
rect 12310 -4060 12340 -4050
rect 12365 -3830 12395 -3820
rect 12365 -3850 12370 -3830
rect 12390 -3850 12395 -3830
rect 12365 -3880 12395 -3850
rect 12365 -3900 12370 -3880
rect 12390 -3900 12395 -3880
rect 12365 -3930 12395 -3900
rect 12365 -3950 12370 -3930
rect 12390 -3950 12395 -3930
rect 12365 -3980 12395 -3950
rect 12365 -4000 12370 -3980
rect 12390 -4000 12395 -3980
rect 12365 -4030 12395 -4000
rect 12365 -4050 12370 -4030
rect 12390 -4050 12395 -4030
rect 12365 -4060 12395 -4050
rect 12420 -3830 12450 -3820
rect 12420 -3850 12425 -3830
rect 12445 -3850 12450 -3830
rect 12420 -3880 12450 -3850
rect 12420 -3900 12425 -3880
rect 12445 -3900 12450 -3880
rect 12420 -3930 12450 -3900
rect 12420 -3950 12425 -3930
rect 12445 -3950 12450 -3930
rect 12420 -3980 12450 -3950
rect 12420 -4000 12425 -3980
rect 12445 -4000 12450 -3980
rect 12420 -4030 12450 -4000
rect 12420 -4050 12425 -4030
rect 12445 -4050 12450 -4030
rect 12420 -4060 12450 -4050
rect 12475 -3830 12505 -3820
rect 12475 -3850 12480 -3830
rect 12500 -3850 12505 -3830
rect 12475 -3880 12505 -3850
rect 12475 -3900 12480 -3880
rect 12500 -3900 12505 -3880
rect 12475 -3930 12505 -3900
rect 12475 -3950 12480 -3930
rect 12500 -3950 12505 -3930
rect 12475 -3980 12505 -3950
rect 12475 -4000 12480 -3980
rect 12500 -4000 12505 -3980
rect 12475 -4030 12505 -4000
rect 12475 -4050 12480 -4030
rect 12500 -4050 12505 -4030
rect 12475 -4060 12505 -4050
rect 12530 -3830 12560 -3820
rect 12530 -3850 12535 -3830
rect 12555 -3850 12560 -3830
rect 12530 -3880 12560 -3850
rect 12530 -3900 12535 -3880
rect 12555 -3900 12560 -3880
rect 12530 -3930 12560 -3900
rect 12530 -3950 12535 -3930
rect 12555 -3950 12560 -3930
rect 12530 -3980 12560 -3950
rect 12530 -4000 12535 -3980
rect 12555 -4000 12560 -3980
rect 12530 -4030 12560 -4000
rect 12530 -4050 12535 -4030
rect 12555 -4050 12560 -4030
rect 12530 -4060 12560 -4050
rect 12585 -3830 12655 -3820
rect 12585 -3850 12590 -3830
rect 12610 -3850 12630 -3830
rect 12650 -3850 12655 -3830
rect 12585 -3880 12655 -3850
rect 12585 -3900 12590 -3880
rect 12610 -3900 12630 -3880
rect 12650 -3900 12655 -3880
rect 12585 -3930 12655 -3900
rect 12585 -3950 12590 -3930
rect 12610 -3950 12630 -3930
rect 12650 -3950 12655 -3930
rect 12585 -3980 12655 -3950
rect 12585 -4000 12590 -3980
rect 12610 -4000 12630 -3980
rect 12650 -4000 12655 -3980
rect 12585 -4030 12655 -4000
rect 12585 -4050 12590 -4030
rect 12610 -4050 12630 -4030
rect 12650 -4050 12655 -4030
rect 12585 -4060 12655 -4050
rect 11175 -4080 11195 -4060
rect 11270 -4080 11290 -4060
rect 11380 -4080 11400 -4060
rect 11490 -4080 11510 -4060
rect 11600 -4080 11620 -4060
rect 11710 -4080 11730 -4060
rect 11820 -4080 11840 -4060
rect 11930 -4080 11950 -4060
rect 12040 -4080 12060 -4060
rect 12150 -4080 12170 -4060
rect 12260 -4080 12280 -4060
rect 12370 -4080 12390 -4060
rect 12480 -4080 12500 -4060
rect 12630 -4080 12650 -4060
rect 11165 -4090 11205 -4080
rect 11165 -4110 11175 -4090
rect 11195 -4110 11205 -4090
rect 11165 -4120 11205 -4110
rect 11260 -4090 11300 -4080
rect 11260 -4110 11270 -4090
rect 11290 -4110 11300 -4090
rect 11260 -4120 11300 -4110
rect 11370 -4090 11410 -4080
rect 11370 -4110 11380 -4090
rect 11400 -4110 11410 -4090
rect 11370 -4120 11410 -4110
rect 11480 -4090 11520 -4080
rect 11480 -4110 11490 -4090
rect 11510 -4110 11520 -4090
rect 11480 -4120 11520 -4110
rect 11590 -4090 11630 -4080
rect 11590 -4110 11600 -4090
rect 11620 -4110 11630 -4090
rect 11590 -4120 11630 -4110
rect 11700 -4090 11740 -4080
rect 11700 -4110 11710 -4090
rect 11730 -4110 11740 -4090
rect 11700 -4120 11740 -4110
rect 11810 -4090 11850 -4080
rect 11810 -4110 11820 -4090
rect 11840 -4110 11850 -4090
rect 11810 -4120 11850 -4110
rect 11920 -4090 11960 -4080
rect 11920 -4110 11930 -4090
rect 11950 -4110 11960 -4090
rect 11920 -4120 11960 -4110
rect 12030 -4090 12070 -4080
rect 12030 -4110 12040 -4090
rect 12060 -4110 12070 -4090
rect 12030 -4120 12070 -4110
rect 12140 -4090 12180 -4080
rect 12140 -4110 12150 -4090
rect 12170 -4110 12180 -4090
rect 12140 -4120 12180 -4110
rect 12250 -4090 12290 -4080
rect 12250 -4110 12260 -4090
rect 12280 -4110 12290 -4090
rect 12250 -4120 12290 -4110
rect 12360 -4090 12400 -4080
rect 12360 -4110 12370 -4090
rect 12390 -4110 12400 -4090
rect 12360 -4120 12400 -4110
rect 12470 -4090 12510 -4080
rect 12470 -4110 12480 -4090
rect 12500 -4110 12510 -4090
rect 12470 -4120 12510 -4110
rect 12620 -4090 12660 -4080
rect 12620 -4110 12630 -4090
rect 12650 -4110 12660 -4090
rect 12620 -4120 12660 -4110
<< viali >>
rect 11640 9030 11660 9050
rect 11760 9030 11780 9050
rect 11880 9030 11900 9050
rect 11210 8970 11230 8990
rect 11470 8970 11490 8990
rect 11580 8985 11600 9005
rect 11700 8985 11720 9005
rect 11820 8985 11840 9005
rect 11940 8985 11960 9005
rect 12090 8960 12110 8980
rect 12210 8960 12230 8980
rect 12330 8960 12350 8980
rect 12450 8960 12470 8980
rect 12570 8960 12590 8980
rect 11340 8855 11360 8860
rect 11340 8835 11360 8855
rect 11760 8830 11780 8850
rect 12150 8830 12170 8850
rect 12211 8830 12229 8850
rect 12270 8830 12290 8850
rect 12390 8830 12410 8850
rect 12510 8830 12530 8850
rect 11350 8600 11370 8620
rect 11470 8600 11490 8620
rect 11590 8600 11610 8620
rect 11710 8600 11730 8620
rect 11830 8600 11850 8620
rect 11950 8600 11970 8620
rect 12070 8600 12090 8620
rect 12190 8600 12210 8620
rect 12310 8600 12330 8620
rect 12430 8600 12450 8620
rect 18850 8600 18870 8620
rect 18970 8600 18990 8620
rect 19090 8600 19110 8620
rect 19210 8600 19230 8620
rect 19330 8600 19350 8620
rect 19450 8600 19470 8620
rect 19570 8600 19590 8620
rect 19690 8600 19710 8620
rect 19810 8600 19830 8620
rect 19930 8600 19950 8620
rect 10590 8185 10610 8205
rect 10910 8185 10930 8205
rect 10990 8185 11010 8205
rect 12960 8265 12980 8285
rect 13070 8265 13090 8285
rect 13180 8265 13200 8285
rect 13290 8265 13310 8285
rect 13400 8265 13420 8285
rect 13510 8265 13530 8285
rect 13620 8265 13640 8285
rect 13730 8265 13750 8285
rect 13840 8265 13860 8285
rect 13950 8265 13970 8285
rect 14060 8265 14080 8285
rect 11290 8130 11310 8150
rect 11410 8130 11430 8150
rect 11530 8130 11550 8150
rect 11650 8130 11670 8150
rect 11770 8130 11790 8150
rect 11831 8130 11849 8150
rect 11890 8130 11910 8150
rect 12010 8130 12030 8150
rect 12130 8130 12150 8150
rect 12250 8130 12270 8150
rect 12370 8130 12390 8150
rect 12490 8130 12510 8150
rect 11350 7920 11370 7940
rect 11470 7920 11490 7940
rect 11590 7920 11610 7940
rect 11710 7920 11730 7940
rect 11830 7920 11850 7940
rect 11950 7920 11970 7940
rect 12070 7920 12090 7940
rect 12190 7920 12210 7940
rect 12310 7920 12330 7940
rect 12430 7920 12450 7940
rect 18090 8185 18110 8205
rect 18410 8185 18430 8205
rect 18490 8185 18510 8205
rect 20455 8265 20475 8285
rect 20565 8265 20585 8285
rect 20675 8265 20695 8285
rect 20785 8265 20805 8285
rect 20895 8265 20915 8285
rect 21005 8265 21025 8285
rect 21115 8265 21135 8285
rect 21225 8265 21245 8285
rect 21335 8265 21355 8285
rect 21445 8265 21465 8285
rect 21555 8265 21575 8285
rect 18790 8130 18810 8150
rect 18910 8130 18930 8150
rect 19030 8130 19050 8150
rect 19150 8130 19170 8150
rect 19270 8130 19290 8150
rect 19331 8130 19349 8150
rect 19390 8130 19410 8150
rect 19510 8130 19530 8150
rect 19630 8130 19650 8150
rect 19750 8130 19770 8150
rect 19870 8130 19890 8150
rect 19990 8130 20010 8150
rect 9745 7645 9765 7665
rect 9855 7645 9875 7665
rect 9965 7645 9985 7665
rect 10075 7645 10095 7665
rect 10185 7645 10205 7665
rect 10295 7645 10315 7665
rect 10405 7645 10425 7665
rect 10515 7645 10535 7665
rect 10625 7645 10645 7665
rect 10735 7645 10755 7665
rect 10845 7645 10865 7665
rect 9800 7475 9820 7495
rect 9910 7475 9930 7495
rect 10020 7475 10040 7495
rect 10130 7475 10150 7495
rect 10240 7475 10260 7495
rect 10350 7475 10370 7495
rect 10460 7475 10480 7495
rect 10570 7475 10590 7495
rect 10680 7475 10700 7495
rect 10790 7475 10810 7495
rect 13015 7895 13035 7915
rect 13071 7895 13089 7915
rect 13125 7895 13145 7915
rect 13235 7895 13255 7915
rect 13345 7895 13365 7915
rect 13455 7895 13475 7915
rect 13565 7895 13585 7915
rect 13675 7895 13695 7915
rect 13785 7895 13805 7915
rect 13895 7895 13915 7915
rect 14005 7895 14025 7915
rect 18850 7920 18870 7940
rect 18970 7920 18990 7940
rect 19090 7920 19110 7940
rect 19210 7920 19230 7940
rect 19330 7920 19350 7940
rect 19450 7920 19470 7940
rect 19570 7920 19590 7940
rect 19690 7920 19710 7940
rect 19810 7920 19830 7940
rect 19930 7920 19950 7940
rect 12960 7645 12980 7665
rect 13070 7645 13090 7665
rect 13180 7645 13200 7665
rect 13290 7645 13310 7665
rect 13400 7645 13420 7665
rect 13510 7645 13530 7665
rect 13620 7645 13640 7665
rect 13730 7645 13750 7665
rect 13840 7645 13860 7665
rect 13950 7645 13970 7665
rect 14060 7645 14080 7665
rect 17245 7645 17265 7665
rect 17355 7645 17375 7665
rect 17465 7645 17485 7665
rect 17575 7645 17595 7665
rect 17685 7645 17705 7665
rect 17795 7645 17815 7665
rect 17905 7645 17925 7665
rect 18015 7645 18035 7665
rect 18125 7645 18145 7665
rect 18235 7645 18255 7665
rect 18345 7645 18365 7665
rect 11290 7450 11310 7470
rect 11410 7450 11430 7470
rect 11530 7450 11550 7470
rect 11650 7450 11670 7470
rect 11770 7450 11790 7470
rect 11831 7450 11849 7470
rect 11890 7450 11910 7470
rect 12010 7450 12030 7470
rect 12130 7450 12150 7470
rect 12250 7450 12270 7470
rect 12370 7450 12390 7470
rect 12490 7450 12510 7470
rect 13015 7475 13035 7495
rect 13125 7475 13145 7495
rect 13235 7475 13255 7495
rect 13345 7475 13365 7495
rect 13455 7475 13475 7495
rect 13565 7475 13585 7495
rect 13675 7475 13695 7495
rect 13785 7475 13805 7495
rect 13895 7475 13915 7495
rect 14005 7475 14025 7495
rect 17300 7475 17320 7495
rect 17410 7475 17430 7495
rect 17520 7475 17540 7495
rect 17630 7475 17650 7495
rect 17740 7475 17760 7495
rect 17850 7475 17870 7495
rect 17960 7475 17980 7495
rect 18070 7475 18090 7495
rect 18180 7475 18200 7495
rect 18290 7475 18310 7495
rect 20510 7895 20530 7915
rect 20566 7895 20584 7915
rect 20620 7895 20640 7915
rect 20730 7895 20750 7915
rect 20840 7895 20860 7915
rect 20950 7895 20970 7915
rect 21060 7895 21080 7915
rect 21170 7895 21190 7915
rect 21280 7895 21300 7915
rect 21390 7895 21410 7915
rect 21500 7895 21520 7915
rect 20455 7645 20475 7665
rect 20565 7645 20585 7665
rect 20675 7645 20695 7665
rect 20785 7645 20805 7665
rect 20895 7645 20915 7665
rect 21005 7645 21025 7665
rect 21115 7645 21135 7665
rect 21225 7645 21245 7665
rect 21335 7645 21355 7665
rect 21445 7645 21465 7665
rect 21555 7645 21575 7665
rect 18790 7450 18810 7470
rect 10821 7415 10839 7435
rect 12986 7415 13004 7435
rect 18910 7450 18930 7470
rect 19030 7450 19050 7470
rect 19150 7450 19170 7470
rect 19270 7450 19290 7470
rect 19331 7450 19349 7470
rect 19390 7450 19410 7470
rect 19510 7450 19530 7470
rect 19630 7450 19650 7470
rect 19750 7450 19770 7470
rect 19870 7450 19890 7470
rect 19990 7450 20010 7470
rect 20510 7475 20530 7495
rect 20620 7475 20640 7495
rect 20730 7475 20750 7495
rect 20840 7475 20860 7495
rect 20950 7475 20970 7495
rect 21060 7475 21080 7495
rect 21170 7475 21190 7495
rect 21280 7475 21300 7495
rect 21390 7475 21410 7495
rect 21500 7475 21520 7495
rect 18321 7415 18339 7435
rect 20481 7415 20499 7435
rect 9810 7350 9835 7375
rect 10645 7350 10670 7375
rect 13155 7350 13180 7375
rect 13990 7350 14015 7375
rect 17310 7350 17335 7375
rect 18145 7350 18170 7375
rect 20650 7350 20675 7375
rect 21485 7350 21510 7375
rect 9810 7290 9835 7315
rect 10645 7290 10670 7315
rect 13155 7290 13180 7315
rect 13990 7290 14015 7315
rect 17310 7290 17335 7315
rect 18145 7290 18170 7315
rect 20650 7290 20675 7315
rect 21485 7290 21510 7315
rect 10821 7255 10839 7275
rect 12986 7255 13004 7275
rect 18321 7255 18339 7275
rect 20481 7255 20499 7275
rect 9800 7195 9820 7215
rect 9910 7195 9930 7215
rect 10020 7195 10040 7215
rect 10130 7195 10150 7215
rect 10240 7195 10260 7215
rect 10350 7195 10370 7215
rect 10460 7195 10480 7215
rect 10570 7195 10590 7215
rect 10680 7195 10700 7215
rect 10790 7195 10810 7215
rect 13015 7195 13035 7215
rect 13125 7195 13145 7215
rect 13235 7195 13255 7215
rect 13345 7195 13365 7215
rect 13455 7195 13475 7215
rect 13565 7195 13585 7215
rect 13675 7195 13695 7215
rect 13785 7195 13805 7215
rect 13895 7195 13915 7215
rect 14005 7195 14025 7215
rect 17300 7195 17320 7215
rect 17410 7195 17430 7215
rect 17520 7195 17540 7215
rect 17630 7195 17650 7215
rect 17740 7195 17760 7215
rect 17850 7195 17870 7215
rect 17960 7195 17980 7215
rect 18070 7195 18090 7215
rect 18180 7195 18200 7215
rect 18290 7195 18310 7215
rect 20510 7195 20530 7215
rect 20620 7195 20640 7215
rect 20730 7195 20750 7215
rect 20840 7195 20860 7215
rect 20950 7195 20970 7215
rect 21060 7195 21080 7215
rect 21170 7195 21190 7215
rect 21280 7195 21300 7215
rect 21390 7195 21410 7215
rect 21500 7195 21520 7215
rect 11340 7155 11360 7175
rect 11450 7155 11470 7175
rect 11560 7155 11580 7175
rect 11670 7155 11690 7175
rect 11780 7155 11800 7175
rect 11890 7155 11910 7175
rect 12000 7155 12020 7175
rect 12110 7155 12130 7175
rect 12220 7155 12240 7175
rect 12330 7155 12350 7175
rect 12440 7155 12460 7175
rect 9745 6975 9763 6995
rect 9855 6975 9873 6995
rect 9965 6975 9983 6995
rect 10075 6975 10093 6995
rect 10185 6975 10203 6995
rect 10295 6975 10313 6995
rect 10405 6975 10423 6995
rect 10515 6975 10533 6995
rect 10625 6975 10643 6995
rect 10735 6975 10753 6995
rect 10845 6975 10863 6995
rect 18840 7155 18860 7175
rect 18950 7155 18970 7175
rect 19060 7155 19080 7175
rect 19170 7155 19190 7175
rect 19280 7155 19300 7175
rect 19390 7155 19410 7175
rect 19500 7155 19520 7175
rect 19610 7155 19630 7175
rect 19720 7155 19740 7175
rect 19830 7155 19850 7175
rect 19940 7155 19960 7175
rect 12962 6975 12980 6995
rect 13072 6975 13090 6995
rect 13182 6975 13200 6995
rect 13292 6975 13310 6995
rect 13402 6975 13420 6995
rect 13512 6975 13530 6995
rect 13622 6975 13640 6995
rect 13732 6975 13750 6995
rect 13842 6975 13860 6995
rect 13952 6975 13970 6995
rect 14062 6975 14080 6995
rect 17245 6975 17263 6995
rect 17355 6975 17373 6995
rect 17465 6975 17483 6995
rect 17575 6975 17593 6995
rect 17685 6975 17703 6995
rect 17795 6975 17813 6995
rect 17905 6975 17923 6995
rect 18015 6975 18033 6995
rect 18125 6975 18143 6995
rect 18235 6975 18253 6995
rect 18345 6975 18363 6995
rect 20457 6975 20475 6995
rect 20567 6975 20585 6995
rect 20677 6975 20695 6995
rect 20787 6975 20805 6995
rect 20897 6975 20915 6995
rect 21007 6975 21025 6995
rect 21117 6975 21135 6995
rect 21227 6975 21245 6995
rect 21337 6975 21355 6995
rect 21447 6975 21465 6995
rect 21557 6975 21575 6995
rect 11395 6935 11415 6955
rect 11505 6935 11525 6955
rect 11615 6935 11635 6955
rect 11725 6935 11745 6955
rect 11835 6935 11855 6955
rect 11945 6935 11965 6955
rect 12055 6935 12075 6955
rect 12165 6935 12185 6955
rect 12275 6935 12295 6955
rect 12385 6935 12405 6955
rect 18895 6935 18915 6955
rect 19005 6935 19025 6955
rect 19115 6935 19135 6955
rect 19225 6935 19245 6955
rect 19335 6935 19355 6955
rect 19445 6935 19465 6955
rect 19555 6935 19575 6955
rect 19665 6935 19685 6955
rect 19775 6935 19795 6955
rect 19885 6935 19905 6955
rect 20555 6880 20575 6900
rect 20665 6880 20685 6900
rect 20775 6880 20795 6900
rect 11095 6735 11115 6755
rect 11200 6750 11220 6770
rect 11315 6735 11335 6755
rect 11420 6750 11440 6770
rect 11243 6690 11260 6710
rect 11535 6735 11555 6755
rect 11650 6750 11670 6770
rect 11463 6690 11480 6710
rect 11610 6690 11627 6710
rect 12135 6735 12155 6755
rect 12240 6750 12260 6770
rect 11825 6690 11845 6710
rect 11876 6690 11893 6710
rect 11955 6690 11975 6710
rect 12355 6735 12375 6755
rect 12460 6750 12480 6770
rect 12283 6690 12300 6710
rect 12575 6735 12595 6755
rect 12690 6750 12710 6770
rect 12503 6690 12520 6710
rect 12650 6690 12667 6710
rect 18595 6735 18615 6755
rect 18700 6750 18720 6770
rect 18815 6735 18835 6755
rect 18920 6750 18940 6770
rect 18743 6690 18760 6710
rect 19035 6735 19055 6755
rect 19150 6750 19170 6770
rect 18963 6690 18980 6710
rect 19110 6690 19127 6710
rect 19635 6735 19655 6755
rect 19740 6750 19760 6770
rect 19325 6690 19345 6710
rect 19376 6690 19393 6710
rect 19455 6690 19475 6710
rect 19855 6735 19875 6755
rect 19960 6750 19980 6770
rect 19783 6690 19800 6710
rect 20075 6735 20095 6755
rect 20190 6750 20210 6770
rect 20003 6690 20020 6710
rect 20150 6690 20167 6710
rect 20571 6655 20591 6675
rect 20625 6660 20645 6680
rect 20720 6660 20740 6680
rect 20520 6605 20540 6625
rect 20810 6605 20830 6625
rect 20476 6545 20496 6565
rect 11112 6470 11129 6490
rect 9770 6415 9795 6440
rect 11315 6470 11335 6490
rect 11535 6470 11555 6490
rect 11830 6470 11850 6490
rect 11880 6470 11900 6490
rect 11928 6470 11945 6490
rect 12152 6470 12169 6490
rect 12355 6470 12375 6490
rect 12575 6470 12595 6490
rect 18612 6470 18629 6490
rect 10780 6415 10805 6440
rect 11155 6410 11175 6430
rect 11260 6410 11280 6430
rect 11370 6410 11390 6430
rect 11480 6410 11500 6430
rect 11590 6410 11610 6430
rect 12195 6410 12215 6430
rect 12300 6410 12320 6430
rect 12410 6410 12430 6430
rect 12520 6410 12540 6430
rect 12630 6410 12650 6430
rect 12995 6415 13020 6440
rect 18815 6470 18835 6490
rect 19035 6470 19055 6490
rect 19330 6470 19350 6490
rect 19380 6470 19400 6490
rect 19428 6470 19445 6490
rect 19652 6470 19669 6490
rect 19855 6470 19875 6490
rect 20075 6470 20095 6490
rect 20570 6545 20590 6565
rect 20854 6545 20874 6565
rect 14005 6415 14030 6440
rect 18655 6410 18675 6430
rect 18760 6410 18780 6430
rect 18870 6410 18890 6430
rect 18980 6410 19000 6430
rect 19090 6410 19110 6430
rect 19695 6410 19715 6430
rect 19800 6410 19820 6430
rect 19910 6410 19930 6430
rect 20020 6410 20040 6430
rect 20130 6410 20150 6430
rect 9775 6310 9795 6330
rect 9975 6310 9995 6330
rect 10175 6310 10195 6330
rect 10375 6310 10395 6330
rect 10575 6310 10595 6330
rect 10676 6310 10694 6330
rect 10775 6310 10795 6330
rect 13005 6310 13025 6330
rect 13106 6310 13124 6330
rect 13205 6310 13225 6330
rect 13405 6310 13425 6330
rect 13605 6310 13625 6330
rect 13805 6310 13825 6330
rect 14005 6310 14025 6330
rect 20533 6325 20553 6345
rect 20797 6325 20817 6345
rect 11325 6210 11345 6230
rect 11435 6210 11455 6230
rect 11545 6210 11565 6230
rect 11655 6210 11675 6230
rect 11765 6210 11785 6230
rect 11820 6210 11840 6230
rect 11875 6210 11895 6230
rect 11985 6210 12005 6230
rect 12095 6210 12115 6230
rect 12205 6210 12225 6230
rect 12315 6210 12335 6230
rect 12425 6210 12445 6230
rect 12535 6210 12555 6230
rect 12605 6225 12625 6245
rect 9875 5960 9895 5980
rect 10075 5960 10095 5980
rect 10275 5960 10295 5980
rect 10475 5960 10495 5980
rect 10675 5960 10695 5980
rect 18825 6250 18845 6270
rect 18935 6250 18955 6270
rect 19045 6250 19065 6270
rect 19155 6250 19175 6270
rect 19265 6250 19285 6270
rect 19320 6250 19340 6270
rect 19375 6250 19395 6270
rect 19485 6250 19505 6270
rect 19595 6250 19615 6270
rect 19705 6250 19725 6270
rect 19815 6250 19835 6270
rect 19925 6250 19945 6270
rect 20035 6250 20055 6270
rect 20105 6265 20125 6285
rect 20455 6265 20475 6285
rect 20570 6265 20590 6285
rect 20760 6265 20780 6285
rect 20875 6265 20895 6285
rect 13105 5960 13125 5980
rect 13305 5960 13325 5980
rect 13505 5960 13525 5980
rect 13705 5960 13725 5980
rect 13905 5960 13925 5980
rect 20610 6205 20630 6225
rect 20665 6205 20685 6225
rect 20720 6205 20740 6225
rect 18675 5930 18695 5950
rect 18770 5930 18790 5950
rect 18880 5930 18900 5950
rect 18990 5930 19010 5950
rect 19100 5930 19120 5950
rect 19210 5930 19230 5950
rect 19320 5930 19340 5950
rect 19430 5930 19450 5950
rect 19540 5930 19560 5950
rect 19650 5930 19670 5950
rect 19760 5930 19780 5950
rect 19870 5930 19890 5950
rect 19980 5930 20000 5950
rect 20130 5930 20150 5950
rect 11175 5890 11195 5910
rect 11270 5890 11290 5910
rect 11380 5890 11400 5910
rect 11490 5890 11510 5910
rect 11600 5890 11620 5910
rect 11710 5890 11730 5910
rect 11820 5890 11840 5910
rect 11930 5890 11950 5910
rect 12040 5890 12060 5910
rect 12150 5890 12170 5910
rect 12260 5890 12280 5910
rect 12370 5890 12390 5910
rect 12480 5890 12500 5910
rect 12630 5890 12650 5910
rect 11640 4490 11660 4510
rect 11760 4490 11780 4510
rect 11880 4490 11900 4510
rect 11210 4430 11230 4450
rect 11470 4430 11490 4450
rect 11580 4445 11600 4465
rect 11700 4445 11720 4465
rect 11820 4445 11840 4465
rect 11940 4445 11960 4465
rect 12090 4420 12110 4440
rect 12210 4420 12230 4440
rect 12330 4420 12350 4440
rect 12450 4420 12470 4440
rect 12570 4420 12590 4440
rect 11340 4315 11360 4320
rect 11340 4295 11360 4315
rect 11760 4290 11780 4310
rect 12150 4290 12170 4310
rect 12211 4290 12229 4310
rect 12270 4290 12290 4310
rect 12390 4290 12410 4310
rect 12510 4290 12530 4310
rect 11370 4180 11390 4200
rect 11480 4180 11500 4200
rect 11590 4180 11610 4200
rect 11700 4180 11720 4200
rect 11810 4180 11830 4200
rect 11920 4180 11940 4200
rect 12030 4180 12050 4200
rect 12140 4180 12160 4200
rect 12250 4180 12270 4200
rect 12360 4180 12380 4200
rect 11315 4060 11335 4080
rect 11370 4060 11390 4080
rect 11425 4060 11445 4080
rect 11535 4060 11555 4080
rect 11645 4060 11665 4080
rect 11755 4060 11775 4080
rect 11865 4060 11885 4080
rect 11975 4060 11995 4080
rect 12085 4060 12105 4080
rect 12195 4060 12215 4080
rect 12305 4060 12325 4080
rect 12415 4060 12435 4080
rect 11320 3935 11340 3955
rect 11425 3935 11445 3955
rect 11535 3935 11555 3955
rect 11645 3935 11665 3955
rect 11755 3935 11775 3955
rect 12060 3935 12080 3955
rect 12165 3935 12185 3955
rect 12275 3935 12295 3955
rect 12385 3935 12405 3955
rect 12495 3935 12515 3955
rect 11277 3875 11294 3895
rect 11370 3875 11390 3895
rect 11480 3875 11500 3895
rect 11700 3875 11720 3895
rect 11810 3875 11830 3895
rect 12017 3875 12034 3895
rect 12220 3875 12240 3895
rect 12440 3875 12460 3895
rect 11408 3755 11425 3775
rect 11628 3755 11645 3775
rect 11775 3755 11792 3775
rect 11260 3695 11280 3715
rect 11365 3695 11385 3715
rect 11480 3695 11500 3715
rect 11585 3695 11605 3715
rect 11700 3695 11720 3715
rect 11815 3695 11835 3715
rect 12000 3705 12020 3725
rect 12148 3755 12165 3775
rect 12220 3705 12240 3725
rect 12368 3755 12385 3775
rect 12515 3755 12532 3775
rect 12440 3705 12460 3725
rect 10220 3610 10240 3630
rect 10330 3610 10350 3630
rect 10440 3610 10460 3630
rect 10550 3610 10570 3630
rect 10660 3610 10680 3630
rect 10770 3610 10790 3630
rect 11350 3600 11370 3620
rect 11470 3600 11490 3620
rect 11590 3600 11610 3620
rect 11710 3600 11730 3620
rect 11830 3600 11850 3620
rect 11950 3600 11970 3620
rect 12070 3600 12090 3620
rect 12190 3600 12210 3620
rect 12310 3600 12330 3620
rect 12430 3600 12450 3620
rect 13010 3610 13030 3630
rect 13120 3610 13140 3630
rect 13230 3610 13250 3630
rect 13340 3610 13360 3630
rect 13450 3610 13470 3630
rect 13560 3610 13580 3630
rect 56 3175 81 3200
rect 1271 3170 1296 3195
rect 56 3115 81 3140
rect 1271 3110 1296 3135
rect 56 3035 81 3060
rect 56 2975 81 3000
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 2340 2930 2365 2955
rect 3090 2955 3110 2975
rect 3145 2955 3165 2975
rect 3275 2955 3295 2975
rect 3455 2955 3475 2975
rect 3635 2955 3655 2975
rect 3815 2955 3835 2975
rect 3995 2955 4015 2975
rect 4175 2955 4195 2975
rect 4355 2955 4375 2975
rect 4535 2955 4555 2975
rect 4715 2955 4735 2975
rect 4845 2955 4865 2975
rect 4895 2955 4915 2975
rect 11290 3130 11310 3150
rect 11410 3130 11430 3150
rect 11530 3130 11550 3150
rect 11650 3130 11670 3150
rect 11770 3130 11790 3150
rect 11831 3130 11849 3150
rect 11890 3130 11910 3150
rect 12010 3130 12030 3150
rect 12130 3130 12150 3150
rect 12250 3130 12270 3150
rect 12370 3130 12390 3150
rect 12490 3130 12510 3150
rect 26350 3600 26370 3620
rect 26470 3600 26490 3620
rect 26590 3600 26610 3620
rect 26710 3600 26730 3620
rect 26830 3600 26850 3620
rect 26950 3600 26970 3620
rect 27070 3600 27090 3620
rect 27190 3600 27210 3620
rect 27310 3600 27330 3620
rect 27430 3600 27450 3620
rect 25590 3185 25610 3205
rect 25910 3185 25930 3205
rect 25990 3185 26010 3205
rect 27955 3265 27975 3285
rect 28065 3265 28085 3285
rect 28175 3265 28195 3285
rect 28285 3265 28305 3285
rect 28395 3265 28415 3285
rect 28505 3265 28525 3285
rect 28615 3265 28635 3285
rect 28725 3265 28745 3285
rect 28835 3265 28855 3285
rect 28945 3265 28965 3285
rect 29055 3265 29075 3285
rect 2340 2870 2365 2895
rect 61 2825 86 2850
rect 734 2825 759 2850
rect 1271 2810 1296 2835
rect 1970 2810 1995 2835
rect 10275 2940 10295 2960
rect 10385 2940 10405 2960
rect 10495 2940 10515 2960
rect 10605 2940 10625 2960
rect 10661 2940 10679 2960
rect 10715 2940 10735 2960
rect 11350 2920 11370 2940
rect 11470 2920 11490 2940
rect 11590 2920 11610 2940
rect 11710 2920 11730 2940
rect 11830 2920 11850 2940
rect 11950 2920 11970 2940
rect 12070 2920 12090 2940
rect 12190 2920 12210 2940
rect 12310 2920 12330 2940
rect 12430 2920 12450 2940
rect 13065 2940 13085 2960
rect 13121 2940 13139 2960
rect 13175 2940 13195 2960
rect 13285 2940 13305 2960
rect 13395 2940 13415 2960
rect 13505 2940 13525 2960
rect 26290 3130 26310 3150
rect 26410 3130 26430 3150
rect 26530 3130 26550 3150
rect 26650 3130 26670 3150
rect 26770 3130 26790 3150
rect 26831 3130 26849 3150
rect 26890 3130 26910 3150
rect 27010 3130 27030 3150
rect 27130 3130 27150 3150
rect 27250 3130 27270 3150
rect 27370 3130 27390 3150
rect 27490 3130 27510 3150
rect 26350 2920 26370 2940
rect 26470 2920 26490 2940
rect 26590 2920 26610 2940
rect 26710 2920 26730 2940
rect 26830 2920 26850 2940
rect 26950 2920 26970 2940
rect 27070 2920 27090 2940
rect 27190 2920 27210 2940
rect 27310 2920 27330 2940
rect 27430 2920 27450 2940
rect 61 2765 86 2790
rect 734 2765 759 2790
rect 3005 2785 3025 2805
rect 3185 2785 3205 2805
rect 3365 2785 3385 2805
rect 3545 2785 3565 2805
rect 3725 2785 3745 2805
rect 3905 2785 3925 2805
rect 4085 2785 4105 2805
rect 4265 2785 4285 2805
rect 4445 2785 4465 2805
rect 4625 2785 4645 2805
rect 4805 2785 4825 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 3365 2725 3385 2745
rect 3545 2725 3565 2745
rect 3725 2725 3745 2745
rect 3905 2725 3925 2745
rect 4085 2725 4105 2745
rect 4265 2725 4285 2745
rect 4445 2725 4465 2745
rect 4625 2725 4645 2745
rect 4805 2725 4825 2745
rect 10220 2680 10240 2700
rect 10330 2680 10350 2700
rect 10440 2680 10460 2700
rect 10550 2680 10570 2700
rect 10660 2680 10680 2700
rect 10770 2680 10790 2700
rect 13010 2680 13030 2700
rect 13120 2680 13140 2700
rect 13230 2680 13250 2700
rect 13340 2680 13360 2700
rect 13450 2680 13470 2700
rect 13560 2680 13580 2700
rect 11290 2450 11310 2470
rect 11410 2450 11430 2470
rect 11530 2450 11550 2470
rect 11650 2450 11670 2470
rect 11770 2450 11790 2470
rect 11831 2450 11849 2470
rect 11890 2450 11910 2470
rect 12010 2450 12030 2470
rect 12130 2450 12150 2470
rect 12250 2450 12270 2470
rect 12370 2450 12390 2470
rect 12490 2450 12510 2470
rect 24745 2645 24765 2665
rect 24855 2645 24875 2665
rect 24965 2645 24985 2665
rect 25075 2645 25095 2665
rect 25185 2645 25205 2665
rect 25295 2645 25315 2665
rect 25405 2645 25425 2665
rect 25515 2645 25535 2665
rect 25625 2645 25645 2665
rect 25735 2645 25755 2665
rect 25845 2645 25865 2665
rect 3275 2355 3295 2375
rect 3365 2350 3385 2370
rect 3455 2355 3475 2375
rect 3815 2355 3835 2375
rect 3895 2355 3915 2375
rect 3995 2355 4015 2375
rect 4175 2355 4195 2375
rect 10275 2410 10295 2430
rect 10385 2410 10405 2430
rect 10495 2410 10515 2430
rect 10605 2410 10625 2430
rect 10715 2410 10735 2430
rect 13065 2410 13085 2430
rect 13175 2410 13195 2430
rect 13285 2410 13305 2430
rect 13395 2410 13415 2430
rect 13505 2410 13525 2430
rect 24800 2475 24820 2495
rect 24910 2475 24930 2495
rect 25020 2475 25040 2495
rect 25130 2475 25150 2495
rect 25240 2475 25260 2495
rect 25350 2475 25370 2495
rect 25460 2475 25480 2495
rect 25570 2475 25590 2495
rect 25680 2475 25700 2495
rect 25790 2475 25810 2495
rect 28010 2895 28030 2915
rect 28066 2895 28084 2915
rect 28120 2895 28140 2915
rect 28230 2895 28250 2915
rect 28340 2895 28360 2915
rect 28450 2895 28470 2915
rect 28560 2895 28580 2915
rect 28670 2895 28690 2915
rect 28780 2895 28800 2915
rect 28890 2895 28910 2915
rect 29000 2895 29020 2915
rect 27955 2645 27975 2665
rect 28065 2645 28085 2665
rect 28175 2645 28195 2665
rect 28285 2645 28305 2665
rect 28395 2645 28415 2665
rect 28505 2645 28525 2665
rect 28615 2645 28635 2665
rect 28725 2645 28745 2665
rect 28835 2645 28855 2665
rect 28945 2645 28965 2665
rect 29055 2645 29075 2665
rect 26290 2450 26310 2470
rect 26410 2450 26430 2470
rect 26530 2450 26550 2470
rect 26650 2450 26670 2470
rect 26770 2450 26790 2470
rect 26831 2450 26849 2470
rect 26890 2450 26910 2470
rect 27010 2450 27030 2470
rect 27130 2450 27150 2470
rect 27250 2450 27270 2470
rect 27370 2450 27390 2470
rect 27490 2450 27510 2470
rect 28010 2475 28030 2495
rect 28120 2475 28140 2495
rect 28230 2475 28250 2495
rect 28340 2475 28360 2495
rect 28450 2475 28470 2495
rect 28560 2475 28580 2495
rect 28670 2475 28690 2495
rect 28780 2475 28800 2495
rect 28890 2475 28910 2495
rect 29000 2475 29020 2495
rect 25821 2415 25839 2435
rect 27981 2415 27999 2435
rect 4535 2355 4555 2375
rect 4715 2355 4735 2375
rect 10775 2365 10795 2385
rect 13035 2350 13055 2370
rect 24810 2350 24835 2375
rect 25645 2350 25670 2375
rect 28150 2350 28175 2375
rect 28985 2350 29010 2375
rect 3635 2310 3655 2330
rect 4355 2310 4375 2330
rect 3455 2265 3475 2285
rect 4535 2265 4555 2285
rect 10275 2290 10295 2310
rect 10385 2290 10405 2310
rect 10495 2290 10515 2310
rect 10605 2290 10625 2310
rect 10715 2290 10735 2310
rect 13065 2290 13085 2310
rect 13175 2290 13195 2310
rect 13285 2290 13305 2310
rect 13395 2290 13415 2310
rect 13505 2290 13525 2310
rect 24810 2290 24835 2315
rect 25645 2290 25670 2315
rect 28150 2290 28175 2315
rect 28985 2290 29010 2315
rect 2755 2070 2775 2090
rect 2875 2070 2895 2090
rect 2995 2070 3015 2090
rect 3115 2070 3135 2090
rect 3235 2070 3255 2090
rect 3355 2070 3375 2090
rect 3475 2070 3495 2090
rect 3595 2070 3615 2090
rect 3715 2070 3735 2090
rect 3835 2070 3855 2090
rect 3995 2070 4015 2090
rect 4155 2070 4175 2090
rect 4275 2070 4295 2090
rect 4395 2070 4415 2090
rect 4515 2070 4535 2090
rect 4635 2070 4655 2090
rect 4755 2070 4775 2090
rect 4875 2070 4895 2090
rect 4995 2070 5015 2090
rect 5115 2070 5135 2090
rect 5235 2070 5255 2090
rect 2630 2025 2650 2045
rect -35 1695 -15 1715
rect 2815 2025 2835 2045
rect 3175 2025 3195 2045
rect 3535 2025 3555 2045
rect 3895 2025 3915 2045
rect 4095 2025 4115 2045
rect 4455 2025 4475 2045
rect 4815 2025 4835 2045
rect 5175 2025 5195 2045
rect 9795 1975 9820 2000
rect 9855 1975 9880 2000
rect 9915 1975 9940 2000
rect 9975 1975 10000 2000
rect 11340 2155 11360 2175
rect 11450 2155 11470 2175
rect 11560 2155 11580 2175
rect 11670 2155 11690 2175
rect 11780 2155 11800 2175
rect 11836 2155 11854 2175
rect 11890 2155 11910 2175
rect 12000 2155 12020 2175
rect 12110 2155 12130 2175
rect 12220 2155 12240 2175
rect 12330 2155 12350 2175
rect 12440 2155 12460 2175
rect 25821 2255 25839 2275
rect 27981 2255 27999 2275
rect 13800 1975 13825 2000
rect 10220 1920 10238 1940
rect 10330 1920 10348 1940
rect 10440 1920 10458 1940
rect 10550 1920 10568 1940
rect 10660 1920 10678 1940
rect 10770 1920 10788 1940
rect 11395 1935 11415 1955
rect 11505 1935 11525 1955
rect 11615 1935 11635 1955
rect 11725 1935 11745 1955
rect 11835 1935 11855 1955
rect 11945 1935 11965 1955
rect 12055 1935 12075 1955
rect 12165 1935 12185 1955
rect 12275 1935 12295 1955
rect 12385 1935 12405 1955
rect 13860 1975 13885 2000
rect 13920 1975 13945 2000
rect 24800 2195 24820 2215
rect 24910 2195 24930 2215
rect 25020 2195 25040 2215
rect 25130 2195 25150 2215
rect 25240 2195 25260 2215
rect 25350 2195 25370 2215
rect 25460 2195 25480 2215
rect 25570 2195 25590 2215
rect 25680 2195 25700 2215
rect 25790 2195 25810 2215
rect 28010 2195 28030 2215
rect 28120 2195 28140 2215
rect 28230 2195 28250 2215
rect 28340 2195 28360 2215
rect 28450 2195 28470 2215
rect 28560 2195 28580 2215
rect 28670 2195 28690 2215
rect 28780 2195 28800 2215
rect 28890 2195 28910 2215
rect 29000 2195 29020 2215
rect 26340 2155 26360 2175
rect 26450 2155 26470 2175
rect 26560 2155 26580 2175
rect 26670 2155 26690 2175
rect 26780 2155 26800 2175
rect 26890 2155 26910 2175
rect 27000 2155 27020 2175
rect 27110 2155 27130 2175
rect 27220 2155 27240 2175
rect 27330 2155 27350 2175
rect 27440 2155 27460 2175
rect 13980 1975 14005 2000
rect 24745 1975 24763 1995
rect 24855 1975 24873 1995
rect 24965 1975 24983 1995
rect 25075 1975 25093 1995
rect 25185 1975 25203 1995
rect 25295 1975 25313 1995
rect 25405 1975 25423 1995
rect 25515 1975 25533 1995
rect 25625 1975 25643 1995
rect 25735 1975 25753 1995
rect 25845 1975 25863 1995
rect 27957 1975 27975 1995
rect 28067 1975 28085 1995
rect 28177 1975 28195 1995
rect 28287 1975 28305 1995
rect 28397 1975 28415 1995
rect 28507 1975 28525 1995
rect 28617 1975 28635 1995
rect 28727 1975 28745 1995
rect 28837 1975 28855 1995
rect 28947 1975 28965 1995
rect 29057 1975 29075 1995
rect 13012 1920 13030 1940
rect 13122 1920 13140 1940
rect 13232 1920 13250 1940
rect 13342 1920 13360 1940
rect 13452 1920 13470 1940
rect 13562 1920 13580 1940
rect 26395 1935 26415 1955
rect 26505 1935 26525 1955
rect 26615 1935 26635 1955
rect 26725 1935 26745 1955
rect 26835 1935 26855 1955
rect 26945 1935 26965 1955
rect 27055 1935 27075 1955
rect 27165 1935 27185 1955
rect 27275 1935 27295 1955
rect 27385 1935 27405 1955
rect 2575 1855 2595 1875
rect 2630 1855 2650 1875
rect 2685 1855 2705 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3055 1855 3075 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3415 1855 3435 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3775 1855 3795 1875
rect 3865 1855 3885 1875
rect 4125 1855 4145 1875
rect 4215 1855 4235 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4575 1855 4595 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 4935 1855 4955 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 28055 1880 28075 1900
rect 28165 1880 28185 1900
rect 28275 1880 28295 1900
rect 3055 1795 3075 1815
rect 3415 1795 3435 1815
rect 3775 1795 3795 1815
rect 4215 1795 4235 1815
rect 4575 1795 4595 1815
rect 4935 1795 4955 1815
rect 3235 1735 3255 1755
rect 3295 1735 3315 1755
rect 3535 1735 3555 1755
rect 3775 1735 3795 1755
rect 4215 1735 4235 1755
rect 4455 1735 4475 1755
rect 4695 1735 4715 1755
rect 4755 1735 4775 1755
rect 11095 1735 11115 1755
rect 11200 1750 11220 1770
rect 3175 1690 3195 1710
rect 3415 1690 3435 1710
rect 3655 1690 3675 1710
rect 4335 1690 4355 1710
rect 4575 1690 4595 1710
rect 4815 1690 4835 1710
rect 10265 1680 10285 1700
rect 10465 1680 10485 1700
rect 10566 1680 10584 1700
rect 10665 1680 10685 1700
rect 3995 1630 4015 1650
rect 11315 1735 11335 1755
rect 11420 1750 11440 1770
rect 11243 1690 11260 1710
rect 11535 1735 11555 1755
rect 11650 1750 11670 1770
rect 11463 1690 11480 1710
rect 11610 1690 11627 1710
rect 12135 1735 12155 1755
rect 12240 1750 12260 1770
rect 11825 1690 11845 1710
rect 11876 1690 11893 1710
rect 11955 1690 11975 1710
rect 12355 1735 12375 1755
rect 12460 1750 12480 1770
rect 12283 1690 12300 1710
rect 12575 1735 12595 1755
rect 12690 1750 12710 1770
rect 12503 1690 12520 1710
rect 12650 1690 12667 1710
rect 26095 1735 26115 1755
rect 26200 1750 26220 1770
rect 13115 1680 13135 1700
rect 13216 1680 13234 1700
rect 13315 1680 13335 1700
rect 13515 1680 13535 1700
rect 3175 1570 3195 1590
rect 9975 1615 10000 1640
rect 4815 1570 4835 1590
rect 3235 1520 3255 1540
rect 3355 1520 3375 1540
rect 3475 1520 3495 1540
rect 3595 1520 3615 1540
rect 3715 1520 3735 1540
rect 4275 1520 4295 1540
rect 4395 1520 4415 1540
rect 4515 1520 4535 1540
rect 4635 1520 4655 1540
rect 4755 1520 4775 1540
rect 2845 1460 2865 1480
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 3925 1460 3945 1480
rect 4065 1460 4085 1480
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 5145 1460 5165 1480
rect 10035 1615 10060 1640
rect 3385 1160 3405 1180
rect 4605 1160 4625 1180
rect 2955 1100 2975 1120
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 3995 1100 4015 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 2915 1015 2935 1035
rect 5120 1015 5140 1035
rect 3005 905 3025 925
rect 3185 905 3205 925
rect 3365 905 3385 925
rect 3545 905 3565 925
rect 3725 905 3745 925
rect 3905 905 3925 925
rect 4085 905 4105 925
rect 4265 905 4285 925
rect 4445 905 4465 925
rect 4625 905 4645 925
rect 4805 905 4825 925
rect 4985 905 5005 925
rect 26315 1735 26335 1755
rect 26420 1750 26440 1770
rect 26243 1690 26260 1710
rect 26535 1735 26555 1755
rect 26650 1750 26670 1770
rect 26463 1690 26480 1710
rect 26610 1690 26627 1710
rect 27135 1735 27155 1755
rect 27240 1750 27260 1770
rect 26825 1690 26845 1710
rect 26876 1690 26893 1710
rect 26955 1690 26975 1710
rect 27355 1735 27375 1755
rect 27460 1750 27480 1770
rect 27283 1690 27300 1710
rect 27575 1735 27595 1755
rect 27690 1750 27710 1770
rect 27503 1690 27520 1710
rect 27650 1690 27667 1710
rect 11112 1470 11129 1490
rect 11315 1470 11335 1490
rect 11535 1470 11555 1490
rect 11830 1470 11850 1490
rect 11880 1470 11900 1490
rect 11928 1470 11945 1490
rect 12152 1470 12169 1490
rect 12355 1470 12375 1490
rect 12575 1470 12595 1490
rect 11155 1410 11175 1430
rect 11260 1410 11280 1430
rect 11370 1410 11390 1430
rect 11480 1410 11500 1430
rect 11590 1410 11610 1430
rect 12195 1410 12215 1430
rect 12300 1410 12320 1430
rect 12410 1410 12430 1430
rect 12520 1410 12540 1430
rect 12630 1410 12650 1430
rect 11325 1210 11345 1230
rect 11435 1210 11455 1230
rect 11545 1210 11565 1230
rect 11655 1210 11675 1230
rect 11765 1210 11785 1230
rect 11820 1210 11840 1230
rect 11875 1210 11895 1230
rect 11985 1210 12005 1230
rect 12095 1210 12115 1230
rect 12205 1210 12225 1230
rect 12315 1210 12335 1230
rect 12425 1210 12445 1230
rect 12535 1210 12555 1230
rect 12605 1225 12625 1245
rect 13740 1615 13765 1640
rect 13800 1615 13825 1640
rect 28071 1655 28091 1675
rect 28125 1660 28145 1680
rect 28220 1660 28240 1680
rect 28020 1605 28040 1625
rect 28310 1605 28330 1625
rect 27976 1545 27996 1565
rect 26112 1470 26129 1490
rect 26315 1470 26335 1490
rect 26535 1470 26555 1490
rect 26830 1470 26850 1490
rect 26880 1470 26900 1490
rect 26928 1470 26945 1490
rect 27152 1470 27169 1490
rect 27355 1470 27375 1490
rect 27575 1470 27595 1490
rect 28070 1545 28090 1565
rect 28354 1545 28374 1565
rect 26155 1410 26175 1430
rect 26260 1410 26280 1430
rect 26370 1410 26390 1430
rect 26480 1410 26500 1430
rect 26590 1410 26610 1430
rect 27195 1410 27215 1430
rect 27300 1410 27320 1430
rect 27410 1410 27430 1430
rect 27520 1410 27540 1430
rect 27630 1410 27650 1430
rect 28033 1325 28053 1345
rect 28297 1325 28317 1345
rect 26325 1250 26345 1270
rect 26435 1250 26455 1270
rect 26545 1250 26565 1270
rect 26655 1250 26675 1270
rect 26765 1250 26785 1270
rect 26820 1250 26840 1270
rect 26875 1250 26895 1270
rect 26985 1250 27005 1270
rect 27095 1250 27115 1270
rect 27205 1250 27225 1270
rect 27315 1250 27335 1270
rect 27425 1250 27445 1270
rect 27535 1250 27555 1270
rect 27605 1265 27625 1285
rect 27955 1265 27975 1285
rect 28070 1265 28090 1285
rect 28260 1265 28280 1285
rect 28375 1265 28395 1285
rect 10365 910 10385 930
rect 10565 910 10585 930
rect 11175 890 11195 910
rect 11270 890 11290 910
rect 11380 890 11400 910
rect 11490 890 11510 910
rect 11600 890 11620 910
rect 11710 890 11730 910
rect 11820 890 11840 910
rect 11930 890 11950 910
rect 12040 890 12060 910
rect 12150 890 12170 910
rect 12260 890 12280 910
rect 12370 890 12390 910
rect 12480 890 12500 910
rect 12630 890 12650 910
rect 13215 910 13235 930
rect 13415 910 13435 930
rect 28110 1205 28130 1225
rect 28165 1205 28185 1225
rect 28220 1205 28240 1225
rect 26175 930 26195 950
rect 26270 930 26290 950
rect 26380 930 26400 950
rect 26490 930 26510 950
rect 26600 930 26620 950
rect 26710 930 26730 950
rect 26820 930 26840 950
rect 26930 930 26950 950
rect 27040 930 27060 950
rect 27150 930 27170 950
rect 27260 930 27280 950
rect 27370 930 27390 950
rect 27480 930 27500 950
rect 27630 930 27650 950
rect 11315 770 11335 790
rect 3140 735 3160 755
rect 3275 735 3295 755
rect 3455 735 3475 755
rect 3635 735 3655 755
rect 3815 735 3835 755
rect 3995 735 4015 755
rect 4175 735 4195 755
rect 4355 735 4375 755
rect 4535 735 4555 755
rect 4715 735 4735 755
rect 4895 735 4915 755
rect 11385 770 11405 790
rect 11455 770 11475 790
rect 11945 775 11965 795
rect 12055 775 12075 795
rect 12165 775 12185 795
rect 12275 775 12295 795
rect 12385 775 12405 795
rect 12495 775 12515 795
rect 12000 655 12020 675
rect 12110 655 12130 675
rect 12220 655 12240 675
rect 12330 655 12350 675
rect 12440 655 12460 675
rect 11350 -1400 11370 -1380
rect 11470 -1400 11490 -1380
rect 11590 -1400 11610 -1380
rect 11710 -1400 11730 -1380
rect 11830 -1400 11850 -1380
rect 11950 -1400 11970 -1380
rect 12070 -1400 12090 -1380
rect 12190 -1400 12210 -1380
rect 12310 -1400 12330 -1380
rect 12430 -1400 12450 -1380
rect 10590 -1815 10610 -1795
rect 10910 -1815 10930 -1795
rect 10990 -1815 11010 -1795
rect 11290 -1870 11310 -1850
rect 11410 -1870 11430 -1850
rect 11530 -1870 11550 -1850
rect 11650 -1870 11670 -1850
rect 11770 -1870 11790 -1850
rect 11831 -1870 11849 -1850
rect 11890 -1870 11910 -1850
rect 12010 -1870 12030 -1850
rect 12130 -1870 12150 -1850
rect 12250 -1870 12270 -1850
rect 12370 -1870 12390 -1850
rect 12490 -1870 12510 -1850
rect 12960 -1990 12980 -1970
rect 13070 -1990 13090 -1970
rect 13180 -1990 13200 -1970
rect 13290 -1990 13310 -1970
rect 13400 -1990 13420 -1970
rect 13510 -1990 13530 -1970
rect 13620 -1990 13640 -1970
rect 13730 -1990 13750 -1970
rect 13840 -1990 13860 -1970
rect 13950 -1990 13970 -1970
rect 14060 -1990 14080 -1970
rect 11350 -2080 11370 -2060
rect 11470 -2080 11490 -2060
rect 11590 -2080 11610 -2060
rect 11710 -2080 11730 -2060
rect 11830 -2080 11850 -2060
rect 11950 -2080 11970 -2060
rect 12070 -2080 12090 -2060
rect 12190 -2080 12210 -2060
rect 12310 -2080 12330 -2060
rect 12430 -2080 12450 -2060
rect 13015 -2360 13035 -2340
rect 13071 -2360 13089 -2340
rect 13125 -2360 13145 -2340
rect 13235 -2360 13255 -2340
rect 13345 -2360 13365 -2340
rect 13455 -2360 13475 -2340
rect 13565 -2360 13585 -2340
rect 13675 -2360 13695 -2340
rect 13785 -2360 13805 -2340
rect 13895 -2360 13915 -2340
rect 14005 -2360 14025 -2340
rect 12960 -2420 12980 -2400
rect 13070 -2420 13090 -2400
rect 13180 -2420 13200 -2400
rect 13290 -2420 13310 -2400
rect 13400 -2420 13420 -2400
rect 13510 -2420 13530 -2400
rect 13620 -2420 13640 -2400
rect 13730 -2420 13750 -2400
rect 13840 -2420 13860 -2400
rect 13950 -2420 13970 -2400
rect 14060 -2420 14080 -2400
rect 11290 -2550 11310 -2530
rect 11410 -2550 11430 -2530
rect 11530 -2550 11550 -2530
rect 11650 -2550 11670 -2530
rect 11770 -2550 11790 -2530
rect 11831 -2550 11849 -2530
rect 11890 -2550 11910 -2530
rect 12010 -2550 12030 -2530
rect 12130 -2550 12150 -2530
rect 12250 -2550 12270 -2530
rect 12370 -2550 12390 -2530
rect 12490 -2550 12510 -2530
rect 13015 -2590 13035 -2570
rect 13125 -2590 13145 -2570
rect 13235 -2590 13255 -2570
rect 13345 -2590 13365 -2570
rect 13455 -2590 13475 -2570
rect 13565 -2590 13585 -2570
rect 13675 -2590 13695 -2570
rect 13785 -2590 13805 -2570
rect 13895 -2590 13915 -2570
rect 14005 -2590 14025 -2570
rect 12985 -2650 13005 -2630
rect 13015 -2710 13035 -2690
rect 13125 -2710 13145 -2690
rect 13235 -2710 13255 -2690
rect 13345 -2710 13365 -2690
rect 13455 -2710 13475 -2690
rect 13565 -2710 13585 -2690
rect 13675 -2710 13695 -2690
rect 13785 -2710 13805 -2690
rect 13895 -2710 13915 -2690
rect 14005 -2710 14025 -2690
rect 11340 -2845 11360 -2825
rect 11450 -2845 11470 -2825
rect 11560 -2845 11580 -2825
rect 11670 -2845 11690 -2825
rect 11780 -2845 11800 -2825
rect 11890 -2845 11910 -2825
rect 12000 -2845 12020 -2825
rect 12110 -2845 12130 -2825
rect 12220 -2845 12240 -2825
rect 12330 -2845 12350 -2825
rect 12440 -2845 12460 -2825
rect 12962 -2930 12980 -2910
rect 13072 -2930 13090 -2910
rect 13182 -2930 13200 -2910
rect 13292 -2930 13310 -2910
rect 13402 -2930 13420 -2910
rect 13512 -2930 13530 -2910
rect 13622 -2930 13640 -2910
rect 13732 -2930 13750 -2910
rect 13842 -2930 13860 -2910
rect 13952 -2930 13970 -2910
rect 14062 -2930 14080 -2910
rect 13005 -2990 13025 -2970
rect 13106 -2990 13124 -2970
rect 13205 -2990 13225 -2970
rect 13405 -2990 13425 -2970
rect 13605 -2990 13625 -2970
rect 13805 -2990 13825 -2970
rect 14005 -2990 14025 -2970
rect 11395 -3065 11415 -3045
rect 11505 -3065 11525 -3045
rect 11615 -3065 11635 -3045
rect 11725 -3065 11745 -3045
rect 11835 -3065 11855 -3045
rect 11945 -3065 11965 -3045
rect 12055 -3065 12075 -3045
rect 12165 -3065 12185 -3045
rect 12275 -3065 12295 -3045
rect 12385 -3065 12405 -3045
rect 11095 -3265 11115 -3245
rect 11200 -3250 11220 -3230
rect 11315 -3265 11335 -3245
rect 11420 -3250 11440 -3230
rect 11243 -3310 11260 -3290
rect 11535 -3265 11555 -3245
rect 11650 -3250 11670 -3230
rect 11463 -3310 11480 -3290
rect 11610 -3310 11627 -3290
rect 12135 -3265 12155 -3245
rect 12240 -3250 12260 -3230
rect 11825 -3310 11845 -3290
rect 11876 -3310 11893 -3290
rect 11955 -3310 11975 -3290
rect 12355 -3265 12375 -3245
rect 12460 -3250 12480 -3230
rect 12283 -3310 12300 -3290
rect 12575 -3265 12595 -3245
rect 12690 -3250 12710 -3230
rect 12503 -3310 12520 -3290
rect 12650 -3310 12667 -3290
rect 13105 -3340 13125 -3320
rect 13305 -3340 13325 -3320
rect 13505 -3340 13525 -3320
rect 13705 -3340 13725 -3320
rect 13905 -3340 13925 -3320
rect 11112 -3530 11129 -3510
rect 11315 -3530 11335 -3510
rect 11535 -3530 11555 -3510
rect 11830 -3530 11850 -3510
rect 11880 -3530 11900 -3510
rect 11928 -3530 11945 -3510
rect 12152 -3530 12169 -3510
rect 12355 -3530 12375 -3510
rect 12575 -3530 12595 -3510
rect 11155 -3590 11175 -3570
rect 11260 -3590 11280 -3570
rect 11370 -3590 11390 -3570
rect 11480 -3590 11500 -3570
rect 11590 -3590 11610 -3570
rect 12195 -3590 12215 -3570
rect 12300 -3590 12320 -3570
rect 12410 -3590 12430 -3570
rect 12520 -3590 12540 -3570
rect 12630 -3590 12650 -3570
rect 11325 -3790 11345 -3770
rect 11435 -3790 11455 -3770
rect 11545 -3790 11565 -3770
rect 11655 -3790 11675 -3770
rect 11765 -3790 11785 -3770
rect 11820 -3790 11840 -3770
rect 11875 -3790 11895 -3770
rect 11985 -3790 12005 -3770
rect 12095 -3790 12115 -3770
rect 12205 -3790 12225 -3770
rect 12315 -3790 12335 -3770
rect 12425 -3790 12445 -3770
rect 12535 -3790 12555 -3770
rect 12605 -3775 12625 -3755
rect 11175 -4110 11195 -4090
rect 11270 -4110 11290 -4090
rect 11380 -4110 11400 -4090
rect 11490 -4110 11510 -4090
rect 11600 -4110 11620 -4090
rect 11710 -4110 11730 -4090
rect 11820 -4110 11840 -4090
rect 11930 -4110 11950 -4090
rect 12040 -4110 12060 -4090
rect 12150 -4110 12170 -4090
rect 12260 -4110 12280 -4090
rect 12370 -4110 12390 -4090
rect 12480 -4110 12500 -4090
rect 12630 -4110 12650 -4090
<< metal1 >>
rect 11632 9055 11668 9060
rect 11632 9025 11635 9055
rect 11665 9025 11668 9055
rect 11632 9020 11668 9025
rect 11752 9055 11788 9060
rect 11752 9025 11755 9055
rect 11785 9025 11788 9055
rect 11752 9020 11788 9025
rect 11872 9055 11908 9060
rect 11872 9025 11875 9055
rect 11905 9025 11908 9055
rect 11872 9020 11908 9025
rect 12080 9055 12120 9060
rect 12080 9025 12085 9055
rect 12115 9025 12120 9055
rect 12080 9020 12120 9025
rect 11570 9010 11610 9015
rect 11200 8995 11240 9000
rect 11200 8965 11205 8995
rect 11235 8965 11240 8995
rect 11200 8960 11240 8965
rect 11460 8995 11500 9000
rect 11460 8965 11465 8995
rect 11495 8965 11500 8995
rect 11570 8980 11575 9010
rect 11605 8980 11610 9010
rect 11570 8975 11610 8980
rect 11690 9010 11730 9015
rect 11690 8980 11695 9010
rect 11725 8980 11730 9010
rect 11690 8975 11730 8980
rect 11810 9010 11850 9015
rect 11810 8980 11815 9010
rect 11845 8980 11850 9010
rect 11810 8975 11850 8980
rect 11930 9010 11970 9015
rect 11930 8980 11935 9010
rect 11965 8980 11970 9010
rect 12090 8990 12110 9020
rect 11930 8975 11970 8980
rect 12080 8985 12120 8990
rect 11460 8960 11500 8965
rect 12080 8955 12085 8985
rect 12115 8955 12120 8985
rect 12080 8950 12120 8955
rect 12200 8985 12240 8990
rect 12200 8955 12205 8985
rect 12235 8955 12240 8985
rect 12200 8950 12240 8955
rect 12320 8985 12360 8990
rect 12320 8955 12325 8985
rect 12355 8955 12360 8985
rect 12320 8950 12360 8955
rect 12440 8985 12480 8990
rect 12440 8955 12445 8985
rect 12475 8955 12480 8985
rect 12440 8950 12480 8955
rect 12560 8985 12600 8990
rect 12560 8955 12565 8985
rect 12595 8955 12600 8985
rect 12560 8950 12600 8955
rect 11330 8860 11370 8865
rect 11330 8830 11335 8860
rect 11365 8830 11370 8860
rect 11330 8825 11370 8830
rect 11750 8855 11790 8860
rect 11750 8825 11755 8855
rect 11785 8825 11790 8855
rect 11340 8770 11360 8825
rect 11750 8820 11790 8825
rect 12140 8855 12180 8860
rect 12140 8825 12145 8855
rect 12175 8825 12180 8855
rect 12140 8820 12180 8825
rect 12203 8850 12237 8860
rect 12203 8830 12211 8850
rect 12229 8830 12237 8850
rect 12203 8820 12237 8830
rect 12260 8855 12300 8860
rect 12260 8825 12265 8855
rect 12295 8825 12300 8855
rect 12260 8820 12300 8825
rect 12380 8855 12420 8860
rect 12380 8825 12385 8855
rect 12415 8825 12420 8855
rect 12380 8820 12420 8825
rect 12500 8855 12540 8860
rect 12500 8825 12505 8855
rect 12535 8825 12540 8855
rect 12500 8820 12540 8825
rect 12210 8770 12230 8820
rect 11330 8765 11370 8770
rect 11330 8735 11335 8765
rect 11365 8735 11370 8765
rect 11330 8730 11370 8735
rect 12200 8765 12240 8770
rect 12200 8735 12205 8765
rect 12235 8735 12240 8765
rect 12200 8730 12240 8735
rect 11340 8625 11380 8630
rect 11340 8595 11345 8625
rect 11375 8595 11380 8625
rect 11340 8590 11380 8595
rect 11460 8625 11500 8630
rect 11460 8595 11465 8625
rect 11495 8595 11500 8625
rect 11460 8590 11500 8595
rect 11580 8625 11620 8630
rect 11580 8595 11585 8625
rect 11615 8595 11620 8625
rect 11580 8590 11620 8595
rect 11700 8625 11740 8630
rect 11700 8595 11705 8625
rect 11735 8595 11740 8625
rect 11700 8590 11740 8595
rect 11820 8625 11860 8630
rect 11820 8595 11825 8625
rect 11855 8595 11860 8625
rect 11820 8590 11860 8595
rect 11940 8625 11980 8630
rect 11940 8595 11945 8625
rect 11975 8595 11980 8625
rect 11940 8590 11980 8595
rect 12060 8625 12100 8630
rect 12060 8595 12065 8625
rect 12095 8595 12100 8625
rect 12060 8590 12100 8595
rect 12180 8625 12220 8630
rect 12180 8595 12185 8625
rect 12215 8595 12220 8625
rect 12180 8590 12220 8595
rect 12300 8625 12340 8630
rect 12300 8595 12305 8625
rect 12335 8595 12340 8625
rect 12300 8590 12340 8595
rect 12420 8625 12460 8630
rect 12420 8595 12425 8625
rect 12455 8595 12460 8625
rect 12420 8590 12460 8595
rect 18840 8625 18880 8630
rect 18840 8595 18845 8625
rect 18875 8595 18880 8625
rect 18840 8590 18880 8595
rect 18960 8625 19000 8630
rect 18960 8595 18965 8625
rect 18995 8595 19000 8625
rect 18960 8590 19000 8595
rect 19080 8625 19120 8630
rect 19080 8595 19085 8625
rect 19115 8595 19120 8625
rect 19080 8590 19120 8595
rect 19200 8625 19240 8630
rect 19200 8595 19205 8625
rect 19235 8595 19240 8625
rect 19200 8590 19240 8595
rect 19320 8625 19360 8630
rect 19320 8595 19325 8625
rect 19355 8595 19360 8625
rect 19320 8590 19360 8595
rect 19440 8625 19480 8630
rect 19440 8595 19445 8625
rect 19475 8595 19480 8625
rect 19440 8590 19480 8595
rect 19560 8625 19600 8630
rect 19560 8595 19565 8625
rect 19595 8595 19600 8625
rect 19560 8590 19600 8595
rect 19680 8625 19720 8630
rect 19680 8595 19685 8625
rect 19715 8595 19720 8625
rect 19680 8590 19720 8595
rect 19800 8625 19840 8630
rect 19800 8595 19805 8625
rect 19835 8595 19840 8625
rect 19800 8590 19840 8595
rect 19920 8625 19960 8630
rect 19920 8595 19925 8625
rect 19955 8595 19960 8625
rect 19920 8590 19960 8595
rect 12950 8290 12990 8295
rect 12950 8260 12955 8290
rect 12985 8260 12990 8290
rect 12950 8255 12990 8260
rect 13060 8290 13100 8295
rect 13060 8260 13065 8290
rect 13095 8260 13100 8290
rect 13060 8255 13100 8260
rect 13170 8290 13210 8295
rect 13170 8260 13175 8290
rect 13205 8260 13210 8290
rect 13170 8255 13210 8260
rect 13280 8290 13320 8295
rect 13280 8260 13285 8290
rect 13315 8260 13320 8290
rect 13280 8255 13320 8260
rect 13390 8290 13430 8295
rect 13390 8260 13395 8290
rect 13425 8260 13430 8290
rect 13390 8255 13430 8260
rect 13500 8290 13540 8295
rect 13500 8260 13505 8290
rect 13535 8260 13540 8290
rect 13500 8255 13540 8260
rect 13610 8290 13650 8295
rect 13610 8260 13615 8290
rect 13645 8260 13650 8290
rect 13610 8255 13650 8260
rect 13720 8290 13760 8295
rect 13720 8260 13725 8290
rect 13755 8260 13760 8290
rect 13720 8255 13760 8260
rect 13830 8290 13870 8295
rect 13830 8260 13835 8290
rect 13865 8260 13870 8290
rect 13830 8255 13870 8260
rect 13940 8290 13980 8295
rect 13940 8260 13945 8290
rect 13975 8260 13980 8290
rect 13940 8255 13980 8260
rect 14050 8290 14090 8295
rect 14050 8260 14055 8290
rect 14085 8260 14090 8290
rect 14050 8255 14090 8260
rect 20445 8290 20485 8295
rect 20445 8260 20450 8290
rect 20480 8260 20485 8290
rect 20445 8255 20485 8260
rect 20555 8290 20595 8295
rect 20555 8260 20560 8290
rect 20590 8260 20595 8290
rect 20555 8255 20595 8260
rect 20665 8290 20705 8295
rect 20665 8260 20670 8290
rect 20700 8260 20705 8290
rect 20665 8255 20705 8260
rect 20775 8290 20815 8295
rect 20775 8260 20780 8290
rect 20810 8260 20815 8290
rect 20775 8255 20815 8260
rect 20885 8290 20925 8295
rect 20885 8260 20890 8290
rect 20920 8260 20925 8290
rect 20885 8255 20925 8260
rect 20995 8290 21035 8295
rect 20995 8260 21000 8290
rect 21030 8260 21035 8290
rect 20995 8255 21035 8260
rect 21105 8290 21145 8295
rect 21105 8260 21110 8290
rect 21140 8260 21145 8290
rect 21105 8255 21145 8260
rect 21215 8290 21255 8295
rect 21215 8260 21220 8290
rect 21250 8260 21255 8290
rect 21215 8255 21255 8260
rect 21325 8290 21365 8295
rect 21325 8260 21330 8290
rect 21360 8260 21365 8290
rect 21325 8255 21365 8260
rect 21435 8290 21475 8295
rect 21435 8260 21440 8290
rect 21470 8260 21475 8290
rect 21435 8255 21475 8260
rect 21545 8290 21585 8295
rect 21545 8260 21550 8290
rect 21580 8260 21585 8290
rect 21545 8255 21585 8260
rect 10580 8210 10620 8215
rect 10580 8180 10585 8210
rect 10615 8180 10620 8210
rect 10580 8175 10620 8180
rect 10905 8205 10940 8215
rect 10905 8185 10910 8205
rect 10930 8185 10940 8205
rect 10905 8175 10940 8185
rect 10980 8210 11015 8215
rect 10980 8180 10985 8210
rect 10980 8175 11015 8180
rect 18080 8210 18120 8215
rect 18080 8180 18085 8210
rect 18115 8180 18120 8210
rect 18080 8175 18120 8180
rect 18405 8205 18440 8215
rect 18405 8185 18410 8205
rect 18430 8185 18440 8205
rect 18405 8175 18440 8185
rect 18480 8210 18515 8215
rect 18480 8180 18485 8210
rect 18480 8175 18515 8180
rect 10910 8160 10930 8175
rect 10900 8155 10940 8160
rect 10900 8125 10905 8155
rect 10935 8125 10940 8155
rect 10900 8120 10940 8125
rect 9735 7670 9775 7675
rect 9735 7640 9740 7670
rect 9770 7640 9775 7670
rect 9735 7635 9775 7640
rect 9845 7670 9885 7675
rect 9845 7640 9850 7670
rect 9880 7640 9885 7670
rect 9845 7635 9885 7640
rect 9955 7670 9995 7675
rect 9955 7640 9960 7670
rect 9990 7640 9995 7670
rect 9955 7635 9995 7640
rect 10065 7670 10105 7675
rect 10065 7640 10070 7670
rect 10100 7640 10105 7670
rect 10065 7635 10105 7640
rect 10175 7670 10215 7675
rect 10175 7640 10180 7670
rect 10210 7640 10215 7670
rect 10175 7635 10215 7640
rect 10285 7670 10325 7675
rect 10285 7640 10290 7670
rect 10320 7640 10325 7670
rect 10285 7635 10325 7640
rect 10395 7670 10435 7675
rect 10395 7640 10400 7670
rect 10430 7640 10435 7670
rect 10395 7635 10435 7640
rect 10505 7670 10545 7675
rect 10505 7640 10510 7670
rect 10540 7640 10545 7670
rect 10505 7635 10545 7640
rect 10615 7670 10655 7675
rect 10615 7640 10620 7670
rect 10650 7640 10655 7670
rect 10615 7635 10655 7640
rect 10725 7670 10765 7675
rect 10725 7640 10730 7670
rect 10760 7640 10765 7670
rect 10725 7635 10765 7640
rect 10835 7670 10875 7675
rect 10835 7640 10840 7670
rect 10870 7640 10875 7670
rect 10835 7635 10875 7640
rect 9790 7500 9830 7505
rect 9790 7470 9795 7500
rect 9825 7470 9830 7500
rect 9790 7465 9830 7470
rect 9900 7500 9940 7505
rect 9900 7470 9905 7500
rect 9935 7470 9940 7500
rect 9900 7465 9940 7470
rect 10010 7500 10050 7505
rect 10010 7470 10015 7500
rect 10045 7470 10050 7500
rect 10010 7465 10050 7470
rect 10120 7500 10160 7505
rect 10120 7470 10125 7500
rect 10155 7470 10160 7500
rect 10120 7465 10160 7470
rect 10230 7500 10270 7505
rect 10230 7470 10235 7500
rect 10265 7470 10270 7500
rect 10230 7465 10270 7470
rect 10340 7500 10380 7505
rect 10340 7470 10345 7500
rect 10375 7470 10380 7500
rect 10340 7465 10380 7470
rect 10450 7500 10490 7505
rect 10450 7470 10455 7500
rect 10485 7470 10490 7500
rect 10450 7465 10490 7470
rect 10560 7500 10600 7505
rect 10560 7470 10565 7500
rect 10595 7470 10600 7500
rect 10560 7465 10600 7470
rect 10670 7500 10710 7505
rect 10670 7470 10675 7500
rect 10705 7470 10710 7500
rect 10670 7465 10710 7470
rect 10780 7500 10820 7505
rect 10780 7470 10785 7500
rect 10815 7470 10820 7500
rect 10990 7480 11010 8175
rect 18410 8160 18430 8175
rect 11280 8150 11320 8160
rect 11280 8130 11290 8150
rect 11310 8130 11320 8150
rect 11280 8120 11320 8130
rect 11400 8150 11440 8160
rect 11400 8130 11410 8150
rect 11430 8130 11440 8150
rect 11400 8120 11440 8130
rect 11520 8150 11560 8160
rect 11520 8130 11530 8150
rect 11550 8130 11560 8150
rect 11520 8120 11560 8130
rect 11640 8150 11680 8160
rect 11640 8130 11650 8150
rect 11670 8130 11680 8150
rect 11640 8120 11680 8130
rect 11760 8150 11800 8160
rect 11760 8130 11770 8150
rect 11790 8130 11800 8150
rect 11760 8120 11800 8130
rect 11823 8155 11857 8160
rect 11823 8125 11826 8155
rect 11854 8125 11857 8155
rect 11823 8120 11857 8125
rect 11880 8150 11920 8160
rect 11880 8130 11890 8150
rect 11910 8130 11920 8150
rect 11880 8120 11920 8130
rect 12000 8150 12040 8160
rect 12000 8130 12010 8150
rect 12030 8130 12040 8150
rect 12000 8120 12040 8130
rect 12120 8150 12160 8160
rect 12120 8130 12130 8150
rect 12150 8130 12160 8150
rect 12120 8120 12160 8130
rect 12240 8150 12280 8160
rect 12240 8130 12250 8150
rect 12270 8130 12280 8150
rect 12240 8120 12280 8130
rect 12360 8150 12400 8160
rect 12360 8130 12370 8150
rect 12390 8130 12400 8150
rect 12360 8120 12400 8130
rect 12480 8150 12520 8160
rect 12480 8130 12490 8150
rect 12510 8130 12520 8150
rect 12480 8120 12520 8130
rect 18400 8155 18440 8160
rect 18400 8125 18405 8155
rect 18435 8125 18440 8155
rect 18400 8120 18440 8125
rect 11290 8105 11310 8120
rect 11280 8100 11320 8105
rect 11280 8070 11285 8100
rect 11315 8070 11320 8100
rect 11280 8065 11320 8070
rect 11410 8060 11430 8120
rect 11530 8105 11550 8120
rect 11520 8100 11560 8105
rect 11520 8070 11525 8100
rect 11555 8070 11560 8100
rect 11520 8065 11560 8070
rect 11650 8060 11670 8120
rect 11770 8105 11790 8120
rect 11760 8100 11800 8105
rect 11760 8070 11765 8100
rect 11795 8070 11800 8100
rect 11760 8065 11800 8070
rect 11890 8060 11910 8120
rect 12010 8105 12030 8120
rect 12000 8100 12040 8105
rect 12000 8070 12005 8100
rect 12035 8070 12040 8100
rect 12000 8065 12040 8070
rect 12130 8060 12150 8120
rect 12250 8105 12270 8120
rect 12240 8100 12280 8105
rect 12240 8070 12245 8100
rect 12275 8070 12280 8100
rect 12240 8065 12280 8070
rect 12370 8060 12390 8120
rect 12490 8105 12510 8120
rect 12480 8100 12520 8105
rect 12480 8070 12485 8100
rect 12515 8070 12520 8100
rect 12480 8065 12520 8070
rect 11400 8055 11440 8060
rect 11400 8025 11405 8055
rect 11435 8025 11440 8055
rect 11400 8020 11440 8025
rect 11640 8055 11680 8060
rect 11640 8025 11645 8055
rect 11675 8025 11680 8055
rect 11640 8020 11680 8025
rect 11880 8055 11920 8060
rect 11880 8025 11885 8055
rect 11915 8025 11920 8055
rect 11880 8020 11920 8025
rect 12120 8055 12160 8060
rect 12120 8025 12125 8055
rect 12155 8025 12160 8055
rect 12120 8020 12160 8025
rect 12360 8055 12400 8060
rect 12360 8025 12365 8055
rect 12395 8025 12400 8055
rect 12360 8020 12400 8025
rect 11410 8005 11430 8020
rect 11340 8000 11380 8005
rect 11340 7970 11345 8000
rect 11375 7970 11380 8000
rect 11340 7965 11380 7970
rect 11400 8000 11440 8005
rect 11400 7970 11405 8000
rect 11435 7970 11440 8000
rect 11400 7965 11440 7970
rect 11580 8000 11620 8005
rect 11580 7970 11585 8000
rect 11615 7970 11620 8000
rect 11580 7965 11620 7970
rect 11820 8000 11860 8005
rect 11820 7970 11825 8000
rect 11855 7970 11860 8000
rect 11820 7965 11860 7970
rect 12060 8000 12100 8005
rect 12060 7970 12065 8000
rect 12095 7970 12100 8000
rect 12060 7965 12100 7970
rect 12300 8000 12340 8005
rect 12300 7970 12305 8000
rect 12335 7970 12340 8000
rect 12300 7965 12340 7970
rect 11350 7950 11370 7965
rect 11590 7950 11610 7965
rect 11830 7950 11850 7965
rect 12070 7950 12090 7965
rect 12310 7950 12330 7965
rect 12490 7950 12510 8065
rect 11340 7940 11380 7950
rect 11340 7920 11350 7940
rect 11370 7920 11380 7940
rect 11340 7910 11380 7920
rect 11460 7945 11500 7950
rect 11460 7915 11465 7945
rect 11495 7915 11500 7945
rect 11460 7910 11500 7915
rect 11580 7940 11620 7950
rect 11580 7920 11590 7940
rect 11610 7920 11620 7940
rect 11580 7910 11620 7920
rect 11700 7945 11740 7950
rect 11700 7915 11705 7945
rect 11735 7915 11740 7945
rect 11700 7910 11740 7915
rect 11820 7940 11860 7950
rect 11820 7920 11830 7940
rect 11850 7920 11860 7940
rect 11820 7910 11860 7920
rect 11940 7945 11980 7950
rect 11940 7915 11945 7945
rect 11975 7915 11980 7945
rect 11940 7910 11980 7915
rect 12060 7940 12100 7950
rect 12060 7920 12070 7940
rect 12090 7920 12100 7940
rect 12060 7910 12100 7920
rect 12180 7945 12220 7950
rect 12180 7915 12185 7945
rect 12215 7915 12220 7945
rect 12180 7910 12220 7915
rect 12300 7940 12340 7950
rect 12300 7920 12310 7940
rect 12330 7920 12340 7940
rect 12300 7910 12340 7920
rect 12420 7945 12460 7950
rect 12420 7915 12425 7945
rect 12455 7915 12460 7945
rect 12420 7910 12460 7915
rect 12480 7945 12520 7950
rect 12480 7915 12485 7945
rect 12515 7915 12520 7945
rect 12480 7910 12520 7915
rect 13005 7920 13045 7925
rect 13005 7890 13010 7920
rect 13040 7890 13045 7920
rect 13005 7885 13045 7890
rect 13063 7915 13097 7925
rect 13063 7895 13071 7915
rect 13089 7895 13097 7915
rect 13063 7885 13097 7895
rect 13115 7920 13155 7925
rect 13115 7890 13120 7920
rect 13150 7890 13155 7920
rect 13115 7885 13155 7890
rect 13225 7920 13265 7925
rect 13225 7890 13230 7920
rect 13260 7890 13265 7920
rect 13225 7885 13265 7890
rect 13335 7920 13375 7925
rect 13335 7890 13340 7920
rect 13370 7890 13375 7920
rect 13335 7885 13375 7890
rect 13445 7920 13485 7925
rect 13445 7890 13450 7920
rect 13480 7890 13485 7920
rect 13445 7885 13485 7890
rect 13555 7920 13595 7925
rect 13555 7890 13560 7920
rect 13590 7890 13595 7920
rect 13555 7885 13595 7890
rect 13665 7920 13705 7925
rect 13665 7890 13670 7920
rect 13700 7890 13705 7920
rect 13665 7885 13705 7890
rect 13775 7920 13815 7925
rect 13775 7890 13780 7920
rect 13810 7890 13815 7920
rect 13775 7885 13815 7890
rect 13885 7920 13925 7925
rect 13885 7890 13890 7920
rect 13920 7890 13925 7920
rect 13885 7885 13925 7890
rect 13995 7920 14035 7925
rect 13995 7890 14000 7920
rect 14030 7890 14035 7920
rect 13995 7885 14035 7890
rect 13070 7836 13090 7885
rect 13060 7830 13100 7836
rect 13060 7800 13065 7830
rect 13095 7800 13100 7830
rect 13060 7780 13100 7800
rect 13060 7750 13065 7780
rect 13095 7750 13100 7780
rect 12690 7730 12730 7735
rect 12690 7700 12695 7730
rect 12725 7700 12730 7730
rect 12690 7695 12730 7700
rect 13060 7730 13100 7750
rect 13060 7700 13065 7730
rect 13095 7700 13100 7730
rect 13060 7695 13100 7700
rect 13680 7830 13720 7836
rect 13680 7800 13685 7830
rect 13715 7800 13720 7830
rect 13680 7780 13720 7800
rect 13680 7750 13685 7780
rect 13715 7750 13720 7780
rect 13680 7730 13720 7750
rect 13680 7700 13685 7730
rect 13715 7700 13720 7730
rect 13680 7695 13720 7700
rect 10780 7465 10820 7470
rect 10980 7475 11020 7480
rect 9800 7380 9820 7465
rect 10980 7445 10985 7475
rect 11015 7445 11020 7475
rect 10813 7440 10847 7445
rect 10980 7440 11020 7445
rect 11280 7470 11320 7480
rect 11280 7450 11290 7470
rect 11310 7450 11320 7470
rect 11280 7440 11320 7450
rect 11400 7470 11440 7480
rect 11400 7450 11410 7470
rect 11430 7450 11440 7470
rect 11400 7440 11440 7450
rect 11520 7470 11560 7480
rect 11520 7450 11530 7470
rect 11550 7450 11560 7470
rect 11520 7440 11560 7450
rect 11640 7470 11680 7480
rect 11640 7450 11650 7470
rect 11670 7450 11680 7470
rect 11640 7440 11680 7450
rect 11760 7470 11800 7480
rect 11760 7450 11770 7470
rect 11790 7450 11800 7470
rect 11760 7440 11800 7450
rect 11823 7475 11857 7480
rect 11823 7445 11826 7475
rect 11854 7445 11857 7475
rect 11823 7440 11857 7445
rect 11880 7470 11920 7480
rect 11880 7450 11890 7470
rect 11910 7450 11920 7470
rect 11880 7440 11920 7450
rect 12000 7470 12040 7480
rect 12000 7450 12010 7470
rect 12030 7450 12040 7470
rect 12000 7440 12040 7450
rect 12120 7470 12160 7480
rect 12120 7450 12130 7470
rect 12150 7450 12160 7470
rect 12120 7440 12160 7450
rect 12240 7470 12280 7480
rect 12240 7450 12250 7470
rect 12270 7450 12280 7470
rect 12240 7440 12280 7450
rect 12360 7470 12400 7480
rect 12360 7450 12370 7470
rect 12390 7450 12400 7470
rect 12360 7440 12400 7450
rect 12480 7470 12520 7480
rect 12480 7450 12490 7470
rect 12510 7450 12520 7470
rect 12480 7440 12520 7450
rect 10813 7410 10816 7440
rect 10844 7410 10847 7440
rect 11290 7425 11310 7440
rect 10813 7405 10847 7410
rect 11280 7420 11320 7425
rect 9800 7345 9805 7380
rect 9840 7345 9845 7380
rect 10635 7345 10640 7380
rect 10675 7345 10680 7380
rect 10635 7320 10680 7345
rect 9800 7285 9805 7320
rect 9840 7285 9845 7320
rect 10635 7285 10640 7320
rect 10675 7285 10680 7320
rect 10820 7285 10840 7405
rect 11280 7390 11285 7420
rect 11315 7390 11320 7420
rect 11280 7385 11320 7390
rect 11410 7380 11430 7440
rect 11530 7425 11550 7440
rect 11520 7420 11560 7425
rect 11520 7390 11525 7420
rect 11555 7390 11560 7420
rect 11520 7385 11560 7390
rect 11650 7380 11670 7440
rect 11770 7425 11790 7440
rect 11760 7420 11800 7425
rect 11760 7390 11765 7420
rect 11795 7390 11800 7420
rect 11760 7385 11800 7390
rect 11400 7375 11440 7380
rect 11400 7345 11405 7375
rect 11435 7345 11440 7375
rect 11400 7340 11440 7345
rect 11640 7375 11680 7380
rect 11640 7345 11645 7375
rect 11675 7345 11680 7375
rect 11640 7340 11680 7345
rect 9800 7225 9820 7285
rect 10813 7280 10847 7285
rect 10813 7250 10816 7280
rect 10844 7250 10847 7280
rect 10813 7245 10847 7250
rect 11440 7280 11480 7285
rect 11440 7250 11445 7280
rect 11475 7250 11480 7280
rect 11440 7245 11480 7250
rect 11660 7280 11700 7285
rect 11660 7250 11665 7280
rect 11695 7250 11700 7280
rect 11660 7245 11700 7250
rect 11330 7235 11370 7240
rect 9790 7220 9830 7225
rect 9790 7190 9795 7220
rect 9825 7190 9830 7220
rect 9790 7185 9830 7190
rect 9900 7220 9940 7225
rect 9900 7190 9905 7220
rect 9935 7190 9940 7220
rect 9900 7185 9940 7190
rect 10010 7220 10050 7225
rect 10010 7190 10015 7220
rect 10045 7190 10050 7220
rect 10010 7185 10050 7190
rect 10120 7220 10160 7225
rect 10120 7190 10125 7220
rect 10155 7190 10160 7220
rect 10120 7185 10160 7190
rect 10230 7220 10270 7225
rect 10230 7190 10235 7220
rect 10265 7190 10270 7220
rect 10230 7185 10270 7190
rect 10340 7220 10380 7225
rect 10340 7190 10345 7220
rect 10375 7190 10380 7220
rect 10340 7185 10380 7190
rect 10450 7220 10490 7225
rect 10450 7190 10455 7220
rect 10485 7190 10490 7220
rect 10450 7185 10490 7190
rect 10560 7220 10600 7225
rect 10560 7190 10565 7220
rect 10595 7190 10600 7220
rect 10560 7185 10600 7190
rect 10670 7220 10710 7225
rect 10670 7190 10675 7220
rect 10705 7190 10710 7220
rect 10670 7185 10710 7190
rect 10780 7220 10820 7225
rect 10780 7190 10785 7220
rect 10815 7190 10820 7220
rect 11330 7205 11335 7235
rect 11365 7205 11370 7235
rect 11330 7200 11370 7205
rect 10780 7185 10820 7190
rect 11340 7185 11360 7200
rect 11450 7185 11470 7245
rect 11550 7235 11590 7240
rect 11550 7205 11555 7235
rect 11585 7205 11590 7235
rect 11550 7200 11590 7205
rect 11560 7185 11580 7200
rect 11670 7185 11690 7245
rect 11770 7240 11790 7385
rect 11890 7380 11910 7440
rect 12010 7425 12030 7440
rect 12000 7420 12040 7425
rect 12000 7390 12005 7420
rect 12035 7390 12040 7420
rect 12000 7385 12040 7390
rect 12130 7380 12150 7440
rect 12250 7425 12270 7440
rect 12240 7420 12280 7425
rect 12240 7390 12245 7420
rect 12275 7390 12280 7420
rect 12240 7385 12280 7390
rect 12370 7380 12390 7440
rect 12490 7425 12510 7440
rect 12480 7420 12520 7425
rect 12480 7390 12485 7420
rect 12515 7390 12520 7420
rect 12480 7385 12520 7390
rect 12700 7380 12720 7695
rect 12950 7670 12990 7675
rect 12950 7640 12955 7670
rect 12985 7640 12990 7670
rect 12950 7635 12990 7640
rect 13060 7670 13100 7675
rect 13060 7640 13065 7670
rect 13095 7640 13100 7670
rect 13060 7635 13100 7640
rect 13170 7670 13210 7675
rect 13170 7640 13175 7670
rect 13205 7640 13210 7670
rect 13170 7635 13210 7640
rect 13280 7670 13320 7675
rect 13280 7640 13285 7670
rect 13315 7640 13320 7670
rect 13280 7635 13320 7640
rect 13390 7670 13430 7675
rect 13390 7640 13395 7670
rect 13425 7640 13430 7670
rect 13390 7635 13430 7640
rect 13500 7670 13540 7675
rect 13500 7640 13505 7670
rect 13535 7640 13540 7670
rect 13500 7635 13540 7640
rect 13610 7670 13650 7675
rect 13610 7640 13615 7670
rect 13645 7640 13650 7670
rect 13610 7635 13650 7640
rect 13720 7670 13760 7675
rect 13720 7640 13725 7670
rect 13755 7640 13760 7670
rect 13720 7635 13760 7640
rect 13830 7670 13870 7675
rect 13830 7640 13835 7670
rect 13865 7640 13870 7670
rect 13830 7635 13870 7640
rect 13940 7670 13980 7675
rect 13940 7640 13945 7670
rect 13975 7640 13980 7670
rect 13940 7635 13980 7640
rect 14050 7670 14090 7675
rect 14050 7640 14055 7670
rect 14085 7640 14090 7670
rect 14050 7635 14090 7640
rect 17235 7670 17275 7675
rect 17235 7640 17240 7670
rect 17270 7640 17275 7670
rect 17235 7635 17275 7640
rect 17345 7670 17385 7675
rect 17345 7640 17350 7670
rect 17380 7640 17385 7670
rect 17345 7635 17385 7640
rect 17455 7670 17495 7675
rect 17455 7640 17460 7670
rect 17490 7640 17495 7670
rect 17455 7635 17495 7640
rect 17565 7670 17605 7675
rect 17565 7640 17570 7670
rect 17600 7640 17605 7670
rect 17565 7635 17605 7640
rect 17675 7670 17715 7675
rect 17675 7640 17680 7670
rect 17710 7640 17715 7670
rect 17675 7635 17715 7640
rect 17785 7670 17825 7675
rect 17785 7640 17790 7670
rect 17820 7640 17825 7670
rect 17785 7635 17825 7640
rect 17895 7670 17935 7675
rect 17895 7640 17900 7670
rect 17930 7640 17935 7670
rect 17895 7635 17935 7640
rect 18005 7670 18045 7675
rect 18005 7640 18010 7670
rect 18040 7640 18045 7670
rect 18005 7635 18045 7640
rect 18115 7670 18155 7675
rect 18115 7640 18120 7670
rect 18150 7640 18155 7670
rect 18115 7635 18155 7640
rect 18225 7670 18265 7675
rect 18225 7640 18230 7670
rect 18260 7640 18265 7670
rect 18225 7635 18265 7640
rect 18335 7670 18375 7675
rect 18335 7640 18340 7670
rect 18370 7640 18375 7670
rect 18335 7635 18375 7640
rect 13005 7500 13045 7505
rect 13005 7470 13010 7500
rect 13040 7470 13045 7500
rect 13005 7465 13045 7470
rect 13115 7500 13155 7505
rect 13115 7470 13120 7500
rect 13150 7470 13155 7500
rect 13115 7465 13155 7470
rect 13225 7500 13265 7505
rect 13225 7470 13230 7500
rect 13260 7470 13265 7500
rect 13225 7465 13265 7470
rect 13335 7500 13375 7505
rect 13335 7470 13340 7500
rect 13370 7470 13375 7500
rect 13335 7465 13375 7470
rect 13445 7500 13485 7505
rect 13445 7470 13450 7500
rect 13480 7470 13485 7500
rect 13445 7465 13485 7470
rect 13555 7500 13595 7505
rect 13555 7470 13560 7500
rect 13590 7470 13595 7500
rect 13555 7465 13595 7470
rect 13665 7500 13705 7505
rect 13665 7470 13670 7500
rect 13700 7470 13705 7500
rect 13665 7465 13705 7470
rect 13775 7500 13815 7505
rect 13775 7470 13780 7500
rect 13810 7470 13815 7500
rect 13775 7465 13815 7470
rect 13885 7500 13925 7505
rect 13885 7470 13890 7500
rect 13920 7470 13925 7500
rect 13885 7465 13925 7470
rect 13995 7500 14035 7505
rect 13995 7470 14000 7500
rect 14030 7470 14035 7500
rect 13995 7465 14035 7470
rect 17290 7500 17330 7505
rect 17290 7470 17295 7500
rect 17325 7470 17330 7500
rect 17290 7465 17330 7470
rect 17400 7500 17440 7505
rect 17400 7470 17405 7500
rect 17435 7470 17440 7500
rect 17400 7465 17440 7470
rect 17510 7500 17550 7505
rect 17510 7470 17515 7500
rect 17545 7470 17550 7500
rect 17510 7465 17550 7470
rect 17620 7500 17660 7505
rect 17620 7470 17625 7500
rect 17655 7470 17660 7500
rect 17620 7465 17660 7470
rect 17730 7500 17770 7505
rect 17730 7470 17735 7500
rect 17765 7470 17770 7500
rect 17730 7465 17770 7470
rect 17840 7500 17880 7505
rect 17840 7470 17845 7500
rect 17875 7470 17880 7500
rect 17840 7465 17880 7470
rect 17950 7500 17990 7505
rect 17950 7470 17955 7500
rect 17985 7470 17990 7500
rect 17950 7465 17990 7470
rect 18060 7500 18100 7505
rect 18060 7470 18065 7500
rect 18095 7470 18100 7500
rect 18060 7465 18100 7470
rect 18170 7500 18210 7505
rect 18170 7470 18175 7500
rect 18205 7470 18210 7500
rect 18170 7465 18210 7470
rect 18280 7500 18320 7505
rect 18280 7470 18285 7500
rect 18315 7470 18320 7500
rect 18490 7480 18510 8175
rect 18780 8150 18820 8160
rect 18780 8130 18790 8150
rect 18810 8130 18820 8150
rect 18780 8120 18820 8130
rect 18900 8150 18940 8160
rect 18900 8130 18910 8150
rect 18930 8130 18940 8150
rect 18900 8120 18940 8130
rect 19020 8150 19060 8160
rect 19020 8130 19030 8150
rect 19050 8130 19060 8150
rect 19020 8120 19060 8130
rect 19140 8150 19180 8160
rect 19140 8130 19150 8150
rect 19170 8130 19180 8150
rect 19140 8120 19180 8130
rect 19260 8150 19300 8160
rect 19260 8130 19270 8150
rect 19290 8130 19300 8150
rect 19260 8120 19300 8130
rect 19323 8155 19357 8160
rect 19323 8125 19326 8155
rect 19354 8125 19357 8155
rect 19323 8120 19357 8125
rect 19380 8150 19420 8160
rect 19380 8130 19390 8150
rect 19410 8130 19420 8150
rect 19380 8120 19420 8130
rect 19500 8150 19540 8160
rect 19500 8130 19510 8150
rect 19530 8130 19540 8150
rect 19500 8120 19540 8130
rect 19620 8150 19660 8160
rect 19620 8130 19630 8150
rect 19650 8130 19660 8150
rect 19620 8120 19660 8130
rect 19740 8150 19780 8160
rect 19740 8130 19750 8150
rect 19770 8130 19780 8150
rect 19740 8120 19780 8130
rect 19860 8150 19900 8160
rect 19860 8130 19870 8150
rect 19890 8130 19900 8150
rect 19860 8120 19900 8130
rect 19980 8150 20020 8160
rect 19980 8130 19990 8150
rect 20010 8130 20020 8150
rect 19980 8120 20020 8130
rect 18790 8105 18810 8120
rect 18780 8100 18820 8105
rect 18780 8070 18785 8100
rect 18815 8070 18820 8100
rect 18780 8065 18820 8070
rect 18910 8060 18930 8120
rect 19030 8105 19050 8120
rect 19020 8100 19060 8105
rect 19020 8070 19025 8100
rect 19055 8070 19060 8100
rect 19020 8065 19060 8070
rect 19150 8060 19170 8120
rect 19270 8105 19290 8120
rect 19260 8100 19300 8105
rect 19260 8070 19265 8100
rect 19295 8070 19300 8100
rect 19260 8065 19300 8070
rect 19390 8060 19410 8120
rect 19510 8105 19530 8120
rect 19500 8100 19540 8105
rect 19500 8070 19505 8100
rect 19535 8070 19540 8100
rect 19500 8065 19540 8070
rect 19630 8060 19650 8120
rect 19750 8105 19770 8120
rect 19740 8100 19780 8105
rect 19740 8070 19745 8100
rect 19775 8070 19780 8100
rect 19740 8065 19780 8070
rect 19870 8060 19890 8120
rect 19990 8105 20010 8120
rect 19980 8100 20020 8105
rect 19980 8070 19985 8100
rect 20015 8070 20020 8100
rect 19980 8065 20020 8070
rect 18900 8055 18940 8060
rect 18900 8025 18905 8055
rect 18935 8025 18940 8055
rect 18900 8020 18940 8025
rect 19140 8055 19180 8060
rect 19140 8025 19145 8055
rect 19175 8025 19180 8055
rect 19140 8020 19180 8025
rect 19380 8055 19420 8060
rect 19380 8025 19385 8055
rect 19415 8025 19420 8055
rect 19380 8020 19420 8025
rect 19620 8055 19660 8060
rect 19620 8025 19625 8055
rect 19655 8025 19660 8055
rect 19620 8020 19660 8025
rect 19860 8055 19900 8060
rect 19860 8025 19865 8055
rect 19895 8025 19900 8055
rect 19860 8020 19900 8025
rect 18910 8005 18930 8020
rect 18840 8000 18880 8005
rect 18840 7970 18845 8000
rect 18875 7970 18880 8000
rect 18840 7965 18880 7970
rect 18900 8000 18940 8005
rect 18900 7970 18905 8000
rect 18935 7970 18940 8000
rect 18900 7965 18940 7970
rect 19080 8000 19120 8005
rect 19080 7970 19085 8000
rect 19115 7970 19120 8000
rect 19080 7965 19120 7970
rect 19320 8000 19360 8005
rect 19320 7970 19325 8000
rect 19355 7970 19360 8000
rect 19320 7965 19360 7970
rect 19560 8000 19600 8005
rect 19560 7970 19565 8000
rect 19595 7970 19600 8000
rect 19560 7965 19600 7970
rect 19800 8000 19840 8005
rect 19800 7970 19805 8000
rect 19835 7970 19840 8000
rect 19800 7965 19840 7970
rect 18850 7950 18870 7965
rect 19090 7950 19110 7965
rect 19330 7950 19350 7965
rect 19570 7950 19590 7965
rect 19810 7950 19830 7965
rect 19990 7950 20010 8065
rect 18840 7940 18880 7950
rect 18840 7920 18850 7940
rect 18870 7920 18880 7940
rect 18840 7910 18880 7920
rect 18960 7945 19000 7950
rect 18960 7915 18965 7945
rect 18995 7915 19000 7945
rect 18960 7910 19000 7915
rect 19080 7940 19120 7950
rect 19080 7920 19090 7940
rect 19110 7920 19120 7940
rect 19080 7910 19120 7920
rect 19200 7945 19240 7950
rect 19200 7915 19205 7945
rect 19235 7915 19240 7945
rect 19200 7910 19240 7915
rect 19320 7940 19360 7950
rect 19320 7920 19330 7940
rect 19350 7920 19360 7940
rect 19320 7910 19360 7920
rect 19440 7945 19480 7950
rect 19440 7915 19445 7945
rect 19475 7915 19480 7945
rect 19440 7910 19480 7915
rect 19560 7940 19600 7950
rect 19560 7920 19570 7940
rect 19590 7920 19600 7940
rect 19560 7910 19600 7920
rect 19680 7945 19720 7950
rect 19680 7915 19685 7945
rect 19715 7915 19720 7945
rect 19680 7910 19720 7915
rect 19800 7940 19840 7950
rect 19800 7920 19810 7940
rect 19830 7920 19840 7940
rect 19800 7910 19840 7920
rect 19920 7945 19960 7950
rect 19920 7915 19925 7945
rect 19955 7915 19960 7945
rect 19920 7910 19960 7915
rect 19980 7945 20020 7950
rect 19980 7915 19985 7945
rect 20015 7915 20020 7945
rect 19980 7910 20020 7915
rect 20500 7920 20540 7925
rect 20500 7890 20505 7920
rect 20535 7890 20540 7920
rect 20500 7885 20540 7890
rect 20558 7915 20592 7925
rect 20558 7895 20566 7915
rect 20584 7895 20592 7915
rect 20558 7885 20592 7895
rect 20610 7920 20650 7925
rect 20610 7890 20615 7920
rect 20645 7890 20650 7920
rect 20610 7885 20650 7890
rect 20720 7920 20760 7925
rect 20720 7890 20725 7920
rect 20755 7890 20760 7920
rect 20720 7885 20760 7890
rect 20830 7920 20870 7925
rect 20830 7890 20835 7920
rect 20865 7890 20870 7920
rect 20830 7885 20870 7890
rect 20940 7920 20980 7925
rect 20940 7890 20945 7920
rect 20975 7890 20980 7920
rect 20940 7885 20980 7890
rect 21050 7920 21090 7925
rect 21050 7890 21055 7920
rect 21085 7890 21090 7920
rect 21050 7885 21090 7890
rect 21160 7920 21200 7925
rect 21160 7890 21165 7920
rect 21195 7890 21200 7920
rect 21160 7885 21200 7890
rect 21270 7920 21310 7925
rect 21270 7890 21275 7920
rect 21305 7890 21310 7920
rect 21270 7885 21310 7890
rect 21380 7920 21420 7925
rect 21380 7890 21385 7920
rect 21415 7890 21420 7920
rect 21380 7885 21420 7890
rect 21490 7920 21530 7925
rect 21490 7890 21495 7920
rect 21525 7890 21530 7920
rect 21490 7885 21530 7890
rect 20565 7836 20585 7885
rect 20555 7830 20595 7836
rect 20555 7800 20560 7830
rect 20590 7800 20595 7830
rect 20555 7780 20595 7800
rect 20555 7750 20560 7780
rect 20590 7750 20595 7780
rect 20190 7730 20230 7735
rect 20190 7700 20195 7730
rect 20225 7700 20230 7730
rect 20190 7695 20230 7700
rect 20555 7730 20595 7750
rect 20555 7700 20560 7730
rect 20590 7700 20595 7730
rect 20555 7695 20595 7700
rect 18280 7465 18320 7470
rect 18480 7475 18520 7480
rect 12978 7440 13012 7445
rect 12978 7410 12981 7440
rect 13009 7410 13012 7440
rect 12978 7405 13012 7410
rect 12985 7380 13005 7405
rect 14005 7380 14025 7465
rect 11880 7375 11920 7380
rect 11880 7345 11885 7375
rect 11915 7345 11920 7375
rect 11880 7340 11920 7345
rect 12120 7375 12160 7380
rect 12120 7345 12125 7375
rect 12155 7345 12160 7375
rect 12120 7340 12160 7345
rect 12360 7375 12400 7380
rect 12360 7345 12365 7375
rect 12395 7345 12400 7375
rect 12360 7340 12400 7345
rect 12690 7375 12730 7380
rect 12690 7345 12695 7375
rect 12725 7345 12730 7375
rect 12690 7340 12730 7345
rect 12975 7375 13015 7380
rect 12975 7345 12980 7375
rect 13010 7345 13015 7375
rect 12975 7340 13015 7345
rect 13145 7345 13150 7380
rect 13185 7345 13190 7380
rect 13979 7345 13985 7380
rect 14020 7345 14025 7380
rect 17300 7380 17320 7465
rect 18480 7445 18485 7475
rect 18515 7445 18520 7475
rect 18313 7440 18347 7445
rect 18480 7440 18520 7445
rect 18780 7470 18820 7480
rect 18780 7450 18790 7470
rect 18810 7450 18820 7470
rect 18780 7440 18820 7450
rect 18900 7470 18940 7480
rect 18900 7450 18910 7470
rect 18930 7450 18940 7470
rect 18900 7440 18940 7450
rect 19020 7470 19060 7480
rect 19020 7450 19030 7470
rect 19050 7450 19060 7470
rect 19020 7440 19060 7450
rect 19140 7470 19180 7480
rect 19140 7450 19150 7470
rect 19170 7450 19180 7470
rect 19140 7440 19180 7450
rect 19260 7470 19300 7480
rect 19260 7450 19270 7470
rect 19290 7450 19300 7470
rect 19260 7440 19300 7450
rect 19323 7475 19357 7480
rect 19323 7445 19326 7475
rect 19354 7445 19357 7475
rect 19323 7440 19357 7445
rect 19380 7470 19420 7480
rect 19380 7450 19390 7470
rect 19410 7450 19420 7470
rect 19380 7440 19420 7450
rect 19500 7470 19540 7480
rect 19500 7450 19510 7470
rect 19530 7450 19540 7470
rect 19500 7440 19540 7450
rect 19620 7470 19660 7480
rect 19620 7450 19630 7470
rect 19650 7450 19660 7470
rect 19620 7440 19660 7450
rect 19740 7470 19780 7480
rect 19740 7450 19750 7470
rect 19770 7450 19780 7470
rect 19740 7440 19780 7450
rect 19860 7470 19900 7480
rect 19860 7450 19870 7470
rect 19890 7450 19900 7470
rect 19860 7440 19900 7450
rect 19980 7470 20020 7480
rect 19980 7450 19990 7470
rect 20010 7450 20020 7470
rect 19980 7440 20020 7450
rect 18313 7410 18316 7440
rect 18344 7410 18347 7440
rect 18790 7425 18810 7440
rect 18313 7405 18347 7410
rect 18780 7420 18820 7425
rect 17300 7345 17305 7380
rect 17340 7345 17345 7380
rect 18135 7345 18140 7380
rect 18175 7345 18180 7380
rect 12120 7285 12140 7340
rect 12815 7325 12855 7330
rect 12815 7295 12820 7325
rect 12850 7295 12855 7325
rect 12815 7290 12855 7295
rect 11880 7280 11920 7285
rect 11880 7250 11885 7280
rect 11915 7250 11920 7280
rect 11880 7245 11920 7250
rect 12100 7280 12140 7285
rect 12100 7250 12105 7280
rect 12135 7250 12140 7280
rect 12100 7245 12140 7250
rect 12320 7280 12360 7285
rect 12320 7250 12325 7280
rect 12355 7250 12360 7280
rect 12320 7245 12360 7250
rect 11770 7235 11810 7240
rect 11770 7205 11775 7235
rect 11805 7205 11810 7235
rect 11770 7200 11810 7205
rect 11780 7185 11800 7200
rect 11890 7185 11910 7245
rect 11990 7235 12030 7240
rect 11990 7205 11995 7235
rect 12025 7205 12030 7235
rect 11990 7200 12030 7205
rect 12000 7185 12020 7200
rect 12110 7185 12130 7245
rect 12210 7235 12250 7240
rect 12210 7205 12215 7235
rect 12245 7205 12250 7235
rect 12210 7200 12250 7205
rect 12220 7185 12240 7200
rect 12330 7185 12350 7245
rect 12430 7235 12470 7240
rect 12430 7205 12435 7235
rect 12465 7205 12470 7235
rect 12430 7200 12470 7205
rect 12440 7185 12460 7200
rect 11330 7175 11370 7185
rect 11330 7155 11340 7175
rect 11360 7155 11370 7175
rect 11330 7145 11370 7155
rect 11440 7175 11480 7185
rect 11440 7155 11450 7175
rect 11470 7155 11480 7175
rect 11440 7145 11480 7155
rect 11550 7175 11590 7185
rect 11550 7155 11560 7175
rect 11580 7155 11590 7175
rect 11550 7145 11590 7155
rect 11660 7175 11700 7185
rect 11660 7155 11670 7175
rect 11690 7155 11700 7175
rect 11660 7145 11700 7155
rect 11770 7175 11810 7185
rect 11770 7155 11780 7175
rect 11800 7155 11810 7175
rect 11770 7145 11810 7155
rect 11880 7175 11920 7185
rect 11880 7155 11890 7175
rect 11910 7155 11920 7175
rect 11880 7145 11920 7155
rect 11990 7175 12030 7185
rect 11990 7155 12000 7175
rect 12020 7155 12030 7175
rect 11990 7145 12030 7155
rect 12100 7175 12140 7185
rect 12100 7155 12110 7175
rect 12130 7155 12140 7175
rect 12100 7145 12140 7155
rect 12210 7175 12250 7185
rect 12210 7155 12220 7175
rect 12240 7155 12250 7175
rect 12210 7145 12250 7155
rect 12320 7175 12360 7185
rect 12320 7155 12330 7175
rect 12350 7155 12360 7175
rect 12320 7145 12360 7155
rect 12430 7175 12470 7185
rect 12430 7155 12440 7175
rect 12460 7155 12470 7175
rect 12430 7145 12470 7155
rect 9735 7000 9775 7005
rect 9735 6970 9740 7000
rect 9770 6970 9775 7000
rect 9735 6965 9775 6970
rect 9845 7000 9885 7005
rect 9845 6970 9850 7000
rect 9880 6970 9885 7000
rect 9845 6965 9885 6970
rect 9955 7000 9995 7005
rect 9955 6970 9960 7000
rect 9990 6970 9995 7000
rect 9955 6965 9995 6970
rect 10065 7000 10105 7005
rect 10065 6970 10070 7000
rect 10100 6970 10105 7000
rect 10065 6965 10105 6970
rect 10175 7000 10215 7005
rect 10175 6970 10180 7000
rect 10210 6970 10215 7000
rect 10175 6965 10215 6970
rect 10285 7000 10325 7005
rect 10285 6970 10290 7000
rect 10320 6970 10325 7000
rect 10285 6965 10325 6970
rect 10395 7000 10435 7005
rect 10395 6970 10400 7000
rect 10430 6970 10435 7000
rect 10395 6965 10435 6970
rect 10505 7000 10545 7005
rect 10505 6970 10510 7000
rect 10540 6970 10545 7000
rect 10505 6965 10545 6970
rect 10615 7000 10655 7005
rect 10615 6970 10620 7000
rect 10650 6970 10655 7000
rect 10615 6965 10655 6970
rect 10725 7000 10765 7005
rect 10725 6970 10730 7000
rect 10760 6970 10765 7000
rect 10725 6965 10765 6970
rect 10835 7000 10875 7005
rect 10835 6970 10840 7000
rect 10870 6970 10875 7000
rect 10835 6965 10875 6970
rect 11385 6960 11425 6965
rect 11385 6930 11390 6960
rect 11420 6930 11425 6960
rect 11385 6925 11425 6930
rect 11495 6955 11535 6965
rect 11495 6935 11505 6955
rect 11525 6935 11535 6955
rect 11495 6925 11535 6935
rect 11605 6960 11645 6965
rect 11605 6930 11610 6960
rect 11640 6930 11645 6960
rect 11605 6925 11645 6930
rect 11715 6955 11755 6965
rect 11715 6935 11725 6955
rect 11745 6935 11755 6955
rect 11715 6925 11755 6935
rect 11825 6960 11865 6965
rect 11825 6930 11830 6960
rect 11860 6930 11865 6960
rect 11825 6925 11865 6930
rect 11935 6955 11975 6965
rect 11935 6935 11945 6955
rect 11965 6935 11975 6955
rect 11935 6925 11975 6935
rect 12045 6960 12085 6965
rect 12045 6930 12050 6960
rect 12080 6930 12085 6960
rect 12045 6925 12085 6930
rect 12155 6955 12195 6965
rect 12155 6935 12165 6955
rect 12185 6935 12195 6955
rect 12155 6925 12195 6935
rect 12245 6960 12305 6965
rect 12245 6930 12270 6960
rect 12300 6930 12305 6960
rect 12245 6925 12305 6930
rect 12375 6955 12415 6965
rect 12375 6935 12385 6955
rect 12405 6935 12415 6955
rect 12375 6925 12415 6935
rect 11505 6910 11525 6925
rect 11725 6910 11745 6925
rect 11945 6910 11965 6925
rect 12165 6910 12185 6925
rect 11495 6905 11555 6910
rect 11495 6875 11500 6905
rect 11530 6875 11555 6905
rect 11495 6870 11555 6875
rect 11715 6905 11755 6910
rect 11715 6875 11720 6905
rect 11750 6875 11755 6905
rect 11715 6870 11755 6875
rect 11935 6905 11975 6910
rect 11935 6875 11940 6905
rect 11970 6875 11975 6905
rect 11935 6870 11975 6875
rect 12155 6905 12195 6910
rect 12155 6875 12160 6905
rect 12190 6875 12195 6905
rect 12155 6870 12195 6875
rect 11190 6850 11230 6855
rect 11190 6820 11195 6850
rect 11225 6820 11230 6850
rect 11190 6815 11230 6820
rect 11410 6850 11450 6855
rect 11410 6820 11415 6850
rect 11445 6820 11450 6850
rect 11410 6815 11450 6820
rect 11200 6780 11220 6815
rect 11420 6780 11440 6815
rect 11190 6770 11230 6780
rect 11085 6760 11125 6765
rect 11085 6730 11090 6760
rect 11120 6730 11125 6760
rect 11190 6750 11200 6770
rect 11220 6750 11230 6770
rect 11410 6770 11450 6780
rect 11190 6740 11230 6750
rect 11305 6760 11345 6765
rect 11085 6725 11125 6730
rect 11305 6730 11310 6760
rect 11340 6730 11345 6760
rect 11410 6750 11420 6770
rect 11440 6750 11450 6770
rect 11535 6765 11555 6870
rect 12245 6855 12265 6925
rect 12385 6910 12405 6925
rect 12375 6905 12415 6910
rect 12375 6875 12380 6905
rect 12410 6875 12415 6905
rect 12375 6870 12415 6875
rect 11640 6850 11680 6855
rect 11640 6820 11645 6850
rect 11675 6820 11680 6850
rect 11640 6815 11680 6820
rect 12230 6850 12270 6855
rect 12230 6820 12235 6850
rect 12265 6820 12270 6850
rect 12230 6815 12270 6820
rect 12450 6850 12490 6855
rect 12450 6820 12455 6850
rect 12485 6820 12490 6850
rect 12450 6815 12490 6820
rect 12680 6850 12720 6855
rect 12680 6820 12685 6850
rect 12715 6820 12720 6850
rect 12680 6815 12720 6820
rect 11650 6780 11670 6815
rect 11820 6805 11860 6810
rect 11640 6770 11680 6780
rect 11820 6775 11825 6805
rect 11855 6775 11860 6805
rect 11820 6770 11860 6775
rect 11940 6805 11980 6810
rect 11940 6775 11945 6805
rect 11975 6775 11980 6805
rect 12240 6780 12260 6815
rect 12460 6780 12480 6815
rect 12690 6780 12710 6815
rect 11940 6770 11980 6775
rect 12230 6770 12270 6780
rect 11410 6740 11450 6750
rect 11525 6760 11565 6765
rect 11305 6725 11345 6730
rect 11525 6730 11530 6760
rect 11560 6730 11565 6760
rect 11640 6750 11650 6770
rect 11670 6750 11680 6770
rect 11640 6740 11680 6750
rect 11525 6725 11565 6730
rect 11830 6720 11850 6770
rect 11950 6720 11970 6770
rect 12125 6760 12165 6765
rect 12125 6730 12130 6760
rect 12160 6730 12165 6760
rect 12230 6750 12240 6770
rect 12260 6750 12270 6770
rect 12450 6770 12490 6780
rect 12230 6740 12270 6750
rect 12345 6760 12385 6765
rect 12125 6725 12165 6730
rect 12345 6730 12350 6760
rect 12380 6730 12385 6760
rect 12450 6750 12460 6770
rect 12480 6750 12490 6770
rect 12680 6770 12720 6780
rect 12450 6740 12490 6750
rect 12565 6760 12605 6765
rect 12345 6725 12385 6730
rect 12565 6730 12570 6760
rect 12600 6730 12605 6760
rect 12680 6750 12690 6770
rect 12710 6750 12720 6770
rect 12680 6740 12720 6750
rect 12565 6725 12605 6730
rect 11237 6715 11269 6720
rect 11237 6685 11240 6715
rect 11266 6685 11269 6715
rect 11237 6680 11269 6685
rect 11457 6715 11489 6720
rect 11457 6685 11460 6715
rect 11486 6685 11489 6715
rect 11457 6680 11489 6685
rect 11601 6715 11633 6720
rect 11601 6685 11604 6715
rect 11630 6685 11633 6715
rect 11601 6680 11633 6685
rect 11820 6710 11850 6720
rect 11820 6690 11825 6710
rect 11845 6690 11850 6710
rect 11820 6680 11850 6690
rect 11867 6715 11899 6720
rect 11867 6685 11870 6715
rect 11896 6685 11899 6715
rect 11867 6680 11899 6685
rect 11950 6710 11980 6720
rect 11950 6690 11955 6710
rect 11975 6690 11980 6710
rect 11950 6680 11980 6690
rect 12277 6715 12309 6720
rect 12277 6685 12280 6715
rect 12306 6685 12309 6715
rect 12277 6680 12309 6685
rect 12497 6715 12529 6720
rect 12497 6685 12500 6715
rect 12526 6685 12529 6715
rect 12497 6680 12529 6685
rect 12641 6715 12673 6720
rect 12641 6685 12644 6715
rect 12670 6685 12673 6715
rect 12641 6680 12673 6685
rect 12825 6575 12845 7290
rect 12985 7285 13005 7340
rect 13145 7320 13190 7345
rect 18135 7320 18180 7345
rect 13145 7285 13150 7320
rect 13185 7285 13190 7320
rect 13980 7285 13985 7320
rect 14020 7285 14025 7320
rect 12978 7280 13012 7285
rect 12978 7250 12981 7280
rect 13009 7250 13012 7280
rect 12978 7245 13012 7250
rect 14005 7225 14025 7285
rect 17300 7285 17305 7320
rect 17340 7285 17345 7320
rect 18135 7285 18140 7320
rect 18175 7285 18180 7320
rect 18320 7285 18340 7405
rect 18780 7390 18785 7420
rect 18815 7390 18820 7420
rect 18780 7385 18820 7390
rect 18910 7380 18930 7440
rect 19030 7425 19050 7440
rect 19020 7420 19060 7425
rect 19020 7390 19025 7420
rect 19055 7390 19060 7420
rect 19020 7385 19060 7390
rect 19150 7380 19170 7440
rect 19270 7425 19290 7440
rect 19260 7420 19300 7425
rect 19260 7390 19265 7420
rect 19295 7390 19300 7420
rect 19260 7385 19300 7390
rect 18900 7375 18940 7380
rect 18900 7345 18905 7375
rect 18935 7345 18940 7375
rect 18900 7340 18940 7345
rect 19140 7375 19180 7380
rect 19140 7345 19145 7375
rect 19175 7345 19180 7375
rect 19140 7340 19180 7345
rect 17300 7225 17320 7285
rect 18313 7280 18347 7285
rect 18313 7250 18316 7280
rect 18344 7250 18347 7280
rect 18313 7245 18347 7250
rect 18940 7280 18980 7285
rect 18940 7250 18945 7280
rect 18975 7250 18980 7280
rect 18940 7245 18980 7250
rect 19160 7280 19200 7285
rect 19160 7250 19165 7280
rect 19195 7250 19200 7280
rect 19160 7245 19200 7250
rect 18830 7235 18870 7240
rect 13005 7220 13045 7225
rect 13005 7190 13010 7220
rect 13040 7190 13045 7220
rect 13005 7185 13045 7190
rect 13115 7220 13155 7225
rect 13115 7190 13120 7220
rect 13150 7190 13155 7220
rect 13115 7185 13155 7190
rect 13225 7220 13265 7225
rect 13225 7190 13230 7220
rect 13260 7190 13265 7220
rect 13225 7185 13265 7190
rect 13335 7220 13375 7225
rect 13335 7190 13340 7220
rect 13370 7190 13375 7220
rect 13335 7185 13375 7190
rect 13445 7220 13485 7225
rect 13445 7190 13450 7220
rect 13480 7190 13485 7220
rect 13445 7185 13485 7190
rect 13555 7220 13595 7225
rect 13555 7190 13560 7220
rect 13590 7190 13595 7220
rect 13555 7185 13595 7190
rect 13665 7220 13705 7225
rect 13665 7190 13670 7220
rect 13700 7190 13705 7220
rect 13665 7185 13705 7190
rect 13775 7220 13815 7225
rect 13775 7190 13780 7220
rect 13810 7190 13815 7220
rect 13775 7185 13815 7190
rect 13885 7220 13925 7225
rect 13885 7190 13890 7220
rect 13920 7190 13925 7220
rect 13885 7185 13925 7190
rect 13995 7220 14035 7225
rect 13995 7190 14000 7220
rect 14030 7190 14035 7220
rect 13995 7185 14035 7190
rect 17290 7220 17330 7225
rect 17290 7190 17295 7220
rect 17325 7190 17330 7220
rect 17290 7185 17330 7190
rect 17400 7220 17440 7225
rect 17400 7190 17405 7220
rect 17435 7190 17440 7220
rect 17400 7185 17440 7190
rect 17510 7220 17550 7225
rect 17510 7190 17515 7220
rect 17545 7190 17550 7220
rect 17510 7185 17550 7190
rect 17620 7220 17660 7225
rect 17620 7190 17625 7220
rect 17655 7190 17660 7220
rect 17620 7185 17660 7190
rect 17730 7220 17770 7225
rect 17730 7190 17735 7220
rect 17765 7190 17770 7220
rect 17730 7185 17770 7190
rect 17840 7220 17880 7225
rect 17840 7190 17845 7220
rect 17875 7190 17880 7220
rect 17840 7185 17880 7190
rect 17950 7220 17990 7225
rect 17950 7190 17955 7220
rect 17985 7190 17990 7220
rect 17950 7185 17990 7190
rect 18060 7220 18100 7225
rect 18060 7190 18065 7220
rect 18095 7190 18100 7220
rect 18060 7185 18100 7190
rect 18170 7220 18210 7225
rect 18170 7190 18175 7220
rect 18205 7190 18210 7220
rect 18170 7185 18210 7190
rect 18280 7220 18320 7225
rect 18280 7190 18285 7220
rect 18315 7190 18320 7220
rect 18830 7205 18835 7235
rect 18865 7205 18870 7235
rect 18830 7200 18870 7205
rect 18280 7185 18320 7190
rect 18840 7185 18860 7200
rect 18950 7185 18970 7245
rect 19050 7235 19090 7240
rect 19050 7205 19055 7235
rect 19085 7205 19090 7235
rect 19050 7200 19090 7205
rect 19060 7185 19080 7200
rect 19170 7185 19190 7245
rect 19270 7240 19290 7385
rect 19390 7380 19410 7440
rect 19510 7425 19530 7440
rect 19500 7420 19540 7425
rect 19500 7390 19505 7420
rect 19535 7390 19540 7420
rect 19500 7385 19540 7390
rect 19630 7380 19650 7440
rect 19750 7425 19770 7440
rect 19740 7420 19780 7425
rect 19740 7390 19745 7420
rect 19775 7390 19780 7420
rect 19740 7385 19780 7390
rect 19870 7380 19890 7440
rect 19990 7425 20010 7440
rect 19980 7420 20020 7425
rect 19980 7390 19985 7420
rect 20015 7390 20020 7420
rect 19980 7385 20020 7390
rect 20200 7380 20220 7695
rect 20445 7670 20485 7675
rect 20445 7640 20450 7670
rect 20480 7640 20485 7670
rect 20445 7635 20485 7640
rect 20555 7670 20595 7675
rect 20555 7640 20560 7670
rect 20590 7640 20595 7670
rect 20555 7635 20595 7640
rect 20665 7670 20705 7675
rect 20665 7640 20670 7670
rect 20700 7640 20705 7670
rect 20665 7635 20705 7640
rect 20775 7670 20815 7675
rect 20775 7640 20780 7670
rect 20810 7640 20815 7670
rect 20775 7635 20815 7640
rect 20885 7670 20925 7675
rect 20885 7640 20890 7670
rect 20920 7640 20925 7670
rect 20885 7635 20925 7640
rect 20995 7670 21035 7675
rect 20995 7640 21000 7670
rect 21030 7640 21035 7670
rect 20995 7635 21035 7640
rect 21105 7670 21145 7675
rect 21105 7640 21110 7670
rect 21140 7640 21145 7670
rect 21105 7635 21145 7640
rect 21215 7670 21255 7675
rect 21215 7640 21220 7670
rect 21250 7640 21255 7670
rect 21215 7635 21255 7640
rect 21325 7670 21365 7675
rect 21325 7640 21330 7670
rect 21360 7640 21365 7670
rect 21325 7635 21365 7640
rect 21435 7670 21475 7675
rect 21435 7640 21440 7670
rect 21470 7640 21475 7670
rect 21435 7635 21475 7640
rect 21545 7670 21585 7675
rect 21545 7640 21550 7670
rect 21580 7640 21585 7670
rect 21545 7635 21585 7640
rect 20500 7500 20540 7505
rect 20500 7470 20505 7500
rect 20535 7470 20540 7500
rect 20500 7465 20540 7470
rect 20610 7500 20650 7505
rect 20610 7470 20615 7500
rect 20645 7470 20650 7500
rect 20610 7465 20650 7470
rect 20720 7500 20760 7505
rect 20720 7470 20725 7500
rect 20755 7470 20760 7500
rect 20720 7465 20760 7470
rect 20830 7500 20870 7505
rect 20830 7470 20835 7500
rect 20865 7470 20870 7500
rect 20830 7465 20870 7470
rect 20940 7500 20980 7505
rect 20940 7470 20945 7500
rect 20975 7470 20980 7500
rect 20940 7465 20980 7470
rect 21050 7500 21090 7505
rect 21050 7470 21055 7500
rect 21085 7470 21090 7500
rect 21050 7465 21090 7470
rect 21160 7500 21200 7505
rect 21160 7470 21165 7500
rect 21195 7470 21200 7500
rect 21160 7465 21200 7470
rect 21270 7500 21310 7505
rect 21270 7470 21275 7500
rect 21305 7470 21310 7500
rect 21270 7465 21310 7470
rect 21380 7500 21420 7505
rect 21380 7470 21385 7500
rect 21415 7470 21420 7500
rect 21380 7465 21420 7470
rect 21490 7500 21530 7505
rect 21490 7470 21495 7500
rect 21525 7470 21530 7500
rect 21490 7465 21530 7470
rect 20473 7440 20507 7445
rect 20473 7410 20476 7440
rect 20504 7410 20507 7440
rect 20473 7405 20507 7410
rect 20480 7380 20500 7405
rect 21500 7380 21520 7465
rect 19380 7375 19420 7380
rect 19380 7345 19385 7375
rect 19415 7345 19420 7375
rect 19380 7340 19420 7345
rect 19620 7375 19660 7380
rect 19620 7345 19625 7375
rect 19655 7345 19660 7375
rect 19620 7340 19660 7345
rect 19860 7375 19900 7380
rect 19860 7345 19865 7375
rect 19895 7345 19900 7375
rect 19860 7340 19900 7345
rect 20190 7375 20230 7380
rect 20190 7345 20195 7375
rect 20225 7345 20230 7375
rect 20190 7340 20230 7345
rect 20470 7375 20510 7380
rect 20470 7345 20475 7375
rect 20505 7345 20510 7375
rect 20470 7340 20510 7345
rect 20640 7345 20645 7380
rect 20680 7345 20685 7380
rect 21474 7345 21480 7380
rect 21515 7345 21520 7380
rect 19620 7285 19640 7340
rect 20315 7325 20355 7330
rect 20315 7295 20320 7325
rect 20350 7295 20355 7325
rect 20315 7290 20355 7295
rect 19380 7280 19420 7285
rect 19380 7250 19385 7280
rect 19415 7250 19420 7280
rect 19380 7245 19420 7250
rect 19600 7280 19640 7285
rect 19600 7250 19605 7280
rect 19635 7250 19640 7280
rect 19600 7245 19640 7250
rect 19820 7280 19860 7285
rect 19820 7250 19825 7280
rect 19855 7250 19860 7280
rect 19820 7245 19860 7250
rect 19270 7235 19310 7240
rect 19270 7205 19275 7235
rect 19305 7205 19310 7235
rect 19270 7200 19310 7205
rect 19280 7185 19300 7200
rect 19390 7185 19410 7245
rect 19490 7235 19530 7240
rect 19490 7205 19495 7235
rect 19525 7205 19530 7235
rect 19490 7200 19530 7205
rect 19500 7185 19520 7200
rect 19610 7185 19630 7245
rect 19710 7235 19750 7240
rect 19710 7205 19715 7235
rect 19745 7205 19750 7235
rect 19710 7200 19750 7205
rect 19720 7185 19740 7200
rect 19830 7185 19850 7245
rect 19930 7235 19970 7240
rect 19930 7205 19935 7235
rect 19965 7205 19970 7235
rect 19930 7200 19970 7205
rect 19940 7185 19960 7200
rect 18830 7175 18870 7185
rect 18830 7155 18840 7175
rect 18860 7155 18870 7175
rect 18830 7145 18870 7155
rect 18940 7175 18980 7185
rect 18940 7155 18950 7175
rect 18970 7155 18980 7175
rect 18940 7145 18980 7155
rect 19050 7175 19090 7185
rect 19050 7155 19060 7175
rect 19080 7155 19090 7175
rect 19050 7145 19090 7155
rect 19160 7175 19200 7185
rect 19160 7155 19170 7175
rect 19190 7155 19200 7175
rect 19160 7145 19200 7155
rect 19270 7175 19310 7185
rect 19270 7155 19280 7175
rect 19300 7155 19310 7175
rect 19270 7145 19310 7155
rect 19380 7175 19420 7185
rect 19380 7155 19390 7175
rect 19410 7155 19420 7175
rect 19380 7145 19420 7155
rect 19490 7175 19530 7185
rect 19490 7155 19500 7175
rect 19520 7155 19530 7175
rect 19490 7145 19530 7155
rect 19600 7175 19640 7185
rect 19600 7155 19610 7175
rect 19630 7155 19640 7175
rect 19600 7145 19640 7155
rect 19710 7175 19750 7185
rect 19710 7155 19720 7175
rect 19740 7155 19750 7175
rect 19710 7145 19750 7155
rect 19820 7175 19860 7185
rect 19820 7155 19830 7175
rect 19850 7155 19860 7175
rect 19820 7145 19860 7155
rect 19930 7175 19970 7185
rect 19930 7155 19940 7175
rect 19960 7155 19970 7175
rect 19930 7145 19970 7155
rect 12950 7000 12990 7005
rect 12950 6970 12955 7000
rect 12985 6970 12990 7000
rect 12950 6965 12990 6970
rect 13060 7000 13100 7005
rect 13060 6970 13065 7000
rect 13095 6970 13100 7000
rect 13060 6965 13100 6970
rect 13170 7000 13210 7005
rect 13170 6970 13175 7000
rect 13205 6970 13210 7000
rect 13170 6965 13210 6970
rect 13280 7000 13320 7005
rect 13280 6970 13285 7000
rect 13315 6970 13320 7000
rect 13280 6965 13320 6970
rect 13390 7000 13430 7005
rect 13390 6970 13395 7000
rect 13425 6970 13430 7000
rect 13390 6965 13430 6970
rect 13500 7000 13540 7005
rect 13500 6970 13505 7000
rect 13535 6970 13540 7000
rect 13500 6965 13540 6970
rect 13610 7000 13650 7005
rect 13610 6970 13615 7000
rect 13645 6970 13650 7000
rect 13610 6965 13650 6970
rect 13720 7000 13760 7005
rect 13720 6970 13725 7000
rect 13755 6970 13760 7000
rect 13720 6965 13760 6970
rect 13830 7000 13870 7005
rect 13830 6970 13835 7000
rect 13865 6970 13870 7000
rect 13830 6965 13870 6970
rect 13940 7000 13980 7005
rect 13940 6970 13945 7000
rect 13975 6970 13980 7000
rect 13940 6965 13980 6970
rect 14050 7000 14090 7005
rect 14050 6970 14055 7000
rect 14085 6970 14090 7000
rect 14050 6965 14090 6970
rect 17235 7000 17275 7005
rect 17235 6970 17240 7000
rect 17270 6970 17275 7000
rect 17235 6965 17275 6970
rect 17345 7000 17385 7005
rect 17345 6970 17350 7000
rect 17380 6970 17385 7000
rect 17345 6965 17385 6970
rect 17455 7000 17495 7005
rect 17455 6970 17460 7000
rect 17490 6970 17495 7000
rect 17455 6965 17495 6970
rect 17565 7000 17605 7005
rect 17565 6970 17570 7000
rect 17600 6970 17605 7000
rect 17565 6965 17605 6970
rect 17675 7000 17715 7005
rect 17675 6970 17680 7000
rect 17710 6970 17715 7000
rect 17675 6965 17715 6970
rect 17785 7000 17825 7005
rect 17785 6970 17790 7000
rect 17820 6970 17825 7000
rect 17785 6965 17825 6970
rect 17895 7000 17935 7005
rect 17895 6970 17900 7000
rect 17930 6970 17935 7000
rect 17895 6965 17935 6970
rect 18005 7000 18045 7005
rect 18005 6970 18010 7000
rect 18040 6970 18045 7000
rect 18005 6965 18045 6970
rect 18115 7000 18155 7005
rect 18115 6970 18120 7000
rect 18150 6970 18155 7000
rect 18115 6965 18155 6970
rect 18225 7000 18265 7005
rect 18225 6970 18230 7000
rect 18260 6970 18265 7000
rect 18225 6965 18265 6970
rect 18335 7000 18375 7005
rect 18335 6970 18340 7000
rect 18370 6970 18375 7000
rect 18335 6965 18375 6970
rect 18885 6960 18925 6965
rect 18885 6930 18890 6960
rect 18920 6930 18925 6960
rect 18885 6925 18925 6930
rect 18995 6955 19035 6965
rect 18995 6935 19005 6955
rect 19025 6935 19035 6955
rect 18995 6925 19035 6935
rect 19105 6960 19145 6965
rect 19105 6930 19110 6960
rect 19140 6930 19145 6960
rect 19105 6925 19145 6930
rect 19215 6955 19255 6965
rect 19215 6935 19225 6955
rect 19245 6935 19255 6955
rect 19215 6925 19255 6935
rect 19325 6960 19365 6965
rect 19325 6930 19330 6960
rect 19360 6930 19365 6960
rect 19325 6925 19365 6930
rect 19435 6955 19475 6965
rect 19435 6935 19445 6955
rect 19465 6935 19475 6955
rect 19435 6925 19475 6935
rect 19545 6960 19585 6965
rect 19545 6930 19550 6960
rect 19580 6930 19585 6960
rect 19545 6925 19585 6930
rect 19655 6955 19695 6965
rect 19655 6935 19665 6955
rect 19685 6935 19695 6955
rect 19655 6925 19695 6935
rect 19745 6960 19805 6965
rect 19745 6930 19770 6960
rect 19800 6930 19805 6960
rect 19745 6925 19805 6930
rect 19875 6955 19915 6965
rect 19875 6935 19885 6955
rect 19905 6935 19915 6955
rect 19875 6925 19915 6935
rect 19005 6910 19025 6925
rect 19225 6910 19245 6925
rect 19445 6910 19465 6925
rect 19665 6910 19685 6925
rect 18995 6905 19055 6910
rect 18995 6875 19000 6905
rect 19030 6875 19055 6905
rect 18995 6870 19055 6875
rect 19215 6905 19255 6910
rect 19215 6875 19220 6905
rect 19250 6875 19255 6905
rect 19215 6870 19255 6875
rect 19435 6905 19475 6910
rect 19435 6875 19440 6905
rect 19470 6875 19475 6905
rect 19435 6870 19475 6875
rect 19655 6905 19695 6910
rect 19655 6875 19660 6905
rect 19690 6875 19695 6905
rect 19655 6870 19695 6875
rect 18690 6850 18730 6855
rect 18690 6820 18695 6850
rect 18725 6820 18730 6850
rect 18690 6815 18730 6820
rect 18910 6850 18950 6855
rect 18910 6820 18915 6850
rect 18945 6820 18950 6850
rect 18910 6815 18950 6820
rect 18700 6780 18720 6815
rect 18920 6780 18940 6815
rect 18690 6770 18730 6780
rect 18585 6760 18625 6765
rect 18585 6730 18590 6760
rect 18620 6730 18625 6760
rect 18690 6750 18700 6770
rect 18720 6750 18730 6770
rect 18910 6770 18950 6780
rect 18690 6740 18730 6750
rect 18805 6760 18845 6765
rect 18585 6725 18625 6730
rect 18805 6730 18810 6760
rect 18840 6730 18845 6760
rect 18910 6750 18920 6770
rect 18940 6750 18950 6770
rect 19035 6765 19055 6870
rect 19745 6855 19765 6925
rect 19885 6910 19905 6925
rect 19875 6905 19915 6910
rect 19875 6875 19880 6905
rect 19910 6875 19915 6905
rect 19875 6870 19915 6875
rect 19140 6850 19180 6855
rect 19140 6820 19145 6850
rect 19175 6820 19180 6850
rect 19140 6815 19180 6820
rect 19730 6850 19770 6855
rect 19730 6820 19735 6850
rect 19765 6820 19770 6850
rect 19730 6815 19770 6820
rect 19950 6850 19990 6855
rect 19950 6820 19955 6850
rect 19985 6820 19990 6850
rect 19950 6815 19990 6820
rect 20180 6850 20220 6855
rect 20180 6820 20185 6850
rect 20215 6820 20220 6850
rect 20180 6815 20220 6820
rect 19150 6780 19170 6815
rect 19320 6805 19360 6810
rect 19140 6770 19180 6780
rect 19320 6775 19325 6805
rect 19355 6775 19360 6805
rect 19320 6770 19360 6775
rect 19440 6805 19480 6810
rect 19440 6775 19445 6805
rect 19475 6775 19480 6805
rect 19740 6780 19760 6815
rect 19960 6780 19980 6815
rect 20190 6780 20210 6815
rect 19440 6770 19480 6775
rect 19730 6770 19770 6780
rect 18910 6740 18950 6750
rect 19025 6760 19065 6765
rect 18805 6725 18845 6730
rect 19025 6730 19030 6760
rect 19060 6730 19065 6760
rect 19140 6750 19150 6770
rect 19170 6750 19180 6770
rect 19140 6740 19180 6750
rect 19025 6725 19065 6730
rect 19330 6720 19350 6770
rect 19450 6720 19470 6770
rect 19625 6760 19665 6765
rect 19625 6730 19630 6760
rect 19660 6730 19665 6760
rect 19730 6750 19740 6770
rect 19760 6750 19770 6770
rect 19950 6770 19990 6780
rect 19730 6740 19770 6750
rect 19845 6760 19885 6765
rect 19625 6725 19665 6730
rect 19845 6730 19850 6760
rect 19880 6730 19885 6760
rect 19950 6750 19960 6770
rect 19980 6750 19990 6770
rect 20180 6770 20220 6780
rect 19950 6740 19990 6750
rect 20065 6760 20105 6765
rect 19845 6725 19885 6730
rect 20065 6730 20070 6760
rect 20100 6730 20105 6760
rect 20180 6750 20190 6770
rect 20210 6750 20220 6770
rect 20180 6740 20220 6750
rect 20065 6725 20105 6730
rect 18737 6715 18769 6720
rect 18737 6685 18740 6715
rect 18766 6685 18769 6715
rect 18737 6680 18769 6685
rect 18957 6715 18989 6720
rect 18957 6685 18960 6715
rect 18986 6685 18989 6715
rect 18957 6680 18989 6685
rect 19101 6715 19133 6720
rect 19101 6685 19104 6715
rect 19130 6685 19133 6715
rect 19101 6680 19133 6685
rect 19320 6710 19350 6720
rect 19320 6690 19325 6710
rect 19345 6690 19350 6710
rect 19320 6680 19350 6690
rect 19367 6715 19399 6720
rect 19367 6685 19370 6715
rect 19396 6685 19399 6715
rect 19367 6680 19399 6685
rect 19450 6710 19480 6720
rect 19450 6690 19455 6710
rect 19475 6690 19480 6710
rect 19450 6680 19480 6690
rect 19777 6715 19809 6720
rect 19777 6685 19780 6715
rect 19806 6685 19809 6715
rect 19777 6680 19809 6685
rect 19997 6715 20029 6720
rect 19997 6685 20000 6715
rect 20026 6685 20029 6715
rect 19997 6680 20029 6685
rect 20141 6715 20173 6720
rect 20141 6685 20144 6715
rect 20170 6685 20173 6715
rect 20141 6680 20173 6685
rect 20325 6575 20345 7290
rect 20480 7285 20500 7340
rect 20640 7320 20685 7345
rect 20640 7285 20645 7320
rect 20680 7285 20685 7320
rect 21475 7285 21480 7320
rect 21515 7285 21520 7320
rect 20473 7280 20507 7285
rect 20473 7250 20476 7280
rect 20504 7250 20507 7280
rect 20473 7245 20507 7250
rect 21500 7225 21520 7285
rect 20500 7220 20540 7225
rect 20500 7190 20505 7220
rect 20535 7190 20540 7220
rect 20500 7185 20540 7190
rect 20610 7220 20650 7225
rect 20610 7190 20615 7220
rect 20645 7190 20650 7220
rect 20610 7185 20650 7190
rect 20720 7220 20760 7225
rect 20720 7190 20725 7220
rect 20755 7190 20760 7220
rect 20720 7185 20760 7190
rect 20830 7220 20870 7225
rect 20830 7190 20835 7220
rect 20865 7190 20870 7220
rect 20830 7185 20870 7190
rect 20940 7220 20980 7225
rect 20940 7190 20945 7220
rect 20975 7190 20980 7220
rect 20940 7185 20980 7190
rect 21050 7220 21090 7225
rect 21050 7190 21055 7220
rect 21085 7190 21090 7220
rect 21050 7185 21090 7190
rect 21160 7220 21200 7225
rect 21160 7190 21165 7220
rect 21195 7190 21200 7220
rect 21160 7185 21200 7190
rect 21270 7220 21310 7225
rect 21270 7190 21275 7220
rect 21305 7190 21310 7220
rect 21270 7185 21310 7190
rect 21380 7220 21420 7225
rect 21380 7190 21385 7220
rect 21415 7190 21420 7220
rect 21380 7185 21420 7190
rect 21490 7220 21530 7225
rect 21490 7190 21495 7220
rect 21525 7190 21530 7220
rect 21490 7185 21530 7190
rect 20445 7000 20485 7005
rect 20445 6970 20450 7000
rect 20480 6970 20485 7000
rect 20445 6965 20485 6970
rect 20555 7000 20595 7005
rect 20555 6970 20560 7000
rect 20590 6970 20595 7000
rect 20555 6965 20595 6970
rect 20665 7000 20705 7005
rect 20665 6970 20670 7000
rect 20700 6970 20705 7000
rect 20665 6965 20705 6970
rect 20775 7000 20815 7005
rect 20775 6970 20780 7000
rect 20810 6970 20815 7000
rect 20775 6965 20815 6970
rect 20885 7000 20925 7005
rect 20885 6970 20890 7000
rect 20920 6970 20925 7000
rect 20885 6965 20925 6970
rect 20995 7000 21035 7005
rect 20995 6970 21000 7000
rect 21030 6970 21035 7000
rect 20995 6965 21035 6970
rect 21105 7000 21145 7005
rect 21105 6970 21110 7000
rect 21140 6970 21145 7000
rect 21105 6965 21145 6970
rect 21215 7000 21255 7005
rect 21215 6970 21220 7000
rect 21250 6970 21255 7000
rect 21215 6965 21255 6970
rect 21325 7000 21365 7005
rect 21325 6970 21330 7000
rect 21360 6970 21365 7000
rect 21325 6965 21365 6970
rect 21435 7000 21475 7005
rect 21435 6970 21440 7000
rect 21470 6970 21475 7000
rect 21435 6965 21475 6970
rect 21545 7000 21585 7005
rect 21545 6970 21550 7000
rect 21580 6970 21585 7000
rect 21545 6965 21585 6970
rect 20545 6905 20585 6910
rect 20545 6875 20550 6905
rect 20580 6875 20585 6905
rect 20545 6870 20585 6875
rect 20655 6905 20695 6910
rect 20655 6875 20660 6905
rect 20690 6875 20695 6905
rect 20655 6870 20695 6875
rect 20765 6905 20805 6910
rect 20765 6875 20770 6905
rect 20800 6875 20805 6905
rect 20765 6870 20805 6875
rect 20566 6680 20598 6685
rect 20566 6650 20570 6680
rect 20596 6650 20598 6680
rect 20615 6680 20655 6690
rect 20615 6660 20625 6680
rect 20645 6660 20655 6680
rect 20615 6650 20655 6660
rect 20710 6680 20750 6690
rect 20710 6660 20720 6680
rect 20740 6660 20750 6680
rect 20710 6650 20750 6660
rect 20566 6645 20598 6650
rect 20510 6630 20550 6635
rect 20510 6600 20515 6630
rect 20545 6600 20550 6630
rect 20510 6595 20550 6600
rect 20570 6575 20590 6645
rect 20625 6635 20645 6650
rect 20720 6635 20740 6650
rect 20616 6630 20656 6635
rect 20616 6600 20621 6630
rect 20651 6600 20656 6630
rect 20616 6595 20656 6600
rect 20710 6630 20750 6635
rect 20710 6600 20715 6630
rect 20745 6600 20750 6630
rect 20710 6595 20750 6600
rect 20800 6630 20840 6635
rect 20800 6600 20805 6630
rect 20835 6600 20840 6630
rect 20800 6595 20840 6600
rect 12815 6570 12855 6575
rect 12815 6540 12820 6570
rect 12850 6540 12855 6570
rect 12815 6535 12855 6540
rect 20315 6570 20355 6575
rect 20315 6540 20320 6570
rect 20350 6540 20355 6570
rect 20315 6535 20355 6540
rect 20471 6570 20503 6575
rect 20471 6540 20475 6570
rect 20501 6540 20503 6570
rect 20471 6535 20503 6540
rect 20560 6565 20600 6575
rect 20560 6545 20570 6565
rect 20590 6545 20600 6565
rect 20560 6535 20600 6545
rect 20847 6570 20879 6575
rect 20847 6540 20849 6570
rect 20875 6540 20879 6570
rect 20847 6535 20879 6540
rect 11106 6495 11138 6500
rect 11106 6465 11109 6495
rect 11135 6465 11138 6495
rect 11106 6460 11138 6465
rect 11305 6495 11345 6500
rect 11305 6465 11310 6495
rect 11340 6465 11345 6495
rect 11305 6460 11345 6465
rect 11525 6495 11565 6500
rect 11525 6465 11530 6495
rect 11560 6465 11565 6495
rect 11525 6460 11565 6465
rect 11825 6490 11855 6500
rect 11825 6470 11830 6490
rect 11850 6470 11855 6490
rect 11825 6460 11855 6470
rect 11875 6490 11905 6500
rect 11875 6470 11880 6490
rect 11900 6470 11905 6490
rect 11875 6460 11905 6470
rect 11922 6495 11954 6500
rect 11922 6465 11925 6495
rect 11951 6465 11954 6495
rect 11922 6460 11954 6465
rect 12146 6495 12178 6500
rect 12146 6465 12149 6495
rect 12175 6465 12178 6495
rect 12146 6460 12178 6465
rect 12345 6495 12385 6500
rect 12345 6465 12350 6495
rect 12380 6465 12385 6495
rect 12345 6460 12385 6465
rect 12565 6495 12605 6500
rect 12565 6465 12570 6495
rect 12600 6465 12605 6495
rect 12565 6460 12605 6465
rect 18606 6495 18638 6500
rect 18606 6465 18609 6495
rect 18635 6465 18638 6495
rect 18606 6460 18638 6465
rect 18805 6495 18845 6500
rect 18805 6465 18810 6495
rect 18840 6465 18845 6495
rect 18805 6460 18845 6465
rect 19025 6495 19065 6500
rect 19025 6465 19030 6495
rect 19060 6465 19065 6495
rect 19025 6460 19065 6465
rect 19325 6490 19355 6500
rect 19325 6470 19330 6490
rect 19350 6470 19355 6490
rect 19325 6460 19355 6470
rect 19375 6490 19405 6500
rect 19375 6470 19380 6490
rect 19400 6470 19405 6490
rect 19375 6460 19405 6470
rect 19422 6495 19454 6500
rect 19422 6465 19425 6495
rect 19451 6465 19454 6495
rect 19422 6460 19454 6465
rect 19646 6495 19678 6500
rect 19646 6465 19649 6495
rect 19675 6465 19678 6495
rect 19646 6460 19678 6465
rect 19845 6495 19885 6500
rect 19845 6465 19850 6495
rect 19880 6465 19885 6495
rect 19845 6460 19885 6465
rect 20065 6495 20105 6500
rect 20065 6465 20070 6495
rect 20100 6465 20105 6495
rect 20065 6460 20105 6465
rect 9760 6410 9765 6445
rect 9800 6410 9805 6445
rect 10770 6410 10775 6445
rect 10810 6410 10815 6445
rect 11145 6435 11185 6440
rect 9775 6340 9795 6410
rect 10780 6395 10800 6410
rect 11145 6405 11150 6435
rect 11180 6405 11185 6435
rect 11145 6400 11185 6405
rect 11250 6435 11290 6440
rect 11250 6405 11255 6435
rect 11285 6405 11290 6435
rect 11250 6400 11290 6405
rect 11360 6435 11400 6440
rect 11360 6405 11365 6435
rect 11395 6405 11400 6435
rect 11360 6400 11400 6405
rect 11470 6435 11510 6440
rect 11470 6405 11475 6435
rect 11505 6405 11510 6435
rect 11470 6400 11510 6405
rect 11580 6435 11620 6440
rect 11580 6405 11585 6435
rect 11615 6405 11620 6435
rect 11580 6400 11620 6405
rect 10665 6390 10705 6395
rect 10665 6360 10670 6390
rect 10700 6360 10705 6390
rect 10665 6355 10705 6360
rect 10770 6390 10810 6395
rect 10770 6360 10775 6390
rect 10805 6360 10810 6390
rect 10770 6355 10810 6360
rect 10675 6340 10695 6355
rect 11830 6350 11850 6460
rect 11810 6345 11850 6350
rect 9765 6335 9805 6340
rect 9765 6305 9770 6335
rect 9800 6305 9805 6335
rect 9765 6300 9805 6305
rect 9965 6335 10005 6340
rect 9965 6305 9970 6335
rect 10000 6305 10005 6335
rect 9965 6300 10005 6305
rect 10165 6335 10205 6340
rect 10165 6305 10170 6335
rect 10200 6305 10205 6335
rect 10165 6300 10205 6305
rect 10365 6335 10405 6340
rect 10365 6305 10370 6335
rect 10400 6305 10405 6335
rect 10365 6300 10405 6305
rect 10565 6335 10605 6340
rect 10565 6305 10570 6335
rect 10600 6305 10605 6335
rect 10565 6300 10605 6305
rect 10668 6330 10702 6340
rect 10668 6310 10676 6330
rect 10694 6310 10702 6330
rect 10668 6300 10702 6310
rect 10765 6335 10805 6340
rect 10765 6305 10770 6335
rect 10800 6305 10805 6335
rect 11810 6315 11815 6345
rect 11845 6315 11850 6345
rect 11810 6310 11850 6315
rect 10765 6300 10805 6305
rect 11315 6295 11355 6300
rect 11315 6265 11320 6295
rect 11350 6265 11355 6295
rect 11315 6260 11355 6265
rect 11325 6240 11345 6260
rect 11820 6240 11840 6310
rect 11880 6300 11900 6460
rect 12185 6435 12225 6440
rect 12185 6405 12190 6435
rect 12220 6405 12225 6435
rect 12185 6400 12225 6405
rect 12290 6435 12330 6440
rect 12290 6405 12295 6435
rect 12325 6405 12330 6435
rect 12290 6400 12330 6405
rect 12400 6435 12440 6440
rect 12400 6405 12405 6435
rect 12435 6405 12440 6435
rect 12400 6400 12440 6405
rect 12510 6435 12550 6440
rect 12510 6405 12515 6435
rect 12545 6405 12550 6435
rect 12510 6400 12550 6405
rect 12620 6435 12660 6440
rect 12620 6405 12625 6435
rect 12655 6405 12660 6435
rect 12985 6410 12990 6445
rect 13025 6410 13030 6445
rect 13995 6410 14000 6445
rect 14035 6410 14040 6445
rect 18645 6435 18685 6440
rect 12620 6400 12660 6405
rect 13000 6395 13020 6410
rect 12990 6390 13030 6395
rect 12990 6360 12995 6390
rect 13025 6360 13030 6390
rect 12990 6355 13030 6360
rect 13095 6390 13135 6395
rect 13095 6360 13100 6390
rect 13130 6360 13135 6390
rect 13095 6355 13135 6360
rect 13105 6340 13125 6355
rect 14005 6340 14025 6410
rect 18645 6405 18650 6435
rect 18680 6405 18685 6435
rect 18645 6400 18685 6405
rect 18750 6435 18790 6440
rect 18750 6405 18755 6435
rect 18785 6405 18790 6435
rect 18750 6400 18790 6405
rect 18860 6435 18900 6440
rect 18860 6405 18865 6435
rect 18895 6405 18900 6435
rect 18860 6400 18900 6405
rect 18970 6435 19010 6440
rect 18970 6405 18975 6435
rect 19005 6405 19010 6435
rect 18970 6400 19010 6405
rect 19080 6435 19120 6440
rect 19080 6405 19085 6435
rect 19115 6405 19120 6435
rect 19080 6400 19120 6405
rect 19330 6390 19350 6460
rect 19310 6385 19350 6390
rect 19310 6355 19315 6385
rect 19345 6355 19350 6385
rect 19310 6350 19350 6355
rect 12995 6335 13035 6340
rect 12995 6305 13000 6335
rect 13030 6305 13035 6335
rect 12995 6300 13035 6305
rect 13098 6330 13132 6340
rect 13098 6310 13106 6330
rect 13124 6310 13132 6330
rect 13098 6300 13132 6310
rect 13195 6335 13235 6340
rect 13195 6305 13200 6335
rect 13230 6305 13235 6335
rect 13195 6300 13235 6305
rect 13395 6335 13435 6340
rect 13395 6305 13400 6335
rect 13430 6305 13435 6335
rect 13395 6300 13435 6305
rect 13595 6335 13635 6340
rect 13595 6305 13600 6335
rect 13630 6305 13635 6335
rect 13595 6300 13635 6305
rect 13795 6335 13835 6340
rect 13795 6305 13800 6335
rect 13830 6305 13835 6335
rect 13795 6300 13835 6305
rect 13995 6335 14035 6340
rect 13995 6305 14000 6335
rect 14030 6305 14035 6335
rect 13995 6300 14035 6305
rect 18815 6335 18855 6340
rect 18815 6305 18820 6335
rect 18850 6305 18855 6335
rect 18815 6300 18855 6305
rect 11880 6295 11920 6300
rect 11880 6265 11885 6295
rect 11915 6265 11920 6295
rect 18825 6280 18845 6300
rect 19320 6280 19340 6350
rect 19380 6340 19400 6460
rect 19685 6435 19725 6440
rect 19685 6405 19690 6435
rect 19720 6405 19725 6435
rect 19685 6400 19725 6405
rect 19790 6435 19830 6440
rect 19790 6405 19795 6435
rect 19825 6405 19830 6435
rect 19790 6400 19830 6405
rect 19900 6435 19940 6440
rect 19900 6405 19905 6435
rect 19935 6405 19940 6435
rect 19900 6400 19940 6405
rect 20010 6435 20050 6440
rect 20010 6405 20015 6435
rect 20045 6405 20050 6435
rect 20010 6400 20050 6405
rect 20120 6435 20160 6440
rect 20120 6405 20125 6435
rect 20155 6405 20160 6435
rect 20120 6400 20160 6405
rect 20526 6350 20558 6355
rect 19380 6335 19420 6340
rect 19380 6305 19385 6335
rect 19415 6305 19420 6335
rect 20526 6320 20528 6350
rect 20554 6320 20558 6350
rect 20526 6315 20558 6320
rect 20792 6350 20824 6355
rect 20792 6320 20796 6350
rect 20822 6320 20824 6350
rect 20792 6315 20824 6320
rect 19380 6300 19420 6305
rect 20095 6290 20135 6295
rect 11880 6260 11920 6265
rect 18815 6270 18855 6280
rect 12595 6250 12635 6255
rect 11315 6230 11355 6240
rect 11315 6210 11325 6230
rect 11345 6210 11355 6230
rect 11315 6200 11355 6210
rect 11425 6235 11465 6240
rect 11425 6205 11430 6235
rect 11460 6205 11465 6235
rect 11425 6200 11465 6205
rect 11535 6235 11575 6240
rect 11535 6205 11540 6235
rect 11570 6205 11575 6235
rect 11535 6200 11575 6205
rect 11645 6235 11685 6240
rect 11645 6205 11650 6235
rect 11680 6205 11685 6235
rect 11645 6200 11685 6205
rect 11755 6235 11795 6240
rect 11755 6205 11760 6235
rect 11790 6205 11795 6235
rect 11755 6200 11795 6205
rect 11815 6230 11845 6240
rect 11815 6210 11820 6230
rect 11840 6210 11845 6230
rect 11815 6200 11845 6210
rect 11865 6235 11905 6240
rect 11865 6205 11870 6235
rect 11900 6205 11905 6235
rect 11865 6200 11905 6205
rect 11975 6235 12015 6240
rect 11975 6205 11980 6235
rect 12010 6205 12015 6235
rect 11975 6200 12015 6205
rect 12085 6235 12125 6240
rect 12085 6205 12090 6235
rect 12120 6205 12125 6235
rect 12085 6200 12125 6205
rect 12195 6235 12235 6240
rect 12195 6205 12200 6235
rect 12230 6205 12235 6235
rect 12195 6200 12235 6205
rect 12305 6235 12345 6240
rect 12305 6205 12310 6235
rect 12340 6205 12345 6235
rect 12305 6200 12345 6205
rect 12415 6235 12455 6240
rect 12415 6205 12420 6235
rect 12450 6205 12455 6235
rect 12415 6200 12455 6205
rect 12525 6235 12565 6240
rect 12525 6205 12530 6235
rect 12560 6205 12565 6235
rect 12595 6220 12600 6250
rect 12630 6220 12635 6250
rect 18815 6250 18825 6270
rect 18845 6250 18855 6270
rect 18815 6240 18855 6250
rect 18925 6275 18965 6280
rect 18925 6245 18930 6275
rect 18960 6245 18965 6275
rect 18925 6240 18965 6245
rect 19035 6275 19075 6280
rect 19035 6245 19040 6275
rect 19070 6245 19075 6275
rect 19035 6240 19075 6245
rect 19145 6275 19185 6280
rect 19145 6245 19150 6275
rect 19180 6245 19185 6275
rect 19145 6240 19185 6245
rect 19255 6275 19295 6280
rect 19255 6245 19260 6275
rect 19290 6245 19295 6275
rect 19255 6240 19295 6245
rect 19315 6270 19345 6280
rect 19315 6250 19320 6270
rect 19340 6250 19345 6270
rect 19315 6240 19345 6250
rect 19365 6275 19405 6280
rect 19365 6245 19370 6275
rect 19400 6245 19405 6275
rect 19365 6240 19405 6245
rect 19475 6275 19515 6280
rect 19475 6245 19480 6275
rect 19510 6245 19515 6275
rect 19475 6240 19515 6245
rect 19585 6275 19625 6280
rect 19585 6245 19590 6275
rect 19620 6245 19625 6275
rect 19585 6240 19625 6245
rect 19695 6275 19735 6280
rect 19695 6245 19700 6275
rect 19730 6245 19735 6275
rect 19695 6240 19735 6245
rect 19805 6275 19845 6280
rect 19805 6245 19810 6275
rect 19840 6245 19845 6275
rect 19805 6240 19845 6245
rect 19915 6275 19955 6280
rect 19915 6245 19920 6275
rect 19950 6245 19955 6275
rect 19915 6240 19955 6245
rect 20025 6275 20065 6280
rect 20025 6245 20030 6275
rect 20060 6245 20065 6275
rect 20095 6260 20100 6290
rect 20130 6260 20135 6290
rect 20095 6255 20135 6260
rect 20445 6290 20485 6295
rect 20445 6260 20450 6290
rect 20480 6260 20485 6290
rect 20445 6255 20485 6260
rect 20560 6290 20600 6295
rect 20560 6260 20565 6290
rect 20595 6260 20600 6290
rect 20560 6255 20600 6260
rect 20655 6290 20695 6295
rect 20655 6260 20660 6290
rect 20690 6260 20695 6290
rect 20655 6255 20695 6260
rect 20750 6290 20790 6295
rect 20750 6260 20755 6290
rect 20785 6260 20790 6290
rect 20750 6255 20790 6260
rect 20865 6290 20905 6295
rect 20865 6260 20870 6290
rect 20900 6260 20905 6290
rect 20865 6255 20905 6260
rect 20025 6240 20065 6245
rect 20665 6235 20685 6255
rect 20875 6235 20895 6255
rect 12595 6215 12635 6220
rect 20600 6230 20640 6235
rect 12525 6200 12565 6205
rect 20600 6200 20605 6230
rect 20635 6200 20640 6230
rect 20600 6195 20640 6200
rect 20660 6230 20690 6235
rect 20660 6195 20690 6200
rect 20710 6230 20750 6235
rect 20710 6200 20715 6230
rect 20745 6200 20750 6230
rect 20710 6195 20750 6200
rect 20865 6230 20905 6235
rect 20865 6200 20870 6230
rect 20900 6200 20905 6230
rect 20865 6195 20905 6200
rect 9865 5985 9905 5990
rect 9865 5955 9870 5985
rect 9900 5955 9905 5985
rect 9865 5950 9905 5955
rect 10065 5985 10105 5990
rect 10065 5955 10070 5985
rect 10100 5955 10105 5985
rect 10065 5950 10105 5955
rect 10265 5985 10305 5990
rect 10265 5955 10270 5985
rect 10300 5955 10305 5985
rect 10265 5950 10305 5955
rect 10465 5985 10505 5990
rect 10465 5955 10470 5985
rect 10500 5955 10505 5985
rect 10465 5950 10505 5955
rect 10665 5985 10705 5990
rect 10665 5955 10670 5985
rect 10700 5955 10705 5985
rect 10665 5950 10705 5955
rect 13095 5985 13135 5990
rect 13095 5955 13100 5985
rect 13130 5955 13135 5985
rect 13095 5950 13135 5955
rect 13295 5985 13335 5990
rect 13295 5955 13300 5985
rect 13330 5955 13335 5985
rect 13295 5950 13335 5955
rect 13495 5985 13535 5990
rect 13495 5955 13500 5985
rect 13530 5955 13535 5985
rect 13495 5950 13535 5955
rect 13695 5985 13735 5990
rect 13695 5955 13700 5985
rect 13730 5955 13735 5985
rect 13695 5950 13735 5955
rect 13895 5985 13935 5990
rect 13895 5955 13900 5985
rect 13930 5955 13935 5985
rect 13895 5950 13935 5955
rect 18665 5955 18705 5960
rect 18665 5925 18670 5955
rect 18700 5925 18705 5955
rect 18665 5920 18705 5925
rect 18760 5955 18800 5960
rect 18760 5925 18765 5955
rect 18795 5925 18800 5955
rect 18760 5920 18800 5925
rect 18870 5955 18910 5960
rect 18870 5925 18875 5955
rect 18905 5925 18910 5955
rect 18870 5920 18910 5925
rect 18980 5955 19020 5960
rect 18980 5925 18985 5955
rect 19015 5925 19020 5955
rect 18980 5920 19020 5925
rect 19090 5955 19130 5960
rect 19090 5925 19095 5955
rect 19125 5925 19130 5955
rect 19090 5920 19130 5925
rect 19200 5955 19240 5960
rect 19200 5925 19205 5955
rect 19235 5925 19240 5955
rect 19200 5920 19240 5925
rect 19310 5955 19350 5960
rect 19310 5925 19315 5955
rect 19345 5925 19350 5955
rect 19310 5920 19350 5925
rect 19420 5955 19460 5960
rect 19420 5925 19425 5955
rect 19455 5925 19460 5955
rect 19420 5920 19460 5925
rect 19530 5955 19570 5960
rect 19530 5925 19535 5955
rect 19565 5925 19570 5955
rect 19530 5920 19570 5925
rect 19640 5955 19680 5960
rect 19640 5925 19645 5955
rect 19675 5925 19680 5955
rect 19640 5920 19680 5925
rect 19750 5955 19790 5960
rect 19750 5925 19755 5955
rect 19785 5925 19790 5955
rect 19750 5920 19790 5925
rect 19860 5955 19900 5960
rect 19860 5925 19865 5955
rect 19895 5925 19900 5955
rect 19860 5920 19900 5925
rect 19970 5955 20010 5960
rect 19970 5925 19975 5955
rect 20005 5925 20010 5955
rect 19970 5920 20010 5925
rect 20120 5955 20160 5960
rect 20120 5925 20125 5955
rect 20155 5925 20160 5955
rect 20120 5920 20160 5925
rect 11165 5915 11205 5920
rect 11165 5885 11170 5915
rect 11200 5885 11205 5915
rect 11165 5880 11205 5885
rect 11260 5915 11300 5920
rect 11260 5885 11265 5915
rect 11295 5885 11300 5915
rect 11260 5880 11300 5885
rect 11370 5915 11410 5920
rect 11370 5885 11375 5915
rect 11405 5885 11410 5915
rect 11370 5880 11410 5885
rect 11480 5915 11520 5920
rect 11480 5885 11485 5915
rect 11515 5885 11520 5915
rect 11480 5880 11520 5885
rect 11590 5915 11630 5920
rect 11590 5885 11595 5915
rect 11625 5885 11630 5915
rect 11590 5880 11630 5885
rect 11700 5915 11740 5920
rect 11700 5885 11705 5915
rect 11735 5885 11740 5915
rect 11700 5880 11740 5885
rect 11810 5915 11850 5920
rect 11810 5885 11815 5915
rect 11845 5885 11850 5915
rect 11810 5880 11850 5885
rect 11920 5915 11960 5920
rect 11920 5885 11925 5915
rect 11955 5885 11960 5915
rect 11920 5880 11960 5885
rect 12030 5915 12070 5920
rect 12030 5885 12035 5915
rect 12065 5885 12070 5915
rect 12030 5880 12070 5885
rect 12140 5915 12180 5920
rect 12140 5885 12145 5915
rect 12175 5885 12180 5915
rect 12140 5880 12180 5885
rect 12250 5915 12290 5920
rect 12250 5885 12255 5915
rect 12285 5885 12290 5915
rect 12250 5880 12290 5885
rect 12360 5915 12400 5920
rect 12360 5885 12365 5915
rect 12395 5885 12400 5915
rect 12360 5880 12400 5885
rect 12470 5915 12510 5920
rect 12470 5885 12475 5915
rect 12505 5885 12510 5915
rect 12470 5880 12510 5885
rect 12620 5915 12660 5920
rect 12620 5885 12625 5915
rect 12655 5885 12660 5915
rect 12620 5880 12660 5885
rect 11632 4515 11668 4520
rect 11632 4485 11635 4515
rect 11665 4485 11668 4515
rect 11632 4480 11668 4485
rect 11752 4515 11788 4520
rect 11752 4485 11755 4515
rect 11785 4485 11788 4515
rect 11752 4480 11788 4485
rect 11872 4515 11908 4520
rect 11872 4485 11875 4515
rect 11905 4485 11908 4515
rect 11872 4480 11908 4485
rect 12080 4515 12120 4520
rect 12080 4485 12085 4515
rect 12115 4485 12120 4515
rect 12080 4480 12120 4485
rect 11570 4470 11610 4475
rect 11200 4455 11240 4460
rect 11200 4425 11205 4455
rect 11235 4425 11240 4455
rect 11200 4420 11240 4425
rect 11460 4455 11500 4460
rect 11460 4425 11465 4455
rect 11495 4425 11500 4455
rect 11570 4440 11575 4470
rect 11605 4440 11610 4470
rect 11570 4435 11610 4440
rect 11690 4470 11730 4475
rect 11690 4440 11695 4470
rect 11725 4440 11730 4470
rect 11690 4435 11730 4440
rect 11810 4470 11850 4475
rect 11810 4440 11815 4470
rect 11845 4440 11850 4470
rect 11810 4435 11850 4440
rect 11930 4470 11970 4475
rect 11930 4440 11935 4470
rect 11965 4440 11970 4470
rect 12090 4450 12110 4480
rect 11930 4435 11970 4440
rect 12080 4445 12120 4450
rect 11460 4420 11500 4425
rect 12080 4415 12085 4445
rect 12115 4415 12120 4445
rect 12080 4410 12120 4415
rect 12200 4445 12240 4450
rect 12200 4415 12205 4445
rect 12235 4415 12240 4445
rect 12200 4410 12240 4415
rect 12320 4445 12360 4450
rect 12320 4415 12325 4445
rect 12355 4415 12360 4445
rect 12320 4410 12360 4415
rect 12440 4445 12480 4450
rect 12440 4415 12445 4445
rect 12475 4415 12480 4445
rect 12440 4410 12480 4415
rect 12560 4445 12600 4450
rect 12560 4415 12565 4445
rect 12595 4415 12600 4445
rect 12560 4410 12600 4415
rect 11330 4320 11370 4325
rect 11050 4315 11090 4320
rect 11050 4285 11055 4315
rect 11085 4285 11090 4315
rect 11330 4290 11335 4320
rect 11365 4290 11370 4320
rect 11330 4285 11370 4290
rect 11750 4315 11790 4320
rect 11750 4285 11755 4315
rect 11785 4285 11790 4315
rect 11050 4280 11090 4285
rect 10210 3635 10250 3640
rect 10210 3605 10215 3635
rect 10245 3605 10250 3635
rect 10210 3600 10250 3605
rect 10320 3635 10360 3640
rect 10320 3605 10325 3635
rect 10355 3605 10360 3635
rect 10320 3600 10360 3605
rect 10430 3635 10470 3640
rect 10430 3605 10435 3635
rect 10465 3605 10470 3635
rect 10430 3600 10470 3605
rect 10540 3635 10580 3640
rect 10540 3605 10545 3635
rect 10575 3605 10580 3635
rect 10540 3600 10580 3605
rect 10650 3635 10690 3640
rect 10650 3605 10655 3635
rect 10685 3605 10690 3635
rect 10650 3600 10690 3605
rect 10760 3635 10800 3640
rect 10760 3605 10765 3635
rect 10795 3605 10800 3635
rect 10760 3600 10800 3605
rect 9899 3555 10040 3560
rect 9899 3550 9905 3555
rect 9895 3530 9905 3550
rect 1261 3525 1301 3530
rect 1261 3495 1266 3525
rect 1296 3495 1301 3525
rect 9899 3525 9905 3530
rect 9935 3525 9955 3555
rect 9985 3525 10005 3555
rect 10035 3525 10040 3555
rect 9899 3520 10040 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3310 1245 3340
rect 1205 3305 1245 3310
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3255 1200 3285
rect 1160 3250 1200 3255
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 46 3110 51 3145
rect 86 3110 91 3145
rect 1170 3105 1190 3250
rect 1160 3100 1200 3105
rect 1160 3070 1165 3100
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 46 2970 51 3005
rect 86 2970 91 3005
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 1215 2855 1235 3305
rect 1271 3200 1291 3490
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 1635 3405 1685 3415
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 1271 3140 1291 3165
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 51 2820 56 2855
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2820 769 2855
rect 1205 2850 1245 2855
rect 1205 2820 1210 2850
rect 1240 2820 1245 2850
rect 2340 2840 2360 2860
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 51 2760 56 2795
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2760 769 2795
rect 1271 2750 1291 2805
rect 2330 2800 2370 2805
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2715 1301 2745
rect 1261 2710 1301 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 952 1710 1302 1870
rect 952 1680 1270 1710
rect 1297 1680 1302 1710
rect 952 1520 1302 1680
rect 1330 1190 1455 1345
rect 1635 1190 1985 2200
rect 2160 1190 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3135 3340 3175 3345
rect 3135 3310 3140 3340
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2735 3240 2775 3245
rect 2735 3210 2740 3240
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3155 2660 3185
rect 2620 3150 2660 3155
rect 2520 2980 2560 2985
rect 2520 2950 2525 2980
rect 2555 2950 2560 2980
rect 2520 2945 2560 2950
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 840 2180 1190
rect 2530 765 2550 2945
rect 2630 2795 2650 3150
rect 2620 2790 2660 2795
rect 2620 2760 2625 2790
rect 2655 2760 2660 2790
rect 2620 2755 2660 2760
rect 2630 2350 2650 2755
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2315 2660 2345
rect 2620 2310 2660 2315
rect 2630 2055 2650 2310
rect 2745 2295 2765 3205
rect 3145 3145 3165 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5360 3335 5400 3340
rect 5360 3305 5365 3335
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 4885 3285 4925 3290
rect 4885 3255 4890 3285
rect 4920 3255 4925 3285
rect 4885 3250 4925 3255
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 3135 3140 3175 3145
rect 3135 3110 3140 3140
rect 3170 3110 3175 3140
rect 3135 3105 3175 3110
rect 4835 3140 4875 3145
rect 4835 3110 4840 3140
rect 4870 3110 4875 3140
rect 4835 3105 4875 3110
rect 3145 2985 3165 3105
rect 3985 3080 4025 3085
rect 3985 3050 3990 3080
rect 4020 3050 4025 3080
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3005 3485 3035
rect 3445 3000 3485 3005
rect 3805 3035 3845 3040
rect 3805 3005 3810 3035
rect 3840 3005 3845 3035
rect 3805 3000 3845 3005
rect 3455 2985 3475 3000
rect 3815 2985 3835 3000
rect 3995 2985 4015 3045
rect 4345 3035 4385 3040
rect 4345 3005 4350 3035
rect 4380 3005 4385 3035
rect 4345 3000 4385 3005
rect 4705 3035 4745 3040
rect 4705 3005 4710 3035
rect 4740 3005 4745 3035
rect 4705 3000 4745 3005
rect 4355 2985 4375 3000
rect 4715 2985 4735 3000
rect 4845 2985 4865 3105
rect 4895 2985 4915 3250
rect 5315 3140 5355 3145
rect 5315 3110 5320 3140
rect 5350 3110 5355 3140
rect 5315 3105 5355 3110
rect 3080 2980 3120 2985
rect 3080 2950 3085 2980
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2950 3305 2980
rect 3265 2945 3305 2950
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2980 3665 2985
rect 3625 2950 3630 2980
rect 3660 2950 3665 2980
rect 3625 2945 3665 2950
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2980 4205 2985
rect 4165 2950 4170 2980
rect 4200 2950 4205 2980
rect 4165 2945 4205 2950
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2980 4565 2985
rect 4525 2950 4530 2980
rect 4560 2950 4565 2980
rect 4525 2945 4565 2950
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 2995 2810 3035 2815
rect 2995 2780 3000 2810
rect 3030 2780 3035 2810
rect 2995 2775 3035 2780
rect 3175 2810 3215 2815
rect 3175 2780 3180 2810
rect 3210 2780 3215 2810
rect 3175 2775 3215 2780
rect 3355 2810 3395 2815
rect 3355 2780 3360 2810
rect 3390 2780 3395 2810
rect 3355 2775 3395 2780
rect 3535 2810 3575 2815
rect 3535 2780 3540 2810
rect 3570 2780 3575 2810
rect 3535 2775 3575 2780
rect 3715 2810 3755 2815
rect 3715 2780 3720 2810
rect 3750 2780 3755 2810
rect 3715 2775 3755 2780
rect 3895 2810 3935 2815
rect 3895 2780 3900 2810
rect 3930 2780 3935 2810
rect 3895 2775 3935 2780
rect 4075 2810 4115 2815
rect 4075 2780 4080 2810
rect 4110 2780 4115 2810
rect 4075 2775 4115 2780
rect 4255 2810 4295 2815
rect 4255 2780 4260 2810
rect 4290 2780 4295 2810
rect 4255 2775 4295 2780
rect 4435 2810 4475 2815
rect 4435 2780 4440 2810
rect 4470 2780 4475 2810
rect 4435 2775 4475 2780
rect 4615 2810 4655 2815
rect 4615 2780 4620 2810
rect 4650 2780 4655 2810
rect 4615 2775 4655 2780
rect 4795 2810 4835 2815
rect 4795 2780 4800 2810
rect 4830 2780 4835 2810
rect 4795 2775 4835 2780
rect 4975 2810 5015 2815
rect 4975 2780 4980 2810
rect 5010 2780 5015 2810
rect 4975 2775 5015 2780
rect 4805 2755 4825 2775
rect 3175 2750 3215 2755
rect 3175 2720 3180 2750
rect 3210 2720 3215 2750
rect 3175 2715 3215 2720
rect 3355 2750 3395 2755
rect 3355 2720 3360 2750
rect 3390 2720 3395 2750
rect 3355 2715 3395 2720
rect 3535 2750 3575 2755
rect 3535 2720 3540 2750
rect 3570 2720 3575 2750
rect 3535 2715 3575 2720
rect 3715 2750 3755 2755
rect 3715 2720 3720 2750
rect 3750 2720 3755 2750
rect 3715 2715 3755 2720
rect 3895 2750 3935 2755
rect 3895 2720 3900 2750
rect 3930 2720 3935 2750
rect 3895 2715 3935 2720
rect 4075 2750 4115 2755
rect 4075 2720 4080 2750
rect 4110 2720 4115 2750
rect 4075 2715 4115 2720
rect 4255 2750 4295 2755
rect 4255 2720 4260 2750
rect 4290 2720 4295 2750
rect 4255 2715 4295 2720
rect 4435 2750 4475 2755
rect 4435 2720 4440 2750
rect 4470 2720 4475 2750
rect 4435 2715 4475 2720
rect 4615 2750 4655 2755
rect 4615 2720 4620 2750
rect 4650 2720 4655 2750
rect 4615 2715 4655 2720
rect 4795 2750 4835 2755
rect 4795 2720 4800 2750
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2375 3395 2380
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3805 2380 3845 2385
rect 3805 2350 3810 2380
rect 3840 2350 3845 2380
rect 3805 2345 3845 2350
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2380 4205 2385
rect 4165 2350 4170 2380
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2260 2775 2290
rect 2735 2255 2775 2260
rect 3275 2205 3295 2345
rect 3355 2340 3395 2345
rect 3455 2295 3475 2345
rect 3625 2335 3665 2340
rect 3625 2305 3630 2335
rect 3660 2305 3665 2335
rect 3625 2300 3665 2305
rect 3445 2290 3485 2295
rect 3445 2260 3450 2290
rect 3480 2260 3485 2290
rect 3445 2255 3485 2260
rect 3265 2200 3305 2205
rect 3265 2170 3270 2200
rect 3300 2170 3305 2200
rect 3265 2165 3305 2170
rect 3635 2155 3655 2300
rect 3815 2250 3835 2345
rect 3805 2245 3845 2250
rect 3805 2215 3810 2245
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 3625 2150 3665 2155
rect 3625 2120 3630 2150
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2065 2785 2095
rect 2745 2060 2785 2065
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2065 2905 2095
rect 2865 2060 2905 2065
rect 2985 2095 3025 2100
rect 2985 2065 2990 2095
rect 3020 2065 3025 2095
rect 2985 2060 3025 2065
rect 3105 2095 3145 2100
rect 3105 2065 3110 2095
rect 3140 2065 3145 2095
rect 3105 2060 3145 2065
rect 3225 2095 3265 2100
rect 3225 2065 3230 2095
rect 3260 2065 3265 2095
rect 3225 2060 3265 2065
rect 3345 2095 3385 2100
rect 3345 2065 3350 2095
rect 3380 2065 3385 2095
rect 3345 2060 3385 2065
rect 3465 2095 3505 2100
rect 3465 2065 3470 2095
rect 3500 2065 3505 2095
rect 3465 2060 3505 2065
rect 3585 2095 3625 2100
rect 3585 2065 3590 2095
rect 3620 2065 3625 2095
rect 3585 2060 3625 2065
rect 3705 2095 3745 2100
rect 3705 2065 3710 2095
rect 3740 2065 3745 2095
rect 3705 2060 3745 2065
rect 3825 2095 3865 2100
rect 3825 2065 3830 2095
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 3895 2055 3915 2345
rect 3995 2205 4015 2345
rect 4345 2335 4385 2340
rect 4345 2305 4350 2335
rect 4380 2305 4385 2335
rect 4345 2300 4385 2305
rect 4535 2295 4555 2345
rect 4525 2290 4565 2295
rect 4525 2260 4530 2290
rect 4560 2260 4565 2290
rect 4525 2255 4565 2260
rect 4715 2205 4735 2345
rect 5270 2290 5310 2295
rect 5270 2260 5275 2290
rect 5305 2260 5310 2290
rect 5270 2255 5310 2260
rect 3985 2200 4025 2205
rect 3985 2170 3990 2200
rect 4020 2170 4025 2200
rect 3985 2165 4025 2170
rect 4705 2200 4745 2205
rect 4705 2170 4710 2200
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2115 4125 2145
rect 4085 2110 4125 2115
rect 3985 2095 4025 2100
rect 3985 2065 3990 2095
rect 4020 2065 4025 2095
rect 3985 2060 4025 2065
rect 4095 2055 4115 2110
rect 4145 2095 4185 2100
rect 4145 2065 4150 2095
rect 4180 2065 4185 2095
rect 4145 2060 4185 2065
rect 4265 2095 4305 2100
rect 4265 2065 4270 2095
rect 4300 2065 4305 2095
rect 4265 2060 4305 2065
rect 4385 2095 4425 2100
rect 4385 2065 4390 2095
rect 4420 2065 4425 2095
rect 4385 2060 4425 2065
rect 4505 2095 4545 2100
rect 4505 2065 4510 2095
rect 4540 2065 4545 2095
rect 4505 2060 4545 2065
rect 4625 2095 4665 2100
rect 4625 2065 4630 2095
rect 4660 2065 4665 2095
rect 4625 2060 4665 2065
rect 4745 2095 4785 2100
rect 4745 2065 4750 2095
rect 4780 2065 4785 2095
rect 4745 2060 4785 2065
rect 4865 2095 4905 2100
rect 4865 2065 4870 2095
rect 4900 2065 4905 2095
rect 4865 2060 4905 2065
rect 4985 2095 5025 2100
rect 4985 2065 4990 2095
rect 5020 2065 5025 2095
rect 4985 2060 5025 2065
rect 5105 2095 5145 2100
rect 5105 2065 5110 2095
rect 5140 2065 5145 2095
rect 5105 2060 5145 2065
rect 5225 2095 5265 2100
rect 5225 2065 5230 2095
rect 5260 2065 5265 2095
rect 5225 2060 5265 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2020 2845 2050
rect 2805 2015 2845 2020
rect 3165 2050 3205 2055
rect 3165 2020 3170 2050
rect 3200 2020 3205 2050
rect 3165 2015 3205 2020
rect 3525 2050 3565 2055
rect 3525 2020 3530 2050
rect 3560 2020 3565 2050
rect 3525 2015 3565 2020
rect 3885 2050 3925 2055
rect 3885 2020 3890 2050
rect 3920 2045 3925 2050
rect 4085 2050 4125 2055
rect 4085 2045 4090 2050
rect 3920 2020 3945 2045
rect 3885 2015 3945 2020
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1850 2965 1880
rect 2925 1845 2965 1850
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1880 3325 1885
rect 3285 1850 3290 1880
rect 3320 1850 3325 1880
rect 3285 1845 3325 1850
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1880 3685 1885
rect 3645 1850 3650 1880
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 2575 1765 2595 1845
rect 2565 1760 2605 1765
rect 2565 1730 2570 1760
rect 2600 1730 2605 1760
rect 2565 1725 2605 1730
rect 2630 1670 2650 1845
rect 2685 1765 2705 1845
rect 2845 1825 2865 1845
rect 3055 1825 3075 1845
rect 3175 1825 3195 1845
rect 2835 1820 2875 1825
rect 2835 1790 2840 1820
rect 2870 1790 2875 1820
rect 2835 1785 2875 1790
rect 3045 1820 3085 1825
rect 3045 1790 3050 1820
rect 3080 1790 3085 1820
rect 3045 1785 3085 1790
rect 3165 1820 3205 1825
rect 3165 1790 3170 1820
rect 3200 1790 3205 1820
rect 3165 1785 3205 1790
rect 2800 1765 2840 1770
rect 3295 1765 3315 1845
rect 3415 1825 3435 1845
rect 3535 1825 3555 1845
rect 3775 1825 3795 1845
rect 3865 1825 3885 1845
rect 3405 1820 3445 1825
rect 3405 1790 3410 1820
rect 3440 1790 3445 1820
rect 3405 1785 3445 1790
rect 3525 1820 3565 1825
rect 3525 1790 3530 1820
rect 3560 1790 3565 1820
rect 3525 1785 3565 1790
rect 3765 1820 3805 1825
rect 3765 1790 3770 1820
rect 3800 1790 3805 1820
rect 3765 1785 3805 1790
rect 3855 1820 3895 1825
rect 3855 1790 3860 1820
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 2675 1760 2715 1765
rect 2675 1730 2680 1760
rect 2710 1730 2715 1760
rect 2800 1735 2805 1765
rect 2835 1735 2840 1765
rect 2800 1730 2840 1735
rect 3225 1760 3265 1765
rect 3225 1730 3230 1760
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 2810 1715 2830 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1730 3325 1760
rect 3285 1725 3325 1730
rect 3415 1720 3435 1785
rect 3525 1760 3565 1765
rect 3525 1730 3530 1760
rect 3560 1730 3565 1760
rect 3525 1725 3565 1730
rect 3765 1760 3805 1765
rect 3765 1730 3770 1760
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 3165 1715 3205 1720
rect 2800 1710 2840 1715
rect 2800 1680 2805 1710
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1685 3205 1715
rect 3165 1680 3205 1685
rect 3405 1715 3445 1720
rect 3405 1685 3410 1715
rect 3440 1685 3445 1715
rect 3405 1680 3445 1685
rect 3645 1715 3685 1720
rect 3645 1685 3650 1715
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 2800 1675 2840 1680
rect 2620 1665 2660 1670
rect 2620 1635 2625 1665
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2630 1045 2650 1630
rect 3165 1595 3205 1600
rect 3165 1565 3170 1595
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1515 2875 1545
rect 2835 1510 2875 1515
rect 3225 1545 3265 1550
rect 3225 1515 3230 1545
rect 3260 1515 3265 1545
rect 3225 1510 3265 1515
rect 3345 1545 3385 1550
rect 3345 1515 3350 1545
rect 3380 1515 3385 1545
rect 3345 1510 3385 1515
rect 3465 1545 3505 1550
rect 3465 1515 3470 1545
rect 3500 1515 3505 1545
rect 3465 1510 3505 1515
rect 3585 1545 3625 1550
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 3705 1545 3745 1550
rect 3705 1515 3710 1545
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 2845 1490 2865 1510
rect 2925 1500 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1470 2930 1500
rect 2960 1470 2965 1500
rect 2925 1465 2965 1470
rect 3045 1500 3085 1505
rect 3045 1470 3050 1500
rect 3080 1470 3085 1500
rect 3045 1465 3085 1470
rect 3165 1500 3205 1505
rect 3165 1470 3170 1500
rect 3200 1470 3205 1500
rect 3165 1465 3205 1470
rect 3285 1500 3325 1505
rect 3285 1470 3290 1500
rect 3320 1470 3325 1500
rect 3285 1465 3325 1470
rect 3525 1500 3565 1505
rect 3525 1470 3530 1500
rect 3560 1470 3565 1500
rect 3525 1465 3565 1470
rect 3645 1500 3685 1505
rect 3645 1470 3650 1500
rect 3680 1470 3685 1500
rect 3645 1465 3685 1470
rect 3765 1500 3805 1505
rect 3765 1470 3770 1500
rect 3800 1470 3805 1500
rect 3925 1490 3945 2015
rect 4065 2020 4090 2045
rect 4120 2020 4125 2050
rect 4065 2015 4125 2020
rect 4445 2050 4485 2055
rect 4445 2020 4450 2050
rect 4480 2020 4485 2050
rect 4445 2015 4485 2020
rect 4805 2050 4845 2055
rect 4805 2020 4810 2050
rect 4840 2020 4845 2050
rect 4805 2015 4845 2020
rect 5165 2050 5205 2055
rect 5165 2020 5170 2050
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 3765 1465 3805 1470
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 3995 1190 4015 1620
rect 4065 1490 4085 2015
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1850 4365 1880
rect 4325 1845 4365 1850
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1880 4725 1885
rect 4685 1850 4690 1880
rect 4720 1850 4725 1880
rect 4685 1845 4725 1850
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1880 5085 1885
rect 5045 1850 5050 1880
rect 5080 1850 5085 1880
rect 5045 1845 5085 1850
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 4125 1825 4145 1845
rect 4215 1825 4235 1845
rect 4455 1825 4475 1845
rect 4575 1825 4595 1845
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1790 4155 1820
rect 4115 1785 4155 1790
rect 4205 1820 4245 1825
rect 4205 1790 4210 1820
rect 4240 1790 4245 1820
rect 4205 1785 4245 1790
rect 4445 1820 4485 1825
rect 4445 1790 4450 1820
rect 4480 1790 4485 1820
rect 4445 1785 4485 1790
rect 4565 1820 4605 1825
rect 4565 1790 4570 1820
rect 4600 1790 4605 1820
rect 4565 1785 4605 1790
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1730 4245 1760
rect 4205 1725 4245 1730
rect 4445 1760 4485 1765
rect 4445 1730 4450 1760
rect 4480 1730 4485 1760
rect 4445 1725 4485 1730
rect 4575 1720 4595 1785
rect 4695 1765 4715 1845
rect 4815 1825 4835 1845
rect 4935 1825 4955 1845
rect 5145 1825 5165 1845
rect 4805 1820 4845 1825
rect 4805 1790 4810 1820
rect 4840 1790 4845 1820
rect 4805 1785 4845 1790
rect 4925 1820 4965 1825
rect 4925 1790 4930 1820
rect 4960 1790 4965 1820
rect 4925 1785 4965 1790
rect 5135 1820 5175 1825
rect 5135 1790 5140 1820
rect 5170 1790 5175 1820
rect 5135 1785 5175 1790
rect 5280 1765 5300 2255
rect 5325 2150 5345 3105
rect 5315 2145 5355 2150
rect 5315 2115 5320 2145
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 5370 1825 5390 3300
rect 5410 3285 5450 3290
rect 5410 3255 5415 3285
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 5360 1820 5400 1825
rect 5360 1790 5365 1820
rect 5395 1790 5400 1820
rect 5360 1785 5400 1790
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1730 4785 1760
rect 4745 1725 4785 1730
rect 5270 1760 5310 1765
rect 5270 1730 5275 1760
rect 5305 1730 5310 1760
rect 5270 1725 5310 1730
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1685 4365 1715
rect 4325 1680 4365 1685
rect 4565 1715 4605 1720
rect 4565 1685 4570 1715
rect 4600 1685 4605 1715
rect 4565 1680 4605 1685
rect 4805 1715 4845 1720
rect 4805 1685 4810 1715
rect 4840 1685 4845 1715
rect 4805 1680 4845 1685
rect 5420 1600 5440 3250
rect 11060 3160 11080 4280
rect 11340 4265 11360 4285
rect 11750 4280 11790 4285
rect 12140 4315 12180 4320
rect 12140 4285 12145 4315
rect 12175 4285 12180 4315
rect 12140 4280 12180 4285
rect 12203 4310 12237 4320
rect 12203 4290 12211 4310
rect 12229 4290 12237 4310
rect 12203 4280 12237 4290
rect 12260 4315 12300 4320
rect 12260 4285 12265 4315
rect 12295 4285 12300 4315
rect 12260 4280 12300 4285
rect 12380 4315 12420 4320
rect 12380 4285 12385 4315
rect 12415 4285 12420 4315
rect 12380 4280 12420 4285
rect 12500 4315 12540 4320
rect 12500 4285 12505 4315
rect 12535 4285 12540 4315
rect 12500 4280 12540 4285
rect 12210 4265 12230 4280
rect 11105 4260 11145 4265
rect 11105 4230 11110 4260
rect 11140 4230 11145 4260
rect 11105 4225 11145 4230
rect 11330 4260 11370 4265
rect 11330 4230 11335 4260
rect 11365 4230 11370 4260
rect 11330 4225 11370 4230
rect 12200 4260 12240 4265
rect 12200 4230 12205 4260
rect 12235 4230 12240 4260
rect 12200 4225 12240 4230
rect 11050 3155 11090 3160
rect 11050 3125 11055 3155
rect 11085 3125 11090 3155
rect 11050 3120 11090 3125
rect 10265 2965 10305 2970
rect 9899 2935 10040 2940
rect 9899 2905 9905 2935
rect 9935 2905 9955 2935
rect 9985 2905 10005 2935
rect 10035 2905 10040 2935
rect 10265 2935 10270 2965
rect 10300 2935 10305 2965
rect 10265 2930 10305 2935
rect 10375 2965 10415 2970
rect 10375 2935 10380 2965
rect 10410 2935 10415 2965
rect 10375 2930 10415 2935
rect 10485 2965 10525 2970
rect 10485 2935 10490 2965
rect 10520 2935 10525 2965
rect 10485 2930 10525 2935
rect 10595 2965 10635 2970
rect 10595 2935 10600 2965
rect 10630 2935 10635 2965
rect 10595 2930 10635 2935
rect 10653 2960 10687 2970
rect 10653 2940 10661 2960
rect 10679 2940 10687 2960
rect 10653 2930 10687 2940
rect 10705 2965 10745 2970
rect 10705 2935 10710 2965
rect 10740 2935 10745 2965
rect 10705 2930 10745 2935
rect 9899 2900 10040 2905
rect 9960 2885 9980 2900
rect 9950 2880 9990 2885
rect 9950 2850 9955 2880
rect 9985 2850 9990 2880
rect 9950 2845 9990 2850
rect 10385 2830 10405 2930
rect 10660 2885 10680 2930
rect 10650 2880 10690 2885
rect 10650 2850 10655 2880
rect 10685 2850 10690 2880
rect 10650 2845 10690 2850
rect 11000 2880 11040 2885
rect 11000 2850 11005 2880
rect 11035 2850 11040 2880
rect 11000 2845 11040 2850
rect 9745 2825 9785 2830
rect 9745 2795 9750 2825
rect 9780 2795 9785 2825
rect 9745 2790 9785 2795
rect 10375 2825 10415 2830
rect 10375 2795 10380 2825
rect 10410 2795 10415 2825
rect 10375 2790 10415 2795
rect 9755 1710 9775 2790
rect 10210 2705 10250 2710
rect 10210 2675 10215 2705
rect 10245 2675 10250 2705
rect 10210 2670 10250 2675
rect 10320 2705 10360 2710
rect 10320 2675 10325 2705
rect 10355 2675 10360 2705
rect 10320 2670 10360 2675
rect 10430 2705 10470 2710
rect 10430 2675 10435 2705
rect 10465 2675 10470 2705
rect 10430 2670 10470 2675
rect 10540 2705 10580 2710
rect 10540 2675 10545 2705
rect 10575 2675 10580 2705
rect 10540 2670 10580 2675
rect 10650 2705 10690 2710
rect 10650 2675 10655 2705
rect 10685 2675 10690 2705
rect 10650 2670 10690 2675
rect 10760 2705 10800 2710
rect 10760 2675 10765 2705
rect 10795 2675 10800 2705
rect 10760 2670 10800 2675
rect 10020 2435 10060 2440
rect 10020 2405 10025 2435
rect 10055 2405 10060 2435
rect 10020 2400 10060 2405
rect 10265 2435 10305 2440
rect 10265 2405 10270 2435
rect 10300 2405 10305 2435
rect 10265 2400 10305 2405
rect 10375 2435 10415 2440
rect 10375 2405 10380 2435
rect 10410 2405 10415 2435
rect 10375 2400 10415 2405
rect 10485 2435 10525 2440
rect 10485 2405 10490 2435
rect 10520 2405 10525 2435
rect 10485 2400 10525 2405
rect 10595 2435 10635 2440
rect 10595 2405 10600 2435
rect 10630 2405 10635 2435
rect 10595 2400 10635 2405
rect 10705 2435 10745 2440
rect 10705 2405 10710 2435
rect 10740 2405 10745 2435
rect 11010 2425 11030 2845
rect 11115 2480 11135 4225
rect 11360 4205 11400 4210
rect 11360 4175 11365 4205
rect 11395 4175 11400 4205
rect 11360 4170 11400 4175
rect 11470 4205 11510 4210
rect 11470 4175 11475 4205
rect 11505 4175 11510 4205
rect 11470 4170 11510 4175
rect 11580 4205 11620 4210
rect 11580 4175 11585 4205
rect 11615 4175 11620 4205
rect 11580 4170 11620 4175
rect 11690 4205 11730 4210
rect 11690 4175 11695 4205
rect 11725 4175 11730 4205
rect 11690 4170 11730 4175
rect 11800 4205 11840 4210
rect 11800 4175 11805 4205
rect 11835 4175 11840 4205
rect 11800 4170 11840 4175
rect 11910 4205 11950 4210
rect 11910 4175 11915 4205
rect 11945 4175 11950 4205
rect 11910 4170 11950 4175
rect 12020 4205 12060 4210
rect 12020 4175 12025 4205
rect 12055 4175 12060 4205
rect 12020 4170 12060 4175
rect 12130 4205 12170 4210
rect 12130 4175 12135 4205
rect 12165 4175 12170 4205
rect 12130 4170 12170 4175
rect 12240 4205 12280 4210
rect 12240 4175 12245 4205
rect 12275 4175 12280 4205
rect 12240 4170 12280 4175
rect 12350 4205 12390 4210
rect 12350 4175 12355 4205
rect 12385 4175 12390 4205
rect 12350 4170 12390 4175
rect 11305 4085 11345 4090
rect 11305 4055 11310 4085
rect 11340 4055 11345 4085
rect 11305 4050 11345 4055
rect 11362 4080 11398 4090
rect 11362 4060 11370 4080
rect 11390 4060 11398 4080
rect 11362 4050 11398 4060
rect 11415 4080 11455 4090
rect 11415 4060 11425 4080
rect 11445 4060 11455 4080
rect 11415 4050 11455 4060
rect 11525 4085 11565 4090
rect 11525 4055 11530 4085
rect 11560 4055 11565 4085
rect 11525 4050 11565 4055
rect 11635 4080 11675 4090
rect 11635 4060 11645 4080
rect 11665 4060 11675 4080
rect 11635 4050 11675 4060
rect 11745 4085 11785 4090
rect 11745 4055 11750 4085
rect 11780 4055 11785 4085
rect 11745 4050 11785 4055
rect 11855 4080 11895 4090
rect 11855 4060 11865 4080
rect 11885 4060 11895 4080
rect 11855 4050 11895 4060
rect 11965 4085 12005 4090
rect 11965 4055 11970 4085
rect 12000 4055 12005 4085
rect 11965 4050 12005 4055
rect 12075 4080 12115 4090
rect 12075 4060 12085 4080
rect 12105 4060 12115 4080
rect 12075 4050 12115 4060
rect 12185 4085 12225 4090
rect 12185 4055 12190 4085
rect 12220 4055 12225 4085
rect 12185 4050 12225 4055
rect 12295 4080 12335 4090
rect 12295 4060 12305 4080
rect 12325 4060 12335 4080
rect 12295 4050 12335 4060
rect 12405 4085 12445 4090
rect 12405 4055 12410 4085
rect 12440 4055 12445 4085
rect 12405 4050 12445 4055
rect 11310 3960 11350 3965
rect 11310 3930 11315 3960
rect 11345 3930 11350 3960
rect 11310 3925 11350 3930
rect 11370 3905 11390 4050
rect 11425 4030 11445 4050
rect 11645 4030 11665 4050
rect 11865 4030 11885 4050
rect 12085 4030 12105 4050
rect 12305 4030 12325 4050
rect 11415 4025 11455 4030
rect 11415 3995 11420 4025
rect 11450 3995 11455 4025
rect 11415 3990 11455 3995
rect 11635 4025 11675 4030
rect 11635 3995 11640 4025
rect 11670 3995 11675 4025
rect 11635 3990 11675 3995
rect 11855 4025 11895 4030
rect 11855 3995 11860 4025
rect 11890 3995 11895 4025
rect 11855 3990 11895 3995
rect 12075 4025 12115 4030
rect 12075 3995 12080 4025
rect 12110 3995 12115 4025
rect 12075 3990 12115 3995
rect 12295 4025 12335 4030
rect 12295 3995 12300 4025
rect 12330 3995 12335 4025
rect 12295 3990 12335 3995
rect 11425 3965 11445 3990
rect 12415 3965 12435 4050
rect 11415 3960 11455 3965
rect 11415 3930 11420 3960
rect 11450 3930 11455 3960
rect 11415 3925 11455 3930
rect 11525 3960 11565 3965
rect 11525 3930 11530 3960
rect 11560 3930 11565 3960
rect 11525 3925 11565 3930
rect 11635 3960 11675 3965
rect 11635 3930 11640 3960
rect 11670 3930 11675 3960
rect 11635 3925 11675 3930
rect 11745 3960 11785 3965
rect 11745 3930 11750 3960
rect 11780 3930 11785 3960
rect 11745 3925 11785 3930
rect 12050 3960 12090 3965
rect 12050 3930 12055 3960
rect 12085 3930 12090 3960
rect 12050 3925 12090 3930
rect 12155 3960 12195 3965
rect 12155 3930 12160 3960
rect 12190 3930 12195 3960
rect 12155 3925 12195 3930
rect 12265 3960 12305 3965
rect 12265 3930 12270 3960
rect 12300 3930 12305 3960
rect 12265 3925 12305 3930
rect 12375 3960 12435 3965
rect 12375 3930 12380 3960
rect 12410 3930 12435 3960
rect 12375 3925 12435 3930
rect 12485 3960 12525 3965
rect 12485 3930 12490 3960
rect 12520 3930 12525 3960
rect 12485 3925 12525 3930
rect 11271 3900 11303 3905
rect 11271 3870 11274 3900
rect 11300 3870 11303 3900
rect 11271 3865 11303 3870
rect 11360 3895 11400 3905
rect 11360 3875 11370 3895
rect 11390 3875 11400 3895
rect 11360 3865 11400 3875
rect 11470 3900 11510 3905
rect 11470 3870 11475 3900
rect 11505 3870 11510 3900
rect 11470 3865 11510 3870
rect 11690 3900 11730 3905
rect 11690 3870 11695 3900
rect 11725 3870 11730 3900
rect 11690 3865 11730 3870
rect 11800 3895 11840 3905
rect 11800 3875 11810 3895
rect 11830 3875 11840 3895
rect 11800 3865 11840 3875
rect 12011 3900 12043 3905
rect 12011 3870 12014 3900
rect 12040 3870 12043 3900
rect 12011 3865 12043 3870
rect 12210 3900 12250 3905
rect 12210 3870 12215 3900
rect 12245 3870 12250 3900
rect 12210 3865 12250 3870
rect 12430 3900 12470 3905
rect 12430 3870 12435 3900
rect 12465 3870 12470 3900
rect 12430 3865 12470 3870
rect 12760 3900 12800 3905
rect 12760 3870 12765 3900
rect 12795 3870 12800 3900
rect 12760 3865 12800 3870
rect 11402 3780 11434 3785
rect 11402 3750 11405 3780
rect 11431 3750 11434 3780
rect 11402 3745 11434 3750
rect 11622 3780 11654 3785
rect 11622 3750 11625 3780
rect 11651 3750 11654 3780
rect 11622 3745 11654 3750
rect 11766 3780 11798 3785
rect 11766 3750 11769 3780
rect 11795 3750 11798 3780
rect 11766 3745 11798 3750
rect 12142 3780 12174 3785
rect 12142 3750 12145 3780
rect 12171 3750 12174 3780
rect 12142 3745 12174 3750
rect 12362 3780 12394 3785
rect 12362 3750 12365 3780
rect 12391 3750 12394 3780
rect 12362 3745 12394 3750
rect 12506 3780 12538 3785
rect 12506 3750 12509 3780
rect 12535 3750 12538 3780
rect 12506 3745 12538 3750
rect 11990 3730 12030 3735
rect 11250 3720 11290 3725
rect 11250 3690 11255 3720
rect 11285 3690 11290 3720
rect 11250 3685 11290 3690
rect 11355 3720 11395 3725
rect 11355 3690 11360 3720
rect 11390 3690 11395 3720
rect 11355 3685 11395 3690
rect 11470 3720 11510 3725
rect 11470 3690 11475 3720
rect 11505 3690 11510 3720
rect 11470 3685 11510 3690
rect 11575 3720 11615 3725
rect 11575 3690 11580 3720
rect 11610 3690 11615 3720
rect 11575 3685 11615 3690
rect 11690 3720 11730 3725
rect 11690 3690 11695 3720
rect 11725 3690 11730 3720
rect 11690 3685 11730 3690
rect 11805 3720 11845 3725
rect 11805 3690 11810 3720
rect 11840 3690 11845 3720
rect 11990 3700 11995 3730
rect 12025 3700 12030 3730
rect 11990 3695 12030 3700
rect 12210 3730 12250 3735
rect 12210 3700 12215 3730
rect 12245 3700 12250 3730
rect 12210 3695 12250 3700
rect 12430 3730 12470 3735
rect 12430 3700 12435 3730
rect 12465 3700 12470 3730
rect 12430 3695 12470 3700
rect 11805 3685 11845 3690
rect 12095 3685 12135 3690
rect 12095 3655 12100 3685
rect 12130 3655 12135 3685
rect 12095 3650 12135 3655
rect 12315 3685 12355 3690
rect 12315 3655 12320 3685
rect 12350 3655 12355 3685
rect 12315 3650 12355 3655
rect 12545 3685 12585 3690
rect 12545 3655 12550 3685
rect 12580 3655 12585 3685
rect 12545 3650 12585 3655
rect 11340 3625 11380 3630
rect 11340 3595 11345 3625
rect 11375 3595 11380 3625
rect 11340 3590 11380 3595
rect 11460 3625 11500 3630
rect 11460 3595 11465 3625
rect 11495 3595 11500 3625
rect 11460 3590 11500 3595
rect 11580 3625 11620 3630
rect 11580 3595 11585 3625
rect 11615 3595 11620 3625
rect 11580 3590 11620 3595
rect 11700 3625 11740 3630
rect 11700 3595 11705 3625
rect 11735 3595 11740 3625
rect 11700 3590 11740 3595
rect 11820 3625 11860 3630
rect 11820 3595 11825 3625
rect 11855 3595 11860 3625
rect 11820 3590 11860 3595
rect 11940 3625 11980 3630
rect 11940 3595 11945 3625
rect 11975 3595 11980 3625
rect 11940 3590 11980 3595
rect 12060 3625 12100 3630
rect 12060 3595 12065 3625
rect 12095 3595 12100 3625
rect 12060 3590 12100 3595
rect 12180 3625 12220 3630
rect 12180 3595 12185 3625
rect 12215 3595 12220 3625
rect 12180 3590 12220 3595
rect 12300 3625 12340 3630
rect 12300 3595 12305 3625
rect 12335 3595 12340 3625
rect 12300 3590 12340 3595
rect 12420 3625 12460 3630
rect 12420 3595 12425 3625
rect 12455 3595 12460 3625
rect 12420 3590 12460 3595
rect 11280 3150 11320 3160
rect 11280 3130 11290 3150
rect 11310 3130 11320 3150
rect 11280 3120 11320 3130
rect 11400 3150 11440 3160
rect 11400 3130 11410 3150
rect 11430 3130 11440 3150
rect 11400 3120 11440 3130
rect 11520 3150 11560 3160
rect 11520 3130 11530 3150
rect 11550 3130 11560 3150
rect 11520 3120 11560 3130
rect 11640 3150 11680 3160
rect 11640 3130 11650 3150
rect 11670 3130 11680 3150
rect 11640 3120 11680 3130
rect 11760 3150 11800 3160
rect 11760 3130 11770 3150
rect 11790 3130 11800 3150
rect 11760 3120 11800 3130
rect 11823 3155 11857 3160
rect 11823 3125 11826 3155
rect 11854 3125 11857 3155
rect 11823 3120 11857 3125
rect 11880 3150 11920 3160
rect 11880 3130 11890 3150
rect 11910 3130 11920 3150
rect 11880 3120 11920 3130
rect 12000 3150 12040 3160
rect 12000 3130 12010 3150
rect 12030 3130 12040 3150
rect 12000 3120 12040 3130
rect 12120 3150 12160 3160
rect 12120 3130 12130 3150
rect 12150 3130 12160 3150
rect 12120 3120 12160 3130
rect 12240 3150 12280 3160
rect 12240 3130 12250 3150
rect 12270 3130 12280 3150
rect 12240 3120 12280 3130
rect 12360 3150 12400 3160
rect 12360 3130 12370 3150
rect 12390 3130 12400 3150
rect 12360 3120 12400 3130
rect 12480 3150 12520 3160
rect 12480 3130 12490 3150
rect 12510 3130 12520 3150
rect 12480 3120 12520 3130
rect 11290 3105 11310 3120
rect 11280 3100 11320 3105
rect 11280 3070 11285 3100
rect 11315 3070 11320 3100
rect 11280 3065 11320 3070
rect 11410 3060 11430 3120
rect 11530 3105 11550 3120
rect 11520 3100 11560 3105
rect 11520 3070 11525 3100
rect 11555 3070 11560 3100
rect 11520 3065 11560 3070
rect 11650 3060 11670 3120
rect 11770 3105 11790 3120
rect 11760 3100 11800 3105
rect 11760 3070 11765 3100
rect 11795 3070 11800 3100
rect 11760 3065 11800 3070
rect 11890 3060 11910 3120
rect 12010 3105 12030 3120
rect 12000 3100 12040 3105
rect 12000 3070 12005 3100
rect 12035 3070 12040 3100
rect 12000 3065 12040 3070
rect 12130 3060 12150 3120
rect 12250 3105 12270 3120
rect 12240 3100 12280 3105
rect 12240 3070 12245 3100
rect 12275 3070 12280 3100
rect 12240 3065 12280 3070
rect 12370 3060 12390 3120
rect 12490 3105 12510 3120
rect 12480 3100 12520 3105
rect 12480 3070 12485 3100
rect 12515 3070 12520 3100
rect 12480 3065 12520 3070
rect 11400 3055 11440 3060
rect 11400 3025 11405 3055
rect 11435 3025 11440 3055
rect 11400 3020 11440 3025
rect 11640 3055 11680 3060
rect 11640 3025 11645 3055
rect 11675 3025 11680 3055
rect 11640 3020 11680 3025
rect 11880 3055 11920 3060
rect 11880 3025 11885 3055
rect 11915 3025 11920 3055
rect 11880 3020 11920 3025
rect 12120 3055 12160 3060
rect 12120 3025 12125 3055
rect 12155 3025 12160 3055
rect 12120 3020 12160 3025
rect 12360 3055 12400 3060
rect 12360 3025 12365 3055
rect 12395 3025 12400 3055
rect 12360 3020 12400 3025
rect 11410 3005 11430 3020
rect 11340 3000 11380 3005
rect 11340 2970 11345 3000
rect 11375 2970 11380 3000
rect 11340 2965 11380 2970
rect 11400 3000 11440 3005
rect 11400 2970 11405 3000
rect 11435 2970 11440 3000
rect 11400 2965 11440 2970
rect 11580 3000 11620 3005
rect 11580 2970 11585 3000
rect 11615 2970 11620 3000
rect 11580 2965 11620 2970
rect 11820 3000 11860 3005
rect 11820 2970 11825 3000
rect 11855 2970 11860 3000
rect 11820 2965 11860 2970
rect 12060 3000 12100 3005
rect 12060 2970 12065 3000
rect 12095 2970 12100 3000
rect 12060 2965 12100 2970
rect 12300 3000 12340 3005
rect 12300 2970 12305 3000
rect 12335 2970 12340 3000
rect 12300 2965 12340 2970
rect 11350 2950 11370 2965
rect 11590 2950 11610 2965
rect 11830 2950 11850 2965
rect 12070 2950 12090 2965
rect 12310 2950 12330 2965
rect 12490 2950 12510 3065
rect 11340 2940 11380 2950
rect 11340 2920 11350 2940
rect 11370 2920 11380 2940
rect 11340 2910 11380 2920
rect 11460 2945 11500 2950
rect 11460 2915 11465 2945
rect 11495 2915 11500 2945
rect 11460 2910 11500 2915
rect 11580 2940 11620 2950
rect 11580 2920 11590 2940
rect 11610 2920 11620 2940
rect 11580 2910 11620 2920
rect 11700 2945 11740 2950
rect 11700 2915 11705 2945
rect 11735 2915 11740 2945
rect 11700 2910 11740 2915
rect 11820 2940 11860 2950
rect 11820 2920 11830 2940
rect 11850 2920 11860 2940
rect 11820 2910 11860 2920
rect 11940 2945 11980 2950
rect 11940 2915 11945 2945
rect 11975 2915 11980 2945
rect 11940 2910 11980 2915
rect 12060 2940 12100 2950
rect 12060 2920 12070 2940
rect 12090 2920 12100 2940
rect 12060 2910 12100 2920
rect 12180 2945 12220 2950
rect 12180 2915 12185 2945
rect 12215 2915 12220 2945
rect 12180 2910 12220 2915
rect 12300 2940 12340 2950
rect 12300 2920 12310 2940
rect 12330 2920 12340 2940
rect 12300 2910 12340 2920
rect 12420 2945 12460 2950
rect 12420 2915 12425 2945
rect 12455 2915 12460 2945
rect 12420 2910 12460 2915
rect 12480 2945 12520 2950
rect 12480 2915 12485 2945
rect 12515 2915 12520 2945
rect 12480 2910 12520 2915
rect 12690 2880 12730 2885
rect 12690 2850 12695 2880
rect 12725 2850 12730 2880
rect 12690 2845 12730 2850
rect 11105 2475 11145 2480
rect 11105 2445 11110 2475
rect 11140 2445 11145 2475
rect 11105 2440 11145 2445
rect 11280 2470 11320 2480
rect 11280 2450 11290 2470
rect 11310 2450 11320 2470
rect 11280 2440 11320 2450
rect 11400 2470 11440 2480
rect 11400 2450 11410 2470
rect 11430 2450 11440 2470
rect 11400 2440 11440 2450
rect 11520 2470 11560 2480
rect 11520 2450 11530 2470
rect 11550 2450 11560 2470
rect 11520 2440 11560 2450
rect 11640 2470 11680 2480
rect 11640 2450 11650 2470
rect 11670 2450 11680 2470
rect 11640 2440 11680 2450
rect 11760 2470 11800 2480
rect 11760 2450 11770 2470
rect 11790 2450 11800 2470
rect 11760 2440 11800 2450
rect 11823 2475 11857 2480
rect 11823 2445 11826 2475
rect 11854 2445 11857 2475
rect 11823 2440 11857 2445
rect 11880 2470 11920 2480
rect 11880 2450 11890 2470
rect 11910 2450 11920 2470
rect 11880 2440 11920 2450
rect 12000 2470 12040 2480
rect 12000 2450 12010 2470
rect 12030 2450 12040 2470
rect 12000 2440 12040 2450
rect 12120 2470 12160 2480
rect 12120 2450 12130 2470
rect 12150 2450 12160 2470
rect 12120 2440 12160 2450
rect 12240 2470 12280 2480
rect 12240 2450 12250 2470
rect 12270 2450 12280 2470
rect 12240 2440 12280 2450
rect 12360 2470 12400 2480
rect 12360 2450 12370 2470
rect 12390 2450 12400 2470
rect 12360 2440 12400 2450
rect 12480 2470 12520 2480
rect 12480 2450 12490 2470
rect 12510 2450 12520 2470
rect 12480 2440 12520 2450
rect 11290 2425 11310 2440
rect 10705 2400 10745 2405
rect 11000 2420 11040 2425
rect 9790 2005 9825 2011
rect 9790 1965 9825 1970
rect 9850 2005 9885 2010
rect 9850 1965 9885 1970
rect 9910 2005 9945 2011
rect 9910 1965 9945 1970
rect 9970 2005 10005 2010
rect 10030 2005 10050 2400
rect 10765 2390 10805 2395
rect 10765 2360 10770 2390
rect 10800 2360 10805 2390
rect 11000 2390 11005 2420
rect 11035 2390 11040 2420
rect 11000 2385 11040 2390
rect 11280 2420 11320 2425
rect 11280 2390 11285 2420
rect 11315 2390 11320 2420
rect 11280 2385 11320 2390
rect 11410 2380 11430 2440
rect 11530 2425 11550 2440
rect 11520 2420 11560 2425
rect 11520 2390 11525 2420
rect 11555 2390 11560 2420
rect 11520 2385 11560 2390
rect 11650 2380 11670 2440
rect 11770 2425 11790 2440
rect 11760 2420 11800 2425
rect 11760 2390 11765 2420
rect 11795 2390 11800 2420
rect 11760 2385 11800 2390
rect 10765 2355 10805 2360
rect 11400 2375 11440 2380
rect 11400 2345 11405 2375
rect 11435 2345 11440 2375
rect 11400 2340 11440 2345
rect 11640 2375 11680 2380
rect 11640 2345 11645 2375
rect 11675 2345 11680 2375
rect 11640 2340 11680 2345
rect 11000 2325 11040 2330
rect 10065 2315 10105 2320
rect 10065 2285 10070 2315
rect 10100 2285 10105 2315
rect 10065 2280 10105 2285
rect 10265 2315 10305 2320
rect 10265 2285 10270 2315
rect 10300 2285 10305 2315
rect 10265 2280 10305 2285
rect 10375 2315 10415 2320
rect 10375 2285 10380 2315
rect 10410 2285 10415 2315
rect 10375 2280 10415 2285
rect 10485 2315 10525 2320
rect 10485 2285 10490 2315
rect 10520 2285 10525 2315
rect 10485 2280 10525 2285
rect 10595 2315 10635 2320
rect 10595 2285 10600 2315
rect 10630 2285 10635 2315
rect 10595 2280 10635 2285
rect 10705 2315 10745 2320
rect 10705 2285 10710 2315
rect 10740 2285 10745 2315
rect 11000 2295 11005 2325
rect 11035 2295 11040 2325
rect 11000 2290 11040 2295
rect 10705 2280 10745 2285
rect 9970 1965 10005 1970
rect 10020 2000 10060 2005
rect 10020 1970 10025 2000
rect 10055 1970 10060 2000
rect 10020 1965 10060 1970
rect 9800 1900 9820 1965
rect 9920 1950 9940 1965
rect 10075 1950 10095 2280
rect 10950 2180 10990 2185
rect 10950 2150 10955 2180
rect 10985 2150 10990 2180
rect 10950 2145 10990 2150
rect 9910 1945 9950 1950
rect 9910 1915 9915 1945
rect 9945 1915 9950 1945
rect 9910 1910 9950 1915
rect 10065 1945 10105 1950
rect 10065 1915 10070 1945
rect 10100 1915 10105 1945
rect 10065 1910 10105 1915
rect 10210 1945 10250 1950
rect 10210 1915 10215 1945
rect 10245 1915 10250 1945
rect 10210 1910 10250 1915
rect 10320 1945 10360 1950
rect 10320 1915 10325 1945
rect 10355 1915 10360 1945
rect 10320 1910 10360 1915
rect 10430 1945 10470 1950
rect 10430 1915 10435 1945
rect 10465 1915 10470 1945
rect 10430 1910 10470 1915
rect 10540 1945 10580 1950
rect 10540 1915 10545 1945
rect 10575 1915 10580 1945
rect 10540 1910 10580 1915
rect 10650 1945 10690 1950
rect 10650 1915 10655 1945
rect 10685 1915 10690 1945
rect 10650 1910 10690 1915
rect 10760 1945 10800 1950
rect 10760 1915 10765 1945
rect 10795 1915 10800 1945
rect 10760 1910 10800 1915
rect 9790 1895 9830 1900
rect 9790 1865 9795 1895
rect 9825 1865 9830 1895
rect 9790 1860 9830 1865
rect 9965 1760 10005 1765
rect 9965 1730 9970 1760
rect 10000 1730 10005 1760
rect 9965 1725 10005 1730
rect 10555 1760 10595 1765
rect 10555 1730 10560 1760
rect 10590 1730 10595 1760
rect 10555 1725 10595 1730
rect 9745 1705 9785 1710
rect 9745 1675 9750 1705
rect 9780 1675 9785 1705
rect 9745 1670 9785 1675
rect 9975 1650 9995 1725
rect 10565 1710 10585 1725
rect 10030 1705 10070 1710
rect 10030 1675 10035 1705
rect 10065 1675 10070 1705
rect 10030 1670 10070 1675
rect 10255 1705 10295 1710
rect 10255 1675 10260 1705
rect 10290 1675 10295 1705
rect 10255 1670 10295 1675
rect 10455 1705 10495 1710
rect 10455 1675 10460 1705
rect 10490 1675 10495 1705
rect 10455 1670 10495 1675
rect 10558 1700 10592 1710
rect 10558 1680 10566 1700
rect 10584 1680 10592 1700
rect 10558 1670 10592 1680
rect 10655 1705 10695 1710
rect 10655 1675 10660 1705
rect 10690 1675 10695 1705
rect 10655 1670 10695 1675
rect 10835 1705 10875 1710
rect 10835 1675 10840 1705
rect 10870 1675 10875 1705
rect 10835 1670 10875 1675
rect 10040 1650 10060 1670
rect 9970 1645 10005 1650
rect 9970 1605 10005 1610
rect 10030 1645 10065 1650
rect 10030 1605 10065 1610
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1565 4845 1595
rect 4805 1560 4845 1565
rect 5410 1595 5450 1600
rect 5410 1565 5415 1595
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1515 4305 1545
rect 4265 1510 4305 1515
rect 4385 1545 4425 1550
rect 4385 1515 4390 1545
rect 4420 1515 4425 1545
rect 4385 1510 4425 1515
rect 4505 1545 4545 1550
rect 4505 1515 4510 1545
rect 4540 1515 4545 1545
rect 4505 1510 4545 1515
rect 4625 1545 4665 1550
rect 4625 1515 4630 1545
rect 4660 1515 4665 1545
rect 4625 1510 4665 1515
rect 4745 1545 4785 1550
rect 4745 1515 4750 1545
rect 4780 1515 4785 1545
rect 4745 1510 4785 1515
rect 5135 1545 5175 1550
rect 5135 1515 5140 1545
rect 5170 1515 5175 1545
rect 5135 1510 5175 1515
rect 4205 1500 4245 1505
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1470 4210 1500
rect 4240 1470 4245 1500
rect 4205 1465 4245 1470
rect 4325 1500 4365 1505
rect 4325 1470 4330 1500
rect 4360 1470 4365 1500
rect 4325 1465 4365 1470
rect 4445 1500 4485 1505
rect 4445 1470 4450 1500
rect 4480 1470 4485 1500
rect 4445 1465 4485 1470
rect 4685 1500 4725 1505
rect 4685 1470 4690 1500
rect 4720 1470 4725 1500
rect 4685 1465 4725 1470
rect 4805 1500 4845 1505
rect 4805 1470 4810 1500
rect 4840 1470 4845 1500
rect 4805 1465 4845 1470
rect 4925 1500 4965 1505
rect 4925 1470 4930 1500
rect 4960 1470 4965 1500
rect 4925 1465 4965 1470
rect 5045 1500 5085 1505
rect 5045 1470 5050 1500
rect 5080 1470 5085 1500
rect 5145 1490 5165 1510
rect 5045 1465 5085 1470
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 10845 1395 10865 1670
rect 10835 1390 10875 1395
rect 10835 1360 10840 1390
rect 10870 1360 10875 1390
rect 10835 1355 10875 1360
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1155 3415 1185
rect 3375 1150 3415 1155
rect 3985 1185 4025 1190
rect 3985 1155 3990 1185
rect 4020 1155 4025 1185
rect 3985 1150 4025 1155
rect 4595 1185 4635 1190
rect 4595 1155 4600 1185
rect 4630 1155 4635 1185
rect 4595 1150 4635 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1095 2985 1125
rect 2945 1090 2985 1095
rect 3025 1125 3065 1130
rect 3025 1095 3030 1125
rect 3060 1095 3065 1125
rect 3025 1090 3065 1095
rect 3105 1125 3145 1130
rect 3105 1095 3110 1125
rect 3140 1095 3145 1125
rect 3105 1090 3145 1095
rect 3185 1125 3225 1130
rect 3185 1095 3190 1125
rect 3220 1095 3225 1125
rect 3185 1090 3225 1095
rect 3265 1125 3305 1130
rect 3265 1095 3270 1125
rect 3300 1095 3305 1125
rect 3265 1090 3305 1095
rect 3345 1125 3385 1130
rect 3345 1095 3350 1125
rect 3380 1095 3385 1125
rect 3345 1090 3385 1095
rect 3425 1125 3465 1130
rect 3425 1095 3430 1125
rect 3460 1095 3465 1125
rect 3425 1090 3465 1095
rect 3505 1125 3545 1130
rect 3505 1095 3510 1125
rect 3540 1095 3545 1125
rect 3505 1090 3545 1095
rect 3585 1125 3625 1130
rect 3585 1095 3590 1125
rect 3620 1095 3625 1125
rect 3585 1090 3625 1095
rect 3665 1125 3705 1130
rect 3665 1095 3670 1125
rect 3700 1095 3705 1125
rect 3665 1090 3705 1095
rect 3745 1125 3785 1130
rect 3745 1095 3750 1125
rect 3780 1095 3785 1125
rect 3745 1090 3785 1095
rect 3825 1125 3865 1130
rect 3825 1095 3830 1125
rect 3860 1095 3865 1125
rect 3825 1090 3865 1095
rect 3905 1125 3945 1130
rect 3905 1095 3910 1125
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1095 4025 1125
rect 3985 1090 4025 1095
rect 4065 1125 4105 1130
rect 4065 1095 4070 1125
rect 4100 1095 4105 1125
rect 4065 1090 4105 1095
rect 4145 1125 4185 1130
rect 4145 1095 4150 1125
rect 4180 1095 4185 1125
rect 4145 1090 4185 1095
rect 4225 1125 4265 1130
rect 4225 1095 4230 1125
rect 4260 1095 4265 1125
rect 4225 1090 4265 1095
rect 4305 1125 4345 1130
rect 4305 1095 4310 1125
rect 4340 1095 4345 1125
rect 4305 1090 4345 1095
rect 4385 1125 4425 1130
rect 4385 1095 4390 1125
rect 4420 1095 4425 1125
rect 4385 1090 4425 1095
rect 4465 1125 4505 1130
rect 4465 1095 4470 1125
rect 4500 1095 4505 1125
rect 4465 1090 4505 1095
rect 4545 1125 4585 1130
rect 4545 1095 4550 1125
rect 4580 1095 4585 1125
rect 4545 1090 4585 1095
rect 4625 1125 4665 1130
rect 4625 1095 4630 1125
rect 4660 1095 4665 1125
rect 4625 1090 4665 1095
rect 4705 1125 4745 1130
rect 4705 1095 4710 1125
rect 4740 1095 4745 1125
rect 4705 1090 4745 1095
rect 4785 1125 4825 1130
rect 4785 1095 4790 1125
rect 4820 1095 4825 1125
rect 4785 1090 4825 1095
rect 4865 1125 4905 1130
rect 4865 1095 4870 1125
rect 4900 1095 4905 1125
rect 4865 1090 4905 1095
rect 4945 1125 4985 1130
rect 4945 1095 4950 1125
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1010 2660 1040
rect 2620 1005 2660 1010
rect 2905 1040 2945 1045
rect 2905 1010 2910 1040
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1010 5150 1040
rect 5110 1005 5150 1010
rect 10355 935 10395 940
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 900 3035 930
rect 2995 895 3035 900
rect 3175 930 3215 935
rect 3175 900 3180 930
rect 3210 900 3215 930
rect 3175 895 3215 900
rect 3355 930 3395 935
rect 3355 900 3360 930
rect 3390 900 3395 930
rect 3355 895 3395 900
rect 3535 930 3575 935
rect 3535 900 3540 930
rect 3570 900 3575 930
rect 3535 895 3575 900
rect 3715 930 3755 935
rect 3715 900 3720 930
rect 3750 900 3755 930
rect 3715 895 3755 900
rect 3895 930 3935 935
rect 3895 900 3900 930
rect 3930 900 3935 930
rect 3895 895 3935 900
rect 4075 930 4115 935
rect 4075 900 4080 930
rect 4110 900 4115 930
rect 4075 895 4115 900
rect 4255 930 4295 935
rect 4255 900 4260 930
rect 4290 900 4295 930
rect 4255 895 4295 900
rect 4435 930 4475 935
rect 4435 900 4440 930
rect 4470 900 4475 930
rect 4435 895 4475 900
rect 4615 930 4655 935
rect 4615 900 4620 930
rect 4650 900 4655 930
rect 4615 895 4655 900
rect 4795 930 4835 935
rect 4795 900 4800 930
rect 4830 900 4835 930
rect 4795 895 4835 900
rect 4975 930 5015 935
rect 4975 900 4980 930
rect 5010 900 5015 930
rect 10355 905 10360 935
rect 10390 905 10395 935
rect 10355 900 10395 905
rect 10555 935 10595 940
rect 10555 905 10560 935
rect 10590 905 10595 935
rect 10555 900 10595 905
rect 4975 895 5015 900
rect 10960 800 10980 2145
rect 11010 1900 11030 2290
rect 11440 2280 11480 2285
rect 11440 2250 11445 2280
rect 11475 2250 11480 2280
rect 11440 2245 11480 2250
rect 11660 2280 11700 2285
rect 11660 2250 11665 2280
rect 11695 2250 11700 2280
rect 11660 2245 11700 2250
rect 11330 2235 11370 2240
rect 11330 2205 11335 2235
rect 11365 2205 11370 2235
rect 11330 2200 11370 2205
rect 11340 2185 11360 2200
rect 11450 2185 11470 2245
rect 11550 2235 11590 2240
rect 11550 2205 11555 2235
rect 11585 2205 11590 2235
rect 11550 2200 11590 2205
rect 11560 2185 11580 2200
rect 11670 2185 11690 2245
rect 11770 2240 11790 2385
rect 11890 2380 11910 2440
rect 12010 2425 12030 2440
rect 12000 2420 12040 2425
rect 12000 2390 12005 2420
rect 12035 2390 12040 2420
rect 12000 2385 12040 2390
rect 12130 2380 12150 2440
rect 12250 2425 12270 2440
rect 12240 2420 12280 2425
rect 12240 2390 12245 2420
rect 12275 2390 12280 2420
rect 12240 2385 12280 2390
rect 12370 2380 12390 2440
rect 12490 2425 12510 2440
rect 12480 2420 12520 2425
rect 12480 2390 12485 2420
rect 12515 2390 12520 2420
rect 12480 2385 12520 2390
rect 12700 2380 12720 2845
rect 11880 2375 11920 2380
rect 11880 2345 11885 2375
rect 11915 2345 11920 2375
rect 11880 2340 11920 2345
rect 12120 2375 12160 2380
rect 12120 2345 12125 2375
rect 12155 2345 12160 2375
rect 12120 2340 12160 2345
rect 12360 2375 12400 2380
rect 12360 2345 12365 2375
rect 12395 2345 12400 2375
rect 12360 2340 12400 2345
rect 12690 2375 12730 2380
rect 12690 2345 12695 2375
rect 12725 2345 12730 2375
rect 12690 2340 12730 2345
rect 12120 2285 12140 2340
rect 12770 2330 12790 3865
rect 12860 3730 12900 3735
rect 12860 3700 12865 3730
rect 12895 3700 12900 3730
rect 12860 3695 12900 3700
rect 12805 3685 12845 3690
rect 12805 3655 12810 3685
rect 12840 3655 12845 3685
rect 12805 3650 12845 3655
rect 12760 2325 12800 2330
rect 12760 2295 12765 2325
rect 12795 2295 12800 2325
rect 12760 2290 12800 2295
rect 11880 2280 11920 2285
rect 11880 2250 11885 2280
rect 11915 2250 11920 2280
rect 11880 2245 11920 2250
rect 12100 2280 12140 2285
rect 12100 2250 12105 2280
rect 12135 2250 12140 2280
rect 12100 2245 12140 2250
rect 12320 2280 12360 2285
rect 12320 2250 12325 2280
rect 12355 2250 12360 2280
rect 12320 2245 12360 2250
rect 11770 2235 11810 2240
rect 11770 2205 11775 2235
rect 11805 2205 11810 2235
rect 11770 2200 11810 2205
rect 11780 2185 11800 2200
rect 11890 2185 11910 2245
rect 11990 2235 12030 2240
rect 11990 2205 11995 2235
rect 12025 2205 12030 2235
rect 11990 2200 12030 2205
rect 12000 2185 12020 2200
rect 12110 2185 12130 2245
rect 12210 2235 12250 2240
rect 12210 2205 12215 2235
rect 12245 2205 12250 2235
rect 12210 2200 12250 2205
rect 12220 2185 12240 2200
rect 12330 2185 12350 2245
rect 12430 2235 12470 2240
rect 12430 2205 12435 2235
rect 12465 2205 12470 2235
rect 12430 2200 12470 2205
rect 12440 2185 12460 2200
rect 11330 2175 11370 2185
rect 11330 2155 11340 2175
rect 11360 2155 11370 2175
rect 11330 2145 11370 2155
rect 11440 2175 11480 2185
rect 11440 2155 11450 2175
rect 11470 2155 11480 2175
rect 11440 2145 11480 2155
rect 11550 2175 11590 2185
rect 11550 2155 11560 2175
rect 11580 2155 11590 2175
rect 11550 2145 11590 2155
rect 11660 2175 11700 2185
rect 11660 2155 11670 2175
rect 11690 2155 11700 2175
rect 11660 2145 11700 2155
rect 11770 2175 11810 2185
rect 11770 2155 11780 2175
rect 11800 2155 11810 2175
rect 11770 2145 11810 2155
rect 11828 2180 11862 2185
rect 11828 2150 11831 2180
rect 11859 2150 11862 2180
rect 11828 2145 11862 2150
rect 11880 2175 11920 2185
rect 11880 2155 11890 2175
rect 11910 2155 11920 2175
rect 11880 2145 11920 2155
rect 11990 2175 12030 2185
rect 11990 2155 12000 2175
rect 12020 2155 12030 2175
rect 11990 2145 12030 2155
rect 12100 2175 12140 2185
rect 12100 2155 12110 2175
rect 12130 2155 12140 2175
rect 12100 2145 12140 2155
rect 12210 2175 12250 2185
rect 12210 2155 12220 2175
rect 12240 2155 12250 2175
rect 12210 2145 12250 2155
rect 12320 2175 12360 2185
rect 12320 2155 12330 2175
rect 12350 2155 12360 2175
rect 12320 2145 12360 2155
rect 12430 2175 12470 2185
rect 12430 2155 12440 2175
rect 12460 2155 12470 2175
rect 12430 2145 12470 2155
rect 11385 1960 11425 1965
rect 11385 1930 11390 1960
rect 11420 1930 11425 1960
rect 11385 1925 11425 1930
rect 11495 1955 11535 1965
rect 11495 1935 11505 1955
rect 11525 1935 11535 1955
rect 11495 1925 11535 1935
rect 11605 1960 11645 1965
rect 11605 1930 11610 1960
rect 11640 1930 11645 1960
rect 11605 1925 11645 1930
rect 11715 1955 11755 1965
rect 11715 1935 11725 1955
rect 11745 1935 11755 1955
rect 11715 1925 11755 1935
rect 11825 1960 11865 1965
rect 11825 1930 11830 1960
rect 11860 1930 11865 1960
rect 11825 1925 11865 1930
rect 11935 1955 11975 1965
rect 11935 1935 11945 1955
rect 11965 1935 11975 1955
rect 11935 1925 11975 1935
rect 12045 1960 12085 1965
rect 12045 1930 12050 1960
rect 12080 1930 12085 1960
rect 12045 1925 12085 1930
rect 12155 1955 12195 1965
rect 12155 1935 12165 1955
rect 12185 1935 12195 1955
rect 12155 1925 12195 1935
rect 12245 1960 12305 1965
rect 12245 1930 12270 1960
rect 12300 1930 12305 1960
rect 12245 1925 12305 1930
rect 12375 1955 12415 1965
rect 12375 1935 12385 1955
rect 12405 1935 12415 1955
rect 12375 1925 12415 1935
rect 11505 1910 11525 1925
rect 11725 1910 11745 1925
rect 11945 1910 11965 1925
rect 12165 1910 12185 1925
rect 11495 1905 11555 1910
rect 11000 1895 11040 1900
rect 11000 1865 11005 1895
rect 11035 1865 11040 1895
rect 11495 1875 11500 1905
rect 11530 1875 11555 1905
rect 11495 1870 11555 1875
rect 11715 1905 11755 1910
rect 11715 1875 11720 1905
rect 11750 1875 11755 1905
rect 11715 1870 11755 1875
rect 11935 1905 11975 1910
rect 11935 1875 11940 1905
rect 11970 1875 11975 1905
rect 11935 1870 11975 1875
rect 12155 1905 12195 1910
rect 12155 1875 12160 1905
rect 12190 1875 12195 1905
rect 12155 1870 12195 1875
rect 11000 1860 11040 1865
rect 11190 1850 11230 1855
rect 11190 1820 11195 1850
rect 11225 1820 11230 1850
rect 11190 1815 11230 1820
rect 11410 1850 11450 1855
rect 11410 1820 11415 1850
rect 11445 1820 11450 1850
rect 11410 1815 11450 1820
rect 11200 1780 11220 1815
rect 11420 1780 11440 1815
rect 11190 1770 11230 1780
rect 11085 1760 11125 1765
rect 11085 1730 11090 1760
rect 11120 1730 11125 1760
rect 11190 1750 11200 1770
rect 11220 1750 11230 1770
rect 11410 1770 11450 1780
rect 11190 1740 11230 1750
rect 11305 1760 11345 1765
rect 11085 1725 11125 1730
rect 11305 1730 11310 1760
rect 11340 1730 11345 1760
rect 11410 1750 11420 1770
rect 11440 1750 11450 1770
rect 11535 1765 11555 1870
rect 12245 1855 12265 1925
rect 12385 1910 12405 1925
rect 12375 1905 12415 1910
rect 12375 1875 12380 1905
rect 12410 1875 12415 1905
rect 12770 1900 12790 2290
rect 12375 1870 12415 1875
rect 12760 1895 12800 1900
rect 12760 1865 12765 1895
rect 12795 1865 12800 1895
rect 12760 1860 12800 1865
rect 11640 1850 11680 1855
rect 11640 1820 11645 1850
rect 11675 1820 11680 1850
rect 11640 1815 11680 1820
rect 12230 1850 12270 1855
rect 12230 1820 12235 1850
rect 12265 1820 12270 1850
rect 12230 1815 12270 1820
rect 12450 1850 12490 1855
rect 12450 1820 12455 1850
rect 12485 1820 12490 1850
rect 12450 1815 12490 1820
rect 12680 1850 12720 1855
rect 12680 1820 12685 1850
rect 12715 1820 12720 1850
rect 12680 1815 12720 1820
rect 11650 1780 11670 1815
rect 11820 1805 11860 1810
rect 11640 1770 11680 1780
rect 11820 1775 11825 1805
rect 11855 1775 11860 1805
rect 11820 1770 11860 1775
rect 11940 1805 11980 1810
rect 11940 1775 11945 1805
rect 11975 1775 11980 1805
rect 12240 1780 12260 1815
rect 12460 1780 12480 1815
rect 12690 1780 12710 1815
rect 11940 1770 11980 1775
rect 12230 1770 12270 1780
rect 11410 1740 11450 1750
rect 11525 1760 11565 1765
rect 11305 1725 11345 1730
rect 11525 1730 11530 1760
rect 11560 1730 11565 1760
rect 11640 1750 11650 1770
rect 11670 1750 11680 1770
rect 11640 1740 11680 1750
rect 11525 1725 11565 1730
rect 11830 1720 11850 1770
rect 11950 1720 11970 1770
rect 12125 1760 12165 1765
rect 12125 1730 12130 1760
rect 12160 1730 12165 1760
rect 12230 1750 12240 1770
rect 12260 1750 12270 1770
rect 12450 1770 12490 1780
rect 12230 1740 12270 1750
rect 12345 1760 12385 1765
rect 12125 1725 12165 1730
rect 12345 1730 12350 1760
rect 12380 1730 12385 1760
rect 12450 1750 12460 1770
rect 12480 1750 12490 1770
rect 12680 1770 12720 1780
rect 12450 1740 12490 1750
rect 12565 1760 12605 1765
rect 12345 1725 12385 1730
rect 12565 1730 12570 1760
rect 12600 1730 12605 1760
rect 12680 1750 12690 1770
rect 12710 1750 12720 1770
rect 12680 1740 12720 1750
rect 12565 1725 12605 1730
rect 11237 1715 11269 1720
rect 11237 1685 11240 1715
rect 11266 1685 11269 1715
rect 11237 1680 11269 1685
rect 11457 1715 11489 1720
rect 11457 1685 11460 1715
rect 11486 1685 11489 1715
rect 11457 1680 11489 1685
rect 11601 1715 11633 1720
rect 11601 1685 11604 1715
rect 11630 1685 11633 1715
rect 11601 1680 11633 1685
rect 11820 1710 11850 1720
rect 11820 1690 11825 1710
rect 11845 1690 11850 1710
rect 11820 1680 11850 1690
rect 11867 1715 11899 1720
rect 11867 1685 11870 1715
rect 11896 1685 11899 1715
rect 11867 1680 11899 1685
rect 11950 1710 11980 1720
rect 11950 1690 11955 1710
rect 11975 1690 11980 1710
rect 11950 1680 11980 1690
rect 12277 1715 12309 1720
rect 12277 1685 12280 1715
rect 12306 1685 12309 1715
rect 12277 1680 12309 1685
rect 12497 1715 12529 1720
rect 12497 1685 12500 1715
rect 12526 1685 12529 1715
rect 12497 1680 12529 1685
rect 12641 1715 12673 1720
rect 12641 1685 12644 1715
rect 12670 1685 12673 1715
rect 12641 1680 12673 1685
rect 11106 1495 11138 1500
rect 11106 1465 11109 1495
rect 11135 1465 11138 1495
rect 11106 1460 11138 1465
rect 11305 1495 11345 1500
rect 11305 1465 11310 1495
rect 11340 1465 11345 1495
rect 11305 1460 11345 1465
rect 11525 1495 11565 1500
rect 11525 1465 11530 1495
rect 11560 1465 11565 1495
rect 11525 1460 11565 1465
rect 11825 1490 11855 1500
rect 11825 1470 11830 1490
rect 11850 1470 11855 1490
rect 11825 1460 11855 1470
rect 11875 1490 11905 1500
rect 11875 1470 11880 1490
rect 11900 1470 11905 1490
rect 11875 1460 11905 1470
rect 11922 1495 11954 1500
rect 11922 1465 11925 1495
rect 11951 1465 11954 1495
rect 11922 1460 11954 1465
rect 12146 1495 12178 1500
rect 12146 1465 12149 1495
rect 12175 1465 12178 1495
rect 12146 1460 12178 1465
rect 12345 1495 12385 1500
rect 12345 1465 12350 1495
rect 12380 1465 12385 1495
rect 12345 1460 12385 1465
rect 12565 1495 12605 1500
rect 12565 1465 12570 1495
rect 12600 1465 12605 1495
rect 12565 1460 12605 1465
rect 11145 1435 11185 1440
rect 11145 1405 11150 1435
rect 11180 1405 11185 1435
rect 11145 1400 11185 1405
rect 11250 1435 11290 1440
rect 11250 1405 11255 1435
rect 11285 1405 11290 1435
rect 11250 1400 11290 1405
rect 11360 1435 11400 1440
rect 11360 1405 11365 1435
rect 11395 1405 11400 1435
rect 11360 1400 11400 1405
rect 11470 1435 11510 1440
rect 11470 1405 11475 1435
rect 11505 1405 11510 1435
rect 11470 1400 11510 1405
rect 11580 1435 11620 1440
rect 11580 1405 11585 1435
rect 11615 1405 11620 1435
rect 11580 1400 11620 1405
rect 11830 1350 11850 1460
rect 11005 1345 11045 1350
rect 11005 1315 11010 1345
rect 11040 1315 11045 1345
rect 11005 1310 11045 1315
rect 11810 1345 11850 1350
rect 11810 1315 11815 1345
rect 11845 1315 11850 1345
rect 11810 1310 11850 1315
rect 11015 860 11035 1310
rect 11315 1295 11355 1300
rect 11315 1265 11320 1295
rect 11350 1265 11355 1295
rect 11315 1260 11355 1265
rect 11325 1240 11345 1260
rect 11820 1240 11840 1310
rect 11880 1300 11900 1460
rect 12185 1435 12225 1440
rect 12185 1405 12190 1435
rect 12220 1405 12225 1435
rect 12185 1400 12225 1405
rect 12290 1435 12330 1440
rect 12290 1405 12295 1435
rect 12325 1405 12330 1435
rect 12290 1400 12330 1405
rect 12400 1435 12440 1440
rect 12400 1405 12405 1435
rect 12435 1405 12440 1435
rect 12400 1400 12440 1405
rect 12510 1435 12550 1440
rect 12510 1405 12515 1435
rect 12545 1405 12550 1435
rect 12510 1400 12550 1405
rect 12620 1435 12660 1440
rect 12620 1405 12625 1435
rect 12655 1405 12660 1435
rect 12620 1400 12660 1405
rect 11880 1295 11920 1300
rect 11880 1265 11885 1295
rect 11915 1265 11920 1295
rect 11880 1260 11920 1265
rect 12815 1255 12835 3650
rect 12595 1250 12635 1255
rect 11315 1230 11355 1240
rect 11315 1210 11325 1230
rect 11345 1210 11355 1230
rect 11315 1200 11355 1210
rect 11425 1235 11465 1240
rect 11425 1205 11430 1235
rect 11460 1205 11465 1235
rect 11425 1200 11465 1205
rect 11535 1235 11575 1240
rect 11535 1205 11540 1235
rect 11570 1205 11575 1235
rect 11535 1200 11575 1205
rect 11645 1235 11685 1240
rect 11645 1205 11650 1235
rect 11680 1205 11685 1235
rect 11645 1200 11685 1205
rect 11755 1235 11795 1240
rect 11755 1205 11760 1235
rect 11790 1205 11795 1235
rect 11755 1200 11795 1205
rect 11815 1230 11845 1240
rect 11815 1210 11820 1230
rect 11840 1210 11845 1230
rect 11815 1200 11845 1210
rect 11865 1235 11905 1240
rect 11865 1205 11870 1235
rect 11900 1205 11905 1235
rect 11865 1200 11905 1205
rect 11975 1235 12015 1240
rect 11975 1205 11980 1235
rect 12010 1205 12015 1235
rect 11975 1200 12015 1205
rect 12085 1235 12125 1240
rect 12085 1205 12090 1235
rect 12120 1205 12125 1235
rect 12085 1200 12125 1205
rect 12195 1235 12235 1240
rect 12195 1205 12200 1235
rect 12230 1205 12235 1235
rect 12195 1200 12235 1205
rect 12305 1235 12345 1240
rect 12305 1205 12310 1235
rect 12340 1205 12345 1235
rect 12305 1200 12345 1205
rect 12415 1235 12455 1240
rect 12415 1205 12420 1235
rect 12450 1205 12455 1235
rect 12415 1200 12455 1205
rect 12525 1235 12565 1240
rect 12525 1205 12530 1235
rect 12560 1205 12565 1235
rect 12595 1220 12600 1250
rect 12630 1220 12635 1250
rect 12595 1215 12635 1220
rect 12805 1250 12845 1255
rect 12805 1220 12810 1250
rect 12840 1220 12845 1250
rect 12805 1215 12845 1220
rect 12525 1200 12565 1205
rect 11165 915 11205 920
rect 11165 885 11170 915
rect 11200 885 11205 915
rect 11165 880 11205 885
rect 11260 915 11300 920
rect 11260 885 11265 915
rect 11295 885 11300 915
rect 11260 880 11300 885
rect 11370 915 11410 920
rect 11370 885 11375 915
rect 11405 885 11410 915
rect 11370 880 11410 885
rect 11480 915 11520 920
rect 11480 885 11485 915
rect 11515 885 11520 915
rect 11480 880 11520 885
rect 11590 915 11630 920
rect 11590 885 11595 915
rect 11625 885 11630 915
rect 11590 880 11630 885
rect 11700 915 11740 920
rect 11700 885 11705 915
rect 11735 885 11740 915
rect 11700 880 11740 885
rect 11810 915 11850 920
rect 11810 885 11815 915
rect 11845 885 11850 915
rect 11810 880 11850 885
rect 11920 915 11960 920
rect 11920 885 11925 915
rect 11955 885 11960 915
rect 11920 880 11960 885
rect 12030 915 12070 920
rect 12030 885 12035 915
rect 12065 885 12070 915
rect 12030 880 12070 885
rect 12140 915 12180 920
rect 12140 885 12145 915
rect 12175 885 12180 915
rect 12140 880 12180 885
rect 12250 915 12290 920
rect 12250 885 12255 915
rect 12285 885 12290 915
rect 12250 880 12290 885
rect 12360 915 12400 920
rect 12360 885 12365 915
rect 12395 885 12400 915
rect 12360 880 12400 885
rect 12470 915 12510 920
rect 12470 885 12475 915
rect 12505 885 12510 915
rect 12470 880 12510 885
rect 12620 915 12660 920
rect 12620 885 12625 915
rect 12655 885 12660 915
rect 12620 880 12660 885
rect 11935 860 11975 865
rect 11005 855 11045 860
rect 11005 825 11010 855
rect 11040 825 11045 855
rect 11005 820 11045 825
rect 11495 855 11535 860
rect 11495 825 11500 855
rect 11530 825 11535 855
rect 11935 830 11940 860
rect 11970 830 11975 860
rect 11935 825 11975 830
rect 12155 860 12195 865
rect 12155 830 12160 860
rect 12190 830 12195 860
rect 12155 825 12195 830
rect 12375 860 12415 865
rect 12375 830 12380 860
rect 12410 830 12415 860
rect 12375 825 12415 830
rect 11495 820 11535 825
rect 11945 805 11965 825
rect 12165 805 12185 825
rect 12385 805 12405 825
rect 12815 805 12835 1215
rect 12870 865 12890 3695
rect 13000 3635 13040 3640
rect 13000 3605 13005 3635
rect 13035 3605 13040 3635
rect 13000 3600 13040 3605
rect 13110 3635 13150 3640
rect 13110 3605 13115 3635
rect 13145 3605 13150 3635
rect 13110 3600 13150 3605
rect 13220 3635 13260 3640
rect 13220 3605 13225 3635
rect 13255 3605 13260 3635
rect 13220 3600 13260 3605
rect 13330 3635 13370 3640
rect 13330 3605 13335 3635
rect 13365 3605 13370 3635
rect 13330 3600 13370 3605
rect 13440 3635 13480 3640
rect 13440 3605 13445 3635
rect 13475 3605 13480 3635
rect 13440 3600 13480 3605
rect 13550 3635 13590 3640
rect 13550 3605 13555 3635
rect 13585 3605 13590 3635
rect 13550 3600 13590 3605
rect 26340 3625 26380 3630
rect 26340 3595 26345 3625
rect 26375 3595 26380 3625
rect 26340 3590 26380 3595
rect 26460 3625 26500 3630
rect 26460 3595 26465 3625
rect 26495 3595 26500 3625
rect 26460 3590 26500 3595
rect 26580 3625 26620 3630
rect 26580 3595 26585 3625
rect 26615 3595 26620 3625
rect 26580 3590 26620 3595
rect 26700 3625 26740 3630
rect 26700 3595 26705 3625
rect 26735 3595 26740 3625
rect 26700 3590 26740 3595
rect 26820 3625 26860 3630
rect 26820 3595 26825 3625
rect 26855 3595 26860 3625
rect 26820 3590 26860 3595
rect 26940 3625 26980 3630
rect 26940 3595 26945 3625
rect 26975 3595 26980 3625
rect 26940 3590 26980 3595
rect 27060 3625 27100 3630
rect 27060 3595 27065 3625
rect 27095 3595 27100 3625
rect 27060 3590 27100 3595
rect 27180 3625 27220 3630
rect 27180 3595 27185 3625
rect 27215 3595 27220 3625
rect 27180 3590 27220 3595
rect 27300 3625 27340 3630
rect 27300 3595 27305 3625
rect 27335 3595 27340 3625
rect 27300 3590 27340 3595
rect 27420 3625 27460 3630
rect 27420 3595 27425 3625
rect 27455 3595 27460 3625
rect 27420 3590 27460 3595
rect 13760 3555 13901 3560
rect 13760 3525 13765 3555
rect 13795 3525 13815 3555
rect 13845 3525 13865 3555
rect 13895 3550 13901 3555
rect 13895 3530 13905 3550
rect 13895 3525 13901 3530
rect 13760 3520 13901 3525
rect 27945 3290 27985 3295
rect 27945 3260 27950 3290
rect 27980 3260 27985 3290
rect 27945 3255 27985 3260
rect 28055 3290 28095 3295
rect 28055 3260 28060 3290
rect 28090 3260 28095 3290
rect 28055 3255 28095 3260
rect 28165 3290 28205 3295
rect 28165 3260 28170 3290
rect 28200 3260 28205 3290
rect 28165 3255 28205 3260
rect 28275 3290 28315 3295
rect 28275 3260 28280 3290
rect 28310 3260 28315 3290
rect 28275 3255 28315 3260
rect 28385 3290 28425 3295
rect 28385 3260 28390 3290
rect 28420 3260 28425 3290
rect 28385 3255 28425 3260
rect 28495 3290 28535 3295
rect 28495 3260 28500 3290
rect 28530 3260 28535 3290
rect 28495 3255 28535 3260
rect 28605 3290 28645 3295
rect 28605 3260 28610 3290
rect 28640 3260 28645 3290
rect 28605 3255 28645 3260
rect 28715 3290 28755 3295
rect 28715 3260 28720 3290
rect 28750 3260 28755 3290
rect 28715 3255 28755 3260
rect 28825 3290 28865 3295
rect 28825 3260 28830 3290
rect 28860 3260 28865 3290
rect 28825 3255 28865 3260
rect 28935 3290 28975 3295
rect 28935 3260 28940 3290
rect 28970 3260 28975 3290
rect 28935 3255 28975 3260
rect 29045 3290 29085 3295
rect 29045 3260 29050 3290
rect 29080 3260 29085 3290
rect 29045 3255 29085 3260
rect 25580 3210 25620 3215
rect 25580 3180 25585 3210
rect 25615 3180 25620 3210
rect 25580 3175 25620 3180
rect 25905 3205 25940 3215
rect 25905 3185 25910 3205
rect 25930 3185 25940 3205
rect 25905 3175 25940 3185
rect 25980 3210 26015 3215
rect 25980 3180 25985 3210
rect 25980 3175 26015 3180
rect 25910 3160 25930 3175
rect 25900 3155 25940 3160
rect 25900 3125 25905 3155
rect 25935 3125 25940 3155
rect 25900 3120 25940 3125
rect 13055 2965 13095 2970
rect 13055 2935 13060 2965
rect 13090 2935 13095 2965
rect 13055 2930 13095 2935
rect 13113 2960 13147 2970
rect 13113 2940 13121 2960
rect 13139 2940 13147 2960
rect 13113 2930 13147 2940
rect 13165 2965 13205 2970
rect 13165 2935 13170 2965
rect 13200 2935 13205 2965
rect 13165 2930 13205 2935
rect 13275 2965 13315 2970
rect 13275 2935 13280 2965
rect 13310 2935 13315 2965
rect 13275 2930 13315 2935
rect 13385 2965 13425 2970
rect 13385 2935 13390 2965
rect 13420 2935 13425 2965
rect 13385 2930 13425 2935
rect 13495 2965 13535 2970
rect 13495 2935 13500 2965
rect 13530 2935 13535 2965
rect 13495 2930 13535 2935
rect 13760 2935 13901 2940
rect 13120 2885 13140 2930
rect 13110 2880 13150 2885
rect 13110 2850 13115 2880
rect 13145 2850 13150 2880
rect 13110 2845 13150 2850
rect 13395 2830 13415 2930
rect 13760 2905 13765 2935
rect 13795 2905 13815 2935
rect 13845 2905 13865 2935
rect 13895 2905 13901 2935
rect 13760 2900 13901 2905
rect 13820 2885 13840 2900
rect 13810 2880 13850 2885
rect 13810 2850 13815 2880
rect 13845 2850 13850 2880
rect 13810 2845 13850 2850
rect 13385 2825 13425 2830
rect 13385 2795 13390 2825
rect 13420 2795 13425 2825
rect 13385 2790 13425 2795
rect 14015 2825 14055 2830
rect 14015 2795 14020 2825
rect 14050 2795 14055 2825
rect 14015 2790 14055 2795
rect 13000 2705 13040 2710
rect 13000 2675 13005 2705
rect 13035 2675 13040 2705
rect 13000 2670 13040 2675
rect 13110 2705 13150 2710
rect 13110 2675 13115 2705
rect 13145 2675 13150 2705
rect 13110 2670 13150 2675
rect 13220 2705 13260 2710
rect 13220 2675 13225 2705
rect 13255 2675 13260 2705
rect 13220 2670 13260 2675
rect 13330 2705 13370 2710
rect 13330 2675 13335 2705
rect 13365 2675 13370 2705
rect 13330 2670 13370 2675
rect 13440 2705 13480 2710
rect 13440 2675 13445 2705
rect 13475 2675 13480 2705
rect 13440 2670 13480 2675
rect 13550 2705 13590 2710
rect 13550 2675 13555 2705
rect 13585 2675 13590 2705
rect 13550 2670 13590 2675
rect 13055 2435 13095 2440
rect 13055 2405 13060 2435
rect 13090 2405 13095 2435
rect 13055 2400 13095 2405
rect 13165 2435 13205 2440
rect 13165 2405 13170 2435
rect 13200 2405 13205 2435
rect 13165 2400 13205 2405
rect 13275 2435 13315 2440
rect 13275 2405 13280 2435
rect 13310 2405 13315 2435
rect 13275 2400 13315 2405
rect 13385 2435 13425 2440
rect 13385 2405 13390 2435
rect 13420 2405 13425 2435
rect 13385 2400 13425 2405
rect 13495 2435 13535 2440
rect 13495 2405 13500 2435
rect 13530 2405 13535 2435
rect 13495 2400 13535 2405
rect 13740 2435 13780 2440
rect 13740 2405 13745 2435
rect 13775 2405 13780 2435
rect 13740 2400 13780 2405
rect 13025 2375 13065 2380
rect 13025 2345 13030 2375
rect 13060 2345 13065 2375
rect 13025 2340 13065 2345
rect 13055 2315 13095 2320
rect 13055 2285 13060 2315
rect 13090 2285 13095 2315
rect 13055 2280 13095 2285
rect 13165 2315 13205 2320
rect 13165 2285 13170 2315
rect 13200 2285 13205 2315
rect 13165 2280 13205 2285
rect 13275 2315 13315 2320
rect 13275 2285 13280 2315
rect 13310 2285 13315 2315
rect 13275 2280 13315 2285
rect 13385 2315 13425 2320
rect 13385 2285 13390 2315
rect 13420 2285 13425 2315
rect 13385 2280 13425 2285
rect 13495 2315 13535 2320
rect 13495 2285 13500 2315
rect 13530 2285 13535 2315
rect 13495 2280 13535 2285
rect 13695 2315 13735 2320
rect 13695 2285 13700 2315
rect 13730 2285 13735 2315
rect 13695 2280 13735 2285
rect 13705 1950 13725 2280
rect 13750 2005 13770 2400
rect 13795 2005 13830 2010
rect 13740 2000 13780 2005
rect 13740 1970 13745 2000
rect 13775 1970 13780 2000
rect 13740 1965 13780 1970
rect 13795 1965 13830 1970
rect 13855 2005 13890 2011
rect 13855 1965 13890 1970
rect 13915 2005 13950 2010
rect 13915 1965 13950 1970
rect 13975 2005 14010 2011
rect 13975 1965 14010 1970
rect 13860 1950 13880 1965
rect 13000 1945 13040 1950
rect 13000 1915 13005 1945
rect 13035 1915 13040 1945
rect 13000 1910 13040 1915
rect 13110 1945 13150 1950
rect 13110 1915 13115 1945
rect 13145 1915 13150 1945
rect 13110 1910 13150 1915
rect 13220 1945 13260 1950
rect 13220 1915 13225 1945
rect 13255 1915 13260 1945
rect 13220 1910 13260 1915
rect 13330 1945 13370 1950
rect 13330 1915 13335 1945
rect 13365 1915 13370 1945
rect 13330 1910 13370 1915
rect 13440 1945 13480 1950
rect 13440 1915 13445 1945
rect 13475 1915 13480 1945
rect 13440 1910 13480 1915
rect 13550 1945 13590 1950
rect 13550 1915 13555 1945
rect 13585 1915 13590 1945
rect 13550 1910 13590 1915
rect 13695 1945 13735 1950
rect 13695 1915 13700 1945
rect 13730 1915 13735 1945
rect 13695 1910 13735 1915
rect 13850 1945 13890 1950
rect 13850 1915 13855 1945
rect 13885 1915 13890 1945
rect 13850 1910 13890 1915
rect 13980 1900 14000 1965
rect 13970 1895 14010 1900
rect 13970 1865 13975 1895
rect 14005 1865 14010 1895
rect 13970 1860 14010 1865
rect 13205 1760 13245 1765
rect 13205 1730 13210 1760
rect 13240 1730 13245 1760
rect 13205 1725 13245 1730
rect 13795 1760 13835 1765
rect 13795 1730 13800 1760
rect 13830 1730 13835 1760
rect 13795 1725 13835 1730
rect 13215 1710 13235 1725
rect 12925 1705 12965 1710
rect 12925 1675 12930 1705
rect 12960 1675 12965 1705
rect 12925 1670 12965 1675
rect 13105 1705 13145 1710
rect 13105 1675 13110 1705
rect 13140 1675 13145 1705
rect 13105 1670 13145 1675
rect 13208 1700 13242 1710
rect 13208 1680 13216 1700
rect 13234 1680 13242 1700
rect 13208 1670 13242 1680
rect 13305 1705 13345 1710
rect 13305 1675 13310 1705
rect 13340 1675 13345 1705
rect 13305 1670 13345 1675
rect 13505 1705 13545 1710
rect 13505 1675 13510 1705
rect 13540 1675 13545 1705
rect 13505 1670 13545 1675
rect 13730 1705 13770 1710
rect 13730 1675 13735 1705
rect 13765 1675 13770 1705
rect 13730 1670 13770 1675
rect 12935 1395 12955 1670
rect 13740 1650 13760 1670
rect 13805 1650 13825 1725
rect 14025 1710 14045 2790
rect 24735 2670 24775 2675
rect 24735 2640 24740 2670
rect 24770 2640 24775 2670
rect 24735 2635 24775 2640
rect 24845 2670 24885 2675
rect 24845 2640 24850 2670
rect 24880 2640 24885 2670
rect 24845 2635 24885 2640
rect 24955 2670 24995 2675
rect 24955 2640 24960 2670
rect 24990 2640 24995 2670
rect 24955 2635 24995 2640
rect 25065 2670 25105 2675
rect 25065 2640 25070 2670
rect 25100 2640 25105 2670
rect 25065 2635 25105 2640
rect 25175 2670 25215 2675
rect 25175 2640 25180 2670
rect 25210 2640 25215 2670
rect 25175 2635 25215 2640
rect 25285 2670 25325 2675
rect 25285 2640 25290 2670
rect 25320 2640 25325 2670
rect 25285 2635 25325 2640
rect 25395 2670 25435 2675
rect 25395 2640 25400 2670
rect 25430 2640 25435 2670
rect 25395 2635 25435 2640
rect 25505 2670 25545 2675
rect 25505 2640 25510 2670
rect 25540 2640 25545 2670
rect 25505 2635 25545 2640
rect 25615 2670 25655 2675
rect 25615 2640 25620 2670
rect 25650 2640 25655 2670
rect 25615 2635 25655 2640
rect 25725 2670 25765 2675
rect 25725 2640 25730 2670
rect 25760 2640 25765 2670
rect 25725 2635 25765 2640
rect 25835 2670 25875 2675
rect 25835 2640 25840 2670
rect 25870 2640 25875 2670
rect 25835 2635 25875 2640
rect 24790 2500 24830 2505
rect 24790 2470 24795 2500
rect 24825 2470 24830 2500
rect 24790 2465 24830 2470
rect 24900 2500 24940 2505
rect 24900 2470 24905 2500
rect 24935 2470 24940 2500
rect 24900 2465 24940 2470
rect 25010 2500 25050 2505
rect 25010 2470 25015 2500
rect 25045 2470 25050 2500
rect 25010 2465 25050 2470
rect 25120 2500 25160 2505
rect 25120 2470 25125 2500
rect 25155 2470 25160 2500
rect 25120 2465 25160 2470
rect 25230 2500 25270 2505
rect 25230 2470 25235 2500
rect 25265 2470 25270 2500
rect 25230 2465 25270 2470
rect 25340 2500 25380 2505
rect 25340 2470 25345 2500
rect 25375 2470 25380 2500
rect 25340 2465 25380 2470
rect 25450 2500 25490 2505
rect 25450 2470 25455 2500
rect 25485 2470 25490 2500
rect 25450 2465 25490 2470
rect 25560 2500 25600 2505
rect 25560 2470 25565 2500
rect 25595 2470 25600 2500
rect 25560 2465 25600 2470
rect 25670 2500 25710 2505
rect 25670 2470 25675 2500
rect 25705 2470 25710 2500
rect 25670 2465 25710 2470
rect 25780 2500 25820 2505
rect 25780 2470 25785 2500
rect 25815 2470 25820 2500
rect 25990 2480 26010 3175
rect 26280 3150 26320 3160
rect 26280 3130 26290 3150
rect 26310 3130 26320 3150
rect 26280 3120 26320 3130
rect 26400 3150 26440 3160
rect 26400 3130 26410 3150
rect 26430 3130 26440 3150
rect 26400 3120 26440 3130
rect 26520 3150 26560 3160
rect 26520 3130 26530 3150
rect 26550 3130 26560 3150
rect 26520 3120 26560 3130
rect 26640 3150 26680 3160
rect 26640 3130 26650 3150
rect 26670 3130 26680 3150
rect 26640 3120 26680 3130
rect 26760 3150 26800 3160
rect 26760 3130 26770 3150
rect 26790 3130 26800 3150
rect 26760 3120 26800 3130
rect 26823 3155 26857 3160
rect 26823 3125 26826 3155
rect 26854 3125 26857 3155
rect 26823 3120 26857 3125
rect 26880 3150 26920 3160
rect 26880 3130 26890 3150
rect 26910 3130 26920 3150
rect 26880 3120 26920 3130
rect 27000 3150 27040 3160
rect 27000 3130 27010 3150
rect 27030 3130 27040 3150
rect 27000 3120 27040 3130
rect 27120 3150 27160 3160
rect 27120 3130 27130 3150
rect 27150 3130 27160 3150
rect 27120 3120 27160 3130
rect 27240 3150 27280 3160
rect 27240 3130 27250 3150
rect 27270 3130 27280 3150
rect 27240 3120 27280 3130
rect 27360 3150 27400 3160
rect 27360 3130 27370 3150
rect 27390 3130 27400 3150
rect 27360 3120 27400 3130
rect 27480 3150 27520 3160
rect 27480 3130 27490 3150
rect 27510 3130 27520 3150
rect 27480 3120 27520 3130
rect 26290 3105 26310 3120
rect 26280 3100 26320 3105
rect 26280 3070 26285 3100
rect 26315 3070 26320 3100
rect 26280 3065 26320 3070
rect 26410 3060 26430 3120
rect 26530 3105 26550 3120
rect 26520 3100 26560 3105
rect 26520 3070 26525 3100
rect 26555 3070 26560 3100
rect 26520 3065 26560 3070
rect 26650 3060 26670 3120
rect 26770 3105 26790 3120
rect 26760 3100 26800 3105
rect 26760 3070 26765 3100
rect 26795 3070 26800 3100
rect 26760 3065 26800 3070
rect 26890 3060 26910 3120
rect 27010 3105 27030 3120
rect 27000 3100 27040 3105
rect 27000 3070 27005 3100
rect 27035 3070 27040 3100
rect 27000 3065 27040 3070
rect 27130 3060 27150 3120
rect 27250 3105 27270 3120
rect 27240 3100 27280 3105
rect 27240 3070 27245 3100
rect 27275 3070 27280 3100
rect 27240 3065 27280 3070
rect 27370 3060 27390 3120
rect 27490 3105 27510 3120
rect 27480 3100 27520 3105
rect 27480 3070 27485 3100
rect 27515 3070 27520 3100
rect 27480 3065 27520 3070
rect 26400 3055 26440 3060
rect 26400 3025 26405 3055
rect 26435 3025 26440 3055
rect 26400 3020 26440 3025
rect 26640 3055 26680 3060
rect 26640 3025 26645 3055
rect 26675 3025 26680 3055
rect 26640 3020 26680 3025
rect 26880 3055 26920 3060
rect 26880 3025 26885 3055
rect 26915 3025 26920 3055
rect 26880 3020 26920 3025
rect 27120 3055 27160 3060
rect 27120 3025 27125 3055
rect 27155 3025 27160 3055
rect 27120 3020 27160 3025
rect 27360 3055 27400 3060
rect 27360 3025 27365 3055
rect 27395 3025 27400 3055
rect 27360 3020 27400 3025
rect 26410 3005 26430 3020
rect 26340 3000 26380 3005
rect 26340 2970 26345 3000
rect 26375 2970 26380 3000
rect 26340 2965 26380 2970
rect 26400 3000 26440 3005
rect 26400 2970 26405 3000
rect 26435 2970 26440 3000
rect 26400 2965 26440 2970
rect 26580 3000 26620 3005
rect 26580 2970 26585 3000
rect 26615 2970 26620 3000
rect 26580 2965 26620 2970
rect 26820 3000 26860 3005
rect 26820 2970 26825 3000
rect 26855 2970 26860 3000
rect 26820 2965 26860 2970
rect 27060 3000 27100 3005
rect 27060 2970 27065 3000
rect 27095 2970 27100 3000
rect 27060 2965 27100 2970
rect 27300 3000 27340 3005
rect 27300 2970 27305 3000
rect 27335 2970 27340 3000
rect 27300 2965 27340 2970
rect 26350 2950 26370 2965
rect 26590 2950 26610 2965
rect 26830 2950 26850 2965
rect 27070 2950 27090 2965
rect 27310 2950 27330 2965
rect 27490 2950 27510 3065
rect 26340 2940 26380 2950
rect 26340 2920 26350 2940
rect 26370 2920 26380 2940
rect 26340 2910 26380 2920
rect 26460 2945 26500 2950
rect 26460 2915 26465 2945
rect 26495 2915 26500 2945
rect 26460 2910 26500 2915
rect 26580 2940 26620 2950
rect 26580 2920 26590 2940
rect 26610 2920 26620 2940
rect 26580 2910 26620 2920
rect 26700 2945 26740 2950
rect 26700 2915 26705 2945
rect 26735 2915 26740 2945
rect 26700 2910 26740 2915
rect 26820 2940 26860 2950
rect 26820 2920 26830 2940
rect 26850 2920 26860 2940
rect 26820 2910 26860 2920
rect 26940 2945 26980 2950
rect 26940 2915 26945 2945
rect 26975 2915 26980 2945
rect 26940 2910 26980 2915
rect 27060 2940 27100 2950
rect 27060 2920 27070 2940
rect 27090 2920 27100 2940
rect 27060 2910 27100 2920
rect 27180 2945 27220 2950
rect 27180 2915 27185 2945
rect 27215 2915 27220 2945
rect 27180 2910 27220 2915
rect 27300 2940 27340 2950
rect 27300 2920 27310 2940
rect 27330 2920 27340 2940
rect 27300 2910 27340 2920
rect 27420 2945 27460 2950
rect 27420 2915 27425 2945
rect 27455 2915 27460 2945
rect 27420 2910 27460 2915
rect 27480 2945 27520 2950
rect 27480 2915 27485 2945
rect 27515 2915 27520 2945
rect 27480 2910 27520 2915
rect 28000 2920 28040 2925
rect 28000 2890 28005 2920
rect 28035 2890 28040 2920
rect 28000 2885 28040 2890
rect 28058 2915 28092 2925
rect 28058 2895 28066 2915
rect 28084 2895 28092 2915
rect 28058 2885 28092 2895
rect 28110 2920 28150 2925
rect 28110 2890 28115 2920
rect 28145 2890 28150 2920
rect 28110 2885 28150 2890
rect 28220 2920 28260 2925
rect 28220 2890 28225 2920
rect 28255 2890 28260 2920
rect 28220 2885 28260 2890
rect 28330 2920 28370 2925
rect 28330 2890 28335 2920
rect 28365 2890 28370 2920
rect 28330 2885 28370 2890
rect 28440 2920 28480 2925
rect 28440 2890 28445 2920
rect 28475 2890 28480 2920
rect 28440 2885 28480 2890
rect 28550 2920 28590 2925
rect 28550 2890 28555 2920
rect 28585 2890 28590 2920
rect 28550 2885 28590 2890
rect 28660 2920 28700 2925
rect 28660 2890 28665 2920
rect 28695 2890 28700 2920
rect 28660 2885 28700 2890
rect 28770 2920 28810 2925
rect 28770 2890 28775 2920
rect 28805 2890 28810 2920
rect 28770 2885 28810 2890
rect 28880 2920 28920 2925
rect 28880 2890 28885 2920
rect 28915 2890 28920 2920
rect 28880 2885 28920 2890
rect 28990 2920 29030 2925
rect 28990 2890 28995 2920
rect 29025 2890 29030 2920
rect 28990 2885 29030 2890
rect 28065 2836 28085 2885
rect 28055 2830 28095 2836
rect 28055 2800 28060 2830
rect 28090 2800 28095 2830
rect 28055 2780 28095 2800
rect 28055 2750 28060 2780
rect 28090 2750 28095 2780
rect 27690 2730 27730 2735
rect 27690 2700 27695 2730
rect 27725 2700 27730 2730
rect 27690 2695 27730 2700
rect 28055 2730 28095 2750
rect 28055 2700 28060 2730
rect 28090 2700 28095 2730
rect 28055 2695 28095 2700
rect 25780 2465 25820 2470
rect 25980 2475 26020 2480
rect 24800 2380 24820 2465
rect 25980 2445 25985 2475
rect 26015 2445 26020 2475
rect 25813 2440 25847 2445
rect 25980 2440 26020 2445
rect 26280 2470 26320 2480
rect 26280 2450 26290 2470
rect 26310 2450 26320 2470
rect 26280 2440 26320 2450
rect 26400 2470 26440 2480
rect 26400 2450 26410 2470
rect 26430 2450 26440 2470
rect 26400 2440 26440 2450
rect 26520 2470 26560 2480
rect 26520 2450 26530 2470
rect 26550 2450 26560 2470
rect 26520 2440 26560 2450
rect 26640 2470 26680 2480
rect 26640 2450 26650 2470
rect 26670 2450 26680 2470
rect 26640 2440 26680 2450
rect 26760 2470 26800 2480
rect 26760 2450 26770 2470
rect 26790 2450 26800 2470
rect 26760 2440 26800 2450
rect 26823 2475 26857 2480
rect 26823 2445 26826 2475
rect 26854 2445 26857 2475
rect 26823 2440 26857 2445
rect 26880 2470 26920 2480
rect 26880 2450 26890 2470
rect 26910 2450 26920 2470
rect 26880 2440 26920 2450
rect 27000 2470 27040 2480
rect 27000 2450 27010 2470
rect 27030 2450 27040 2470
rect 27000 2440 27040 2450
rect 27120 2470 27160 2480
rect 27120 2450 27130 2470
rect 27150 2450 27160 2470
rect 27120 2440 27160 2450
rect 27240 2470 27280 2480
rect 27240 2450 27250 2470
rect 27270 2450 27280 2470
rect 27240 2440 27280 2450
rect 27360 2470 27400 2480
rect 27360 2450 27370 2470
rect 27390 2450 27400 2470
rect 27360 2440 27400 2450
rect 27480 2470 27520 2480
rect 27480 2450 27490 2470
rect 27510 2450 27520 2470
rect 27480 2440 27520 2450
rect 25813 2410 25816 2440
rect 25844 2410 25847 2440
rect 26290 2425 26310 2440
rect 25813 2405 25847 2410
rect 26280 2420 26320 2425
rect 24800 2345 24805 2380
rect 24840 2345 24845 2380
rect 25635 2345 25640 2380
rect 25675 2345 25680 2380
rect 25635 2320 25680 2345
rect 24800 2285 24805 2320
rect 24840 2285 24845 2320
rect 25635 2285 25640 2320
rect 25675 2285 25680 2320
rect 25820 2285 25840 2405
rect 26280 2390 26285 2420
rect 26315 2390 26320 2420
rect 26280 2385 26320 2390
rect 26410 2380 26430 2440
rect 26530 2425 26550 2440
rect 26520 2420 26560 2425
rect 26520 2390 26525 2420
rect 26555 2390 26560 2420
rect 26520 2385 26560 2390
rect 26650 2380 26670 2440
rect 26770 2425 26790 2440
rect 26760 2420 26800 2425
rect 26760 2390 26765 2420
rect 26795 2390 26800 2420
rect 26760 2385 26800 2390
rect 26400 2375 26440 2380
rect 26400 2345 26405 2375
rect 26435 2345 26440 2375
rect 26400 2340 26440 2345
rect 26640 2375 26680 2380
rect 26640 2345 26645 2375
rect 26675 2345 26680 2375
rect 26640 2340 26680 2345
rect 24800 2225 24820 2285
rect 25813 2280 25847 2285
rect 25813 2250 25816 2280
rect 25844 2250 25847 2280
rect 25813 2245 25847 2250
rect 26440 2280 26480 2285
rect 26440 2250 26445 2280
rect 26475 2250 26480 2280
rect 26440 2245 26480 2250
rect 26660 2280 26700 2285
rect 26660 2250 26665 2280
rect 26695 2250 26700 2280
rect 26660 2245 26700 2250
rect 26330 2235 26370 2240
rect 24790 2220 24830 2225
rect 24790 2190 24795 2220
rect 24825 2190 24830 2220
rect 24790 2185 24830 2190
rect 24900 2220 24940 2225
rect 24900 2190 24905 2220
rect 24935 2190 24940 2220
rect 24900 2185 24940 2190
rect 25010 2220 25050 2225
rect 25010 2190 25015 2220
rect 25045 2190 25050 2220
rect 25010 2185 25050 2190
rect 25120 2220 25160 2225
rect 25120 2190 25125 2220
rect 25155 2190 25160 2220
rect 25120 2185 25160 2190
rect 25230 2220 25270 2225
rect 25230 2190 25235 2220
rect 25265 2190 25270 2220
rect 25230 2185 25270 2190
rect 25340 2220 25380 2225
rect 25340 2190 25345 2220
rect 25375 2190 25380 2220
rect 25340 2185 25380 2190
rect 25450 2220 25490 2225
rect 25450 2190 25455 2220
rect 25485 2190 25490 2220
rect 25450 2185 25490 2190
rect 25560 2220 25600 2225
rect 25560 2190 25565 2220
rect 25595 2190 25600 2220
rect 25560 2185 25600 2190
rect 25670 2220 25710 2225
rect 25670 2190 25675 2220
rect 25705 2190 25710 2220
rect 25670 2185 25710 2190
rect 25780 2220 25820 2225
rect 25780 2190 25785 2220
rect 25815 2190 25820 2220
rect 26330 2205 26335 2235
rect 26365 2205 26370 2235
rect 26330 2200 26370 2205
rect 25780 2185 25820 2190
rect 26340 2185 26360 2200
rect 26450 2185 26470 2245
rect 26550 2235 26590 2240
rect 26550 2205 26555 2235
rect 26585 2205 26590 2235
rect 26550 2200 26590 2205
rect 26560 2185 26580 2200
rect 26670 2185 26690 2245
rect 26770 2240 26790 2385
rect 26890 2380 26910 2440
rect 27010 2425 27030 2440
rect 27000 2420 27040 2425
rect 27000 2390 27005 2420
rect 27035 2390 27040 2420
rect 27000 2385 27040 2390
rect 27130 2380 27150 2440
rect 27250 2425 27270 2440
rect 27240 2420 27280 2425
rect 27240 2390 27245 2420
rect 27275 2390 27280 2420
rect 27240 2385 27280 2390
rect 27370 2380 27390 2440
rect 27490 2425 27510 2440
rect 27480 2420 27520 2425
rect 27480 2390 27485 2420
rect 27515 2390 27520 2420
rect 27480 2385 27520 2390
rect 27700 2380 27720 2695
rect 27945 2670 27985 2675
rect 27945 2640 27950 2670
rect 27980 2640 27985 2670
rect 27945 2635 27985 2640
rect 28055 2670 28095 2675
rect 28055 2640 28060 2670
rect 28090 2640 28095 2670
rect 28055 2635 28095 2640
rect 28165 2670 28205 2675
rect 28165 2640 28170 2670
rect 28200 2640 28205 2670
rect 28165 2635 28205 2640
rect 28275 2670 28315 2675
rect 28275 2640 28280 2670
rect 28310 2640 28315 2670
rect 28275 2635 28315 2640
rect 28385 2670 28425 2675
rect 28385 2640 28390 2670
rect 28420 2640 28425 2670
rect 28385 2635 28425 2640
rect 28495 2670 28535 2675
rect 28495 2640 28500 2670
rect 28530 2640 28535 2670
rect 28495 2635 28535 2640
rect 28605 2670 28645 2675
rect 28605 2640 28610 2670
rect 28640 2640 28645 2670
rect 28605 2635 28645 2640
rect 28715 2670 28755 2675
rect 28715 2640 28720 2670
rect 28750 2640 28755 2670
rect 28715 2635 28755 2640
rect 28825 2670 28865 2675
rect 28825 2640 28830 2670
rect 28860 2640 28865 2670
rect 28825 2635 28865 2640
rect 28935 2670 28975 2675
rect 28935 2640 28940 2670
rect 28970 2640 28975 2670
rect 28935 2635 28975 2640
rect 29045 2670 29085 2675
rect 29045 2640 29050 2670
rect 29080 2640 29085 2670
rect 29045 2635 29085 2640
rect 28000 2500 28040 2505
rect 28000 2470 28005 2500
rect 28035 2470 28040 2500
rect 28000 2465 28040 2470
rect 28110 2500 28150 2505
rect 28110 2470 28115 2500
rect 28145 2470 28150 2500
rect 28110 2465 28150 2470
rect 28220 2500 28260 2505
rect 28220 2470 28225 2500
rect 28255 2470 28260 2500
rect 28220 2465 28260 2470
rect 28330 2500 28370 2505
rect 28330 2470 28335 2500
rect 28365 2470 28370 2500
rect 28330 2465 28370 2470
rect 28440 2500 28480 2505
rect 28440 2470 28445 2500
rect 28475 2470 28480 2500
rect 28440 2465 28480 2470
rect 28550 2500 28590 2505
rect 28550 2470 28555 2500
rect 28585 2470 28590 2500
rect 28550 2465 28590 2470
rect 28660 2500 28700 2505
rect 28660 2470 28665 2500
rect 28695 2470 28700 2500
rect 28660 2465 28700 2470
rect 28770 2500 28810 2505
rect 28770 2470 28775 2500
rect 28805 2470 28810 2500
rect 28770 2465 28810 2470
rect 28880 2500 28920 2505
rect 28880 2470 28885 2500
rect 28915 2470 28920 2500
rect 28880 2465 28920 2470
rect 28990 2500 29030 2505
rect 28990 2470 28995 2500
rect 29025 2470 29030 2500
rect 28990 2465 29030 2470
rect 27973 2440 28007 2445
rect 27973 2410 27976 2440
rect 28004 2410 28007 2440
rect 27973 2405 28007 2410
rect 27980 2380 28000 2405
rect 29000 2380 29020 2465
rect 26880 2375 26920 2380
rect 26880 2345 26885 2375
rect 26915 2345 26920 2375
rect 26880 2340 26920 2345
rect 27120 2375 27160 2380
rect 27120 2345 27125 2375
rect 27155 2345 27160 2375
rect 27120 2340 27160 2345
rect 27360 2375 27400 2380
rect 27360 2345 27365 2375
rect 27395 2345 27400 2375
rect 27360 2340 27400 2345
rect 27690 2375 27730 2380
rect 27690 2345 27695 2375
rect 27725 2345 27730 2375
rect 27690 2340 27730 2345
rect 27970 2375 28010 2380
rect 27970 2345 27975 2375
rect 28005 2345 28010 2375
rect 27970 2340 28010 2345
rect 28140 2345 28145 2380
rect 28180 2345 28185 2380
rect 28974 2345 28980 2380
rect 29015 2345 29020 2380
rect 27120 2285 27140 2340
rect 27815 2325 27855 2330
rect 27815 2295 27820 2325
rect 27850 2295 27855 2325
rect 27815 2290 27855 2295
rect 26880 2280 26920 2285
rect 26880 2250 26885 2280
rect 26915 2250 26920 2280
rect 26880 2245 26920 2250
rect 27100 2280 27140 2285
rect 27100 2250 27105 2280
rect 27135 2250 27140 2280
rect 27100 2245 27140 2250
rect 27320 2280 27360 2285
rect 27320 2250 27325 2280
rect 27355 2250 27360 2280
rect 27320 2245 27360 2250
rect 26770 2235 26810 2240
rect 26770 2205 26775 2235
rect 26805 2205 26810 2235
rect 26770 2200 26810 2205
rect 26780 2185 26800 2200
rect 26890 2185 26910 2245
rect 26990 2235 27030 2240
rect 26990 2205 26995 2235
rect 27025 2205 27030 2235
rect 26990 2200 27030 2205
rect 27000 2185 27020 2200
rect 27110 2185 27130 2245
rect 27210 2235 27250 2240
rect 27210 2205 27215 2235
rect 27245 2205 27250 2235
rect 27210 2200 27250 2205
rect 27220 2185 27240 2200
rect 27330 2185 27350 2245
rect 27430 2235 27470 2240
rect 27430 2205 27435 2235
rect 27465 2205 27470 2235
rect 27430 2200 27470 2205
rect 27440 2185 27460 2200
rect 26330 2175 26370 2185
rect 26330 2155 26340 2175
rect 26360 2155 26370 2175
rect 26330 2145 26370 2155
rect 26440 2175 26480 2185
rect 26440 2155 26450 2175
rect 26470 2155 26480 2175
rect 26440 2145 26480 2155
rect 26550 2175 26590 2185
rect 26550 2155 26560 2175
rect 26580 2155 26590 2175
rect 26550 2145 26590 2155
rect 26660 2175 26700 2185
rect 26660 2155 26670 2175
rect 26690 2155 26700 2175
rect 26660 2145 26700 2155
rect 26770 2175 26810 2185
rect 26770 2155 26780 2175
rect 26800 2155 26810 2175
rect 26770 2145 26810 2155
rect 26880 2175 26920 2185
rect 26880 2155 26890 2175
rect 26910 2155 26920 2175
rect 26880 2145 26920 2155
rect 26990 2175 27030 2185
rect 26990 2155 27000 2175
rect 27020 2155 27030 2175
rect 26990 2145 27030 2155
rect 27100 2175 27140 2185
rect 27100 2155 27110 2175
rect 27130 2155 27140 2175
rect 27100 2145 27140 2155
rect 27210 2175 27250 2185
rect 27210 2155 27220 2175
rect 27240 2155 27250 2175
rect 27210 2145 27250 2155
rect 27320 2175 27360 2185
rect 27320 2155 27330 2175
rect 27350 2155 27360 2175
rect 27320 2145 27360 2155
rect 27430 2175 27470 2185
rect 27430 2155 27440 2175
rect 27460 2155 27470 2175
rect 27430 2145 27470 2155
rect 24735 2000 24775 2005
rect 24735 1970 24740 2000
rect 24770 1970 24775 2000
rect 24735 1965 24775 1970
rect 24845 2000 24885 2005
rect 24845 1970 24850 2000
rect 24880 1970 24885 2000
rect 24845 1965 24885 1970
rect 24955 2000 24995 2005
rect 24955 1970 24960 2000
rect 24990 1970 24995 2000
rect 24955 1965 24995 1970
rect 25065 2000 25105 2005
rect 25065 1970 25070 2000
rect 25100 1970 25105 2000
rect 25065 1965 25105 1970
rect 25175 2000 25215 2005
rect 25175 1970 25180 2000
rect 25210 1970 25215 2000
rect 25175 1965 25215 1970
rect 25285 2000 25325 2005
rect 25285 1970 25290 2000
rect 25320 1970 25325 2000
rect 25285 1965 25325 1970
rect 25395 2000 25435 2005
rect 25395 1970 25400 2000
rect 25430 1970 25435 2000
rect 25395 1965 25435 1970
rect 25505 2000 25545 2005
rect 25505 1970 25510 2000
rect 25540 1970 25545 2000
rect 25505 1965 25545 1970
rect 25615 2000 25655 2005
rect 25615 1970 25620 2000
rect 25650 1970 25655 2000
rect 25615 1965 25655 1970
rect 25725 2000 25765 2005
rect 25725 1970 25730 2000
rect 25760 1970 25765 2000
rect 25725 1965 25765 1970
rect 25835 2000 25875 2005
rect 25835 1970 25840 2000
rect 25870 1970 25875 2000
rect 25835 1965 25875 1970
rect 26385 1960 26425 1965
rect 26385 1930 26390 1960
rect 26420 1930 26425 1960
rect 26385 1925 26425 1930
rect 26495 1955 26535 1965
rect 26495 1935 26505 1955
rect 26525 1935 26535 1955
rect 26495 1925 26535 1935
rect 26605 1960 26645 1965
rect 26605 1930 26610 1960
rect 26640 1930 26645 1960
rect 26605 1925 26645 1930
rect 26715 1955 26755 1965
rect 26715 1935 26725 1955
rect 26745 1935 26755 1955
rect 26715 1925 26755 1935
rect 26825 1960 26865 1965
rect 26825 1930 26830 1960
rect 26860 1930 26865 1960
rect 26825 1925 26865 1930
rect 26935 1955 26975 1965
rect 26935 1935 26945 1955
rect 26965 1935 26975 1955
rect 26935 1925 26975 1935
rect 27045 1960 27085 1965
rect 27045 1930 27050 1960
rect 27080 1930 27085 1960
rect 27045 1925 27085 1930
rect 27155 1955 27195 1965
rect 27155 1935 27165 1955
rect 27185 1935 27195 1955
rect 27155 1925 27195 1935
rect 27245 1960 27305 1965
rect 27245 1930 27270 1960
rect 27300 1930 27305 1960
rect 27245 1925 27305 1930
rect 27375 1955 27415 1965
rect 27375 1935 27385 1955
rect 27405 1935 27415 1955
rect 27375 1925 27415 1935
rect 26505 1910 26525 1925
rect 26725 1910 26745 1925
rect 26945 1910 26965 1925
rect 27165 1910 27185 1925
rect 26495 1905 26555 1910
rect 26495 1875 26500 1905
rect 26530 1875 26555 1905
rect 26495 1870 26555 1875
rect 26715 1905 26755 1910
rect 26715 1875 26720 1905
rect 26750 1875 26755 1905
rect 26715 1870 26755 1875
rect 26935 1905 26975 1910
rect 26935 1875 26940 1905
rect 26970 1875 26975 1905
rect 26935 1870 26975 1875
rect 27155 1905 27195 1910
rect 27155 1875 27160 1905
rect 27190 1875 27195 1905
rect 27155 1870 27195 1875
rect 26190 1850 26230 1855
rect 26190 1820 26195 1850
rect 26225 1820 26230 1850
rect 26190 1815 26230 1820
rect 26410 1850 26450 1855
rect 26410 1820 26415 1850
rect 26445 1820 26450 1850
rect 26410 1815 26450 1820
rect 26200 1780 26220 1815
rect 26420 1780 26440 1815
rect 26190 1770 26230 1780
rect 26085 1760 26125 1765
rect 26085 1730 26090 1760
rect 26120 1730 26125 1760
rect 26190 1750 26200 1770
rect 26220 1750 26230 1770
rect 26410 1770 26450 1780
rect 26190 1740 26230 1750
rect 26305 1760 26345 1765
rect 26085 1725 26125 1730
rect 26305 1730 26310 1760
rect 26340 1730 26345 1760
rect 26410 1750 26420 1770
rect 26440 1750 26450 1770
rect 26535 1765 26555 1870
rect 27245 1855 27265 1925
rect 27385 1910 27405 1925
rect 27375 1905 27415 1910
rect 27375 1875 27380 1905
rect 27410 1875 27415 1905
rect 27375 1870 27415 1875
rect 26640 1850 26680 1855
rect 26640 1820 26645 1850
rect 26675 1820 26680 1850
rect 26640 1815 26680 1820
rect 27230 1850 27270 1855
rect 27230 1820 27235 1850
rect 27265 1820 27270 1850
rect 27230 1815 27270 1820
rect 27450 1850 27490 1855
rect 27450 1820 27455 1850
rect 27485 1820 27490 1850
rect 27450 1815 27490 1820
rect 27680 1850 27720 1855
rect 27680 1820 27685 1850
rect 27715 1820 27720 1850
rect 27680 1815 27720 1820
rect 26650 1780 26670 1815
rect 26820 1805 26860 1810
rect 26640 1770 26680 1780
rect 26820 1775 26825 1805
rect 26855 1775 26860 1805
rect 26820 1770 26860 1775
rect 26940 1805 26980 1810
rect 26940 1775 26945 1805
rect 26975 1775 26980 1805
rect 27240 1780 27260 1815
rect 27460 1780 27480 1815
rect 27690 1780 27710 1815
rect 26940 1770 26980 1775
rect 27230 1770 27270 1780
rect 26410 1740 26450 1750
rect 26525 1760 26565 1765
rect 26305 1725 26345 1730
rect 26525 1730 26530 1760
rect 26560 1730 26565 1760
rect 26640 1750 26650 1770
rect 26670 1750 26680 1770
rect 26640 1740 26680 1750
rect 26525 1725 26565 1730
rect 26830 1720 26850 1770
rect 26950 1720 26970 1770
rect 27125 1760 27165 1765
rect 27125 1730 27130 1760
rect 27160 1730 27165 1760
rect 27230 1750 27240 1770
rect 27260 1750 27270 1770
rect 27450 1770 27490 1780
rect 27230 1740 27270 1750
rect 27345 1760 27385 1765
rect 27125 1725 27165 1730
rect 27345 1730 27350 1760
rect 27380 1730 27385 1760
rect 27450 1750 27460 1770
rect 27480 1750 27490 1770
rect 27680 1770 27720 1780
rect 27450 1740 27490 1750
rect 27565 1760 27605 1765
rect 27345 1725 27385 1730
rect 27565 1730 27570 1760
rect 27600 1730 27605 1760
rect 27680 1750 27690 1770
rect 27710 1750 27720 1770
rect 27680 1740 27720 1750
rect 27565 1725 27605 1730
rect 26237 1715 26269 1720
rect 14015 1705 14055 1710
rect 14015 1675 14020 1705
rect 14050 1675 14055 1705
rect 26237 1685 26240 1715
rect 26266 1685 26269 1715
rect 26237 1680 26269 1685
rect 26457 1715 26489 1720
rect 26457 1685 26460 1715
rect 26486 1685 26489 1715
rect 26457 1680 26489 1685
rect 26601 1715 26633 1720
rect 26601 1685 26604 1715
rect 26630 1685 26633 1715
rect 26601 1680 26633 1685
rect 26820 1710 26850 1720
rect 26820 1690 26825 1710
rect 26845 1690 26850 1710
rect 26820 1680 26850 1690
rect 26867 1715 26899 1720
rect 26867 1685 26870 1715
rect 26896 1685 26899 1715
rect 26867 1680 26899 1685
rect 26950 1710 26980 1720
rect 26950 1690 26955 1710
rect 26975 1690 26980 1710
rect 26950 1680 26980 1690
rect 27277 1715 27309 1720
rect 27277 1685 27280 1715
rect 27306 1685 27309 1715
rect 27277 1680 27309 1685
rect 27497 1715 27529 1720
rect 27497 1685 27500 1715
rect 27526 1685 27529 1715
rect 27497 1680 27529 1685
rect 27641 1715 27673 1720
rect 27641 1685 27644 1715
rect 27670 1685 27673 1715
rect 27641 1680 27673 1685
rect 14015 1670 14055 1675
rect 13735 1645 13770 1650
rect 13735 1605 13770 1610
rect 13795 1645 13830 1650
rect 13795 1605 13830 1610
rect 27825 1575 27845 2290
rect 27980 2285 28000 2340
rect 28140 2320 28185 2345
rect 28140 2285 28145 2320
rect 28180 2285 28185 2320
rect 28975 2285 28980 2320
rect 29015 2285 29020 2320
rect 27973 2280 28007 2285
rect 27973 2250 27976 2280
rect 28004 2250 28007 2280
rect 27973 2245 28007 2250
rect 29000 2225 29020 2285
rect 28000 2220 28040 2225
rect 28000 2190 28005 2220
rect 28035 2190 28040 2220
rect 28000 2185 28040 2190
rect 28110 2220 28150 2225
rect 28110 2190 28115 2220
rect 28145 2190 28150 2220
rect 28110 2185 28150 2190
rect 28220 2220 28260 2225
rect 28220 2190 28225 2220
rect 28255 2190 28260 2220
rect 28220 2185 28260 2190
rect 28330 2220 28370 2225
rect 28330 2190 28335 2220
rect 28365 2190 28370 2220
rect 28330 2185 28370 2190
rect 28440 2220 28480 2225
rect 28440 2190 28445 2220
rect 28475 2190 28480 2220
rect 28440 2185 28480 2190
rect 28550 2220 28590 2225
rect 28550 2190 28555 2220
rect 28585 2190 28590 2220
rect 28550 2185 28590 2190
rect 28660 2220 28700 2225
rect 28660 2190 28665 2220
rect 28695 2190 28700 2220
rect 28660 2185 28700 2190
rect 28770 2220 28810 2225
rect 28770 2190 28775 2220
rect 28805 2190 28810 2220
rect 28770 2185 28810 2190
rect 28880 2220 28920 2225
rect 28880 2190 28885 2220
rect 28915 2190 28920 2220
rect 28880 2185 28920 2190
rect 28990 2220 29030 2225
rect 28990 2190 28995 2220
rect 29025 2190 29030 2220
rect 28990 2185 29030 2190
rect 27945 2000 27985 2005
rect 27945 1970 27950 2000
rect 27980 1970 27985 2000
rect 27945 1965 27985 1970
rect 28055 2000 28095 2005
rect 28055 1970 28060 2000
rect 28090 1970 28095 2000
rect 28055 1965 28095 1970
rect 28165 2000 28205 2005
rect 28165 1970 28170 2000
rect 28200 1970 28205 2000
rect 28165 1965 28205 1970
rect 28275 2000 28315 2005
rect 28275 1970 28280 2000
rect 28310 1970 28315 2000
rect 28275 1965 28315 1970
rect 28385 2000 28425 2005
rect 28385 1970 28390 2000
rect 28420 1970 28425 2000
rect 28385 1965 28425 1970
rect 28495 2000 28535 2005
rect 28495 1970 28500 2000
rect 28530 1970 28535 2000
rect 28495 1965 28535 1970
rect 28605 2000 28645 2005
rect 28605 1970 28610 2000
rect 28640 1970 28645 2000
rect 28605 1965 28645 1970
rect 28715 2000 28755 2005
rect 28715 1970 28720 2000
rect 28750 1970 28755 2000
rect 28715 1965 28755 1970
rect 28825 2000 28865 2005
rect 28825 1970 28830 2000
rect 28860 1970 28865 2000
rect 28825 1965 28865 1970
rect 28935 2000 28975 2005
rect 28935 1970 28940 2000
rect 28970 1970 28975 2000
rect 28935 1965 28975 1970
rect 29045 2000 29085 2005
rect 29045 1970 29050 2000
rect 29080 1970 29085 2000
rect 29045 1965 29085 1970
rect 28045 1905 28085 1910
rect 28045 1875 28050 1905
rect 28080 1875 28085 1905
rect 28045 1870 28085 1875
rect 28155 1905 28195 1910
rect 28155 1875 28160 1905
rect 28190 1875 28195 1905
rect 28155 1870 28195 1875
rect 28265 1905 28305 1910
rect 28265 1875 28270 1905
rect 28300 1875 28305 1905
rect 28265 1870 28305 1875
rect 28066 1680 28098 1685
rect 28066 1650 28070 1680
rect 28096 1650 28098 1680
rect 28115 1680 28155 1690
rect 28115 1660 28125 1680
rect 28145 1660 28155 1680
rect 28115 1650 28155 1660
rect 28210 1680 28250 1690
rect 28210 1660 28220 1680
rect 28240 1660 28250 1680
rect 28210 1650 28250 1660
rect 28066 1645 28098 1650
rect 28010 1630 28050 1635
rect 28010 1600 28015 1630
rect 28045 1600 28050 1630
rect 28010 1595 28050 1600
rect 28070 1575 28090 1645
rect 28125 1635 28145 1650
rect 28220 1635 28240 1650
rect 28116 1630 28156 1635
rect 28116 1600 28121 1630
rect 28151 1600 28156 1630
rect 28116 1595 28156 1600
rect 28210 1630 28250 1635
rect 28210 1600 28215 1630
rect 28245 1600 28250 1630
rect 28210 1595 28250 1600
rect 28300 1630 28340 1635
rect 28300 1600 28305 1630
rect 28335 1600 28340 1630
rect 28300 1595 28340 1600
rect 27815 1570 27855 1575
rect 27815 1540 27820 1570
rect 27850 1540 27855 1570
rect 27815 1535 27855 1540
rect 27971 1570 28003 1575
rect 27971 1540 27975 1570
rect 28001 1540 28003 1570
rect 27971 1535 28003 1540
rect 28060 1565 28100 1575
rect 28060 1545 28070 1565
rect 28090 1545 28100 1565
rect 28060 1535 28100 1545
rect 28347 1570 28379 1575
rect 28347 1540 28349 1570
rect 28375 1540 28379 1570
rect 28347 1535 28379 1540
rect 26106 1495 26138 1500
rect 26106 1465 26109 1495
rect 26135 1465 26138 1495
rect 26106 1460 26138 1465
rect 26305 1495 26345 1500
rect 26305 1465 26310 1495
rect 26340 1465 26345 1495
rect 26305 1460 26345 1465
rect 26525 1495 26565 1500
rect 26525 1465 26530 1495
rect 26560 1465 26565 1495
rect 26525 1460 26565 1465
rect 26825 1490 26855 1500
rect 26825 1470 26830 1490
rect 26850 1470 26855 1490
rect 26825 1460 26855 1470
rect 26875 1490 26905 1500
rect 26875 1470 26880 1490
rect 26900 1470 26905 1490
rect 26875 1460 26905 1470
rect 26922 1495 26954 1500
rect 26922 1465 26925 1495
rect 26951 1465 26954 1495
rect 26922 1460 26954 1465
rect 27146 1495 27178 1500
rect 27146 1465 27149 1495
rect 27175 1465 27178 1495
rect 27146 1460 27178 1465
rect 27345 1495 27385 1500
rect 27345 1465 27350 1495
rect 27380 1465 27385 1495
rect 27345 1460 27385 1465
rect 27565 1495 27605 1500
rect 27565 1465 27570 1495
rect 27600 1465 27605 1495
rect 27565 1460 27605 1465
rect 26145 1435 26185 1440
rect 26145 1405 26150 1435
rect 26180 1405 26185 1435
rect 26145 1400 26185 1405
rect 26250 1435 26290 1440
rect 26250 1405 26255 1435
rect 26285 1405 26290 1435
rect 26250 1400 26290 1405
rect 26360 1435 26400 1440
rect 26360 1405 26365 1435
rect 26395 1405 26400 1435
rect 26360 1400 26400 1405
rect 26470 1435 26510 1440
rect 26470 1405 26475 1435
rect 26505 1405 26510 1435
rect 26470 1400 26510 1405
rect 26580 1435 26620 1440
rect 26580 1405 26585 1435
rect 26615 1405 26620 1435
rect 26580 1400 26620 1405
rect 12925 1390 12965 1395
rect 26830 1390 26850 1460
rect 12925 1360 12930 1390
rect 12960 1360 12965 1390
rect 12925 1355 12965 1360
rect 26810 1385 26850 1390
rect 26810 1355 26815 1385
rect 26845 1355 26850 1385
rect 26810 1350 26850 1355
rect 26315 1335 26355 1340
rect 26315 1305 26320 1335
rect 26350 1305 26355 1335
rect 26315 1300 26355 1305
rect 26325 1280 26345 1300
rect 26820 1280 26840 1350
rect 26880 1340 26900 1460
rect 27185 1435 27225 1440
rect 27185 1405 27190 1435
rect 27220 1405 27225 1435
rect 27185 1400 27225 1405
rect 27290 1435 27330 1440
rect 27290 1405 27295 1435
rect 27325 1405 27330 1435
rect 27290 1400 27330 1405
rect 27400 1435 27440 1440
rect 27400 1405 27405 1435
rect 27435 1405 27440 1435
rect 27400 1400 27440 1405
rect 27510 1435 27550 1440
rect 27510 1405 27515 1435
rect 27545 1405 27550 1435
rect 27510 1400 27550 1405
rect 27620 1435 27660 1440
rect 27620 1405 27625 1435
rect 27655 1405 27660 1435
rect 27620 1400 27660 1405
rect 28026 1350 28058 1355
rect 26880 1335 26920 1340
rect 26880 1305 26885 1335
rect 26915 1305 26920 1335
rect 28026 1320 28028 1350
rect 28054 1320 28058 1350
rect 28026 1315 28058 1320
rect 28292 1350 28324 1355
rect 28292 1320 28296 1350
rect 28322 1320 28324 1350
rect 28292 1315 28324 1320
rect 26880 1300 26920 1305
rect 27595 1290 27635 1295
rect 26315 1270 26355 1280
rect 26315 1250 26325 1270
rect 26345 1250 26355 1270
rect 26315 1240 26355 1250
rect 26425 1275 26465 1280
rect 26425 1245 26430 1275
rect 26460 1245 26465 1275
rect 26425 1240 26465 1245
rect 26535 1275 26575 1280
rect 26535 1245 26540 1275
rect 26570 1245 26575 1275
rect 26535 1240 26575 1245
rect 26645 1275 26685 1280
rect 26645 1245 26650 1275
rect 26680 1245 26685 1275
rect 26645 1240 26685 1245
rect 26755 1275 26795 1280
rect 26755 1245 26760 1275
rect 26790 1245 26795 1275
rect 26755 1240 26795 1245
rect 26815 1270 26845 1280
rect 26815 1250 26820 1270
rect 26840 1250 26845 1270
rect 26815 1240 26845 1250
rect 26865 1275 26905 1280
rect 26865 1245 26870 1275
rect 26900 1245 26905 1275
rect 26865 1240 26905 1245
rect 26975 1275 27015 1280
rect 26975 1245 26980 1275
rect 27010 1245 27015 1275
rect 26975 1240 27015 1245
rect 27085 1275 27125 1280
rect 27085 1245 27090 1275
rect 27120 1245 27125 1275
rect 27085 1240 27125 1245
rect 27195 1275 27235 1280
rect 27195 1245 27200 1275
rect 27230 1245 27235 1275
rect 27195 1240 27235 1245
rect 27305 1275 27345 1280
rect 27305 1245 27310 1275
rect 27340 1245 27345 1275
rect 27305 1240 27345 1245
rect 27415 1275 27455 1280
rect 27415 1245 27420 1275
rect 27450 1245 27455 1275
rect 27415 1240 27455 1245
rect 27525 1275 27565 1280
rect 27525 1245 27530 1275
rect 27560 1245 27565 1275
rect 27595 1260 27600 1290
rect 27630 1260 27635 1290
rect 27595 1255 27635 1260
rect 27945 1290 27985 1295
rect 27945 1260 27950 1290
rect 27980 1260 27985 1290
rect 27945 1255 27985 1260
rect 28060 1290 28100 1295
rect 28060 1260 28065 1290
rect 28095 1260 28100 1290
rect 28060 1255 28100 1260
rect 28155 1290 28195 1295
rect 28155 1260 28160 1290
rect 28190 1260 28195 1290
rect 28155 1255 28195 1260
rect 28250 1290 28290 1295
rect 28250 1260 28255 1290
rect 28285 1260 28290 1290
rect 28250 1255 28290 1260
rect 28365 1290 28405 1295
rect 28365 1260 28370 1290
rect 28400 1260 28405 1290
rect 28365 1255 28405 1260
rect 27525 1240 27565 1245
rect 28165 1235 28185 1255
rect 28375 1235 28395 1255
rect 28100 1230 28140 1235
rect 28100 1200 28105 1230
rect 28135 1200 28140 1230
rect 28100 1195 28140 1200
rect 28160 1230 28190 1235
rect 28160 1195 28190 1200
rect 28210 1230 28250 1235
rect 28210 1200 28215 1230
rect 28245 1200 28250 1230
rect 28210 1195 28250 1200
rect 28365 1230 28405 1235
rect 28365 1200 28370 1230
rect 28400 1200 28405 1230
rect 28365 1195 28405 1200
rect 26165 955 26205 960
rect 13205 935 13245 940
rect 13205 905 13210 935
rect 13240 905 13245 935
rect 13205 900 13245 905
rect 13405 935 13445 940
rect 13405 905 13410 935
rect 13440 905 13445 935
rect 26165 925 26170 955
rect 26200 925 26205 955
rect 26165 920 26205 925
rect 26260 955 26300 960
rect 26260 925 26265 955
rect 26295 925 26300 955
rect 26260 920 26300 925
rect 26370 955 26410 960
rect 26370 925 26375 955
rect 26405 925 26410 955
rect 26370 920 26410 925
rect 26480 955 26520 960
rect 26480 925 26485 955
rect 26515 925 26520 955
rect 26480 920 26520 925
rect 26590 955 26630 960
rect 26590 925 26595 955
rect 26625 925 26630 955
rect 26590 920 26630 925
rect 26700 955 26740 960
rect 26700 925 26705 955
rect 26735 925 26740 955
rect 26700 920 26740 925
rect 26810 955 26850 960
rect 26810 925 26815 955
rect 26845 925 26850 955
rect 26810 920 26850 925
rect 26920 955 26960 960
rect 26920 925 26925 955
rect 26955 925 26960 955
rect 26920 920 26960 925
rect 27030 955 27070 960
rect 27030 925 27035 955
rect 27065 925 27070 955
rect 27030 920 27070 925
rect 27140 955 27180 960
rect 27140 925 27145 955
rect 27175 925 27180 955
rect 27140 920 27180 925
rect 27250 955 27290 960
rect 27250 925 27255 955
rect 27285 925 27290 955
rect 27250 920 27290 925
rect 27360 955 27400 960
rect 27360 925 27365 955
rect 27395 925 27400 955
rect 27360 920 27400 925
rect 27470 955 27510 960
rect 27470 925 27475 955
rect 27505 925 27510 955
rect 27470 920 27510 925
rect 27620 955 27660 960
rect 27620 925 27625 955
rect 27655 925 27660 955
rect 27620 920 27660 925
rect 13405 900 13445 905
rect 12860 860 12900 865
rect 12860 830 12865 860
rect 12895 830 12900 860
rect 12860 825 12900 830
rect 10950 795 10990 800
rect 10950 765 10955 795
rect 10985 765 10990 795
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 730 2560 760
rect 2520 725 2560 730
rect 3130 760 3170 765
rect 3130 730 3135 760
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 730 3665 760
rect 3625 725 3665 730
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 760 4025 765
rect 3985 730 3990 760
rect 4020 730 4025 760
rect 3985 725 4025 730
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 760 4385 765
rect 4345 730 4350 760
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 730 4565 760
rect 4525 725 4565 730
rect 4705 760 4745 765
rect 4705 730 4710 760
rect 4740 730 4745 760
rect 4705 725 4745 730
rect 4885 760 4925 765
rect 10950 760 10990 765
rect 11305 795 11345 800
rect 11305 765 11310 795
rect 11340 765 11345 795
rect 11305 760 11345 765
rect 11375 795 11415 800
rect 11375 765 11380 795
rect 11410 765 11415 795
rect 11375 760 11415 765
rect 11445 795 11485 800
rect 11445 765 11450 795
rect 11480 765 11485 795
rect 11935 795 11975 805
rect 11935 775 11945 795
rect 11965 775 11975 795
rect 11935 765 11975 775
rect 12045 800 12085 805
rect 12045 770 12050 800
rect 12080 770 12085 800
rect 12045 765 12085 770
rect 12155 795 12195 805
rect 12155 775 12165 795
rect 12185 775 12195 795
rect 12155 765 12195 775
rect 12265 800 12305 805
rect 12265 770 12270 800
rect 12300 770 12305 800
rect 12265 765 12305 770
rect 12375 795 12415 805
rect 12375 775 12385 795
rect 12405 775 12415 795
rect 12375 765 12415 775
rect 12485 800 12525 805
rect 12485 770 12490 800
rect 12520 770 12525 800
rect 12485 765 12525 770
rect 12805 800 12845 805
rect 12805 770 12810 800
rect 12840 770 12845 800
rect 12805 765 12845 770
rect 11445 760 11485 765
rect 4885 730 4890 760
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3275 295 3295 725
rect 3455 710 3475 725
rect 3815 710 3835 725
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 675 3485 705
rect 3445 670 3485 675
rect 3805 705 3845 710
rect 3805 675 3810 705
rect 3840 675 3845 705
rect 3805 670 3845 675
rect 3815 295 3835 670
rect 3995 295 4015 725
rect 4175 710 4195 725
rect 4165 705 4205 710
rect 4165 675 4170 705
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 4715 295 4735 725
rect 11990 680 12030 685
rect 11990 650 11995 680
rect 12025 650 12030 680
rect 11990 645 12030 650
rect 12100 680 12140 685
rect 12100 650 12105 680
rect 12135 650 12140 680
rect 12100 645 12140 650
rect 12210 680 12250 685
rect 12210 650 12215 680
rect 12245 650 12250 680
rect 12210 645 12250 650
rect 12320 680 12360 685
rect 12320 650 12325 680
rect 12355 650 12360 680
rect 12320 645 12360 650
rect 12430 680 12470 685
rect 12430 650 12435 680
rect 12465 650 12470 680
rect 12430 645 12470 650
rect 11340 -1375 11380 -1370
rect 11340 -1405 11345 -1375
rect 11375 -1405 11380 -1375
rect 11340 -1410 11380 -1405
rect 11460 -1375 11500 -1370
rect 11460 -1405 11465 -1375
rect 11495 -1405 11500 -1375
rect 11460 -1410 11500 -1405
rect 11580 -1375 11620 -1370
rect 11580 -1405 11585 -1375
rect 11615 -1405 11620 -1375
rect 11580 -1410 11620 -1405
rect 11700 -1375 11740 -1370
rect 11700 -1405 11705 -1375
rect 11735 -1405 11740 -1375
rect 11700 -1410 11740 -1405
rect 11820 -1375 11860 -1370
rect 11820 -1405 11825 -1375
rect 11855 -1405 11860 -1375
rect 11820 -1410 11860 -1405
rect 11940 -1375 11980 -1370
rect 11940 -1405 11945 -1375
rect 11975 -1405 11980 -1375
rect 11940 -1410 11980 -1405
rect 12060 -1375 12100 -1370
rect 12060 -1405 12065 -1375
rect 12095 -1405 12100 -1375
rect 12060 -1410 12100 -1405
rect 12180 -1375 12220 -1370
rect 12180 -1405 12185 -1375
rect 12215 -1405 12220 -1375
rect 12180 -1410 12220 -1405
rect 12300 -1375 12340 -1370
rect 12300 -1405 12305 -1375
rect 12335 -1405 12340 -1375
rect 12300 -1410 12340 -1405
rect 12420 -1375 12460 -1370
rect 12420 -1405 12425 -1375
rect 12455 -1405 12460 -1375
rect 12420 -1410 12460 -1405
rect 10580 -1790 10620 -1785
rect 10580 -1820 10585 -1790
rect 10615 -1820 10620 -1790
rect 10580 -1825 10620 -1820
rect 10905 -1795 10940 -1785
rect 10905 -1815 10910 -1795
rect 10930 -1815 10940 -1795
rect 10905 -1825 10940 -1815
rect 10980 -1790 11015 -1785
rect 10980 -1820 10985 -1790
rect 10980 -1825 11015 -1820
rect 10910 -1840 10930 -1825
rect 10900 -1845 10940 -1840
rect 10900 -1875 10905 -1845
rect 10935 -1875 10940 -1845
rect 10900 -1880 10940 -1875
rect 10990 -2520 11010 -1825
rect 11280 -1850 11320 -1840
rect 11280 -1870 11290 -1850
rect 11310 -1870 11320 -1850
rect 11280 -1880 11320 -1870
rect 11400 -1850 11440 -1840
rect 11400 -1870 11410 -1850
rect 11430 -1870 11440 -1850
rect 11400 -1880 11440 -1870
rect 11520 -1850 11560 -1840
rect 11520 -1870 11530 -1850
rect 11550 -1870 11560 -1850
rect 11520 -1880 11560 -1870
rect 11640 -1850 11680 -1840
rect 11640 -1870 11650 -1850
rect 11670 -1870 11680 -1850
rect 11640 -1880 11680 -1870
rect 11760 -1850 11800 -1840
rect 11760 -1870 11770 -1850
rect 11790 -1870 11800 -1850
rect 11760 -1880 11800 -1870
rect 11823 -1845 11857 -1840
rect 11823 -1875 11826 -1845
rect 11854 -1875 11857 -1845
rect 11823 -1880 11857 -1875
rect 11880 -1850 11920 -1840
rect 11880 -1870 11890 -1850
rect 11910 -1870 11920 -1850
rect 11880 -1880 11920 -1870
rect 12000 -1850 12040 -1840
rect 12000 -1870 12010 -1850
rect 12030 -1870 12040 -1850
rect 12000 -1880 12040 -1870
rect 12120 -1850 12160 -1840
rect 12120 -1870 12130 -1850
rect 12150 -1870 12160 -1850
rect 12120 -1880 12160 -1870
rect 12240 -1850 12280 -1840
rect 12240 -1870 12250 -1850
rect 12270 -1870 12280 -1850
rect 12240 -1880 12280 -1870
rect 12360 -1850 12400 -1840
rect 12360 -1870 12370 -1850
rect 12390 -1870 12400 -1850
rect 12360 -1880 12400 -1870
rect 12480 -1850 12520 -1840
rect 12480 -1870 12490 -1850
rect 12510 -1870 12520 -1850
rect 12480 -1880 12520 -1870
rect 11290 -1895 11310 -1880
rect 11280 -1900 11320 -1895
rect 11280 -1930 11285 -1900
rect 11315 -1930 11320 -1900
rect 11280 -1935 11320 -1930
rect 11410 -1940 11430 -1880
rect 11530 -1895 11550 -1880
rect 11520 -1900 11560 -1895
rect 11520 -1930 11525 -1900
rect 11555 -1930 11560 -1900
rect 11520 -1935 11560 -1930
rect 11650 -1940 11670 -1880
rect 11770 -1895 11790 -1880
rect 11760 -1900 11800 -1895
rect 11760 -1930 11765 -1900
rect 11795 -1930 11800 -1900
rect 11760 -1935 11800 -1930
rect 11890 -1940 11910 -1880
rect 12010 -1895 12030 -1880
rect 12000 -1900 12040 -1895
rect 12000 -1930 12005 -1900
rect 12035 -1930 12040 -1900
rect 12000 -1935 12040 -1930
rect 12130 -1940 12150 -1880
rect 12250 -1895 12270 -1880
rect 12240 -1900 12280 -1895
rect 12240 -1930 12245 -1900
rect 12275 -1930 12280 -1900
rect 12240 -1935 12280 -1930
rect 12370 -1940 12390 -1880
rect 12490 -1895 12510 -1880
rect 12480 -1900 12520 -1895
rect 12480 -1930 12485 -1900
rect 12515 -1930 12520 -1900
rect 12480 -1935 12520 -1930
rect 11400 -1945 11440 -1940
rect 11400 -1975 11405 -1945
rect 11435 -1975 11440 -1945
rect 11400 -1980 11440 -1975
rect 11640 -1945 11680 -1940
rect 11640 -1975 11645 -1945
rect 11675 -1975 11680 -1945
rect 11640 -1980 11680 -1975
rect 11880 -1945 11920 -1940
rect 11880 -1975 11885 -1945
rect 11915 -1975 11920 -1945
rect 11880 -1980 11920 -1975
rect 12120 -1945 12160 -1940
rect 12120 -1975 12125 -1945
rect 12155 -1975 12160 -1945
rect 12120 -1980 12160 -1975
rect 12360 -1945 12400 -1940
rect 12360 -1975 12365 -1945
rect 12395 -1975 12400 -1945
rect 12360 -1980 12400 -1975
rect 11410 -1995 11430 -1980
rect 11340 -2000 11380 -1995
rect 11340 -2030 11345 -2000
rect 11375 -2030 11380 -2000
rect 11340 -2035 11380 -2030
rect 11400 -2000 11440 -1995
rect 11400 -2030 11405 -2000
rect 11435 -2030 11440 -2000
rect 11400 -2035 11440 -2030
rect 11580 -2000 11620 -1995
rect 11580 -2030 11585 -2000
rect 11615 -2030 11620 -2000
rect 11580 -2035 11620 -2030
rect 11820 -2000 11860 -1995
rect 11820 -2030 11825 -2000
rect 11855 -2030 11860 -2000
rect 11820 -2035 11860 -2030
rect 12060 -2000 12100 -1995
rect 12060 -2030 12065 -2000
rect 12095 -2030 12100 -2000
rect 12060 -2035 12100 -2030
rect 12300 -2000 12340 -1995
rect 12300 -2030 12305 -2000
rect 12335 -2030 12340 -2000
rect 12300 -2035 12340 -2030
rect 11350 -2050 11370 -2035
rect 11590 -2050 11610 -2035
rect 11830 -2050 11850 -2035
rect 12070 -2050 12090 -2035
rect 12310 -2050 12330 -2035
rect 12490 -2050 12510 -1935
rect 12950 -1965 12990 -1960
rect 12950 -1995 12955 -1965
rect 12985 -1995 12990 -1965
rect 12950 -2000 12990 -1995
rect 13060 -1965 13100 -1960
rect 13060 -1995 13065 -1965
rect 13095 -1995 13100 -1965
rect 13060 -2000 13100 -1995
rect 13170 -1965 13210 -1960
rect 13170 -1995 13175 -1965
rect 13205 -1995 13210 -1965
rect 13170 -2000 13210 -1995
rect 13280 -1965 13320 -1960
rect 13280 -1995 13285 -1965
rect 13315 -1995 13320 -1965
rect 13280 -2000 13320 -1995
rect 13390 -1965 13430 -1960
rect 13390 -1995 13395 -1965
rect 13425 -1995 13430 -1965
rect 13390 -2000 13430 -1995
rect 13500 -1965 13540 -1960
rect 13500 -1995 13505 -1965
rect 13535 -1995 13540 -1965
rect 13500 -2000 13540 -1995
rect 13610 -1965 13650 -1960
rect 13610 -1995 13615 -1965
rect 13645 -1995 13650 -1965
rect 13610 -2000 13650 -1995
rect 13720 -1965 13760 -1960
rect 13720 -1995 13725 -1965
rect 13755 -1995 13760 -1965
rect 13720 -2000 13760 -1995
rect 13830 -1965 13870 -1960
rect 13830 -1995 13835 -1965
rect 13865 -1995 13870 -1965
rect 13830 -2000 13870 -1995
rect 13940 -1965 13980 -1960
rect 13940 -1995 13945 -1965
rect 13975 -1995 13980 -1965
rect 13940 -2000 13980 -1995
rect 14050 -1965 14090 -1960
rect 14050 -1995 14055 -1965
rect 14085 -1995 14090 -1965
rect 14050 -2000 14090 -1995
rect 11340 -2060 11380 -2050
rect 11340 -2080 11350 -2060
rect 11370 -2080 11380 -2060
rect 11340 -2090 11380 -2080
rect 11460 -2055 11500 -2050
rect 11460 -2085 11465 -2055
rect 11495 -2085 11500 -2055
rect 11460 -2090 11500 -2085
rect 11580 -2060 11620 -2050
rect 11580 -2080 11590 -2060
rect 11610 -2080 11620 -2060
rect 11580 -2090 11620 -2080
rect 11700 -2055 11740 -2050
rect 11700 -2085 11705 -2055
rect 11735 -2085 11740 -2055
rect 11700 -2090 11740 -2085
rect 11820 -2060 11860 -2050
rect 11820 -2080 11830 -2060
rect 11850 -2080 11860 -2060
rect 11820 -2090 11860 -2080
rect 11940 -2055 11980 -2050
rect 11940 -2085 11945 -2055
rect 11975 -2085 11980 -2055
rect 11940 -2090 11980 -2085
rect 12060 -2060 12100 -2050
rect 12060 -2080 12070 -2060
rect 12090 -2080 12100 -2060
rect 12060 -2090 12100 -2080
rect 12180 -2055 12220 -2050
rect 12180 -2085 12185 -2055
rect 12215 -2085 12220 -2055
rect 12180 -2090 12220 -2085
rect 12300 -2060 12340 -2050
rect 12300 -2080 12310 -2060
rect 12330 -2080 12340 -2060
rect 12300 -2090 12340 -2080
rect 12420 -2055 12460 -2050
rect 12420 -2085 12425 -2055
rect 12455 -2085 12460 -2055
rect 12420 -2090 12460 -2085
rect 12480 -2055 12520 -2050
rect 12480 -2085 12485 -2055
rect 12515 -2085 12520 -2055
rect 12480 -2090 12520 -2085
rect 12690 -2270 12730 -2265
rect 12690 -2300 12695 -2270
rect 12725 -2300 12730 -2270
rect 12690 -2305 12730 -2300
rect 10980 -2525 11020 -2520
rect 10980 -2555 10985 -2525
rect 11015 -2555 11020 -2525
rect 10980 -2560 11020 -2555
rect 11280 -2530 11320 -2520
rect 11280 -2550 11290 -2530
rect 11310 -2550 11320 -2530
rect 11280 -2560 11320 -2550
rect 11400 -2530 11440 -2520
rect 11400 -2550 11410 -2530
rect 11430 -2550 11440 -2530
rect 11400 -2560 11440 -2550
rect 11520 -2530 11560 -2520
rect 11520 -2550 11530 -2530
rect 11550 -2550 11560 -2530
rect 11520 -2560 11560 -2550
rect 11640 -2530 11680 -2520
rect 11640 -2550 11650 -2530
rect 11670 -2550 11680 -2530
rect 11640 -2560 11680 -2550
rect 11760 -2530 11800 -2520
rect 11760 -2550 11770 -2530
rect 11790 -2550 11800 -2530
rect 11760 -2560 11800 -2550
rect 11823 -2525 11857 -2520
rect 11823 -2555 11826 -2525
rect 11854 -2555 11857 -2525
rect 11823 -2560 11857 -2555
rect 11880 -2530 11920 -2520
rect 11880 -2550 11890 -2530
rect 11910 -2550 11920 -2530
rect 11880 -2560 11920 -2550
rect 12000 -2530 12040 -2520
rect 12000 -2550 12010 -2530
rect 12030 -2550 12040 -2530
rect 12000 -2560 12040 -2550
rect 12120 -2530 12160 -2520
rect 12120 -2550 12130 -2530
rect 12150 -2550 12160 -2530
rect 12120 -2560 12160 -2550
rect 12240 -2530 12280 -2520
rect 12240 -2550 12250 -2530
rect 12270 -2550 12280 -2530
rect 12240 -2560 12280 -2550
rect 12360 -2530 12400 -2520
rect 12360 -2550 12370 -2530
rect 12390 -2550 12400 -2530
rect 12360 -2560 12400 -2550
rect 12480 -2530 12520 -2520
rect 12480 -2550 12490 -2530
rect 12510 -2550 12520 -2530
rect 12480 -2560 12520 -2550
rect 11290 -2575 11310 -2560
rect 11280 -2580 11320 -2575
rect 11280 -2610 11285 -2580
rect 11315 -2610 11320 -2580
rect 11280 -2615 11320 -2610
rect 11410 -2620 11430 -2560
rect 11530 -2575 11550 -2560
rect 11520 -2580 11560 -2575
rect 11520 -2610 11525 -2580
rect 11555 -2610 11560 -2580
rect 11520 -2615 11560 -2610
rect 11650 -2620 11670 -2560
rect 11770 -2575 11790 -2560
rect 11760 -2580 11800 -2575
rect 11760 -2610 11765 -2580
rect 11795 -2610 11800 -2580
rect 11760 -2615 11800 -2610
rect 11400 -2625 11440 -2620
rect 11400 -2655 11405 -2625
rect 11435 -2655 11440 -2625
rect 11400 -2660 11440 -2655
rect 11640 -2625 11680 -2620
rect 11640 -2655 11645 -2625
rect 11675 -2655 11680 -2625
rect 11640 -2660 11680 -2655
rect 11440 -2720 11480 -2715
rect 11440 -2750 11445 -2720
rect 11475 -2750 11480 -2720
rect 11440 -2755 11480 -2750
rect 11660 -2720 11700 -2715
rect 11660 -2750 11665 -2720
rect 11695 -2750 11700 -2720
rect 11660 -2755 11700 -2750
rect 11330 -2765 11370 -2760
rect 11330 -2795 11335 -2765
rect 11365 -2795 11370 -2765
rect 11330 -2800 11370 -2795
rect 11340 -2815 11360 -2800
rect 11450 -2815 11470 -2755
rect 11550 -2765 11590 -2760
rect 11550 -2795 11555 -2765
rect 11585 -2795 11590 -2765
rect 11550 -2800 11590 -2795
rect 11560 -2815 11580 -2800
rect 11670 -2815 11690 -2755
rect 11770 -2760 11790 -2615
rect 11890 -2620 11910 -2560
rect 12010 -2575 12030 -2560
rect 12000 -2580 12040 -2575
rect 12000 -2610 12005 -2580
rect 12035 -2610 12040 -2580
rect 12000 -2615 12040 -2610
rect 12130 -2620 12150 -2560
rect 12250 -2575 12270 -2560
rect 12240 -2580 12280 -2575
rect 12240 -2610 12245 -2580
rect 12275 -2610 12280 -2580
rect 12240 -2615 12280 -2610
rect 12370 -2620 12390 -2560
rect 12490 -2575 12510 -2560
rect 12480 -2580 12520 -2575
rect 12480 -2610 12485 -2580
rect 12515 -2610 12520 -2580
rect 12480 -2615 12520 -2610
rect 12700 -2620 12720 -2305
rect 13005 -2335 13045 -2330
rect 13005 -2365 13010 -2335
rect 13040 -2365 13045 -2335
rect 13005 -2370 13045 -2365
rect 13063 -2340 13097 -2330
rect 13063 -2360 13071 -2340
rect 13089 -2360 13097 -2340
rect 13063 -2370 13097 -2360
rect 13115 -2335 13155 -2330
rect 13115 -2365 13120 -2335
rect 13150 -2365 13155 -2335
rect 13115 -2370 13155 -2365
rect 13225 -2335 13265 -2330
rect 13225 -2365 13230 -2335
rect 13260 -2365 13265 -2335
rect 13225 -2370 13265 -2365
rect 13335 -2335 13375 -2330
rect 13335 -2365 13340 -2335
rect 13370 -2365 13375 -2335
rect 13335 -2370 13375 -2365
rect 13445 -2335 13485 -2330
rect 13445 -2365 13450 -2335
rect 13480 -2365 13485 -2335
rect 13445 -2370 13485 -2365
rect 13555 -2335 13595 -2330
rect 13555 -2365 13560 -2335
rect 13590 -2365 13595 -2335
rect 13555 -2370 13595 -2365
rect 13665 -2335 13705 -2330
rect 13665 -2365 13670 -2335
rect 13700 -2365 13705 -2335
rect 13665 -2370 13705 -2365
rect 13775 -2335 13815 -2330
rect 13775 -2365 13780 -2335
rect 13810 -2365 13815 -2335
rect 13775 -2370 13815 -2365
rect 13885 -2335 13925 -2330
rect 13885 -2365 13890 -2335
rect 13920 -2365 13925 -2335
rect 13885 -2370 13925 -2365
rect 13995 -2335 14035 -2330
rect 13995 -2365 14000 -2335
rect 14030 -2365 14035 -2335
rect 13995 -2370 14035 -2365
rect 12950 -2395 12990 -2390
rect 12950 -2425 12955 -2395
rect 12985 -2425 12990 -2395
rect 12950 -2430 12990 -2425
rect 13060 -2395 13100 -2390
rect 13060 -2425 13065 -2395
rect 13095 -2425 13100 -2395
rect 13060 -2430 13100 -2425
rect 13170 -2395 13210 -2390
rect 13170 -2425 13175 -2395
rect 13205 -2425 13210 -2395
rect 13170 -2430 13210 -2425
rect 13280 -2395 13320 -2390
rect 13280 -2425 13285 -2395
rect 13315 -2425 13320 -2395
rect 13280 -2430 13320 -2425
rect 13390 -2395 13430 -2390
rect 13390 -2425 13395 -2395
rect 13425 -2425 13430 -2395
rect 13390 -2430 13430 -2425
rect 13500 -2395 13540 -2390
rect 13500 -2425 13505 -2395
rect 13535 -2425 13540 -2395
rect 13500 -2430 13540 -2425
rect 13610 -2395 13650 -2390
rect 13610 -2425 13615 -2395
rect 13645 -2425 13650 -2395
rect 13610 -2430 13650 -2425
rect 13720 -2395 13760 -2390
rect 13720 -2425 13725 -2395
rect 13755 -2425 13760 -2395
rect 13720 -2430 13760 -2425
rect 13830 -2395 13870 -2390
rect 13830 -2425 13835 -2395
rect 13865 -2425 13870 -2395
rect 13830 -2430 13870 -2425
rect 13940 -2395 13980 -2390
rect 13940 -2425 13945 -2395
rect 13975 -2425 13980 -2395
rect 13940 -2430 13980 -2425
rect 14050 -2395 14090 -2390
rect 14050 -2425 14055 -2395
rect 14085 -2425 14090 -2395
rect 14050 -2430 14090 -2425
rect 13005 -2565 13045 -2560
rect 13005 -2595 13010 -2565
rect 13040 -2595 13045 -2565
rect 13005 -2600 13045 -2595
rect 13115 -2565 13155 -2560
rect 13115 -2595 13120 -2565
rect 13150 -2595 13155 -2565
rect 13115 -2600 13155 -2595
rect 13225 -2565 13265 -2560
rect 13225 -2595 13230 -2565
rect 13260 -2595 13265 -2565
rect 13225 -2600 13265 -2595
rect 13335 -2565 13375 -2560
rect 13335 -2595 13340 -2565
rect 13370 -2595 13375 -2565
rect 13335 -2600 13375 -2595
rect 13445 -2565 13485 -2560
rect 13445 -2595 13450 -2565
rect 13480 -2595 13485 -2565
rect 13445 -2600 13485 -2595
rect 13555 -2565 13595 -2560
rect 13555 -2595 13560 -2565
rect 13590 -2595 13595 -2565
rect 13555 -2600 13595 -2595
rect 13665 -2565 13705 -2560
rect 13665 -2595 13670 -2565
rect 13700 -2595 13705 -2565
rect 13665 -2600 13705 -2595
rect 13775 -2565 13815 -2560
rect 13775 -2595 13780 -2565
rect 13810 -2595 13815 -2565
rect 13775 -2600 13815 -2595
rect 13885 -2565 13925 -2560
rect 13885 -2595 13890 -2565
rect 13920 -2595 13925 -2565
rect 13885 -2600 13925 -2595
rect 13995 -2565 14035 -2560
rect 13995 -2595 14000 -2565
rect 14030 -2595 14035 -2565
rect 13995 -2600 14035 -2595
rect 11880 -2625 11920 -2620
rect 11880 -2655 11885 -2625
rect 11915 -2655 11920 -2625
rect 11880 -2660 11920 -2655
rect 12120 -2625 12160 -2620
rect 12120 -2655 12125 -2625
rect 12155 -2655 12160 -2625
rect 12120 -2660 12160 -2655
rect 12360 -2625 12400 -2620
rect 12360 -2655 12365 -2625
rect 12395 -2655 12400 -2625
rect 12360 -2660 12400 -2655
rect 12690 -2625 12730 -2620
rect 12690 -2655 12695 -2625
rect 12725 -2655 12730 -2625
rect 12690 -2660 12730 -2655
rect 12975 -2625 13015 -2620
rect 12975 -2655 12980 -2625
rect 13010 -2655 13015 -2625
rect 12975 -2660 13015 -2655
rect 12120 -2715 12140 -2660
rect 13005 -2685 13045 -2680
rect 13005 -2715 13010 -2685
rect 13040 -2715 13045 -2685
rect 11880 -2720 11920 -2715
rect 11880 -2750 11885 -2720
rect 11915 -2750 11920 -2720
rect 11880 -2755 11920 -2750
rect 12100 -2720 12140 -2715
rect 12100 -2750 12105 -2720
rect 12135 -2750 12140 -2720
rect 12100 -2755 12140 -2750
rect 12320 -2720 12360 -2715
rect 13005 -2720 13045 -2715
rect 13115 -2685 13155 -2680
rect 13115 -2715 13120 -2685
rect 13150 -2715 13155 -2685
rect 13115 -2720 13155 -2715
rect 13225 -2685 13265 -2680
rect 13225 -2715 13230 -2685
rect 13260 -2715 13265 -2685
rect 13225 -2720 13265 -2715
rect 13335 -2685 13375 -2680
rect 13335 -2715 13340 -2685
rect 13370 -2715 13375 -2685
rect 13335 -2720 13375 -2715
rect 13445 -2685 13485 -2680
rect 13445 -2715 13450 -2685
rect 13480 -2715 13485 -2685
rect 13445 -2720 13485 -2715
rect 13555 -2685 13595 -2680
rect 13555 -2715 13560 -2685
rect 13590 -2715 13595 -2685
rect 13555 -2720 13595 -2715
rect 13665 -2685 13705 -2680
rect 13665 -2715 13670 -2685
rect 13700 -2715 13705 -2685
rect 13665 -2720 13705 -2715
rect 13775 -2685 13815 -2680
rect 13775 -2715 13780 -2685
rect 13810 -2715 13815 -2685
rect 13775 -2720 13815 -2715
rect 13885 -2685 13925 -2680
rect 13885 -2715 13890 -2685
rect 13920 -2715 13925 -2685
rect 13885 -2720 13925 -2715
rect 13995 -2685 14035 -2680
rect 13995 -2715 14000 -2685
rect 14030 -2715 14035 -2685
rect 13995 -2720 14035 -2715
rect 12320 -2750 12325 -2720
rect 12355 -2750 12360 -2720
rect 12320 -2755 12360 -2750
rect 11770 -2765 11810 -2760
rect 11770 -2795 11775 -2765
rect 11805 -2795 11810 -2765
rect 11770 -2800 11810 -2795
rect 11780 -2815 11800 -2800
rect 11890 -2815 11910 -2755
rect 11990 -2765 12030 -2760
rect 11990 -2795 11995 -2765
rect 12025 -2795 12030 -2765
rect 11990 -2800 12030 -2795
rect 12000 -2815 12020 -2800
rect 12110 -2815 12130 -2755
rect 12210 -2765 12250 -2760
rect 12210 -2795 12215 -2765
rect 12245 -2795 12250 -2765
rect 12210 -2800 12250 -2795
rect 12220 -2815 12240 -2800
rect 12330 -2815 12350 -2755
rect 12430 -2765 12470 -2760
rect 12430 -2795 12435 -2765
rect 12465 -2795 12470 -2765
rect 12430 -2800 12470 -2795
rect 12440 -2815 12460 -2800
rect 11330 -2825 11370 -2815
rect 11330 -2845 11340 -2825
rect 11360 -2845 11370 -2825
rect 11330 -2855 11370 -2845
rect 11440 -2825 11480 -2815
rect 11440 -2845 11450 -2825
rect 11470 -2845 11480 -2825
rect 11440 -2855 11480 -2845
rect 11550 -2825 11590 -2815
rect 11550 -2845 11560 -2825
rect 11580 -2845 11590 -2825
rect 11550 -2855 11590 -2845
rect 11660 -2825 11700 -2815
rect 11660 -2845 11670 -2825
rect 11690 -2845 11700 -2825
rect 11660 -2855 11700 -2845
rect 11770 -2825 11810 -2815
rect 11770 -2845 11780 -2825
rect 11800 -2845 11810 -2825
rect 11770 -2855 11810 -2845
rect 11880 -2825 11920 -2815
rect 11880 -2845 11890 -2825
rect 11910 -2845 11920 -2825
rect 11880 -2855 11920 -2845
rect 11990 -2825 12030 -2815
rect 11990 -2845 12000 -2825
rect 12020 -2845 12030 -2825
rect 11990 -2855 12030 -2845
rect 12100 -2825 12140 -2815
rect 12100 -2845 12110 -2825
rect 12130 -2845 12140 -2825
rect 12100 -2855 12140 -2845
rect 12210 -2825 12250 -2815
rect 12210 -2845 12220 -2825
rect 12240 -2845 12250 -2825
rect 12210 -2855 12250 -2845
rect 12320 -2825 12360 -2815
rect 12320 -2845 12330 -2825
rect 12350 -2845 12360 -2825
rect 12320 -2855 12360 -2845
rect 12430 -2825 12470 -2815
rect 12430 -2845 12440 -2825
rect 12460 -2845 12470 -2825
rect 12430 -2855 12470 -2845
rect 12950 -2905 12990 -2900
rect 12950 -2935 12955 -2905
rect 12985 -2935 12990 -2905
rect 12950 -2940 12990 -2935
rect 13060 -2905 13100 -2900
rect 13060 -2935 13065 -2905
rect 13095 -2935 13100 -2905
rect 13060 -2940 13100 -2935
rect 13170 -2905 13210 -2900
rect 13170 -2935 13175 -2905
rect 13205 -2935 13210 -2905
rect 13170 -2940 13210 -2935
rect 13280 -2905 13320 -2900
rect 13280 -2935 13285 -2905
rect 13315 -2935 13320 -2905
rect 13280 -2940 13320 -2935
rect 13390 -2905 13430 -2900
rect 13390 -2935 13395 -2905
rect 13425 -2935 13430 -2905
rect 13390 -2940 13430 -2935
rect 13500 -2905 13540 -2900
rect 13500 -2935 13505 -2905
rect 13535 -2935 13540 -2905
rect 13500 -2940 13540 -2935
rect 13610 -2905 13650 -2900
rect 13610 -2935 13615 -2905
rect 13645 -2935 13650 -2905
rect 13610 -2940 13650 -2935
rect 13720 -2905 13760 -2900
rect 13720 -2935 13725 -2905
rect 13755 -2935 13760 -2905
rect 13720 -2940 13760 -2935
rect 13830 -2905 13870 -2900
rect 13830 -2935 13835 -2905
rect 13865 -2935 13870 -2905
rect 13830 -2940 13870 -2935
rect 13940 -2905 13980 -2900
rect 13940 -2935 13945 -2905
rect 13975 -2935 13980 -2905
rect 13940 -2940 13980 -2935
rect 14050 -2905 14090 -2900
rect 14050 -2935 14055 -2905
rect 14085 -2935 14090 -2905
rect 14050 -2940 14090 -2935
rect 12995 -2965 13035 -2960
rect 12995 -2995 13000 -2965
rect 13030 -2995 13035 -2965
rect 12995 -3000 13035 -2995
rect 13098 -2970 13132 -2960
rect 13098 -2990 13106 -2970
rect 13124 -2990 13132 -2970
rect 13098 -3000 13132 -2990
rect 13195 -2965 13235 -2960
rect 13195 -2995 13200 -2965
rect 13230 -2995 13235 -2965
rect 13195 -3000 13235 -2995
rect 13395 -2965 13435 -2960
rect 13395 -2995 13400 -2965
rect 13430 -2995 13435 -2965
rect 13395 -3000 13435 -2995
rect 13595 -2965 13635 -2960
rect 13595 -2995 13600 -2965
rect 13630 -2995 13635 -2965
rect 13595 -3000 13635 -2995
rect 13795 -2965 13835 -2960
rect 13795 -2995 13800 -2965
rect 13830 -2995 13835 -2965
rect 13795 -3000 13835 -2995
rect 13995 -2965 14035 -2960
rect 13995 -2995 14000 -2965
rect 14030 -2995 14035 -2965
rect 13995 -3000 14035 -2995
rect 11385 -3040 11425 -3035
rect 11385 -3070 11390 -3040
rect 11420 -3070 11425 -3040
rect 11385 -3075 11425 -3070
rect 11495 -3045 11535 -3035
rect 11495 -3065 11505 -3045
rect 11525 -3065 11535 -3045
rect 11495 -3075 11535 -3065
rect 11605 -3040 11645 -3035
rect 11605 -3070 11610 -3040
rect 11640 -3070 11645 -3040
rect 11605 -3075 11645 -3070
rect 11715 -3045 11755 -3035
rect 11715 -3065 11725 -3045
rect 11745 -3065 11755 -3045
rect 11715 -3075 11755 -3065
rect 11825 -3040 11865 -3035
rect 11825 -3070 11830 -3040
rect 11860 -3070 11865 -3040
rect 11825 -3075 11865 -3070
rect 11935 -3045 11975 -3035
rect 11935 -3065 11945 -3045
rect 11965 -3065 11975 -3045
rect 11935 -3075 11975 -3065
rect 12045 -3040 12085 -3035
rect 12045 -3070 12050 -3040
rect 12080 -3070 12085 -3040
rect 12045 -3075 12085 -3070
rect 12155 -3045 12195 -3035
rect 12155 -3065 12165 -3045
rect 12185 -3065 12195 -3045
rect 12155 -3075 12195 -3065
rect 12245 -3040 12305 -3035
rect 12245 -3070 12270 -3040
rect 12300 -3070 12305 -3040
rect 12245 -3075 12305 -3070
rect 12375 -3045 12415 -3035
rect 12375 -3065 12385 -3045
rect 12405 -3065 12415 -3045
rect 12375 -3075 12415 -3065
rect 11505 -3090 11525 -3075
rect 11725 -3090 11745 -3075
rect 11945 -3090 11965 -3075
rect 12165 -3090 12185 -3075
rect 11495 -3095 11555 -3090
rect 11495 -3125 11500 -3095
rect 11530 -3125 11555 -3095
rect 11495 -3130 11555 -3125
rect 11715 -3095 11755 -3090
rect 11715 -3125 11720 -3095
rect 11750 -3125 11755 -3095
rect 11715 -3130 11755 -3125
rect 11935 -3095 11975 -3090
rect 11935 -3125 11940 -3095
rect 11970 -3125 11975 -3095
rect 11935 -3130 11975 -3125
rect 12155 -3095 12195 -3090
rect 12155 -3125 12160 -3095
rect 12190 -3125 12195 -3095
rect 12155 -3130 12195 -3125
rect 11190 -3150 11230 -3145
rect 11190 -3180 11195 -3150
rect 11225 -3180 11230 -3150
rect 11190 -3185 11230 -3180
rect 11410 -3150 11450 -3145
rect 11410 -3180 11415 -3150
rect 11445 -3180 11450 -3150
rect 11410 -3185 11450 -3180
rect 11200 -3220 11220 -3185
rect 11420 -3220 11440 -3185
rect 11190 -3230 11230 -3220
rect 11085 -3240 11125 -3235
rect 11085 -3270 11090 -3240
rect 11120 -3270 11125 -3240
rect 11190 -3250 11200 -3230
rect 11220 -3250 11230 -3230
rect 11410 -3230 11450 -3220
rect 11190 -3260 11230 -3250
rect 11305 -3240 11345 -3235
rect 11085 -3275 11125 -3270
rect 11305 -3270 11310 -3240
rect 11340 -3270 11345 -3240
rect 11410 -3250 11420 -3230
rect 11440 -3250 11450 -3230
rect 11535 -3235 11555 -3130
rect 12245 -3145 12265 -3075
rect 12385 -3090 12405 -3075
rect 12375 -3095 12415 -3090
rect 12375 -3125 12380 -3095
rect 12410 -3125 12415 -3095
rect 12375 -3130 12415 -3125
rect 11640 -3150 11680 -3145
rect 11640 -3180 11645 -3150
rect 11675 -3180 11680 -3150
rect 11640 -3185 11680 -3180
rect 12230 -3150 12270 -3145
rect 12230 -3180 12235 -3150
rect 12265 -3180 12270 -3150
rect 12230 -3185 12270 -3180
rect 12450 -3150 12490 -3145
rect 12450 -3180 12455 -3150
rect 12485 -3180 12490 -3150
rect 12450 -3185 12490 -3180
rect 12680 -3150 12720 -3145
rect 12680 -3180 12685 -3150
rect 12715 -3180 12720 -3150
rect 12680 -3185 12720 -3180
rect 11650 -3220 11670 -3185
rect 11820 -3195 11860 -3190
rect 11640 -3230 11680 -3220
rect 11820 -3225 11825 -3195
rect 11855 -3225 11860 -3195
rect 11820 -3230 11860 -3225
rect 11940 -3195 11980 -3190
rect 11940 -3225 11945 -3195
rect 11975 -3225 11980 -3195
rect 12240 -3220 12260 -3185
rect 12460 -3220 12480 -3185
rect 12690 -3220 12710 -3185
rect 11940 -3230 11980 -3225
rect 12230 -3230 12270 -3220
rect 11410 -3260 11450 -3250
rect 11525 -3240 11565 -3235
rect 11305 -3275 11345 -3270
rect 11525 -3270 11530 -3240
rect 11560 -3270 11565 -3240
rect 11640 -3250 11650 -3230
rect 11670 -3250 11680 -3230
rect 11640 -3260 11680 -3250
rect 11525 -3275 11565 -3270
rect 11830 -3280 11850 -3230
rect 11950 -3280 11970 -3230
rect 12125 -3240 12165 -3235
rect 12125 -3270 12130 -3240
rect 12160 -3270 12165 -3240
rect 12230 -3250 12240 -3230
rect 12260 -3250 12270 -3230
rect 12450 -3230 12490 -3220
rect 12230 -3260 12270 -3250
rect 12345 -3240 12385 -3235
rect 12125 -3275 12165 -3270
rect 12345 -3270 12350 -3240
rect 12380 -3270 12385 -3240
rect 12450 -3250 12460 -3230
rect 12480 -3250 12490 -3230
rect 12680 -3230 12720 -3220
rect 12450 -3260 12490 -3250
rect 12565 -3240 12605 -3235
rect 12345 -3275 12385 -3270
rect 12565 -3270 12570 -3240
rect 12600 -3270 12605 -3240
rect 12680 -3250 12690 -3230
rect 12710 -3250 12720 -3230
rect 12680 -3260 12720 -3250
rect 12565 -3275 12605 -3270
rect 11237 -3285 11269 -3280
rect 11237 -3315 11240 -3285
rect 11266 -3315 11269 -3285
rect 11237 -3320 11269 -3315
rect 11457 -3285 11489 -3280
rect 11457 -3315 11460 -3285
rect 11486 -3315 11489 -3285
rect 11457 -3320 11489 -3315
rect 11601 -3285 11633 -3280
rect 11601 -3315 11604 -3285
rect 11630 -3315 11633 -3285
rect 11601 -3320 11633 -3315
rect 11820 -3290 11850 -3280
rect 11820 -3310 11825 -3290
rect 11845 -3310 11850 -3290
rect 11820 -3320 11850 -3310
rect 11867 -3285 11899 -3280
rect 11867 -3315 11870 -3285
rect 11896 -3315 11899 -3285
rect 11867 -3320 11899 -3315
rect 11950 -3290 11980 -3280
rect 11950 -3310 11955 -3290
rect 11975 -3310 11980 -3290
rect 11950 -3320 11980 -3310
rect 12277 -3285 12309 -3280
rect 12277 -3315 12280 -3285
rect 12306 -3315 12309 -3285
rect 12277 -3320 12309 -3315
rect 12497 -3285 12529 -3280
rect 12497 -3315 12500 -3285
rect 12526 -3315 12529 -3285
rect 12497 -3320 12529 -3315
rect 12641 -3285 12673 -3280
rect 12641 -3315 12644 -3285
rect 12670 -3315 12673 -3285
rect 12641 -3320 12673 -3315
rect 13095 -3315 13135 -3310
rect 13095 -3345 13100 -3315
rect 13130 -3345 13135 -3315
rect 13095 -3350 13135 -3345
rect 13295 -3315 13335 -3310
rect 13295 -3345 13300 -3315
rect 13330 -3345 13335 -3315
rect 13295 -3350 13335 -3345
rect 13495 -3315 13535 -3310
rect 13495 -3345 13500 -3315
rect 13530 -3345 13535 -3315
rect 13495 -3350 13535 -3345
rect 13695 -3315 13735 -3310
rect 13695 -3345 13700 -3315
rect 13730 -3345 13735 -3315
rect 13695 -3350 13735 -3345
rect 13895 -3315 13935 -3310
rect 13895 -3345 13900 -3315
rect 13930 -3345 13935 -3315
rect 13895 -3350 13935 -3345
rect 11106 -3505 11138 -3500
rect 11106 -3535 11109 -3505
rect 11135 -3535 11138 -3505
rect 11106 -3540 11138 -3535
rect 11305 -3505 11345 -3500
rect 11305 -3535 11310 -3505
rect 11340 -3535 11345 -3505
rect 11305 -3540 11345 -3535
rect 11525 -3505 11565 -3500
rect 11525 -3535 11530 -3505
rect 11560 -3535 11565 -3505
rect 11525 -3540 11565 -3535
rect 11825 -3510 11855 -3500
rect 11825 -3530 11830 -3510
rect 11850 -3530 11855 -3510
rect 11825 -3540 11855 -3530
rect 11875 -3510 11905 -3500
rect 11875 -3530 11880 -3510
rect 11900 -3530 11905 -3510
rect 11875 -3540 11905 -3530
rect 11922 -3505 11954 -3500
rect 11922 -3535 11925 -3505
rect 11951 -3535 11954 -3505
rect 11922 -3540 11954 -3535
rect 12146 -3505 12178 -3500
rect 12146 -3535 12149 -3505
rect 12175 -3535 12178 -3505
rect 12146 -3540 12178 -3535
rect 12345 -3505 12385 -3500
rect 12345 -3535 12350 -3505
rect 12380 -3535 12385 -3505
rect 12345 -3540 12385 -3535
rect 12565 -3505 12605 -3500
rect 12565 -3535 12570 -3505
rect 12600 -3535 12605 -3505
rect 12565 -3540 12605 -3535
rect 11145 -3565 11185 -3560
rect 11145 -3595 11150 -3565
rect 11180 -3595 11185 -3565
rect 11145 -3600 11185 -3595
rect 11250 -3565 11290 -3560
rect 11250 -3595 11255 -3565
rect 11285 -3595 11290 -3565
rect 11250 -3600 11290 -3595
rect 11360 -3565 11400 -3560
rect 11360 -3595 11365 -3565
rect 11395 -3595 11400 -3565
rect 11360 -3600 11400 -3595
rect 11470 -3565 11510 -3560
rect 11470 -3595 11475 -3565
rect 11505 -3595 11510 -3565
rect 11470 -3600 11510 -3595
rect 11580 -3565 11620 -3560
rect 11580 -3595 11585 -3565
rect 11615 -3595 11620 -3565
rect 11580 -3600 11620 -3595
rect 11830 -3650 11850 -3540
rect 11810 -3655 11850 -3650
rect 11810 -3685 11815 -3655
rect 11845 -3685 11850 -3655
rect 11810 -3690 11850 -3685
rect 11315 -3705 11355 -3700
rect 11315 -3735 11320 -3705
rect 11350 -3735 11355 -3705
rect 11315 -3740 11355 -3735
rect 11325 -3760 11345 -3740
rect 11820 -3760 11840 -3690
rect 11880 -3700 11900 -3540
rect 12185 -3565 12225 -3560
rect 12185 -3595 12190 -3565
rect 12220 -3595 12225 -3565
rect 12185 -3600 12225 -3595
rect 12290 -3565 12330 -3560
rect 12290 -3595 12295 -3565
rect 12325 -3595 12330 -3565
rect 12290 -3600 12330 -3595
rect 12400 -3565 12440 -3560
rect 12400 -3595 12405 -3565
rect 12435 -3595 12440 -3565
rect 12400 -3600 12440 -3595
rect 12510 -3565 12550 -3560
rect 12510 -3595 12515 -3565
rect 12545 -3595 12550 -3565
rect 12510 -3600 12550 -3595
rect 12620 -3565 12660 -3560
rect 12620 -3595 12625 -3565
rect 12655 -3595 12660 -3565
rect 12620 -3600 12660 -3595
rect 11880 -3705 11920 -3700
rect 11880 -3735 11885 -3705
rect 11915 -3735 11920 -3705
rect 11880 -3740 11920 -3735
rect 12595 -3750 12635 -3745
rect 11315 -3770 11355 -3760
rect 11315 -3790 11325 -3770
rect 11345 -3790 11355 -3770
rect 11315 -3800 11355 -3790
rect 11425 -3765 11465 -3760
rect 11425 -3795 11430 -3765
rect 11460 -3795 11465 -3765
rect 11425 -3800 11465 -3795
rect 11535 -3765 11575 -3760
rect 11535 -3795 11540 -3765
rect 11570 -3795 11575 -3765
rect 11535 -3800 11575 -3795
rect 11645 -3765 11685 -3760
rect 11645 -3795 11650 -3765
rect 11680 -3795 11685 -3765
rect 11645 -3800 11685 -3795
rect 11755 -3765 11795 -3760
rect 11755 -3795 11760 -3765
rect 11790 -3795 11795 -3765
rect 11755 -3800 11795 -3795
rect 11815 -3770 11845 -3760
rect 11815 -3790 11820 -3770
rect 11840 -3790 11845 -3770
rect 11815 -3800 11845 -3790
rect 11865 -3765 11905 -3760
rect 11865 -3795 11870 -3765
rect 11900 -3795 11905 -3765
rect 11865 -3800 11905 -3795
rect 11975 -3765 12015 -3760
rect 11975 -3795 11980 -3765
rect 12010 -3795 12015 -3765
rect 11975 -3800 12015 -3795
rect 12085 -3765 12125 -3760
rect 12085 -3795 12090 -3765
rect 12120 -3795 12125 -3765
rect 12085 -3800 12125 -3795
rect 12195 -3765 12235 -3760
rect 12195 -3795 12200 -3765
rect 12230 -3795 12235 -3765
rect 12195 -3800 12235 -3795
rect 12305 -3765 12345 -3760
rect 12305 -3795 12310 -3765
rect 12340 -3795 12345 -3765
rect 12305 -3800 12345 -3795
rect 12415 -3765 12455 -3760
rect 12415 -3795 12420 -3765
rect 12450 -3795 12455 -3765
rect 12415 -3800 12455 -3795
rect 12525 -3765 12565 -3760
rect 12525 -3795 12530 -3765
rect 12560 -3795 12565 -3765
rect 12595 -3780 12600 -3750
rect 12630 -3780 12635 -3750
rect 12595 -3785 12635 -3780
rect 12525 -3800 12565 -3795
rect 11165 -4085 11205 -4080
rect 11165 -4115 11170 -4085
rect 11200 -4115 11205 -4085
rect 11165 -4120 11205 -4115
rect 11260 -4085 11300 -4080
rect 11260 -4115 11265 -4085
rect 11295 -4115 11300 -4085
rect 11260 -4120 11300 -4115
rect 11370 -4085 11410 -4080
rect 11370 -4115 11375 -4085
rect 11405 -4115 11410 -4085
rect 11370 -4120 11410 -4115
rect 11480 -4085 11520 -4080
rect 11480 -4115 11485 -4085
rect 11515 -4115 11520 -4085
rect 11480 -4120 11520 -4115
rect 11590 -4085 11630 -4080
rect 11590 -4115 11595 -4085
rect 11625 -4115 11630 -4085
rect 11590 -4120 11630 -4115
rect 11700 -4085 11740 -4080
rect 11700 -4115 11705 -4085
rect 11735 -4115 11740 -4085
rect 11700 -4120 11740 -4115
rect 11810 -4085 11850 -4080
rect 11810 -4115 11815 -4085
rect 11845 -4115 11850 -4085
rect 11810 -4120 11850 -4115
rect 11920 -4085 11960 -4080
rect 11920 -4115 11925 -4085
rect 11955 -4115 11960 -4085
rect 11920 -4120 11960 -4115
rect 12030 -4085 12070 -4080
rect 12030 -4115 12035 -4085
rect 12065 -4115 12070 -4085
rect 12030 -4120 12070 -4115
rect 12140 -4085 12180 -4080
rect 12140 -4115 12145 -4085
rect 12175 -4115 12180 -4085
rect 12140 -4120 12180 -4115
rect 12250 -4085 12290 -4080
rect 12250 -4115 12255 -4085
rect 12285 -4115 12290 -4085
rect 12250 -4120 12290 -4115
rect 12360 -4085 12400 -4080
rect 12360 -4115 12365 -4085
rect 12395 -4115 12400 -4085
rect 12360 -4120 12400 -4115
rect 12470 -4085 12510 -4080
rect 12470 -4115 12475 -4085
rect 12505 -4115 12510 -4085
rect 12470 -4120 12510 -4115
rect 12620 -4085 12660 -4080
rect 12620 -4115 12625 -4085
rect 12655 -4115 12660 -4085
rect 12620 -4120 12660 -4115
<< via1 >>
rect 11635 9050 11665 9055
rect 11635 9030 11640 9050
rect 11640 9030 11660 9050
rect 11660 9030 11665 9050
rect 11635 9025 11665 9030
rect 11755 9050 11785 9055
rect 11755 9030 11760 9050
rect 11760 9030 11780 9050
rect 11780 9030 11785 9050
rect 11755 9025 11785 9030
rect 11875 9050 11905 9055
rect 11875 9030 11880 9050
rect 11880 9030 11900 9050
rect 11900 9030 11905 9050
rect 11875 9025 11905 9030
rect 12085 9025 12115 9055
rect 11205 8990 11235 8995
rect 11205 8970 11210 8990
rect 11210 8970 11230 8990
rect 11230 8970 11235 8990
rect 11205 8965 11235 8970
rect 11465 8990 11495 8995
rect 11465 8970 11470 8990
rect 11470 8970 11490 8990
rect 11490 8970 11495 8990
rect 11465 8965 11495 8970
rect 11575 9005 11605 9010
rect 11575 8985 11580 9005
rect 11580 8985 11600 9005
rect 11600 8985 11605 9005
rect 11575 8980 11605 8985
rect 11695 9005 11725 9010
rect 11695 8985 11700 9005
rect 11700 8985 11720 9005
rect 11720 8985 11725 9005
rect 11695 8980 11725 8985
rect 11815 9005 11845 9010
rect 11815 8985 11820 9005
rect 11820 8985 11840 9005
rect 11840 8985 11845 9005
rect 11815 8980 11845 8985
rect 11935 9005 11965 9010
rect 11935 8985 11940 9005
rect 11940 8985 11960 9005
rect 11960 8985 11965 9005
rect 11935 8980 11965 8985
rect 12085 8980 12115 8985
rect 12085 8960 12090 8980
rect 12090 8960 12110 8980
rect 12110 8960 12115 8980
rect 12085 8955 12115 8960
rect 12205 8980 12235 8985
rect 12205 8960 12210 8980
rect 12210 8960 12230 8980
rect 12230 8960 12235 8980
rect 12205 8955 12235 8960
rect 12325 8980 12355 8985
rect 12325 8960 12330 8980
rect 12330 8960 12350 8980
rect 12350 8960 12355 8980
rect 12325 8955 12355 8960
rect 12445 8980 12475 8985
rect 12445 8960 12450 8980
rect 12450 8960 12470 8980
rect 12470 8960 12475 8980
rect 12445 8955 12475 8960
rect 12565 8980 12595 8985
rect 12565 8960 12570 8980
rect 12570 8960 12590 8980
rect 12590 8960 12595 8980
rect 12565 8955 12595 8960
rect 11335 8835 11340 8860
rect 11340 8835 11360 8860
rect 11360 8835 11365 8860
rect 11335 8830 11365 8835
rect 11755 8850 11785 8855
rect 11755 8830 11760 8850
rect 11760 8830 11780 8850
rect 11780 8830 11785 8850
rect 11755 8825 11785 8830
rect 12145 8850 12175 8855
rect 12145 8830 12150 8850
rect 12150 8830 12170 8850
rect 12170 8830 12175 8850
rect 12145 8825 12175 8830
rect 12265 8850 12295 8855
rect 12265 8830 12270 8850
rect 12270 8830 12290 8850
rect 12290 8830 12295 8850
rect 12265 8825 12295 8830
rect 12385 8850 12415 8855
rect 12385 8830 12390 8850
rect 12390 8830 12410 8850
rect 12410 8830 12415 8850
rect 12385 8825 12415 8830
rect 12505 8850 12535 8855
rect 12505 8830 12510 8850
rect 12510 8830 12530 8850
rect 12530 8830 12535 8850
rect 12505 8825 12535 8830
rect 11335 8735 11365 8765
rect 12205 8735 12235 8765
rect 11345 8620 11375 8625
rect 11345 8600 11350 8620
rect 11350 8600 11370 8620
rect 11370 8600 11375 8620
rect 11345 8595 11375 8600
rect 11465 8620 11495 8625
rect 11465 8600 11470 8620
rect 11470 8600 11490 8620
rect 11490 8600 11495 8620
rect 11465 8595 11495 8600
rect 11585 8620 11615 8625
rect 11585 8600 11590 8620
rect 11590 8600 11610 8620
rect 11610 8600 11615 8620
rect 11585 8595 11615 8600
rect 11705 8620 11735 8625
rect 11705 8600 11710 8620
rect 11710 8600 11730 8620
rect 11730 8600 11735 8620
rect 11705 8595 11735 8600
rect 11825 8620 11855 8625
rect 11825 8600 11830 8620
rect 11830 8600 11850 8620
rect 11850 8600 11855 8620
rect 11825 8595 11855 8600
rect 11945 8620 11975 8625
rect 11945 8600 11950 8620
rect 11950 8600 11970 8620
rect 11970 8600 11975 8620
rect 11945 8595 11975 8600
rect 12065 8620 12095 8625
rect 12065 8600 12070 8620
rect 12070 8600 12090 8620
rect 12090 8600 12095 8620
rect 12065 8595 12095 8600
rect 12185 8620 12215 8625
rect 12185 8600 12190 8620
rect 12190 8600 12210 8620
rect 12210 8600 12215 8620
rect 12185 8595 12215 8600
rect 12305 8620 12335 8625
rect 12305 8600 12310 8620
rect 12310 8600 12330 8620
rect 12330 8600 12335 8620
rect 12305 8595 12335 8600
rect 12425 8620 12455 8625
rect 12425 8600 12430 8620
rect 12430 8600 12450 8620
rect 12450 8600 12455 8620
rect 12425 8595 12455 8600
rect 18845 8620 18875 8625
rect 18845 8600 18850 8620
rect 18850 8600 18870 8620
rect 18870 8600 18875 8620
rect 18845 8595 18875 8600
rect 18965 8620 18995 8625
rect 18965 8600 18970 8620
rect 18970 8600 18990 8620
rect 18990 8600 18995 8620
rect 18965 8595 18995 8600
rect 19085 8620 19115 8625
rect 19085 8600 19090 8620
rect 19090 8600 19110 8620
rect 19110 8600 19115 8620
rect 19085 8595 19115 8600
rect 19205 8620 19235 8625
rect 19205 8600 19210 8620
rect 19210 8600 19230 8620
rect 19230 8600 19235 8620
rect 19205 8595 19235 8600
rect 19325 8620 19355 8625
rect 19325 8600 19330 8620
rect 19330 8600 19350 8620
rect 19350 8600 19355 8620
rect 19325 8595 19355 8600
rect 19445 8620 19475 8625
rect 19445 8600 19450 8620
rect 19450 8600 19470 8620
rect 19470 8600 19475 8620
rect 19445 8595 19475 8600
rect 19565 8620 19595 8625
rect 19565 8600 19570 8620
rect 19570 8600 19590 8620
rect 19590 8600 19595 8620
rect 19565 8595 19595 8600
rect 19685 8620 19715 8625
rect 19685 8600 19690 8620
rect 19690 8600 19710 8620
rect 19710 8600 19715 8620
rect 19685 8595 19715 8600
rect 19805 8620 19835 8625
rect 19805 8600 19810 8620
rect 19810 8600 19830 8620
rect 19830 8600 19835 8620
rect 19805 8595 19835 8600
rect 19925 8620 19955 8625
rect 19925 8600 19930 8620
rect 19930 8600 19950 8620
rect 19950 8600 19955 8620
rect 19925 8595 19955 8600
rect 12955 8285 12985 8290
rect 12955 8265 12960 8285
rect 12960 8265 12980 8285
rect 12980 8265 12985 8285
rect 12955 8260 12985 8265
rect 13065 8285 13095 8290
rect 13065 8265 13070 8285
rect 13070 8265 13090 8285
rect 13090 8265 13095 8285
rect 13065 8260 13095 8265
rect 13175 8285 13205 8290
rect 13175 8265 13180 8285
rect 13180 8265 13200 8285
rect 13200 8265 13205 8285
rect 13175 8260 13205 8265
rect 13285 8285 13315 8290
rect 13285 8265 13290 8285
rect 13290 8265 13310 8285
rect 13310 8265 13315 8285
rect 13285 8260 13315 8265
rect 13395 8285 13425 8290
rect 13395 8265 13400 8285
rect 13400 8265 13420 8285
rect 13420 8265 13425 8285
rect 13395 8260 13425 8265
rect 13505 8285 13535 8290
rect 13505 8265 13510 8285
rect 13510 8265 13530 8285
rect 13530 8265 13535 8285
rect 13505 8260 13535 8265
rect 13615 8285 13645 8290
rect 13615 8265 13620 8285
rect 13620 8265 13640 8285
rect 13640 8265 13645 8285
rect 13615 8260 13645 8265
rect 13725 8285 13755 8290
rect 13725 8265 13730 8285
rect 13730 8265 13750 8285
rect 13750 8265 13755 8285
rect 13725 8260 13755 8265
rect 13835 8285 13865 8290
rect 13835 8265 13840 8285
rect 13840 8265 13860 8285
rect 13860 8265 13865 8285
rect 13835 8260 13865 8265
rect 13945 8285 13975 8290
rect 13945 8265 13950 8285
rect 13950 8265 13970 8285
rect 13970 8265 13975 8285
rect 13945 8260 13975 8265
rect 14055 8285 14085 8290
rect 14055 8265 14060 8285
rect 14060 8265 14080 8285
rect 14080 8265 14085 8285
rect 14055 8260 14085 8265
rect 20450 8285 20480 8290
rect 20450 8265 20455 8285
rect 20455 8265 20475 8285
rect 20475 8265 20480 8285
rect 20450 8260 20480 8265
rect 20560 8285 20590 8290
rect 20560 8265 20565 8285
rect 20565 8265 20585 8285
rect 20585 8265 20590 8285
rect 20560 8260 20590 8265
rect 20670 8285 20700 8290
rect 20670 8265 20675 8285
rect 20675 8265 20695 8285
rect 20695 8265 20700 8285
rect 20670 8260 20700 8265
rect 20780 8285 20810 8290
rect 20780 8265 20785 8285
rect 20785 8265 20805 8285
rect 20805 8265 20810 8285
rect 20780 8260 20810 8265
rect 20890 8285 20920 8290
rect 20890 8265 20895 8285
rect 20895 8265 20915 8285
rect 20915 8265 20920 8285
rect 20890 8260 20920 8265
rect 21000 8285 21030 8290
rect 21000 8265 21005 8285
rect 21005 8265 21025 8285
rect 21025 8265 21030 8285
rect 21000 8260 21030 8265
rect 21110 8285 21140 8290
rect 21110 8265 21115 8285
rect 21115 8265 21135 8285
rect 21135 8265 21140 8285
rect 21110 8260 21140 8265
rect 21220 8285 21250 8290
rect 21220 8265 21225 8285
rect 21225 8265 21245 8285
rect 21245 8265 21250 8285
rect 21220 8260 21250 8265
rect 21330 8285 21360 8290
rect 21330 8265 21335 8285
rect 21335 8265 21355 8285
rect 21355 8265 21360 8285
rect 21330 8260 21360 8265
rect 21440 8285 21470 8290
rect 21440 8265 21445 8285
rect 21445 8265 21465 8285
rect 21465 8265 21470 8285
rect 21440 8260 21470 8265
rect 21550 8285 21580 8290
rect 21550 8265 21555 8285
rect 21555 8265 21575 8285
rect 21575 8265 21580 8285
rect 21550 8260 21580 8265
rect 10585 8205 10615 8210
rect 10585 8185 10590 8205
rect 10590 8185 10610 8205
rect 10610 8185 10615 8205
rect 10585 8180 10615 8185
rect 10985 8205 11015 8210
rect 10985 8185 10990 8205
rect 10990 8185 11010 8205
rect 11010 8185 11015 8205
rect 10985 8180 11015 8185
rect 18085 8205 18115 8210
rect 18085 8185 18090 8205
rect 18090 8185 18110 8205
rect 18110 8185 18115 8205
rect 18085 8180 18115 8185
rect 18485 8205 18515 8210
rect 18485 8185 18490 8205
rect 18490 8185 18510 8205
rect 18510 8185 18515 8205
rect 18485 8180 18515 8185
rect 10905 8125 10935 8155
rect 9740 7665 9770 7670
rect 9740 7645 9745 7665
rect 9745 7645 9765 7665
rect 9765 7645 9770 7665
rect 9740 7640 9770 7645
rect 9850 7665 9880 7670
rect 9850 7645 9855 7665
rect 9855 7645 9875 7665
rect 9875 7645 9880 7665
rect 9850 7640 9880 7645
rect 9960 7665 9990 7670
rect 9960 7645 9965 7665
rect 9965 7645 9985 7665
rect 9985 7645 9990 7665
rect 9960 7640 9990 7645
rect 10070 7665 10100 7670
rect 10070 7645 10075 7665
rect 10075 7645 10095 7665
rect 10095 7645 10100 7665
rect 10070 7640 10100 7645
rect 10180 7665 10210 7670
rect 10180 7645 10185 7665
rect 10185 7645 10205 7665
rect 10205 7645 10210 7665
rect 10180 7640 10210 7645
rect 10290 7665 10320 7670
rect 10290 7645 10295 7665
rect 10295 7645 10315 7665
rect 10315 7645 10320 7665
rect 10290 7640 10320 7645
rect 10400 7665 10430 7670
rect 10400 7645 10405 7665
rect 10405 7645 10425 7665
rect 10425 7645 10430 7665
rect 10400 7640 10430 7645
rect 10510 7665 10540 7670
rect 10510 7645 10515 7665
rect 10515 7645 10535 7665
rect 10535 7645 10540 7665
rect 10510 7640 10540 7645
rect 10620 7665 10650 7670
rect 10620 7645 10625 7665
rect 10625 7645 10645 7665
rect 10645 7645 10650 7665
rect 10620 7640 10650 7645
rect 10730 7665 10760 7670
rect 10730 7645 10735 7665
rect 10735 7645 10755 7665
rect 10755 7645 10760 7665
rect 10730 7640 10760 7645
rect 10840 7665 10870 7670
rect 10840 7645 10845 7665
rect 10845 7645 10865 7665
rect 10865 7645 10870 7665
rect 10840 7640 10870 7645
rect 9795 7495 9825 7500
rect 9795 7475 9800 7495
rect 9800 7475 9820 7495
rect 9820 7475 9825 7495
rect 9795 7470 9825 7475
rect 9905 7495 9935 7500
rect 9905 7475 9910 7495
rect 9910 7475 9930 7495
rect 9930 7475 9935 7495
rect 9905 7470 9935 7475
rect 10015 7495 10045 7500
rect 10015 7475 10020 7495
rect 10020 7475 10040 7495
rect 10040 7475 10045 7495
rect 10015 7470 10045 7475
rect 10125 7495 10155 7500
rect 10125 7475 10130 7495
rect 10130 7475 10150 7495
rect 10150 7475 10155 7495
rect 10125 7470 10155 7475
rect 10235 7495 10265 7500
rect 10235 7475 10240 7495
rect 10240 7475 10260 7495
rect 10260 7475 10265 7495
rect 10235 7470 10265 7475
rect 10345 7495 10375 7500
rect 10345 7475 10350 7495
rect 10350 7475 10370 7495
rect 10370 7475 10375 7495
rect 10345 7470 10375 7475
rect 10455 7495 10485 7500
rect 10455 7475 10460 7495
rect 10460 7475 10480 7495
rect 10480 7475 10485 7495
rect 10455 7470 10485 7475
rect 10565 7495 10595 7500
rect 10565 7475 10570 7495
rect 10570 7475 10590 7495
rect 10590 7475 10595 7495
rect 10565 7470 10595 7475
rect 10675 7495 10705 7500
rect 10675 7475 10680 7495
rect 10680 7475 10700 7495
rect 10700 7475 10705 7495
rect 10675 7470 10705 7475
rect 10785 7495 10815 7500
rect 10785 7475 10790 7495
rect 10790 7475 10810 7495
rect 10810 7475 10815 7495
rect 10785 7470 10815 7475
rect 11826 8150 11854 8155
rect 11826 8130 11831 8150
rect 11831 8130 11849 8150
rect 11849 8130 11854 8150
rect 11826 8125 11854 8130
rect 18405 8125 18435 8155
rect 11285 8070 11315 8100
rect 11525 8070 11555 8100
rect 11765 8070 11795 8100
rect 12005 8070 12035 8100
rect 12245 8070 12275 8100
rect 12485 8070 12515 8100
rect 11405 8025 11435 8055
rect 11645 8025 11675 8055
rect 11885 8025 11915 8055
rect 12125 8025 12155 8055
rect 12365 8025 12395 8055
rect 11345 7970 11375 8000
rect 11405 7970 11435 8000
rect 11585 7970 11615 8000
rect 11825 7970 11855 8000
rect 12065 7970 12095 8000
rect 12305 7970 12335 8000
rect 11465 7940 11495 7945
rect 11465 7920 11470 7940
rect 11470 7920 11490 7940
rect 11490 7920 11495 7940
rect 11465 7915 11495 7920
rect 11705 7940 11735 7945
rect 11705 7920 11710 7940
rect 11710 7920 11730 7940
rect 11730 7920 11735 7940
rect 11705 7915 11735 7920
rect 11945 7940 11975 7945
rect 11945 7920 11950 7940
rect 11950 7920 11970 7940
rect 11970 7920 11975 7940
rect 11945 7915 11975 7920
rect 12185 7940 12215 7945
rect 12185 7920 12190 7940
rect 12190 7920 12210 7940
rect 12210 7920 12215 7940
rect 12185 7915 12215 7920
rect 12425 7940 12455 7945
rect 12425 7920 12430 7940
rect 12430 7920 12450 7940
rect 12450 7920 12455 7940
rect 12425 7915 12455 7920
rect 12485 7915 12515 7945
rect 13010 7915 13040 7920
rect 13010 7895 13015 7915
rect 13015 7895 13035 7915
rect 13035 7895 13040 7915
rect 13010 7890 13040 7895
rect 13120 7915 13150 7920
rect 13120 7895 13125 7915
rect 13125 7895 13145 7915
rect 13145 7895 13150 7915
rect 13120 7890 13150 7895
rect 13230 7915 13260 7920
rect 13230 7895 13235 7915
rect 13235 7895 13255 7915
rect 13255 7895 13260 7915
rect 13230 7890 13260 7895
rect 13340 7915 13370 7920
rect 13340 7895 13345 7915
rect 13345 7895 13365 7915
rect 13365 7895 13370 7915
rect 13340 7890 13370 7895
rect 13450 7915 13480 7920
rect 13450 7895 13455 7915
rect 13455 7895 13475 7915
rect 13475 7895 13480 7915
rect 13450 7890 13480 7895
rect 13560 7915 13590 7920
rect 13560 7895 13565 7915
rect 13565 7895 13585 7915
rect 13585 7895 13590 7915
rect 13560 7890 13590 7895
rect 13670 7915 13700 7920
rect 13670 7895 13675 7915
rect 13675 7895 13695 7915
rect 13695 7895 13700 7915
rect 13670 7890 13700 7895
rect 13780 7915 13810 7920
rect 13780 7895 13785 7915
rect 13785 7895 13805 7915
rect 13805 7895 13810 7915
rect 13780 7890 13810 7895
rect 13890 7915 13920 7920
rect 13890 7895 13895 7915
rect 13895 7895 13915 7915
rect 13915 7895 13920 7915
rect 13890 7890 13920 7895
rect 14000 7915 14030 7920
rect 14000 7895 14005 7915
rect 14005 7895 14025 7915
rect 14025 7895 14030 7915
rect 14000 7890 14030 7895
rect 13065 7800 13095 7830
rect 13065 7750 13095 7780
rect 12695 7700 12725 7730
rect 13065 7700 13095 7730
rect 13685 7800 13715 7830
rect 13685 7750 13715 7780
rect 13685 7700 13715 7730
rect 10985 7445 11015 7475
rect 11826 7470 11854 7475
rect 11826 7450 11831 7470
rect 11831 7450 11849 7470
rect 11849 7450 11854 7470
rect 11826 7445 11854 7450
rect 10816 7435 10844 7440
rect 10816 7415 10821 7435
rect 10821 7415 10839 7435
rect 10839 7415 10844 7435
rect 10816 7410 10844 7415
rect 9805 7375 9840 7380
rect 9805 7350 9810 7375
rect 9810 7350 9835 7375
rect 9835 7350 9840 7375
rect 9805 7345 9840 7350
rect 10640 7375 10675 7380
rect 10640 7350 10645 7375
rect 10645 7350 10670 7375
rect 10670 7350 10675 7375
rect 10640 7345 10675 7350
rect 9805 7315 9840 7320
rect 9805 7290 9810 7315
rect 9810 7290 9835 7315
rect 9835 7290 9840 7315
rect 9805 7285 9840 7290
rect 10640 7315 10675 7320
rect 10640 7290 10645 7315
rect 10645 7290 10670 7315
rect 10670 7290 10675 7315
rect 10640 7285 10675 7290
rect 11285 7390 11315 7420
rect 11525 7390 11555 7420
rect 11765 7390 11795 7420
rect 11405 7345 11435 7375
rect 11645 7345 11675 7375
rect 10816 7275 10844 7280
rect 10816 7255 10821 7275
rect 10821 7255 10839 7275
rect 10839 7255 10844 7275
rect 10816 7250 10844 7255
rect 11445 7250 11475 7280
rect 11665 7250 11695 7280
rect 9795 7215 9825 7220
rect 9795 7195 9800 7215
rect 9800 7195 9820 7215
rect 9820 7195 9825 7215
rect 9795 7190 9825 7195
rect 9905 7215 9935 7220
rect 9905 7195 9910 7215
rect 9910 7195 9930 7215
rect 9930 7195 9935 7215
rect 9905 7190 9935 7195
rect 10015 7215 10045 7220
rect 10015 7195 10020 7215
rect 10020 7195 10040 7215
rect 10040 7195 10045 7215
rect 10015 7190 10045 7195
rect 10125 7215 10155 7220
rect 10125 7195 10130 7215
rect 10130 7195 10150 7215
rect 10150 7195 10155 7215
rect 10125 7190 10155 7195
rect 10235 7215 10265 7220
rect 10235 7195 10240 7215
rect 10240 7195 10260 7215
rect 10260 7195 10265 7215
rect 10235 7190 10265 7195
rect 10345 7215 10375 7220
rect 10345 7195 10350 7215
rect 10350 7195 10370 7215
rect 10370 7195 10375 7215
rect 10345 7190 10375 7195
rect 10455 7215 10485 7220
rect 10455 7195 10460 7215
rect 10460 7195 10480 7215
rect 10480 7195 10485 7215
rect 10455 7190 10485 7195
rect 10565 7215 10595 7220
rect 10565 7195 10570 7215
rect 10570 7195 10590 7215
rect 10590 7195 10595 7215
rect 10565 7190 10595 7195
rect 10675 7215 10705 7220
rect 10675 7195 10680 7215
rect 10680 7195 10700 7215
rect 10700 7195 10705 7215
rect 10675 7190 10705 7195
rect 10785 7215 10815 7220
rect 10785 7195 10790 7215
rect 10790 7195 10810 7215
rect 10810 7195 10815 7215
rect 10785 7190 10815 7195
rect 11335 7205 11365 7235
rect 11555 7205 11585 7235
rect 12005 7390 12035 7420
rect 12245 7390 12275 7420
rect 12485 7390 12515 7420
rect 12955 7665 12985 7670
rect 12955 7645 12960 7665
rect 12960 7645 12980 7665
rect 12980 7645 12985 7665
rect 12955 7640 12985 7645
rect 13065 7665 13095 7670
rect 13065 7645 13070 7665
rect 13070 7645 13090 7665
rect 13090 7645 13095 7665
rect 13065 7640 13095 7645
rect 13175 7665 13205 7670
rect 13175 7645 13180 7665
rect 13180 7645 13200 7665
rect 13200 7645 13205 7665
rect 13175 7640 13205 7645
rect 13285 7665 13315 7670
rect 13285 7645 13290 7665
rect 13290 7645 13310 7665
rect 13310 7645 13315 7665
rect 13285 7640 13315 7645
rect 13395 7665 13425 7670
rect 13395 7645 13400 7665
rect 13400 7645 13420 7665
rect 13420 7645 13425 7665
rect 13395 7640 13425 7645
rect 13505 7665 13535 7670
rect 13505 7645 13510 7665
rect 13510 7645 13530 7665
rect 13530 7645 13535 7665
rect 13505 7640 13535 7645
rect 13615 7665 13645 7670
rect 13615 7645 13620 7665
rect 13620 7645 13640 7665
rect 13640 7645 13645 7665
rect 13615 7640 13645 7645
rect 13725 7665 13755 7670
rect 13725 7645 13730 7665
rect 13730 7645 13750 7665
rect 13750 7645 13755 7665
rect 13725 7640 13755 7645
rect 13835 7665 13865 7670
rect 13835 7645 13840 7665
rect 13840 7645 13860 7665
rect 13860 7645 13865 7665
rect 13835 7640 13865 7645
rect 13945 7665 13975 7670
rect 13945 7645 13950 7665
rect 13950 7645 13970 7665
rect 13970 7645 13975 7665
rect 13945 7640 13975 7645
rect 14055 7665 14085 7670
rect 14055 7645 14060 7665
rect 14060 7645 14080 7665
rect 14080 7645 14085 7665
rect 14055 7640 14085 7645
rect 17240 7665 17270 7670
rect 17240 7645 17245 7665
rect 17245 7645 17265 7665
rect 17265 7645 17270 7665
rect 17240 7640 17270 7645
rect 17350 7665 17380 7670
rect 17350 7645 17355 7665
rect 17355 7645 17375 7665
rect 17375 7645 17380 7665
rect 17350 7640 17380 7645
rect 17460 7665 17490 7670
rect 17460 7645 17465 7665
rect 17465 7645 17485 7665
rect 17485 7645 17490 7665
rect 17460 7640 17490 7645
rect 17570 7665 17600 7670
rect 17570 7645 17575 7665
rect 17575 7645 17595 7665
rect 17595 7645 17600 7665
rect 17570 7640 17600 7645
rect 17680 7665 17710 7670
rect 17680 7645 17685 7665
rect 17685 7645 17705 7665
rect 17705 7645 17710 7665
rect 17680 7640 17710 7645
rect 17790 7665 17820 7670
rect 17790 7645 17795 7665
rect 17795 7645 17815 7665
rect 17815 7645 17820 7665
rect 17790 7640 17820 7645
rect 17900 7665 17930 7670
rect 17900 7645 17905 7665
rect 17905 7645 17925 7665
rect 17925 7645 17930 7665
rect 17900 7640 17930 7645
rect 18010 7665 18040 7670
rect 18010 7645 18015 7665
rect 18015 7645 18035 7665
rect 18035 7645 18040 7665
rect 18010 7640 18040 7645
rect 18120 7665 18150 7670
rect 18120 7645 18125 7665
rect 18125 7645 18145 7665
rect 18145 7645 18150 7665
rect 18120 7640 18150 7645
rect 18230 7665 18260 7670
rect 18230 7645 18235 7665
rect 18235 7645 18255 7665
rect 18255 7645 18260 7665
rect 18230 7640 18260 7645
rect 18340 7665 18370 7670
rect 18340 7645 18345 7665
rect 18345 7645 18365 7665
rect 18365 7645 18370 7665
rect 18340 7640 18370 7645
rect 13010 7495 13040 7500
rect 13010 7475 13015 7495
rect 13015 7475 13035 7495
rect 13035 7475 13040 7495
rect 13010 7470 13040 7475
rect 13120 7495 13150 7500
rect 13120 7475 13125 7495
rect 13125 7475 13145 7495
rect 13145 7475 13150 7495
rect 13120 7470 13150 7475
rect 13230 7495 13260 7500
rect 13230 7475 13235 7495
rect 13235 7475 13255 7495
rect 13255 7475 13260 7495
rect 13230 7470 13260 7475
rect 13340 7495 13370 7500
rect 13340 7475 13345 7495
rect 13345 7475 13365 7495
rect 13365 7475 13370 7495
rect 13340 7470 13370 7475
rect 13450 7495 13480 7500
rect 13450 7475 13455 7495
rect 13455 7475 13475 7495
rect 13475 7475 13480 7495
rect 13450 7470 13480 7475
rect 13560 7495 13590 7500
rect 13560 7475 13565 7495
rect 13565 7475 13585 7495
rect 13585 7475 13590 7495
rect 13560 7470 13590 7475
rect 13670 7495 13700 7500
rect 13670 7475 13675 7495
rect 13675 7475 13695 7495
rect 13695 7475 13700 7495
rect 13670 7470 13700 7475
rect 13780 7495 13810 7500
rect 13780 7475 13785 7495
rect 13785 7475 13805 7495
rect 13805 7475 13810 7495
rect 13780 7470 13810 7475
rect 13890 7495 13920 7500
rect 13890 7475 13895 7495
rect 13895 7475 13915 7495
rect 13915 7475 13920 7495
rect 13890 7470 13920 7475
rect 14000 7495 14030 7500
rect 14000 7475 14005 7495
rect 14005 7475 14025 7495
rect 14025 7475 14030 7495
rect 14000 7470 14030 7475
rect 17295 7495 17325 7500
rect 17295 7475 17300 7495
rect 17300 7475 17320 7495
rect 17320 7475 17325 7495
rect 17295 7470 17325 7475
rect 17405 7495 17435 7500
rect 17405 7475 17410 7495
rect 17410 7475 17430 7495
rect 17430 7475 17435 7495
rect 17405 7470 17435 7475
rect 17515 7495 17545 7500
rect 17515 7475 17520 7495
rect 17520 7475 17540 7495
rect 17540 7475 17545 7495
rect 17515 7470 17545 7475
rect 17625 7495 17655 7500
rect 17625 7475 17630 7495
rect 17630 7475 17650 7495
rect 17650 7475 17655 7495
rect 17625 7470 17655 7475
rect 17735 7495 17765 7500
rect 17735 7475 17740 7495
rect 17740 7475 17760 7495
rect 17760 7475 17765 7495
rect 17735 7470 17765 7475
rect 17845 7495 17875 7500
rect 17845 7475 17850 7495
rect 17850 7475 17870 7495
rect 17870 7475 17875 7495
rect 17845 7470 17875 7475
rect 17955 7495 17985 7500
rect 17955 7475 17960 7495
rect 17960 7475 17980 7495
rect 17980 7475 17985 7495
rect 17955 7470 17985 7475
rect 18065 7495 18095 7500
rect 18065 7475 18070 7495
rect 18070 7475 18090 7495
rect 18090 7475 18095 7495
rect 18065 7470 18095 7475
rect 18175 7495 18205 7500
rect 18175 7475 18180 7495
rect 18180 7475 18200 7495
rect 18200 7475 18205 7495
rect 18175 7470 18205 7475
rect 18285 7495 18315 7500
rect 18285 7475 18290 7495
rect 18290 7475 18310 7495
rect 18310 7475 18315 7495
rect 18285 7470 18315 7475
rect 19326 8150 19354 8155
rect 19326 8130 19331 8150
rect 19331 8130 19349 8150
rect 19349 8130 19354 8150
rect 19326 8125 19354 8130
rect 18785 8070 18815 8100
rect 19025 8070 19055 8100
rect 19265 8070 19295 8100
rect 19505 8070 19535 8100
rect 19745 8070 19775 8100
rect 19985 8070 20015 8100
rect 18905 8025 18935 8055
rect 19145 8025 19175 8055
rect 19385 8025 19415 8055
rect 19625 8025 19655 8055
rect 19865 8025 19895 8055
rect 18845 7970 18875 8000
rect 18905 7970 18935 8000
rect 19085 7970 19115 8000
rect 19325 7970 19355 8000
rect 19565 7970 19595 8000
rect 19805 7970 19835 8000
rect 18965 7940 18995 7945
rect 18965 7920 18970 7940
rect 18970 7920 18990 7940
rect 18990 7920 18995 7940
rect 18965 7915 18995 7920
rect 19205 7940 19235 7945
rect 19205 7920 19210 7940
rect 19210 7920 19230 7940
rect 19230 7920 19235 7940
rect 19205 7915 19235 7920
rect 19445 7940 19475 7945
rect 19445 7920 19450 7940
rect 19450 7920 19470 7940
rect 19470 7920 19475 7940
rect 19445 7915 19475 7920
rect 19685 7940 19715 7945
rect 19685 7920 19690 7940
rect 19690 7920 19710 7940
rect 19710 7920 19715 7940
rect 19685 7915 19715 7920
rect 19925 7940 19955 7945
rect 19925 7920 19930 7940
rect 19930 7920 19950 7940
rect 19950 7920 19955 7940
rect 19925 7915 19955 7920
rect 19985 7915 20015 7945
rect 20505 7915 20535 7920
rect 20505 7895 20510 7915
rect 20510 7895 20530 7915
rect 20530 7895 20535 7915
rect 20505 7890 20535 7895
rect 20615 7915 20645 7920
rect 20615 7895 20620 7915
rect 20620 7895 20640 7915
rect 20640 7895 20645 7915
rect 20615 7890 20645 7895
rect 20725 7915 20755 7920
rect 20725 7895 20730 7915
rect 20730 7895 20750 7915
rect 20750 7895 20755 7915
rect 20725 7890 20755 7895
rect 20835 7915 20865 7920
rect 20835 7895 20840 7915
rect 20840 7895 20860 7915
rect 20860 7895 20865 7915
rect 20835 7890 20865 7895
rect 20945 7915 20975 7920
rect 20945 7895 20950 7915
rect 20950 7895 20970 7915
rect 20970 7895 20975 7915
rect 20945 7890 20975 7895
rect 21055 7915 21085 7920
rect 21055 7895 21060 7915
rect 21060 7895 21080 7915
rect 21080 7895 21085 7915
rect 21055 7890 21085 7895
rect 21165 7915 21195 7920
rect 21165 7895 21170 7915
rect 21170 7895 21190 7915
rect 21190 7895 21195 7915
rect 21165 7890 21195 7895
rect 21275 7915 21305 7920
rect 21275 7895 21280 7915
rect 21280 7895 21300 7915
rect 21300 7895 21305 7915
rect 21275 7890 21305 7895
rect 21385 7915 21415 7920
rect 21385 7895 21390 7915
rect 21390 7895 21410 7915
rect 21410 7895 21415 7915
rect 21385 7890 21415 7895
rect 21495 7915 21525 7920
rect 21495 7895 21500 7915
rect 21500 7895 21520 7915
rect 21520 7895 21525 7915
rect 21495 7890 21525 7895
rect 20560 7800 20590 7830
rect 20560 7750 20590 7780
rect 20195 7700 20225 7730
rect 20560 7700 20590 7730
rect 12981 7435 13009 7440
rect 12981 7415 12986 7435
rect 12986 7415 13004 7435
rect 13004 7415 13009 7435
rect 12981 7410 13009 7415
rect 11885 7345 11915 7375
rect 12125 7345 12155 7375
rect 12365 7345 12395 7375
rect 12695 7345 12725 7375
rect 12980 7345 13010 7375
rect 13150 7375 13185 7380
rect 13150 7350 13155 7375
rect 13155 7350 13180 7375
rect 13180 7350 13185 7375
rect 13150 7345 13185 7350
rect 13985 7375 14020 7380
rect 13985 7350 13990 7375
rect 13990 7350 14015 7375
rect 14015 7350 14020 7375
rect 13985 7345 14020 7350
rect 18485 7445 18515 7475
rect 19326 7470 19354 7475
rect 19326 7450 19331 7470
rect 19331 7450 19349 7470
rect 19349 7450 19354 7470
rect 19326 7445 19354 7450
rect 18316 7435 18344 7440
rect 18316 7415 18321 7435
rect 18321 7415 18339 7435
rect 18339 7415 18344 7435
rect 18316 7410 18344 7415
rect 17305 7375 17340 7380
rect 17305 7350 17310 7375
rect 17310 7350 17335 7375
rect 17335 7350 17340 7375
rect 17305 7345 17340 7350
rect 18140 7375 18175 7380
rect 18140 7350 18145 7375
rect 18145 7350 18170 7375
rect 18170 7350 18175 7375
rect 18140 7345 18175 7350
rect 12820 7295 12850 7325
rect 11885 7250 11915 7280
rect 12105 7250 12135 7280
rect 12325 7250 12355 7280
rect 11775 7205 11805 7235
rect 11995 7205 12025 7235
rect 12215 7205 12245 7235
rect 12435 7205 12465 7235
rect 9740 6995 9770 7000
rect 9740 6975 9745 6995
rect 9745 6975 9763 6995
rect 9763 6975 9770 6995
rect 9740 6970 9770 6975
rect 9850 6995 9880 7000
rect 9850 6975 9855 6995
rect 9855 6975 9873 6995
rect 9873 6975 9880 6995
rect 9850 6970 9880 6975
rect 9960 6995 9990 7000
rect 9960 6975 9965 6995
rect 9965 6975 9983 6995
rect 9983 6975 9990 6995
rect 9960 6970 9990 6975
rect 10070 6995 10100 7000
rect 10070 6975 10075 6995
rect 10075 6975 10093 6995
rect 10093 6975 10100 6995
rect 10070 6970 10100 6975
rect 10180 6995 10210 7000
rect 10180 6975 10185 6995
rect 10185 6975 10203 6995
rect 10203 6975 10210 6995
rect 10180 6970 10210 6975
rect 10290 6995 10320 7000
rect 10290 6975 10295 6995
rect 10295 6975 10313 6995
rect 10313 6975 10320 6995
rect 10290 6970 10320 6975
rect 10400 6995 10430 7000
rect 10400 6975 10405 6995
rect 10405 6975 10423 6995
rect 10423 6975 10430 6995
rect 10400 6970 10430 6975
rect 10510 6995 10540 7000
rect 10510 6975 10515 6995
rect 10515 6975 10533 6995
rect 10533 6975 10540 6995
rect 10510 6970 10540 6975
rect 10620 6995 10650 7000
rect 10620 6975 10625 6995
rect 10625 6975 10643 6995
rect 10643 6975 10650 6995
rect 10620 6970 10650 6975
rect 10730 6995 10760 7000
rect 10730 6975 10735 6995
rect 10735 6975 10753 6995
rect 10753 6975 10760 6995
rect 10730 6970 10760 6975
rect 10840 6995 10870 7000
rect 10840 6975 10845 6995
rect 10845 6975 10863 6995
rect 10863 6975 10870 6995
rect 10840 6970 10870 6975
rect 11390 6955 11420 6960
rect 11390 6935 11395 6955
rect 11395 6935 11415 6955
rect 11415 6935 11420 6955
rect 11390 6930 11420 6935
rect 11610 6955 11640 6960
rect 11610 6935 11615 6955
rect 11615 6935 11635 6955
rect 11635 6935 11640 6955
rect 11610 6930 11640 6935
rect 11830 6955 11860 6960
rect 11830 6935 11835 6955
rect 11835 6935 11855 6955
rect 11855 6935 11860 6955
rect 11830 6930 11860 6935
rect 12050 6955 12080 6960
rect 12050 6935 12055 6955
rect 12055 6935 12075 6955
rect 12075 6935 12080 6955
rect 12050 6930 12080 6935
rect 12270 6955 12300 6960
rect 12270 6935 12275 6955
rect 12275 6935 12295 6955
rect 12295 6935 12300 6955
rect 12270 6930 12300 6935
rect 11500 6875 11530 6905
rect 11720 6875 11750 6905
rect 11940 6875 11970 6905
rect 12160 6875 12190 6905
rect 11195 6820 11225 6850
rect 11415 6820 11445 6850
rect 11090 6755 11120 6760
rect 11090 6735 11095 6755
rect 11095 6735 11115 6755
rect 11115 6735 11120 6755
rect 11090 6730 11120 6735
rect 11310 6755 11340 6760
rect 11310 6735 11315 6755
rect 11315 6735 11335 6755
rect 11335 6735 11340 6755
rect 11310 6730 11340 6735
rect 12380 6875 12410 6905
rect 11645 6820 11675 6850
rect 12235 6820 12265 6850
rect 12455 6820 12485 6850
rect 12685 6820 12715 6850
rect 11825 6775 11855 6805
rect 11945 6775 11975 6805
rect 11530 6755 11560 6760
rect 11530 6735 11535 6755
rect 11535 6735 11555 6755
rect 11555 6735 11560 6755
rect 11530 6730 11560 6735
rect 12130 6755 12160 6760
rect 12130 6735 12135 6755
rect 12135 6735 12155 6755
rect 12155 6735 12160 6755
rect 12130 6730 12160 6735
rect 12350 6755 12380 6760
rect 12350 6735 12355 6755
rect 12355 6735 12375 6755
rect 12375 6735 12380 6755
rect 12350 6730 12380 6735
rect 12570 6755 12600 6760
rect 12570 6735 12575 6755
rect 12575 6735 12595 6755
rect 12595 6735 12600 6755
rect 12570 6730 12600 6735
rect 11240 6710 11266 6715
rect 11240 6690 11243 6710
rect 11243 6690 11260 6710
rect 11260 6690 11266 6710
rect 11240 6685 11266 6690
rect 11460 6710 11486 6715
rect 11460 6690 11463 6710
rect 11463 6690 11480 6710
rect 11480 6690 11486 6710
rect 11460 6685 11486 6690
rect 11604 6710 11630 6715
rect 11604 6690 11610 6710
rect 11610 6690 11627 6710
rect 11627 6690 11630 6710
rect 11604 6685 11630 6690
rect 11870 6710 11896 6715
rect 11870 6690 11876 6710
rect 11876 6690 11893 6710
rect 11893 6690 11896 6710
rect 11870 6685 11896 6690
rect 12280 6710 12306 6715
rect 12280 6690 12283 6710
rect 12283 6690 12300 6710
rect 12300 6690 12306 6710
rect 12280 6685 12306 6690
rect 12500 6710 12526 6715
rect 12500 6690 12503 6710
rect 12503 6690 12520 6710
rect 12520 6690 12526 6710
rect 12500 6685 12526 6690
rect 12644 6710 12670 6715
rect 12644 6690 12650 6710
rect 12650 6690 12667 6710
rect 12667 6690 12670 6710
rect 12644 6685 12670 6690
rect 13150 7315 13185 7320
rect 13150 7290 13155 7315
rect 13155 7290 13180 7315
rect 13180 7290 13185 7315
rect 13150 7285 13185 7290
rect 13985 7315 14020 7320
rect 13985 7290 13990 7315
rect 13990 7290 14015 7315
rect 14015 7290 14020 7315
rect 13985 7285 14020 7290
rect 12981 7275 13009 7280
rect 12981 7255 12986 7275
rect 12986 7255 13004 7275
rect 13004 7255 13009 7275
rect 12981 7250 13009 7255
rect 17305 7315 17340 7320
rect 17305 7290 17310 7315
rect 17310 7290 17335 7315
rect 17335 7290 17340 7315
rect 17305 7285 17340 7290
rect 18140 7315 18175 7320
rect 18140 7290 18145 7315
rect 18145 7290 18170 7315
rect 18170 7290 18175 7315
rect 18140 7285 18175 7290
rect 18785 7390 18815 7420
rect 19025 7390 19055 7420
rect 19265 7390 19295 7420
rect 18905 7345 18935 7375
rect 19145 7345 19175 7375
rect 18316 7275 18344 7280
rect 18316 7255 18321 7275
rect 18321 7255 18339 7275
rect 18339 7255 18344 7275
rect 18316 7250 18344 7255
rect 18945 7250 18975 7280
rect 19165 7250 19195 7280
rect 13010 7215 13040 7220
rect 13010 7195 13015 7215
rect 13015 7195 13035 7215
rect 13035 7195 13040 7215
rect 13010 7190 13040 7195
rect 13120 7215 13150 7220
rect 13120 7195 13125 7215
rect 13125 7195 13145 7215
rect 13145 7195 13150 7215
rect 13120 7190 13150 7195
rect 13230 7215 13260 7220
rect 13230 7195 13235 7215
rect 13235 7195 13255 7215
rect 13255 7195 13260 7215
rect 13230 7190 13260 7195
rect 13340 7215 13370 7220
rect 13340 7195 13345 7215
rect 13345 7195 13365 7215
rect 13365 7195 13370 7215
rect 13340 7190 13370 7195
rect 13450 7215 13480 7220
rect 13450 7195 13455 7215
rect 13455 7195 13475 7215
rect 13475 7195 13480 7215
rect 13450 7190 13480 7195
rect 13560 7215 13590 7220
rect 13560 7195 13565 7215
rect 13565 7195 13585 7215
rect 13585 7195 13590 7215
rect 13560 7190 13590 7195
rect 13670 7215 13700 7220
rect 13670 7195 13675 7215
rect 13675 7195 13695 7215
rect 13695 7195 13700 7215
rect 13670 7190 13700 7195
rect 13780 7215 13810 7220
rect 13780 7195 13785 7215
rect 13785 7195 13805 7215
rect 13805 7195 13810 7215
rect 13780 7190 13810 7195
rect 13890 7215 13920 7220
rect 13890 7195 13895 7215
rect 13895 7195 13915 7215
rect 13915 7195 13920 7215
rect 13890 7190 13920 7195
rect 14000 7215 14030 7220
rect 14000 7195 14005 7215
rect 14005 7195 14025 7215
rect 14025 7195 14030 7215
rect 14000 7190 14030 7195
rect 17295 7215 17325 7220
rect 17295 7195 17300 7215
rect 17300 7195 17320 7215
rect 17320 7195 17325 7215
rect 17295 7190 17325 7195
rect 17405 7215 17435 7220
rect 17405 7195 17410 7215
rect 17410 7195 17430 7215
rect 17430 7195 17435 7215
rect 17405 7190 17435 7195
rect 17515 7215 17545 7220
rect 17515 7195 17520 7215
rect 17520 7195 17540 7215
rect 17540 7195 17545 7215
rect 17515 7190 17545 7195
rect 17625 7215 17655 7220
rect 17625 7195 17630 7215
rect 17630 7195 17650 7215
rect 17650 7195 17655 7215
rect 17625 7190 17655 7195
rect 17735 7215 17765 7220
rect 17735 7195 17740 7215
rect 17740 7195 17760 7215
rect 17760 7195 17765 7215
rect 17735 7190 17765 7195
rect 17845 7215 17875 7220
rect 17845 7195 17850 7215
rect 17850 7195 17870 7215
rect 17870 7195 17875 7215
rect 17845 7190 17875 7195
rect 17955 7215 17985 7220
rect 17955 7195 17960 7215
rect 17960 7195 17980 7215
rect 17980 7195 17985 7215
rect 17955 7190 17985 7195
rect 18065 7215 18095 7220
rect 18065 7195 18070 7215
rect 18070 7195 18090 7215
rect 18090 7195 18095 7215
rect 18065 7190 18095 7195
rect 18175 7215 18205 7220
rect 18175 7195 18180 7215
rect 18180 7195 18200 7215
rect 18200 7195 18205 7215
rect 18175 7190 18205 7195
rect 18285 7215 18315 7220
rect 18285 7195 18290 7215
rect 18290 7195 18310 7215
rect 18310 7195 18315 7215
rect 18285 7190 18315 7195
rect 18835 7205 18865 7235
rect 19055 7205 19085 7235
rect 19505 7390 19535 7420
rect 19745 7390 19775 7420
rect 19985 7390 20015 7420
rect 20450 7665 20480 7670
rect 20450 7645 20455 7665
rect 20455 7645 20475 7665
rect 20475 7645 20480 7665
rect 20450 7640 20480 7645
rect 20560 7665 20590 7670
rect 20560 7645 20565 7665
rect 20565 7645 20585 7665
rect 20585 7645 20590 7665
rect 20560 7640 20590 7645
rect 20670 7665 20700 7670
rect 20670 7645 20675 7665
rect 20675 7645 20695 7665
rect 20695 7645 20700 7665
rect 20670 7640 20700 7645
rect 20780 7665 20810 7670
rect 20780 7645 20785 7665
rect 20785 7645 20805 7665
rect 20805 7645 20810 7665
rect 20780 7640 20810 7645
rect 20890 7665 20920 7670
rect 20890 7645 20895 7665
rect 20895 7645 20915 7665
rect 20915 7645 20920 7665
rect 20890 7640 20920 7645
rect 21000 7665 21030 7670
rect 21000 7645 21005 7665
rect 21005 7645 21025 7665
rect 21025 7645 21030 7665
rect 21000 7640 21030 7645
rect 21110 7665 21140 7670
rect 21110 7645 21115 7665
rect 21115 7645 21135 7665
rect 21135 7645 21140 7665
rect 21110 7640 21140 7645
rect 21220 7665 21250 7670
rect 21220 7645 21225 7665
rect 21225 7645 21245 7665
rect 21245 7645 21250 7665
rect 21220 7640 21250 7645
rect 21330 7665 21360 7670
rect 21330 7645 21335 7665
rect 21335 7645 21355 7665
rect 21355 7645 21360 7665
rect 21330 7640 21360 7645
rect 21440 7665 21470 7670
rect 21440 7645 21445 7665
rect 21445 7645 21465 7665
rect 21465 7645 21470 7665
rect 21440 7640 21470 7645
rect 21550 7665 21580 7670
rect 21550 7645 21555 7665
rect 21555 7645 21575 7665
rect 21575 7645 21580 7665
rect 21550 7640 21580 7645
rect 20505 7495 20535 7500
rect 20505 7475 20510 7495
rect 20510 7475 20530 7495
rect 20530 7475 20535 7495
rect 20505 7470 20535 7475
rect 20615 7495 20645 7500
rect 20615 7475 20620 7495
rect 20620 7475 20640 7495
rect 20640 7475 20645 7495
rect 20615 7470 20645 7475
rect 20725 7495 20755 7500
rect 20725 7475 20730 7495
rect 20730 7475 20750 7495
rect 20750 7475 20755 7495
rect 20725 7470 20755 7475
rect 20835 7495 20865 7500
rect 20835 7475 20840 7495
rect 20840 7475 20860 7495
rect 20860 7475 20865 7495
rect 20835 7470 20865 7475
rect 20945 7495 20975 7500
rect 20945 7475 20950 7495
rect 20950 7475 20970 7495
rect 20970 7475 20975 7495
rect 20945 7470 20975 7475
rect 21055 7495 21085 7500
rect 21055 7475 21060 7495
rect 21060 7475 21080 7495
rect 21080 7475 21085 7495
rect 21055 7470 21085 7475
rect 21165 7495 21195 7500
rect 21165 7475 21170 7495
rect 21170 7475 21190 7495
rect 21190 7475 21195 7495
rect 21165 7470 21195 7475
rect 21275 7495 21305 7500
rect 21275 7475 21280 7495
rect 21280 7475 21300 7495
rect 21300 7475 21305 7495
rect 21275 7470 21305 7475
rect 21385 7495 21415 7500
rect 21385 7475 21390 7495
rect 21390 7475 21410 7495
rect 21410 7475 21415 7495
rect 21385 7470 21415 7475
rect 21495 7495 21525 7500
rect 21495 7475 21500 7495
rect 21500 7475 21520 7495
rect 21520 7475 21525 7495
rect 21495 7470 21525 7475
rect 20476 7435 20504 7440
rect 20476 7415 20481 7435
rect 20481 7415 20499 7435
rect 20499 7415 20504 7435
rect 20476 7410 20504 7415
rect 19385 7345 19415 7375
rect 19625 7345 19655 7375
rect 19865 7345 19895 7375
rect 20195 7345 20225 7375
rect 20475 7345 20505 7375
rect 20645 7375 20680 7380
rect 20645 7350 20650 7375
rect 20650 7350 20675 7375
rect 20675 7350 20680 7375
rect 20645 7345 20680 7350
rect 21480 7375 21515 7380
rect 21480 7350 21485 7375
rect 21485 7350 21510 7375
rect 21510 7350 21515 7375
rect 21480 7345 21515 7350
rect 20320 7295 20350 7325
rect 19385 7250 19415 7280
rect 19605 7250 19635 7280
rect 19825 7250 19855 7280
rect 19275 7205 19305 7235
rect 19495 7205 19525 7235
rect 19715 7205 19745 7235
rect 19935 7205 19965 7235
rect 12955 6995 12985 7000
rect 12955 6975 12962 6995
rect 12962 6975 12980 6995
rect 12980 6975 12985 6995
rect 12955 6970 12985 6975
rect 13065 6995 13095 7000
rect 13065 6975 13072 6995
rect 13072 6975 13090 6995
rect 13090 6975 13095 6995
rect 13065 6970 13095 6975
rect 13175 6995 13205 7000
rect 13175 6975 13182 6995
rect 13182 6975 13200 6995
rect 13200 6975 13205 6995
rect 13175 6970 13205 6975
rect 13285 6995 13315 7000
rect 13285 6975 13292 6995
rect 13292 6975 13310 6995
rect 13310 6975 13315 6995
rect 13285 6970 13315 6975
rect 13395 6995 13425 7000
rect 13395 6975 13402 6995
rect 13402 6975 13420 6995
rect 13420 6975 13425 6995
rect 13395 6970 13425 6975
rect 13505 6995 13535 7000
rect 13505 6975 13512 6995
rect 13512 6975 13530 6995
rect 13530 6975 13535 6995
rect 13505 6970 13535 6975
rect 13615 6995 13645 7000
rect 13615 6975 13622 6995
rect 13622 6975 13640 6995
rect 13640 6975 13645 6995
rect 13615 6970 13645 6975
rect 13725 6995 13755 7000
rect 13725 6975 13732 6995
rect 13732 6975 13750 6995
rect 13750 6975 13755 6995
rect 13725 6970 13755 6975
rect 13835 6995 13865 7000
rect 13835 6975 13842 6995
rect 13842 6975 13860 6995
rect 13860 6975 13865 6995
rect 13835 6970 13865 6975
rect 13945 6995 13975 7000
rect 13945 6975 13952 6995
rect 13952 6975 13970 6995
rect 13970 6975 13975 6995
rect 13945 6970 13975 6975
rect 14055 6995 14085 7000
rect 14055 6975 14062 6995
rect 14062 6975 14080 6995
rect 14080 6975 14085 6995
rect 14055 6970 14085 6975
rect 17240 6995 17270 7000
rect 17240 6975 17245 6995
rect 17245 6975 17263 6995
rect 17263 6975 17270 6995
rect 17240 6970 17270 6975
rect 17350 6995 17380 7000
rect 17350 6975 17355 6995
rect 17355 6975 17373 6995
rect 17373 6975 17380 6995
rect 17350 6970 17380 6975
rect 17460 6995 17490 7000
rect 17460 6975 17465 6995
rect 17465 6975 17483 6995
rect 17483 6975 17490 6995
rect 17460 6970 17490 6975
rect 17570 6995 17600 7000
rect 17570 6975 17575 6995
rect 17575 6975 17593 6995
rect 17593 6975 17600 6995
rect 17570 6970 17600 6975
rect 17680 6995 17710 7000
rect 17680 6975 17685 6995
rect 17685 6975 17703 6995
rect 17703 6975 17710 6995
rect 17680 6970 17710 6975
rect 17790 6995 17820 7000
rect 17790 6975 17795 6995
rect 17795 6975 17813 6995
rect 17813 6975 17820 6995
rect 17790 6970 17820 6975
rect 17900 6995 17930 7000
rect 17900 6975 17905 6995
rect 17905 6975 17923 6995
rect 17923 6975 17930 6995
rect 17900 6970 17930 6975
rect 18010 6995 18040 7000
rect 18010 6975 18015 6995
rect 18015 6975 18033 6995
rect 18033 6975 18040 6995
rect 18010 6970 18040 6975
rect 18120 6995 18150 7000
rect 18120 6975 18125 6995
rect 18125 6975 18143 6995
rect 18143 6975 18150 6995
rect 18120 6970 18150 6975
rect 18230 6995 18260 7000
rect 18230 6975 18235 6995
rect 18235 6975 18253 6995
rect 18253 6975 18260 6995
rect 18230 6970 18260 6975
rect 18340 6995 18370 7000
rect 18340 6975 18345 6995
rect 18345 6975 18363 6995
rect 18363 6975 18370 6995
rect 18340 6970 18370 6975
rect 18890 6955 18920 6960
rect 18890 6935 18895 6955
rect 18895 6935 18915 6955
rect 18915 6935 18920 6955
rect 18890 6930 18920 6935
rect 19110 6955 19140 6960
rect 19110 6935 19115 6955
rect 19115 6935 19135 6955
rect 19135 6935 19140 6955
rect 19110 6930 19140 6935
rect 19330 6955 19360 6960
rect 19330 6935 19335 6955
rect 19335 6935 19355 6955
rect 19355 6935 19360 6955
rect 19330 6930 19360 6935
rect 19550 6955 19580 6960
rect 19550 6935 19555 6955
rect 19555 6935 19575 6955
rect 19575 6935 19580 6955
rect 19550 6930 19580 6935
rect 19770 6955 19800 6960
rect 19770 6935 19775 6955
rect 19775 6935 19795 6955
rect 19795 6935 19800 6955
rect 19770 6930 19800 6935
rect 19000 6875 19030 6905
rect 19220 6875 19250 6905
rect 19440 6875 19470 6905
rect 19660 6875 19690 6905
rect 18695 6820 18725 6850
rect 18915 6820 18945 6850
rect 18590 6755 18620 6760
rect 18590 6735 18595 6755
rect 18595 6735 18615 6755
rect 18615 6735 18620 6755
rect 18590 6730 18620 6735
rect 18810 6755 18840 6760
rect 18810 6735 18815 6755
rect 18815 6735 18835 6755
rect 18835 6735 18840 6755
rect 18810 6730 18840 6735
rect 19880 6875 19910 6905
rect 19145 6820 19175 6850
rect 19735 6820 19765 6850
rect 19955 6820 19985 6850
rect 20185 6820 20215 6850
rect 19325 6775 19355 6805
rect 19445 6775 19475 6805
rect 19030 6755 19060 6760
rect 19030 6735 19035 6755
rect 19035 6735 19055 6755
rect 19055 6735 19060 6755
rect 19030 6730 19060 6735
rect 19630 6755 19660 6760
rect 19630 6735 19635 6755
rect 19635 6735 19655 6755
rect 19655 6735 19660 6755
rect 19630 6730 19660 6735
rect 19850 6755 19880 6760
rect 19850 6735 19855 6755
rect 19855 6735 19875 6755
rect 19875 6735 19880 6755
rect 19850 6730 19880 6735
rect 20070 6755 20100 6760
rect 20070 6735 20075 6755
rect 20075 6735 20095 6755
rect 20095 6735 20100 6755
rect 20070 6730 20100 6735
rect 18740 6710 18766 6715
rect 18740 6690 18743 6710
rect 18743 6690 18760 6710
rect 18760 6690 18766 6710
rect 18740 6685 18766 6690
rect 18960 6710 18986 6715
rect 18960 6690 18963 6710
rect 18963 6690 18980 6710
rect 18980 6690 18986 6710
rect 18960 6685 18986 6690
rect 19104 6710 19130 6715
rect 19104 6690 19110 6710
rect 19110 6690 19127 6710
rect 19127 6690 19130 6710
rect 19104 6685 19130 6690
rect 19370 6710 19396 6715
rect 19370 6690 19376 6710
rect 19376 6690 19393 6710
rect 19393 6690 19396 6710
rect 19370 6685 19396 6690
rect 19780 6710 19806 6715
rect 19780 6690 19783 6710
rect 19783 6690 19800 6710
rect 19800 6690 19806 6710
rect 19780 6685 19806 6690
rect 20000 6710 20026 6715
rect 20000 6690 20003 6710
rect 20003 6690 20020 6710
rect 20020 6690 20026 6710
rect 20000 6685 20026 6690
rect 20144 6710 20170 6715
rect 20144 6690 20150 6710
rect 20150 6690 20167 6710
rect 20167 6690 20170 6710
rect 20144 6685 20170 6690
rect 20645 7315 20680 7320
rect 20645 7290 20650 7315
rect 20650 7290 20675 7315
rect 20675 7290 20680 7315
rect 20645 7285 20680 7290
rect 21480 7315 21515 7320
rect 21480 7290 21485 7315
rect 21485 7290 21510 7315
rect 21510 7290 21515 7315
rect 21480 7285 21515 7290
rect 20476 7275 20504 7280
rect 20476 7255 20481 7275
rect 20481 7255 20499 7275
rect 20499 7255 20504 7275
rect 20476 7250 20504 7255
rect 20505 7215 20535 7220
rect 20505 7195 20510 7215
rect 20510 7195 20530 7215
rect 20530 7195 20535 7215
rect 20505 7190 20535 7195
rect 20615 7215 20645 7220
rect 20615 7195 20620 7215
rect 20620 7195 20640 7215
rect 20640 7195 20645 7215
rect 20615 7190 20645 7195
rect 20725 7215 20755 7220
rect 20725 7195 20730 7215
rect 20730 7195 20750 7215
rect 20750 7195 20755 7215
rect 20725 7190 20755 7195
rect 20835 7215 20865 7220
rect 20835 7195 20840 7215
rect 20840 7195 20860 7215
rect 20860 7195 20865 7215
rect 20835 7190 20865 7195
rect 20945 7215 20975 7220
rect 20945 7195 20950 7215
rect 20950 7195 20970 7215
rect 20970 7195 20975 7215
rect 20945 7190 20975 7195
rect 21055 7215 21085 7220
rect 21055 7195 21060 7215
rect 21060 7195 21080 7215
rect 21080 7195 21085 7215
rect 21055 7190 21085 7195
rect 21165 7215 21195 7220
rect 21165 7195 21170 7215
rect 21170 7195 21190 7215
rect 21190 7195 21195 7215
rect 21165 7190 21195 7195
rect 21275 7215 21305 7220
rect 21275 7195 21280 7215
rect 21280 7195 21300 7215
rect 21300 7195 21305 7215
rect 21275 7190 21305 7195
rect 21385 7215 21415 7220
rect 21385 7195 21390 7215
rect 21390 7195 21410 7215
rect 21410 7195 21415 7215
rect 21385 7190 21415 7195
rect 21495 7215 21525 7220
rect 21495 7195 21500 7215
rect 21500 7195 21520 7215
rect 21520 7195 21525 7215
rect 21495 7190 21525 7195
rect 20450 6995 20480 7000
rect 20450 6975 20457 6995
rect 20457 6975 20475 6995
rect 20475 6975 20480 6995
rect 20450 6970 20480 6975
rect 20560 6995 20590 7000
rect 20560 6975 20567 6995
rect 20567 6975 20585 6995
rect 20585 6975 20590 6995
rect 20560 6970 20590 6975
rect 20670 6995 20700 7000
rect 20670 6975 20677 6995
rect 20677 6975 20695 6995
rect 20695 6975 20700 6995
rect 20670 6970 20700 6975
rect 20780 6995 20810 7000
rect 20780 6975 20787 6995
rect 20787 6975 20805 6995
rect 20805 6975 20810 6995
rect 20780 6970 20810 6975
rect 20890 6995 20920 7000
rect 20890 6975 20897 6995
rect 20897 6975 20915 6995
rect 20915 6975 20920 6995
rect 20890 6970 20920 6975
rect 21000 6995 21030 7000
rect 21000 6975 21007 6995
rect 21007 6975 21025 6995
rect 21025 6975 21030 6995
rect 21000 6970 21030 6975
rect 21110 6995 21140 7000
rect 21110 6975 21117 6995
rect 21117 6975 21135 6995
rect 21135 6975 21140 6995
rect 21110 6970 21140 6975
rect 21220 6995 21250 7000
rect 21220 6975 21227 6995
rect 21227 6975 21245 6995
rect 21245 6975 21250 6995
rect 21220 6970 21250 6975
rect 21330 6995 21360 7000
rect 21330 6975 21337 6995
rect 21337 6975 21355 6995
rect 21355 6975 21360 6995
rect 21330 6970 21360 6975
rect 21440 6995 21470 7000
rect 21440 6975 21447 6995
rect 21447 6975 21465 6995
rect 21465 6975 21470 6995
rect 21440 6970 21470 6975
rect 21550 6995 21580 7000
rect 21550 6975 21557 6995
rect 21557 6975 21575 6995
rect 21575 6975 21580 6995
rect 21550 6970 21580 6975
rect 20550 6900 20580 6905
rect 20550 6880 20555 6900
rect 20555 6880 20575 6900
rect 20575 6880 20580 6900
rect 20550 6875 20580 6880
rect 20660 6900 20690 6905
rect 20660 6880 20665 6900
rect 20665 6880 20685 6900
rect 20685 6880 20690 6900
rect 20660 6875 20690 6880
rect 20770 6900 20800 6905
rect 20770 6880 20775 6900
rect 20775 6880 20795 6900
rect 20795 6880 20800 6900
rect 20770 6875 20800 6880
rect 20570 6675 20596 6680
rect 20570 6655 20571 6675
rect 20571 6655 20591 6675
rect 20591 6655 20596 6675
rect 20570 6650 20596 6655
rect 20515 6625 20545 6630
rect 20515 6605 20520 6625
rect 20520 6605 20540 6625
rect 20540 6605 20545 6625
rect 20515 6600 20545 6605
rect 20621 6600 20651 6630
rect 20715 6600 20745 6630
rect 20805 6625 20835 6630
rect 20805 6605 20810 6625
rect 20810 6605 20830 6625
rect 20830 6605 20835 6625
rect 20805 6600 20835 6605
rect 12820 6540 12850 6570
rect 20320 6540 20350 6570
rect 20475 6565 20501 6570
rect 20475 6545 20476 6565
rect 20476 6545 20496 6565
rect 20496 6545 20501 6565
rect 20475 6540 20501 6545
rect 20849 6565 20875 6570
rect 20849 6545 20854 6565
rect 20854 6545 20874 6565
rect 20874 6545 20875 6565
rect 20849 6540 20875 6545
rect 11109 6490 11135 6495
rect 11109 6470 11112 6490
rect 11112 6470 11129 6490
rect 11129 6470 11135 6490
rect 11109 6465 11135 6470
rect 11310 6490 11340 6495
rect 11310 6470 11315 6490
rect 11315 6470 11335 6490
rect 11335 6470 11340 6490
rect 11310 6465 11340 6470
rect 11530 6490 11560 6495
rect 11530 6470 11535 6490
rect 11535 6470 11555 6490
rect 11555 6470 11560 6490
rect 11530 6465 11560 6470
rect 11925 6490 11951 6495
rect 11925 6470 11928 6490
rect 11928 6470 11945 6490
rect 11945 6470 11951 6490
rect 11925 6465 11951 6470
rect 12149 6490 12175 6495
rect 12149 6470 12152 6490
rect 12152 6470 12169 6490
rect 12169 6470 12175 6490
rect 12149 6465 12175 6470
rect 12350 6490 12380 6495
rect 12350 6470 12355 6490
rect 12355 6470 12375 6490
rect 12375 6470 12380 6490
rect 12350 6465 12380 6470
rect 12570 6490 12600 6495
rect 12570 6470 12575 6490
rect 12575 6470 12595 6490
rect 12595 6470 12600 6490
rect 12570 6465 12600 6470
rect 18609 6490 18635 6495
rect 18609 6470 18612 6490
rect 18612 6470 18629 6490
rect 18629 6470 18635 6490
rect 18609 6465 18635 6470
rect 18810 6490 18840 6495
rect 18810 6470 18815 6490
rect 18815 6470 18835 6490
rect 18835 6470 18840 6490
rect 18810 6465 18840 6470
rect 19030 6490 19060 6495
rect 19030 6470 19035 6490
rect 19035 6470 19055 6490
rect 19055 6470 19060 6490
rect 19030 6465 19060 6470
rect 19425 6490 19451 6495
rect 19425 6470 19428 6490
rect 19428 6470 19445 6490
rect 19445 6470 19451 6490
rect 19425 6465 19451 6470
rect 19649 6490 19675 6495
rect 19649 6470 19652 6490
rect 19652 6470 19669 6490
rect 19669 6470 19675 6490
rect 19649 6465 19675 6470
rect 19850 6490 19880 6495
rect 19850 6470 19855 6490
rect 19855 6470 19875 6490
rect 19875 6470 19880 6490
rect 19850 6465 19880 6470
rect 20070 6490 20100 6495
rect 20070 6470 20075 6490
rect 20075 6470 20095 6490
rect 20095 6470 20100 6490
rect 20070 6465 20100 6470
rect 9765 6440 9800 6445
rect 9765 6415 9770 6440
rect 9770 6415 9795 6440
rect 9795 6415 9800 6440
rect 9765 6410 9800 6415
rect 10775 6440 10810 6445
rect 10775 6415 10780 6440
rect 10780 6415 10805 6440
rect 10805 6415 10810 6440
rect 10775 6410 10810 6415
rect 11150 6430 11180 6435
rect 11150 6410 11155 6430
rect 11155 6410 11175 6430
rect 11175 6410 11180 6430
rect 11150 6405 11180 6410
rect 11255 6430 11285 6435
rect 11255 6410 11260 6430
rect 11260 6410 11280 6430
rect 11280 6410 11285 6430
rect 11255 6405 11285 6410
rect 11365 6430 11395 6435
rect 11365 6410 11370 6430
rect 11370 6410 11390 6430
rect 11390 6410 11395 6430
rect 11365 6405 11395 6410
rect 11475 6430 11505 6435
rect 11475 6410 11480 6430
rect 11480 6410 11500 6430
rect 11500 6410 11505 6430
rect 11475 6405 11505 6410
rect 11585 6430 11615 6435
rect 11585 6410 11590 6430
rect 11590 6410 11610 6430
rect 11610 6410 11615 6430
rect 11585 6405 11615 6410
rect 10670 6360 10700 6390
rect 10775 6360 10805 6390
rect 9770 6330 9800 6335
rect 9770 6310 9775 6330
rect 9775 6310 9795 6330
rect 9795 6310 9800 6330
rect 9770 6305 9800 6310
rect 9970 6330 10000 6335
rect 9970 6310 9975 6330
rect 9975 6310 9995 6330
rect 9995 6310 10000 6330
rect 9970 6305 10000 6310
rect 10170 6330 10200 6335
rect 10170 6310 10175 6330
rect 10175 6310 10195 6330
rect 10195 6310 10200 6330
rect 10170 6305 10200 6310
rect 10370 6330 10400 6335
rect 10370 6310 10375 6330
rect 10375 6310 10395 6330
rect 10395 6310 10400 6330
rect 10370 6305 10400 6310
rect 10570 6330 10600 6335
rect 10570 6310 10575 6330
rect 10575 6310 10595 6330
rect 10595 6310 10600 6330
rect 10570 6305 10600 6310
rect 10770 6330 10800 6335
rect 10770 6310 10775 6330
rect 10775 6310 10795 6330
rect 10795 6310 10800 6330
rect 10770 6305 10800 6310
rect 11815 6315 11845 6345
rect 11320 6265 11350 6295
rect 12190 6430 12220 6435
rect 12190 6410 12195 6430
rect 12195 6410 12215 6430
rect 12215 6410 12220 6430
rect 12190 6405 12220 6410
rect 12295 6430 12325 6435
rect 12295 6410 12300 6430
rect 12300 6410 12320 6430
rect 12320 6410 12325 6430
rect 12295 6405 12325 6410
rect 12405 6430 12435 6435
rect 12405 6410 12410 6430
rect 12410 6410 12430 6430
rect 12430 6410 12435 6430
rect 12405 6405 12435 6410
rect 12515 6430 12545 6435
rect 12515 6410 12520 6430
rect 12520 6410 12540 6430
rect 12540 6410 12545 6430
rect 12515 6405 12545 6410
rect 12625 6430 12655 6435
rect 12625 6410 12630 6430
rect 12630 6410 12650 6430
rect 12650 6410 12655 6430
rect 12625 6405 12655 6410
rect 12990 6440 13025 6445
rect 12990 6415 12995 6440
rect 12995 6415 13020 6440
rect 13020 6415 13025 6440
rect 12990 6410 13025 6415
rect 14000 6440 14035 6445
rect 14000 6415 14005 6440
rect 14005 6415 14030 6440
rect 14030 6415 14035 6440
rect 14000 6410 14035 6415
rect 12995 6360 13025 6390
rect 13100 6360 13130 6390
rect 18650 6430 18680 6435
rect 18650 6410 18655 6430
rect 18655 6410 18675 6430
rect 18675 6410 18680 6430
rect 18650 6405 18680 6410
rect 18755 6430 18785 6435
rect 18755 6410 18760 6430
rect 18760 6410 18780 6430
rect 18780 6410 18785 6430
rect 18755 6405 18785 6410
rect 18865 6430 18895 6435
rect 18865 6410 18870 6430
rect 18870 6410 18890 6430
rect 18890 6410 18895 6430
rect 18865 6405 18895 6410
rect 18975 6430 19005 6435
rect 18975 6410 18980 6430
rect 18980 6410 19000 6430
rect 19000 6410 19005 6430
rect 18975 6405 19005 6410
rect 19085 6430 19115 6435
rect 19085 6410 19090 6430
rect 19090 6410 19110 6430
rect 19110 6410 19115 6430
rect 19085 6405 19115 6410
rect 19315 6355 19345 6385
rect 13000 6330 13030 6335
rect 13000 6310 13005 6330
rect 13005 6310 13025 6330
rect 13025 6310 13030 6330
rect 13000 6305 13030 6310
rect 13200 6330 13230 6335
rect 13200 6310 13205 6330
rect 13205 6310 13225 6330
rect 13225 6310 13230 6330
rect 13200 6305 13230 6310
rect 13400 6330 13430 6335
rect 13400 6310 13405 6330
rect 13405 6310 13425 6330
rect 13425 6310 13430 6330
rect 13400 6305 13430 6310
rect 13600 6330 13630 6335
rect 13600 6310 13605 6330
rect 13605 6310 13625 6330
rect 13625 6310 13630 6330
rect 13600 6305 13630 6310
rect 13800 6330 13830 6335
rect 13800 6310 13805 6330
rect 13805 6310 13825 6330
rect 13825 6310 13830 6330
rect 13800 6305 13830 6310
rect 14000 6330 14030 6335
rect 14000 6310 14005 6330
rect 14005 6310 14025 6330
rect 14025 6310 14030 6330
rect 14000 6305 14030 6310
rect 18820 6305 18850 6335
rect 11885 6265 11915 6295
rect 19690 6430 19720 6435
rect 19690 6410 19695 6430
rect 19695 6410 19715 6430
rect 19715 6410 19720 6430
rect 19690 6405 19720 6410
rect 19795 6430 19825 6435
rect 19795 6410 19800 6430
rect 19800 6410 19820 6430
rect 19820 6410 19825 6430
rect 19795 6405 19825 6410
rect 19905 6430 19935 6435
rect 19905 6410 19910 6430
rect 19910 6410 19930 6430
rect 19930 6410 19935 6430
rect 19905 6405 19935 6410
rect 20015 6430 20045 6435
rect 20015 6410 20020 6430
rect 20020 6410 20040 6430
rect 20040 6410 20045 6430
rect 20015 6405 20045 6410
rect 20125 6430 20155 6435
rect 20125 6410 20130 6430
rect 20130 6410 20150 6430
rect 20150 6410 20155 6430
rect 20125 6405 20155 6410
rect 19385 6305 19415 6335
rect 20528 6345 20554 6350
rect 20528 6325 20533 6345
rect 20533 6325 20553 6345
rect 20553 6325 20554 6345
rect 20528 6320 20554 6325
rect 20796 6345 20822 6350
rect 20796 6325 20797 6345
rect 20797 6325 20817 6345
rect 20817 6325 20822 6345
rect 20796 6320 20822 6325
rect 11430 6230 11460 6235
rect 11430 6210 11435 6230
rect 11435 6210 11455 6230
rect 11455 6210 11460 6230
rect 11430 6205 11460 6210
rect 11540 6230 11570 6235
rect 11540 6210 11545 6230
rect 11545 6210 11565 6230
rect 11565 6210 11570 6230
rect 11540 6205 11570 6210
rect 11650 6230 11680 6235
rect 11650 6210 11655 6230
rect 11655 6210 11675 6230
rect 11675 6210 11680 6230
rect 11650 6205 11680 6210
rect 11760 6230 11790 6235
rect 11760 6210 11765 6230
rect 11765 6210 11785 6230
rect 11785 6210 11790 6230
rect 11760 6205 11790 6210
rect 11870 6230 11900 6235
rect 11870 6210 11875 6230
rect 11875 6210 11895 6230
rect 11895 6210 11900 6230
rect 11870 6205 11900 6210
rect 11980 6230 12010 6235
rect 11980 6210 11985 6230
rect 11985 6210 12005 6230
rect 12005 6210 12010 6230
rect 11980 6205 12010 6210
rect 12090 6230 12120 6235
rect 12090 6210 12095 6230
rect 12095 6210 12115 6230
rect 12115 6210 12120 6230
rect 12090 6205 12120 6210
rect 12200 6230 12230 6235
rect 12200 6210 12205 6230
rect 12205 6210 12225 6230
rect 12225 6210 12230 6230
rect 12200 6205 12230 6210
rect 12310 6230 12340 6235
rect 12310 6210 12315 6230
rect 12315 6210 12335 6230
rect 12335 6210 12340 6230
rect 12310 6205 12340 6210
rect 12420 6230 12450 6235
rect 12420 6210 12425 6230
rect 12425 6210 12445 6230
rect 12445 6210 12450 6230
rect 12420 6205 12450 6210
rect 12530 6230 12560 6235
rect 12530 6210 12535 6230
rect 12535 6210 12555 6230
rect 12555 6210 12560 6230
rect 12530 6205 12560 6210
rect 12600 6245 12630 6250
rect 12600 6225 12605 6245
rect 12605 6225 12625 6245
rect 12625 6225 12630 6245
rect 12600 6220 12630 6225
rect 18930 6270 18960 6275
rect 18930 6250 18935 6270
rect 18935 6250 18955 6270
rect 18955 6250 18960 6270
rect 18930 6245 18960 6250
rect 19040 6270 19070 6275
rect 19040 6250 19045 6270
rect 19045 6250 19065 6270
rect 19065 6250 19070 6270
rect 19040 6245 19070 6250
rect 19150 6270 19180 6275
rect 19150 6250 19155 6270
rect 19155 6250 19175 6270
rect 19175 6250 19180 6270
rect 19150 6245 19180 6250
rect 19260 6270 19290 6275
rect 19260 6250 19265 6270
rect 19265 6250 19285 6270
rect 19285 6250 19290 6270
rect 19260 6245 19290 6250
rect 19370 6270 19400 6275
rect 19370 6250 19375 6270
rect 19375 6250 19395 6270
rect 19395 6250 19400 6270
rect 19370 6245 19400 6250
rect 19480 6270 19510 6275
rect 19480 6250 19485 6270
rect 19485 6250 19505 6270
rect 19505 6250 19510 6270
rect 19480 6245 19510 6250
rect 19590 6270 19620 6275
rect 19590 6250 19595 6270
rect 19595 6250 19615 6270
rect 19615 6250 19620 6270
rect 19590 6245 19620 6250
rect 19700 6270 19730 6275
rect 19700 6250 19705 6270
rect 19705 6250 19725 6270
rect 19725 6250 19730 6270
rect 19700 6245 19730 6250
rect 19810 6270 19840 6275
rect 19810 6250 19815 6270
rect 19815 6250 19835 6270
rect 19835 6250 19840 6270
rect 19810 6245 19840 6250
rect 19920 6270 19950 6275
rect 19920 6250 19925 6270
rect 19925 6250 19945 6270
rect 19945 6250 19950 6270
rect 19920 6245 19950 6250
rect 20030 6270 20060 6275
rect 20030 6250 20035 6270
rect 20035 6250 20055 6270
rect 20055 6250 20060 6270
rect 20030 6245 20060 6250
rect 20100 6285 20130 6290
rect 20100 6265 20105 6285
rect 20105 6265 20125 6285
rect 20125 6265 20130 6285
rect 20100 6260 20130 6265
rect 20450 6285 20480 6290
rect 20450 6265 20455 6285
rect 20455 6265 20475 6285
rect 20475 6265 20480 6285
rect 20450 6260 20480 6265
rect 20565 6285 20595 6290
rect 20565 6265 20570 6285
rect 20570 6265 20590 6285
rect 20590 6265 20595 6285
rect 20565 6260 20595 6265
rect 20660 6260 20690 6290
rect 20755 6285 20785 6290
rect 20755 6265 20760 6285
rect 20760 6265 20780 6285
rect 20780 6265 20785 6285
rect 20755 6260 20785 6265
rect 20870 6285 20900 6290
rect 20870 6265 20875 6285
rect 20875 6265 20895 6285
rect 20895 6265 20900 6285
rect 20870 6260 20900 6265
rect 20605 6225 20635 6230
rect 20605 6205 20610 6225
rect 20610 6205 20630 6225
rect 20630 6205 20635 6225
rect 20605 6200 20635 6205
rect 20660 6225 20690 6230
rect 20660 6205 20665 6225
rect 20665 6205 20685 6225
rect 20685 6205 20690 6225
rect 20660 6200 20690 6205
rect 20715 6225 20745 6230
rect 20715 6205 20720 6225
rect 20720 6205 20740 6225
rect 20740 6205 20745 6225
rect 20715 6200 20745 6205
rect 20870 6200 20900 6230
rect 9870 5980 9900 5985
rect 9870 5960 9875 5980
rect 9875 5960 9895 5980
rect 9895 5960 9900 5980
rect 9870 5955 9900 5960
rect 10070 5980 10100 5985
rect 10070 5960 10075 5980
rect 10075 5960 10095 5980
rect 10095 5960 10100 5980
rect 10070 5955 10100 5960
rect 10270 5980 10300 5985
rect 10270 5960 10275 5980
rect 10275 5960 10295 5980
rect 10295 5960 10300 5980
rect 10270 5955 10300 5960
rect 10470 5980 10500 5985
rect 10470 5960 10475 5980
rect 10475 5960 10495 5980
rect 10495 5960 10500 5980
rect 10470 5955 10500 5960
rect 10670 5980 10700 5985
rect 10670 5960 10675 5980
rect 10675 5960 10695 5980
rect 10695 5960 10700 5980
rect 10670 5955 10700 5960
rect 13100 5980 13130 5985
rect 13100 5960 13105 5980
rect 13105 5960 13125 5980
rect 13125 5960 13130 5980
rect 13100 5955 13130 5960
rect 13300 5980 13330 5985
rect 13300 5960 13305 5980
rect 13305 5960 13325 5980
rect 13325 5960 13330 5980
rect 13300 5955 13330 5960
rect 13500 5980 13530 5985
rect 13500 5960 13505 5980
rect 13505 5960 13525 5980
rect 13525 5960 13530 5980
rect 13500 5955 13530 5960
rect 13700 5980 13730 5985
rect 13700 5960 13705 5980
rect 13705 5960 13725 5980
rect 13725 5960 13730 5980
rect 13700 5955 13730 5960
rect 13900 5980 13930 5985
rect 13900 5960 13905 5980
rect 13905 5960 13925 5980
rect 13925 5960 13930 5980
rect 13900 5955 13930 5960
rect 18670 5950 18700 5955
rect 18670 5930 18675 5950
rect 18675 5930 18695 5950
rect 18695 5930 18700 5950
rect 18670 5925 18700 5930
rect 18765 5950 18795 5955
rect 18765 5930 18770 5950
rect 18770 5930 18790 5950
rect 18790 5930 18795 5950
rect 18765 5925 18795 5930
rect 18875 5950 18905 5955
rect 18875 5930 18880 5950
rect 18880 5930 18900 5950
rect 18900 5930 18905 5950
rect 18875 5925 18905 5930
rect 18985 5950 19015 5955
rect 18985 5930 18990 5950
rect 18990 5930 19010 5950
rect 19010 5930 19015 5950
rect 18985 5925 19015 5930
rect 19095 5950 19125 5955
rect 19095 5930 19100 5950
rect 19100 5930 19120 5950
rect 19120 5930 19125 5950
rect 19095 5925 19125 5930
rect 19205 5950 19235 5955
rect 19205 5930 19210 5950
rect 19210 5930 19230 5950
rect 19230 5930 19235 5950
rect 19205 5925 19235 5930
rect 19315 5950 19345 5955
rect 19315 5930 19320 5950
rect 19320 5930 19340 5950
rect 19340 5930 19345 5950
rect 19315 5925 19345 5930
rect 19425 5950 19455 5955
rect 19425 5930 19430 5950
rect 19430 5930 19450 5950
rect 19450 5930 19455 5950
rect 19425 5925 19455 5930
rect 19535 5950 19565 5955
rect 19535 5930 19540 5950
rect 19540 5930 19560 5950
rect 19560 5930 19565 5950
rect 19535 5925 19565 5930
rect 19645 5950 19675 5955
rect 19645 5930 19650 5950
rect 19650 5930 19670 5950
rect 19670 5930 19675 5950
rect 19645 5925 19675 5930
rect 19755 5950 19785 5955
rect 19755 5930 19760 5950
rect 19760 5930 19780 5950
rect 19780 5930 19785 5950
rect 19755 5925 19785 5930
rect 19865 5950 19895 5955
rect 19865 5930 19870 5950
rect 19870 5930 19890 5950
rect 19890 5930 19895 5950
rect 19865 5925 19895 5930
rect 19975 5950 20005 5955
rect 19975 5930 19980 5950
rect 19980 5930 20000 5950
rect 20000 5930 20005 5950
rect 19975 5925 20005 5930
rect 20125 5950 20155 5955
rect 20125 5930 20130 5950
rect 20130 5930 20150 5950
rect 20150 5930 20155 5950
rect 20125 5925 20155 5930
rect 11170 5910 11200 5915
rect 11170 5890 11175 5910
rect 11175 5890 11195 5910
rect 11195 5890 11200 5910
rect 11170 5885 11200 5890
rect 11265 5910 11295 5915
rect 11265 5890 11270 5910
rect 11270 5890 11290 5910
rect 11290 5890 11295 5910
rect 11265 5885 11295 5890
rect 11375 5910 11405 5915
rect 11375 5890 11380 5910
rect 11380 5890 11400 5910
rect 11400 5890 11405 5910
rect 11375 5885 11405 5890
rect 11485 5910 11515 5915
rect 11485 5890 11490 5910
rect 11490 5890 11510 5910
rect 11510 5890 11515 5910
rect 11485 5885 11515 5890
rect 11595 5910 11625 5915
rect 11595 5890 11600 5910
rect 11600 5890 11620 5910
rect 11620 5890 11625 5910
rect 11595 5885 11625 5890
rect 11705 5910 11735 5915
rect 11705 5890 11710 5910
rect 11710 5890 11730 5910
rect 11730 5890 11735 5910
rect 11705 5885 11735 5890
rect 11815 5910 11845 5915
rect 11815 5890 11820 5910
rect 11820 5890 11840 5910
rect 11840 5890 11845 5910
rect 11815 5885 11845 5890
rect 11925 5910 11955 5915
rect 11925 5890 11930 5910
rect 11930 5890 11950 5910
rect 11950 5890 11955 5910
rect 11925 5885 11955 5890
rect 12035 5910 12065 5915
rect 12035 5890 12040 5910
rect 12040 5890 12060 5910
rect 12060 5890 12065 5910
rect 12035 5885 12065 5890
rect 12145 5910 12175 5915
rect 12145 5890 12150 5910
rect 12150 5890 12170 5910
rect 12170 5890 12175 5910
rect 12145 5885 12175 5890
rect 12255 5910 12285 5915
rect 12255 5890 12260 5910
rect 12260 5890 12280 5910
rect 12280 5890 12285 5910
rect 12255 5885 12285 5890
rect 12365 5910 12395 5915
rect 12365 5890 12370 5910
rect 12370 5890 12390 5910
rect 12390 5890 12395 5910
rect 12365 5885 12395 5890
rect 12475 5910 12505 5915
rect 12475 5890 12480 5910
rect 12480 5890 12500 5910
rect 12500 5890 12505 5910
rect 12475 5885 12505 5890
rect 12625 5910 12655 5915
rect 12625 5890 12630 5910
rect 12630 5890 12650 5910
rect 12650 5890 12655 5910
rect 12625 5885 12655 5890
rect 11635 4510 11665 4515
rect 11635 4490 11640 4510
rect 11640 4490 11660 4510
rect 11660 4490 11665 4510
rect 11635 4485 11665 4490
rect 11755 4510 11785 4515
rect 11755 4490 11760 4510
rect 11760 4490 11780 4510
rect 11780 4490 11785 4510
rect 11755 4485 11785 4490
rect 11875 4510 11905 4515
rect 11875 4490 11880 4510
rect 11880 4490 11900 4510
rect 11900 4490 11905 4510
rect 11875 4485 11905 4490
rect 12085 4485 12115 4515
rect 11205 4450 11235 4455
rect 11205 4430 11210 4450
rect 11210 4430 11230 4450
rect 11230 4430 11235 4450
rect 11205 4425 11235 4430
rect 11465 4450 11495 4455
rect 11465 4430 11470 4450
rect 11470 4430 11490 4450
rect 11490 4430 11495 4450
rect 11465 4425 11495 4430
rect 11575 4465 11605 4470
rect 11575 4445 11580 4465
rect 11580 4445 11600 4465
rect 11600 4445 11605 4465
rect 11575 4440 11605 4445
rect 11695 4465 11725 4470
rect 11695 4445 11700 4465
rect 11700 4445 11720 4465
rect 11720 4445 11725 4465
rect 11695 4440 11725 4445
rect 11815 4465 11845 4470
rect 11815 4445 11820 4465
rect 11820 4445 11840 4465
rect 11840 4445 11845 4465
rect 11815 4440 11845 4445
rect 11935 4465 11965 4470
rect 11935 4445 11940 4465
rect 11940 4445 11960 4465
rect 11960 4445 11965 4465
rect 11935 4440 11965 4445
rect 12085 4440 12115 4445
rect 12085 4420 12090 4440
rect 12090 4420 12110 4440
rect 12110 4420 12115 4440
rect 12085 4415 12115 4420
rect 12205 4440 12235 4445
rect 12205 4420 12210 4440
rect 12210 4420 12230 4440
rect 12230 4420 12235 4440
rect 12205 4415 12235 4420
rect 12325 4440 12355 4445
rect 12325 4420 12330 4440
rect 12330 4420 12350 4440
rect 12350 4420 12355 4440
rect 12325 4415 12355 4420
rect 12445 4440 12475 4445
rect 12445 4420 12450 4440
rect 12450 4420 12470 4440
rect 12470 4420 12475 4440
rect 12445 4415 12475 4420
rect 12565 4440 12595 4445
rect 12565 4420 12570 4440
rect 12570 4420 12590 4440
rect 12590 4420 12595 4440
rect 12565 4415 12595 4420
rect 11055 4285 11085 4315
rect 11335 4295 11340 4320
rect 11340 4295 11360 4320
rect 11360 4295 11365 4320
rect 11335 4290 11365 4295
rect 11755 4310 11785 4315
rect 11755 4290 11760 4310
rect 11760 4290 11780 4310
rect 11780 4290 11785 4310
rect 11755 4285 11785 4290
rect 10215 3630 10245 3635
rect 10215 3610 10220 3630
rect 10220 3610 10240 3630
rect 10240 3610 10245 3630
rect 10215 3605 10245 3610
rect 10325 3630 10355 3635
rect 10325 3610 10330 3630
rect 10330 3610 10350 3630
rect 10350 3610 10355 3630
rect 10325 3605 10355 3610
rect 10435 3630 10465 3635
rect 10435 3610 10440 3630
rect 10440 3610 10460 3630
rect 10460 3610 10465 3630
rect 10435 3605 10465 3610
rect 10545 3630 10575 3635
rect 10545 3610 10550 3630
rect 10550 3610 10570 3630
rect 10570 3610 10575 3630
rect 10545 3605 10575 3610
rect 10655 3630 10685 3635
rect 10655 3610 10660 3630
rect 10660 3610 10680 3630
rect 10680 3610 10685 3630
rect 10655 3605 10685 3610
rect 10765 3630 10795 3635
rect 10765 3610 10770 3630
rect 10770 3610 10790 3630
rect 10790 3610 10795 3630
rect 10765 3605 10795 3610
rect 1266 3495 1296 3525
rect 9905 3525 9935 3555
rect 9955 3525 9985 3555
rect 10005 3525 10035 3555
rect -10 3415 20 3445
rect 945 3415 975 3445
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1210 3310 1240 3340
rect 1165 3255 1195 3285
rect 51 3200 86 3205
rect 51 3175 56 3200
rect 56 3175 81 3200
rect 81 3175 86 3200
rect 51 3170 86 3175
rect 51 3140 86 3145
rect 51 3115 56 3140
rect 56 3115 81 3140
rect 81 3115 86 3140
rect 51 3110 86 3115
rect 1165 3070 1195 3100
rect 51 3060 86 3065
rect 51 3035 56 3060
rect 56 3035 81 3060
rect 81 3035 86 3060
rect 51 3030 86 3035
rect 51 3000 86 3005
rect 51 2975 56 3000
rect 56 2975 81 3000
rect 81 2975 86 3000
rect 51 2970 86 2975
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 4445 3465 4475 3495
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 1266 3195 1301 3200
rect 1266 3170 1271 3195
rect 1271 3170 1296 3195
rect 1296 3170 1301 3195
rect 1266 3165 1301 3170
rect 1266 3135 1301 3140
rect 1266 3110 1271 3135
rect 1271 3110 1296 3135
rect 1296 3110 1301 3135
rect 1266 3105 1301 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 56 2850 91 2855
rect 56 2825 61 2850
rect 61 2825 86 2850
rect 86 2825 91 2850
rect 56 2820 91 2825
rect 729 2850 764 2855
rect 729 2825 734 2850
rect 734 2825 759 2850
rect 759 2825 764 2850
rect 729 2820 764 2825
rect 1210 2820 1240 2850
rect 1266 2835 1301 2840
rect 1266 2810 1271 2835
rect 1271 2810 1296 2835
rect 1296 2810 1301 2835
rect 1266 2805 1301 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 56 2790 91 2795
rect 56 2765 61 2790
rect 61 2765 86 2790
rect 86 2765 91 2790
rect 56 2760 91 2765
rect 729 2790 764 2795
rect 729 2765 734 2790
rect 734 2765 759 2790
rect 759 2765 764 2790
rect 729 2760 764 2765
rect 1266 2715 1296 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1297 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 2740 3210 2770 3240
rect 2625 3155 2655 3185
rect 2525 2950 2555 2980
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2625 2760 2655 2790
rect 2625 2315 2655 2345
rect 5145 3415 5175 3445
rect 5365 3305 5395 3335
rect 4890 3255 4920 3285
rect 4445 3155 4475 3185
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 3990 3050 4020 3080
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 5320 3110 5350 3140
rect 3085 2975 3115 2980
rect 3085 2955 3090 2975
rect 3090 2955 3110 2975
rect 3110 2955 3115 2975
rect 3085 2950 3115 2955
rect 3270 2975 3300 2980
rect 3270 2955 3275 2975
rect 3275 2955 3295 2975
rect 3295 2955 3300 2975
rect 3270 2950 3300 2955
rect 3630 2975 3660 2980
rect 3630 2955 3635 2975
rect 3635 2955 3655 2975
rect 3655 2955 3660 2975
rect 3630 2950 3660 2955
rect 4170 2975 4200 2980
rect 4170 2955 4175 2975
rect 4175 2955 4195 2975
rect 4195 2955 4200 2975
rect 4170 2950 4200 2955
rect 4530 2975 4560 2980
rect 4530 2955 4535 2975
rect 4535 2955 4555 2975
rect 4555 2955 4560 2975
rect 4530 2950 4560 2955
rect 3000 2805 3030 2810
rect 3000 2785 3005 2805
rect 3005 2785 3025 2805
rect 3025 2785 3030 2805
rect 3000 2780 3030 2785
rect 3180 2805 3210 2810
rect 3180 2785 3185 2805
rect 3185 2785 3205 2805
rect 3205 2785 3210 2805
rect 3180 2780 3210 2785
rect 3360 2805 3390 2810
rect 3360 2785 3365 2805
rect 3365 2785 3385 2805
rect 3385 2785 3390 2805
rect 3360 2780 3390 2785
rect 3540 2805 3570 2810
rect 3540 2785 3545 2805
rect 3545 2785 3565 2805
rect 3565 2785 3570 2805
rect 3540 2780 3570 2785
rect 3720 2805 3750 2810
rect 3720 2785 3725 2805
rect 3725 2785 3745 2805
rect 3745 2785 3750 2805
rect 3720 2780 3750 2785
rect 3900 2805 3930 2810
rect 3900 2785 3905 2805
rect 3905 2785 3925 2805
rect 3925 2785 3930 2805
rect 3900 2780 3930 2785
rect 4080 2805 4110 2810
rect 4080 2785 4085 2805
rect 4085 2785 4105 2805
rect 4105 2785 4110 2805
rect 4080 2780 4110 2785
rect 4260 2805 4290 2810
rect 4260 2785 4265 2805
rect 4265 2785 4285 2805
rect 4285 2785 4290 2805
rect 4260 2780 4290 2785
rect 4440 2805 4470 2810
rect 4440 2785 4445 2805
rect 4445 2785 4465 2805
rect 4465 2785 4470 2805
rect 4440 2780 4470 2785
rect 4620 2805 4650 2810
rect 4620 2785 4625 2805
rect 4625 2785 4645 2805
rect 4645 2785 4650 2805
rect 4620 2780 4650 2785
rect 4800 2805 4830 2810
rect 4800 2785 4805 2805
rect 4805 2785 4825 2805
rect 4825 2785 4830 2805
rect 4800 2780 4830 2785
rect 4980 2805 5010 2810
rect 4980 2785 4985 2805
rect 4985 2785 5005 2805
rect 5005 2785 5010 2805
rect 4980 2780 5010 2785
rect 3180 2745 3210 2750
rect 3180 2725 3185 2745
rect 3185 2725 3205 2745
rect 3205 2725 3210 2745
rect 3180 2720 3210 2725
rect 3360 2745 3390 2750
rect 3360 2725 3365 2745
rect 3365 2725 3385 2745
rect 3385 2725 3390 2745
rect 3360 2720 3390 2725
rect 3540 2745 3570 2750
rect 3540 2725 3545 2745
rect 3545 2725 3565 2745
rect 3565 2725 3570 2745
rect 3540 2720 3570 2725
rect 3720 2745 3750 2750
rect 3720 2725 3725 2745
rect 3725 2725 3745 2745
rect 3745 2725 3750 2745
rect 3720 2720 3750 2725
rect 3900 2745 3930 2750
rect 3900 2725 3905 2745
rect 3905 2725 3925 2745
rect 3925 2725 3930 2745
rect 3900 2720 3930 2725
rect 4080 2745 4110 2750
rect 4080 2725 4085 2745
rect 4085 2725 4105 2745
rect 4105 2725 4110 2745
rect 4080 2720 4110 2725
rect 4260 2745 4290 2750
rect 4260 2725 4265 2745
rect 4265 2725 4285 2745
rect 4285 2725 4290 2745
rect 4260 2720 4290 2725
rect 4440 2745 4470 2750
rect 4440 2725 4445 2745
rect 4445 2725 4465 2745
rect 4465 2725 4470 2745
rect 4440 2720 4470 2725
rect 4620 2745 4650 2750
rect 4620 2725 4625 2745
rect 4625 2725 4645 2745
rect 4645 2725 4650 2745
rect 4620 2720 4650 2725
rect 4800 2745 4830 2750
rect 4800 2725 4805 2745
rect 4805 2725 4825 2745
rect 4825 2725 4830 2745
rect 4800 2720 4830 2725
rect 3360 2370 3390 2375
rect 3360 2350 3365 2370
rect 3365 2350 3385 2370
rect 3385 2350 3390 2370
rect 3360 2345 3390 2350
rect 3810 2375 3840 2380
rect 3810 2355 3815 2375
rect 3815 2355 3835 2375
rect 3835 2355 3840 2375
rect 3810 2350 3840 2355
rect 4170 2375 4200 2380
rect 4170 2355 4175 2375
rect 4175 2355 4195 2375
rect 4195 2355 4200 2375
rect 4170 2350 4200 2355
rect 2740 2260 2770 2290
rect 3630 2330 3660 2335
rect 3630 2310 3635 2330
rect 3635 2310 3655 2330
rect 3655 2310 3660 2330
rect 3630 2305 3660 2310
rect 3450 2285 3480 2290
rect 3450 2265 3455 2285
rect 3455 2265 3475 2285
rect 3475 2265 3480 2285
rect 3450 2260 3480 2265
rect 3270 2170 3300 2200
rect 3810 2215 3840 2245
rect 3630 2120 3660 2150
rect 2750 2090 2780 2095
rect 2750 2070 2755 2090
rect 2755 2070 2775 2090
rect 2775 2070 2780 2090
rect 2750 2065 2780 2070
rect 2870 2090 2900 2095
rect 2870 2070 2875 2090
rect 2875 2070 2895 2090
rect 2895 2070 2900 2090
rect 2870 2065 2900 2070
rect 2990 2090 3020 2095
rect 2990 2070 2995 2090
rect 2995 2070 3015 2090
rect 3015 2070 3020 2090
rect 2990 2065 3020 2070
rect 3110 2090 3140 2095
rect 3110 2070 3115 2090
rect 3115 2070 3135 2090
rect 3135 2070 3140 2090
rect 3110 2065 3140 2070
rect 3230 2090 3260 2095
rect 3230 2070 3235 2090
rect 3235 2070 3255 2090
rect 3255 2070 3260 2090
rect 3230 2065 3260 2070
rect 3350 2090 3380 2095
rect 3350 2070 3355 2090
rect 3355 2070 3375 2090
rect 3375 2070 3380 2090
rect 3350 2065 3380 2070
rect 3470 2090 3500 2095
rect 3470 2070 3475 2090
rect 3475 2070 3495 2090
rect 3495 2070 3500 2090
rect 3470 2065 3500 2070
rect 3590 2090 3620 2095
rect 3590 2070 3595 2090
rect 3595 2070 3615 2090
rect 3615 2070 3620 2090
rect 3590 2065 3620 2070
rect 3710 2090 3740 2095
rect 3710 2070 3715 2090
rect 3715 2070 3735 2090
rect 3735 2070 3740 2090
rect 3710 2065 3740 2070
rect 3830 2090 3860 2095
rect 3830 2070 3835 2090
rect 3835 2070 3855 2090
rect 3855 2070 3860 2090
rect 3830 2065 3860 2070
rect 4350 2330 4380 2335
rect 4350 2310 4355 2330
rect 4355 2310 4375 2330
rect 4375 2310 4380 2330
rect 4350 2305 4380 2310
rect 4530 2285 4560 2290
rect 4530 2265 4535 2285
rect 4535 2265 4555 2285
rect 4555 2265 4560 2285
rect 4530 2260 4560 2265
rect 5275 2260 5305 2290
rect 3990 2170 4020 2200
rect 4710 2170 4740 2200
rect 4090 2115 4120 2145
rect 3990 2090 4020 2095
rect 3990 2070 3995 2090
rect 3995 2070 4015 2090
rect 4015 2070 4020 2090
rect 3990 2065 4020 2070
rect 4150 2090 4180 2095
rect 4150 2070 4155 2090
rect 4155 2070 4175 2090
rect 4175 2070 4180 2090
rect 4150 2065 4180 2070
rect 4270 2090 4300 2095
rect 4270 2070 4275 2090
rect 4275 2070 4295 2090
rect 4295 2070 4300 2090
rect 4270 2065 4300 2070
rect 4390 2090 4420 2095
rect 4390 2070 4395 2090
rect 4395 2070 4415 2090
rect 4415 2070 4420 2090
rect 4390 2065 4420 2070
rect 4510 2090 4540 2095
rect 4510 2070 4515 2090
rect 4515 2070 4535 2090
rect 4535 2070 4540 2090
rect 4510 2065 4540 2070
rect 4630 2090 4660 2095
rect 4630 2070 4635 2090
rect 4635 2070 4655 2090
rect 4655 2070 4660 2090
rect 4630 2065 4660 2070
rect 4750 2090 4780 2095
rect 4750 2070 4755 2090
rect 4755 2070 4775 2090
rect 4775 2070 4780 2090
rect 4750 2065 4780 2070
rect 4870 2090 4900 2095
rect 4870 2070 4875 2090
rect 4875 2070 4895 2090
rect 4895 2070 4900 2090
rect 4870 2065 4900 2070
rect 4990 2090 5020 2095
rect 4990 2070 4995 2090
rect 4995 2070 5015 2090
rect 5015 2070 5020 2090
rect 4990 2065 5020 2070
rect 5110 2090 5140 2095
rect 5110 2070 5115 2090
rect 5115 2070 5135 2090
rect 5135 2070 5140 2090
rect 5110 2065 5140 2070
rect 5230 2090 5260 2095
rect 5230 2070 5235 2090
rect 5235 2070 5255 2090
rect 5255 2070 5260 2090
rect 5230 2065 5260 2070
rect 2625 2045 2655 2050
rect 2625 2025 2630 2045
rect 2630 2025 2650 2045
rect 2650 2025 2655 2045
rect 2625 2020 2655 2025
rect 2810 2045 2840 2050
rect 2810 2025 2815 2045
rect 2815 2025 2835 2045
rect 2835 2025 2840 2045
rect 2810 2020 2840 2025
rect 3170 2045 3200 2050
rect 3170 2025 3175 2045
rect 3175 2025 3195 2045
rect 3195 2025 3200 2045
rect 3170 2020 3200 2025
rect 3530 2045 3560 2050
rect 3530 2025 3535 2045
rect 3535 2025 3555 2045
rect 3555 2025 3560 2045
rect 3530 2020 3560 2025
rect 3890 2045 3920 2050
rect 4090 2045 4120 2050
rect 3890 2025 3895 2045
rect 3895 2025 3915 2045
rect 3915 2025 3920 2045
rect 3890 2020 3920 2025
rect 2930 1875 2960 1880
rect 2930 1855 2935 1875
rect 2935 1855 2955 1875
rect 2955 1855 2960 1875
rect 2930 1850 2960 1855
rect 3290 1875 3320 1880
rect 3290 1855 3295 1875
rect 3295 1855 3315 1875
rect 3315 1855 3320 1875
rect 3290 1850 3320 1855
rect 3650 1875 3680 1880
rect 3650 1855 3655 1875
rect 3655 1855 3675 1875
rect 3675 1855 3680 1875
rect 3650 1850 3680 1855
rect 2570 1730 2600 1760
rect 2840 1790 2870 1820
rect 3050 1815 3080 1820
rect 3050 1795 3055 1815
rect 3055 1795 3075 1815
rect 3075 1795 3080 1815
rect 3050 1790 3080 1795
rect 3170 1790 3200 1820
rect 3410 1815 3440 1820
rect 3410 1795 3415 1815
rect 3415 1795 3435 1815
rect 3435 1795 3440 1815
rect 3410 1790 3440 1795
rect 3530 1790 3560 1820
rect 3770 1815 3800 1820
rect 3770 1795 3775 1815
rect 3775 1795 3795 1815
rect 3795 1795 3800 1815
rect 3770 1790 3800 1795
rect 3860 1790 3890 1820
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3230 1755 3260 1760
rect 3230 1735 3235 1755
rect 3235 1735 3255 1755
rect 3255 1735 3260 1755
rect 3230 1730 3260 1735
rect 3290 1755 3320 1760
rect 3290 1735 3295 1755
rect 3295 1735 3315 1755
rect 3315 1735 3320 1755
rect 3290 1730 3320 1735
rect 3530 1755 3560 1760
rect 3530 1735 3535 1755
rect 3535 1735 3555 1755
rect 3555 1735 3560 1755
rect 3530 1730 3560 1735
rect 3770 1755 3800 1760
rect 3770 1735 3775 1755
rect 3775 1735 3795 1755
rect 3795 1735 3800 1755
rect 3770 1730 3800 1735
rect 2805 1680 2835 1710
rect 3170 1710 3200 1715
rect 3170 1690 3175 1710
rect 3175 1690 3195 1710
rect 3195 1690 3200 1710
rect 3170 1685 3200 1690
rect 3410 1710 3440 1715
rect 3410 1690 3415 1710
rect 3415 1690 3435 1710
rect 3435 1690 3440 1710
rect 3410 1685 3440 1690
rect 3650 1710 3680 1715
rect 3650 1690 3655 1710
rect 3655 1690 3675 1710
rect 3675 1690 3680 1710
rect 3650 1685 3680 1690
rect 2625 1635 2655 1665
rect 3170 1590 3200 1595
rect 3170 1570 3175 1590
rect 3175 1570 3195 1590
rect 3195 1570 3200 1590
rect 3170 1565 3200 1570
rect 2840 1515 2870 1545
rect 3230 1540 3260 1545
rect 3230 1520 3235 1540
rect 3235 1520 3255 1540
rect 3255 1520 3260 1540
rect 3230 1515 3260 1520
rect 3350 1540 3380 1545
rect 3350 1520 3355 1540
rect 3355 1520 3375 1540
rect 3375 1520 3380 1540
rect 3350 1515 3380 1520
rect 3470 1540 3500 1545
rect 3470 1520 3475 1540
rect 3475 1520 3495 1540
rect 3495 1520 3500 1540
rect 3470 1515 3500 1520
rect 3590 1540 3620 1545
rect 3590 1520 3595 1540
rect 3595 1520 3615 1540
rect 3615 1520 3620 1540
rect 3590 1515 3620 1520
rect 3710 1540 3740 1545
rect 3710 1520 3715 1540
rect 3715 1520 3735 1540
rect 3735 1520 3740 1540
rect 3710 1515 3740 1520
rect 2930 1495 2960 1500
rect 2930 1475 2935 1495
rect 2935 1475 2955 1495
rect 2955 1475 2960 1495
rect 2930 1470 2960 1475
rect 3050 1495 3080 1500
rect 3050 1475 3055 1495
rect 3055 1475 3075 1495
rect 3075 1475 3080 1495
rect 3050 1470 3080 1475
rect 3170 1495 3200 1500
rect 3170 1475 3175 1495
rect 3175 1475 3195 1495
rect 3195 1475 3200 1495
rect 3170 1470 3200 1475
rect 3290 1495 3320 1500
rect 3290 1475 3295 1495
rect 3295 1475 3315 1495
rect 3315 1475 3320 1495
rect 3290 1470 3320 1475
rect 3530 1495 3560 1500
rect 3530 1475 3535 1495
rect 3535 1475 3555 1495
rect 3555 1475 3560 1495
rect 3530 1470 3560 1475
rect 3650 1495 3680 1500
rect 3650 1475 3655 1495
rect 3655 1475 3675 1495
rect 3675 1475 3680 1495
rect 3650 1470 3680 1475
rect 3770 1495 3800 1500
rect 3770 1475 3775 1495
rect 3775 1475 3795 1495
rect 3795 1475 3800 1495
rect 3770 1470 3800 1475
rect 4090 2025 4095 2045
rect 4095 2025 4115 2045
rect 4115 2025 4120 2045
rect 4090 2020 4120 2025
rect 4450 2045 4480 2050
rect 4450 2025 4455 2045
rect 4455 2025 4475 2045
rect 4475 2025 4480 2045
rect 4450 2020 4480 2025
rect 4810 2045 4840 2050
rect 4810 2025 4815 2045
rect 4815 2025 4835 2045
rect 4835 2025 4840 2045
rect 4810 2020 4840 2025
rect 5170 2045 5200 2050
rect 5170 2025 5175 2045
rect 5175 2025 5195 2045
rect 5195 2025 5200 2045
rect 5170 2020 5200 2025
rect 4330 1875 4360 1880
rect 4330 1855 4335 1875
rect 4335 1855 4355 1875
rect 4355 1855 4360 1875
rect 4330 1850 4360 1855
rect 4690 1875 4720 1880
rect 4690 1855 4695 1875
rect 4695 1855 4715 1875
rect 4715 1855 4720 1875
rect 4690 1850 4720 1855
rect 5050 1875 5080 1880
rect 5050 1855 5055 1875
rect 5055 1855 5075 1875
rect 5075 1855 5080 1875
rect 5050 1850 5080 1855
rect 4120 1790 4150 1820
rect 4210 1815 4240 1820
rect 4210 1795 4215 1815
rect 4215 1795 4235 1815
rect 4235 1795 4240 1815
rect 4210 1790 4240 1795
rect 4450 1790 4480 1820
rect 4570 1815 4600 1820
rect 4570 1795 4575 1815
rect 4575 1795 4595 1815
rect 4595 1795 4600 1815
rect 4570 1790 4600 1795
rect 4210 1755 4240 1760
rect 4210 1735 4215 1755
rect 4215 1735 4235 1755
rect 4235 1735 4240 1755
rect 4210 1730 4240 1735
rect 4450 1755 4480 1760
rect 4450 1735 4455 1755
rect 4455 1735 4475 1755
rect 4475 1735 4480 1755
rect 4450 1730 4480 1735
rect 4810 1790 4840 1820
rect 4930 1815 4960 1820
rect 4930 1795 4935 1815
rect 4935 1795 4955 1815
rect 4955 1795 4960 1815
rect 4930 1790 4960 1795
rect 5140 1790 5170 1820
rect 5320 2115 5350 2145
rect 5415 3255 5445 3285
rect 5365 1790 5395 1820
rect 4690 1755 4720 1760
rect 4690 1735 4695 1755
rect 4695 1735 4715 1755
rect 4715 1735 4720 1755
rect 4690 1730 4720 1735
rect 4750 1755 4780 1760
rect 4750 1735 4755 1755
rect 4755 1735 4775 1755
rect 4775 1735 4780 1755
rect 4750 1730 4780 1735
rect 5275 1730 5305 1760
rect 4330 1710 4360 1715
rect 4330 1690 4335 1710
rect 4335 1690 4355 1710
rect 4355 1690 4360 1710
rect 4330 1685 4360 1690
rect 4570 1710 4600 1715
rect 4570 1690 4575 1710
rect 4575 1690 4595 1710
rect 4595 1690 4600 1710
rect 4570 1685 4600 1690
rect 4810 1710 4840 1715
rect 4810 1690 4815 1710
rect 4815 1690 4835 1710
rect 4835 1690 4840 1710
rect 4810 1685 4840 1690
rect 12145 4310 12175 4315
rect 12145 4290 12150 4310
rect 12150 4290 12170 4310
rect 12170 4290 12175 4310
rect 12145 4285 12175 4290
rect 12265 4310 12295 4315
rect 12265 4290 12270 4310
rect 12270 4290 12290 4310
rect 12290 4290 12295 4310
rect 12265 4285 12295 4290
rect 12385 4310 12415 4315
rect 12385 4290 12390 4310
rect 12390 4290 12410 4310
rect 12410 4290 12415 4310
rect 12385 4285 12415 4290
rect 12505 4310 12535 4315
rect 12505 4290 12510 4310
rect 12510 4290 12530 4310
rect 12530 4290 12535 4310
rect 12505 4285 12535 4290
rect 11110 4230 11140 4260
rect 11335 4230 11365 4260
rect 12205 4230 12235 4260
rect 11055 3125 11085 3155
rect 9905 2905 9935 2935
rect 9955 2905 9985 2935
rect 10005 2905 10035 2935
rect 10270 2960 10300 2965
rect 10270 2940 10275 2960
rect 10275 2940 10295 2960
rect 10295 2940 10300 2960
rect 10270 2935 10300 2940
rect 10380 2960 10410 2965
rect 10380 2940 10385 2960
rect 10385 2940 10405 2960
rect 10405 2940 10410 2960
rect 10380 2935 10410 2940
rect 10490 2960 10520 2965
rect 10490 2940 10495 2960
rect 10495 2940 10515 2960
rect 10515 2940 10520 2960
rect 10490 2935 10520 2940
rect 10600 2960 10630 2965
rect 10600 2940 10605 2960
rect 10605 2940 10625 2960
rect 10625 2940 10630 2960
rect 10600 2935 10630 2940
rect 10710 2960 10740 2965
rect 10710 2940 10715 2960
rect 10715 2940 10735 2960
rect 10735 2940 10740 2960
rect 10710 2935 10740 2940
rect 9955 2850 9985 2880
rect 10655 2850 10685 2880
rect 11005 2850 11035 2880
rect 9750 2795 9780 2825
rect 10380 2795 10410 2825
rect 10215 2700 10245 2705
rect 10215 2680 10220 2700
rect 10220 2680 10240 2700
rect 10240 2680 10245 2700
rect 10215 2675 10245 2680
rect 10325 2700 10355 2705
rect 10325 2680 10330 2700
rect 10330 2680 10350 2700
rect 10350 2680 10355 2700
rect 10325 2675 10355 2680
rect 10435 2700 10465 2705
rect 10435 2680 10440 2700
rect 10440 2680 10460 2700
rect 10460 2680 10465 2700
rect 10435 2675 10465 2680
rect 10545 2700 10575 2705
rect 10545 2680 10550 2700
rect 10550 2680 10570 2700
rect 10570 2680 10575 2700
rect 10545 2675 10575 2680
rect 10655 2700 10685 2705
rect 10655 2680 10660 2700
rect 10660 2680 10680 2700
rect 10680 2680 10685 2700
rect 10655 2675 10685 2680
rect 10765 2700 10795 2705
rect 10765 2680 10770 2700
rect 10770 2680 10790 2700
rect 10790 2680 10795 2700
rect 10765 2675 10795 2680
rect 10025 2405 10055 2435
rect 10270 2430 10300 2435
rect 10270 2410 10275 2430
rect 10275 2410 10295 2430
rect 10295 2410 10300 2430
rect 10270 2405 10300 2410
rect 10380 2430 10410 2435
rect 10380 2410 10385 2430
rect 10385 2410 10405 2430
rect 10405 2410 10410 2430
rect 10380 2405 10410 2410
rect 10490 2430 10520 2435
rect 10490 2410 10495 2430
rect 10495 2410 10515 2430
rect 10515 2410 10520 2430
rect 10490 2405 10520 2410
rect 10600 2430 10630 2435
rect 10600 2410 10605 2430
rect 10605 2410 10625 2430
rect 10625 2410 10630 2430
rect 10600 2405 10630 2410
rect 10710 2430 10740 2435
rect 10710 2410 10715 2430
rect 10715 2410 10735 2430
rect 10735 2410 10740 2430
rect 10710 2405 10740 2410
rect 11365 4200 11395 4205
rect 11365 4180 11370 4200
rect 11370 4180 11390 4200
rect 11390 4180 11395 4200
rect 11365 4175 11395 4180
rect 11475 4200 11505 4205
rect 11475 4180 11480 4200
rect 11480 4180 11500 4200
rect 11500 4180 11505 4200
rect 11475 4175 11505 4180
rect 11585 4200 11615 4205
rect 11585 4180 11590 4200
rect 11590 4180 11610 4200
rect 11610 4180 11615 4200
rect 11585 4175 11615 4180
rect 11695 4200 11725 4205
rect 11695 4180 11700 4200
rect 11700 4180 11720 4200
rect 11720 4180 11725 4200
rect 11695 4175 11725 4180
rect 11805 4200 11835 4205
rect 11805 4180 11810 4200
rect 11810 4180 11830 4200
rect 11830 4180 11835 4200
rect 11805 4175 11835 4180
rect 11915 4200 11945 4205
rect 11915 4180 11920 4200
rect 11920 4180 11940 4200
rect 11940 4180 11945 4200
rect 11915 4175 11945 4180
rect 12025 4200 12055 4205
rect 12025 4180 12030 4200
rect 12030 4180 12050 4200
rect 12050 4180 12055 4200
rect 12025 4175 12055 4180
rect 12135 4200 12165 4205
rect 12135 4180 12140 4200
rect 12140 4180 12160 4200
rect 12160 4180 12165 4200
rect 12135 4175 12165 4180
rect 12245 4200 12275 4205
rect 12245 4180 12250 4200
rect 12250 4180 12270 4200
rect 12270 4180 12275 4200
rect 12245 4175 12275 4180
rect 12355 4200 12385 4205
rect 12355 4180 12360 4200
rect 12360 4180 12380 4200
rect 12380 4180 12385 4200
rect 12355 4175 12385 4180
rect 11310 4080 11340 4085
rect 11310 4060 11315 4080
rect 11315 4060 11335 4080
rect 11335 4060 11340 4080
rect 11310 4055 11340 4060
rect 11530 4080 11560 4085
rect 11530 4060 11535 4080
rect 11535 4060 11555 4080
rect 11555 4060 11560 4080
rect 11530 4055 11560 4060
rect 11750 4080 11780 4085
rect 11750 4060 11755 4080
rect 11755 4060 11775 4080
rect 11775 4060 11780 4080
rect 11750 4055 11780 4060
rect 11970 4080 12000 4085
rect 11970 4060 11975 4080
rect 11975 4060 11995 4080
rect 11995 4060 12000 4080
rect 11970 4055 12000 4060
rect 12190 4080 12220 4085
rect 12190 4060 12195 4080
rect 12195 4060 12215 4080
rect 12215 4060 12220 4080
rect 12190 4055 12220 4060
rect 12410 4080 12440 4085
rect 12410 4060 12415 4080
rect 12415 4060 12435 4080
rect 12435 4060 12440 4080
rect 12410 4055 12440 4060
rect 11315 3955 11345 3960
rect 11315 3935 11320 3955
rect 11320 3935 11340 3955
rect 11340 3935 11345 3955
rect 11315 3930 11345 3935
rect 11420 3995 11450 4025
rect 11640 3995 11670 4025
rect 11860 3995 11890 4025
rect 12080 3995 12110 4025
rect 12300 3995 12330 4025
rect 11420 3955 11450 3960
rect 11420 3935 11425 3955
rect 11425 3935 11445 3955
rect 11445 3935 11450 3955
rect 11420 3930 11450 3935
rect 11530 3955 11560 3960
rect 11530 3935 11535 3955
rect 11535 3935 11555 3955
rect 11555 3935 11560 3955
rect 11530 3930 11560 3935
rect 11640 3955 11670 3960
rect 11640 3935 11645 3955
rect 11645 3935 11665 3955
rect 11665 3935 11670 3955
rect 11640 3930 11670 3935
rect 11750 3955 11780 3960
rect 11750 3935 11755 3955
rect 11755 3935 11775 3955
rect 11775 3935 11780 3955
rect 11750 3930 11780 3935
rect 12055 3955 12085 3960
rect 12055 3935 12060 3955
rect 12060 3935 12080 3955
rect 12080 3935 12085 3955
rect 12055 3930 12085 3935
rect 12160 3955 12190 3960
rect 12160 3935 12165 3955
rect 12165 3935 12185 3955
rect 12185 3935 12190 3955
rect 12160 3930 12190 3935
rect 12270 3955 12300 3960
rect 12270 3935 12275 3955
rect 12275 3935 12295 3955
rect 12295 3935 12300 3955
rect 12270 3930 12300 3935
rect 12380 3955 12410 3960
rect 12380 3935 12385 3955
rect 12385 3935 12405 3955
rect 12405 3935 12410 3955
rect 12380 3930 12410 3935
rect 12490 3955 12520 3960
rect 12490 3935 12495 3955
rect 12495 3935 12515 3955
rect 12515 3935 12520 3955
rect 12490 3930 12520 3935
rect 11274 3895 11300 3900
rect 11274 3875 11277 3895
rect 11277 3875 11294 3895
rect 11294 3875 11300 3895
rect 11274 3870 11300 3875
rect 11475 3895 11505 3900
rect 11475 3875 11480 3895
rect 11480 3875 11500 3895
rect 11500 3875 11505 3895
rect 11475 3870 11505 3875
rect 11695 3895 11725 3900
rect 11695 3875 11700 3895
rect 11700 3875 11720 3895
rect 11720 3875 11725 3895
rect 11695 3870 11725 3875
rect 12014 3895 12040 3900
rect 12014 3875 12017 3895
rect 12017 3875 12034 3895
rect 12034 3875 12040 3895
rect 12014 3870 12040 3875
rect 12215 3895 12245 3900
rect 12215 3875 12220 3895
rect 12220 3875 12240 3895
rect 12240 3875 12245 3895
rect 12215 3870 12245 3875
rect 12435 3895 12465 3900
rect 12435 3875 12440 3895
rect 12440 3875 12460 3895
rect 12460 3875 12465 3895
rect 12435 3870 12465 3875
rect 12765 3870 12795 3900
rect 11405 3775 11431 3780
rect 11405 3755 11408 3775
rect 11408 3755 11425 3775
rect 11425 3755 11431 3775
rect 11405 3750 11431 3755
rect 11625 3775 11651 3780
rect 11625 3755 11628 3775
rect 11628 3755 11645 3775
rect 11645 3755 11651 3775
rect 11625 3750 11651 3755
rect 11769 3775 11795 3780
rect 11769 3755 11775 3775
rect 11775 3755 11792 3775
rect 11792 3755 11795 3775
rect 11769 3750 11795 3755
rect 12145 3775 12171 3780
rect 12145 3755 12148 3775
rect 12148 3755 12165 3775
rect 12165 3755 12171 3775
rect 12145 3750 12171 3755
rect 12365 3775 12391 3780
rect 12365 3755 12368 3775
rect 12368 3755 12385 3775
rect 12385 3755 12391 3775
rect 12365 3750 12391 3755
rect 12509 3775 12535 3780
rect 12509 3755 12515 3775
rect 12515 3755 12532 3775
rect 12532 3755 12535 3775
rect 12509 3750 12535 3755
rect 11255 3715 11285 3720
rect 11255 3695 11260 3715
rect 11260 3695 11280 3715
rect 11280 3695 11285 3715
rect 11255 3690 11285 3695
rect 11360 3715 11390 3720
rect 11360 3695 11365 3715
rect 11365 3695 11385 3715
rect 11385 3695 11390 3715
rect 11360 3690 11390 3695
rect 11475 3715 11505 3720
rect 11475 3695 11480 3715
rect 11480 3695 11500 3715
rect 11500 3695 11505 3715
rect 11475 3690 11505 3695
rect 11580 3715 11610 3720
rect 11580 3695 11585 3715
rect 11585 3695 11605 3715
rect 11605 3695 11610 3715
rect 11580 3690 11610 3695
rect 11695 3715 11725 3720
rect 11695 3695 11700 3715
rect 11700 3695 11720 3715
rect 11720 3695 11725 3715
rect 11695 3690 11725 3695
rect 11810 3715 11840 3720
rect 11810 3695 11815 3715
rect 11815 3695 11835 3715
rect 11835 3695 11840 3715
rect 11810 3690 11840 3695
rect 11995 3725 12025 3730
rect 11995 3705 12000 3725
rect 12000 3705 12020 3725
rect 12020 3705 12025 3725
rect 11995 3700 12025 3705
rect 12215 3725 12245 3730
rect 12215 3705 12220 3725
rect 12220 3705 12240 3725
rect 12240 3705 12245 3725
rect 12215 3700 12245 3705
rect 12435 3725 12465 3730
rect 12435 3705 12440 3725
rect 12440 3705 12460 3725
rect 12460 3705 12465 3725
rect 12435 3700 12465 3705
rect 12100 3655 12130 3685
rect 12320 3655 12350 3685
rect 12550 3655 12580 3685
rect 11345 3620 11375 3625
rect 11345 3600 11350 3620
rect 11350 3600 11370 3620
rect 11370 3600 11375 3620
rect 11345 3595 11375 3600
rect 11465 3620 11495 3625
rect 11465 3600 11470 3620
rect 11470 3600 11490 3620
rect 11490 3600 11495 3620
rect 11465 3595 11495 3600
rect 11585 3620 11615 3625
rect 11585 3600 11590 3620
rect 11590 3600 11610 3620
rect 11610 3600 11615 3620
rect 11585 3595 11615 3600
rect 11705 3620 11735 3625
rect 11705 3600 11710 3620
rect 11710 3600 11730 3620
rect 11730 3600 11735 3620
rect 11705 3595 11735 3600
rect 11825 3620 11855 3625
rect 11825 3600 11830 3620
rect 11830 3600 11850 3620
rect 11850 3600 11855 3620
rect 11825 3595 11855 3600
rect 11945 3620 11975 3625
rect 11945 3600 11950 3620
rect 11950 3600 11970 3620
rect 11970 3600 11975 3620
rect 11945 3595 11975 3600
rect 12065 3620 12095 3625
rect 12065 3600 12070 3620
rect 12070 3600 12090 3620
rect 12090 3600 12095 3620
rect 12065 3595 12095 3600
rect 12185 3620 12215 3625
rect 12185 3600 12190 3620
rect 12190 3600 12210 3620
rect 12210 3600 12215 3620
rect 12185 3595 12215 3600
rect 12305 3620 12335 3625
rect 12305 3600 12310 3620
rect 12310 3600 12330 3620
rect 12330 3600 12335 3620
rect 12305 3595 12335 3600
rect 12425 3620 12455 3625
rect 12425 3600 12430 3620
rect 12430 3600 12450 3620
rect 12450 3600 12455 3620
rect 12425 3595 12455 3600
rect 11826 3150 11854 3155
rect 11826 3130 11831 3150
rect 11831 3130 11849 3150
rect 11849 3130 11854 3150
rect 11826 3125 11854 3130
rect 11285 3070 11315 3100
rect 11525 3070 11555 3100
rect 11765 3070 11795 3100
rect 12005 3070 12035 3100
rect 12245 3070 12275 3100
rect 12485 3070 12515 3100
rect 11405 3025 11435 3055
rect 11645 3025 11675 3055
rect 11885 3025 11915 3055
rect 12125 3025 12155 3055
rect 12365 3025 12395 3055
rect 11345 2970 11375 3000
rect 11405 2970 11435 3000
rect 11585 2970 11615 3000
rect 11825 2970 11855 3000
rect 12065 2970 12095 3000
rect 12305 2970 12335 3000
rect 11465 2940 11495 2945
rect 11465 2920 11470 2940
rect 11470 2920 11490 2940
rect 11490 2920 11495 2940
rect 11465 2915 11495 2920
rect 11705 2940 11735 2945
rect 11705 2920 11710 2940
rect 11710 2920 11730 2940
rect 11730 2920 11735 2940
rect 11705 2915 11735 2920
rect 11945 2940 11975 2945
rect 11945 2920 11950 2940
rect 11950 2920 11970 2940
rect 11970 2920 11975 2940
rect 11945 2915 11975 2920
rect 12185 2940 12215 2945
rect 12185 2920 12190 2940
rect 12190 2920 12210 2940
rect 12210 2920 12215 2940
rect 12185 2915 12215 2920
rect 12425 2940 12455 2945
rect 12425 2920 12430 2940
rect 12430 2920 12450 2940
rect 12450 2920 12455 2940
rect 12425 2915 12455 2920
rect 12485 2915 12515 2945
rect 12695 2850 12725 2880
rect 11110 2445 11140 2475
rect 11826 2470 11854 2475
rect 11826 2450 11831 2470
rect 11831 2450 11849 2470
rect 11849 2450 11854 2470
rect 11826 2445 11854 2450
rect 9790 2000 9825 2005
rect 9790 1975 9795 2000
rect 9795 1975 9820 2000
rect 9820 1975 9825 2000
rect 9790 1970 9825 1975
rect 9850 2000 9885 2005
rect 9850 1975 9855 2000
rect 9855 1975 9880 2000
rect 9880 1975 9885 2000
rect 9850 1970 9885 1975
rect 9910 2000 9945 2005
rect 9910 1975 9915 2000
rect 9915 1975 9940 2000
rect 9940 1975 9945 2000
rect 9910 1970 9945 1975
rect 10770 2385 10800 2390
rect 10770 2365 10775 2385
rect 10775 2365 10795 2385
rect 10795 2365 10800 2385
rect 10770 2360 10800 2365
rect 11005 2390 11035 2420
rect 11285 2390 11315 2420
rect 11525 2390 11555 2420
rect 11765 2390 11795 2420
rect 11405 2345 11435 2375
rect 11645 2345 11675 2375
rect 10070 2285 10100 2315
rect 10270 2310 10300 2315
rect 10270 2290 10275 2310
rect 10275 2290 10295 2310
rect 10295 2290 10300 2310
rect 10270 2285 10300 2290
rect 10380 2310 10410 2315
rect 10380 2290 10385 2310
rect 10385 2290 10405 2310
rect 10405 2290 10410 2310
rect 10380 2285 10410 2290
rect 10490 2310 10520 2315
rect 10490 2290 10495 2310
rect 10495 2290 10515 2310
rect 10515 2290 10520 2310
rect 10490 2285 10520 2290
rect 10600 2310 10630 2315
rect 10600 2290 10605 2310
rect 10605 2290 10625 2310
rect 10625 2290 10630 2310
rect 10600 2285 10630 2290
rect 10710 2310 10740 2315
rect 10710 2290 10715 2310
rect 10715 2290 10735 2310
rect 10735 2290 10740 2310
rect 10710 2285 10740 2290
rect 11005 2295 11035 2325
rect 9970 2000 10005 2005
rect 9970 1975 9975 2000
rect 9975 1975 10000 2000
rect 10000 1975 10005 2000
rect 9970 1970 10005 1975
rect 10025 1970 10055 2000
rect 10955 2150 10985 2180
rect 9915 1915 9945 1945
rect 10070 1915 10100 1945
rect 10215 1940 10245 1945
rect 10215 1920 10220 1940
rect 10220 1920 10238 1940
rect 10238 1920 10245 1940
rect 10215 1915 10245 1920
rect 10325 1940 10355 1945
rect 10325 1920 10330 1940
rect 10330 1920 10348 1940
rect 10348 1920 10355 1940
rect 10325 1915 10355 1920
rect 10435 1940 10465 1945
rect 10435 1920 10440 1940
rect 10440 1920 10458 1940
rect 10458 1920 10465 1940
rect 10435 1915 10465 1920
rect 10545 1940 10575 1945
rect 10545 1920 10550 1940
rect 10550 1920 10568 1940
rect 10568 1920 10575 1940
rect 10545 1915 10575 1920
rect 10655 1940 10685 1945
rect 10655 1920 10660 1940
rect 10660 1920 10678 1940
rect 10678 1920 10685 1940
rect 10655 1915 10685 1920
rect 10765 1940 10795 1945
rect 10765 1920 10770 1940
rect 10770 1920 10788 1940
rect 10788 1920 10795 1940
rect 10765 1915 10795 1920
rect 9795 1865 9825 1895
rect 9970 1730 10000 1760
rect 10560 1730 10590 1760
rect 9750 1675 9780 1705
rect 10035 1675 10065 1705
rect 10260 1700 10290 1705
rect 10260 1680 10265 1700
rect 10265 1680 10285 1700
rect 10285 1680 10290 1700
rect 10260 1675 10290 1680
rect 10460 1700 10490 1705
rect 10460 1680 10465 1700
rect 10465 1680 10485 1700
rect 10485 1680 10490 1700
rect 10460 1675 10490 1680
rect 10660 1700 10690 1705
rect 10660 1680 10665 1700
rect 10665 1680 10685 1700
rect 10685 1680 10690 1700
rect 10660 1675 10690 1680
rect 10840 1675 10870 1705
rect 9970 1640 10005 1645
rect 9970 1615 9975 1640
rect 9975 1615 10000 1640
rect 10000 1615 10005 1640
rect 9970 1610 10005 1615
rect 10030 1640 10065 1645
rect 10030 1615 10035 1640
rect 10035 1615 10060 1640
rect 10060 1615 10065 1640
rect 10030 1610 10065 1615
rect 4810 1590 4840 1595
rect 4810 1570 4815 1590
rect 4815 1570 4835 1590
rect 4835 1570 4840 1590
rect 4810 1565 4840 1570
rect 5415 1565 5445 1595
rect 4270 1540 4300 1545
rect 4270 1520 4275 1540
rect 4275 1520 4295 1540
rect 4295 1520 4300 1540
rect 4270 1515 4300 1520
rect 4390 1540 4420 1545
rect 4390 1520 4395 1540
rect 4395 1520 4415 1540
rect 4415 1520 4420 1540
rect 4390 1515 4420 1520
rect 4510 1540 4540 1545
rect 4510 1520 4515 1540
rect 4515 1520 4535 1540
rect 4535 1520 4540 1540
rect 4510 1515 4540 1520
rect 4630 1540 4660 1545
rect 4630 1520 4635 1540
rect 4635 1520 4655 1540
rect 4655 1520 4660 1540
rect 4630 1515 4660 1520
rect 4750 1540 4780 1545
rect 4750 1520 4755 1540
rect 4755 1520 4775 1540
rect 4775 1520 4780 1540
rect 4750 1515 4780 1520
rect 5140 1515 5170 1545
rect 4210 1495 4240 1500
rect 4210 1475 4215 1495
rect 4215 1475 4235 1495
rect 4235 1475 4240 1495
rect 4210 1470 4240 1475
rect 4330 1495 4360 1500
rect 4330 1475 4335 1495
rect 4335 1475 4355 1495
rect 4355 1475 4360 1495
rect 4330 1470 4360 1475
rect 4450 1495 4480 1500
rect 4450 1475 4455 1495
rect 4455 1475 4475 1495
rect 4475 1475 4480 1495
rect 4450 1470 4480 1475
rect 4690 1495 4720 1500
rect 4690 1475 4695 1495
rect 4695 1475 4715 1495
rect 4715 1475 4720 1495
rect 4690 1470 4720 1475
rect 4810 1495 4840 1500
rect 4810 1475 4815 1495
rect 4815 1475 4835 1495
rect 4835 1475 4840 1495
rect 4810 1470 4840 1475
rect 4930 1495 4960 1500
rect 4930 1475 4935 1495
rect 4935 1475 4955 1495
rect 4955 1475 4960 1495
rect 4930 1470 4960 1475
rect 5050 1495 5080 1500
rect 5050 1475 5055 1495
rect 5055 1475 5075 1495
rect 5075 1475 5080 1495
rect 5050 1470 5080 1475
rect 10840 1360 10870 1390
rect 3380 1180 3410 1185
rect 3380 1160 3385 1180
rect 3385 1160 3405 1180
rect 3405 1160 3410 1180
rect 3380 1155 3410 1160
rect 3990 1155 4020 1185
rect 4600 1180 4630 1185
rect 4600 1160 4605 1180
rect 4605 1160 4625 1180
rect 4625 1160 4630 1180
rect 4600 1155 4630 1160
rect 2950 1120 2980 1125
rect 2950 1100 2955 1120
rect 2955 1100 2975 1120
rect 2975 1100 2980 1120
rect 2950 1095 2980 1100
rect 3030 1120 3060 1125
rect 3030 1100 3035 1120
rect 3035 1100 3055 1120
rect 3055 1100 3060 1120
rect 3030 1095 3060 1100
rect 3110 1120 3140 1125
rect 3110 1100 3115 1120
rect 3115 1100 3135 1120
rect 3135 1100 3140 1120
rect 3110 1095 3140 1100
rect 3190 1120 3220 1125
rect 3190 1100 3195 1120
rect 3195 1100 3215 1120
rect 3215 1100 3220 1120
rect 3190 1095 3220 1100
rect 3270 1120 3300 1125
rect 3270 1100 3275 1120
rect 3275 1100 3295 1120
rect 3295 1100 3300 1120
rect 3270 1095 3300 1100
rect 3350 1120 3380 1125
rect 3350 1100 3355 1120
rect 3355 1100 3375 1120
rect 3375 1100 3380 1120
rect 3350 1095 3380 1100
rect 3430 1120 3460 1125
rect 3430 1100 3435 1120
rect 3435 1100 3455 1120
rect 3455 1100 3460 1120
rect 3430 1095 3460 1100
rect 3510 1120 3540 1125
rect 3510 1100 3515 1120
rect 3515 1100 3535 1120
rect 3535 1100 3540 1120
rect 3510 1095 3540 1100
rect 3590 1120 3620 1125
rect 3590 1100 3595 1120
rect 3595 1100 3615 1120
rect 3615 1100 3620 1120
rect 3590 1095 3620 1100
rect 3670 1120 3700 1125
rect 3670 1100 3675 1120
rect 3675 1100 3695 1120
rect 3695 1100 3700 1120
rect 3670 1095 3700 1100
rect 3750 1120 3780 1125
rect 3750 1100 3755 1120
rect 3755 1100 3775 1120
rect 3775 1100 3780 1120
rect 3750 1095 3780 1100
rect 3830 1120 3860 1125
rect 3830 1100 3835 1120
rect 3835 1100 3855 1120
rect 3855 1100 3860 1120
rect 3830 1095 3860 1100
rect 3910 1120 3940 1125
rect 3910 1100 3915 1120
rect 3915 1100 3935 1120
rect 3935 1100 3940 1120
rect 3910 1095 3940 1100
rect 3990 1120 4020 1125
rect 3990 1100 3995 1120
rect 3995 1100 4015 1120
rect 4015 1100 4020 1120
rect 3990 1095 4020 1100
rect 4070 1120 4100 1125
rect 4070 1100 4075 1120
rect 4075 1100 4095 1120
rect 4095 1100 4100 1120
rect 4070 1095 4100 1100
rect 4150 1120 4180 1125
rect 4150 1100 4155 1120
rect 4155 1100 4175 1120
rect 4175 1100 4180 1120
rect 4150 1095 4180 1100
rect 4230 1120 4260 1125
rect 4230 1100 4235 1120
rect 4235 1100 4255 1120
rect 4255 1100 4260 1120
rect 4230 1095 4260 1100
rect 4310 1120 4340 1125
rect 4310 1100 4315 1120
rect 4315 1100 4335 1120
rect 4335 1100 4340 1120
rect 4310 1095 4340 1100
rect 4390 1120 4420 1125
rect 4390 1100 4395 1120
rect 4395 1100 4415 1120
rect 4415 1100 4420 1120
rect 4390 1095 4420 1100
rect 4470 1120 4500 1125
rect 4470 1100 4475 1120
rect 4475 1100 4495 1120
rect 4495 1100 4500 1120
rect 4470 1095 4500 1100
rect 4550 1120 4580 1125
rect 4550 1100 4555 1120
rect 4555 1100 4575 1120
rect 4575 1100 4580 1120
rect 4550 1095 4580 1100
rect 4630 1120 4660 1125
rect 4630 1100 4635 1120
rect 4635 1100 4655 1120
rect 4655 1100 4660 1120
rect 4630 1095 4660 1100
rect 4710 1120 4740 1125
rect 4710 1100 4715 1120
rect 4715 1100 4735 1120
rect 4735 1100 4740 1120
rect 4710 1095 4740 1100
rect 4790 1120 4820 1125
rect 4790 1100 4795 1120
rect 4795 1100 4815 1120
rect 4815 1100 4820 1120
rect 4790 1095 4820 1100
rect 4870 1120 4900 1125
rect 4870 1100 4875 1120
rect 4875 1100 4895 1120
rect 4895 1100 4900 1120
rect 4870 1095 4900 1100
rect 4950 1120 4980 1125
rect 4950 1100 4955 1120
rect 4955 1100 4975 1120
rect 4975 1100 4980 1120
rect 4950 1095 4980 1100
rect 2625 1010 2655 1040
rect 2910 1035 2940 1040
rect 2910 1015 2915 1035
rect 2915 1015 2935 1035
rect 2935 1015 2940 1035
rect 2910 1010 2940 1015
rect 5115 1035 5145 1040
rect 5115 1015 5120 1035
rect 5120 1015 5140 1035
rect 5140 1015 5145 1035
rect 5115 1010 5145 1015
rect 3000 925 3030 930
rect 3000 905 3005 925
rect 3005 905 3025 925
rect 3025 905 3030 925
rect 3000 900 3030 905
rect 3180 925 3210 930
rect 3180 905 3185 925
rect 3185 905 3205 925
rect 3205 905 3210 925
rect 3180 900 3210 905
rect 3360 925 3390 930
rect 3360 905 3365 925
rect 3365 905 3385 925
rect 3385 905 3390 925
rect 3360 900 3390 905
rect 3540 925 3570 930
rect 3540 905 3545 925
rect 3545 905 3565 925
rect 3565 905 3570 925
rect 3540 900 3570 905
rect 3720 925 3750 930
rect 3720 905 3725 925
rect 3725 905 3745 925
rect 3745 905 3750 925
rect 3720 900 3750 905
rect 3900 925 3930 930
rect 3900 905 3905 925
rect 3905 905 3925 925
rect 3925 905 3930 925
rect 3900 900 3930 905
rect 4080 925 4110 930
rect 4080 905 4085 925
rect 4085 905 4105 925
rect 4105 905 4110 925
rect 4080 900 4110 905
rect 4260 925 4290 930
rect 4260 905 4265 925
rect 4265 905 4285 925
rect 4285 905 4290 925
rect 4260 900 4290 905
rect 4440 925 4470 930
rect 4440 905 4445 925
rect 4445 905 4465 925
rect 4465 905 4470 925
rect 4440 900 4470 905
rect 4620 925 4650 930
rect 4620 905 4625 925
rect 4625 905 4645 925
rect 4645 905 4650 925
rect 4620 900 4650 905
rect 4800 925 4830 930
rect 4800 905 4805 925
rect 4805 905 4825 925
rect 4825 905 4830 925
rect 4800 900 4830 905
rect 4980 925 5010 930
rect 4980 905 4985 925
rect 4985 905 5005 925
rect 5005 905 5010 925
rect 4980 900 5010 905
rect 10360 930 10390 935
rect 10360 910 10365 930
rect 10365 910 10385 930
rect 10385 910 10390 930
rect 10360 905 10390 910
rect 10560 930 10590 935
rect 10560 910 10565 930
rect 10565 910 10585 930
rect 10585 910 10590 930
rect 10560 905 10590 910
rect 11445 2250 11475 2280
rect 11665 2250 11695 2280
rect 11335 2205 11365 2235
rect 11555 2205 11585 2235
rect 12005 2390 12035 2420
rect 12245 2390 12275 2420
rect 12485 2390 12515 2420
rect 11885 2345 11915 2375
rect 12125 2345 12155 2375
rect 12365 2345 12395 2375
rect 12695 2345 12725 2375
rect 12865 3700 12895 3730
rect 12810 3655 12840 3685
rect 12765 2295 12795 2325
rect 11885 2250 11915 2280
rect 12105 2250 12135 2280
rect 12325 2250 12355 2280
rect 11775 2205 11805 2235
rect 11995 2205 12025 2235
rect 12215 2205 12245 2235
rect 12435 2205 12465 2235
rect 11831 2175 11859 2180
rect 11831 2155 11836 2175
rect 11836 2155 11854 2175
rect 11854 2155 11859 2175
rect 11831 2150 11859 2155
rect 11390 1955 11420 1960
rect 11390 1935 11395 1955
rect 11395 1935 11415 1955
rect 11415 1935 11420 1955
rect 11390 1930 11420 1935
rect 11610 1955 11640 1960
rect 11610 1935 11615 1955
rect 11615 1935 11635 1955
rect 11635 1935 11640 1955
rect 11610 1930 11640 1935
rect 11830 1955 11860 1960
rect 11830 1935 11835 1955
rect 11835 1935 11855 1955
rect 11855 1935 11860 1955
rect 11830 1930 11860 1935
rect 12050 1955 12080 1960
rect 12050 1935 12055 1955
rect 12055 1935 12075 1955
rect 12075 1935 12080 1955
rect 12050 1930 12080 1935
rect 12270 1955 12300 1960
rect 12270 1935 12275 1955
rect 12275 1935 12295 1955
rect 12295 1935 12300 1955
rect 12270 1930 12300 1935
rect 11005 1865 11035 1895
rect 11500 1875 11530 1905
rect 11720 1875 11750 1905
rect 11940 1875 11970 1905
rect 12160 1875 12190 1905
rect 11195 1820 11225 1850
rect 11415 1820 11445 1850
rect 11090 1755 11120 1760
rect 11090 1735 11095 1755
rect 11095 1735 11115 1755
rect 11115 1735 11120 1755
rect 11090 1730 11120 1735
rect 11310 1755 11340 1760
rect 11310 1735 11315 1755
rect 11315 1735 11335 1755
rect 11335 1735 11340 1755
rect 11310 1730 11340 1735
rect 12380 1875 12410 1905
rect 12765 1865 12795 1895
rect 11645 1820 11675 1850
rect 12235 1820 12265 1850
rect 12455 1820 12485 1850
rect 12685 1820 12715 1850
rect 11825 1775 11855 1805
rect 11945 1775 11975 1805
rect 11530 1755 11560 1760
rect 11530 1735 11535 1755
rect 11535 1735 11555 1755
rect 11555 1735 11560 1755
rect 11530 1730 11560 1735
rect 12130 1755 12160 1760
rect 12130 1735 12135 1755
rect 12135 1735 12155 1755
rect 12155 1735 12160 1755
rect 12130 1730 12160 1735
rect 12350 1755 12380 1760
rect 12350 1735 12355 1755
rect 12355 1735 12375 1755
rect 12375 1735 12380 1755
rect 12350 1730 12380 1735
rect 12570 1755 12600 1760
rect 12570 1735 12575 1755
rect 12575 1735 12595 1755
rect 12595 1735 12600 1755
rect 12570 1730 12600 1735
rect 11240 1710 11266 1715
rect 11240 1690 11243 1710
rect 11243 1690 11260 1710
rect 11260 1690 11266 1710
rect 11240 1685 11266 1690
rect 11460 1710 11486 1715
rect 11460 1690 11463 1710
rect 11463 1690 11480 1710
rect 11480 1690 11486 1710
rect 11460 1685 11486 1690
rect 11604 1710 11630 1715
rect 11604 1690 11610 1710
rect 11610 1690 11627 1710
rect 11627 1690 11630 1710
rect 11604 1685 11630 1690
rect 11870 1710 11896 1715
rect 11870 1690 11876 1710
rect 11876 1690 11893 1710
rect 11893 1690 11896 1710
rect 11870 1685 11896 1690
rect 12280 1710 12306 1715
rect 12280 1690 12283 1710
rect 12283 1690 12300 1710
rect 12300 1690 12306 1710
rect 12280 1685 12306 1690
rect 12500 1710 12526 1715
rect 12500 1690 12503 1710
rect 12503 1690 12520 1710
rect 12520 1690 12526 1710
rect 12500 1685 12526 1690
rect 12644 1710 12670 1715
rect 12644 1690 12650 1710
rect 12650 1690 12667 1710
rect 12667 1690 12670 1710
rect 12644 1685 12670 1690
rect 11109 1490 11135 1495
rect 11109 1470 11112 1490
rect 11112 1470 11129 1490
rect 11129 1470 11135 1490
rect 11109 1465 11135 1470
rect 11310 1490 11340 1495
rect 11310 1470 11315 1490
rect 11315 1470 11335 1490
rect 11335 1470 11340 1490
rect 11310 1465 11340 1470
rect 11530 1490 11560 1495
rect 11530 1470 11535 1490
rect 11535 1470 11555 1490
rect 11555 1470 11560 1490
rect 11530 1465 11560 1470
rect 11925 1490 11951 1495
rect 11925 1470 11928 1490
rect 11928 1470 11945 1490
rect 11945 1470 11951 1490
rect 11925 1465 11951 1470
rect 12149 1490 12175 1495
rect 12149 1470 12152 1490
rect 12152 1470 12169 1490
rect 12169 1470 12175 1490
rect 12149 1465 12175 1470
rect 12350 1490 12380 1495
rect 12350 1470 12355 1490
rect 12355 1470 12375 1490
rect 12375 1470 12380 1490
rect 12350 1465 12380 1470
rect 12570 1490 12600 1495
rect 12570 1470 12575 1490
rect 12575 1470 12595 1490
rect 12595 1470 12600 1490
rect 12570 1465 12600 1470
rect 11150 1430 11180 1435
rect 11150 1410 11155 1430
rect 11155 1410 11175 1430
rect 11175 1410 11180 1430
rect 11150 1405 11180 1410
rect 11255 1430 11285 1435
rect 11255 1410 11260 1430
rect 11260 1410 11280 1430
rect 11280 1410 11285 1430
rect 11255 1405 11285 1410
rect 11365 1430 11395 1435
rect 11365 1410 11370 1430
rect 11370 1410 11390 1430
rect 11390 1410 11395 1430
rect 11365 1405 11395 1410
rect 11475 1430 11505 1435
rect 11475 1410 11480 1430
rect 11480 1410 11500 1430
rect 11500 1410 11505 1430
rect 11475 1405 11505 1410
rect 11585 1430 11615 1435
rect 11585 1410 11590 1430
rect 11590 1410 11610 1430
rect 11610 1410 11615 1430
rect 11585 1405 11615 1410
rect 11010 1315 11040 1345
rect 11815 1315 11845 1345
rect 11320 1265 11350 1295
rect 12190 1430 12220 1435
rect 12190 1410 12195 1430
rect 12195 1410 12215 1430
rect 12215 1410 12220 1430
rect 12190 1405 12220 1410
rect 12295 1430 12325 1435
rect 12295 1410 12300 1430
rect 12300 1410 12320 1430
rect 12320 1410 12325 1430
rect 12295 1405 12325 1410
rect 12405 1430 12435 1435
rect 12405 1410 12410 1430
rect 12410 1410 12430 1430
rect 12430 1410 12435 1430
rect 12405 1405 12435 1410
rect 12515 1430 12545 1435
rect 12515 1410 12520 1430
rect 12520 1410 12540 1430
rect 12540 1410 12545 1430
rect 12515 1405 12545 1410
rect 12625 1430 12655 1435
rect 12625 1410 12630 1430
rect 12630 1410 12650 1430
rect 12650 1410 12655 1430
rect 12625 1405 12655 1410
rect 11885 1265 11915 1295
rect 11430 1230 11460 1235
rect 11430 1210 11435 1230
rect 11435 1210 11455 1230
rect 11455 1210 11460 1230
rect 11430 1205 11460 1210
rect 11540 1230 11570 1235
rect 11540 1210 11545 1230
rect 11545 1210 11565 1230
rect 11565 1210 11570 1230
rect 11540 1205 11570 1210
rect 11650 1230 11680 1235
rect 11650 1210 11655 1230
rect 11655 1210 11675 1230
rect 11675 1210 11680 1230
rect 11650 1205 11680 1210
rect 11760 1230 11790 1235
rect 11760 1210 11765 1230
rect 11765 1210 11785 1230
rect 11785 1210 11790 1230
rect 11760 1205 11790 1210
rect 11870 1230 11900 1235
rect 11870 1210 11875 1230
rect 11875 1210 11895 1230
rect 11895 1210 11900 1230
rect 11870 1205 11900 1210
rect 11980 1230 12010 1235
rect 11980 1210 11985 1230
rect 11985 1210 12005 1230
rect 12005 1210 12010 1230
rect 11980 1205 12010 1210
rect 12090 1230 12120 1235
rect 12090 1210 12095 1230
rect 12095 1210 12115 1230
rect 12115 1210 12120 1230
rect 12090 1205 12120 1210
rect 12200 1230 12230 1235
rect 12200 1210 12205 1230
rect 12205 1210 12225 1230
rect 12225 1210 12230 1230
rect 12200 1205 12230 1210
rect 12310 1230 12340 1235
rect 12310 1210 12315 1230
rect 12315 1210 12335 1230
rect 12335 1210 12340 1230
rect 12310 1205 12340 1210
rect 12420 1230 12450 1235
rect 12420 1210 12425 1230
rect 12425 1210 12445 1230
rect 12445 1210 12450 1230
rect 12420 1205 12450 1210
rect 12530 1230 12560 1235
rect 12530 1210 12535 1230
rect 12535 1210 12555 1230
rect 12555 1210 12560 1230
rect 12530 1205 12560 1210
rect 12600 1245 12630 1250
rect 12600 1225 12605 1245
rect 12605 1225 12625 1245
rect 12625 1225 12630 1245
rect 12600 1220 12630 1225
rect 12810 1220 12840 1250
rect 11170 910 11200 915
rect 11170 890 11175 910
rect 11175 890 11195 910
rect 11195 890 11200 910
rect 11170 885 11200 890
rect 11265 910 11295 915
rect 11265 890 11270 910
rect 11270 890 11290 910
rect 11290 890 11295 910
rect 11265 885 11295 890
rect 11375 910 11405 915
rect 11375 890 11380 910
rect 11380 890 11400 910
rect 11400 890 11405 910
rect 11375 885 11405 890
rect 11485 910 11515 915
rect 11485 890 11490 910
rect 11490 890 11510 910
rect 11510 890 11515 910
rect 11485 885 11515 890
rect 11595 910 11625 915
rect 11595 890 11600 910
rect 11600 890 11620 910
rect 11620 890 11625 910
rect 11595 885 11625 890
rect 11705 910 11735 915
rect 11705 890 11710 910
rect 11710 890 11730 910
rect 11730 890 11735 910
rect 11705 885 11735 890
rect 11815 910 11845 915
rect 11815 890 11820 910
rect 11820 890 11840 910
rect 11840 890 11845 910
rect 11815 885 11845 890
rect 11925 910 11955 915
rect 11925 890 11930 910
rect 11930 890 11950 910
rect 11950 890 11955 910
rect 11925 885 11955 890
rect 12035 910 12065 915
rect 12035 890 12040 910
rect 12040 890 12060 910
rect 12060 890 12065 910
rect 12035 885 12065 890
rect 12145 910 12175 915
rect 12145 890 12150 910
rect 12150 890 12170 910
rect 12170 890 12175 910
rect 12145 885 12175 890
rect 12255 910 12285 915
rect 12255 890 12260 910
rect 12260 890 12280 910
rect 12280 890 12285 910
rect 12255 885 12285 890
rect 12365 910 12395 915
rect 12365 890 12370 910
rect 12370 890 12390 910
rect 12390 890 12395 910
rect 12365 885 12395 890
rect 12475 910 12505 915
rect 12475 890 12480 910
rect 12480 890 12500 910
rect 12500 890 12505 910
rect 12475 885 12505 890
rect 12625 910 12655 915
rect 12625 890 12630 910
rect 12630 890 12650 910
rect 12650 890 12655 910
rect 12625 885 12655 890
rect 11010 825 11040 855
rect 11500 825 11530 855
rect 11940 830 11970 860
rect 12160 830 12190 860
rect 12380 830 12410 860
rect 13005 3630 13035 3635
rect 13005 3610 13010 3630
rect 13010 3610 13030 3630
rect 13030 3610 13035 3630
rect 13005 3605 13035 3610
rect 13115 3630 13145 3635
rect 13115 3610 13120 3630
rect 13120 3610 13140 3630
rect 13140 3610 13145 3630
rect 13115 3605 13145 3610
rect 13225 3630 13255 3635
rect 13225 3610 13230 3630
rect 13230 3610 13250 3630
rect 13250 3610 13255 3630
rect 13225 3605 13255 3610
rect 13335 3630 13365 3635
rect 13335 3610 13340 3630
rect 13340 3610 13360 3630
rect 13360 3610 13365 3630
rect 13335 3605 13365 3610
rect 13445 3630 13475 3635
rect 13445 3610 13450 3630
rect 13450 3610 13470 3630
rect 13470 3610 13475 3630
rect 13445 3605 13475 3610
rect 13555 3630 13585 3635
rect 13555 3610 13560 3630
rect 13560 3610 13580 3630
rect 13580 3610 13585 3630
rect 13555 3605 13585 3610
rect 26345 3620 26375 3625
rect 26345 3600 26350 3620
rect 26350 3600 26370 3620
rect 26370 3600 26375 3620
rect 26345 3595 26375 3600
rect 26465 3620 26495 3625
rect 26465 3600 26470 3620
rect 26470 3600 26490 3620
rect 26490 3600 26495 3620
rect 26465 3595 26495 3600
rect 26585 3620 26615 3625
rect 26585 3600 26590 3620
rect 26590 3600 26610 3620
rect 26610 3600 26615 3620
rect 26585 3595 26615 3600
rect 26705 3620 26735 3625
rect 26705 3600 26710 3620
rect 26710 3600 26730 3620
rect 26730 3600 26735 3620
rect 26705 3595 26735 3600
rect 26825 3620 26855 3625
rect 26825 3600 26830 3620
rect 26830 3600 26850 3620
rect 26850 3600 26855 3620
rect 26825 3595 26855 3600
rect 26945 3620 26975 3625
rect 26945 3600 26950 3620
rect 26950 3600 26970 3620
rect 26970 3600 26975 3620
rect 26945 3595 26975 3600
rect 27065 3620 27095 3625
rect 27065 3600 27070 3620
rect 27070 3600 27090 3620
rect 27090 3600 27095 3620
rect 27065 3595 27095 3600
rect 27185 3620 27215 3625
rect 27185 3600 27190 3620
rect 27190 3600 27210 3620
rect 27210 3600 27215 3620
rect 27185 3595 27215 3600
rect 27305 3620 27335 3625
rect 27305 3600 27310 3620
rect 27310 3600 27330 3620
rect 27330 3600 27335 3620
rect 27305 3595 27335 3600
rect 27425 3620 27455 3625
rect 27425 3600 27430 3620
rect 27430 3600 27450 3620
rect 27450 3600 27455 3620
rect 27425 3595 27455 3600
rect 13765 3525 13795 3555
rect 13815 3525 13845 3555
rect 13865 3525 13895 3555
rect 27950 3285 27980 3290
rect 27950 3265 27955 3285
rect 27955 3265 27975 3285
rect 27975 3265 27980 3285
rect 27950 3260 27980 3265
rect 28060 3285 28090 3290
rect 28060 3265 28065 3285
rect 28065 3265 28085 3285
rect 28085 3265 28090 3285
rect 28060 3260 28090 3265
rect 28170 3285 28200 3290
rect 28170 3265 28175 3285
rect 28175 3265 28195 3285
rect 28195 3265 28200 3285
rect 28170 3260 28200 3265
rect 28280 3285 28310 3290
rect 28280 3265 28285 3285
rect 28285 3265 28305 3285
rect 28305 3265 28310 3285
rect 28280 3260 28310 3265
rect 28390 3285 28420 3290
rect 28390 3265 28395 3285
rect 28395 3265 28415 3285
rect 28415 3265 28420 3285
rect 28390 3260 28420 3265
rect 28500 3285 28530 3290
rect 28500 3265 28505 3285
rect 28505 3265 28525 3285
rect 28525 3265 28530 3285
rect 28500 3260 28530 3265
rect 28610 3285 28640 3290
rect 28610 3265 28615 3285
rect 28615 3265 28635 3285
rect 28635 3265 28640 3285
rect 28610 3260 28640 3265
rect 28720 3285 28750 3290
rect 28720 3265 28725 3285
rect 28725 3265 28745 3285
rect 28745 3265 28750 3285
rect 28720 3260 28750 3265
rect 28830 3285 28860 3290
rect 28830 3265 28835 3285
rect 28835 3265 28855 3285
rect 28855 3265 28860 3285
rect 28830 3260 28860 3265
rect 28940 3285 28970 3290
rect 28940 3265 28945 3285
rect 28945 3265 28965 3285
rect 28965 3265 28970 3285
rect 28940 3260 28970 3265
rect 29050 3285 29080 3290
rect 29050 3265 29055 3285
rect 29055 3265 29075 3285
rect 29075 3265 29080 3285
rect 29050 3260 29080 3265
rect 25585 3205 25615 3210
rect 25585 3185 25590 3205
rect 25590 3185 25610 3205
rect 25610 3185 25615 3205
rect 25585 3180 25615 3185
rect 25985 3205 26015 3210
rect 25985 3185 25990 3205
rect 25990 3185 26010 3205
rect 26010 3185 26015 3205
rect 25985 3180 26015 3185
rect 25905 3125 25935 3155
rect 13060 2960 13090 2965
rect 13060 2940 13065 2960
rect 13065 2940 13085 2960
rect 13085 2940 13090 2960
rect 13060 2935 13090 2940
rect 13170 2960 13200 2965
rect 13170 2940 13175 2960
rect 13175 2940 13195 2960
rect 13195 2940 13200 2960
rect 13170 2935 13200 2940
rect 13280 2960 13310 2965
rect 13280 2940 13285 2960
rect 13285 2940 13305 2960
rect 13305 2940 13310 2960
rect 13280 2935 13310 2940
rect 13390 2960 13420 2965
rect 13390 2940 13395 2960
rect 13395 2940 13415 2960
rect 13415 2940 13420 2960
rect 13390 2935 13420 2940
rect 13500 2960 13530 2965
rect 13500 2940 13505 2960
rect 13505 2940 13525 2960
rect 13525 2940 13530 2960
rect 13500 2935 13530 2940
rect 13115 2850 13145 2880
rect 13765 2905 13795 2935
rect 13815 2905 13845 2935
rect 13865 2905 13895 2935
rect 13815 2850 13845 2880
rect 13390 2795 13420 2825
rect 14020 2795 14050 2825
rect 13005 2700 13035 2705
rect 13005 2680 13010 2700
rect 13010 2680 13030 2700
rect 13030 2680 13035 2700
rect 13005 2675 13035 2680
rect 13115 2700 13145 2705
rect 13115 2680 13120 2700
rect 13120 2680 13140 2700
rect 13140 2680 13145 2700
rect 13115 2675 13145 2680
rect 13225 2700 13255 2705
rect 13225 2680 13230 2700
rect 13230 2680 13250 2700
rect 13250 2680 13255 2700
rect 13225 2675 13255 2680
rect 13335 2700 13365 2705
rect 13335 2680 13340 2700
rect 13340 2680 13360 2700
rect 13360 2680 13365 2700
rect 13335 2675 13365 2680
rect 13445 2700 13475 2705
rect 13445 2680 13450 2700
rect 13450 2680 13470 2700
rect 13470 2680 13475 2700
rect 13445 2675 13475 2680
rect 13555 2700 13585 2705
rect 13555 2680 13560 2700
rect 13560 2680 13580 2700
rect 13580 2680 13585 2700
rect 13555 2675 13585 2680
rect 13060 2430 13090 2435
rect 13060 2410 13065 2430
rect 13065 2410 13085 2430
rect 13085 2410 13090 2430
rect 13060 2405 13090 2410
rect 13170 2430 13200 2435
rect 13170 2410 13175 2430
rect 13175 2410 13195 2430
rect 13195 2410 13200 2430
rect 13170 2405 13200 2410
rect 13280 2430 13310 2435
rect 13280 2410 13285 2430
rect 13285 2410 13305 2430
rect 13305 2410 13310 2430
rect 13280 2405 13310 2410
rect 13390 2430 13420 2435
rect 13390 2410 13395 2430
rect 13395 2410 13415 2430
rect 13415 2410 13420 2430
rect 13390 2405 13420 2410
rect 13500 2430 13530 2435
rect 13500 2410 13505 2430
rect 13505 2410 13525 2430
rect 13525 2410 13530 2430
rect 13500 2405 13530 2410
rect 13745 2405 13775 2435
rect 13030 2370 13060 2375
rect 13030 2350 13035 2370
rect 13035 2350 13055 2370
rect 13055 2350 13060 2370
rect 13030 2345 13060 2350
rect 13060 2310 13090 2315
rect 13060 2290 13065 2310
rect 13065 2290 13085 2310
rect 13085 2290 13090 2310
rect 13060 2285 13090 2290
rect 13170 2310 13200 2315
rect 13170 2290 13175 2310
rect 13175 2290 13195 2310
rect 13195 2290 13200 2310
rect 13170 2285 13200 2290
rect 13280 2310 13310 2315
rect 13280 2290 13285 2310
rect 13285 2290 13305 2310
rect 13305 2290 13310 2310
rect 13280 2285 13310 2290
rect 13390 2310 13420 2315
rect 13390 2290 13395 2310
rect 13395 2290 13415 2310
rect 13415 2290 13420 2310
rect 13390 2285 13420 2290
rect 13500 2310 13530 2315
rect 13500 2290 13505 2310
rect 13505 2290 13525 2310
rect 13525 2290 13530 2310
rect 13500 2285 13530 2290
rect 13700 2285 13730 2315
rect 13745 1970 13775 2000
rect 13795 2000 13830 2005
rect 13795 1975 13800 2000
rect 13800 1975 13825 2000
rect 13825 1975 13830 2000
rect 13795 1970 13830 1975
rect 13855 2000 13890 2005
rect 13855 1975 13860 2000
rect 13860 1975 13885 2000
rect 13885 1975 13890 2000
rect 13855 1970 13890 1975
rect 13915 2000 13950 2005
rect 13915 1975 13920 2000
rect 13920 1975 13945 2000
rect 13945 1975 13950 2000
rect 13915 1970 13950 1975
rect 13975 2000 14010 2005
rect 13975 1975 13980 2000
rect 13980 1975 14005 2000
rect 14005 1975 14010 2000
rect 13975 1970 14010 1975
rect 13005 1940 13035 1945
rect 13005 1920 13012 1940
rect 13012 1920 13030 1940
rect 13030 1920 13035 1940
rect 13005 1915 13035 1920
rect 13115 1940 13145 1945
rect 13115 1920 13122 1940
rect 13122 1920 13140 1940
rect 13140 1920 13145 1940
rect 13115 1915 13145 1920
rect 13225 1940 13255 1945
rect 13225 1920 13232 1940
rect 13232 1920 13250 1940
rect 13250 1920 13255 1940
rect 13225 1915 13255 1920
rect 13335 1940 13365 1945
rect 13335 1920 13342 1940
rect 13342 1920 13360 1940
rect 13360 1920 13365 1940
rect 13335 1915 13365 1920
rect 13445 1940 13475 1945
rect 13445 1920 13452 1940
rect 13452 1920 13470 1940
rect 13470 1920 13475 1940
rect 13445 1915 13475 1920
rect 13555 1940 13585 1945
rect 13555 1920 13562 1940
rect 13562 1920 13580 1940
rect 13580 1920 13585 1940
rect 13555 1915 13585 1920
rect 13700 1915 13730 1945
rect 13855 1915 13885 1945
rect 13975 1865 14005 1895
rect 13210 1730 13240 1760
rect 13800 1730 13830 1760
rect 12930 1675 12960 1705
rect 13110 1700 13140 1705
rect 13110 1680 13115 1700
rect 13115 1680 13135 1700
rect 13135 1680 13140 1700
rect 13110 1675 13140 1680
rect 13310 1700 13340 1705
rect 13310 1680 13315 1700
rect 13315 1680 13335 1700
rect 13335 1680 13340 1700
rect 13310 1675 13340 1680
rect 13510 1700 13540 1705
rect 13510 1680 13515 1700
rect 13515 1680 13535 1700
rect 13535 1680 13540 1700
rect 13510 1675 13540 1680
rect 13735 1675 13765 1705
rect 24740 2665 24770 2670
rect 24740 2645 24745 2665
rect 24745 2645 24765 2665
rect 24765 2645 24770 2665
rect 24740 2640 24770 2645
rect 24850 2665 24880 2670
rect 24850 2645 24855 2665
rect 24855 2645 24875 2665
rect 24875 2645 24880 2665
rect 24850 2640 24880 2645
rect 24960 2665 24990 2670
rect 24960 2645 24965 2665
rect 24965 2645 24985 2665
rect 24985 2645 24990 2665
rect 24960 2640 24990 2645
rect 25070 2665 25100 2670
rect 25070 2645 25075 2665
rect 25075 2645 25095 2665
rect 25095 2645 25100 2665
rect 25070 2640 25100 2645
rect 25180 2665 25210 2670
rect 25180 2645 25185 2665
rect 25185 2645 25205 2665
rect 25205 2645 25210 2665
rect 25180 2640 25210 2645
rect 25290 2665 25320 2670
rect 25290 2645 25295 2665
rect 25295 2645 25315 2665
rect 25315 2645 25320 2665
rect 25290 2640 25320 2645
rect 25400 2665 25430 2670
rect 25400 2645 25405 2665
rect 25405 2645 25425 2665
rect 25425 2645 25430 2665
rect 25400 2640 25430 2645
rect 25510 2665 25540 2670
rect 25510 2645 25515 2665
rect 25515 2645 25535 2665
rect 25535 2645 25540 2665
rect 25510 2640 25540 2645
rect 25620 2665 25650 2670
rect 25620 2645 25625 2665
rect 25625 2645 25645 2665
rect 25645 2645 25650 2665
rect 25620 2640 25650 2645
rect 25730 2665 25760 2670
rect 25730 2645 25735 2665
rect 25735 2645 25755 2665
rect 25755 2645 25760 2665
rect 25730 2640 25760 2645
rect 25840 2665 25870 2670
rect 25840 2645 25845 2665
rect 25845 2645 25865 2665
rect 25865 2645 25870 2665
rect 25840 2640 25870 2645
rect 24795 2495 24825 2500
rect 24795 2475 24800 2495
rect 24800 2475 24820 2495
rect 24820 2475 24825 2495
rect 24795 2470 24825 2475
rect 24905 2495 24935 2500
rect 24905 2475 24910 2495
rect 24910 2475 24930 2495
rect 24930 2475 24935 2495
rect 24905 2470 24935 2475
rect 25015 2495 25045 2500
rect 25015 2475 25020 2495
rect 25020 2475 25040 2495
rect 25040 2475 25045 2495
rect 25015 2470 25045 2475
rect 25125 2495 25155 2500
rect 25125 2475 25130 2495
rect 25130 2475 25150 2495
rect 25150 2475 25155 2495
rect 25125 2470 25155 2475
rect 25235 2495 25265 2500
rect 25235 2475 25240 2495
rect 25240 2475 25260 2495
rect 25260 2475 25265 2495
rect 25235 2470 25265 2475
rect 25345 2495 25375 2500
rect 25345 2475 25350 2495
rect 25350 2475 25370 2495
rect 25370 2475 25375 2495
rect 25345 2470 25375 2475
rect 25455 2495 25485 2500
rect 25455 2475 25460 2495
rect 25460 2475 25480 2495
rect 25480 2475 25485 2495
rect 25455 2470 25485 2475
rect 25565 2495 25595 2500
rect 25565 2475 25570 2495
rect 25570 2475 25590 2495
rect 25590 2475 25595 2495
rect 25565 2470 25595 2475
rect 25675 2495 25705 2500
rect 25675 2475 25680 2495
rect 25680 2475 25700 2495
rect 25700 2475 25705 2495
rect 25675 2470 25705 2475
rect 25785 2495 25815 2500
rect 25785 2475 25790 2495
rect 25790 2475 25810 2495
rect 25810 2475 25815 2495
rect 25785 2470 25815 2475
rect 26826 3150 26854 3155
rect 26826 3130 26831 3150
rect 26831 3130 26849 3150
rect 26849 3130 26854 3150
rect 26826 3125 26854 3130
rect 26285 3070 26315 3100
rect 26525 3070 26555 3100
rect 26765 3070 26795 3100
rect 27005 3070 27035 3100
rect 27245 3070 27275 3100
rect 27485 3070 27515 3100
rect 26405 3025 26435 3055
rect 26645 3025 26675 3055
rect 26885 3025 26915 3055
rect 27125 3025 27155 3055
rect 27365 3025 27395 3055
rect 26345 2970 26375 3000
rect 26405 2970 26435 3000
rect 26585 2970 26615 3000
rect 26825 2970 26855 3000
rect 27065 2970 27095 3000
rect 27305 2970 27335 3000
rect 26465 2940 26495 2945
rect 26465 2920 26470 2940
rect 26470 2920 26490 2940
rect 26490 2920 26495 2940
rect 26465 2915 26495 2920
rect 26705 2940 26735 2945
rect 26705 2920 26710 2940
rect 26710 2920 26730 2940
rect 26730 2920 26735 2940
rect 26705 2915 26735 2920
rect 26945 2940 26975 2945
rect 26945 2920 26950 2940
rect 26950 2920 26970 2940
rect 26970 2920 26975 2940
rect 26945 2915 26975 2920
rect 27185 2940 27215 2945
rect 27185 2920 27190 2940
rect 27190 2920 27210 2940
rect 27210 2920 27215 2940
rect 27185 2915 27215 2920
rect 27425 2940 27455 2945
rect 27425 2920 27430 2940
rect 27430 2920 27450 2940
rect 27450 2920 27455 2940
rect 27425 2915 27455 2920
rect 27485 2915 27515 2945
rect 28005 2915 28035 2920
rect 28005 2895 28010 2915
rect 28010 2895 28030 2915
rect 28030 2895 28035 2915
rect 28005 2890 28035 2895
rect 28115 2915 28145 2920
rect 28115 2895 28120 2915
rect 28120 2895 28140 2915
rect 28140 2895 28145 2915
rect 28115 2890 28145 2895
rect 28225 2915 28255 2920
rect 28225 2895 28230 2915
rect 28230 2895 28250 2915
rect 28250 2895 28255 2915
rect 28225 2890 28255 2895
rect 28335 2915 28365 2920
rect 28335 2895 28340 2915
rect 28340 2895 28360 2915
rect 28360 2895 28365 2915
rect 28335 2890 28365 2895
rect 28445 2915 28475 2920
rect 28445 2895 28450 2915
rect 28450 2895 28470 2915
rect 28470 2895 28475 2915
rect 28445 2890 28475 2895
rect 28555 2915 28585 2920
rect 28555 2895 28560 2915
rect 28560 2895 28580 2915
rect 28580 2895 28585 2915
rect 28555 2890 28585 2895
rect 28665 2915 28695 2920
rect 28665 2895 28670 2915
rect 28670 2895 28690 2915
rect 28690 2895 28695 2915
rect 28665 2890 28695 2895
rect 28775 2915 28805 2920
rect 28775 2895 28780 2915
rect 28780 2895 28800 2915
rect 28800 2895 28805 2915
rect 28775 2890 28805 2895
rect 28885 2915 28915 2920
rect 28885 2895 28890 2915
rect 28890 2895 28910 2915
rect 28910 2895 28915 2915
rect 28885 2890 28915 2895
rect 28995 2915 29025 2920
rect 28995 2895 29000 2915
rect 29000 2895 29020 2915
rect 29020 2895 29025 2915
rect 28995 2890 29025 2895
rect 28060 2800 28090 2830
rect 28060 2750 28090 2780
rect 27695 2700 27725 2730
rect 28060 2700 28090 2730
rect 25985 2445 26015 2475
rect 26826 2470 26854 2475
rect 26826 2450 26831 2470
rect 26831 2450 26849 2470
rect 26849 2450 26854 2470
rect 26826 2445 26854 2450
rect 25816 2435 25844 2440
rect 25816 2415 25821 2435
rect 25821 2415 25839 2435
rect 25839 2415 25844 2435
rect 25816 2410 25844 2415
rect 24805 2375 24840 2380
rect 24805 2350 24810 2375
rect 24810 2350 24835 2375
rect 24835 2350 24840 2375
rect 24805 2345 24840 2350
rect 25640 2375 25675 2380
rect 25640 2350 25645 2375
rect 25645 2350 25670 2375
rect 25670 2350 25675 2375
rect 25640 2345 25675 2350
rect 24805 2315 24840 2320
rect 24805 2290 24810 2315
rect 24810 2290 24835 2315
rect 24835 2290 24840 2315
rect 24805 2285 24840 2290
rect 25640 2315 25675 2320
rect 25640 2290 25645 2315
rect 25645 2290 25670 2315
rect 25670 2290 25675 2315
rect 25640 2285 25675 2290
rect 26285 2390 26315 2420
rect 26525 2390 26555 2420
rect 26765 2390 26795 2420
rect 26405 2345 26435 2375
rect 26645 2345 26675 2375
rect 25816 2275 25844 2280
rect 25816 2255 25821 2275
rect 25821 2255 25839 2275
rect 25839 2255 25844 2275
rect 25816 2250 25844 2255
rect 26445 2250 26475 2280
rect 26665 2250 26695 2280
rect 24795 2215 24825 2220
rect 24795 2195 24800 2215
rect 24800 2195 24820 2215
rect 24820 2195 24825 2215
rect 24795 2190 24825 2195
rect 24905 2215 24935 2220
rect 24905 2195 24910 2215
rect 24910 2195 24930 2215
rect 24930 2195 24935 2215
rect 24905 2190 24935 2195
rect 25015 2215 25045 2220
rect 25015 2195 25020 2215
rect 25020 2195 25040 2215
rect 25040 2195 25045 2215
rect 25015 2190 25045 2195
rect 25125 2215 25155 2220
rect 25125 2195 25130 2215
rect 25130 2195 25150 2215
rect 25150 2195 25155 2215
rect 25125 2190 25155 2195
rect 25235 2215 25265 2220
rect 25235 2195 25240 2215
rect 25240 2195 25260 2215
rect 25260 2195 25265 2215
rect 25235 2190 25265 2195
rect 25345 2215 25375 2220
rect 25345 2195 25350 2215
rect 25350 2195 25370 2215
rect 25370 2195 25375 2215
rect 25345 2190 25375 2195
rect 25455 2215 25485 2220
rect 25455 2195 25460 2215
rect 25460 2195 25480 2215
rect 25480 2195 25485 2215
rect 25455 2190 25485 2195
rect 25565 2215 25595 2220
rect 25565 2195 25570 2215
rect 25570 2195 25590 2215
rect 25590 2195 25595 2215
rect 25565 2190 25595 2195
rect 25675 2215 25705 2220
rect 25675 2195 25680 2215
rect 25680 2195 25700 2215
rect 25700 2195 25705 2215
rect 25675 2190 25705 2195
rect 25785 2215 25815 2220
rect 25785 2195 25790 2215
rect 25790 2195 25810 2215
rect 25810 2195 25815 2215
rect 25785 2190 25815 2195
rect 26335 2205 26365 2235
rect 26555 2205 26585 2235
rect 27005 2390 27035 2420
rect 27245 2390 27275 2420
rect 27485 2390 27515 2420
rect 27950 2665 27980 2670
rect 27950 2645 27955 2665
rect 27955 2645 27975 2665
rect 27975 2645 27980 2665
rect 27950 2640 27980 2645
rect 28060 2665 28090 2670
rect 28060 2645 28065 2665
rect 28065 2645 28085 2665
rect 28085 2645 28090 2665
rect 28060 2640 28090 2645
rect 28170 2665 28200 2670
rect 28170 2645 28175 2665
rect 28175 2645 28195 2665
rect 28195 2645 28200 2665
rect 28170 2640 28200 2645
rect 28280 2665 28310 2670
rect 28280 2645 28285 2665
rect 28285 2645 28305 2665
rect 28305 2645 28310 2665
rect 28280 2640 28310 2645
rect 28390 2665 28420 2670
rect 28390 2645 28395 2665
rect 28395 2645 28415 2665
rect 28415 2645 28420 2665
rect 28390 2640 28420 2645
rect 28500 2665 28530 2670
rect 28500 2645 28505 2665
rect 28505 2645 28525 2665
rect 28525 2645 28530 2665
rect 28500 2640 28530 2645
rect 28610 2665 28640 2670
rect 28610 2645 28615 2665
rect 28615 2645 28635 2665
rect 28635 2645 28640 2665
rect 28610 2640 28640 2645
rect 28720 2665 28750 2670
rect 28720 2645 28725 2665
rect 28725 2645 28745 2665
rect 28745 2645 28750 2665
rect 28720 2640 28750 2645
rect 28830 2665 28860 2670
rect 28830 2645 28835 2665
rect 28835 2645 28855 2665
rect 28855 2645 28860 2665
rect 28830 2640 28860 2645
rect 28940 2665 28970 2670
rect 28940 2645 28945 2665
rect 28945 2645 28965 2665
rect 28965 2645 28970 2665
rect 28940 2640 28970 2645
rect 29050 2665 29080 2670
rect 29050 2645 29055 2665
rect 29055 2645 29075 2665
rect 29075 2645 29080 2665
rect 29050 2640 29080 2645
rect 28005 2495 28035 2500
rect 28005 2475 28010 2495
rect 28010 2475 28030 2495
rect 28030 2475 28035 2495
rect 28005 2470 28035 2475
rect 28115 2495 28145 2500
rect 28115 2475 28120 2495
rect 28120 2475 28140 2495
rect 28140 2475 28145 2495
rect 28115 2470 28145 2475
rect 28225 2495 28255 2500
rect 28225 2475 28230 2495
rect 28230 2475 28250 2495
rect 28250 2475 28255 2495
rect 28225 2470 28255 2475
rect 28335 2495 28365 2500
rect 28335 2475 28340 2495
rect 28340 2475 28360 2495
rect 28360 2475 28365 2495
rect 28335 2470 28365 2475
rect 28445 2495 28475 2500
rect 28445 2475 28450 2495
rect 28450 2475 28470 2495
rect 28470 2475 28475 2495
rect 28445 2470 28475 2475
rect 28555 2495 28585 2500
rect 28555 2475 28560 2495
rect 28560 2475 28580 2495
rect 28580 2475 28585 2495
rect 28555 2470 28585 2475
rect 28665 2495 28695 2500
rect 28665 2475 28670 2495
rect 28670 2475 28690 2495
rect 28690 2475 28695 2495
rect 28665 2470 28695 2475
rect 28775 2495 28805 2500
rect 28775 2475 28780 2495
rect 28780 2475 28800 2495
rect 28800 2475 28805 2495
rect 28775 2470 28805 2475
rect 28885 2495 28915 2500
rect 28885 2475 28890 2495
rect 28890 2475 28910 2495
rect 28910 2475 28915 2495
rect 28885 2470 28915 2475
rect 28995 2495 29025 2500
rect 28995 2475 29000 2495
rect 29000 2475 29020 2495
rect 29020 2475 29025 2495
rect 28995 2470 29025 2475
rect 27976 2435 28004 2440
rect 27976 2415 27981 2435
rect 27981 2415 27999 2435
rect 27999 2415 28004 2435
rect 27976 2410 28004 2415
rect 26885 2345 26915 2375
rect 27125 2345 27155 2375
rect 27365 2345 27395 2375
rect 27695 2345 27725 2375
rect 27975 2345 28005 2375
rect 28145 2375 28180 2380
rect 28145 2350 28150 2375
rect 28150 2350 28175 2375
rect 28175 2350 28180 2375
rect 28145 2345 28180 2350
rect 28980 2375 29015 2380
rect 28980 2350 28985 2375
rect 28985 2350 29010 2375
rect 29010 2350 29015 2375
rect 28980 2345 29015 2350
rect 27820 2295 27850 2325
rect 26885 2250 26915 2280
rect 27105 2250 27135 2280
rect 27325 2250 27355 2280
rect 26775 2205 26805 2235
rect 26995 2205 27025 2235
rect 27215 2205 27245 2235
rect 27435 2205 27465 2235
rect 24740 1995 24770 2000
rect 24740 1975 24745 1995
rect 24745 1975 24763 1995
rect 24763 1975 24770 1995
rect 24740 1970 24770 1975
rect 24850 1995 24880 2000
rect 24850 1975 24855 1995
rect 24855 1975 24873 1995
rect 24873 1975 24880 1995
rect 24850 1970 24880 1975
rect 24960 1995 24990 2000
rect 24960 1975 24965 1995
rect 24965 1975 24983 1995
rect 24983 1975 24990 1995
rect 24960 1970 24990 1975
rect 25070 1995 25100 2000
rect 25070 1975 25075 1995
rect 25075 1975 25093 1995
rect 25093 1975 25100 1995
rect 25070 1970 25100 1975
rect 25180 1995 25210 2000
rect 25180 1975 25185 1995
rect 25185 1975 25203 1995
rect 25203 1975 25210 1995
rect 25180 1970 25210 1975
rect 25290 1995 25320 2000
rect 25290 1975 25295 1995
rect 25295 1975 25313 1995
rect 25313 1975 25320 1995
rect 25290 1970 25320 1975
rect 25400 1995 25430 2000
rect 25400 1975 25405 1995
rect 25405 1975 25423 1995
rect 25423 1975 25430 1995
rect 25400 1970 25430 1975
rect 25510 1995 25540 2000
rect 25510 1975 25515 1995
rect 25515 1975 25533 1995
rect 25533 1975 25540 1995
rect 25510 1970 25540 1975
rect 25620 1995 25650 2000
rect 25620 1975 25625 1995
rect 25625 1975 25643 1995
rect 25643 1975 25650 1995
rect 25620 1970 25650 1975
rect 25730 1995 25760 2000
rect 25730 1975 25735 1995
rect 25735 1975 25753 1995
rect 25753 1975 25760 1995
rect 25730 1970 25760 1975
rect 25840 1995 25870 2000
rect 25840 1975 25845 1995
rect 25845 1975 25863 1995
rect 25863 1975 25870 1995
rect 25840 1970 25870 1975
rect 26390 1955 26420 1960
rect 26390 1935 26395 1955
rect 26395 1935 26415 1955
rect 26415 1935 26420 1955
rect 26390 1930 26420 1935
rect 26610 1955 26640 1960
rect 26610 1935 26615 1955
rect 26615 1935 26635 1955
rect 26635 1935 26640 1955
rect 26610 1930 26640 1935
rect 26830 1955 26860 1960
rect 26830 1935 26835 1955
rect 26835 1935 26855 1955
rect 26855 1935 26860 1955
rect 26830 1930 26860 1935
rect 27050 1955 27080 1960
rect 27050 1935 27055 1955
rect 27055 1935 27075 1955
rect 27075 1935 27080 1955
rect 27050 1930 27080 1935
rect 27270 1955 27300 1960
rect 27270 1935 27275 1955
rect 27275 1935 27295 1955
rect 27295 1935 27300 1955
rect 27270 1930 27300 1935
rect 26500 1875 26530 1905
rect 26720 1875 26750 1905
rect 26940 1875 26970 1905
rect 27160 1875 27190 1905
rect 26195 1820 26225 1850
rect 26415 1820 26445 1850
rect 26090 1755 26120 1760
rect 26090 1735 26095 1755
rect 26095 1735 26115 1755
rect 26115 1735 26120 1755
rect 26090 1730 26120 1735
rect 26310 1755 26340 1760
rect 26310 1735 26315 1755
rect 26315 1735 26335 1755
rect 26335 1735 26340 1755
rect 26310 1730 26340 1735
rect 27380 1875 27410 1905
rect 26645 1820 26675 1850
rect 27235 1820 27265 1850
rect 27455 1820 27485 1850
rect 27685 1820 27715 1850
rect 26825 1775 26855 1805
rect 26945 1775 26975 1805
rect 26530 1755 26560 1760
rect 26530 1735 26535 1755
rect 26535 1735 26555 1755
rect 26555 1735 26560 1755
rect 26530 1730 26560 1735
rect 27130 1755 27160 1760
rect 27130 1735 27135 1755
rect 27135 1735 27155 1755
rect 27155 1735 27160 1755
rect 27130 1730 27160 1735
rect 27350 1755 27380 1760
rect 27350 1735 27355 1755
rect 27355 1735 27375 1755
rect 27375 1735 27380 1755
rect 27350 1730 27380 1735
rect 27570 1755 27600 1760
rect 27570 1735 27575 1755
rect 27575 1735 27595 1755
rect 27595 1735 27600 1755
rect 27570 1730 27600 1735
rect 14020 1675 14050 1705
rect 26240 1710 26266 1715
rect 26240 1690 26243 1710
rect 26243 1690 26260 1710
rect 26260 1690 26266 1710
rect 26240 1685 26266 1690
rect 26460 1710 26486 1715
rect 26460 1690 26463 1710
rect 26463 1690 26480 1710
rect 26480 1690 26486 1710
rect 26460 1685 26486 1690
rect 26604 1710 26630 1715
rect 26604 1690 26610 1710
rect 26610 1690 26627 1710
rect 26627 1690 26630 1710
rect 26604 1685 26630 1690
rect 26870 1710 26896 1715
rect 26870 1690 26876 1710
rect 26876 1690 26893 1710
rect 26893 1690 26896 1710
rect 26870 1685 26896 1690
rect 27280 1710 27306 1715
rect 27280 1690 27283 1710
rect 27283 1690 27300 1710
rect 27300 1690 27306 1710
rect 27280 1685 27306 1690
rect 27500 1710 27526 1715
rect 27500 1690 27503 1710
rect 27503 1690 27520 1710
rect 27520 1690 27526 1710
rect 27500 1685 27526 1690
rect 27644 1710 27670 1715
rect 27644 1690 27650 1710
rect 27650 1690 27667 1710
rect 27667 1690 27670 1710
rect 27644 1685 27670 1690
rect 13735 1640 13770 1645
rect 13735 1615 13740 1640
rect 13740 1615 13765 1640
rect 13765 1615 13770 1640
rect 13735 1610 13770 1615
rect 13795 1640 13830 1645
rect 13795 1615 13800 1640
rect 13800 1615 13825 1640
rect 13825 1615 13830 1640
rect 13795 1610 13830 1615
rect 28145 2315 28180 2320
rect 28145 2290 28150 2315
rect 28150 2290 28175 2315
rect 28175 2290 28180 2315
rect 28145 2285 28180 2290
rect 28980 2315 29015 2320
rect 28980 2290 28985 2315
rect 28985 2290 29010 2315
rect 29010 2290 29015 2315
rect 28980 2285 29015 2290
rect 27976 2275 28004 2280
rect 27976 2255 27981 2275
rect 27981 2255 27999 2275
rect 27999 2255 28004 2275
rect 27976 2250 28004 2255
rect 28005 2215 28035 2220
rect 28005 2195 28010 2215
rect 28010 2195 28030 2215
rect 28030 2195 28035 2215
rect 28005 2190 28035 2195
rect 28115 2215 28145 2220
rect 28115 2195 28120 2215
rect 28120 2195 28140 2215
rect 28140 2195 28145 2215
rect 28115 2190 28145 2195
rect 28225 2215 28255 2220
rect 28225 2195 28230 2215
rect 28230 2195 28250 2215
rect 28250 2195 28255 2215
rect 28225 2190 28255 2195
rect 28335 2215 28365 2220
rect 28335 2195 28340 2215
rect 28340 2195 28360 2215
rect 28360 2195 28365 2215
rect 28335 2190 28365 2195
rect 28445 2215 28475 2220
rect 28445 2195 28450 2215
rect 28450 2195 28470 2215
rect 28470 2195 28475 2215
rect 28445 2190 28475 2195
rect 28555 2215 28585 2220
rect 28555 2195 28560 2215
rect 28560 2195 28580 2215
rect 28580 2195 28585 2215
rect 28555 2190 28585 2195
rect 28665 2215 28695 2220
rect 28665 2195 28670 2215
rect 28670 2195 28690 2215
rect 28690 2195 28695 2215
rect 28665 2190 28695 2195
rect 28775 2215 28805 2220
rect 28775 2195 28780 2215
rect 28780 2195 28800 2215
rect 28800 2195 28805 2215
rect 28775 2190 28805 2195
rect 28885 2215 28915 2220
rect 28885 2195 28890 2215
rect 28890 2195 28910 2215
rect 28910 2195 28915 2215
rect 28885 2190 28915 2195
rect 28995 2215 29025 2220
rect 28995 2195 29000 2215
rect 29000 2195 29020 2215
rect 29020 2195 29025 2215
rect 28995 2190 29025 2195
rect 27950 1995 27980 2000
rect 27950 1975 27957 1995
rect 27957 1975 27975 1995
rect 27975 1975 27980 1995
rect 27950 1970 27980 1975
rect 28060 1995 28090 2000
rect 28060 1975 28067 1995
rect 28067 1975 28085 1995
rect 28085 1975 28090 1995
rect 28060 1970 28090 1975
rect 28170 1995 28200 2000
rect 28170 1975 28177 1995
rect 28177 1975 28195 1995
rect 28195 1975 28200 1995
rect 28170 1970 28200 1975
rect 28280 1995 28310 2000
rect 28280 1975 28287 1995
rect 28287 1975 28305 1995
rect 28305 1975 28310 1995
rect 28280 1970 28310 1975
rect 28390 1995 28420 2000
rect 28390 1975 28397 1995
rect 28397 1975 28415 1995
rect 28415 1975 28420 1995
rect 28390 1970 28420 1975
rect 28500 1995 28530 2000
rect 28500 1975 28507 1995
rect 28507 1975 28525 1995
rect 28525 1975 28530 1995
rect 28500 1970 28530 1975
rect 28610 1995 28640 2000
rect 28610 1975 28617 1995
rect 28617 1975 28635 1995
rect 28635 1975 28640 1995
rect 28610 1970 28640 1975
rect 28720 1995 28750 2000
rect 28720 1975 28727 1995
rect 28727 1975 28745 1995
rect 28745 1975 28750 1995
rect 28720 1970 28750 1975
rect 28830 1995 28860 2000
rect 28830 1975 28837 1995
rect 28837 1975 28855 1995
rect 28855 1975 28860 1995
rect 28830 1970 28860 1975
rect 28940 1995 28970 2000
rect 28940 1975 28947 1995
rect 28947 1975 28965 1995
rect 28965 1975 28970 1995
rect 28940 1970 28970 1975
rect 29050 1995 29080 2000
rect 29050 1975 29057 1995
rect 29057 1975 29075 1995
rect 29075 1975 29080 1995
rect 29050 1970 29080 1975
rect 28050 1900 28080 1905
rect 28050 1880 28055 1900
rect 28055 1880 28075 1900
rect 28075 1880 28080 1900
rect 28050 1875 28080 1880
rect 28160 1900 28190 1905
rect 28160 1880 28165 1900
rect 28165 1880 28185 1900
rect 28185 1880 28190 1900
rect 28160 1875 28190 1880
rect 28270 1900 28300 1905
rect 28270 1880 28275 1900
rect 28275 1880 28295 1900
rect 28295 1880 28300 1900
rect 28270 1875 28300 1880
rect 28070 1675 28096 1680
rect 28070 1655 28071 1675
rect 28071 1655 28091 1675
rect 28091 1655 28096 1675
rect 28070 1650 28096 1655
rect 28015 1625 28045 1630
rect 28015 1605 28020 1625
rect 28020 1605 28040 1625
rect 28040 1605 28045 1625
rect 28015 1600 28045 1605
rect 28121 1600 28151 1630
rect 28215 1600 28245 1630
rect 28305 1625 28335 1630
rect 28305 1605 28310 1625
rect 28310 1605 28330 1625
rect 28330 1605 28335 1625
rect 28305 1600 28335 1605
rect 27820 1540 27850 1570
rect 27975 1565 28001 1570
rect 27975 1545 27976 1565
rect 27976 1545 27996 1565
rect 27996 1545 28001 1565
rect 27975 1540 28001 1545
rect 28349 1565 28375 1570
rect 28349 1545 28354 1565
rect 28354 1545 28374 1565
rect 28374 1545 28375 1565
rect 28349 1540 28375 1545
rect 26109 1490 26135 1495
rect 26109 1470 26112 1490
rect 26112 1470 26129 1490
rect 26129 1470 26135 1490
rect 26109 1465 26135 1470
rect 26310 1490 26340 1495
rect 26310 1470 26315 1490
rect 26315 1470 26335 1490
rect 26335 1470 26340 1490
rect 26310 1465 26340 1470
rect 26530 1490 26560 1495
rect 26530 1470 26535 1490
rect 26535 1470 26555 1490
rect 26555 1470 26560 1490
rect 26530 1465 26560 1470
rect 26925 1490 26951 1495
rect 26925 1470 26928 1490
rect 26928 1470 26945 1490
rect 26945 1470 26951 1490
rect 26925 1465 26951 1470
rect 27149 1490 27175 1495
rect 27149 1470 27152 1490
rect 27152 1470 27169 1490
rect 27169 1470 27175 1490
rect 27149 1465 27175 1470
rect 27350 1490 27380 1495
rect 27350 1470 27355 1490
rect 27355 1470 27375 1490
rect 27375 1470 27380 1490
rect 27350 1465 27380 1470
rect 27570 1490 27600 1495
rect 27570 1470 27575 1490
rect 27575 1470 27595 1490
rect 27595 1470 27600 1490
rect 27570 1465 27600 1470
rect 26150 1430 26180 1435
rect 26150 1410 26155 1430
rect 26155 1410 26175 1430
rect 26175 1410 26180 1430
rect 26150 1405 26180 1410
rect 26255 1430 26285 1435
rect 26255 1410 26260 1430
rect 26260 1410 26280 1430
rect 26280 1410 26285 1430
rect 26255 1405 26285 1410
rect 26365 1430 26395 1435
rect 26365 1410 26370 1430
rect 26370 1410 26390 1430
rect 26390 1410 26395 1430
rect 26365 1405 26395 1410
rect 26475 1430 26505 1435
rect 26475 1410 26480 1430
rect 26480 1410 26500 1430
rect 26500 1410 26505 1430
rect 26475 1405 26505 1410
rect 26585 1430 26615 1435
rect 26585 1410 26590 1430
rect 26590 1410 26610 1430
rect 26610 1410 26615 1430
rect 26585 1405 26615 1410
rect 12930 1360 12960 1390
rect 26815 1355 26845 1385
rect 26320 1305 26350 1335
rect 27190 1430 27220 1435
rect 27190 1410 27195 1430
rect 27195 1410 27215 1430
rect 27215 1410 27220 1430
rect 27190 1405 27220 1410
rect 27295 1430 27325 1435
rect 27295 1410 27300 1430
rect 27300 1410 27320 1430
rect 27320 1410 27325 1430
rect 27295 1405 27325 1410
rect 27405 1430 27435 1435
rect 27405 1410 27410 1430
rect 27410 1410 27430 1430
rect 27430 1410 27435 1430
rect 27405 1405 27435 1410
rect 27515 1430 27545 1435
rect 27515 1410 27520 1430
rect 27520 1410 27540 1430
rect 27540 1410 27545 1430
rect 27515 1405 27545 1410
rect 27625 1430 27655 1435
rect 27625 1410 27630 1430
rect 27630 1410 27650 1430
rect 27650 1410 27655 1430
rect 27625 1405 27655 1410
rect 26885 1305 26915 1335
rect 28028 1345 28054 1350
rect 28028 1325 28033 1345
rect 28033 1325 28053 1345
rect 28053 1325 28054 1345
rect 28028 1320 28054 1325
rect 28296 1345 28322 1350
rect 28296 1325 28297 1345
rect 28297 1325 28317 1345
rect 28317 1325 28322 1345
rect 28296 1320 28322 1325
rect 26430 1270 26460 1275
rect 26430 1250 26435 1270
rect 26435 1250 26455 1270
rect 26455 1250 26460 1270
rect 26430 1245 26460 1250
rect 26540 1270 26570 1275
rect 26540 1250 26545 1270
rect 26545 1250 26565 1270
rect 26565 1250 26570 1270
rect 26540 1245 26570 1250
rect 26650 1270 26680 1275
rect 26650 1250 26655 1270
rect 26655 1250 26675 1270
rect 26675 1250 26680 1270
rect 26650 1245 26680 1250
rect 26760 1270 26790 1275
rect 26760 1250 26765 1270
rect 26765 1250 26785 1270
rect 26785 1250 26790 1270
rect 26760 1245 26790 1250
rect 26870 1270 26900 1275
rect 26870 1250 26875 1270
rect 26875 1250 26895 1270
rect 26895 1250 26900 1270
rect 26870 1245 26900 1250
rect 26980 1270 27010 1275
rect 26980 1250 26985 1270
rect 26985 1250 27005 1270
rect 27005 1250 27010 1270
rect 26980 1245 27010 1250
rect 27090 1270 27120 1275
rect 27090 1250 27095 1270
rect 27095 1250 27115 1270
rect 27115 1250 27120 1270
rect 27090 1245 27120 1250
rect 27200 1270 27230 1275
rect 27200 1250 27205 1270
rect 27205 1250 27225 1270
rect 27225 1250 27230 1270
rect 27200 1245 27230 1250
rect 27310 1270 27340 1275
rect 27310 1250 27315 1270
rect 27315 1250 27335 1270
rect 27335 1250 27340 1270
rect 27310 1245 27340 1250
rect 27420 1270 27450 1275
rect 27420 1250 27425 1270
rect 27425 1250 27445 1270
rect 27445 1250 27450 1270
rect 27420 1245 27450 1250
rect 27530 1270 27560 1275
rect 27530 1250 27535 1270
rect 27535 1250 27555 1270
rect 27555 1250 27560 1270
rect 27530 1245 27560 1250
rect 27600 1285 27630 1290
rect 27600 1265 27605 1285
rect 27605 1265 27625 1285
rect 27625 1265 27630 1285
rect 27600 1260 27630 1265
rect 27950 1285 27980 1290
rect 27950 1265 27955 1285
rect 27955 1265 27975 1285
rect 27975 1265 27980 1285
rect 27950 1260 27980 1265
rect 28065 1285 28095 1290
rect 28065 1265 28070 1285
rect 28070 1265 28090 1285
rect 28090 1265 28095 1285
rect 28065 1260 28095 1265
rect 28160 1260 28190 1290
rect 28255 1285 28285 1290
rect 28255 1265 28260 1285
rect 28260 1265 28280 1285
rect 28280 1265 28285 1285
rect 28255 1260 28285 1265
rect 28370 1285 28400 1290
rect 28370 1265 28375 1285
rect 28375 1265 28395 1285
rect 28395 1265 28400 1285
rect 28370 1260 28400 1265
rect 28105 1225 28135 1230
rect 28105 1205 28110 1225
rect 28110 1205 28130 1225
rect 28130 1205 28135 1225
rect 28105 1200 28135 1205
rect 28160 1225 28190 1230
rect 28160 1205 28165 1225
rect 28165 1205 28185 1225
rect 28185 1205 28190 1225
rect 28160 1200 28190 1205
rect 28215 1225 28245 1230
rect 28215 1205 28220 1225
rect 28220 1205 28240 1225
rect 28240 1205 28245 1225
rect 28215 1200 28245 1205
rect 28370 1200 28400 1230
rect 13210 930 13240 935
rect 13210 910 13215 930
rect 13215 910 13235 930
rect 13235 910 13240 930
rect 13210 905 13240 910
rect 13410 930 13440 935
rect 13410 910 13415 930
rect 13415 910 13435 930
rect 13435 910 13440 930
rect 13410 905 13440 910
rect 26170 950 26200 955
rect 26170 930 26175 950
rect 26175 930 26195 950
rect 26195 930 26200 950
rect 26170 925 26200 930
rect 26265 950 26295 955
rect 26265 930 26270 950
rect 26270 930 26290 950
rect 26290 930 26295 950
rect 26265 925 26295 930
rect 26375 950 26405 955
rect 26375 930 26380 950
rect 26380 930 26400 950
rect 26400 930 26405 950
rect 26375 925 26405 930
rect 26485 950 26515 955
rect 26485 930 26490 950
rect 26490 930 26510 950
rect 26510 930 26515 950
rect 26485 925 26515 930
rect 26595 950 26625 955
rect 26595 930 26600 950
rect 26600 930 26620 950
rect 26620 930 26625 950
rect 26595 925 26625 930
rect 26705 950 26735 955
rect 26705 930 26710 950
rect 26710 930 26730 950
rect 26730 930 26735 950
rect 26705 925 26735 930
rect 26815 950 26845 955
rect 26815 930 26820 950
rect 26820 930 26840 950
rect 26840 930 26845 950
rect 26815 925 26845 930
rect 26925 950 26955 955
rect 26925 930 26930 950
rect 26930 930 26950 950
rect 26950 930 26955 950
rect 26925 925 26955 930
rect 27035 950 27065 955
rect 27035 930 27040 950
rect 27040 930 27060 950
rect 27060 930 27065 950
rect 27035 925 27065 930
rect 27145 950 27175 955
rect 27145 930 27150 950
rect 27150 930 27170 950
rect 27170 930 27175 950
rect 27145 925 27175 930
rect 27255 950 27285 955
rect 27255 930 27260 950
rect 27260 930 27280 950
rect 27280 930 27285 950
rect 27255 925 27285 930
rect 27365 950 27395 955
rect 27365 930 27370 950
rect 27370 930 27390 950
rect 27390 930 27395 950
rect 27365 925 27395 930
rect 27475 950 27505 955
rect 27475 930 27480 950
rect 27480 930 27500 950
rect 27500 930 27505 950
rect 27475 925 27505 930
rect 27625 950 27655 955
rect 27625 930 27630 950
rect 27630 930 27650 950
rect 27650 930 27655 950
rect 27625 925 27655 930
rect 12865 830 12895 860
rect 10955 765 10985 795
rect 2525 730 2555 760
rect 3135 755 3165 760
rect 3135 735 3140 755
rect 3140 735 3160 755
rect 3160 735 3165 755
rect 3135 730 3165 735
rect 3630 755 3660 760
rect 3630 735 3635 755
rect 3635 735 3655 755
rect 3655 735 3660 755
rect 3630 730 3660 735
rect 3990 755 4020 760
rect 3990 735 3995 755
rect 3995 735 4015 755
rect 4015 735 4020 755
rect 3990 730 4020 735
rect 4350 755 4380 760
rect 4350 735 4355 755
rect 4355 735 4375 755
rect 4375 735 4380 755
rect 4350 730 4380 735
rect 4530 755 4560 760
rect 4530 735 4535 755
rect 4535 735 4555 755
rect 4555 735 4560 755
rect 4530 730 4560 735
rect 4710 755 4740 760
rect 4710 735 4715 755
rect 4715 735 4735 755
rect 4735 735 4740 755
rect 4710 730 4740 735
rect 11310 790 11340 795
rect 11310 770 11315 790
rect 11315 770 11335 790
rect 11335 770 11340 790
rect 11310 765 11340 770
rect 11380 790 11410 795
rect 11380 770 11385 790
rect 11385 770 11405 790
rect 11405 770 11410 790
rect 11380 765 11410 770
rect 11450 790 11480 795
rect 11450 770 11455 790
rect 11455 770 11475 790
rect 11475 770 11480 790
rect 11450 765 11480 770
rect 12050 795 12080 800
rect 12050 775 12055 795
rect 12055 775 12075 795
rect 12075 775 12080 795
rect 12050 770 12080 775
rect 12270 795 12300 800
rect 12270 775 12275 795
rect 12275 775 12295 795
rect 12295 775 12300 795
rect 12270 770 12300 775
rect 12490 795 12520 800
rect 12490 775 12495 795
rect 12495 775 12515 795
rect 12515 775 12520 795
rect 12490 770 12520 775
rect 12810 770 12840 800
rect 4890 755 4920 760
rect 4890 735 4895 755
rect 4895 735 4915 755
rect 4915 735 4920 755
rect 4890 730 4920 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 11995 675 12025 680
rect 11995 655 12000 675
rect 12000 655 12020 675
rect 12020 655 12025 675
rect 11995 650 12025 655
rect 12105 675 12135 680
rect 12105 655 12110 675
rect 12110 655 12130 675
rect 12130 655 12135 675
rect 12105 650 12135 655
rect 12215 675 12245 680
rect 12215 655 12220 675
rect 12220 655 12240 675
rect 12240 655 12245 675
rect 12215 650 12245 655
rect 12325 675 12355 680
rect 12325 655 12330 675
rect 12330 655 12350 675
rect 12350 655 12355 675
rect 12325 650 12355 655
rect 12435 675 12465 680
rect 12435 655 12440 675
rect 12440 655 12460 675
rect 12460 655 12465 675
rect 12435 650 12465 655
rect 11345 -1380 11375 -1375
rect 11345 -1400 11350 -1380
rect 11350 -1400 11370 -1380
rect 11370 -1400 11375 -1380
rect 11345 -1405 11375 -1400
rect 11465 -1380 11495 -1375
rect 11465 -1400 11470 -1380
rect 11470 -1400 11490 -1380
rect 11490 -1400 11495 -1380
rect 11465 -1405 11495 -1400
rect 11585 -1380 11615 -1375
rect 11585 -1400 11590 -1380
rect 11590 -1400 11610 -1380
rect 11610 -1400 11615 -1380
rect 11585 -1405 11615 -1400
rect 11705 -1380 11735 -1375
rect 11705 -1400 11710 -1380
rect 11710 -1400 11730 -1380
rect 11730 -1400 11735 -1380
rect 11705 -1405 11735 -1400
rect 11825 -1380 11855 -1375
rect 11825 -1400 11830 -1380
rect 11830 -1400 11850 -1380
rect 11850 -1400 11855 -1380
rect 11825 -1405 11855 -1400
rect 11945 -1380 11975 -1375
rect 11945 -1400 11950 -1380
rect 11950 -1400 11970 -1380
rect 11970 -1400 11975 -1380
rect 11945 -1405 11975 -1400
rect 12065 -1380 12095 -1375
rect 12065 -1400 12070 -1380
rect 12070 -1400 12090 -1380
rect 12090 -1400 12095 -1380
rect 12065 -1405 12095 -1400
rect 12185 -1380 12215 -1375
rect 12185 -1400 12190 -1380
rect 12190 -1400 12210 -1380
rect 12210 -1400 12215 -1380
rect 12185 -1405 12215 -1400
rect 12305 -1380 12335 -1375
rect 12305 -1400 12310 -1380
rect 12310 -1400 12330 -1380
rect 12330 -1400 12335 -1380
rect 12305 -1405 12335 -1400
rect 12425 -1380 12455 -1375
rect 12425 -1400 12430 -1380
rect 12430 -1400 12450 -1380
rect 12450 -1400 12455 -1380
rect 12425 -1405 12455 -1400
rect 10585 -1795 10615 -1790
rect 10585 -1815 10590 -1795
rect 10590 -1815 10610 -1795
rect 10610 -1815 10615 -1795
rect 10585 -1820 10615 -1815
rect 10985 -1795 11015 -1790
rect 10985 -1815 10990 -1795
rect 10990 -1815 11010 -1795
rect 11010 -1815 11015 -1795
rect 10985 -1820 11015 -1815
rect 10905 -1875 10935 -1845
rect 11826 -1850 11854 -1845
rect 11826 -1870 11831 -1850
rect 11831 -1870 11849 -1850
rect 11849 -1870 11854 -1850
rect 11826 -1875 11854 -1870
rect 11285 -1930 11315 -1900
rect 11525 -1930 11555 -1900
rect 11765 -1930 11795 -1900
rect 12005 -1930 12035 -1900
rect 12245 -1930 12275 -1900
rect 12485 -1930 12515 -1900
rect 11405 -1975 11435 -1945
rect 11645 -1975 11675 -1945
rect 11885 -1975 11915 -1945
rect 12125 -1975 12155 -1945
rect 12365 -1975 12395 -1945
rect 11345 -2030 11375 -2000
rect 11405 -2030 11435 -2000
rect 11585 -2030 11615 -2000
rect 11825 -2030 11855 -2000
rect 12065 -2030 12095 -2000
rect 12305 -2030 12335 -2000
rect 12955 -1970 12985 -1965
rect 12955 -1990 12960 -1970
rect 12960 -1990 12980 -1970
rect 12980 -1990 12985 -1970
rect 12955 -1995 12985 -1990
rect 13065 -1970 13095 -1965
rect 13065 -1990 13070 -1970
rect 13070 -1990 13090 -1970
rect 13090 -1990 13095 -1970
rect 13065 -1995 13095 -1990
rect 13175 -1970 13205 -1965
rect 13175 -1990 13180 -1970
rect 13180 -1990 13200 -1970
rect 13200 -1990 13205 -1970
rect 13175 -1995 13205 -1990
rect 13285 -1970 13315 -1965
rect 13285 -1990 13290 -1970
rect 13290 -1990 13310 -1970
rect 13310 -1990 13315 -1970
rect 13285 -1995 13315 -1990
rect 13395 -1970 13425 -1965
rect 13395 -1990 13400 -1970
rect 13400 -1990 13420 -1970
rect 13420 -1990 13425 -1970
rect 13395 -1995 13425 -1990
rect 13505 -1970 13535 -1965
rect 13505 -1990 13510 -1970
rect 13510 -1990 13530 -1970
rect 13530 -1990 13535 -1970
rect 13505 -1995 13535 -1990
rect 13615 -1970 13645 -1965
rect 13615 -1990 13620 -1970
rect 13620 -1990 13640 -1970
rect 13640 -1990 13645 -1970
rect 13615 -1995 13645 -1990
rect 13725 -1970 13755 -1965
rect 13725 -1990 13730 -1970
rect 13730 -1990 13750 -1970
rect 13750 -1990 13755 -1970
rect 13725 -1995 13755 -1990
rect 13835 -1970 13865 -1965
rect 13835 -1990 13840 -1970
rect 13840 -1990 13860 -1970
rect 13860 -1990 13865 -1970
rect 13835 -1995 13865 -1990
rect 13945 -1970 13975 -1965
rect 13945 -1990 13950 -1970
rect 13950 -1990 13970 -1970
rect 13970 -1990 13975 -1970
rect 13945 -1995 13975 -1990
rect 14055 -1970 14085 -1965
rect 14055 -1990 14060 -1970
rect 14060 -1990 14080 -1970
rect 14080 -1990 14085 -1970
rect 14055 -1995 14085 -1990
rect 11465 -2060 11495 -2055
rect 11465 -2080 11470 -2060
rect 11470 -2080 11490 -2060
rect 11490 -2080 11495 -2060
rect 11465 -2085 11495 -2080
rect 11705 -2060 11735 -2055
rect 11705 -2080 11710 -2060
rect 11710 -2080 11730 -2060
rect 11730 -2080 11735 -2060
rect 11705 -2085 11735 -2080
rect 11945 -2060 11975 -2055
rect 11945 -2080 11950 -2060
rect 11950 -2080 11970 -2060
rect 11970 -2080 11975 -2060
rect 11945 -2085 11975 -2080
rect 12185 -2060 12215 -2055
rect 12185 -2080 12190 -2060
rect 12190 -2080 12210 -2060
rect 12210 -2080 12215 -2060
rect 12185 -2085 12215 -2080
rect 12425 -2060 12455 -2055
rect 12425 -2080 12430 -2060
rect 12430 -2080 12450 -2060
rect 12450 -2080 12455 -2060
rect 12425 -2085 12455 -2080
rect 12485 -2085 12515 -2055
rect 12695 -2300 12725 -2270
rect 10985 -2555 11015 -2525
rect 11826 -2530 11854 -2525
rect 11826 -2550 11831 -2530
rect 11831 -2550 11849 -2530
rect 11849 -2550 11854 -2530
rect 11826 -2555 11854 -2550
rect 11285 -2610 11315 -2580
rect 11525 -2610 11555 -2580
rect 11765 -2610 11795 -2580
rect 11405 -2655 11435 -2625
rect 11645 -2655 11675 -2625
rect 11445 -2750 11475 -2720
rect 11665 -2750 11695 -2720
rect 11335 -2795 11365 -2765
rect 11555 -2795 11585 -2765
rect 12005 -2610 12035 -2580
rect 12245 -2610 12275 -2580
rect 12485 -2610 12515 -2580
rect 13010 -2340 13040 -2335
rect 13010 -2360 13015 -2340
rect 13015 -2360 13035 -2340
rect 13035 -2360 13040 -2340
rect 13010 -2365 13040 -2360
rect 13120 -2340 13150 -2335
rect 13120 -2360 13125 -2340
rect 13125 -2360 13145 -2340
rect 13145 -2360 13150 -2340
rect 13120 -2365 13150 -2360
rect 13230 -2340 13260 -2335
rect 13230 -2360 13235 -2340
rect 13235 -2360 13255 -2340
rect 13255 -2360 13260 -2340
rect 13230 -2365 13260 -2360
rect 13340 -2340 13370 -2335
rect 13340 -2360 13345 -2340
rect 13345 -2360 13365 -2340
rect 13365 -2360 13370 -2340
rect 13340 -2365 13370 -2360
rect 13450 -2340 13480 -2335
rect 13450 -2360 13455 -2340
rect 13455 -2360 13475 -2340
rect 13475 -2360 13480 -2340
rect 13450 -2365 13480 -2360
rect 13560 -2340 13590 -2335
rect 13560 -2360 13565 -2340
rect 13565 -2360 13585 -2340
rect 13585 -2360 13590 -2340
rect 13560 -2365 13590 -2360
rect 13670 -2340 13700 -2335
rect 13670 -2360 13675 -2340
rect 13675 -2360 13695 -2340
rect 13695 -2360 13700 -2340
rect 13670 -2365 13700 -2360
rect 13780 -2340 13810 -2335
rect 13780 -2360 13785 -2340
rect 13785 -2360 13805 -2340
rect 13805 -2360 13810 -2340
rect 13780 -2365 13810 -2360
rect 13890 -2340 13920 -2335
rect 13890 -2360 13895 -2340
rect 13895 -2360 13915 -2340
rect 13915 -2360 13920 -2340
rect 13890 -2365 13920 -2360
rect 14000 -2340 14030 -2335
rect 14000 -2360 14005 -2340
rect 14005 -2360 14025 -2340
rect 14025 -2360 14030 -2340
rect 14000 -2365 14030 -2360
rect 12955 -2400 12985 -2395
rect 12955 -2420 12960 -2400
rect 12960 -2420 12980 -2400
rect 12980 -2420 12985 -2400
rect 12955 -2425 12985 -2420
rect 13065 -2400 13095 -2395
rect 13065 -2420 13070 -2400
rect 13070 -2420 13090 -2400
rect 13090 -2420 13095 -2400
rect 13065 -2425 13095 -2420
rect 13175 -2400 13205 -2395
rect 13175 -2420 13180 -2400
rect 13180 -2420 13200 -2400
rect 13200 -2420 13205 -2400
rect 13175 -2425 13205 -2420
rect 13285 -2400 13315 -2395
rect 13285 -2420 13290 -2400
rect 13290 -2420 13310 -2400
rect 13310 -2420 13315 -2400
rect 13285 -2425 13315 -2420
rect 13395 -2400 13425 -2395
rect 13395 -2420 13400 -2400
rect 13400 -2420 13420 -2400
rect 13420 -2420 13425 -2400
rect 13395 -2425 13425 -2420
rect 13505 -2400 13535 -2395
rect 13505 -2420 13510 -2400
rect 13510 -2420 13530 -2400
rect 13530 -2420 13535 -2400
rect 13505 -2425 13535 -2420
rect 13615 -2400 13645 -2395
rect 13615 -2420 13620 -2400
rect 13620 -2420 13640 -2400
rect 13640 -2420 13645 -2400
rect 13615 -2425 13645 -2420
rect 13725 -2400 13755 -2395
rect 13725 -2420 13730 -2400
rect 13730 -2420 13750 -2400
rect 13750 -2420 13755 -2400
rect 13725 -2425 13755 -2420
rect 13835 -2400 13865 -2395
rect 13835 -2420 13840 -2400
rect 13840 -2420 13860 -2400
rect 13860 -2420 13865 -2400
rect 13835 -2425 13865 -2420
rect 13945 -2400 13975 -2395
rect 13945 -2420 13950 -2400
rect 13950 -2420 13970 -2400
rect 13970 -2420 13975 -2400
rect 13945 -2425 13975 -2420
rect 14055 -2400 14085 -2395
rect 14055 -2420 14060 -2400
rect 14060 -2420 14080 -2400
rect 14080 -2420 14085 -2400
rect 14055 -2425 14085 -2420
rect 13010 -2570 13040 -2565
rect 13010 -2590 13015 -2570
rect 13015 -2590 13035 -2570
rect 13035 -2590 13040 -2570
rect 13010 -2595 13040 -2590
rect 13120 -2570 13150 -2565
rect 13120 -2590 13125 -2570
rect 13125 -2590 13145 -2570
rect 13145 -2590 13150 -2570
rect 13120 -2595 13150 -2590
rect 13230 -2570 13260 -2565
rect 13230 -2590 13235 -2570
rect 13235 -2590 13255 -2570
rect 13255 -2590 13260 -2570
rect 13230 -2595 13260 -2590
rect 13340 -2570 13370 -2565
rect 13340 -2590 13345 -2570
rect 13345 -2590 13365 -2570
rect 13365 -2590 13370 -2570
rect 13340 -2595 13370 -2590
rect 13450 -2570 13480 -2565
rect 13450 -2590 13455 -2570
rect 13455 -2590 13475 -2570
rect 13475 -2590 13480 -2570
rect 13450 -2595 13480 -2590
rect 13560 -2570 13590 -2565
rect 13560 -2590 13565 -2570
rect 13565 -2590 13585 -2570
rect 13585 -2590 13590 -2570
rect 13560 -2595 13590 -2590
rect 13670 -2570 13700 -2565
rect 13670 -2590 13675 -2570
rect 13675 -2590 13695 -2570
rect 13695 -2590 13700 -2570
rect 13670 -2595 13700 -2590
rect 13780 -2570 13810 -2565
rect 13780 -2590 13785 -2570
rect 13785 -2590 13805 -2570
rect 13805 -2590 13810 -2570
rect 13780 -2595 13810 -2590
rect 13890 -2570 13920 -2565
rect 13890 -2590 13895 -2570
rect 13895 -2590 13915 -2570
rect 13915 -2590 13920 -2570
rect 13890 -2595 13920 -2590
rect 14000 -2570 14030 -2565
rect 14000 -2590 14005 -2570
rect 14005 -2590 14025 -2570
rect 14025 -2590 14030 -2570
rect 14000 -2595 14030 -2590
rect 11885 -2655 11915 -2625
rect 12125 -2655 12155 -2625
rect 12365 -2655 12395 -2625
rect 12695 -2655 12725 -2625
rect 12980 -2630 13010 -2625
rect 12980 -2650 12985 -2630
rect 12985 -2650 13005 -2630
rect 13005 -2650 13010 -2630
rect 12980 -2655 13010 -2650
rect 13010 -2690 13040 -2685
rect 13010 -2710 13015 -2690
rect 13015 -2710 13035 -2690
rect 13035 -2710 13040 -2690
rect 13010 -2715 13040 -2710
rect 11885 -2750 11915 -2720
rect 12105 -2750 12135 -2720
rect 13120 -2690 13150 -2685
rect 13120 -2710 13125 -2690
rect 13125 -2710 13145 -2690
rect 13145 -2710 13150 -2690
rect 13120 -2715 13150 -2710
rect 13230 -2690 13260 -2685
rect 13230 -2710 13235 -2690
rect 13235 -2710 13255 -2690
rect 13255 -2710 13260 -2690
rect 13230 -2715 13260 -2710
rect 13340 -2690 13370 -2685
rect 13340 -2710 13345 -2690
rect 13345 -2710 13365 -2690
rect 13365 -2710 13370 -2690
rect 13340 -2715 13370 -2710
rect 13450 -2690 13480 -2685
rect 13450 -2710 13455 -2690
rect 13455 -2710 13475 -2690
rect 13475 -2710 13480 -2690
rect 13450 -2715 13480 -2710
rect 13560 -2690 13590 -2685
rect 13560 -2710 13565 -2690
rect 13565 -2710 13585 -2690
rect 13585 -2710 13590 -2690
rect 13560 -2715 13590 -2710
rect 13670 -2690 13700 -2685
rect 13670 -2710 13675 -2690
rect 13675 -2710 13695 -2690
rect 13695 -2710 13700 -2690
rect 13670 -2715 13700 -2710
rect 13780 -2690 13810 -2685
rect 13780 -2710 13785 -2690
rect 13785 -2710 13805 -2690
rect 13805 -2710 13810 -2690
rect 13780 -2715 13810 -2710
rect 13890 -2690 13920 -2685
rect 13890 -2710 13895 -2690
rect 13895 -2710 13915 -2690
rect 13915 -2710 13920 -2690
rect 13890 -2715 13920 -2710
rect 14000 -2690 14030 -2685
rect 14000 -2710 14005 -2690
rect 14005 -2710 14025 -2690
rect 14025 -2710 14030 -2690
rect 14000 -2715 14030 -2710
rect 12325 -2750 12355 -2720
rect 11775 -2795 11805 -2765
rect 11995 -2795 12025 -2765
rect 12215 -2795 12245 -2765
rect 12435 -2795 12465 -2765
rect 12955 -2910 12985 -2905
rect 12955 -2930 12962 -2910
rect 12962 -2930 12980 -2910
rect 12980 -2930 12985 -2910
rect 12955 -2935 12985 -2930
rect 13065 -2910 13095 -2905
rect 13065 -2930 13072 -2910
rect 13072 -2930 13090 -2910
rect 13090 -2930 13095 -2910
rect 13065 -2935 13095 -2930
rect 13175 -2910 13205 -2905
rect 13175 -2930 13182 -2910
rect 13182 -2930 13200 -2910
rect 13200 -2930 13205 -2910
rect 13175 -2935 13205 -2930
rect 13285 -2910 13315 -2905
rect 13285 -2930 13292 -2910
rect 13292 -2930 13310 -2910
rect 13310 -2930 13315 -2910
rect 13285 -2935 13315 -2930
rect 13395 -2910 13425 -2905
rect 13395 -2930 13402 -2910
rect 13402 -2930 13420 -2910
rect 13420 -2930 13425 -2910
rect 13395 -2935 13425 -2930
rect 13505 -2910 13535 -2905
rect 13505 -2930 13512 -2910
rect 13512 -2930 13530 -2910
rect 13530 -2930 13535 -2910
rect 13505 -2935 13535 -2930
rect 13615 -2910 13645 -2905
rect 13615 -2930 13622 -2910
rect 13622 -2930 13640 -2910
rect 13640 -2930 13645 -2910
rect 13615 -2935 13645 -2930
rect 13725 -2910 13755 -2905
rect 13725 -2930 13732 -2910
rect 13732 -2930 13750 -2910
rect 13750 -2930 13755 -2910
rect 13725 -2935 13755 -2930
rect 13835 -2910 13865 -2905
rect 13835 -2930 13842 -2910
rect 13842 -2930 13860 -2910
rect 13860 -2930 13865 -2910
rect 13835 -2935 13865 -2930
rect 13945 -2910 13975 -2905
rect 13945 -2930 13952 -2910
rect 13952 -2930 13970 -2910
rect 13970 -2930 13975 -2910
rect 13945 -2935 13975 -2930
rect 14055 -2910 14085 -2905
rect 14055 -2930 14062 -2910
rect 14062 -2930 14080 -2910
rect 14080 -2930 14085 -2910
rect 14055 -2935 14085 -2930
rect 13000 -2970 13030 -2965
rect 13000 -2990 13005 -2970
rect 13005 -2990 13025 -2970
rect 13025 -2990 13030 -2970
rect 13000 -2995 13030 -2990
rect 13200 -2970 13230 -2965
rect 13200 -2990 13205 -2970
rect 13205 -2990 13225 -2970
rect 13225 -2990 13230 -2970
rect 13200 -2995 13230 -2990
rect 13400 -2970 13430 -2965
rect 13400 -2990 13405 -2970
rect 13405 -2990 13425 -2970
rect 13425 -2990 13430 -2970
rect 13400 -2995 13430 -2990
rect 13600 -2970 13630 -2965
rect 13600 -2990 13605 -2970
rect 13605 -2990 13625 -2970
rect 13625 -2990 13630 -2970
rect 13600 -2995 13630 -2990
rect 13800 -2970 13830 -2965
rect 13800 -2990 13805 -2970
rect 13805 -2990 13825 -2970
rect 13825 -2990 13830 -2970
rect 13800 -2995 13830 -2990
rect 14000 -2970 14030 -2965
rect 14000 -2990 14005 -2970
rect 14005 -2990 14025 -2970
rect 14025 -2990 14030 -2970
rect 14000 -2995 14030 -2990
rect 11390 -3045 11420 -3040
rect 11390 -3065 11395 -3045
rect 11395 -3065 11415 -3045
rect 11415 -3065 11420 -3045
rect 11390 -3070 11420 -3065
rect 11610 -3045 11640 -3040
rect 11610 -3065 11615 -3045
rect 11615 -3065 11635 -3045
rect 11635 -3065 11640 -3045
rect 11610 -3070 11640 -3065
rect 11830 -3045 11860 -3040
rect 11830 -3065 11835 -3045
rect 11835 -3065 11855 -3045
rect 11855 -3065 11860 -3045
rect 11830 -3070 11860 -3065
rect 12050 -3045 12080 -3040
rect 12050 -3065 12055 -3045
rect 12055 -3065 12075 -3045
rect 12075 -3065 12080 -3045
rect 12050 -3070 12080 -3065
rect 12270 -3045 12300 -3040
rect 12270 -3065 12275 -3045
rect 12275 -3065 12295 -3045
rect 12295 -3065 12300 -3045
rect 12270 -3070 12300 -3065
rect 11500 -3125 11530 -3095
rect 11720 -3125 11750 -3095
rect 11940 -3125 11970 -3095
rect 12160 -3125 12190 -3095
rect 11195 -3180 11225 -3150
rect 11415 -3180 11445 -3150
rect 11090 -3245 11120 -3240
rect 11090 -3265 11095 -3245
rect 11095 -3265 11115 -3245
rect 11115 -3265 11120 -3245
rect 11090 -3270 11120 -3265
rect 11310 -3245 11340 -3240
rect 11310 -3265 11315 -3245
rect 11315 -3265 11335 -3245
rect 11335 -3265 11340 -3245
rect 11310 -3270 11340 -3265
rect 12380 -3125 12410 -3095
rect 11645 -3180 11675 -3150
rect 12235 -3180 12265 -3150
rect 12455 -3180 12485 -3150
rect 12685 -3180 12715 -3150
rect 11825 -3225 11855 -3195
rect 11945 -3225 11975 -3195
rect 11530 -3245 11560 -3240
rect 11530 -3265 11535 -3245
rect 11535 -3265 11555 -3245
rect 11555 -3265 11560 -3245
rect 11530 -3270 11560 -3265
rect 12130 -3245 12160 -3240
rect 12130 -3265 12135 -3245
rect 12135 -3265 12155 -3245
rect 12155 -3265 12160 -3245
rect 12130 -3270 12160 -3265
rect 12350 -3245 12380 -3240
rect 12350 -3265 12355 -3245
rect 12355 -3265 12375 -3245
rect 12375 -3265 12380 -3245
rect 12350 -3270 12380 -3265
rect 12570 -3245 12600 -3240
rect 12570 -3265 12575 -3245
rect 12575 -3265 12595 -3245
rect 12595 -3265 12600 -3245
rect 12570 -3270 12600 -3265
rect 11240 -3290 11266 -3285
rect 11240 -3310 11243 -3290
rect 11243 -3310 11260 -3290
rect 11260 -3310 11266 -3290
rect 11240 -3315 11266 -3310
rect 11460 -3290 11486 -3285
rect 11460 -3310 11463 -3290
rect 11463 -3310 11480 -3290
rect 11480 -3310 11486 -3290
rect 11460 -3315 11486 -3310
rect 11604 -3290 11630 -3285
rect 11604 -3310 11610 -3290
rect 11610 -3310 11627 -3290
rect 11627 -3310 11630 -3290
rect 11604 -3315 11630 -3310
rect 11870 -3290 11896 -3285
rect 11870 -3310 11876 -3290
rect 11876 -3310 11893 -3290
rect 11893 -3310 11896 -3290
rect 11870 -3315 11896 -3310
rect 12280 -3290 12306 -3285
rect 12280 -3310 12283 -3290
rect 12283 -3310 12300 -3290
rect 12300 -3310 12306 -3290
rect 12280 -3315 12306 -3310
rect 12500 -3290 12526 -3285
rect 12500 -3310 12503 -3290
rect 12503 -3310 12520 -3290
rect 12520 -3310 12526 -3290
rect 12500 -3315 12526 -3310
rect 12644 -3290 12670 -3285
rect 12644 -3310 12650 -3290
rect 12650 -3310 12667 -3290
rect 12667 -3310 12670 -3290
rect 12644 -3315 12670 -3310
rect 13100 -3320 13130 -3315
rect 13100 -3340 13105 -3320
rect 13105 -3340 13125 -3320
rect 13125 -3340 13130 -3320
rect 13100 -3345 13130 -3340
rect 13300 -3320 13330 -3315
rect 13300 -3340 13305 -3320
rect 13305 -3340 13325 -3320
rect 13325 -3340 13330 -3320
rect 13300 -3345 13330 -3340
rect 13500 -3320 13530 -3315
rect 13500 -3340 13505 -3320
rect 13505 -3340 13525 -3320
rect 13525 -3340 13530 -3320
rect 13500 -3345 13530 -3340
rect 13700 -3320 13730 -3315
rect 13700 -3340 13705 -3320
rect 13705 -3340 13725 -3320
rect 13725 -3340 13730 -3320
rect 13700 -3345 13730 -3340
rect 13900 -3320 13930 -3315
rect 13900 -3340 13905 -3320
rect 13905 -3340 13925 -3320
rect 13925 -3340 13930 -3320
rect 13900 -3345 13930 -3340
rect 11109 -3510 11135 -3505
rect 11109 -3530 11112 -3510
rect 11112 -3530 11129 -3510
rect 11129 -3530 11135 -3510
rect 11109 -3535 11135 -3530
rect 11310 -3510 11340 -3505
rect 11310 -3530 11315 -3510
rect 11315 -3530 11335 -3510
rect 11335 -3530 11340 -3510
rect 11310 -3535 11340 -3530
rect 11530 -3510 11560 -3505
rect 11530 -3530 11535 -3510
rect 11535 -3530 11555 -3510
rect 11555 -3530 11560 -3510
rect 11530 -3535 11560 -3530
rect 11925 -3510 11951 -3505
rect 11925 -3530 11928 -3510
rect 11928 -3530 11945 -3510
rect 11945 -3530 11951 -3510
rect 11925 -3535 11951 -3530
rect 12149 -3510 12175 -3505
rect 12149 -3530 12152 -3510
rect 12152 -3530 12169 -3510
rect 12169 -3530 12175 -3510
rect 12149 -3535 12175 -3530
rect 12350 -3510 12380 -3505
rect 12350 -3530 12355 -3510
rect 12355 -3530 12375 -3510
rect 12375 -3530 12380 -3510
rect 12350 -3535 12380 -3530
rect 12570 -3510 12600 -3505
rect 12570 -3530 12575 -3510
rect 12575 -3530 12595 -3510
rect 12595 -3530 12600 -3510
rect 12570 -3535 12600 -3530
rect 11150 -3570 11180 -3565
rect 11150 -3590 11155 -3570
rect 11155 -3590 11175 -3570
rect 11175 -3590 11180 -3570
rect 11150 -3595 11180 -3590
rect 11255 -3570 11285 -3565
rect 11255 -3590 11260 -3570
rect 11260 -3590 11280 -3570
rect 11280 -3590 11285 -3570
rect 11255 -3595 11285 -3590
rect 11365 -3570 11395 -3565
rect 11365 -3590 11370 -3570
rect 11370 -3590 11390 -3570
rect 11390 -3590 11395 -3570
rect 11365 -3595 11395 -3590
rect 11475 -3570 11505 -3565
rect 11475 -3590 11480 -3570
rect 11480 -3590 11500 -3570
rect 11500 -3590 11505 -3570
rect 11475 -3595 11505 -3590
rect 11585 -3570 11615 -3565
rect 11585 -3590 11590 -3570
rect 11590 -3590 11610 -3570
rect 11610 -3590 11615 -3570
rect 11585 -3595 11615 -3590
rect 11815 -3685 11845 -3655
rect 11320 -3735 11350 -3705
rect 12190 -3570 12220 -3565
rect 12190 -3590 12195 -3570
rect 12195 -3590 12215 -3570
rect 12215 -3590 12220 -3570
rect 12190 -3595 12220 -3590
rect 12295 -3570 12325 -3565
rect 12295 -3590 12300 -3570
rect 12300 -3590 12320 -3570
rect 12320 -3590 12325 -3570
rect 12295 -3595 12325 -3590
rect 12405 -3570 12435 -3565
rect 12405 -3590 12410 -3570
rect 12410 -3590 12430 -3570
rect 12430 -3590 12435 -3570
rect 12405 -3595 12435 -3590
rect 12515 -3570 12545 -3565
rect 12515 -3590 12520 -3570
rect 12520 -3590 12540 -3570
rect 12540 -3590 12545 -3570
rect 12515 -3595 12545 -3590
rect 12625 -3570 12655 -3565
rect 12625 -3590 12630 -3570
rect 12630 -3590 12650 -3570
rect 12650 -3590 12655 -3570
rect 12625 -3595 12655 -3590
rect 11885 -3735 11915 -3705
rect 11430 -3770 11460 -3765
rect 11430 -3790 11435 -3770
rect 11435 -3790 11455 -3770
rect 11455 -3790 11460 -3770
rect 11430 -3795 11460 -3790
rect 11540 -3770 11570 -3765
rect 11540 -3790 11545 -3770
rect 11545 -3790 11565 -3770
rect 11565 -3790 11570 -3770
rect 11540 -3795 11570 -3790
rect 11650 -3770 11680 -3765
rect 11650 -3790 11655 -3770
rect 11655 -3790 11675 -3770
rect 11675 -3790 11680 -3770
rect 11650 -3795 11680 -3790
rect 11760 -3770 11790 -3765
rect 11760 -3790 11765 -3770
rect 11765 -3790 11785 -3770
rect 11785 -3790 11790 -3770
rect 11760 -3795 11790 -3790
rect 11870 -3770 11900 -3765
rect 11870 -3790 11875 -3770
rect 11875 -3790 11895 -3770
rect 11895 -3790 11900 -3770
rect 11870 -3795 11900 -3790
rect 11980 -3770 12010 -3765
rect 11980 -3790 11985 -3770
rect 11985 -3790 12005 -3770
rect 12005 -3790 12010 -3770
rect 11980 -3795 12010 -3790
rect 12090 -3770 12120 -3765
rect 12090 -3790 12095 -3770
rect 12095 -3790 12115 -3770
rect 12115 -3790 12120 -3770
rect 12090 -3795 12120 -3790
rect 12200 -3770 12230 -3765
rect 12200 -3790 12205 -3770
rect 12205 -3790 12225 -3770
rect 12225 -3790 12230 -3770
rect 12200 -3795 12230 -3790
rect 12310 -3770 12340 -3765
rect 12310 -3790 12315 -3770
rect 12315 -3790 12335 -3770
rect 12335 -3790 12340 -3770
rect 12310 -3795 12340 -3790
rect 12420 -3770 12450 -3765
rect 12420 -3790 12425 -3770
rect 12425 -3790 12445 -3770
rect 12445 -3790 12450 -3770
rect 12420 -3795 12450 -3790
rect 12530 -3770 12560 -3765
rect 12530 -3790 12535 -3770
rect 12535 -3790 12555 -3770
rect 12555 -3790 12560 -3770
rect 12530 -3795 12560 -3790
rect 12600 -3755 12630 -3750
rect 12600 -3775 12605 -3755
rect 12605 -3775 12625 -3755
rect 12625 -3775 12630 -3755
rect 12600 -3780 12630 -3775
rect 11170 -4090 11200 -4085
rect 11170 -4110 11175 -4090
rect 11175 -4110 11195 -4090
rect 11195 -4110 11200 -4090
rect 11170 -4115 11200 -4110
rect 11265 -4090 11295 -4085
rect 11265 -4110 11270 -4090
rect 11270 -4110 11290 -4090
rect 11290 -4110 11295 -4090
rect 11265 -4115 11295 -4110
rect 11375 -4090 11405 -4085
rect 11375 -4110 11380 -4090
rect 11380 -4110 11400 -4090
rect 11400 -4110 11405 -4090
rect 11375 -4115 11405 -4110
rect 11485 -4090 11515 -4085
rect 11485 -4110 11490 -4090
rect 11490 -4110 11510 -4090
rect 11510 -4110 11515 -4090
rect 11485 -4115 11515 -4110
rect 11595 -4090 11625 -4085
rect 11595 -4110 11600 -4090
rect 11600 -4110 11620 -4090
rect 11620 -4110 11625 -4090
rect 11595 -4115 11625 -4110
rect 11705 -4090 11735 -4085
rect 11705 -4110 11710 -4090
rect 11710 -4110 11730 -4090
rect 11730 -4110 11735 -4090
rect 11705 -4115 11735 -4110
rect 11815 -4090 11845 -4085
rect 11815 -4110 11820 -4090
rect 11820 -4110 11840 -4090
rect 11840 -4110 11845 -4090
rect 11815 -4115 11845 -4110
rect 11925 -4090 11955 -4085
rect 11925 -4110 11930 -4090
rect 11930 -4110 11950 -4090
rect 11950 -4110 11955 -4090
rect 11925 -4115 11955 -4110
rect 12035 -4090 12065 -4085
rect 12035 -4110 12040 -4090
rect 12040 -4110 12060 -4090
rect 12060 -4110 12065 -4090
rect 12035 -4115 12065 -4110
rect 12145 -4090 12175 -4085
rect 12145 -4110 12150 -4090
rect 12150 -4110 12170 -4090
rect 12170 -4110 12175 -4090
rect 12145 -4115 12175 -4110
rect 12255 -4090 12285 -4085
rect 12255 -4110 12260 -4090
rect 12260 -4110 12280 -4090
rect 12280 -4110 12285 -4090
rect 12255 -4115 12285 -4110
rect 12365 -4090 12395 -4085
rect 12365 -4110 12370 -4090
rect 12370 -4110 12390 -4090
rect 12390 -4110 12395 -4090
rect 12365 -4115 12395 -4110
rect 12475 -4090 12505 -4085
rect 12475 -4110 12480 -4090
rect 12480 -4110 12500 -4090
rect 12500 -4110 12505 -4090
rect 12475 -4115 12505 -4110
rect 12625 -4090 12655 -4085
rect 12625 -4110 12630 -4090
rect 12630 -4110 12650 -4090
rect 12650 -4110 12655 -4090
rect 12625 -4115 12655 -4110
<< metal2 >>
rect 11632 9055 11668 9060
rect 11632 9025 11635 9055
rect 11665 9050 11668 9055
rect 11752 9055 11788 9060
rect 11752 9050 11755 9055
rect 11665 9030 11755 9050
rect 11665 9025 11668 9030
rect 11632 9020 11668 9025
rect 11752 9025 11755 9030
rect 11785 9050 11788 9055
rect 11872 9055 11908 9060
rect 11872 9050 11875 9055
rect 11785 9030 11875 9050
rect 11785 9025 11788 9030
rect 11752 9020 11788 9025
rect 11872 9025 11875 9030
rect 11905 9050 11908 9055
rect 12080 9055 12120 9060
rect 12080 9050 12085 9055
rect 11905 9030 12085 9050
rect 11905 9025 11908 9030
rect 11872 9020 11908 9025
rect 12080 9025 12085 9030
rect 12115 9025 12120 9055
rect 12080 9020 12120 9025
rect 11570 9010 11610 9015
rect 11570 9000 11575 9010
rect 11200 8995 11240 9000
rect 11200 8965 11205 8995
rect 11235 8965 11240 8995
rect 11200 8960 11240 8965
rect 11460 8995 11575 9000
rect 11460 8965 11465 8995
rect 11495 8980 11575 8995
rect 11605 9005 11610 9010
rect 11690 9010 11730 9015
rect 11690 9005 11695 9010
rect 11605 8985 11695 9005
rect 11605 8980 11610 8985
rect 11495 8965 11500 8980
rect 11570 8975 11610 8980
rect 11690 8980 11695 8985
rect 11725 9005 11730 9010
rect 11810 9010 11850 9015
rect 11810 9005 11815 9010
rect 11725 8985 11815 9005
rect 11725 8980 11730 8985
rect 11690 8975 11730 8980
rect 11810 8980 11815 8985
rect 11845 9005 11850 9010
rect 11930 9010 11970 9015
rect 11930 9005 11935 9010
rect 11845 8985 11935 9005
rect 11845 8980 11850 8985
rect 11810 8975 11850 8980
rect 11930 8980 11935 8985
rect 11965 8980 11970 9010
rect 11930 8975 11970 8980
rect 12080 8985 12120 8990
rect 11460 8960 11500 8965
rect 12080 8955 12085 8985
rect 12115 8980 12120 8985
rect 12200 8985 12240 8990
rect 12200 8980 12205 8985
rect 12115 8960 12205 8980
rect 12115 8955 12120 8960
rect 12080 8950 12120 8955
rect 12200 8955 12205 8960
rect 12235 8980 12240 8985
rect 12320 8985 12360 8990
rect 12320 8980 12325 8985
rect 12235 8960 12325 8980
rect 12235 8955 12240 8960
rect 12200 8950 12240 8955
rect 12320 8955 12325 8960
rect 12355 8980 12360 8985
rect 12440 8985 12480 8990
rect 12440 8980 12445 8985
rect 12355 8960 12445 8980
rect 12355 8955 12360 8960
rect 12320 8950 12360 8955
rect 12440 8955 12445 8960
rect 12475 8980 12480 8985
rect 12560 8985 12600 8990
rect 12560 8980 12565 8985
rect 12475 8960 12565 8980
rect 12475 8955 12480 8960
rect 12440 8950 12480 8955
rect 12560 8955 12565 8960
rect 12595 8955 12600 8985
rect 12560 8950 12600 8955
rect 11330 8860 11370 8865
rect 11330 8830 11335 8860
rect 11365 8830 11370 8860
rect 11330 8825 11370 8830
rect 11750 8855 11790 8860
rect 11750 8825 11755 8855
rect 11785 8850 11790 8855
rect 12140 8855 12180 8860
rect 12140 8850 12145 8855
rect 11785 8830 12145 8850
rect 11785 8825 11790 8830
rect 11750 8820 11790 8825
rect 12140 8825 12145 8830
rect 12175 8850 12180 8855
rect 12260 8855 12300 8860
rect 12260 8850 12265 8855
rect 12175 8830 12265 8850
rect 12175 8825 12180 8830
rect 12140 8820 12180 8825
rect 12260 8825 12265 8830
rect 12295 8850 12300 8855
rect 12380 8855 12420 8860
rect 12380 8850 12385 8855
rect 12295 8830 12385 8850
rect 12295 8825 12300 8830
rect 12260 8820 12300 8825
rect 12380 8825 12385 8830
rect 12415 8850 12420 8855
rect 12500 8855 12540 8860
rect 12500 8850 12505 8855
rect 12415 8830 12505 8850
rect 12415 8825 12420 8830
rect 12380 8820 12420 8825
rect 12500 8825 12505 8830
rect 12535 8825 12540 8855
rect 12500 8820 12540 8825
rect 11330 8765 11370 8770
rect 11330 8735 11335 8765
rect 11365 8760 11370 8765
rect 12200 8765 12240 8770
rect 12200 8760 12205 8765
rect 11365 8740 12205 8760
rect 11365 8735 11370 8740
rect 11330 8730 11370 8735
rect 12200 8735 12205 8740
rect 12235 8735 12240 8765
rect 12200 8730 12240 8735
rect 11340 8625 11380 8630
rect 11340 8595 11345 8625
rect 11375 8620 11380 8625
rect 11460 8625 11500 8630
rect 11460 8620 11465 8625
rect 11375 8600 11465 8620
rect 11375 8595 11380 8600
rect 11340 8590 11380 8595
rect 11460 8595 11465 8600
rect 11495 8620 11500 8625
rect 11580 8625 11620 8630
rect 11580 8620 11585 8625
rect 11495 8600 11585 8620
rect 11495 8595 11500 8600
rect 11460 8590 11500 8595
rect 11580 8595 11585 8600
rect 11615 8620 11620 8625
rect 11700 8625 11740 8630
rect 11700 8620 11705 8625
rect 11615 8600 11705 8620
rect 11615 8595 11620 8600
rect 11580 8590 11620 8595
rect 11700 8595 11705 8600
rect 11735 8620 11740 8625
rect 11820 8625 11860 8630
rect 11820 8620 11825 8625
rect 11735 8600 11825 8620
rect 11735 8595 11740 8600
rect 11700 8590 11740 8595
rect 11820 8595 11825 8600
rect 11855 8620 11860 8625
rect 11940 8625 11980 8630
rect 11940 8620 11945 8625
rect 11855 8600 11945 8620
rect 11855 8595 11860 8600
rect 11820 8590 11860 8595
rect 11940 8595 11945 8600
rect 11975 8620 11980 8625
rect 12060 8625 12100 8630
rect 12060 8620 12065 8625
rect 11975 8600 12065 8620
rect 11975 8595 11980 8600
rect 11940 8590 11980 8595
rect 12060 8595 12065 8600
rect 12095 8620 12100 8625
rect 12180 8625 12220 8630
rect 12180 8620 12185 8625
rect 12095 8600 12185 8620
rect 12095 8595 12100 8600
rect 12060 8590 12100 8595
rect 12180 8595 12185 8600
rect 12215 8620 12220 8625
rect 12300 8625 12340 8630
rect 12300 8620 12305 8625
rect 12215 8600 12305 8620
rect 12215 8595 12220 8600
rect 12180 8590 12220 8595
rect 12300 8595 12305 8600
rect 12335 8620 12340 8625
rect 12420 8625 12460 8630
rect 12420 8620 12425 8625
rect 12335 8600 12425 8620
rect 12335 8595 12340 8600
rect 12300 8590 12340 8595
rect 12420 8595 12425 8600
rect 12455 8595 12460 8625
rect 12420 8590 12460 8595
rect 18840 8625 18880 8630
rect 18840 8595 18845 8625
rect 18875 8620 18880 8625
rect 18960 8625 19000 8630
rect 18960 8620 18965 8625
rect 18875 8600 18965 8620
rect 18875 8595 18880 8600
rect 18840 8590 18880 8595
rect 18960 8595 18965 8600
rect 18995 8620 19000 8625
rect 19080 8625 19120 8630
rect 19080 8620 19085 8625
rect 18995 8600 19085 8620
rect 18995 8595 19000 8600
rect 18960 8590 19000 8595
rect 19080 8595 19085 8600
rect 19115 8620 19120 8625
rect 19200 8625 19240 8630
rect 19200 8620 19205 8625
rect 19115 8600 19205 8620
rect 19115 8595 19120 8600
rect 19080 8590 19120 8595
rect 19200 8595 19205 8600
rect 19235 8620 19240 8625
rect 19320 8625 19360 8630
rect 19320 8620 19325 8625
rect 19235 8600 19325 8620
rect 19235 8595 19240 8600
rect 19200 8590 19240 8595
rect 19320 8595 19325 8600
rect 19355 8620 19360 8625
rect 19440 8625 19480 8630
rect 19440 8620 19445 8625
rect 19355 8600 19445 8620
rect 19355 8595 19360 8600
rect 19320 8590 19360 8595
rect 19440 8595 19445 8600
rect 19475 8620 19480 8625
rect 19560 8625 19600 8630
rect 19560 8620 19565 8625
rect 19475 8600 19565 8620
rect 19475 8595 19480 8600
rect 19440 8590 19480 8595
rect 19560 8595 19565 8600
rect 19595 8620 19600 8625
rect 19680 8625 19720 8630
rect 19680 8620 19685 8625
rect 19595 8600 19685 8620
rect 19595 8595 19600 8600
rect 19560 8590 19600 8595
rect 19680 8595 19685 8600
rect 19715 8620 19720 8625
rect 19800 8625 19840 8630
rect 19800 8620 19805 8625
rect 19715 8600 19805 8620
rect 19715 8595 19720 8600
rect 19680 8590 19720 8595
rect 19800 8595 19805 8600
rect 19835 8620 19840 8625
rect 19920 8625 19960 8630
rect 19920 8620 19925 8625
rect 19835 8600 19925 8620
rect 19835 8595 19840 8600
rect 19800 8590 19840 8595
rect 19920 8595 19925 8600
rect 19955 8595 19960 8625
rect 19920 8590 19960 8595
rect 12950 8290 12990 8295
rect 12950 8260 12955 8290
rect 12985 8285 12990 8290
rect 13060 8290 13100 8295
rect 13060 8285 13065 8290
rect 12985 8265 13065 8285
rect 12985 8260 12990 8265
rect 12950 8255 12990 8260
rect 13060 8260 13065 8265
rect 13095 8285 13100 8290
rect 13170 8290 13210 8295
rect 13170 8285 13175 8290
rect 13095 8265 13175 8285
rect 13095 8260 13100 8265
rect 13060 8255 13100 8260
rect 13170 8260 13175 8265
rect 13205 8285 13210 8290
rect 13280 8290 13320 8295
rect 13280 8285 13285 8290
rect 13205 8265 13285 8285
rect 13205 8260 13210 8265
rect 13170 8255 13210 8260
rect 13280 8260 13285 8265
rect 13315 8285 13320 8290
rect 13390 8290 13430 8295
rect 13390 8285 13395 8290
rect 13315 8265 13395 8285
rect 13315 8260 13320 8265
rect 13280 8255 13320 8260
rect 13390 8260 13395 8265
rect 13425 8285 13430 8290
rect 13500 8290 13540 8295
rect 13500 8285 13505 8290
rect 13425 8265 13505 8285
rect 13425 8260 13430 8265
rect 13390 8255 13430 8260
rect 13500 8260 13505 8265
rect 13535 8285 13540 8290
rect 13610 8290 13650 8295
rect 13610 8285 13615 8290
rect 13535 8265 13615 8285
rect 13535 8260 13540 8265
rect 13500 8255 13540 8260
rect 13610 8260 13615 8265
rect 13645 8285 13650 8290
rect 13720 8290 13760 8295
rect 13720 8285 13725 8290
rect 13645 8265 13725 8285
rect 13645 8260 13650 8265
rect 13610 8255 13650 8260
rect 13720 8260 13725 8265
rect 13755 8285 13760 8290
rect 13830 8290 13870 8295
rect 13830 8285 13835 8290
rect 13755 8265 13835 8285
rect 13755 8260 13760 8265
rect 13720 8255 13760 8260
rect 13830 8260 13835 8265
rect 13865 8285 13870 8290
rect 13940 8290 13980 8295
rect 13940 8285 13945 8290
rect 13865 8265 13945 8285
rect 13865 8260 13870 8265
rect 13830 8255 13870 8260
rect 13940 8260 13945 8265
rect 13975 8285 13980 8290
rect 14050 8290 14090 8295
rect 14050 8285 14055 8290
rect 13975 8265 14055 8285
rect 13975 8260 13980 8265
rect 13940 8255 13980 8260
rect 14050 8260 14055 8265
rect 14085 8260 14090 8290
rect 14050 8255 14090 8260
rect 20445 8290 20485 8295
rect 20445 8260 20450 8290
rect 20480 8285 20485 8290
rect 20555 8290 20595 8295
rect 20555 8285 20560 8290
rect 20480 8265 20560 8285
rect 20480 8260 20485 8265
rect 20445 8255 20485 8260
rect 20555 8260 20560 8265
rect 20590 8285 20595 8290
rect 20665 8290 20705 8295
rect 20665 8285 20670 8290
rect 20590 8265 20670 8285
rect 20590 8260 20595 8265
rect 20555 8255 20595 8260
rect 20665 8260 20670 8265
rect 20700 8285 20705 8290
rect 20775 8290 20815 8295
rect 20775 8285 20780 8290
rect 20700 8265 20780 8285
rect 20700 8260 20705 8265
rect 20665 8255 20705 8260
rect 20775 8260 20780 8265
rect 20810 8285 20815 8290
rect 20885 8290 20925 8295
rect 20885 8285 20890 8290
rect 20810 8265 20890 8285
rect 20810 8260 20815 8265
rect 20775 8255 20815 8260
rect 20885 8260 20890 8265
rect 20920 8285 20925 8290
rect 20995 8290 21035 8295
rect 20995 8285 21000 8290
rect 20920 8265 21000 8285
rect 20920 8260 20925 8265
rect 20885 8255 20925 8260
rect 20995 8260 21000 8265
rect 21030 8285 21035 8290
rect 21105 8290 21145 8295
rect 21105 8285 21110 8290
rect 21030 8265 21110 8285
rect 21030 8260 21035 8265
rect 20995 8255 21035 8260
rect 21105 8260 21110 8265
rect 21140 8285 21145 8290
rect 21215 8290 21255 8295
rect 21215 8285 21220 8290
rect 21140 8265 21220 8285
rect 21140 8260 21145 8265
rect 21105 8255 21145 8260
rect 21215 8260 21220 8265
rect 21250 8285 21255 8290
rect 21325 8290 21365 8295
rect 21325 8285 21330 8290
rect 21250 8265 21330 8285
rect 21250 8260 21255 8265
rect 21215 8255 21255 8260
rect 21325 8260 21330 8265
rect 21360 8285 21365 8290
rect 21435 8290 21475 8295
rect 21435 8285 21440 8290
rect 21360 8265 21440 8285
rect 21360 8260 21365 8265
rect 21325 8255 21365 8260
rect 21435 8260 21440 8265
rect 21470 8285 21475 8290
rect 21545 8290 21585 8295
rect 21545 8285 21550 8290
rect 21470 8265 21550 8285
rect 21470 8260 21475 8265
rect 21435 8255 21475 8260
rect 21545 8260 21550 8265
rect 21580 8260 21585 8290
rect 21545 8255 21585 8260
rect 10580 8210 10620 8215
rect 10580 8180 10585 8210
rect 10615 8205 10620 8210
rect 10980 8210 11015 8215
rect 10980 8205 10985 8210
rect 10615 8185 10985 8205
rect 10615 8180 10620 8185
rect 10580 8175 10620 8180
rect 10980 8180 10985 8185
rect 10980 8175 11015 8180
rect 18080 8210 18120 8215
rect 18080 8180 18085 8210
rect 18115 8205 18120 8210
rect 18480 8210 18515 8215
rect 18480 8205 18485 8210
rect 18115 8185 18485 8205
rect 18115 8180 18120 8185
rect 18080 8175 18120 8180
rect 18480 8180 18485 8185
rect 18480 8175 18515 8180
rect 10900 8155 10940 8160
rect 10900 8125 10905 8155
rect 10935 8150 10940 8155
rect 11823 8155 11857 8160
rect 11823 8150 11826 8155
rect 10935 8130 11826 8150
rect 10935 8125 10940 8130
rect 10900 8120 10940 8125
rect 11823 8125 11826 8130
rect 11854 8125 11857 8155
rect 11823 8120 11857 8125
rect 18400 8155 18440 8160
rect 18400 8125 18405 8155
rect 18435 8150 18440 8155
rect 19323 8155 19357 8160
rect 19323 8150 19326 8155
rect 18435 8130 19326 8150
rect 18435 8125 18440 8130
rect 18400 8120 18440 8125
rect 19323 8125 19326 8130
rect 19354 8125 19357 8155
rect 19323 8120 19357 8125
rect 11280 8100 11320 8105
rect 11280 8070 11285 8100
rect 11315 8095 11320 8100
rect 11520 8100 11560 8105
rect 11520 8095 11525 8100
rect 11315 8075 11525 8095
rect 11315 8070 11320 8075
rect 11280 8065 11320 8070
rect 11520 8070 11525 8075
rect 11555 8095 11560 8100
rect 11760 8100 11800 8105
rect 11760 8095 11765 8100
rect 11555 8075 11765 8095
rect 11555 8070 11560 8075
rect 11520 8065 11560 8070
rect 11760 8070 11765 8075
rect 11795 8095 11800 8100
rect 12000 8100 12040 8105
rect 12000 8095 12005 8100
rect 11795 8075 12005 8095
rect 11795 8070 11800 8075
rect 11760 8065 11800 8070
rect 12000 8070 12005 8075
rect 12035 8095 12040 8100
rect 12240 8100 12280 8105
rect 12240 8095 12245 8100
rect 12035 8075 12245 8095
rect 12035 8070 12040 8075
rect 12000 8065 12040 8070
rect 12240 8070 12245 8075
rect 12275 8095 12280 8100
rect 12480 8100 12520 8105
rect 12480 8095 12485 8100
rect 12275 8075 12485 8095
rect 12275 8070 12280 8075
rect 12240 8065 12280 8070
rect 12480 8070 12485 8075
rect 12515 8070 12520 8100
rect 12480 8065 12520 8070
rect 18780 8100 18820 8105
rect 18780 8070 18785 8100
rect 18815 8095 18820 8100
rect 19020 8100 19060 8105
rect 19020 8095 19025 8100
rect 18815 8075 19025 8095
rect 18815 8070 18820 8075
rect 18780 8065 18820 8070
rect 19020 8070 19025 8075
rect 19055 8095 19060 8100
rect 19260 8100 19300 8105
rect 19260 8095 19265 8100
rect 19055 8075 19265 8095
rect 19055 8070 19060 8075
rect 19020 8065 19060 8070
rect 19260 8070 19265 8075
rect 19295 8095 19300 8100
rect 19500 8100 19540 8105
rect 19500 8095 19505 8100
rect 19295 8075 19505 8095
rect 19295 8070 19300 8075
rect 19260 8065 19300 8070
rect 19500 8070 19505 8075
rect 19535 8095 19540 8100
rect 19740 8100 19780 8105
rect 19740 8095 19745 8100
rect 19535 8075 19745 8095
rect 19535 8070 19540 8075
rect 19500 8065 19540 8070
rect 19740 8070 19745 8075
rect 19775 8095 19780 8100
rect 19980 8100 20020 8105
rect 19980 8095 19985 8100
rect 19775 8075 19985 8095
rect 19775 8070 19780 8075
rect 19740 8065 19780 8070
rect 19980 8070 19985 8075
rect 20015 8070 20020 8100
rect 19980 8065 20020 8070
rect 11400 8055 11440 8060
rect 11400 8025 11405 8055
rect 11435 8050 11440 8055
rect 11640 8055 11680 8060
rect 11640 8050 11645 8055
rect 11435 8030 11645 8050
rect 11435 8025 11440 8030
rect 11400 8020 11440 8025
rect 11640 8025 11645 8030
rect 11675 8050 11680 8055
rect 11880 8055 11920 8060
rect 11880 8050 11885 8055
rect 11675 8030 11885 8050
rect 11675 8025 11680 8030
rect 11640 8020 11680 8025
rect 11880 8025 11885 8030
rect 11915 8050 11920 8055
rect 12120 8055 12160 8060
rect 12120 8050 12125 8055
rect 11915 8030 12125 8050
rect 11915 8025 11920 8030
rect 11880 8020 11920 8025
rect 12120 8025 12125 8030
rect 12155 8050 12160 8055
rect 12360 8055 12400 8060
rect 12360 8050 12365 8055
rect 12155 8030 12365 8050
rect 12155 8025 12160 8030
rect 12120 8020 12160 8025
rect 12360 8025 12365 8030
rect 12395 8025 12400 8055
rect 12360 8020 12400 8025
rect 18900 8055 18940 8060
rect 18900 8025 18905 8055
rect 18935 8050 18940 8055
rect 19140 8055 19180 8060
rect 19140 8050 19145 8055
rect 18935 8030 19145 8050
rect 18935 8025 18940 8030
rect 18900 8020 18940 8025
rect 19140 8025 19145 8030
rect 19175 8050 19180 8055
rect 19380 8055 19420 8060
rect 19380 8050 19385 8055
rect 19175 8030 19385 8050
rect 19175 8025 19180 8030
rect 19140 8020 19180 8025
rect 19380 8025 19385 8030
rect 19415 8050 19420 8055
rect 19620 8055 19660 8060
rect 19620 8050 19625 8055
rect 19415 8030 19625 8050
rect 19415 8025 19420 8030
rect 19380 8020 19420 8025
rect 19620 8025 19625 8030
rect 19655 8050 19660 8055
rect 19860 8055 19900 8060
rect 19860 8050 19865 8055
rect 19655 8030 19865 8050
rect 19655 8025 19660 8030
rect 19620 8020 19660 8025
rect 19860 8025 19865 8030
rect 19895 8025 19900 8055
rect 19860 8020 19900 8025
rect 11340 8000 11380 8005
rect 11340 7970 11345 8000
rect 11375 7995 11380 8000
rect 11400 8000 11440 8005
rect 11400 7995 11405 8000
rect 11375 7975 11405 7995
rect 11375 7970 11380 7975
rect 11340 7965 11380 7970
rect 11400 7970 11405 7975
rect 11435 7995 11440 8000
rect 11580 8000 11620 8005
rect 11580 7995 11585 8000
rect 11435 7975 11585 7995
rect 11435 7970 11440 7975
rect 11400 7965 11440 7970
rect 11580 7970 11585 7975
rect 11615 7995 11620 8000
rect 11820 8000 11860 8005
rect 11820 7995 11825 8000
rect 11615 7975 11825 7995
rect 11615 7970 11620 7975
rect 11580 7965 11620 7970
rect 11820 7970 11825 7975
rect 11855 7995 11860 8000
rect 12060 8000 12100 8005
rect 12060 7995 12065 8000
rect 11855 7975 12065 7995
rect 11855 7970 11860 7975
rect 11820 7965 11860 7970
rect 12060 7970 12065 7975
rect 12095 7995 12100 8000
rect 12300 8000 12340 8005
rect 12300 7995 12305 8000
rect 12095 7975 12305 7995
rect 12095 7970 12100 7975
rect 12060 7965 12100 7970
rect 12300 7970 12305 7975
rect 12335 7970 12340 8000
rect 12300 7965 12340 7970
rect 18840 8000 18880 8005
rect 18840 7970 18845 8000
rect 18875 7995 18880 8000
rect 18900 8000 18940 8005
rect 18900 7995 18905 8000
rect 18875 7975 18905 7995
rect 18875 7970 18880 7975
rect 18840 7965 18880 7970
rect 18900 7970 18905 7975
rect 18935 7995 18940 8000
rect 19080 8000 19120 8005
rect 19080 7995 19085 8000
rect 18935 7975 19085 7995
rect 18935 7970 18940 7975
rect 18900 7965 18940 7970
rect 19080 7970 19085 7975
rect 19115 7995 19120 8000
rect 19320 8000 19360 8005
rect 19320 7995 19325 8000
rect 19115 7975 19325 7995
rect 19115 7970 19120 7975
rect 19080 7965 19120 7970
rect 19320 7970 19325 7975
rect 19355 7995 19360 8000
rect 19560 8000 19600 8005
rect 19560 7995 19565 8000
rect 19355 7975 19565 7995
rect 19355 7970 19360 7975
rect 19320 7965 19360 7970
rect 19560 7970 19565 7975
rect 19595 7995 19600 8000
rect 19800 8000 19840 8005
rect 19800 7995 19805 8000
rect 19595 7975 19805 7995
rect 19595 7970 19600 7975
rect 19560 7965 19600 7970
rect 19800 7970 19805 7975
rect 19835 7970 19840 8000
rect 19800 7965 19840 7970
rect 11460 7945 11500 7950
rect 11460 7915 11465 7945
rect 11495 7940 11500 7945
rect 11700 7945 11740 7950
rect 11700 7940 11705 7945
rect 11495 7920 11705 7940
rect 11495 7915 11500 7920
rect 11460 7910 11500 7915
rect 11700 7915 11705 7920
rect 11735 7940 11740 7945
rect 11940 7945 11980 7950
rect 11940 7940 11945 7945
rect 11735 7920 11945 7940
rect 11735 7915 11740 7920
rect 11700 7910 11740 7915
rect 11940 7915 11945 7920
rect 11975 7940 11980 7945
rect 12180 7945 12220 7950
rect 12180 7940 12185 7945
rect 11975 7920 12185 7940
rect 11975 7915 11980 7920
rect 11940 7910 11980 7915
rect 12180 7915 12185 7920
rect 12215 7940 12220 7945
rect 12420 7945 12460 7950
rect 12420 7940 12425 7945
rect 12215 7920 12425 7940
rect 12215 7915 12220 7920
rect 12180 7910 12220 7915
rect 12420 7915 12425 7920
rect 12455 7940 12460 7945
rect 12480 7945 12520 7950
rect 12480 7940 12485 7945
rect 12455 7920 12485 7940
rect 12455 7915 12460 7920
rect 12420 7910 12460 7915
rect 12480 7915 12485 7920
rect 12515 7915 12520 7945
rect 18960 7945 19000 7950
rect 12480 7910 12520 7915
rect 13005 7920 13045 7925
rect 13005 7890 13010 7920
rect 13040 7915 13045 7920
rect 13115 7920 13155 7925
rect 13115 7915 13120 7920
rect 13040 7895 13120 7915
rect 13040 7890 13045 7895
rect 13005 7885 13045 7890
rect 13115 7890 13120 7895
rect 13150 7915 13155 7920
rect 13225 7920 13265 7925
rect 13225 7915 13230 7920
rect 13150 7895 13230 7915
rect 13150 7890 13155 7895
rect 13115 7885 13155 7890
rect 13225 7890 13230 7895
rect 13260 7915 13265 7920
rect 13335 7920 13375 7925
rect 13335 7915 13340 7920
rect 13260 7895 13340 7915
rect 13260 7890 13265 7895
rect 13225 7885 13265 7890
rect 13335 7890 13340 7895
rect 13370 7915 13375 7920
rect 13445 7920 13485 7925
rect 13445 7915 13450 7920
rect 13370 7895 13450 7915
rect 13370 7890 13375 7895
rect 13335 7885 13375 7890
rect 13445 7890 13450 7895
rect 13480 7915 13485 7920
rect 13555 7920 13595 7925
rect 13555 7915 13560 7920
rect 13480 7895 13560 7915
rect 13480 7890 13485 7895
rect 13445 7885 13485 7890
rect 13555 7890 13560 7895
rect 13590 7915 13595 7920
rect 13665 7920 13705 7925
rect 13665 7915 13670 7920
rect 13590 7895 13670 7915
rect 13590 7890 13595 7895
rect 13555 7885 13595 7890
rect 13665 7890 13670 7895
rect 13700 7915 13705 7920
rect 13775 7920 13815 7925
rect 13775 7915 13780 7920
rect 13700 7895 13780 7915
rect 13700 7890 13705 7895
rect 13665 7885 13705 7890
rect 13775 7890 13780 7895
rect 13810 7915 13815 7920
rect 13885 7920 13925 7925
rect 13885 7915 13890 7920
rect 13810 7895 13890 7915
rect 13810 7890 13815 7895
rect 13775 7885 13815 7890
rect 13885 7890 13890 7895
rect 13920 7915 13925 7920
rect 13995 7920 14035 7925
rect 13995 7915 14000 7920
rect 13920 7895 14000 7915
rect 13920 7890 13925 7895
rect 13885 7885 13925 7890
rect 13995 7890 14000 7895
rect 14030 7890 14035 7920
rect 18960 7915 18965 7945
rect 18995 7940 19000 7945
rect 19200 7945 19240 7950
rect 19200 7940 19205 7945
rect 18995 7920 19205 7940
rect 18995 7915 19000 7920
rect 18960 7910 19000 7915
rect 19200 7915 19205 7920
rect 19235 7940 19240 7945
rect 19440 7945 19480 7950
rect 19440 7940 19445 7945
rect 19235 7920 19445 7940
rect 19235 7915 19240 7920
rect 19200 7910 19240 7915
rect 19440 7915 19445 7920
rect 19475 7940 19480 7945
rect 19680 7945 19720 7950
rect 19680 7940 19685 7945
rect 19475 7920 19685 7940
rect 19475 7915 19480 7920
rect 19440 7910 19480 7915
rect 19680 7915 19685 7920
rect 19715 7940 19720 7945
rect 19920 7945 19960 7950
rect 19920 7940 19925 7945
rect 19715 7920 19925 7940
rect 19715 7915 19720 7920
rect 19680 7910 19720 7915
rect 19920 7915 19925 7920
rect 19955 7940 19960 7945
rect 19980 7945 20020 7950
rect 19980 7940 19985 7945
rect 19955 7920 19985 7940
rect 19955 7915 19960 7920
rect 19920 7910 19960 7915
rect 19980 7915 19985 7920
rect 20015 7915 20020 7945
rect 19980 7910 20020 7915
rect 20500 7920 20540 7925
rect 13995 7885 14035 7890
rect 20500 7890 20505 7920
rect 20535 7915 20540 7920
rect 20610 7920 20650 7925
rect 20610 7915 20615 7920
rect 20535 7895 20615 7915
rect 20535 7890 20540 7895
rect 20500 7885 20540 7890
rect 20610 7890 20615 7895
rect 20645 7915 20650 7920
rect 20720 7920 20760 7925
rect 20720 7915 20725 7920
rect 20645 7895 20725 7915
rect 20645 7890 20650 7895
rect 20610 7885 20650 7890
rect 20720 7890 20725 7895
rect 20755 7915 20760 7920
rect 20830 7920 20870 7925
rect 20830 7915 20835 7920
rect 20755 7895 20835 7915
rect 20755 7890 20760 7895
rect 20720 7885 20760 7890
rect 20830 7890 20835 7895
rect 20865 7915 20870 7920
rect 20940 7920 20980 7925
rect 20940 7915 20945 7920
rect 20865 7895 20945 7915
rect 20865 7890 20870 7895
rect 20830 7885 20870 7890
rect 20940 7890 20945 7895
rect 20975 7915 20980 7920
rect 21050 7920 21090 7925
rect 21050 7915 21055 7920
rect 20975 7895 21055 7915
rect 20975 7890 20980 7895
rect 20940 7885 20980 7890
rect 21050 7890 21055 7895
rect 21085 7915 21090 7920
rect 21160 7920 21200 7925
rect 21160 7915 21165 7920
rect 21085 7895 21165 7915
rect 21085 7890 21090 7895
rect 21050 7885 21090 7890
rect 21160 7890 21165 7895
rect 21195 7915 21200 7920
rect 21270 7920 21310 7925
rect 21270 7915 21275 7920
rect 21195 7895 21275 7915
rect 21195 7890 21200 7895
rect 21160 7885 21200 7890
rect 21270 7890 21275 7895
rect 21305 7915 21310 7920
rect 21380 7920 21420 7925
rect 21380 7915 21385 7920
rect 21305 7895 21385 7915
rect 21305 7890 21310 7895
rect 21270 7885 21310 7890
rect 21380 7890 21385 7895
rect 21415 7915 21420 7920
rect 21490 7920 21530 7925
rect 21490 7915 21495 7920
rect 21415 7895 21495 7915
rect 21415 7890 21420 7895
rect 21380 7885 21420 7890
rect 21490 7890 21495 7895
rect 21525 7890 21530 7920
rect 21490 7885 21530 7890
rect 13060 7830 13100 7836
rect 13060 7800 13065 7830
rect 13095 7800 13100 7830
rect 13060 7780 13100 7800
rect 13060 7750 13065 7780
rect 13095 7750 13100 7780
rect 12690 7730 12730 7735
rect 12690 7700 12695 7730
rect 12725 7725 12730 7730
rect 13060 7730 13100 7750
rect 13060 7725 13065 7730
rect 12725 7705 13065 7725
rect 12725 7700 12730 7705
rect 12690 7695 12730 7700
rect 13060 7700 13065 7705
rect 13095 7700 13100 7730
rect 13060 7695 13100 7700
rect 13680 7830 13720 7836
rect 13680 7800 13685 7830
rect 13715 7800 13720 7830
rect 13680 7780 13720 7800
rect 13680 7750 13685 7780
rect 13715 7775 13720 7780
rect 20555 7830 20595 7836
rect 20555 7800 20560 7830
rect 20590 7800 20595 7830
rect 20555 7780 20595 7800
rect 13715 7755 14385 7775
rect 13715 7750 13720 7755
rect 13680 7730 13720 7750
rect 20555 7750 20560 7780
rect 20590 7750 20595 7780
rect 13680 7700 13685 7730
rect 13715 7700 13720 7730
rect 13680 7695 13720 7700
rect 20190 7730 20230 7735
rect 20190 7700 20195 7730
rect 20225 7725 20230 7730
rect 20555 7730 20595 7750
rect 20555 7725 20560 7730
rect 20225 7705 20560 7725
rect 20225 7700 20230 7705
rect 20190 7695 20230 7700
rect 20555 7700 20560 7705
rect 20590 7700 20595 7730
rect 20555 7695 20595 7700
rect 9735 7670 9775 7675
rect 9735 7640 9740 7670
rect 9770 7665 9775 7670
rect 9845 7670 9885 7675
rect 9845 7665 9850 7670
rect 9770 7645 9850 7665
rect 9770 7640 9775 7645
rect 9735 7635 9775 7640
rect 9845 7640 9850 7645
rect 9880 7665 9885 7670
rect 9955 7670 9995 7675
rect 9955 7665 9960 7670
rect 9880 7645 9960 7665
rect 9880 7640 9885 7645
rect 9845 7635 9885 7640
rect 9955 7640 9960 7645
rect 9990 7665 9995 7670
rect 10065 7670 10105 7675
rect 10065 7665 10070 7670
rect 9990 7645 10070 7665
rect 9990 7640 9995 7645
rect 9955 7635 9995 7640
rect 10065 7640 10070 7645
rect 10100 7665 10105 7670
rect 10175 7670 10215 7675
rect 10175 7665 10180 7670
rect 10100 7645 10180 7665
rect 10100 7640 10105 7645
rect 10065 7635 10105 7640
rect 10175 7640 10180 7645
rect 10210 7665 10215 7670
rect 10285 7670 10325 7675
rect 10285 7665 10290 7670
rect 10210 7645 10290 7665
rect 10210 7640 10215 7645
rect 10175 7635 10215 7640
rect 10285 7640 10290 7645
rect 10320 7665 10325 7670
rect 10395 7670 10435 7675
rect 10395 7665 10400 7670
rect 10320 7645 10400 7665
rect 10320 7640 10325 7645
rect 10285 7635 10325 7640
rect 10395 7640 10400 7645
rect 10430 7665 10435 7670
rect 10505 7670 10545 7675
rect 10505 7665 10510 7670
rect 10430 7645 10510 7665
rect 10430 7640 10435 7645
rect 10395 7635 10435 7640
rect 10505 7640 10510 7645
rect 10540 7665 10545 7670
rect 10615 7670 10655 7675
rect 10615 7665 10620 7670
rect 10540 7645 10620 7665
rect 10540 7640 10545 7645
rect 10505 7635 10545 7640
rect 10615 7640 10620 7645
rect 10650 7665 10655 7670
rect 10725 7670 10765 7675
rect 10725 7665 10730 7670
rect 10650 7645 10730 7665
rect 10650 7640 10655 7645
rect 10615 7635 10655 7640
rect 10725 7640 10730 7645
rect 10760 7665 10765 7670
rect 10835 7670 10875 7675
rect 10835 7665 10840 7670
rect 10760 7645 10840 7665
rect 10760 7640 10765 7645
rect 10725 7635 10765 7640
rect 10835 7640 10840 7645
rect 10870 7640 10875 7670
rect 10835 7635 10875 7640
rect 12950 7670 12990 7675
rect 12950 7640 12955 7670
rect 12985 7665 12990 7670
rect 13060 7670 13100 7675
rect 13060 7665 13065 7670
rect 12985 7645 13065 7665
rect 12985 7640 12990 7645
rect 12950 7635 12990 7640
rect 13060 7640 13065 7645
rect 13095 7665 13100 7670
rect 13170 7670 13210 7675
rect 13170 7665 13175 7670
rect 13095 7645 13175 7665
rect 13095 7640 13100 7645
rect 13060 7635 13100 7640
rect 13170 7640 13175 7645
rect 13205 7665 13210 7670
rect 13280 7670 13320 7675
rect 13280 7665 13285 7670
rect 13205 7645 13285 7665
rect 13205 7640 13210 7645
rect 13170 7635 13210 7640
rect 13280 7640 13285 7645
rect 13315 7665 13320 7670
rect 13390 7670 13430 7675
rect 13390 7665 13395 7670
rect 13315 7645 13395 7665
rect 13315 7640 13320 7645
rect 13280 7635 13320 7640
rect 13390 7640 13395 7645
rect 13425 7665 13430 7670
rect 13500 7670 13540 7675
rect 13500 7665 13505 7670
rect 13425 7645 13505 7665
rect 13425 7640 13430 7645
rect 13390 7635 13430 7640
rect 13500 7640 13505 7645
rect 13535 7665 13540 7670
rect 13610 7670 13650 7675
rect 13610 7665 13615 7670
rect 13535 7645 13615 7665
rect 13535 7640 13540 7645
rect 13500 7635 13540 7640
rect 13610 7640 13615 7645
rect 13645 7665 13650 7670
rect 13720 7670 13760 7675
rect 13720 7665 13725 7670
rect 13645 7645 13725 7665
rect 13645 7640 13650 7645
rect 13610 7635 13650 7640
rect 13720 7640 13725 7645
rect 13755 7665 13760 7670
rect 13830 7670 13870 7675
rect 13830 7665 13835 7670
rect 13755 7645 13835 7665
rect 13755 7640 13760 7645
rect 13720 7635 13760 7640
rect 13830 7640 13835 7645
rect 13865 7665 13870 7670
rect 13940 7670 13980 7675
rect 13940 7665 13945 7670
rect 13865 7645 13945 7665
rect 13865 7640 13870 7645
rect 13830 7635 13870 7640
rect 13940 7640 13945 7645
rect 13975 7665 13980 7670
rect 14050 7670 14090 7675
rect 14050 7665 14055 7670
rect 13975 7645 14055 7665
rect 13975 7640 13980 7645
rect 13940 7635 13980 7640
rect 14050 7640 14055 7645
rect 14085 7640 14090 7670
rect 14050 7635 14090 7640
rect 17235 7670 17275 7675
rect 17235 7640 17240 7670
rect 17270 7665 17275 7670
rect 17345 7670 17385 7675
rect 17345 7665 17350 7670
rect 17270 7645 17350 7665
rect 17270 7640 17275 7645
rect 17235 7635 17275 7640
rect 17345 7640 17350 7645
rect 17380 7665 17385 7670
rect 17455 7670 17495 7675
rect 17455 7665 17460 7670
rect 17380 7645 17460 7665
rect 17380 7640 17385 7645
rect 17345 7635 17385 7640
rect 17455 7640 17460 7645
rect 17490 7665 17495 7670
rect 17565 7670 17605 7675
rect 17565 7665 17570 7670
rect 17490 7645 17570 7665
rect 17490 7640 17495 7645
rect 17455 7635 17495 7640
rect 17565 7640 17570 7645
rect 17600 7665 17605 7670
rect 17675 7670 17715 7675
rect 17675 7665 17680 7670
rect 17600 7645 17680 7665
rect 17600 7640 17605 7645
rect 17565 7635 17605 7640
rect 17675 7640 17680 7645
rect 17710 7665 17715 7670
rect 17785 7670 17825 7675
rect 17785 7665 17790 7670
rect 17710 7645 17790 7665
rect 17710 7640 17715 7645
rect 17675 7635 17715 7640
rect 17785 7640 17790 7645
rect 17820 7665 17825 7670
rect 17895 7670 17935 7675
rect 17895 7665 17900 7670
rect 17820 7645 17900 7665
rect 17820 7640 17825 7645
rect 17785 7635 17825 7640
rect 17895 7640 17900 7645
rect 17930 7665 17935 7670
rect 18005 7670 18045 7675
rect 18005 7665 18010 7670
rect 17930 7645 18010 7665
rect 17930 7640 17935 7645
rect 17895 7635 17935 7640
rect 18005 7640 18010 7645
rect 18040 7665 18045 7670
rect 18115 7670 18155 7675
rect 18115 7665 18120 7670
rect 18040 7645 18120 7665
rect 18040 7640 18045 7645
rect 18005 7635 18045 7640
rect 18115 7640 18120 7645
rect 18150 7665 18155 7670
rect 18225 7670 18265 7675
rect 18225 7665 18230 7670
rect 18150 7645 18230 7665
rect 18150 7640 18155 7645
rect 18115 7635 18155 7640
rect 18225 7640 18230 7645
rect 18260 7665 18265 7670
rect 18335 7670 18375 7675
rect 18335 7665 18340 7670
rect 18260 7645 18340 7665
rect 18260 7640 18265 7645
rect 18225 7635 18265 7640
rect 18335 7640 18340 7645
rect 18370 7640 18375 7670
rect 18335 7635 18375 7640
rect 20445 7670 20485 7675
rect 20445 7640 20450 7670
rect 20480 7665 20485 7670
rect 20555 7670 20595 7675
rect 20555 7665 20560 7670
rect 20480 7645 20560 7665
rect 20480 7640 20485 7645
rect 20445 7635 20485 7640
rect 20555 7640 20560 7645
rect 20590 7665 20595 7670
rect 20665 7670 20705 7675
rect 20665 7665 20670 7670
rect 20590 7645 20670 7665
rect 20590 7640 20595 7645
rect 20555 7635 20595 7640
rect 20665 7640 20670 7645
rect 20700 7665 20705 7670
rect 20775 7670 20815 7675
rect 20775 7665 20780 7670
rect 20700 7645 20780 7665
rect 20700 7640 20705 7645
rect 20665 7635 20705 7640
rect 20775 7640 20780 7645
rect 20810 7665 20815 7670
rect 20885 7670 20925 7675
rect 20885 7665 20890 7670
rect 20810 7645 20890 7665
rect 20810 7640 20815 7645
rect 20775 7635 20815 7640
rect 20885 7640 20890 7645
rect 20920 7665 20925 7670
rect 20995 7670 21035 7675
rect 20995 7665 21000 7670
rect 20920 7645 21000 7665
rect 20920 7640 20925 7645
rect 20885 7635 20925 7640
rect 20995 7640 21000 7645
rect 21030 7665 21035 7670
rect 21105 7670 21145 7675
rect 21105 7665 21110 7670
rect 21030 7645 21110 7665
rect 21030 7640 21035 7645
rect 20995 7635 21035 7640
rect 21105 7640 21110 7645
rect 21140 7665 21145 7670
rect 21215 7670 21255 7675
rect 21215 7665 21220 7670
rect 21140 7645 21220 7665
rect 21140 7640 21145 7645
rect 21105 7635 21145 7640
rect 21215 7640 21220 7645
rect 21250 7665 21255 7670
rect 21325 7670 21365 7675
rect 21325 7665 21330 7670
rect 21250 7645 21330 7665
rect 21250 7640 21255 7645
rect 21215 7635 21255 7640
rect 21325 7640 21330 7645
rect 21360 7665 21365 7670
rect 21435 7670 21475 7675
rect 21435 7665 21440 7670
rect 21360 7645 21440 7665
rect 21360 7640 21365 7645
rect 21325 7635 21365 7640
rect 21435 7640 21440 7645
rect 21470 7665 21475 7670
rect 21545 7670 21585 7675
rect 21545 7665 21550 7670
rect 21470 7645 21550 7665
rect 21470 7640 21475 7645
rect 21435 7635 21475 7640
rect 21545 7640 21550 7645
rect 21580 7640 21585 7670
rect 21545 7635 21585 7640
rect 9790 7500 9830 7505
rect 9790 7470 9795 7500
rect 9825 7495 9830 7500
rect 9900 7500 9940 7505
rect 9900 7495 9905 7500
rect 9825 7475 9905 7495
rect 9825 7470 9830 7475
rect 9790 7465 9830 7470
rect 9900 7470 9905 7475
rect 9935 7495 9940 7500
rect 10010 7500 10050 7505
rect 10010 7495 10015 7500
rect 9935 7475 10015 7495
rect 9935 7470 9940 7475
rect 9900 7465 9940 7470
rect 10010 7470 10015 7475
rect 10045 7495 10050 7500
rect 10120 7500 10160 7505
rect 10120 7495 10125 7500
rect 10045 7475 10125 7495
rect 10045 7470 10050 7475
rect 10010 7465 10050 7470
rect 10120 7470 10125 7475
rect 10155 7495 10160 7500
rect 10230 7500 10270 7505
rect 10230 7495 10235 7500
rect 10155 7475 10235 7495
rect 10155 7470 10160 7475
rect 10120 7465 10160 7470
rect 10230 7470 10235 7475
rect 10265 7495 10270 7500
rect 10340 7500 10380 7505
rect 10340 7495 10345 7500
rect 10265 7475 10345 7495
rect 10265 7470 10270 7475
rect 10230 7465 10270 7470
rect 10340 7470 10345 7475
rect 10375 7495 10380 7500
rect 10450 7500 10490 7505
rect 10450 7495 10455 7500
rect 10375 7475 10455 7495
rect 10375 7470 10380 7475
rect 10340 7465 10380 7470
rect 10450 7470 10455 7475
rect 10485 7495 10490 7500
rect 10560 7500 10600 7505
rect 10560 7495 10565 7500
rect 10485 7475 10565 7495
rect 10485 7470 10490 7475
rect 10450 7465 10490 7470
rect 10560 7470 10565 7475
rect 10595 7495 10600 7500
rect 10670 7500 10710 7505
rect 10670 7495 10675 7500
rect 10595 7475 10675 7495
rect 10595 7470 10600 7475
rect 10560 7465 10600 7470
rect 10670 7470 10675 7475
rect 10705 7495 10710 7500
rect 10780 7500 10820 7505
rect 10780 7495 10785 7500
rect 10705 7475 10785 7495
rect 10705 7470 10710 7475
rect 10670 7465 10710 7470
rect 10780 7470 10785 7475
rect 10815 7470 10820 7500
rect 13005 7500 13045 7505
rect 10780 7465 10820 7470
rect 10980 7475 11020 7480
rect 10980 7445 10985 7475
rect 11015 7470 11020 7475
rect 11823 7475 11857 7480
rect 11823 7470 11826 7475
rect 11015 7450 11826 7470
rect 11015 7445 11020 7450
rect 10813 7440 10847 7445
rect 10980 7440 11020 7445
rect 11823 7445 11826 7450
rect 11854 7445 11857 7475
rect 13005 7470 13010 7500
rect 13040 7495 13045 7500
rect 13115 7500 13155 7505
rect 13115 7495 13120 7500
rect 13040 7475 13120 7495
rect 13040 7470 13045 7475
rect 13005 7465 13045 7470
rect 13115 7470 13120 7475
rect 13150 7495 13155 7500
rect 13225 7500 13265 7505
rect 13225 7495 13230 7500
rect 13150 7475 13230 7495
rect 13150 7470 13155 7475
rect 13115 7465 13155 7470
rect 13225 7470 13230 7475
rect 13260 7495 13265 7500
rect 13335 7500 13375 7505
rect 13335 7495 13340 7500
rect 13260 7475 13340 7495
rect 13260 7470 13265 7475
rect 13225 7465 13265 7470
rect 13335 7470 13340 7475
rect 13370 7495 13375 7500
rect 13445 7500 13485 7505
rect 13445 7495 13450 7500
rect 13370 7475 13450 7495
rect 13370 7470 13375 7475
rect 13335 7465 13375 7470
rect 13445 7470 13450 7475
rect 13480 7495 13485 7500
rect 13555 7500 13595 7505
rect 13555 7495 13560 7500
rect 13480 7475 13560 7495
rect 13480 7470 13485 7475
rect 13445 7465 13485 7470
rect 13555 7470 13560 7475
rect 13590 7495 13595 7500
rect 13665 7500 13705 7505
rect 13665 7495 13670 7500
rect 13590 7475 13670 7495
rect 13590 7470 13595 7475
rect 13555 7465 13595 7470
rect 13665 7470 13670 7475
rect 13700 7495 13705 7500
rect 13775 7500 13815 7505
rect 13775 7495 13780 7500
rect 13700 7475 13780 7495
rect 13700 7470 13705 7475
rect 13665 7465 13705 7470
rect 13775 7470 13780 7475
rect 13810 7495 13815 7500
rect 13885 7500 13925 7505
rect 13885 7495 13890 7500
rect 13810 7475 13890 7495
rect 13810 7470 13815 7475
rect 13775 7465 13815 7470
rect 13885 7470 13890 7475
rect 13920 7495 13925 7500
rect 13995 7500 14035 7505
rect 13995 7495 14000 7500
rect 13920 7475 14000 7495
rect 13920 7470 13925 7475
rect 13885 7465 13925 7470
rect 13995 7470 14000 7475
rect 14030 7470 14035 7500
rect 13995 7465 14035 7470
rect 17290 7500 17330 7505
rect 17290 7470 17295 7500
rect 17325 7495 17330 7500
rect 17400 7500 17440 7505
rect 17400 7495 17405 7500
rect 17325 7475 17405 7495
rect 17325 7470 17330 7475
rect 17290 7465 17330 7470
rect 17400 7470 17405 7475
rect 17435 7495 17440 7500
rect 17510 7500 17550 7505
rect 17510 7495 17515 7500
rect 17435 7475 17515 7495
rect 17435 7470 17440 7475
rect 17400 7465 17440 7470
rect 17510 7470 17515 7475
rect 17545 7495 17550 7500
rect 17620 7500 17660 7505
rect 17620 7495 17625 7500
rect 17545 7475 17625 7495
rect 17545 7470 17550 7475
rect 17510 7465 17550 7470
rect 17620 7470 17625 7475
rect 17655 7495 17660 7500
rect 17730 7500 17770 7505
rect 17730 7495 17735 7500
rect 17655 7475 17735 7495
rect 17655 7470 17660 7475
rect 17620 7465 17660 7470
rect 17730 7470 17735 7475
rect 17765 7495 17770 7500
rect 17840 7500 17880 7505
rect 17840 7495 17845 7500
rect 17765 7475 17845 7495
rect 17765 7470 17770 7475
rect 17730 7465 17770 7470
rect 17840 7470 17845 7475
rect 17875 7495 17880 7500
rect 17950 7500 17990 7505
rect 17950 7495 17955 7500
rect 17875 7475 17955 7495
rect 17875 7470 17880 7475
rect 17840 7465 17880 7470
rect 17950 7470 17955 7475
rect 17985 7495 17990 7500
rect 18060 7500 18100 7505
rect 18060 7495 18065 7500
rect 17985 7475 18065 7495
rect 17985 7470 17990 7475
rect 17950 7465 17990 7470
rect 18060 7470 18065 7475
rect 18095 7495 18100 7500
rect 18170 7500 18210 7505
rect 18170 7495 18175 7500
rect 18095 7475 18175 7495
rect 18095 7470 18100 7475
rect 18060 7465 18100 7470
rect 18170 7470 18175 7475
rect 18205 7495 18210 7500
rect 18280 7500 18320 7505
rect 18280 7495 18285 7500
rect 18205 7475 18285 7495
rect 18205 7470 18210 7475
rect 18170 7465 18210 7470
rect 18280 7470 18285 7475
rect 18315 7470 18320 7500
rect 20500 7500 20540 7505
rect 18280 7465 18320 7470
rect 18480 7475 18520 7480
rect 18480 7445 18485 7475
rect 18515 7470 18520 7475
rect 19323 7475 19357 7480
rect 19323 7470 19326 7475
rect 18515 7450 19326 7470
rect 18515 7445 18520 7450
rect 11823 7440 11857 7445
rect 12978 7440 13012 7445
rect 10813 7410 10816 7440
rect 10844 7425 10847 7440
rect 10844 7420 11320 7425
rect 10844 7410 11285 7420
rect 10813 7405 11285 7410
rect 11280 7390 11285 7405
rect 11315 7415 11320 7420
rect 11520 7420 11560 7425
rect 11520 7415 11525 7420
rect 11315 7395 11525 7415
rect 11315 7390 11320 7395
rect 11280 7385 11320 7390
rect 11520 7390 11525 7395
rect 11555 7415 11560 7420
rect 11760 7420 11800 7425
rect 11760 7415 11765 7420
rect 11555 7395 11765 7415
rect 11555 7390 11560 7395
rect 11520 7385 11560 7390
rect 11760 7390 11765 7395
rect 11795 7415 11800 7420
rect 12000 7420 12040 7425
rect 12000 7415 12005 7420
rect 11795 7395 12005 7415
rect 11795 7390 11800 7395
rect 11760 7385 11800 7390
rect 12000 7390 12005 7395
rect 12035 7415 12040 7420
rect 12240 7420 12280 7425
rect 12240 7415 12245 7420
rect 12035 7395 12245 7415
rect 12035 7390 12040 7395
rect 12000 7385 12040 7390
rect 12240 7390 12245 7395
rect 12275 7415 12280 7420
rect 12480 7420 12520 7425
rect 12480 7415 12485 7420
rect 12275 7395 12485 7415
rect 12275 7390 12280 7395
rect 12240 7385 12280 7390
rect 12480 7390 12485 7395
rect 12515 7390 12520 7420
rect 12978 7410 12981 7440
rect 13009 7410 13012 7440
rect 12978 7405 13012 7410
rect 18313 7440 18347 7445
rect 18480 7440 18520 7445
rect 19323 7445 19326 7450
rect 19354 7445 19357 7475
rect 20500 7470 20505 7500
rect 20535 7495 20540 7500
rect 20610 7500 20650 7505
rect 20610 7495 20615 7500
rect 20535 7475 20615 7495
rect 20535 7470 20540 7475
rect 20500 7465 20540 7470
rect 20610 7470 20615 7475
rect 20645 7495 20650 7500
rect 20720 7500 20760 7505
rect 20720 7495 20725 7500
rect 20645 7475 20725 7495
rect 20645 7470 20650 7475
rect 20610 7465 20650 7470
rect 20720 7470 20725 7475
rect 20755 7495 20760 7500
rect 20830 7500 20870 7505
rect 20830 7495 20835 7500
rect 20755 7475 20835 7495
rect 20755 7470 20760 7475
rect 20720 7465 20760 7470
rect 20830 7470 20835 7475
rect 20865 7495 20870 7500
rect 20940 7500 20980 7505
rect 20940 7495 20945 7500
rect 20865 7475 20945 7495
rect 20865 7470 20870 7475
rect 20830 7465 20870 7470
rect 20940 7470 20945 7475
rect 20975 7495 20980 7500
rect 21050 7500 21090 7505
rect 21050 7495 21055 7500
rect 20975 7475 21055 7495
rect 20975 7470 20980 7475
rect 20940 7465 20980 7470
rect 21050 7470 21055 7475
rect 21085 7495 21090 7500
rect 21160 7500 21200 7505
rect 21160 7495 21165 7500
rect 21085 7475 21165 7495
rect 21085 7470 21090 7475
rect 21050 7465 21090 7470
rect 21160 7470 21165 7475
rect 21195 7495 21200 7500
rect 21270 7500 21310 7505
rect 21270 7495 21275 7500
rect 21195 7475 21275 7495
rect 21195 7470 21200 7475
rect 21160 7465 21200 7470
rect 21270 7470 21275 7475
rect 21305 7495 21310 7500
rect 21380 7500 21420 7505
rect 21380 7495 21385 7500
rect 21305 7475 21385 7495
rect 21305 7470 21310 7475
rect 21270 7465 21310 7470
rect 21380 7470 21385 7475
rect 21415 7495 21420 7500
rect 21490 7500 21530 7505
rect 21490 7495 21495 7500
rect 21415 7475 21495 7495
rect 21415 7470 21420 7475
rect 21380 7465 21420 7470
rect 21490 7470 21495 7475
rect 21525 7470 21530 7500
rect 21490 7465 21530 7470
rect 19323 7440 19357 7445
rect 20473 7440 20507 7445
rect 18313 7410 18316 7440
rect 18344 7425 18347 7440
rect 18344 7420 18820 7425
rect 18344 7410 18785 7420
rect 18313 7405 18785 7410
rect 12480 7385 12520 7390
rect 18780 7390 18785 7405
rect 18815 7415 18820 7420
rect 19020 7420 19060 7425
rect 19020 7415 19025 7420
rect 18815 7395 19025 7415
rect 18815 7390 18820 7395
rect 18780 7385 18820 7390
rect 19020 7390 19025 7395
rect 19055 7415 19060 7420
rect 19260 7420 19300 7425
rect 19260 7415 19265 7420
rect 19055 7395 19265 7415
rect 19055 7390 19060 7395
rect 19020 7385 19060 7390
rect 19260 7390 19265 7395
rect 19295 7415 19300 7420
rect 19500 7420 19540 7425
rect 19500 7415 19505 7420
rect 19295 7395 19505 7415
rect 19295 7390 19300 7395
rect 19260 7385 19300 7390
rect 19500 7390 19505 7395
rect 19535 7415 19540 7420
rect 19740 7420 19780 7425
rect 19740 7415 19745 7420
rect 19535 7395 19745 7415
rect 19535 7390 19540 7395
rect 19500 7385 19540 7390
rect 19740 7390 19745 7395
rect 19775 7415 19780 7420
rect 19980 7420 20020 7425
rect 19980 7415 19985 7420
rect 19775 7395 19985 7415
rect 19775 7390 19780 7395
rect 19740 7385 19780 7390
rect 19980 7390 19985 7395
rect 20015 7390 20020 7420
rect 20473 7410 20476 7440
rect 20504 7410 20507 7440
rect 20473 7405 20507 7410
rect 19980 7385 20020 7390
rect 9800 7345 9805 7380
rect 9840 7345 9845 7380
rect 10635 7345 10640 7380
rect 10675 7345 10680 7380
rect 11400 7375 11440 7380
rect 11400 7345 11405 7375
rect 11435 7370 11440 7375
rect 11640 7375 11680 7380
rect 11640 7370 11645 7375
rect 11435 7350 11645 7370
rect 11435 7345 11440 7350
rect 11400 7340 11440 7345
rect 11640 7345 11645 7350
rect 11675 7370 11680 7375
rect 11880 7375 11920 7380
rect 11880 7370 11885 7375
rect 11675 7350 11885 7370
rect 11675 7345 11680 7350
rect 11640 7340 11680 7345
rect 11880 7345 11885 7350
rect 11915 7370 11920 7375
rect 12120 7375 12160 7380
rect 12120 7370 12125 7375
rect 11915 7350 12125 7370
rect 11915 7345 11920 7350
rect 11880 7340 11920 7345
rect 12120 7345 12125 7350
rect 12155 7370 12160 7375
rect 12360 7375 12400 7380
rect 12360 7370 12365 7375
rect 12155 7350 12365 7370
rect 12155 7345 12160 7350
rect 12120 7340 12160 7345
rect 12360 7345 12365 7350
rect 12395 7370 12400 7375
rect 12690 7375 12730 7380
rect 12690 7370 12695 7375
rect 12395 7350 12695 7370
rect 12395 7345 12400 7350
rect 12360 7340 12400 7345
rect 12690 7345 12695 7350
rect 12725 7370 12730 7375
rect 12975 7375 13015 7380
rect 12975 7370 12980 7375
rect 12725 7350 12980 7370
rect 12725 7345 12730 7350
rect 12690 7340 12730 7345
rect 12975 7345 12980 7350
rect 13010 7345 13015 7375
rect 13145 7345 13150 7380
rect 13185 7345 13190 7380
rect 13979 7345 13985 7380
rect 14020 7345 14025 7380
rect 17300 7345 17305 7380
rect 17340 7345 17345 7380
rect 18135 7345 18140 7380
rect 18175 7345 18180 7380
rect 18900 7375 18940 7380
rect 18900 7345 18905 7375
rect 18935 7370 18940 7375
rect 19140 7375 19180 7380
rect 19140 7370 19145 7375
rect 18935 7350 19145 7370
rect 18935 7345 18940 7350
rect 12975 7340 13015 7345
rect 18900 7340 18940 7345
rect 19140 7345 19145 7350
rect 19175 7370 19180 7375
rect 19380 7375 19420 7380
rect 19380 7370 19385 7375
rect 19175 7350 19385 7370
rect 19175 7345 19180 7350
rect 19140 7340 19180 7345
rect 19380 7345 19385 7350
rect 19415 7370 19420 7375
rect 19620 7375 19660 7380
rect 19620 7370 19625 7375
rect 19415 7350 19625 7370
rect 19415 7345 19420 7350
rect 19380 7340 19420 7345
rect 19620 7345 19625 7350
rect 19655 7370 19660 7375
rect 19860 7375 19900 7380
rect 19860 7370 19865 7375
rect 19655 7350 19865 7370
rect 19655 7345 19660 7350
rect 19620 7340 19660 7345
rect 19860 7345 19865 7350
rect 19895 7370 19900 7375
rect 20190 7375 20230 7380
rect 20190 7370 20195 7375
rect 19895 7350 20195 7370
rect 19895 7345 19900 7350
rect 19860 7340 19900 7345
rect 20190 7345 20195 7350
rect 20225 7370 20230 7375
rect 20470 7375 20510 7380
rect 20470 7370 20475 7375
rect 20225 7350 20475 7370
rect 20225 7345 20230 7350
rect 20190 7340 20230 7345
rect 20470 7345 20475 7350
rect 20505 7345 20510 7375
rect 20640 7345 20645 7380
rect 20680 7345 20685 7380
rect 21474 7345 21480 7380
rect 21515 7345 21520 7380
rect 20470 7340 20510 7345
rect 12815 7325 12855 7330
rect 12815 7320 12820 7325
rect 9800 7285 9805 7320
rect 9840 7285 9845 7320
rect 10635 7285 10640 7320
rect 10675 7300 12820 7320
rect 10675 7285 10680 7300
rect 12815 7295 12820 7300
rect 12850 7320 12855 7325
rect 20315 7325 20355 7330
rect 20315 7320 20320 7325
rect 12850 7300 13150 7320
rect 12850 7295 12855 7300
rect 12815 7290 12855 7295
rect 13145 7285 13150 7300
rect 13185 7285 13190 7320
rect 13980 7285 13985 7320
rect 14020 7285 14025 7320
rect 17300 7285 17305 7320
rect 17340 7285 17345 7320
rect 18135 7285 18140 7320
rect 18175 7300 20320 7320
rect 18175 7285 18180 7300
rect 20315 7295 20320 7300
rect 20350 7320 20355 7325
rect 20350 7300 20645 7320
rect 20350 7295 20355 7300
rect 20315 7290 20355 7295
rect 20640 7285 20645 7300
rect 20680 7285 20685 7320
rect 21475 7285 21480 7320
rect 21515 7285 21520 7320
rect 10813 7280 10847 7285
rect 10813 7250 10816 7280
rect 10844 7250 10847 7280
rect 10813 7245 10847 7250
rect 11440 7280 11480 7285
rect 11440 7250 11445 7280
rect 11475 7275 11480 7280
rect 11660 7280 11700 7285
rect 11660 7275 11665 7280
rect 11475 7255 11665 7275
rect 11475 7250 11480 7255
rect 11440 7245 11480 7250
rect 11660 7250 11665 7255
rect 11695 7275 11700 7280
rect 11880 7280 11920 7285
rect 11880 7275 11885 7280
rect 11695 7255 11885 7275
rect 11695 7250 11700 7255
rect 11660 7245 11700 7250
rect 11880 7250 11885 7255
rect 11915 7275 11920 7280
rect 12100 7280 12140 7285
rect 12100 7275 12105 7280
rect 11915 7255 12105 7275
rect 11915 7250 11920 7255
rect 11880 7245 11920 7250
rect 12100 7250 12105 7255
rect 12135 7275 12140 7280
rect 12320 7280 12360 7285
rect 12320 7275 12325 7280
rect 12135 7255 12325 7275
rect 12135 7250 12140 7255
rect 12100 7245 12140 7250
rect 12320 7250 12325 7255
rect 12355 7250 12360 7280
rect 12320 7245 12360 7250
rect 12978 7280 13012 7285
rect 12978 7250 12981 7280
rect 13009 7250 13012 7280
rect 12978 7245 13012 7250
rect 18313 7280 18347 7285
rect 18313 7250 18316 7280
rect 18344 7250 18347 7280
rect 18313 7245 18347 7250
rect 18940 7280 18980 7285
rect 18940 7250 18945 7280
rect 18975 7275 18980 7280
rect 19160 7280 19200 7285
rect 19160 7275 19165 7280
rect 18975 7255 19165 7275
rect 18975 7250 18980 7255
rect 18940 7245 18980 7250
rect 19160 7250 19165 7255
rect 19195 7275 19200 7280
rect 19380 7280 19420 7285
rect 19380 7275 19385 7280
rect 19195 7255 19385 7275
rect 19195 7250 19200 7255
rect 19160 7245 19200 7250
rect 19380 7250 19385 7255
rect 19415 7275 19420 7280
rect 19600 7280 19640 7285
rect 19600 7275 19605 7280
rect 19415 7255 19605 7275
rect 19415 7250 19420 7255
rect 19380 7245 19420 7250
rect 19600 7250 19605 7255
rect 19635 7275 19640 7280
rect 19820 7280 19860 7285
rect 19820 7275 19825 7280
rect 19635 7255 19825 7275
rect 19635 7250 19640 7255
rect 19600 7245 19640 7250
rect 19820 7250 19825 7255
rect 19855 7250 19860 7280
rect 19820 7245 19860 7250
rect 20473 7280 20507 7285
rect 20473 7250 20476 7280
rect 20504 7250 20507 7280
rect 20473 7245 20507 7250
rect 11330 7235 11370 7240
rect 9790 7220 9830 7225
rect 9790 7190 9795 7220
rect 9825 7215 9830 7220
rect 9900 7220 9940 7225
rect 9900 7215 9905 7220
rect 9825 7195 9905 7215
rect 9825 7190 9830 7195
rect 9790 7185 9830 7190
rect 9900 7190 9905 7195
rect 9935 7215 9940 7220
rect 10010 7220 10050 7225
rect 10010 7215 10015 7220
rect 9935 7195 10015 7215
rect 9935 7190 9940 7195
rect 9900 7185 9940 7190
rect 10010 7190 10015 7195
rect 10045 7215 10050 7220
rect 10120 7220 10160 7225
rect 10120 7215 10125 7220
rect 10045 7195 10125 7215
rect 10045 7190 10050 7195
rect 10010 7185 10050 7190
rect 10120 7190 10125 7195
rect 10155 7215 10160 7220
rect 10230 7220 10270 7225
rect 10230 7215 10235 7220
rect 10155 7195 10235 7215
rect 10155 7190 10160 7195
rect 10120 7185 10160 7190
rect 10230 7190 10235 7195
rect 10265 7215 10270 7220
rect 10340 7220 10380 7225
rect 10340 7215 10345 7220
rect 10265 7195 10345 7215
rect 10265 7190 10270 7195
rect 10230 7185 10270 7190
rect 10340 7190 10345 7195
rect 10375 7215 10380 7220
rect 10450 7220 10490 7225
rect 10450 7215 10455 7220
rect 10375 7195 10455 7215
rect 10375 7190 10380 7195
rect 10340 7185 10380 7190
rect 10450 7190 10455 7195
rect 10485 7215 10490 7220
rect 10560 7220 10600 7225
rect 10560 7215 10565 7220
rect 10485 7195 10565 7215
rect 10485 7190 10490 7195
rect 10450 7185 10490 7190
rect 10560 7190 10565 7195
rect 10595 7215 10600 7220
rect 10670 7220 10710 7225
rect 10670 7215 10675 7220
rect 10595 7195 10675 7215
rect 10595 7190 10600 7195
rect 10560 7185 10600 7190
rect 10670 7190 10675 7195
rect 10705 7215 10710 7220
rect 10780 7220 10820 7225
rect 10780 7215 10785 7220
rect 10705 7195 10785 7215
rect 10705 7190 10710 7195
rect 10670 7185 10710 7190
rect 10780 7190 10785 7195
rect 10815 7190 10820 7220
rect 11330 7205 11335 7235
rect 11365 7230 11370 7235
rect 11550 7235 11590 7240
rect 11550 7230 11555 7235
rect 11365 7210 11555 7230
rect 11365 7205 11370 7210
rect 11330 7200 11370 7205
rect 11550 7205 11555 7210
rect 11585 7230 11590 7235
rect 11770 7235 11810 7240
rect 11770 7230 11775 7235
rect 11585 7210 11775 7230
rect 11585 7205 11590 7210
rect 11550 7200 11590 7205
rect 11770 7205 11775 7210
rect 11805 7230 11810 7235
rect 11990 7235 12030 7240
rect 11990 7230 11995 7235
rect 11805 7210 11995 7230
rect 11805 7205 11810 7210
rect 11770 7200 11810 7205
rect 11990 7205 11995 7210
rect 12025 7230 12030 7235
rect 12210 7235 12250 7240
rect 12210 7230 12215 7235
rect 12025 7210 12215 7230
rect 12025 7205 12030 7210
rect 11990 7200 12030 7205
rect 12210 7205 12215 7210
rect 12245 7230 12250 7235
rect 12430 7235 12470 7240
rect 12430 7230 12435 7235
rect 12245 7210 12435 7230
rect 12245 7205 12250 7210
rect 12210 7200 12250 7205
rect 12430 7205 12435 7210
rect 12465 7205 12470 7235
rect 18830 7235 18870 7240
rect 12430 7200 12470 7205
rect 13005 7220 13045 7225
rect 10780 7185 10820 7190
rect 13005 7190 13010 7220
rect 13040 7215 13045 7220
rect 13115 7220 13155 7225
rect 13115 7215 13120 7220
rect 13040 7195 13120 7215
rect 13040 7190 13045 7195
rect 13005 7185 13045 7190
rect 13115 7190 13120 7195
rect 13150 7215 13155 7220
rect 13225 7220 13265 7225
rect 13225 7215 13230 7220
rect 13150 7195 13230 7215
rect 13150 7190 13155 7195
rect 13115 7185 13155 7190
rect 13225 7190 13230 7195
rect 13260 7215 13265 7220
rect 13335 7220 13375 7225
rect 13335 7215 13340 7220
rect 13260 7195 13340 7215
rect 13260 7190 13265 7195
rect 13225 7185 13265 7190
rect 13335 7190 13340 7195
rect 13370 7215 13375 7220
rect 13445 7220 13485 7225
rect 13445 7215 13450 7220
rect 13370 7195 13450 7215
rect 13370 7190 13375 7195
rect 13335 7185 13375 7190
rect 13445 7190 13450 7195
rect 13480 7215 13485 7220
rect 13555 7220 13595 7225
rect 13555 7215 13560 7220
rect 13480 7195 13560 7215
rect 13480 7190 13485 7195
rect 13445 7185 13485 7190
rect 13555 7190 13560 7195
rect 13590 7215 13595 7220
rect 13665 7220 13705 7225
rect 13665 7215 13670 7220
rect 13590 7195 13670 7215
rect 13590 7190 13595 7195
rect 13555 7185 13595 7190
rect 13665 7190 13670 7195
rect 13700 7215 13705 7220
rect 13775 7220 13815 7225
rect 13775 7215 13780 7220
rect 13700 7195 13780 7215
rect 13700 7190 13705 7195
rect 13665 7185 13705 7190
rect 13775 7190 13780 7195
rect 13810 7215 13815 7220
rect 13885 7220 13925 7225
rect 13885 7215 13890 7220
rect 13810 7195 13890 7215
rect 13810 7190 13815 7195
rect 13775 7185 13815 7190
rect 13885 7190 13890 7195
rect 13920 7215 13925 7220
rect 13995 7220 14035 7225
rect 13995 7215 14000 7220
rect 13920 7195 14000 7215
rect 13920 7190 13925 7195
rect 13885 7185 13925 7190
rect 13995 7190 14000 7195
rect 14030 7190 14035 7220
rect 13995 7185 14035 7190
rect 17290 7220 17330 7225
rect 17290 7190 17295 7220
rect 17325 7215 17330 7220
rect 17400 7220 17440 7225
rect 17400 7215 17405 7220
rect 17325 7195 17405 7215
rect 17325 7190 17330 7195
rect 17290 7185 17330 7190
rect 17400 7190 17405 7195
rect 17435 7215 17440 7220
rect 17510 7220 17550 7225
rect 17510 7215 17515 7220
rect 17435 7195 17515 7215
rect 17435 7190 17440 7195
rect 17400 7185 17440 7190
rect 17510 7190 17515 7195
rect 17545 7215 17550 7220
rect 17620 7220 17660 7225
rect 17620 7215 17625 7220
rect 17545 7195 17625 7215
rect 17545 7190 17550 7195
rect 17510 7185 17550 7190
rect 17620 7190 17625 7195
rect 17655 7215 17660 7220
rect 17730 7220 17770 7225
rect 17730 7215 17735 7220
rect 17655 7195 17735 7215
rect 17655 7190 17660 7195
rect 17620 7185 17660 7190
rect 17730 7190 17735 7195
rect 17765 7215 17770 7220
rect 17840 7220 17880 7225
rect 17840 7215 17845 7220
rect 17765 7195 17845 7215
rect 17765 7190 17770 7195
rect 17730 7185 17770 7190
rect 17840 7190 17845 7195
rect 17875 7215 17880 7220
rect 17950 7220 17990 7225
rect 17950 7215 17955 7220
rect 17875 7195 17955 7215
rect 17875 7190 17880 7195
rect 17840 7185 17880 7190
rect 17950 7190 17955 7195
rect 17985 7215 17990 7220
rect 18060 7220 18100 7225
rect 18060 7215 18065 7220
rect 17985 7195 18065 7215
rect 17985 7190 17990 7195
rect 17950 7185 17990 7190
rect 18060 7190 18065 7195
rect 18095 7215 18100 7220
rect 18170 7220 18210 7225
rect 18170 7215 18175 7220
rect 18095 7195 18175 7215
rect 18095 7190 18100 7195
rect 18060 7185 18100 7190
rect 18170 7190 18175 7195
rect 18205 7215 18210 7220
rect 18280 7220 18320 7225
rect 18280 7215 18285 7220
rect 18205 7195 18285 7215
rect 18205 7190 18210 7195
rect 18170 7185 18210 7190
rect 18280 7190 18285 7195
rect 18315 7190 18320 7220
rect 18830 7205 18835 7235
rect 18865 7230 18870 7235
rect 19050 7235 19090 7240
rect 19050 7230 19055 7235
rect 18865 7210 19055 7230
rect 18865 7205 18870 7210
rect 18830 7200 18870 7205
rect 19050 7205 19055 7210
rect 19085 7230 19090 7235
rect 19270 7235 19310 7240
rect 19270 7230 19275 7235
rect 19085 7210 19275 7230
rect 19085 7205 19090 7210
rect 19050 7200 19090 7205
rect 19270 7205 19275 7210
rect 19305 7230 19310 7235
rect 19490 7235 19530 7240
rect 19490 7230 19495 7235
rect 19305 7210 19495 7230
rect 19305 7205 19310 7210
rect 19270 7200 19310 7205
rect 19490 7205 19495 7210
rect 19525 7230 19530 7235
rect 19710 7235 19750 7240
rect 19710 7230 19715 7235
rect 19525 7210 19715 7230
rect 19525 7205 19530 7210
rect 19490 7200 19530 7205
rect 19710 7205 19715 7210
rect 19745 7230 19750 7235
rect 19930 7235 19970 7240
rect 19930 7230 19935 7235
rect 19745 7210 19935 7230
rect 19745 7205 19750 7210
rect 19710 7200 19750 7205
rect 19930 7205 19935 7210
rect 19965 7205 19970 7235
rect 19930 7200 19970 7205
rect 20500 7220 20540 7225
rect 18280 7185 18320 7190
rect 20500 7190 20505 7220
rect 20535 7215 20540 7220
rect 20610 7220 20650 7225
rect 20610 7215 20615 7220
rect 20535 7195 20615 7215
rect 20535 7190 20540 7195
rect 20500 7185 20540 7190
rect 20610 7190 20615 7195
rect 20645 7215 20650 7220
rect 20720 7220 20760 7225
rect 20720 7215 20725 7220
rect 20645 7195 20725 7215
rect 20645 7190 20650 7195
rect 20610 7185 20650 7190
rect 20720 7190 20725 7195
rect 20755 7215 20760 7220
rect 20830 7220 20870 7225
rect 20830 7215 20835 7220
rect 20755 7195 20835 7215
rect 20755 7190 20760 7195
rect 20720 7185 20760 7190
rect 20830 7190 20835 7195
rect 20865 7215 20870 7220
rect 20940 7220 20980 7225
rect 20940 7215 20945 7220
rect 20865 7195 20945 7215
rect 20865 7190 20870 7195
rect 20830 7185 20870 7190
rect 20940 7190 20945 7195
rect 20975 7215 20980 7220
rect 21050 7220 21090 7225
rect 21050 7215 21055 7220
rect 20975 7195 21055 7215
rect 20975 7190 20980 7195
rect 20940 7185 20980 7190
rect 21050 7190 21055 7195
rect 21085 7215 21090 7220
rect 21160 7220 21200 7225
rect 21160 7215 21165 7220
rect 21085 7195 21165 7215
rect 21085 7190 21090 7195
rect 21050 7185 21090 7190
rect 21160 7190 21165 7195
rect 21195 7215 21200 7220
rect 21270 7220 21310 7225
rect 21270 7215 21275 7220
rect 21195 7195 21275 7215
rect 21195 7190 21200 7195
rect 21160 7185 21200 7190
rect 21270 7190 21275 7195
rect 21305 7215 21310 7220
rect 21380 7220 21420 7225
rect 21380 7215 21385 7220
rect 21305 7195 21385 7215
rect 21305 7190 21310 7195
rect 21270 7185 21310 7190
rect 21380 7190 21385 7195
rect 21415 7215 21420 7220
rect 21490 7220 21530 7225
rect 21490 7215 21495 7220
rect 21415 7195 21495 7215
rect 21415 7190 21420 7195
rect 21380 7185 21420 7190
rect 21490 7190 21495 7195
rect 21525 7190 21530 7220
rect 21490 7185 21530 7190
rect 9735 7000 9775 7005
rect 9735 6970 9740 7000
rect 9770 6995 9775 7000
rect 9845 7000 9885 7005
rect 9845 6995 9850 7000
rect 9770 6975 9850 6995
rect 9770 6970 9775 6975
rect 9735 6965 9775 6970
rect 9845 6970 9850 6975
rect 9880 6995 9885 7000
rect 9955 7000 9995 7005
rect 9955 6995 9960 7000
rect 9880 6975 9960 6995
rect 9880 6970 9885 6975
rect 9845 6965 9885 6970
rect 9955 6970 9960 6975
rect 9990 6995 9995 7000
rect 10065 7000 10105 7005
rect 10065 6995 10070 7000
rect 9990 6975 10070 6995
rect 9990 6970 9995 6975
rect 9955 6965 9995 6970
rect 10065 6970 10070 6975
rect 10100 6995 10105 7000
rect 10175 7000 10215 7005
rect 10175 6995 10180 7000
rect 10100 6975 10180 6995
rect 10100 6970 10105 6975
rect 10065 6965 10105 6970
rect 10175 6970 10180 6975
rect 10210 6995 10215 7000
rect 10285 7000 10325 7005
rect 10285 6995 10290 7000
rect 10210 6975 10290 6995
rect 10210 6970 10215 6975
rect 10175 6965 10215 6970
rect 10285 6970 10290 6975
rect 10320 6995 10325 7000
rect 10395 7000 10435 7005
rect 10395 6995 10400 7000
rect 10320 6975 10400 6995
rect 10320 6970 10325 6975
rect 10285 6965 10325 6970
rect 10395 6970 10400 6975
rect 10430 6995 10435 7000
rect 10505 7000 10545 7005
rect 10505 6995 10510 7000
rect 10430 6975 10510 6995
rect 10430 6970 10435 6975
rect 10395 6965 10435 6970
rect 10505 6970 10510 6975
rect 10540 6995 10545 7000
rect 10615 7000 10655 7005
rect 10615 6995 10620 7000
rect 10540 6975 10620 6995
rect 10540 6970 10545 6975
rect 10505 6965 10545 6970
rect 10615 6970 10620 6975
rect 10650 6995 10655 7000
rect 10725 7000 10765 7005
rect 10725 6995 10730 7000
rect 10650 6975 10730 6995
rect 10650 6970 10655 6975
rect 10615 6965 10655 6970
rect 10725 6970 10730 6975
rect 10760 6995 10765 7000
rect 10835 7000 10875 7005
rect 10835 6995 10840 7000
rect 10760 6975 10840 6995
rect 10760 6970 10765 6975
rect 10725 6965 10765 6970
rect 10835 6970 10840 6975
rect 10870 6970 10875 7000
rect 10835 6965 10875 6970
rect 12950 7000 12990 7005
rect 12950 6970 12955 7000
rect 12985 6995 12990 7000
rect 13060 7000 13100 7005
rect 13060 6995 13065 7000
rect 12985 6975 13065 6995
rect 12985 6970 12990 6975
rect 12950 6965 12990 6970
rect 13060 6970 13065 6975
rect 13095 6995 13100 7000
rect 13170 7000 13210 7005
rect 13170 6995 13175 7000
rect 13095 6975 13175 6995
rect 13095 6970 13100 6975
rect 13060 6965 13100 6970
rect 13170 6970 13175 6975
rect 13205 6995 13210 7000
rect 13280 7000 13320 7005
rect 13280 6995 13285 7000
rect 13205 6975 13285 6995
rect 13205 6970 13210 6975
rect 13170 6965 13210 6970
rect 13280 6970 13285 6975
rect 13315 6995 13320 7000
rect 13390 7000 13430 7005
rect 13390 6995 13395 7000
rect 13315 6975 13395 6995
rect 13315 6970 13320 6975
rect 13280 6965 13320 6970
rect 13390 6970 13395 6975
rect 13425 6995 13430 7000
rect 13500 7000 13540 7005
rect 13500 6995 13505 7000
rect 13425 6975 13505 6995
rect 13425 6970 13430 6975
rect 13390 6965 13430 6970
rect 13500 6970 13505 6975
rect 13535 6995 13540 7000
rect 13610 7000 13650 7005
rect 13610 6995 13615 7000
rect 13535 6975 13615 6995
rect 13535 6970 13540 6975
rect 13500 6965 13540 6970
rect 13610 6970 13615 6975
rect 13645 6995 13650 7000
rect 13720 7000 13760 7005
rect 13720 6995 13725 7000
rect 13645 6975 13725 6995
rect 13645 6970 13650 6975
rect 13610 6965 13650 6970
rect 13720 6970 13725 6975
rect 13755 6995 13760 7000
rect 13830 7000 13870 7005
rect 13830 6995 13835 7000
rect 13755 6975 13835 6995
rect 13755 6970 13760 6975
rect 13720 6965 13760 6970
rect 13830 6970 13835 6975
rect 13865 6995 13870 7000
rect 13940 7000 13980 7005
rect 13940 6995 13945 7000
rect 13865 6975 13945 6995
rect 13865 6970 13870 6975
rect 13830 6965 13870 6970
rect 13940 6970 13945 6975
rect 13975 6995 13980 7000
rect 14050 7000 14090 7005
rect 14050 6995 14055 7000
rect 13975 6975 14055 6995
rect 13975 6970 13980 6975
rect 13940 6965 13980 6970
rect 14050 6970 14055 6975
rect 14085 6970 14090 7000
rect 14050 6965 14090 6970
rect 17235 7000 17275 7005
rect 17235 6970 17240 7000
rect 17270 6995 17275 7000
rect 17345 7000 17385 7005
rect 17345 6995 17350 7000
rect 17270 6975 17350 6995
rect 17270 6970 17275 6975
rect 17235 6965 17275 6970
rect 17345 6970 17350 6975
rect 17380 6995 17385 7000
rect 17455 7000 17495 7005
rect 17455 6995 17460 7000
rect 17380 6975 17460 6995
rect 17380 6970 17385 6975
rect 17345 6965 17385 6970
rect 17455 6970 17460 6975
rect 17490 6995 17495 7000
rect 17565 7000 17605 7005
rect 17565 6995 17570 7000
rect 17490 6975 17570 6995
rect 17490 6970 17495 6975
rect 17455 6965 17495 6970
rect 17565 6970 17570 6975
rect 17600 6995 17605 7000
rect 17675 7000 17715 7005
rect 17675 6995 17680 7000
rect 17600 6975 17680 6995
rect 17600 6970 17605 6975
rect 17565 6965 17605 6970
rect 17675 6970 17680 6975
rect 17710 6995 17715 7000
rect 17785 7000 17825 7005
rect 17785 6995 17790 7000
rect 17710 6975 17790 6995
rect 17710 6970 17715 6975
rect 17675 6965 17715 6970
rect 17785 6970 17790 6975
rect 17820 6995 17825 7000
rect 17895 7000 17935 7005
rect 17895 6995 17900 7000
rect 17820 6975 17900 6995
rect 17820 6970 17825 6975
rect 17785 6965 17825 6970
rect 17895 6970 17900 6975
rect 17930 6995 17935 7000
rect 18005 7000 18045 7005
rect 18005 6995 18010 7000
rect 17930 6975 18010 6995
rect 17930 6970 17935 6975
rect 17895 6965 17935 6970
rect 18005 6970 18010 6975
rect 18040 6995 18045 7000
rect 18115 7000 18155 7005
rect 18115 6995 18120 7000
rect 18040 6975 18120 6995
rect 18040 6970 18045 6975
rect 18005 6965 18045 6970
rect 18115 6970 18120 6975
rect 18150 6995 18155 7000
rect 18225 7000 18265 7005
rect 18225 6995 18230 7000
rect 18150 6975 18230 6995
rect 18150 6970 18155 6975
rect 18115 6965 18155 6970
rect 18225 6970 18230 6975
rect 18260 6995 18265 7000
rect 18335 7000 18375 7005
rect 18335 6995 18340 7000
rect 18260 6975 18340 6995
rect 18260 6970 18265 6975
rect 18225 6965 18265 6970
rect 18335 6970 18340 6975
rect 18370 6970 18375 7000
rect 18335 6965 18375 6970
rect 20445 7000 20485 7005
rect 20445 6970 20450 7000
rect 20480 6995 20485 7000
rect 20555 7000 20595 7005
rect 20555 6995 20560 7000
rect 20480 6975 20560 6995
rect 20480 6970 20485 6975
rect 20445 6965 20485 6970
rect 20555 6970 20560 6975
rect 20590 6995 20595 7000
rect 20665 7000 20705 7005
rect 20665 6995 20670 7000
rect 20590 6975 20670 6995
rect 20590 6970 20595 6975
rect 20555 6965 20595 6970
rect 20665 6970 20670 6975
rect 20700 6995 20705 7000
rect 20775 7000 20815 7005
rect 20775 6995 20780 7000
rect 20700 6975 20780 6995
rect 20700 6970 20705 6975
rect 20665 6965 20705 6970
rect 20775 6970 20780 6975
rect 20810 6995 20815 7000
rect 20885 7000 20925 7005
rect 20885 6995 20890 7000
rect 20810 6975 20890 6995
rect 20810 6970 20815 6975
rect 20775 6965 20815 6970
rect 20885 6970 20890 6975
rect 20920 6995 20925 7000
rect 20995 7000 21035 7005
rect 20995 6995 21000 7000
rect 20920 6975 21000 6995
rect 20920 6970 20925 6975
rect 20885 6965 20925 6970
rect 20995 6970 21000 6975
rect 21030 6995 21035 7000
rect 21105 7000 21145 7005
rect 21105 6995 21110 7000
rect 21030 6975 21110 6995
rect 21030 6970 21035 6975
rect 20995 6965 21035 6970
rect 21105 6970 21110 6975
rect 21140 6995 21145 7000
rect 21215 7000 21255 7005
rect 21215 6995 21220 7000
rect 21140 6975 21220 6995
rect 21140 6970 21145 6975
rect 21105 6965 21145 6970
rect 21215 6970 21220 6975
rect 21250 6995 21255 7000
rect 21325 7000 21365 7005
rect 21325 6995 21330 7000
rect 21250 6975 21330 6995
rect 21250 6970 21255 6975
rect 21215 6965 21255 6970
rect 21325 6970 21330 6975
rect 21360 6995 21365 7000
rect 21435 7000 21475 7005
rect 21435 6995 21440 7000
rect 21360 6975 21440 6995
rect 21360 6970 21365 6975
rect 21325 6965 21365 6970
rect 21435 6970 21440 6975
rect 21470 6995 21475 7000
rect 21545 7000 21585 7005
rect 21545 6995 21550 7000
rect 21470 6975 21550 6995
rect 21470 6970 21475 6975
rect 21435 6965 21475 6970
rect 21545 6970 21550 6975
rect 21580 6970 21585 7000
rect 21545 6965 21585 6970
rect 11385 6960 11425 6965
rect 11385 6930 11390 6960
rect 11420 6955 11425 6960
rect 11605 6960 11645 6965
rect 11605 6955 11610 6960
rect 11420 6935 11610 6955
rect 11420 6930 11425 6935
rect 11385 6925 11425 6930
rect 11605 6930 11610 6935
rect 11640 6955 11645 6960
rect 11825 6960 11865 6965
rect 11825 6955 11830 6960
rect 11640 6935 11830 6955
rect 11640 6930 11645 6935
rect 11605 6925 11645 6930
rect 11825 6930 11830 6935
rect 11860 6955 11865 6960
rect 12045 6960 12085 6965
rect 12045 6955 12050 6960
rect 11860 6935 12050 6955
rect 11860 6930 11865 6935
rect 11825 6925 11865 6930
rect 12045 6930 12050 6935
rect 12080 6955 12085 6960
rect 12265 6960 12305 6965
rect 12265 6955 12270 6960
rect 12080 6935 12270 6955
rect 12080 6930 12085 6935
rect 12045 6925 12085 6930
rect 12265 6930 12270 6935
rect 12300 6930 12305 6960
rect 12265 6925 12305 6930
rect 18885 6960 18925 6965
rect 18885 6930 18890 6960
rect 18920 6955 18925 6960
rect 19105 6960 19145 6965
rect 19105 6955 19110 6960
rect 18920 6935 19110 6955
rect 18920 6930 18925 6935
rect 18885 6925 18925 6930
rect 19105 6930 19110 6935
rect 19140 6955 19145 6960
rect 19325 6960 19365 6965
rect 19325 6955 19330 6960
rect 19140 6935 19330 6955
rect 19140 6930 19145 6935
rect 19105 6925 19145 6930
rect 19325 6930 19330 6935
rect 19360 6955 19365 6960
rect 19545 6960 19585 6965
rect 19545 6955 19550 6960
rect 19360 6935 19550 6955
rect 19360 6930 19365 6935
rect 19325 6925 19365 6930
rect 19545 6930 19550 6935
rect 19580 6955 19585 6960
rect 19765 6960 19805 6965
rect 19765 6955 19770 6960
rect 19580 6935 19770 6955
rect 19580 6930 19585 6935
rect 19545 6925 19585 6930
rect 19765 6930 19770 6935
rect 19800 6930 19805 6960
rect 19765 6925 19805 6930
rect 11495 6905 11535 6910
rect 11495 6875 11500 6905
rect 11530 6900 11535 6905
rect 11715 6905 11755 6910
rect 11715 6900 11720 6905
rect 11530 6880 11720 6900
rect 11530 6875 11535 6880
rect 11495 6870 11535 6875
rect 11715 6875 11720 6880
rect 11750 6900 11755 6905
rect 11935 6905 11975 6910
rect 11935 6900 11940 6905
rect 11750 6880 11940 6900
rect 11750 6875 11755 6880
rect 11715 6870 11755 6875
rect 11935 6875 11940 6880
rect 11970 6900 11975 6905
rect 12155 6905 12195 6910
rect 12155 6900 12160 6905
rect 11970 6880 12160 6900
rect 11970 6875 11975 6880
rect 11935 6870 11975 6875
rect 12155 6875 12160 6880
rect 12190 6900 12195 6905
rect 12375 6905 12415 6910
rect 12375 6900 12380 6905
rect 12190 6880 12380 6900
rect 12190 6875 12195 6880
rect 12155 6870 12195 6875
rect 12375 6875 12380 6880
rect 12410 6875 12415 6905
rect 12375 6870 12415 6875
rect 18995 6905 19035 6910
rect 18995 6875 19000 6905
rect 19030 6900 19035 6905
rect 19215 6905 19255 6910
rect 19215 6900 19220 6905
rect 19030 6880 19220 6900
rect 19030 6875 19035 6880
rect 18995 6870 19035 6875
rect 19215 6875 19220 6880
rect 19250 6900 19255 6905
rect 19435 6905 19475 6910
rect 19435 6900 19440 6905
rect 19250 6880 19440 6900
rect 19250 6875 19255 6880
rect 19215 6870 19255 6875
rect 19435 6875 19440 6880
rect 19470 6900 19475 6905
rect 19655 6905 19695 6910
rect 19655 6900 19660 6905
rect 19470 6880 19660 6900
rect 19470 6875 19475 6880
rect 19435 6870 19475 6875
rect 19655 6875 19660 6880
rect 19690 6900 19695 6905
rect 19875 6905 19915 6910
rect 19875 6900 19880 6905
rect 19690 6880 19880 6900
rect 19690 6875 19695 6880
rect 19655 6870 19695 6875
rect 19875 6875 19880 6880
rect 19910 6875 19915 6905
rect 19875 6870 19915 6875
rect 20545 6905 20585 6910
rect 20545 6875 20550 6905
rect 20580 6900 20585 6905
rect 20655 6905 20695 6910
rect 20655 6900 20660 6905
rect 20580 6880 20660 6900
rect 20580 6875 20585 6880
rect 20545 6870 20585 6875
rect 20655 6875 20660 6880
rect 20690 6900 20695 6905
rect 20765 6905 20805 6910
rect 20765 6900 20770 6905
rect 20690 6880 20770 6900
rect 20690 6875 20695 6880
rect 20655 6870 20695 6875
rect 20765 6875 20770 6880
rect 20800 6875 20805 6905
rect 20765 6870 20805 6875
rect 11190 6850 11230 6855
rect 11190 6820 11195 6850
rect 11225 6845 11230 6850
rect 11410 6850 11450 6855
rect 11410 6845 11415 6850
rect 11225 6825 11415 6845
rect 11225 6820 11230 6825
rect 11190 6815 11230 6820
rect 11410 6820 11415 6825
rect 11445 6845 11450 6850
rect 11640 6850 11680 6855
rect 11640 6845 11645 6850
rect 11445 6825 11645 6845
rect 11445 6820 11450 6825
rect 11410 6815 11450 6820
rect 11640 6820 11645 6825
rect 11675 6845 11680 6850
rect 12230 6850 12270 6855
rect 12230 6845 12235 6850
rect 11675 6825 12235 6845
rect 11675 6820 11680 6825
rect 11640 6815 11680 6820
rect 12230 6820 12235 6825
rect 12265 6845 12270 6850
rect 12450 6850 12490 6855
rect 12450 6845 12455 6850
rect 12265 6825 12455 6845
rect 12265 6820 12270 6825
rect 12230 6815 12270 6820
rect 12450 6820 12455 6825
rect 12485 6845 12490 6850
rect 12680 6850 12720 6855
rect 12680 6845 12685 6850
rect 12485 6825 12685 6845
rect 12485 6820 12490 6825
rect 12450 6815 12490 6820
rect 12680 6820 12685 6825
rect 12715 6820 12720 6850
rect 12680 6815 12720 6820
rect 18690 6850 18730 6855
rect 18690 6820 18695 6850
rect 18725 6845 18730 6850
rect 18910 6850 18950 6855
rect 18910 6845 18915 6850
rect 18725 6825 18915 6845
rect 18725 6820 18730 6825
rect 18690 6815 18730 6820
rect 18910 6820 18915 6825
rect 18945 6845 18950 6850
rect 19140 6850 19180 6855
rect 19140 6845 19145 6850
rect 18945 6825 19145 6845
rect 18945 6820 18950 6825
rect 18910 6815 18950 6820
rect 19140 6820 19145 6825
rect 19175 6845 19180 6850
rect 19730 6850 19770 6855
rect 19730 6845 19735 6850
rect 19175 6825 19735 6845
rect 19175 6820 19180 6825
rect 19140 6815 19180 6820
rect 19730 6820 19735 6825
rect 19765 6845 19770 6850
rect 19950 6850 19990 6855
rect 19950 6845 19955 6850
rect 19765 6825 19955 6845
rect 19765 6820 19770 6825
rect 19730 6815 19770 6820
rect 19950 6820 19955 6825
rect 19985 6845 19990 6850
rect 20180 6850 20220 6855
rect 20180 6845 20185 6850
rect 19985 6825 20185 6845
rect 19985 6820 19990 6825
rect 19950 6815 19990 6820
rect 20180 6820 20185 6825
rect 20215 6820 20220 6850
rect 20180 6815 20220 6820
rect 11820 6805 11860 6810
rect 11820 6775 11825 6805
rect 11855 6800 11860 6805
rect 11940 6805 11980 6810
rect 11940 6800 11945 6805
rect 11855 6780 11945 6800
rect 11855 6775 11860 6780
rect 11820 6770 11860 6775
rect 11940 6775 11945 6780
rect 11975 6775 11980 6805
rect 11940 6770 11980 6775
rect 19320 6805 19360 6810
rect 19320 6775 19325 6805
rect 19355 6800 19360 6805
rect 19440 6805 19480 6810
rect 19440 6800 19445 6805
rect 19355 6780 19445 6800
rect 19355 6775 19360 6780
rect 19320 6770 19360 6775
rect 19440 6775 19445 6780
rect 19475 6775 19480 6805
rect 19440 6770 19480 6775
rect 11085 6760 11125 6765
rect 11085 6730 11090 6760
rect 11120 6755 11125 6760
rect 11305 6760 11345 6765
rect 11305 6755 11310 6760
rect 11120 6735 11310 6755
rect 11120 6730 11125 6735
rect 11085 6725 11125 6730
rect 11305 6730 11310 6735
rect 11340 6755 11345 6760
rect 11525 6760 11565 6765
rect 11525 6755 11530 6760
rect 11340 6735 11530 6755
rect 11340 6730 11345 6735
rect 11305 6725 11345 6730
rect 11525 6730 11530 6735
rect 11560 6755 11565 6760
rect 12125 6760 12165 6765
rect 12125 6755 12130 6760
rect 11560 6735 12130 6755
rect 11560 6730 11565 6735
rect 11525 6725 11565 6730
rect 12125 6730 12130 6735
rect 12160 6755 12165 6760
rect 12345 6760 12385 6765
rect 12345 6755 12350 6760
rect 12160 6735 12350 6755
rect 12160 6730 12165 6735
rect 12125 6725 12165 6730
rect 12345 6730 12350 6735
rect 12380 6755 12385 6760
rect 12565 6760 12605 6765
rect 12565 6755 12570 6760
rect 12380 6735 12570 6755
rect 12380 6730 12385 6735
rect 12345 6725 12385 6730
rect 12565 6730 12570 6735
rect 12600 6730 12605 6760
rect 12565 6725 12605 6730
rect 18585 6760 18625 6765
rect 18585 6730 18590 6760
rect 18620 6755 18625 6760
rect 18805 6760 18845 6765
rect 18805 6755 18810 6760
rect 18620 6735 18810 6755
rect 18620 6730 18625 6735
rect 18585 6725 18625 6730
rect 18805 6730 18810 6735
rect 18840 6755 18845 6760
rect 19025 6760 19065 6765
rect 19025 6755 19030 6760
rect 18840 6735 19030 6755
rect 18840 6730 18845 6735
rect 18805 6725 18845 6730
rect 19025 6730 19030 6735
rect 19060 6755 19065 6760
rect 19625 6760 19665 6765
rect 19625 6755 19630 6760
rect 19060 6735 19630 6755
rect 19060 6730 19065 6735
rect 19025 6725 19065 6730
rect 19625 6730 19630 6735
rect 19660 6755 19665 6760
rect 19845 6760 19885 6765
rect 19845 6755 19850 6760
rect 19660 6735 19850 6755
rect 19660 6730 19665 6735
rect 19625 6725 19665 6730
rect 19845 6730 19850 6735
rect 19880 6755 19885 6760
rect 20065 6760 20105 6765
rect 20065 6755 20070 6760
rect 19880 6735 20070 6755
rect 19880 6730 19885 6735
rect 19845 6725 19885 6730
rect 20065 6730 20070 6735
rect 20100 6730 20105 6760
rect 20065 6725 20105 6730
rect 11237 6715 11269 6720
rect 11237 6710 11240 6715
rect 10910 6690 11240 6710
rect 11237 6685 11240 6690
rect 11266 6710 11269 6715
rect 11457 6715 11489 6720
rect 11457 6710 11460 6715
rect 11266 6690 11460 6710
rect 11266 6685 11269 6690
rect 11237 6680 11269 6685
rect 11457 6685 11460 6690
rect 11486 6710 11489 6715
rect 11601 6715 11633 6720
rect 11601 6710 11604 6715
rect 11486 6690 11604 6710
rect 11486 6685 11489 6690
rect 11457 6680 11489 6685
rect 11601 6685 11604 6690
rect 11630 6710 11633 6715
rect 11867 6715 11899 6720
rect 11867 6710 11870 6715
rect 11630 6690 11870 6710
rect 11630 6685 11633 6690
rect 11601 6680 11633 6685
rect 11867 6685 11870 6690
rect 11896 6710 11899 6715
rect 12277 6715 12309 6720
rect 12277 6710 12280 6715
rect 11896 6690 12280 6710
rect 11896 6685 11899 6690
rect 11867 6680 11899 6685
rect 12277 6685 12280 6690
rect 12306 6710 12309 6715
rect 12497 6715 12529 6720
rect 12497 6710 12500 6715
rect 12306 6690 12500 6710
rect 12306 6685 12309 6690
rect 12277 6680 12309 6685
rect 12497 6685 12500 6690
rect 12526 6710 12529 6715
rect 12641 6715 12673 6720
rect 12641 6710 12644 6715
rect 12526 6690 12644 6710
rect 12526 6685 12529 6690
rect 12497 6680 12529 6685
rect 12641 6685 12644 6690
rect 12670 6685 12673 6715
rect 18737 6715 18769 6720
rect 18737 6710 18740 6715
rect 18410 6690 18740 6710
rect 12641 6680 12673 6685
rect 18737 6685 18740 6690
rect 18766 6710 18769 6715
rect 18957 6715 18989 6720
rect 18957 6710 18960 6715
rect 18766 6690 18960 6710
rect 18766 6685 18769 6690
rect 18737 6680 18769 6685
rect 18957 6685 18960 6690
rect 18986 6710 18989 6715
rect 19101 6715 19133 6720
rect 19101 6710 19104 6715
rect 18986 6690 19104 6710
rect 18986 6685 18989 6690
rect 18957 6680 18989 6685
rect 19101 6685 19104 6690
rect 19130 6710 19133 6715
rect 19367 6715 19399 6720
rect 19367 6710 19370 6715
rect 19130 6690 19370 6710
rect 19130 6685 19133 6690
rect 19101 6680 19133 6685
rect 19367 6685 19370 6690
rect 19396 6710 19399 6715
rect 19777 6715 19809 6720
rect 19777 6710 19780 6715
rect 19396 6690 19780 6710
rect 19396 6685 19399 6690
rect 19367 6680 19399 6685
rect 19777 6685 19780 6690
rect 19806 6710 19809 6715
rect 19997 6715 20029 6720
rect 19997 6710 20000 6715
rect 19806 6690 20000 6710
rect 19806 6685 19809 6690
rect 19777 6680 19809 6685
rect 19997 6685 20000 6690
rect 20026 6710 20029 6715
rect 20141 6715 20173 6720
rect 20141 6710 20144 6715
rect 20026 6690 20144 6710
rect 20026 6685 20029 6690
rect 19997 6680 20029 6685
rect 20141 6685 20144 6690
rect 20170 6685 20173 6715
rect 20141 6680 20173 6685
rect 20566 6680 20598 6685
rect 20566 6650 20570 6680
rect 20596 6650 20598 6680
rect 20566 6645 20598 6650
rect 20510 6630 20550 6635
rect 20510 6600 20515 6630
rect 20545 6625 20550 6630
rect 20616 6630 20656 6635
rect 20616 6625 20621 6630
rect 20545 6605 20621 6625
rect 20545 6600 20550 6605
rect 20510 6595 20550 6600
rect 20616 6600 20621 6605
rect 20651 6600 20656 6630
rect 20616 6595 20656 6600
rect 20710 6630 20750 6635
rect 20710 6600 20715 6630
rect 20745 6625 20750 6630
rect 20800 6630 20840 6635
rect 20800 6625 20805 6630
rect 20745 6605 20805 6625
rect 20745 6600 20750 6605
rect 20710 6595 20750 6600
rect 20800 6600 20805 6605
rect 20835 6600 20840 6630
rect 20800 6595 20840 6600
rect 12815 6570 12855 6575
rect 12815 6540 12820 6570
rect 12850 6540 12855 6570
rect 12815 6535 12855 6540
rect 20315 6570 20355 6575
rect 20315 6540 20320 6570
rect 20350 6565 20355 6570
rect 20471 6570 20503 6575
rect 20471 6565 20475 6570
rect 20350 6545 20475 6565
rect 20350 6540 20355 6545
rect 20315 6535 20355 6540
rect 20471 6540 20475 6545
rect 20501 6565 20503 6570
rect 20847 6570 20879 6575
rect 20847 6565 20849 6570
rect 20501 6545 20849 6565
rect 20501 6540 20503 6545
rect 20471 6535 20503 6540
rect 20847 6540 20849 6545
rect 20875 6540 20879 6570
rect 20847 6535 20879 6540
rect 11106 6495 11138 6500
rect 11106 6490 11109 6495
rect 10910 6470 11109 6490
rect 11106 6465 11109 6470
rect 11135 6490 11138 6495
rect 11305 6495 11345 6500
rect 11305 6490 11310 6495
rect 11135 6470 11310 6490
rect 11135 6465 11138 6470
rect 11106 6460 11138 6465
rect 11305 6465 11310 6470
rect 11340 6490 11345 6495
rect 11525 6495 11565 6500
rect 11525 6490 11530 6495
rect 11340 6470 11530 6490
rect 11340 6465 11345 6470
rect 11305 6460 11345 6465
rect 11525 6465 11530 6470
rect 11560 6490 11565 6495
rect 11922 6495 11954 6500
rect 11922 6490 11925 6495
rect 11560 6470 11925 6490
rect 11560 6465 11565 6470
rect 11525 6460 11565 6465
rect 11922 6465 11925 6470
rect 11951 6490 11954 6495
rect 12146 6495 12178 6500
rect 12146 6490 12149 6495
rect 11951 6470 12149 6490
rect 11951 6465 11954 6470
rect 11922 6460 11954 6465
rect 12146 6465 12149 6470
rect 12175 6490 12178 6495
rect 12345 6495 12385 6500
rect 12345 6490 12350 6495
rect 12175 6470 12350 6490
rect 12175 6465 12178 6470
rect 12146 6460 12178 6465
rect 12345 6465 12350 6470
rect 12380 6490 12385 6495
rect 12565 6495 12605 6500
rect 12565 6490 12570 6495
rect 12380 6470 12570 6490
rect 12380 6465 12385 6470
rect 12345 6460 12385 6465
rect 12565 6465 12570 6470
rect 12600 6465 12605 6495
rect 18606 6495 18638 6500
rect 18606 6490 18609 6495
rect 18410 6470 18609 6490
rect 12565 6460 12605 6465
rect 18606 6465 18609 6470
rect 18635 6490 18638 6495
rect 18805 6495 18845 6500
rect 18805 6490 18810 6495
rect 18635 6470 18810 6490
rect 18635 6465 18638 6470
rect 18606 6460 18638 6465
rect 18805 6465 18810 6470
rect 18840 6490 18845 6495
rect 19025 6495 19065 6500
rect 19025 6490 19030 6495
rect 18840 6470 19030 6490
rect 18840 6465 18845 6470
rect 18805 6460 18845 6465
rect 19025 6465 19030 6470
rect 19060 6490 19065 6495
rect 19422 6495 19454 6500
rect 19422 6490 19425 6495
rect 19060 6470 19425 6490
rect 19060 6465 19065 6470
rect 19025 6460 19065 6465
rect 19422 6465 19425 6470
rect 19451 6490 19454 6495
rect 19646 6495 19678 6500
rect 19646 6490 19649 6495
rect 19451 6470 19649 6490
rect 19451 6465 19454 6470
rect 19422 6460 19454 6465
rect 19646 6465 19649 6470
rect 19675 6490 19678 6495
rect 19845 6495 19885 6500
rect 19845 6490 19850 6495
rect 19675 6470 19850 6490
rect 19675 6465 19678 6470
rect 19646 6460 19678 6465
rect 19845 6465 19850 6470
rect 19880 6490 19885 6495
rect 20065 6495 20105 6500
rect 20065 6490 20070 6495
rect 19880 6470 20070 6490
rect 19880 6465 19885 6470
rect 19845 6460 19885 6465
rect 20065 6465 20070 6470
rect 20100 6465 20105 6495
rect 20065 6460 20105 6465
rect 9760 6410 9765 6445
rect 9800 6410 9805 6445
rect 10770 6410 10775 6445
rect 10810 6410 10815 6445
rect 11145 6435 11185 6440
rect 11145 6405 11150 6435
rect 11180 6430 11185 6435
rect 11250 6435 11290 6440
rect 11250 6430 11255 6435
rect 11180 6410 11255 6430
rect 11180 6405 11185 6410
rect 11145 6400 11185 6405
rect 11250 6405 11255 6410
rect 11285 6430 11290 6435
rect 11360 6435 11400 6440
rect 11360 6430 11365 6435
rect 11285 6410 11365 6430
rect 11285 6405 11290 6410
rect 11250 6400 11290 6405
rect 11360 6405 11365 6410
rect 11395 6430 11400 6435
rect 11470 6435 11510 6440
rect 11470 6430 11475 6435
rect 11395 6410 11475 6430
rect 11395 6405 11400 6410
rect 11360 6400 11400 6405
rect 11470 6405 11475 6410
rect 11505 6430 11510 6435
rect 11580 6435 11620 6440
rect 11580 6430 11585 6435
rect 11505 6410 11585 6430
rect 11505 6405 11510 6410
rect 11470 6400 11510 6405
rect 11580 6405 11585 6410
rect 11615 6430 11620 6435
rect 12185 6435 12225 6440
rect 12185 6430 12190 6435
rect 11615 6410 12190 6430
rect 11615 6405 11620 6410
rect 11580 6400 11620 6405
rect 12185 6405 12190 6410
rect 12220 6430 12225 6435
rect 12290 6435 12330 6440
rect 12290 6430 12295 6435
rect 12220 6410 12295 6430
rect 12220 6405 12225 6410
rect 12185 6400 12225 6405
rect 12290 6405 12295 6410
rect 12325 6430 12330 6435
rect 12400 6435 12440 6440
rect 12400 6430 12405 6435
rect 12325 6410 12405 6430
rect 12325 6405 12330 6410
rect 12290 6400 12330 6405
rect 12400 6405 12405 6410
rect 12435 6430 12440 6435
rect 12510 6435 12550 6440
rect 12510 6430 12515 6435
rect 12435 6410 12515 6430
rect 12435 6405 12440 6410
rect 12400 6400 12440 6405
rect 12510 6405 12515 6410
rect 12545 6430 12550 6435
rect 12620 6435 12660 6440
rect 12620 6430 12625 6435
rect 12545 6410 12625 6430
rect 12545 6405 12550 6410
rect 12510 6400 12550 6405
rect 12620 6405 12625 6410
rect 12655 6405 12660 6435
rect 12985 6410 12990 6445
rect 13025 6410 13030 6445
rect 13995 6410 14000 6445
rect 14035 6410 14040 6445
rect 18645 6435 18685 6440
rect 12620 6400 12660 6405
rect 18645 6405 18650 6435
rect 18680 6430 18685 6435
rect 18750 6435 18790 6440
rect 18750 6430 18755 6435
rect 18680 6410 18755 6430
rect 18680 6405 18685 6410
rect 18645 6400 18685 6405
rect 18750 6405 18755 6410
rect 18785 6430 18790 6435
rect 18860 6435 18900 6440
rect 18860 6430 18865 6435
rect 18785 6410 18865 6430
rect 18785 6405 18790 6410
rect 18750 6400 18790 6405
rect 18860 6405 18865 6410
rect 18895 6430 18900 6435
rect 18970 6435 19010 6440
rect 18970 6430 18975 6435
rect 18895 6410 18975 6430
rect 18895 6405 18900 6410
rect 18860 6400 18900 6405
rect 18970 6405 18975 6410
rect 19005 6430 19010 6435
rect 19080 6435 19120 6440
rect 19080 6430 19085 6435
rect 19005 6410 19085 6430
rect 19005 6405 19010 6410
rect 18970 6400 19010 6405
rect 19080 6405 19085 6410
rect 19115 6430 19120 6435
rect 19685 6435 19725 6440
rect 19685 6430 19690 6435
rect 19115 6410 19690 6430
rect 19115 6405 19120 6410
rect 19080 6400 19120 6405
rect 19685 6405 19690 6410
rect 19720 6430 19725 6435
rect 19790 6435 19830 6440
rect 19790 6430 19795 6435
rect 19720 6410 19795 6430
rect 19720 6405 19725 6410
rect 19685 6400 19725 6405
rect 19790 6405 19795 6410
rect 19825 6430 19830 6435
rect 19900 6435 19940 6440
rect 19900 6430 19905 6435
rect 19825 6410 19905 6430
rect 19825 6405 19830 6410
rect 19790 6400 19830 6405
rect 19900 6405 19905 6410
rect 19935 6430 19940 6435
rect 20010 6435 20050 6440
rect 20010 6430 20015 6435
rect 19935 6410 20015 6430
rect 19935 6405 19940 6410
rect 19900 6400 19940 6405
rect 20010 6405 20015 6410
rect 20045 6430 20050 6435
rect 20120 6435 20160 6440
rect 20120 6430 20125 6435
rect 20045 6410 20125 6430
rect 20045 6405 20050 6410
rect 20010 6400 20050 6405
rect 20120 6405 20125 6410
rect 20155 6405 20160 6435
rect 20120 6400 20160 6405
rect 10665 6390 10705 6395
rect 10665 6360 10670 6390
rect 10700 6385 10705 6390
rect 10770 6390 10810 6395
rect 10770 6385 10775 6390
rect 10700 6365 10775 6385
rect 10700 6360 10705 6365
rect 10665 6355 10705 6360
rect 10770 6360 10775 6365
rect 10805 6385 10810 6390
rect 12990 6390 13030 6395
rect 12990 6385 12995 6390
rect 10805 6365 12995 6385
rect 10805 6360 10810 6365
rect 10770 6355 10810 6360
rect 12990 6360 12995 6365
rect 13025 6385 13030 6390
rect 13095 6390 13135 6395
rect 13095 6385 13100 6390
rect 13025 6365 13100 6385
rect 13025 6360 13030 6365
rect 12990 6355 13030 6360
rect 13095 6360 13100 6365
rect 13130 6360 13135 6390
rect 13095 6355 13135 6360
rect 19310 6385 19350 6390
rect 19310 6355 19315 6385
rect 19345 6355 19350 6385
rect 19310 6350 19350 6355
rect 20526 6350 20558 6355
rect 11810 6345 11850 6350
rect 20526 6345 20528 6350
rect 9765 6335 9805 6340
rect 9765 6305 9770 6335
rect 9800 6330 9805 6335
rect 9965 6335 10005 6340
rect 9965 6330 9970 6335
rect 9800 6310 9970 6330
rect 9800 6305 9805 6310
rect 9765 6300 9805 6305
rect 9965 6305 9970 6310
rect 10000 6330 10005 6335
rect 10165 6335 10205 6340
rect 10165 6330 10170 6335
rect 10000 6310 10170 6330
rect 10000 6305 10005 6310
rect 9965 6300 10005 6305
rect 10165 6305 10170 6310
rect 10200 6330 10205 6335
rect 10365 6335 10405 6340
rect 10365 6330 10370 6335
rect 10200 6310 10370 6330
rect 10200 6305 10205 6310
rect 10165 6300 10205 6305
rect 10365 6305 10370 6310
rect 10400 6330 10405 6335
rect 10565 6335 10605 6340
rect 10565 6330 10570 6335
rect 10400 6310 10570 6330
rect 10400 6305 10405 6310
rect 10365 6300 10405 6305
rect 10565 6305 10570 6310
rect 10600 6330 10605 6335
rect 10765 6335 10805 6340
rect 10765 6330 10770 6335
rect 10600 6310 10770 6330
rect 10600 6305 10605 6310
rect 10565 6300 10605 6305
rect 10765 6305 10770 6310
rect 10800 6305 10805 6335
rect 11810 6315 11815 6345
rect 11845 6315 11850 6345
rect 11810 6310 11850 6315
rect 12995 6335 13035 6340
rect 10765 6300 10805 6305
rect 12995 6305 13000 6335
rect 13030 6330 13035 6335
rect 13195 6335 13235 6340
rect 13195 6330 13200 6335
rect 13030 6310 13200 6330
rect 13030 6305 13035 6310
rect 12995 6300 13035 6305
rect 13195 6305 13200 6310
rect 13230 6330 13235 6335
rect 13395 6335 13435 6340
rect 13395 6330 13400 6335
rect 13230 6310 13400 6330
rect 13230 6305 13235 6310
rect 13195 6300 13235 6305
rect 13395 6305 13400 6310
rect 13430 6330 13435 6335
rect 13595 6335 13635 6340
rect 13595 6330 13600 6335
rect 13430 6310 13600 6330
rect 13430 6305 13435 6310
rect 13395 6300 13435 6305
rect 13595 6305 13600 6310
rect 13630 6330 13635 6335
rect 13795 6335 13835 6340
rect 13795 6330 13800 6335
rect 13630 6310 13800 6330
rect 13630 6305 13635 6310
rect 13595 6300 13635 6305
rect 13795 6305 13800 6310
rect 13830 6330 13835 6335
rect 13995 6335 14035 6340
rect 13995 6330 14000 6335
rect 13830 6310 14000 6330
rect 13830 6305 13835 6310
rect 13795 6300 13835 6305
rect 13995 6305 14000 6310
rect 14030 6305 14035 6335
rect 13995 6300 14035 6305
rect 18815 6335 18855 6340
rect 18815 6305 18820 6335
rect 18850 6330 18855 6335
rect 19380 6335 19420 6340
rect 19380 6330 19385 6335
rect 18850 6310 19385 6330
rect 18850 6305 18855 6310
rect 18815 6300 18855 6305
rect 19380 6305 19385 6310
rect 19415 6305 19420 6335
rect 20525 6325 20528 6345
rect 20526 6320 20528 6325
rect 20554 6345 20558 6350
rect 20792 6350 20824 6355
rect 20792 6345 20796 6350
rect 20554 6325 20796 6345
rect 20554 6320 20558 6325
rect 20526 6315 20558 6320
rect 20792 6320 20796 6325
rect 20822 6345 20824 6350
rect 20822 6325 20825 6345
rect 20822 6320 20824 6325
rect 20792 6315 20824 6320
rect 19380 6300 19420 6305
rect 11315 6295 11355 6300
rect 11315 6265 11320 6295
rect 11350 6290 11355 6295
rect 11880 6295 11920 6300
rect 11880 6290 11885 6295
rect 11350 6270 11885 6290
rect 11350 6265 11355 6270
rect 11315 6260 11355 6265
rect 11880 6265 11885 6270
rect 11915 6265 11920 6295
rect 20095 6290 20135 6295
rect 11880 6260 11920 6265
rect 18925 6275 18965 6280
rect 12595 6250 12635 6255
rect 11425 6235 11465 6240
rect 11425 6205 11430 6235
rect 11460 6230 11465 6235
rect 11535 6235 11575 6240
rect 11535 6230 11540 6235
rect 11460 6210 11540 6230
rect 11460 6205 11465 6210
rect 11425 6200 11465 6205
rect 11535 6205 11540 6210
rect 11570 6230 11575 6235
rect 11645 6235 11685 6240
rect 11645 6230 11650 6235
rect 11570 6210 11650 6230
rect 11570 6205 11575 6210
rect 11535 6200 11575 6205
rect 11645 6205 11650 6210
rect 11680 6230 11685 6235
rect 11755 6235 11795 6240
rect 11755 6230 11760 6235
rect 11680 6210 11760 6230
rect 11680 6205 11685 6210
rect 11645 6200 11685 6205
rect 11755 6205 11760 6210
rect 11790 6230 11795 6235
rect 11865 6235 11905 6240
rect 11865 6230 11870 6235
rect 11790 6210 11870 6230
rect 11790 6205 11795 6210
rect 11755 6200 11795 6205
rect 11865 6205 11870 6210
rect 11900 6230 11905 6235
rect 11975 6235 12015 6240
rect 11975 6230 11980 6235
rect 11900 6210 11980 6230
rect 11900 6205 11905 6210
rect 11865 6200 11905 6205
rect 11975 6205 11980 6210
rect 12010 6230 12015 6235
rect 12085 6235 12125 6240
rect 12085 6230 12090 6235
rect 12010 6210 12090 6230
rect 12010 6205 12015 6210
rect 11975 6200 12015 6205
rect 12085 6205 12090 6210
rect 12120 6230 12125 6235
rect 12195 6235 12235 6240
rect 12195 6230 12200 6235
rect 12120 6210 12200 6230
rect 12120 6205 12125 6210
rect 12085 6200 12125 6205
rect 12195 6205 12200 6210
rect 12230 6230 12235 6235
rect 12305 6235 12345 6240
rect 12305 6230 12310 6235
rect 12230 6210 12310 6230
rect 12230 6205 12235 6210
rect 12195 6200 12235 6205
rect 12305 6205 12310 6210
rect 12340 6230 12345 6235
rect 12415 6235 12455 6240
rect 12415 6230 12420 6235
rect 12340 6210 12420 6230
rect 12340 6205 12345 6210
rect 12305 6200 12345 6205
rect 12415 6205 12420 6210
rect 12450 6230 12455 6235
rect 12525 6235 12565 6240
rect 12525 6230 12530 6235
rect 12450 6210 12530 6230
rect 12450 6205 12455 6210
rect 12415 6200 12455 6205
rect 12525 6205 12530 6210
rect 12560 6205 12565 6235
rect 12595 6220 12600 6250
rect 12630 6245 12635 6250
rect 18925 6245 18930 6275
rect 18960 6270 18965 6275
rect 19035 6275 19075 6280
rect 19035 6270 19040 6275
rect 18960 6250 19040 6270
rect 18960 6245 18965 6250
rect 12630 6225 12695 6245
rect 18925 6240 18965 6245
rect 19035 6245 19040 6250
rect 19070 6270 19075 6275
rect 19145 6275 19185 6280
rect 19145 6270 19150 6275
rect 19070 6250 19150 6270
rect 19070 6245 19075 6250
rect 19035 6240 19075 6245
rect 19145 6245 19150 6250
rect 19180 6270 19185 6275
rect 19255 6275 19295 6280
rect 19255 6270 19260 6275
rect 19180 6250 19260 6270
rect 19180 6245 19185 6250
rect 19145 6240 19185 6245
rect 19255 6245 19260 6250
rect 19290 6270 19295 6275
rect 19365 6275 19405 6280
rect 19365 6270 19370 6275
rect 19290 6250 19370 6270
rect 19290 6245 19295 6250
rect 19255 6240 19295 6245
rect 19365 6245 19370 6250
rect 19400 6270 19405 6275
rect 19475 6275 19515 6280
rect 19475 6270 19480 6275
rect 19400 6250 19480 6270
rect 19400 6245 19405 6250
rect 19365 6240 19405 6245
rect 19475 6245 19480 6250
rect 19510 6270 19515 6275
rect 19585 6275 19625 6280
rect 19585 6270 19590 6275
rect 19510 6250 19590 6270
rect 19510 6245 19515 6250
rect 19475 6240 19515 6245
rect 19585 6245 19590 6250
rect 19620 6270 19625 6275
rect 19695 6275 19735 6280
rect 19695 6270 19700 6275
rect 19620 6250 19700 6270
rect 19620 6245 19625 6250
rect 19585 6240 19625 6245
rect 19695 6245 19700 6250
rect 19730 6270 19735 6275
rect 19805 6275 19845 6280
rect 19805 6270 19810 6275
rect 19730 6250 19810 6270
rect 19730 6245 19735 6250
rect 19695 6240 19735 6245
rect 19805 6245 19810 6250
rect 19840 6270 19845 6275
rect 19915 6275 19955 6280
rect 19915 6270 19920 6275
rect 19840 6250 19920 6270
rect 19840 6245 19845 6250
rect 19805 6240 19845 6245
rect 19915 6245 19920 6250
rect 19950 6270 19955 6275
rect 20025 6275 20065 6280
rect 20025 6270 20030 6275
rect 19950 6250 20030 6270
rect 19950 6245 19955 6250
rect 19915 6240 19955 6245
rect 20025 6245 20030 6250
rect 20060 6245 20065 6275
rect 20095 6260 20100 6290
rect 20130 6285 20135 6290
rect 20445 6290 20485 6295
rect 20445 6285 20450 6290
rect 20130 6265 20450 6285
rect 20130 6260 20135 6265
rect 20095 6255 20135 6260
rect 20445 6260 20450 6265
rect 20480 6285 20485 6290
rect 20560 6290 20600 6295
rect 20560 6285 20565 6290
rect 20480 6265 20565 6285
rect 20480 6260 20485 6265
rect 20445 6255 20485 6260
rect 20560 6260 20565 6265
rect 20595 6260 20600 6290
rect 20560 6255 20600 6260
rect 20655 6290 20695 6295
rect 20655 6260 20660 6290
rect 20690 6285 20695 6290
rect 20750 6290 20790 6295
rect 20750 6285 20755 6290
rect 20690 6265 20755 6285
rect 20690 6260 20695 6265
rect 20655 6255 20695 6260
rect 20750 6260 20755 6265
rect 20785 6260 20790 6290
rect 20750 6255 20790 6260
rect 20865 6290 20905 6295
rect 20865 6260 20870 6290
rect 20900 6260 20905 6290
rect 20865 6255 20905 6260
rect 20025 6240 20065 6245
rect 20600 6230 20640 6235
rect 12630 6220 12635 6225
rect 12595 6215 12635 6220
rect 12525 6200 12565 6205
rect 20600 6200 20605 6230
rect 20635 6225 20640 6230
rect 20660 6230 20690 6235
rect 20635 6205 20660 6225
rect 20635 6200 20640 6205
rect 20600 6195 20640 6200
rect 20660 6195 20690 6200
rect 20710 6230 20750 6235
rect 20710 6200 20715 6230
rect 20745 6225 20750 6230
rect 20865 6230 20905 6235
rect 20865 6225 20870 6230
rect 20745 6205 20870 6225
rect 20745 6200 20750 6205
rect 20710 6195 20750 6200
rect 20865 6200 20870 6205
rect 20900 6200 20905 6230
rect 20865 6195 20905 6200
rect 9865 5985 9905 5990
rect 9865 5955 9870 5985
rect 9900 5980 9905 5985
rect 10065 5985 10105 5990
rect 10065 5980 10070 5985
rect 9900 5960 10070 5980
rect 9900 5955 9905 5960
rect 9865 5950 9905 5955
rect 10065 5955 10070 5960
rect 10100 5980 10105 5985
rect 10265 5985 10305 5990
rect 10265 5980 10270 5985
rect 10100 5960 10270 5980
rect 10100 5955 10105 5960
rect 10065 5950 10105 5955
rect 10265 5955 10270 5960
rect 10300 5980 10305 5985
rect 10465 5985 10505 5990
rect 10465 5980 10470 5985
rect 10300 5960 10470 5980
rect 10300 5955 10305 5960
rect 10265 5950 10305 5955
rect 10465 5955 10470 5960
rect 10500 5980 10505 5985
rect 10665 5985 10705 5990
rect 10665 5980 10670 5985
rect 10500 5960 10670 5980
rect 10500 5955 10505 5960
rect 10465 5950 10505 5955
rect 10665 5955 10670 5960
rect 10700 5955 10705 5985
rect 10665 5950 10705 5955
rect 13095 5985 13135 5990
rect 13095 5955 13100 5985
rect 13130 5980 13135 5985
rect 13295 5985 13335 5990
rect 13295 5980 13300 5985
rect 13130 5960 13300 5980
rect 13130 5955 13135 5960
rect 13095 5950 13135 5955
rect 13295 5955 13300 5960
rect 13330 5980 13335 5985
rect 13495 5985 13535 5990
rect 13495 5980 13500 5985
rect 13330 5960 13500 5980
rect 13330 5955 13335 5960
rect 13295 5950 13335 5955
rect 13495 5955 13500 5960
rect 13530 5980 13535 5985
rect 13695 5985 13735 5990
rect 13695 5980 13700 5985
rect 13530 5960 13700 5980
rect 13530 5955 13535 5960
rect 13495 5950 13535 5955
rect 13695 5955 13700 5960
rect 13730 5980 13735 5985
rect 13895 5985 13935 5990
rect 13895 5980 13900 5985
rect 13730 5960 13900 5980
rect 13730 5955 13735 5960
rect 13695 5950 13735 5955
rect 13895 5955 13900 5960
rect 13930 5955 13935 5985
rect 13895 5950 13935 5955
rect 18665 5955 18705 5960
rect 18665 5925 18670 5955
rect 18700 5950 18705 5955
rect 18760 5955 18800 5960
rect 18760 5950 18765 5955
rect 18700 5930 18765 5950
rect 18700 5925 18705 5930
rect 18665 5920 18705 5925
rect 18760 5925 18765 5930
rect 18795 5950 18800 5955
rect 18870 5955 18910 5960
rect 18870 5950 18875 5955
rect 18795 5930 18875 5950
rect 18795 5925 18800 5930
rect 18760 5920 18800 5925
rect 18870 5925 18875 5930
rect 18905 5950 18910 5955
rect 18980 5955 19020 5960
rect 18980 5950 18985 5955
rect 18905 5930 18985 5950
rect 18905 5925 18910 5930
rect 18870 5920 18910 5925
rect 18980 5925 18985 5930
rect 19015 5950 19020 5955
rect 19090 5955 19130 5960
rect 19090 5950 19095 5955
rect 19015 5930 19095 5950
rect 19015 5925 19020 5930
rect 18980 5920 19020 5925
rect 19090 5925 19095 5930
rect 19125 5950 19130 5955
rect 19200 5955 19240 5960
rect 19200 5950 19205 5955
rect 19125 5930 19205 5950
rect 19125 5925 19130 5930
rect 19090 5920 19130 5925
rect 19200 5925 19205 5930
rect 19235 5950 19240 5955
rect 19310 5955 19350 5960
rect 19310 5950 19315 5955
rect 19235 5930 19315 5950
rect 19235 5925 19240 5930
rect 19200 5920 19240 5925
rect 19310 5925 19315 5930
rect 19345 5950 19350 5955
rect 19420 5955 19460 5960
rect 19420 5950 19425 5955
rect 19345 5930 19425 5950
rect 19345 5925 19350 5930
rect 19310 5920 19350 5925
rect 19420 5925 19425 5930
rect 19455 5950 19460 5955
rect 19530 5955 19570 5960
rect 19530 5950 19535 5955
rect 19455 5930 19535 5950
rect 19455 5925 19460 5930
rect 19420 5920 19460 5925
rect 19530 5925 19535 5930
rect 19565 5950 19570 5955
rect 19640 5955 19680 5960
rect 19640 5950 19645 5955
rect 19565 5930 19645 5950
rect 19565 5925 19570 5930
rect 19530 5920 19570 5925
rect 19640 5925 19645 5930
rect 19675 5950 19680 5955
rect 19750 5955 19790 5960
rect 19750 5950 19755 5955
rect 19675 5930 19755 5950
rect 19675 5925 19680 5930
rect 19640 5920 19680 5925
rect 19750 5925 19755 5930
rect 19785 5950 19790 5955
rect 19860 5955 19900 5960
rect 19860 5950 19865 5955
rect 19785 5930 19865 5950
rect 19785 5925 19790 5930
rect 19750 5920 19790 5925
rect 19860 5925 19865 5930
rect 19895 5950 19900 5955
rect 19970 5955 20010 5960
rect 19970 5950 19975 5955
rect 19895 5930 19975 5950
rect 19895 5925 19900 5930
rect 19860 5920 19900 5925
rect 19970 5925 19975 5930
rect 20005 5950 20010 5955
rect 20120 5955 20160 5960
rect 20120 5950 20125 5955
rect 20005 5930 20125 5950
rect 20005 5925 20010 5930
rect 19970 5920 20010 5925
rect 20120 5925 20125 5930
rect 20155 5925 20160 5955
rect 20120 5920 20160 5925
rect 11165 5915 11205 5920
rect 11165 5885 11170 5915
rect 11200 5910 11205 5915
rect 11260 5915 11300 5920
rect 11260 5910 11265 5915
rect 11200 5890 11265 5910
rect 11200 5885 11205 5890
rect 11165 5880 11205 5885
rect 11260 5885 11265 5890
rect 11295 5910 11300 5915
rect 11370 5915 11410 5920
rect 11370 5910 11375 5915
rect 11295 5890 11375 5910
rect 11295 5885 11300 5890
rect 11260 5880 11300 5885
rect 11370 5885 11375 5890
rect 11405 5910 11410 5915
rect 11480 5915 11520 5920
rect 11480 5910 11485 5915
rect 11405 5890 11485 5910
rect 11405 5885 11410 5890
rect 11370 5880 11410 5885
rect 11480 5885 11485 5890
rect 11515 5910 11520 5915
rect 11590 5915 11630 5920
rect 11590 5910 11595 5915
rect 11515 5890 11595 5910
rect 11515 5885 11520 5890
rect 11480 5880 11520 5885
rect 11590 5885 11595 5890
rect 11625 5910 11630 5915
rect 11700 5915 11740 5920
rect 11700 5910 11705 5915
rect 11625 5890 11705 5910
rect 11625 5885 11630 5890
rect 11590 5880 11630 5885
rect 11700 5885 11705 5890
rect 11735 5910 11740 5915
rect 11810 5915 11850 5920
rect 11810 5910 11815 5915
rect 11735 5890 11815 5910
rect 11735 5885 11740 5890
rect 11700 5880 11740 5885
rect 11810 5885 11815 5890
rect 11845 5910 11850 5915
rect 11920 5915 11960 5920
rect 11920 5910 11925 5915
rect 11845 5890 11925 5910
rect 11845 5885 11850 5890
rect 11810 5880 11850 5885
rect 11920 5885 11925 5890
rect 11955 5910 11960 5915
rect 12030 5915 12070 5920
rect 12030 5910 12035 5915
rect 11955 5890 12035 5910
rect 11955 5885 11960 5890
rect 11920 5880 11960 5885
rect 12030 5885 12035 5890
rect 12065 5910 12070 5915
rect 12140 5915 12180 5920
rect 12140 5910 12145 5915
rect 12065 5890 12145 5910
rect 12065 5885 12070 5890
rect 12030 5880 12070 5885
rect 12140 5885 12145 5890
rect 12175 5910 12180 5915
rect 12250 5915 12290 5920
rect 12250 5910 12255 5915
rect 12175 5890 12255 5910
rect 12175 5885 12180 5890
rect 12140 5880 12180 5885
rect 12250 5885 12255 5890
rect 12285 5910 12290 5915
rect 12360 5915 12400 5920
rect 12360 5910 12365 5915
rect 12285 5890 12365 5910
rect 12285 5885 12290 5890
rect 12250 5880 12290 5885
rect 12360 5885 12365 5890
rect 12395 5910 12400 5915
rect 12470 5915 12510 5920
rect 12470 5910 12475 5915
rect 12395 5890 12475 5910
rect 12395 5885 12400 5890
rect 12360 5880 12400 5885
rect 12470 5885 12475 5890
rect 12505 5910 12510 5915
rect 12620 5915 12660 5920
rect 12620 5910 12625 5915
rect 12505 5890 12625 5910
rect 12505 5885 12510 5890
rect 12470 5880 12510 5885
rect 12620 5885 12625 5890
rect 12655 5885 12660 5915
rect 12620 5880 12660 5885
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect 11632 4515 11668 4520
rect 11632 4485 11635 4515
rect 11665 4510 11668 4515
rect 11752 4515 11788 4520
rect 11752 4510 11755 4515
rect 11665 4490 11755 4510
rect 11665 4485 11668 4490
rect 11632 4480 11668 4485
rect 11752 4485 11755 4490
rect 11785 4510 11788 4515
rect 11872 4515 11908 4520
rect 11872 4510 11875 4515
rect 11785 4490 11875 4510
rect 11785 4485 11788 4490
rect 11752 4480 11788 4485
rect 11872 4485 11875 4490
rect 11905 4510 11908 4515
rect 12080 4515 12120 4520
rect 12080 4510 12085 4515
rect 11905 4490 12085 4510
rect 11905 4485 11908 4490
rect 11872 4480 11908 4485
rect 12080 4485 12085 4490
rect 12115 4485 12120 4515
rect 12080 4480 12120 4485
rect 11570 4470 11610 4475
rect 11570 4460 11575 4470
rect 11200 4455 11240 4460
rect 11200 4425 11205 4455
rect 11235 4425 11240 4455
rect 11200 4420 11240 4425
rect 11460 4455 11575 4460
rect 11460 4425 11465 4455
rect 11495 4440 11575 4455
rect 11605 4465 11610 4470
rect 11690 4470 11730 4475
rect 11690 4465 11695 4470
rect 11605 4445 11695 4465
rect 11605 4440 11610 4445
rect 11495 4425 11500 4440
rect 11570 4435 11610 4440
rect 11690 4440 11695 4445
rect 11725 4465 11730 4470
rect 11810 4470 11850 4475
rect 11810 4465 11815 4470
rect 11725 4445 11815 4465
rect 11725 4440 11730 4445
rect 11690 4435 11730 4440
rect 11810 4440 11815 4445
rect 11845 4465 11850 4470
rect 11930 4470 11970 4475
rect 11930 4465 11935 4470
rect 11845 4445 11935 4465
rect 11845 4440 11850 4445
rect 11810 4435 11850 4440
rect 11930 4440 11935 4445
rect 11965 4440 11970 4470
rect 11930 4435 11970 4440
rect 12080 4445 12120 4450
rect 11460 4420 11500 4425
rect 12080 4415 12085 4445
rect 12115 4440 12120 4445
rect 12200 4445 12240 4450
rect 12200 4440 12205 4445
rect 12115 4420 12205 4440
rect 12115 4415 12120 4420
rect 12080 4410 12120 4415
rect 12200 4415 12205 4420
rect 12235 4440 12240 4445
rect 12320 4445 12360 4450
rect 12320 4440 12325 4445
rect 12235 4420 12325 4440
rect 12235 4415 12240 4420
rect 12200 4410 12240 4415
rect 12320 4415 12325 4420
rect 12355 4440 12360 4445
rect 12440 4445 12480 4450
rect 12440 4440 12445 4445
rect 12355 4420 12445 4440
rect 12355 4415 12360 4420
rect 12320 4410 12360 4415
rect 12440 4415 12445 4420
rect 12475 4440 12480 4445
rect 12560 4445 12600 4450
rect 12560 4440 12565 4445
rect 12475 4420 12565 4440
rect 12475 4415 12480 4420
rect 12440 4410 12480 4415
rect 12560 4415 12565 4420
rect 12595 4415 12600 4445
rect 12560 4410 12600 4415
rect 11330 4320 11370 4325
rect 11050 4315 11090 4320
rect 11050 4285 11055 4315
rect 11085 4310 11090 4315
rect 11330 4310 11335 4320
rect 11085 4290 11335 4310
rect 11365 4310 11370 4320
rect 11750 4315 11790 4320
rect 11750 4310 11755 4315
rect 11365 4290 11755 4310
rect 11085 4285 11090 4290
rect 11330 4285 11370 4290
rect 11750 4285 11755 4290
rect 11785 4310 11790 4315
rect 12140 4315 12180 4320
rect 12140 4310 12145 4315
rect 11785 4290 12145 4310
rect 11785 4285 11790 4290
rect 11050 4280 11090 4285
rect 11750 4280 11790 4285
rect 12140 4285 12145 4290
rect 12175 4310 12180 4315
rect 12260 4315 12300 4320
rect 12260 4310 12265 4315
rect 12175 4290 12265 4310
rect 12175 4285 12180 4290
rect 12140 4280 12180 4285
rect 12260 4285 12265 4290
rect 12295 4310 12300 4315
rect 12380 4315 12420 4320
rect 12380 4310 12385 4315
rect 12295 4290 12385 4310
rect 12295 4285 12300 4290
rect 12260 4280 12300 4285
rect 12380 4285 12385 4290
rect 12415 4310 12420 4315
rect 12500 4315 12540 4320
rect 12500 4310 12505 4315
rect 12415 4290 12505 4310
rect 12415 4285 12420 4290
rect 12380 4280 12420 4285
rect 12500 4285 12505 4290
rect 12535 4285 12540 4315
rect 12500 4280 12540 4285
rect 11105 4260 11145 4265
rect 11105 4230 11110 4260
rect 11140 4255 11145 4260
rect 11330 4260 11370 4265
rect 11330 4255 11335 4260
rect 11140 4235 11335 4255
rect 11140 4230 11145 4235
rect 11105 4225 11145 4230
rect 11330 4230 11335 4235
rect 11365 4255 11370 4260
rect 12200 4260 12240 4265
rect 12200 4255 12205 4260
rect 11365 4235 12205 4255
rect 11365 4230 11370 4235
rect 11330 4225 11370 4230
rect 12200 4230 12205 4235
rect 12235 4230 12240 4260
rect 12200 4225 12240 4230
rect 11360 4205 11400 4210
rect 11360 4175 11365 4205
rect 11395 4200 11400 4205
rect 11470 4205 11510 4210
rect 11470 4200 11475 4205
rect 11395 4180 11475 4200
rect 11395 4175 11400 4180
rect 11360 4170 11400 4175
rect 11470 4175 11475 4180
rect 11505 4200 11510 4205
rect 11580 4205 11620 4210
rect 11580 4200 11585 4205
rect 11505 4180 11585 4200
rect 11505 4175 11510 4180
rect 11470 4170 11510 4175
rect 11580 4175 11585 4180
rect 11615 4200 11620 4205
rect 11690 4205 11730 4210
rect 11690 4200 11695 4205
rect 11615 4180 11695 4200
rect 11615 4175 11620 4180
rect 11580 4170 11620 4175
rect 11690 4175 11695 4180
rect 11725 4200 11730 4205
rect 11800 4205 11840 4210
rect 11800 4200 11805 4205
rect 11725 4180 11805 4200
rect 11725 4175 11730 4180
rect 11690 4170 11730 4175
rect 11800 4175 11805 4180
rect 11835 4200 11840 4205
rect 11910 4205 11950 4210
rect 11910 4200 11915 4205
rect 11835 4180 11915 4200
rect 11835 4175 11840 4180
rect 11800 4170 11840 4175
rect 11910 4175 11915 4180
rect 11945 4200 11950 4205
rect 12020 4205 12060 4210
rect 12020 4200 12025 4205
rect 11945 4180 12025 4200
rect 11945 4175 11950 4180
rect 11910 4170 11950 4175
rect 12020 4175 12025 4180
rect 12055 4200 12060 4205
rect 12130 4205 12170 4210
rect 12130 4200 12135 4205
rect 12055 4180 12135 4200
rect 12055 4175 12060 4180
rect 12020 4170 12060 4175
rect 12130 4175 12135 4180
rect 12165 4200 12170 4205
rect 12240 4205 12280 4210
rect 12240 4200 12245 4205
rect 12165 4180 12245 4200
rect 12165 4175 12170 4180
rect 12130 4170 12170 4175
rect 12240 4175 12245 4180
rect 12275 4200 12280 4205
rect 12350 4205 12390 4210
rect 12350 4200 12355 4205
rect 12275 4180 12355 4200
rect 12275 4175 12280 4180
rect 12240 4170 12280 4175
rect 12350 4175 12355 4180
rect 12385 4175 12390 4205
rect 12350 4170 12390 4175
rect 11305 4085 11345 4090
rect 11305 4055 11310 4085
rect 11340 4080 11345 4085
rect 11525 4085 11565 4090
rect 11525 4080 11530 4085
rect 11340 4060 11530 4080
rect 11340 4055 11345 4060
rect 11305 4050 11345 4055
rect 11525 4055 11530 4060
rect 11560 4080 11565 4085
rect 11745 4085 11785 4090
rect 11745 4080 11750 4085
rect 11560 4060 11750 4080
rect 11560 4055 11565 4060
rect 11525 4050 11565 4055
rect 11745 4055 11750 4060
rect 11780 4080 11785 4085
rect 11965 4085 12005 4090
rect 11965 4080 11970 4085
rect 11780 4060 11970 4080
rect 11780 4055 11785 4060
rect 11745 4050 11785 4055
rect 11965 4055 11970 4060
rect 12000 4080 12005 4085
rect 12185 4085 12225 4090
rect 12185 4080 12190 4085
rect 12000 4060 12190 4080
rect 12000 4055 12005 4060
rect 11965 4050 12005 4055
rect 12185 4055 12190 4060
rect 12220 4080 12225 4085
rect 12405 4085 12445 4090
rect 12405 4080 12410 4085
rect 12220 4060 12410 4080
rect 12220 4055 12225 4060
rect 12185 4050 12225 4055
rect 12405 4055 12410 4060
rect 12440 4055 12445 4085
rect 12405 4050 12445 4055
rect 11415 4025 11455 4030
rect 11415 3995 11420 4025
rect 11450 4020 11455 4025
rect 11635 4025 11675 4030
rect 11635 4020 11640 4025
rect 11450 4000 11640 4020
rect 11450 3995 11455 4000
rect 11415 3990 11455 3995
rect 11635 3995 11640 4000
rect 11670 4020 11675 4025
rect 11855 4025 11895 4030
rect 11855 4020 11860 4025
rect 11670 4000 11860 4020
rect 11670 3995 11675 4000
rect 11635 3990 11675 3995
rect 11855 3995 11860 4000
rect 11890 4020 11895 4025
rect 12075 4025 12115 4030
rect 12075 4020 12080 4025
rect 11890 4000 12080 4020
rect 11890 3995 11895 4000
rect 11855 3990 11895 3995
rect 12075 3995 12080 4000
rect 12110 4020 12115 4025
rect 12295 4025 12335 4030
rect 12295 4020 12300 4025
rect 12110 4000 12300 4020
rect 12110 3995 12115 4000
rect 12075 3990 12115 3995
rect 12295 3995 12300 4000
rect 12330 3995 12335 4025
rect 12295 3990 12335 3995
rect 11310 3960 11350 3965
rect 11310 3930 11315 3960
rect 11345 3955 11350 3960
rect 11415 3960 11455 3965
rect 11415 3955 11420 3960
rect 11345 3935 11420 3955
rect 11345 3930 11350 3935
rect 11310 3925 11350 3930
rect 11415 3930 11420 3935
rect 11450 3955 11455 3960
rect 11525 3960 11565 3965
rect 11525 3955 11530 3960
rect 11450 3935 11530 3955
rect 11450 3930 11455 3935
rect 11415 3925 11455 3930
rect 11525 3930 11530 3935
rect 11560 3955 11565 3960
rect 11635 3960 11675 3965
rect 11635 3955 11640 3960
rect 11560 3935 11640 3955
rect 11560 3930 11565 3935
rect 11525 3925 11565 3930
rect 11635 3930 11640 3935
rect 11670 3955 11675 3960
rect 11745 3960 11785 3965
rect 11745 3955 11750 3960
rect 11670 3935 11750 3955
rect 11670 3930 11675 3935
rect 11635 3925 11675 3930
rect 11745 3930 11750 3935
rect 11780 3930 11785 3960
rect 11745 3925 11785 3930
rect 12050 3960 12090 3965
rect 12050 3930 12055 3960
rect 12085 3955 12090 3960
rect 12155 3960 12195 3965
rect 12155 3955 12160 3960
rect 12085 3935 12160 3955
rect 12085 3930 12090 3935
rect 12050 3925 12090 3930
rect 12155 3930 12160 3935
rect 12190 3955 12195 3960
rect 12265 3960 12305 3965
rect 12265 3955 12270 3960
rect 12190 3935 12270 3955
rect 12190 3930 12195 3935
rect 12155 3925 12195 3930
rect 12265 3930 12270 3935
rect 12300 3955 12305 3960
rect 12375 3960 12415 3965
rect 12375 3955 12380 3960
rect 12300 3935 12380 3955
rect 12300 3930 12305 3935
rect 12265 3925 12305 3930
rect 12375 3930 12380 3935
rect 12410 3955 12415 3960
rect 12485 3960 12525 3965
rect 12485 3955 12490 3960
rect 12410 3935 12490 3955
rect 12410 3930 12415 3935
rect 12375 3925 12415 3930
rect 12485 3930 12490 3935
rect 12520 3930 12525 3960
rect 12485 3925 12525 3930
rect 11271 3900 11303 3905
rect 11271 3870 11274 3900
rect 11300 3895 11303 3900
rect 11470 3900 11510 3905
rect 11470 3895 11475 3900
rect 11300 3875 11475 3895
rect 11300 3870 11303 3875
rect 11271 3865 11303 3870
rect 11470 3870 11475 3875
rect 11505 3895 11510 3900
rect 11690 3900 11730 3905
rect 11690 3895 11695 3900
rect 11505 3875 11695 3895
rect 11505 3870 11510 3875
rect 11470 3865 11510 3870
rect 11690 3870 11695 3875
rect 11725 3895 11730 3900
rect 12011 3900 12043 3905
rect 12011 3895 12014 3900
rect 11725 3875 12014 3895
rect 11725 3870 11730 3875
rect 11690 3865 11730 3870
rect 12011 3870 12014 3875
rect 12040 3895 12043 3900
rect 12210 3900 12250 3905
rect 12210 3895 12215 3900
rect 12040 3875 12215 3895
rect 12040 3870 12043 3875
rect 12011 3865 12043 3870
rect 12210 3870 12215 3875
rect 12245 3895 12250 3900
rect 12430 3900 12470 3905
rect 12430 3895 12435 3900
rect 12245 3875 12435 3895
rect 12245 3870 12250 3875
rect 12210 3865 12250 3870
rect 12430 3870 12435 3875
rect 12465 3895 12470 3900
rect 12760 3900 12800 3905
rect 12760 3895 12765 3900
rect 12465 3875 12765 3895
rect 12465 3870 12470 3875
rect 12430 3865 12470 3870
rect 12760 3870 12765 3875
rect 12795 3870 12800 3900
rect 12760 3865 12800 3870
rect 11402 3780 11434 3785
rect 11402 3775 11405 3780
rect 10625 3755 11405 3775
rect 11402 3750 11405 3755
rect 11431 3775 11434 3780
rect 11622 3780 11654 3785
rect 11622 3775 11625 3780
rect 11431 3755 11625 3775
rect 11431 3750 11434 3755
rect 11402 3745 11434 3750
rect 11622 3750 11625 3755
rect 11651 3775 11654 3780
rect 11766 3780 11798 3785
rect 11766 3775 11769 3780
rect 11651 3755 11769 3775
rect 11651 3750 11654 3755
rect 11622 3745 11654 3750
rect 11766 3750 11769 3755
rect 11795 3775 11798 3780
rect 12142 3780 12174 3785
rect 12142 3775 12145 3780
rect 11795 3755 12145 3775
rect 11795 3750 11798 3755
rect 11766 3745 11798 3750
rect 12142 3750 12145 3755
rect 12171 3775 12174 3780
rect 12362 3780 12394 3785
rect 12362 3775 12365 3780
rect 12171 3755 12365 3775
rect 12171 3750 12174 3755
rect 12142 3745 12174 3750
rect 12362 3750 12365 3755
rect 12391 3775 12394 3780
rect 12506 3780 12538 3785
rect 12506 3775 12509 3780
rect 12391 3755 12509 3775
rect 12391 3750 12394 3755
rect 12362 3745 12394 3750
rect 12506 3750 12509 3755
rect 12535 3750 12538 3780
rect 12506 3745 12538 3750
rect 11990 3730 12030 3735
rect 11250 3720 11290 3725
rect 11250 3690 11255 3720
rect 11285 3715 11290 3720
rect 11355 3720 11395 3725
rect 11355 3715 11360 3720
rect 11285 3695 11360 3715
rect 11285 3690 11290 3695
rect 11250 3685 11290 3690
rect 11355 3690 11360 3695
rect 11390 3715 11395 3720
rect 11470 3720 11510 3725
rect 11470 3715 11475 3720
rect 11390 3695 11475 3715
rect 11390 3690 11395 3695
rect 11355 3685 11395 3690
rect 11470 3690 11475 3695
rect 11505 3715 11510 3720
rect 11575 3720 11615 3725
rect 11575 3715 11580 3720
rect 11505 3695 11580 3715
rect 11505 3690 11510 3695
rect 11470 3685 11510 3690
rect 11575 3690 11580 3695
rect 11610 3715 11615 3720
rect 11690 3720 11730 3725
rect 11690 3715 11695 3720
rect 11610 3695 11695 3715
rect 11610 3690 11615 3695
rect 11575 3685 11615 3690
rect 11690 3690 11695 3695
rect 11725 3715 11730 3720
rect 11805 3720 11845 3725
rect 11805 3715 11810 3720
rect 11725 3695 11810 3715
rect 11725 3690 11730 3695
rect 11690 3685 11730 3690
rect 11805 3690 11810 3695
rect 11840 3690 11845 3720
rect 11990 3700 11995 3730
rect 12025 3725 12030 3730
rect 12210 3730 12250 3735
rect 12210 3725 12215 3730
rect 12025 3705 12215 3725
rect 12025 3700 12030 3705
rect 11990 3695 12030 3700
rect 12210 3700 12215 3705
rect 12245 3725 12250 3730
rect 12430 3730 12470 3735
rect 12430 3725 12435 3730
rect 12245 3705 12435 3725
rect 12245 3700 12250 3705
rect 12210 3695 12250 3700
rect 12430 3700 12435 3705
rect 12465 3725 12470 3730
rect 12860 3730 12900 3735
rect 12860 3725 12865 3730
rect 12465 3705 12865 3725
rect 12465 3700 12470 3705
rect 12430 3695 12470 3700
rect 12860 3700 12865 3705
rect 12895 3700 12900 3730
rect 12860 3695 12900 3700
rect 11805 3685 11845 3690
rect 12095 3685 12135 3690
rect 12095 3655 12100 3685
rect 12130 3680 12135 3685
rect 12315 3685 12355 3690
rect 12315 3680 12320 3685
rect 12130 3660 12320 3680
rect 12130 3655 12135 3660
rect 12095 3650 12135 3655
rect 12315 3655 12320 3660
rect 12350 3680 12355 3685
rect 12545 3685 12585 3690
rect 12545 3680 12550 3685
rect 12350 3660 12550 3680
rect 12350 3655 12355 3660
rect 12315 3650 12355 3655
rect 12545 3655 12550 3660
rect 12580 3680 12585 3685
rect 12805 3685 12845 3690
rect 12805 3680 12810 3685
rect 12580 3660 12810 3680
rect 12580 3655 12585 3660
rect 12545 3650 12585 3655
rect 12805 3655 12810 3660
rect 12840 3655 12845 3685
rect 12805 3650 12845 3655
rect 10210 3635 10250 3640
rect 10210 3605 10215 3635
rect 10245 3630 10250 3635
rect 10320 3635 10360 3640
rect 10320 3630 10325 3635
rect 10245 3610 10325 3630
rect 10245 3605 10250 3610
rect 10210 3600 10250 3605
rect 10320 3605 10325 3610
rect 10355 3630 10360 3635
rect 10430 3635 10470 3640
rect 10430 3630 10435 3635
rect 10355 3610 10435 3630
rect 10355 3605 10360 3610
rect 10320 3600 10360 3605
rect 10430 3605 10435 3610
rect 10465 3630 10470 3635
rect 10540 3635 10580 3640
rect 10540 3630 10545 3635
rect 10465 3610 10545 3630
rect 10465 3605 10470 3610
rect 10430 3600 10470 3605
rect 10540 3605 10545 3610
rect 10575 3630 10580 3635
rect 10650 3635 10690 3640
rect 10650 3630 10655 3635
rect 10575 3610 10655 3630
rect 10575 3605 10580 3610
rect 10540 3600 10580 3605
rect 10650 3605 10655 3610
rect 10685 3630 10690 3635
rect 10760 3635 10800 3640
rect 10760 3630 10765 3635
rect 10685 3610 10765 3630
rect 10685 3605 10690 3610
rect 10650 3600 10690 3605
rect 10760 3605 10765 3610
rect 10795 3605 10800 3635
rect 13000 3635 13040 3640
rect 10760 3600 10800 3605
rect 11340 3625 11380 3630
rect 11340 3595 11345 3625
rect 11375 3620 11380 3625
rect 11460 3625 11500 3630
rect 11460 3620 11465 3625
rect 11375 3600 11465 3620
rect 11375 3595 11380 3600
rect 11340 3590 11380 3595
rect 11460 3595 11465 3600
rect 11495 3620 11500 3625
rect 11580 3625 11620 3630
rect 11580 3620 11585 3625
rect 11495 3600 11585 3620
rect 11495 3595 11500 3600
rect 11460 3590 11500 3595
rect 11580 3595 11585 3600
rect 11615 3620 11620 3625
rect 11700 3625 11740 3630
rect 11700 3620 11705 3625
rect 11615 3600 11705 3620
rect 11615 3595 11620 3600
rect 11580 3590 11620 3595
rect 11700 3595 11705 3600
rect 11735 3620 11740 3625
rect 11820 3625 11860 3630
rect 11820 3620 11825 3625
rect 11735 3600 11825 3620
rect 11735 3595 11740 3600
rect 11700 3590 11740 3595
rect 11820 3595 11825 3600
rect 11855 3620 11860 3625
rect 11940 3625 11980 3630
rect 11940 3620 11945 3625
rect 11855 3600 11945 3620
rect 11855 3595 11860 3600
rect 11820 3590 11860 3595
rect 11940 3595 11945 3600
rect 11975 3620 11980 3625
rect 12060 3625 12100 3630
rect 12060 3620 12065 3625
rect 11975 3600 12065 3620
rect 11975 3595 11980 3600
rect 11940 3590 11980 3595
rect 12060 3595 12065 3600
rect 12095 3620 12100 3625
rect 12180 3625 12220 3630
rect 12180 3620 12185 3625
rect 12095 3600 12185 3620
rect 12095 3595 12100 3600
rect 12060 3590 12100 3595
rect 12180 3595 12185 3600
rect 12215 3620 12220 3625
rect 12300 3625 12340 3630
rect 12300 3620 12305 3625
rect 12215 3600 12305 3620
rect 12215 3595 12220 3600
rect 12180 3590 12220 3595
rect 12300 3595 12305 3600
rect 12335 3620 12340 3625
rect 12420 3625 12460 3630
rect 12420 3620 12425 3625
rect 12335 3600 12425 3620
rect 12335 3595 12340 3600
rect 12300 3590 12340 3595
rect 12420 3595 12425 3600
rect 12455 3595 12460 3625
rect 13000 3605 13005 3635
rect 13035 3630 13040 3635
rect 13110 3635 13150 3640
rect 13110 3630 13115 3635
rect 13035 3610 13115 3630
rect 13035 3605 13040 3610
rect 13000 3600 13040 3605
rect 13110 3605 13115 3610
rect 13145 3630 13150 3635
rect 13220 3635 13260 3640
rect 13220 3630 13225 3635
rect 13145 3610 13225 3630
rect 13145 3605 13150 3610
rect 13110 3600 13150 3605
rect 13220 3605 13225 3610
rect 13255 3630 13260 3635
rect 13330 3635 13370 3640
rect 13330 3630 13335 3635
rect 13255 3610 13335 3630
rect 13255 3605 13260 3610
rect 13220 3600 13260 3605
rect 13330 3605 13335 3610
rect 13365 3630 13370 3635
rect 13440 3635 13480 3640
rect 13440 3630 13445 3635
rect 13365 3610 13445 3630
rect 13365 3605 13370 3610
rect 13330 3600 13370 3605
rect 13440 3605 13445 3610
rect 13475 3630 13480 3635
rect 13550 3635 13590 3640
rect 13550 3630 13555 3635
rect 13475 3610 13555 3630
rect 13475 3605 13480 3610
rect 13440 3600 13480 3605
rect 13550 3605 13555 3610
rect 13585 3605 13590 3635
rect 13550 3600 13590 3605
rect 26340 3625 26380 3630
rect 12420 3590 12460 3595
rect 26340 3595 26345 3625
rect 26375 3620 26380 3625
rect 26460 3625 26500 3630
rect 26460 3620 26465 3625
rect 26375 3600 26465 3620
rect 26375 3595 26380 3600
rect 26340 3590 26380 3595
rect 26460 3595 26465 3600
rect 26495 3620 26500 3625
rect 26580 3625 26620 3630
rect 26580 3620 26585 3625
rect 26495 3600 26585 3620
rect 26495 3595 26500 3600
rect 26460 3590 26500 3595
rect 26580 3595 26585 3600
rect 26615 3620 26620 3625
rect 26700 3625 26740 3630
rect 26700 3620 26705 3625
rect 26615 3600 26705 3620
rect 26615 3595 26620 3600
rect 26580 3590 26620 3595
rect 26700 3595 26705 3600
rect 26735 3620 26740 3625
rect 26820 3625 26860 3630
rect 26820 3620 26825 3625
rect 26735 3600 26825 3620
rect 26735 3595 26740 3600
rect 26700 3590 26740 3595
rect 26820 3595 26825 3600
rect 26855 3620 26860 3625
rect 26940 3625 26980 3630
rect 26940 3620 26945 3625
rect 26855 3600 26945 3620
rect 26855 3595 26860 3600
rect 26820 3590 26860 3595
rect 26940 3595 26945 3600
rect 26975 3620 26980 3625
rect 27060 3625 27100 3630
rect 27060 3620 27065 3625
rect 26975 3600 27065 3620
rect 26975 3595 26980 3600
rect 26940 3590 26980 3595
rect 27060 3595 27065 3600
rect 27095 3620 27100 3625
rect 27180 3625 27220 3630
rect 27180 3620 27185 3625
rect 27095 3600 27185 3620
rect 27095 3595 27100 3600
rect 27060 3590 27100 3595
rect 27180 3595 27185 3600
rect 27215 3620 27220 3625
rect 27300 3625 27340 3630
rect 27300 3620 27305 3625
rect 27215 3600 27305 3620
rect 27215 3595 27220 3600
rect 27180 3590 27220 3595
rect 27300 3595 27305 3600
rect 27335 3620 27340 3625
rect 27420 3625 27460 3630
rect 27420 3620 27425 3625
rect 27335 3600 27425 3620
rect 27335 3595 27340 3600
rect 27300 3590 27340 3595
rect 27420 3595 27425 3600
rect 27455 3595 27460 3625
rect 27420 3590 27460 3595
rect 9899 3555 10040 3560
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 1261 3525 1301 3530
rect 1261 3520 1266 3525
rect -75 3500 1266 3520
rect -75 3495 -70 3500
rect -110 3490 -70 3495
rect 1261 3495 1266 3500
rect 1296 3495 1301 3525
rect 9899 3525 9905 3555
rect 9935 3525 9955 3555
rect 9985 3525 10005 3555
rect 10035 3525 10040 3555
rect 9899 3520 10040 3525
rect 13760 3555 13901 3560
rect 13760 3525 13765 3555
rect 13795 3525 13815 3555
rect 13845 3525 13865 3555
rect 13895 3525 13901 3555
rect 13760 3520 13901 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3440 5185 3445
rect 5550 3445 5590 3450
rect 5550 3440 5555 3445
rect 5175 3420 5555 3440
rect 5175 3415 5185 3420
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect 5550 3415 5555 3420
rect 5585 3415 5590 3445
rect 5550 3410 5590 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3335 1245 3340
rect 3135 3340 3175 3345
rect 3135 3335 3140 3340
rect 1240 3315 3140 3335
rect 1240 3310 1245 3315
rect 1205 3305 1245 3310
rect 3135 3310 3140 3315
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5360 3335 5400 3340
rect 5360 3330 5365 3335
rect 3425 3310 5365 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5360 3305 5365 3310
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 27945 3290 27985 3295
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3280 1200 3285
rect 4885 3285 4925 3290
rect 4885 3280 4890 3285
rect 1195 3260 4890 3280
rect 1195 3255 1200 3260
rect 1160 3250 1200 3255
rect 4885 3255 4890 3260
rect 4920 3280 4925 3285
rect 5410 3285 5450 3290
rect 5410 3280 5415 3285
rect 4920 3260 5415 3280
rect 4920 3255 4925 3260
rect 4885 3250 4925 3255
rect 5410 3255 5415 3260
rect 5445 3255 5450 3285
rect 27945 3260 27950 3290
rect 27980 3285 27985 3290
rect 28055 3290 28095 3295
rect 28055 3285 28060 3290
rect 27980 3265 28060 3285
rect 27980 3260 27985 3265
rect 27945 3255 27985 3260
rect 28055 3260 28060 3265
rect 28090 3285 28095 3290
rect 28165 3290 28205 3295
rect 28165 3285 28170 3290
rect 28090 3265 28170 3285
rect 28090 3260 28095 3265
rect 28055 3255 28095 3260
rect 28165 3260 28170 3265
rect 28200 3285 28205 3290
rect 28275 3290 28315 3295
rect 28275 3285 28280 3290
rect 28200 3265 28280 3285
rect 28200 3260 28205 3265
rect 28165 3255 28205 3260
rect 28275 3260 28280 3265
rect 28310 3285 28315 3290
rect 28385 3290 28425 3295
rect 28385 3285 28390 3290
rect 28310 3265 28390 3285
rect 28310 3260 28315 3265
rect 28275 3255 28315 3260
rect 28385 3260 28390 3265
rect 28420 3285 28425 3290
rect 28495 3290 28535 3295
rect 28495 3285 28500 3290
rect 28420 3265 28500 3285
rect 28420 3260 28425 3265
rect 28385 3255 28425 3260
rect 28495 3260 28500 3265
rect 28530 3285 28535 3290
rect 28605 3290 28645 3295
rect 28605 3285 28610 3290
rect 28530 3265 28610 3285
rect 28530 3260 28535 3265
rect 28495 3255 28535 3260
rect 28605 3260 28610 3265
rect 28640 3285 28645 3290
rect 28715 3290 28755 3295
rect 28715 3285 28720 3290
rect 28640 3265 28720 3285
rect 28640 3260 28645 3265
rect 28605 3255 28645 3260
rect 28715 3260 28720 3265
rect 28750 3285 28755 3290
rect 28825 3290 28865 3295
rect 28825 3285 28830 3290
rect 28750 3265 28830 3285
rect 28750 3260 28755 3265
rect 28715 3255 28755 3260
rect 28825 3260 28830 3265
rect 28860 3285 28865 3290
rect 28935 3290 28975 3295
rect 28935 3285 28940 3290
rect 28860 3265 28940 3285
rect 28860 3260 28865 3265
rect 28825 3255 28865 3260
rect 28935 3260 28940 3265
rect 28970 3285 28975 3290
rect 29045 3290 29085 3295
rect 29045 3285 29050 3290
rect 28970 3265 29050 3285
rect 28970 3260 28975 3265
rect 28935 3255 28975 3260
rect 29045 3260 29050 3265
rect 29080 3260 29085 3290
rect 29045 3255 29085 3260
rect 5410 3250 5450 3255
rect 2735 3240 2775 3245
rect 2735 3235 2740 3240
rect 46 3215 2740 3235
rect 46 3205 91 3215
rect 2735 3210 2740 3215
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 25580 3210 25620 3215
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3180 2660 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2655 3160 4445 3180
rect 2655 3155 2660 3160
rect 2620 3150 2660 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 25580 3180 25585 3210
rect 25615 3205 25620 3210
rect 25980 3210 26015 3215
rect 25980 3205 25985 3210
rect 25615 3185 25985 3205
rect 25615 3180 25620 3185
rect 25580 3175 25620 3180
rect 25980 3180 25985 3185
rect 25980 3175 26015 3180
rect 4440 3150 4480 3155
rect 11050 3155 11090 3160
rect -110 3140 -70 3145
rect -110 3110 -105 3140
rect -75 3135 -70 3140
rect 46 3135 51 3145
rect -75 3115 51 3135
rect -75 3110 -70 3115
rect 46 3110 51 3115
rect 86 3110 91 3145
rect 3135 3140 3175 3145
rect -110 3105 -70 3110
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 3135 3110 3140 3140
rect 3170 3135 3175 3140
rect 4835 3140 4875 3145
rect 4835 3135 4840 3140
rect 3170 3115 4840 3135
rect 3170 3110 3175 3115
rect 3135 3105 3175 3110
rect 4835 3110 4840 3115
rect 4870 3135 4875 3140
rect 5315 3140 5355 3145
rect 5315 3135 5320 3140
rect 4870 3115 5320 3135
rect 4870 3110 4875 3115
rect 4835 3105 4875 3110
rect 5315 3110 5320 3115
rect 5350 3110 5355 3140
rect 11050 3125 11055 3155
rect 11085 3150 11090 3155
rect 11823 3155 11857 3160
rect 11823 3150 11826 3155
rect 11085 3130 11826 3150
rect 11085 3125 11090 3130
rect 11050 3120 11090 3125
rect 11823 3125 11826 3130
rect 11854 3125 11857 3155
rect 11823 3120 11857 3125
rect 25900 3155 25940 3160
rect 25900 3125 25905 3155
rect 25935 3150 25940 3155
rect 26823 3155 26857 3160
rect 26823 3150 26826 3155
rect 25935 3130 26826 3150
rect 25935 3125 25940 3130
rect 25900 3120 25940 3125
rect 26823 3125 26826 3130
rect 26854 3125 26857 3155
rect 26823 3120 26857 3125
rect 5315 3105 5355 3110
rect 1160 3100 1200 3105
rect 1160 3095 1165 3100
rect 46 3075 1165 3095
rect 46 3065 91 3075
rect 1160 3070 1165 3075
rect 1195 3070 1200 3100
rect 11280 3100 11320 3105
rect 1160 3065 1200 3070
rect 3985 3080 4025 3085
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 3985 3050 3990 3080
rect 4020 3075 4025 3080
rect 4020 3055 6100 3075
rect 11280 3070 11285 3100
rect 11315 3095 11320 3100
rect 11520 3100 11560 3105
rect 11520 3095 11525 3100
rect 11315 3075 11525 3095
rect 11315 3070 11320 3075
rect 11280 3065 11320 3070
rect 11520 3070 11525 3075
rect 11555 3095 11560 3100
rect 11760 3100 11800 3105
rect 11760 3095 11765 3100
rect 11555 3075 11765 3095
rect 11555 3070 11560 3075
rect 11520 3065 11560 3070
rect 11760 3070 11765 3075
rect 11795 3095 11800 3100
rect 12000 3100 12040 3105
rect 12000 3095 12005 3100
rect 11795 3075 12005 3095
rect 11795 3070 11800 3075
rect 11760 3065 11800 3070
rect 12000 3070 12005 3075
rect 12035 3095 12040 3100
rect 12240 3100 12280 3105
rect 12240 3095 12245 3100
rect 12035 3075 12245 3095
rect 12035 3070 12040 3075
rect 12000 3065 12040 3070
rect 12240 3070 12245 3075
rect 12275 3095 12280 3100
rect 12480 3100 12520 3105
rect 12480 3095 12485 3100
rect 12275 3075 12485 3095
rect 12275 3070 12280 3075
rect 12240 3065 12280 3070
rect 12480 3070 12485 3075
rect 12515 3070 12520 3100
rect 12480 3065 12520 3070
rect 26280 3100 26320 3105
rect 26280 3070 26285 3100
rect 26315 3095 26320 3100
rect 26520 3100 26560 3105
rect 26520 3095 26525 3100
rect 26315 3075 26525 3095
rect 26315 3070 26320 3075
rect 26280 3065 26320 3070
rect 26520 3070 26525 3075
rect 26555 3095 26560 3100
rect 26760 3100 26800 3105
rect 26760 3095 26765 3100
rect 26555 3075 26765 3095
rect 26555 3070 26560 3075
rect 26520 3065 26560 3070
rect 26760 3070 26765 3075
rect 26795 3095 26800 3100
rect 27000 3100 27040 3105
rect 27000 3095 27005 3100
rect 26795 3075 27005 3095
rect 26795 3070 26800 3075
rect 26760 3065 26800 3070
rect 27000 3070 27005 3075
rect 27035 3095 27040 3100
rect 27240 3100 27280 3105
rect 27240 3095 27245 3100
rect 27035 3075 27245 3095
rect 27035 3070 27040 3075
rect 27000 3065 27040 3070
rect 27240 3070 27245 3075
rect 27275 3095 27280 3100
rect 27480 3100 27520 3105
rect 27480 3095 27485 3100
rect 27275 3075 27485 3095
rect 27275 3070 27280 3075
rect 27240 3065 27280 3070
rect 27480 3070 27485 3075
rect 27515 3070 27520 3100
rect 27480 3065 27520 3070
rect 11400 3055 11440 3060
rect 4020 3050 4025 3055
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3030 3485 3035
rect 3805 3035 3845 3040
rect 3805 3030 3810 3035
rect 3480 3010 3810 3030
rect 3480 3005 3485 3010
rect -110 3000 -70 3005
rect -110 2970 -105 3000
rect -75 2995 -70 3000
rect 46 2995 51 3005
rect -75 2975 51 2995
rect -75 2970 -70 2975
rect 46 2970 51 2975
rect 86 2970 91 3005
rect 3445 3000 3485 3005
rect 3805 3005 3810 3010
rect 3840 3030 3845 3035
rect 4345 3035 4385 3040
rect 4345 3030 4350 3035
rect 3840 3010 4350 3030
rect 3840 3005 3845 3010
rect 3805 3000 3845 3005
rect 4345 3005 4350 3010
rect 4380 3030 4385 3035
rect 4705 3035 4745 3040
rect 4705 3030 4710 3035
rect 4380 3010 4710 3030
rect 4380 3005 4385 3010
rect 4345 3000 4385 3005
rect 4705 3005 4710 3010
rect 4740 3030 4745 3035
rect 4740 3010 6100 3030
rect 11400 3025 11405 3055
rect 11435 3050 11440 3055
rect 11640 3055 11680 3060
rect 11640 3050 11645 3055
rect 11435 3030 11645 3050
rect 11435 3025 11440 3030
rect 11400 3020 11440 3025
rect 11640 3025 11645 3030
rect 11675 3050 11680 3055
rect 11880 3055 11920 3060
rect 11880 3050 11885 3055
rect 11675 3030 11885 3050
rect 11675 3025 11680 3030
rect 11640 3020 11680 3025
rect 11880 3025 11885 3030
rect 11915 3050 11920 3055
rect 12120 3055 12160 3060
rect 12120 3050 12125 3055
rect 11915 3030 12125 3050
rect 11915 3025 11920 3030
rect 11880 3020 11920 3025
rect 12120 3025 12125 3030
rect 12155 3050 12160 3055
rect 12360 3055 12400 3060
rect 12360 3050 12365 3055
rect 12155 3030 12365 3050
rect 12155 3025 12160 3030
rect 12120 3020 12160 3025
rect 12360 3025 12365 3030
rect 12395 3025 12400 3055
rect 12360 3020 12400 3025
rect 26400 3055 26440 3060
rect 26400 3025 26405 3055
rect 26435 3050 26440 3055
rect 26640 3055 26680 3060
rect 26640 3050 26645 3055
rect 26435 3030 26645 3050
rect 26435 3025 26440 3030
rect 26400 3020 26440 3025
rect 26640 3025 26645 3030
rect 26675 3050 26680 3055
rect 26880 3055 26920 3060
rect 26880 3050 26885 3055
rect 26675 3030 26885 3050
rect 26675 3025 26680 3030
rect 26640 3020 26680 3025
rect 26880 3025 26885 3030
rect 26915 3050 26920 3055
rect 27120 3055 27160 3060
rect 27120 3050 27125 3055
rect 26915 3030 27125 3050
rect 26915 3025 26920 3030
rect 26880 3020 26920 3025
rect 27120 3025 27125 3030
rect 27155 3050 27160 3055
rect 27360 3055 27400 3060
rect 27360 3050 27365 3055
rect 27155 3030 27365 3050
rect 27155 3025 27160 3030
rect 27120 3020 27160 3025
rect 27360 3025 27365 3030
rect 27395 3025 27400 3055
rect 27360 3020 27400 3025
rect 4740 3005 4745 3010
rect 4705 3000 4745 3005
rect 11340 3000 11380 3005
rect 2520 2980 2560 2985
rect -110 2965 -70 2970
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2520 2950 2525 2980
rect 2555 2975 2560 2980
rect 3080 2980 3120 2985
rect 3080 2975 3085 2980
rect 2555 2955 3085 2975
rect 2555 2950 2560 2955
rect 2520 2945 2560 2950
rect 3080 2950 3085 2955
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2975 3305 2980
rect 3625 2980 3665 2985
rect 3625 2975 3630 2980
rect 3300 2955 3630 2975
rect 3300 2950 3305 2955
rect 3265 2945 3305 2950
rect 3625 2950 3630 2955
rect 3660 2975 3665 2980
rect 4165 2980 4205 2985
rect 4165 2975 4170 2980
rect 3660 2955 4170 2975
rect 3660 2950 3665 2955
rect 3625 2945 3665 2950
rect 4165 2950 4170 2955
rect 4200 2975 4205 2980
rect 4525 2980 4565 2985
rect 4525 2975 4530 2980
rect 4200 2955 4530 2975
rect 4200 2950 4205 2955
rect 4165 2945 4205 2950
rect 4525 2950 4530 2955
rect 4560 2975 4565 2980
rect 4560 2955 6100 2975
rect 11340 2970 11345 3000
rect 11375 2995 11380 3000
rect 11400 3000 11440 3005
rect 11400 2995 11405 3000
rect 11375 2975 11405 2995
rect 11375 2970 11380 2975
rect 10265 2965 10305 2970
rect 4560 2950 4565 2955
rect 4525 2945 4565 2950
rect 2425 2920 2465 2925
rect 9899 2935 10040 2940
rect -110 2910 -70 2915
rect -110 2880 -105 2910
rect -75 2905 -70 2910
rect 905 2910 1125 2920
rect 905 2905 920 2910
rect -75 2885 920 2905
rect -75 2880 -70 2885
rect -110 2875 -70 2880
rect 905 2880 920 2885
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 9899 2905 9905 2935
rect 9935 2905 9955 2935
rect 9985 2905 10005 2935
rect 10035 2905 10040 2935
rect 10265 2935 10270 2965
rect 10300 2960 10305 2965
rect 10375 2965 10415 2970
rect 10375 2960 10380 2965
rect 10300 2940 10380 2960
rect 10300 2935 10305 2940
rect 10265 2930 10305 2935
rect 10375 2935 10380 2940
rect 10410 2960 10415 2965
rect 10485 2965 10525 2970
rect 10485 2960 10490 2965
rect 10410 2940 10490 2960
rect 10410 2935 10415 2940
rect 10375 2930 10415 2935
rect 10485 2935 10490 2940
rect 10520 2960 10525 2965
rect 10595 2965 10635 2970
rect 10595 2960 10600 2965
rect 10520 2940 10600 2960
rect 10520 2935 10525 2940
rect 10485 2930 10525 2935
rect 10595 2935 10600 2940
rect 10630 2960 10635 2965
rect 10705 2965 10745 2970
rect 11340 2965 11380 2970
rect 11400 2970 11405 2975
rect 11435 2995 11440 3000
rect 11580 3000 11620 3005
rect 11580 2995 11585 3000
rect 11435 2975 11585 2995
rect 11435 2970 11440 2975
rect 11400 2965 11440 2970
rect 11580 2970 11585 2975
rect 11615 2995 11620 3000
rect 11820 3000 11860 3005
rect 11820 2995 11825 3000
rect 11615 2975 11825 2995
rect 11615 2970 11620 2975
rect 11580 2965 11620 2970
rect 11820 2970 11825 2975
rect 11855 2995 11860 3000
rect 12060 3000 12100 3005
rect 12060 2995 12065 3000
rect 11855 2975 12065 2995
rect 11855 2970 11860 2975
rect 11820 2965 11860 2970
rect 12060 2970 12065 2975
rect 12095 2995 12100 3000
rect 12300 3000 12340 3005
rect 12300 2995 12305 3000
rect 12095 2975 12305 2995
rect 12095 2970 12100 2975
rect 12060 2965 12100 2970
rect 12300 2970 12305 2975
rect 12335 2970 12340 3000
rect 26340 3000 26380 3005
rect 26340 2970 26345 3000
rect 26375 2995 26380 3000
rect 26400 3000 26440 3005
rect 26400 2995 26405 3000
rect 26375 2975 26405 2995
rect 26375 2970 26380 2975
rect 12300 2965 12340 2970
rect 13055 2965 13095 2970
rect 10705 2960 10710 2965
rect 10630 2940 10710 2960
rect 10630 2935 10635 2940
rect 10595 2930 10635 2935
rect 10705 2935 10710 2940
rect 10740 2935 10745 2965
rect 10705 2930 10745 2935
rect 11460 2945 11500 2950
rect 11460 2915 11465 2945
rect 11495 2940 11500 2945
rect 11700 2945 11740 2950
rect 11700 2940 11705 2945
rect 11495 2920 11705 2940
rect 11495 2915 11500 2920
rect 11460 2910 11500 2915
rect 11700 2915 11705 2920
rect 11735 2940 11740 2945
rect 11940 2945 11980 2950
rect 11940 2940 11945 2945
rect 11735 2920 11945 2940
rect 11735 2915 11740 2920
rect 11700 2910 11740 2915
rect 11940 2915 11945 2920
rect 11975 2940 11980 2945
rect 12180 2945 12220 2950
rect 12180 2940 12185 2945
rect 11975 2920 12185 2940
rect 11975 2915 11980 2920
rect 11940 2910 11980 2915
rect 12180 2915 12185 2920
rect 12215 2940 12220 2945
rect 12420 2945 12460 2950
rect 12420 2940 12425 2945
rect 12215 2920 12425 2940
rect 12215 2915 12220 2920
rect 12180 2910 12220 2915
rect 12420 2915 12425 2920
rect 12455 2940 12460 2945
rect 12480 2945 12520 2950
rect 12480 2940 12485 2945
rect 12455 2920 12485 2940
rect 12455 2915 12460 2920
rect 12420 2910 12460 2915
rect 12480 2915 12485 2920
rect 12515 2915 12520 2945
rect 13055 2935 13060 2965
rect 13090 2960 13095 2965
rect 13165 2965 13205 2970
rect 13165 2960 13170 2965
rect 13090 2940 13170 2960
rect 13090 2935 13095 2940
rect 13055 2930 13095 2935
rect 13165 2935 13170 2940
rect 13200 2960 13205 2965
rect 13275 2965 13315 2970
rect 13275 2960 13280 2965
rect 13200 2940 13280 2960
rect 13200 2935 13205 2940
rect 13165 2930 13205 2935
rect 13275 2935 13280 2940
rect 13310 2960 13315 2965
rect 13385 2965 13425 2970
rect 13385 2960 13390 2965
rect 13310 2940 13390 2960
rect 13310 2935 13315 2940
rect 13275 2930 13315 2935
rect 13385 2935 13390 2940
rect 13420 2960 13425 2965
rect 13495 2965 13535 2970
rect 26340 2965 26380 2970
rect 26400 2970 26405 2975
rect 26435 2995 26440 3000
rect 26580 3000 26620 3005
rect 26580 2995 26585 3000
rect 26435 2975 26585 2995
rect 26435 2970 26440 2975
rect 26400 2965 26440 2970
rect 26580 2970 26585 2975
rect 26615 2995 26620 3000
rect 26820 3000 26860 3005
rect 26820 2995 26825 3000
rect 26615 2975 26825 2995
rect 26615 2970 26620 2975
rect 26580 2965 26620 2970
rect 26820 2970 26825 2975
rect 26855 2995 26860 3000
rect 27060 3000 27100 3005
rect 27060 2995 27065 3000
rect 26855 2975 27065 2995
rect 26855 2970 26860 2975
rect 26820 2965 26860 2970
rect 27060 2970 27065 2975
rect 27095 2995 27100 3000
rect 27300 3000 27340 3005
rect 27300 2995 27305 3000
rect 27095 2975 27305 2995
rect 27095 2970 27100 2975
rect 27060 2965 27100 2970
rect 27300 2970 27305 2975
rect 27335 2970 27340 3000
rect 27300 2965 27340 2970
rect 13495 2960 13500 2965
rect 13420 2940 13500 2960
rect 13420 2935 13425 2940
rect 13385 2930 13425 2935
rect 13495 2935 13500 2940
rect 13530 2935 13535 2965
rect 26460 2945 26500 2950
rect 13495 2930 13535 2935
rect 13760 2935 13901 2940
rect 12480 2910 12520 2915
rect 905 2870 1125 2880
rect 2330 2900 2375 2905
rect 9899 2900 10040 2905
rect 13760 2905 13765 2935
rect 13795 2905 13815 2935
rect 13845 2905 13865 2935
rect 13895 2905 13901 2935
rect 26460 2915 26465 2945
rect 26495 2940 26500 2945
rect 26700 2945 26740 2950
rect 26700 2940 26705 2945
rect 26495 2920 26705 2940
rect 26495 2915 26500 2920
rect 26460 2910 26500 2915
rect 26700 2915 26705 2920
rect 26735 2940 26740 2945
rect 26940 2945 26980 2950
rect 26940 2940 26945 2945
rect 26735 2920 26945 2940
rect 26735 2915 26740 2920
rect 26700 2910 26740 2915
rect 26940 2915 26945 2920
rect 26975 2940 26980 2945
rect 27180 2945 27220 2950
rect 27180 2940 27185 2945
rect 26975 2920 27185 2940
rect 26975 2915 26980 2920
rect 26940 2910 26980 2915
rect 27180 2915 27185 2920
rect 27215 2940 27220 2945
rect 27420 2945 27460 2950
rect 27420 2940 27425 2945
rect 27215 2920 27425 2940
rect 27215 2915 27220 2920
rect 27180 2910 27220 2915
rect 27420 2915 27425 2920
rect 27455 2940 27460 2945
rect 27480 2945 27520 2950
rect 27480 2940 27485 2945
rect 27455 2920 27485 2940
rect 27455 2915 27460 2920
rect 27420 2910 27460 2915
rect 27480 2915 27485 2920
rect 27515 2915 27520 2945
rect 27480 2910 27520 2915
rect 28000 2920 28040 2925
rect 13760 2900 13901 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 28000 2890 28005 2920
rect 28035 2915 28040 2920
rect 28110 2920 28150 2925
rect 28110 2915 28115 2920
rect 28035 2895 28115 2915
rect 28035 2890 28040 2895
rect 28000 2885 28040 2890
rect 28110 2890 28115 2895
rect 28145 2915 28150 2920
rect 28220 2920 28260 2925
rect 28220 2915 28225 2920
rect 28145 2895 28225 2915
rect 28145 2890 28150 2895
rect 28110 2885 28150 2890
rect 28220 2890 28225 2895
rect 28255 2915 28260 2920
rect 28330 2920 28370 2925
rect 28330 2915 28335 2920
rect 28255 2895 28335 2915
rect 28255 2890 28260 2895
rect 28220 2885 28260 2890
rect 28330 2890 28335 2895
rect 28365 2915 28370 2920
rect 28440 2920 28480 2925
rect 28440 2915 28445 2920
rect 28365 2895 28445 2915
rect 28365 2890 28370 2895
rect 28330 2885 28370 2890
rect 28440 2890 28445 2895
rect 28475 2915 28480 2920
rect 28550 2920 28590 2925
rect 28550 2915 28555 2920
rect 28475 2895 28555 2915
rect 28475 2890 28480 2895
rect 28440 2885 28480 2890
rect 28550 2890 28555 2895
rect 28585 2915 28590 2920
rect 28660 2920 28700 2925
rect 28660 2915 28665 2920
rect 28585 2895 28665 2915
rect 28585 2890 28590 2895
rect 28550 2885 28590 2890
rect 28660 2890 28665 2895
rect 28695 2915 28700 2920
rect 28770 2920 28810 2925
rect 28770 2915 28775 2920
rect 28695 2895 28775 2915
rect 28695 2890 28700 2895
rect 28660 2885 28700 2890
rect 28770 2890 28775 2895
rect 28805 2915 28810 2920
rect 28880 2920 28920 2925
rect 28880 2915 28885 2920
rect 28805 2895 28885 2915
rect 28805 2890 28810 2895
rect 28770 2885 28810 2890
rect 28880 2890 28885 2895
rect 28915 2915 28920 2920
rect 28990 2920 29030 2925
rect 28990 2915 28995 2920
rect 28915 2895 28995 2915
rect 28915 2890 28920 2895
rect 28880 2885 28920 2890
rect 28990 2890 28995 2895
rect 29025 2890 29030 2920
rect 28990 2885 29030 2890
rect 2330 2860 2375 2865
rect 9950 2880 9990 2885
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 51 2850 56 2855
rect -25 2830 56 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 51 2820 56 2830
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2845 769 2855
rect 1205 2850 1245 2855
rect 1205 2845 1210 2850
rect 764 2825 1210 2845
rect 764 2820 769 2825
rect 1205 2820 1210 2825
rect 1240 2820 1245 2850
rect 9950 2850 9955 2880
rect 9985 2875 9990 2880
rect 10650 2880 10690 2885
rect 10650 2875 10655 2880
rect 9985 2855 10655 2875
rect 9985 2850 9990 2855
rect 9950 2845 9990 2850
rect 10650 2850 10655 2855
rect 10685 2875 10690 2880
rect 11000 2880 11040 2885
rect 11000 2875 11005 2880
rect 10685 2855 11005 2875
rect 10685 2850 10690 2855
rect 10650 2845 10690 2850
rect 11000 2850 11005 2855
rect 11035 2850 11040 2880
rect 11000 2845 11040 2850
rect 12690 2880 12730 2885
rect 12690 2850 12695 2880
rect 12725 2875 12730 2880
rect 13110 2880 13150 2885
rect 13110 2875 13115 2880
rect 12725 2855 13115 2875
rect 12725 2850 12730 2855
rect 12690 2845 12730 2850
rect 13110 2850 13115 2855
rect 13145 2875 13150 2880
rect 13810 2880 13850 2885
rect 13810 2875 13815 2880
rect 13145 2855 13815 2875
rect 13145 2850 13150 2855
rect 13110 2845 13150 2850
rect 13810 2850 13815 2855
rect 13845 2850 13850 2880
rect 13810 2845 13850 2850
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 28055 2830 28095 2836
rect 9745 2825 9785 2830
rect 2330 2800 2370 2805
rect 2995 2810 3035 2815
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 51 2785 56 2795
rect 20 2765 56 2785
rect -15 2760 25 2765
rect 51 2760 56 2765
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2785 769 2795
rect 2620 2790 2660 2795
rect 2620 2785 2625 2790
rect 764 2765 2625 2785
rect 764 2760 769 2765
rect 2620 2760 2625 2765
rect 2655 2760 2660 2790
rect 2995 2780 3000 2810
rect 3030 2805 3035 2810
rect 3175 2810 3215 2815
rect 3175 2805 3180 2810
rect 3030 2785 3180 2805
rect 3030 2780 3035 2785
rect 2995 2775 3035 2780
rect 3175 2780 3180 2785
rect 3210 2805 3215 2810
rect 3355 2810 3395 2815
rect 3355 2805 3360 2810
rect 3210 2785 3360 2805
rect 3210 2780 3215 2785
rect 3175 2775 3215 2780
rect 3355 2780 3360 2785
rect 3390 2805 3395 2810
rect 3535 2810 3575 2815
rect 3535 2805 3540 2810
rect 3390 2785 3540 2805
rect 3390 2780 3395 2785
rect 3355 2775 3395 2780
rect 3535 2780 3540 2785
rect 3570 2805 3575 2810
rect 3715 2810 3755 2815
rect 3715 2805 3720 2810
rect 3570 2785 3720 2805
rect 3570 2780 3575 2785
rect 3535 2775 3575 2780
rect 3715 2780 3720 2785
rect 3750 2805 3755 2810
rect 3895 2810 3935 2815
rect 3895 2805 3900 2810
rect 3750 2785 3900 2805
rect 3750 2780 3755 2785
rect 3715 2775 3755 2780
rect 3895 2780 3900 2785
rect 3930 2805 3935 2810
rect 4075 2810 4115 2815
rect 4075 2805 4080 2810
rect 3930 2785 4080 2805
rect 3930 2780 3935 2785
rect 3895 2775 3935 2780
rect 4075 2780 4080 2785
rect 4110 2805 4115 2810
rect 4255 2810 4295 2815
rect 4255 2805 4260 2810
rect 4110 2785 4260 2805
rect 4110 2780 4115 2785
rect 4075 2775 4115 2780
rect 4255 2780 4260 2785
rect 4290 2805 4295 2810
rect 4435 2810 4475 2815
rect 4435 2805 4440 2810
rect 4290 2785 4440 2805
rect 4290 2780 4295 2785
rect 4255 2775 4295 2780
rect 4435 2780 4440 2785
rect 4470 2805 4475 2810
rect 4615 2810 4655 2815
rect 4615 2805 4620 2810
rect 4470 2785 4620 2805
rect 4470 2780 4475 2785
rect 4435 2775 4475 2780
rect 4615 2780 4620 2785
rect 4650 2805 4655 2810
rect 4795 2810 4835 2815
rect 4795 2805 4800 2810
rect 4650 2785 4800 2805
rect 4650 2780 4655 2785
rect 4615 2775 4655 2780
rect 4795 2780 4800 2785
rect 4830 2805 4835 2810
rect 4975 2810 5015 2815
rect 4975 2805 4980 2810
rect 4830 2785 4980 2805
rect 4830 2780 4835 2785
rect 4795 2775 4835 2780
rect 4975 2780 4980 2785
rect 5010 2805 5015 2810
rect 5550 2810 5590 2815
rect 5550 2805 5555 2810
rect 5010 2785 5555 2805
rect 5010 2780 5015 2785
rect 4975 2775 5015 2780
rect 5550 2780 5555 2785
rect 5585 2780 5590 2810
rect 9745 2795 9750 2825
rect 9780 2820 9785 2825
rect 10375 2825 10415 2830
rect 10375 2820 10380 2825
rect 9780 2800 10380 2820
rect 9780 2795 9785 2800
rect 9745 2790 9785 2795
rect 10375 2795 10380 2800
rect 10410 2795 10415 2825
rect 10375 2790 10415 2795
rect 13385 2825 13425 2830
rect 13385 2795 13390 2825
rect 13420 2820 13425 2825
rect 14015 2825 14055 2830
rect 14015 2820 14020 2825
rect 13420 2800 14020 2820
rect 13420 2795 13425 2800
rect 13385 2790 13425 2795
rect 14015 2795 14020 2800
rect 14050 2795 14055 2825
rect 14015 2790 14055 2795
rect 28055 2800 28060 2830
rect 28090 2800 28095 2830
rect 5550 2775 5590 2780
rect 28055 2780 28095 2800
rect 2620 2755 2660 2760
rect 3175 2750 3215 2755
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2740 1301 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1296 2720 2155 2740
rect 1296 2715 1301 2720
rect 1261 2710 1301 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 3175 2720 3180 2750
rect 3210 2745 3215 2750
rect 3355 2750 3395 2755
rect 3355 2745 3360 2750
rect 3210 2725 3360 2745
rect 3210 2720 3215 2725
rect 3175 2715 3215 2720
rect 3355 2720 3360 2725
rect 3390 2745 3395 2750
rect 3535 2750 3575 2755
rect 3535 2745 3540 2750
rect 3390 2725 3540 2745
rect 3390 2720 3395 2725
rect 3355 2715 3395 2720
rect 3535 2720 3540 2725
rect 3570 2745 3575 2750
rect 3715 2750 3755 2755
rect 3715 2745 3720 2750
rect 3570 2725 3720 2745
rect 3570 2720 3575 2725
rect 3535 2715 3575 2720
rect 3715 2720 3720 2725
rect 3750 2745 3755 2750
rect 3895 2750 3935 2755
rect 3895 2745 3900 2750
rect 3750 2725 3900 2745
rect 3750 2720 3755 2725
rect 3715 2715 3755 2720
rect 3895 2720 3900 2725
rect 3930 2745 3935 2750
rect 4075 2750 4115 2755
rect 4075 2745 4080 2750
rect 3930 2725 4080 2745
rect 3930 2720 3935 2725
rect 3895 2715 3935 2720
rect 4075 2720 4080 2725
rect 4110 2745 4115 2750
rect 4255 2750 4295 2755
rect 4255 2745 4260 2750
rect 4110 2725 4260 2745
rect 4110 2720 4115 2725
rect 4075 2715 4115 2720
rect 4255 2720 4260 2725
rect 4290 2745 4295 2750
rect 4435 2750 4475 2755
rect 4435 2745 4440 2750
rect 4290 2725 4440 2745
rect 4290 2720 4295 2725
rect 4255 2715 4295 2720
rect 4435 2720 4440 2725
rect 4470 2745 4475 2750
rect 4615 2750 4655 2755
rect 4615 2745 4620 2750
rect 4470 2725 4620 2745
rect 4470 2720 4475 2725
rect 4435 2715 4475 2720
rect 4615 2720 4620 2725
rect 4650 2745 4655 2750
rect 4795 2750 4835 2755
rect 4795 2745 4800 2750
rect 4650 2725 4800 2745
rect 4650 2720 4655 2725
rect 4615 2715 4655 2720
rect 4795 2720 4800 2725
rect 4830 2720 4835 2750
rect 28055 2750 28060 2780
rect 28090 2750 28095 2780
rect 4795 2715 4835 2720
rect 27690 2730 27730 2735
rect 2150 2710 2190 2715
rect 10210 2705 10250 2710
rect 10210 2675 10215 2705
rect 10245 2700 10250 2705
rect 10320 2705 10360 2710
rect 10320 2700 10325 2705
rect 10245 2680 10325 2700
rect 10245 2675 10250 2680
rect 10210 2670 10250 2675
rect 10320 2675 10325 2680
rect 10355 2700 10360 2705
rect 10430 2705 10470 2710
rect 10430 2700 10435 2705
rect 10355 2680 10435 2700
rect 10355 2675 10360 2680
rect 10320 2670 10360 2675
rect 10430 2675 10435 2680
rect 10465 2700 10470 2705
rect 10540 2705 10580 2710
rect 10540 2700 10545 2705
rect 10465 2680 10545 2700
rect 10465 2675 10470 2680
rect 10430 2670 10470 2675
rect 10540 2675 10545 2680
rect 10575 2700 10580 2705
rect 10650 2705 10690 2710
rect 10650 2700 10655 2705
rect 10575 2680 10655 2700
rect 10575 2675 10580 2680
rect 10540 2670 10580 2675
rect 10650 2675 10655 2680
rect 10685 2700 10690 2705
rect 10760 2705 10800 2710
rect 10760 2700 10765 2705
rect 10685 2680 10765 2700
rect 10685 2675 10690 2680
rect 10650 2670 10690 2675
rect 10760 2675 10765 2680
rect 10795 2675 10800 2705
rect 10760 2670 10800 2675
rect 13000 2705 13040 2710
rect 13000 2675 13005 2705
rect 13035 2700 13040 2705
rect 13110 2705 13150 2710
rect 13110 2700 13115 2705
rect 13035 2680 13115 2700
rect 13035 2675 13040 2680
rect 13000 2670 13040 2675
rect 13110 2675 13115 2680
rect 13145 2700 13150 2705
rect 13220 2705 13260 2710
rect 13220 2700 13225 2705
rect 13145 2680 13225 2700
rect 13145 2675 13150 2680
rect 13110 2670 13150 2675
rect 13220 2675 13225 2680
rect 13255 2700 13260 2705
rect 13330 2705 13370 2710
rect 13330 2700 13335 2705
rect 13255 2680 13335 2700
rect 13255 2675 13260 2680
rect 13220 2670 13260 2675
rect 13330 2675 13335 2680
rect 13365 2700 13370 2705
rect 13440 2705 13480 2710
rect 13440 2700 13445 2705
rect 13365 2680 13445 2700
rect 13365 2675 13370 2680
rect 13330 2670 13370 2675
rect 13440 2675 13445 2680
rect 13475 2700 13480 2705
rect 13550 2705 13590 2710
rect 13550 2700 13555 2705
rect 13475 2680 13555 2700
rect 13475 2675 13480 2680
rect 13440 2670 13480 2675
rect 13550 2675 13555 2680
rect 13585 2675 13590 2705
rect 27690 2700 27695 2730
rect 27725 2725 27730 2730
rect 28055 2730 28095 2750
rect 28055 2725 28060 2730
rect 27725 2705 28060 2725
rect 27725 2700 27730 2705
rect 27690 2695 27730 2700
rect 28055 2700 28060 2705
rect 28090 2700 28095 2730
rect 28055 2695 28095 2700
rect 13550 2670 13590 2675
rect 24735 2670 24775 2675
rect 24735 2640 24740 2670
rect 24770 2665 24775 2670
rect 24845 2670 24885 2675
rect 24845 2665 24850 2670
rect 24770 2645 24850 2665
rect 24770 2640 24775 2645
rect 24735 2635 24775 2640
rect 24845 2640 24850 2645
rect 24880 2665 24885 2670
rect 24955 2670 24995 2675
rect 24955 2665 24960 2670
rect 24880 2645 24960 2665
rect 24880 2640 24885 2645
rect 24845 2635 24885 2640
rect 24955 2640 24960 2645
rect 24990 2665 24995 2670
rect 25065 2670 25105 2675
rect 25065 2665 25070 2670
rect 24990 2645 25070 2665
rect 24990 2640 24995 2645
rect 24955 2635 24995 2640
rect 25065 2640 25070 2645
rect 25100 2665 25105 2670
rect 25175 2670 25215 2675
rect 25175 2665 25180 2670
rect 25100 2645 25180 2665
rect 25100 2640 25105 2645
rect 25065 2635 25105 2640
rect 25175 2640 25180 2645
rect 25210 2665 25215 2670
rect 25285 2670 25325 2675
rect 25285 2665 25290 2670
rect 25210 2645 25290 2665
rect 25210 2640 25215 2645
rect 25175 2635 25215 2640
rect 25285 2640 25290 2645
rect 25320 2665 25325 2670
rect 25395 2670 25435 2675
rect 25395 2665 25400 2670
rect 25320 2645 25400 2665
rect 25320 2640 25325 2645
rect 25285 2635 25325 2640
rect 25395 2640 25400 2645
rect 25430 2665 25435 2670
rect 25505 2670 25545 2675
rect 25505 2665 25510 2670
rect 25430 2645 25510 2665
rect 25430 2640 25435 2645
rect 25395 2635 25435 2640
rect 25505 2640 25510 2645
rect 25540 2665 25545 2670
rect 25615 2670 25655 2675
rect 25615 2665 25620 2670
rect 25540 2645 25620 2665
rect 25540 2640 25545 2645
rect 25505 2635 25545 2640
rect 25615 2640 25620 2645
rect 25650 2665 25655 2670
rect 25725 2670 25765 2675
rect 25725 2665 25730 2670
rect 25650 2645 25730 2665
rect 25650 2640 25655 2645
rect 25615 2635 25655 2640
rect 25725 2640 25730 2645
rect 25760 2665 25765 2670
rect 25835 2670 25875 2675
rect 25835 2665 25840 2670
rect 25760 2645 25840 2665
rect 25760 2640 25765 2645
rect 25725 2635 25765 2640
rect 25835 2640 25840 2645
rect 25870 2640 25875 2670
rect 25835 2635 25875 2640
rect 27945 2670 27985 2675
rect 27945 2640 27950 2670
rect 27980 2665 27985 2670
rect 28055 2670 28095 2675
rect 28055 2665 28060 2670
rect 27980 2645 28060 2665
rect 27980 2640 27985 2645
rect 27945 2635 27985 2640
rect 28055 2640 28060 2645
rect 28090 2665 28095 2670
rect 28165 2670 28205 2675
rect 28165 2665 28170 2670
rect 28090 2645 28170 2665
rect 28090 2640 28095 2645
rect 28055 2635 28095 2640
rect 28165 2640 28170 2645
rect 28200 2665 28205 2670
rect 28275 2670 28315 2675
rect 28275 2665 28280 2670
rect 28200 2645 28280 2665
rect 28200 2640 28205 2645
rect 28165 2635 28205 2640
rect 28275 2640 28280 2645
rect 28310 2665 28315 2670
rect 28385 2670 28425 2675
rect 28385 2665 28390 2670
rect 28310 2645 28390 2665
rect 28310 2640 28315 2645
rect 28275 2635 28315 2640
rect 28385 2640 28390 2645
rect 28420 2665 28425 2670
rect 28495 2670 28535 2675
rect 28495 2665 28500 2670
rect 28420 2645 28500 2665
rect 28420 2640 28425 2645
rect 28385 2635 28425 2640
rect 28495 2640 28500 2645
rect 28530 2665 28535 2670
rect 28605 2670 28645 2675
rect 28605 2665 28610 2670
rect 28530 2645 28610 2665
rect 28530 2640 28535 2645
rect 28495 2635 28535 2640
rect 28605 2640 28610 2645
rect 28640 2665 28645 2670
rect 28715 2670 28755 2675
rect 28715 2665 28720 2670
rect 28640 2645 28720 2665
rect 28640 2640 28645 2645
rect 28605 2635 28645 2640
rect 28715 2640 28720 2645
rect 28750 2665 28755 2670
rect 28825 2670 28865 2675
rect 28825 2665 28830 2670
rect 28750 2645 28830 2665
rect 28750 2640 28755 2645
rect 28715 2635 28755 2640
rect 28825 2640 28830 2645
rect 28860 2665 28865 2670
rect 28935 2670 28975 2675
rect 28935 2665 28940 2670
rect 28860 2645 28940 2665
rect 28860 2640 28865 2645
rect 28825 2635 28865 2640
rect 28935 2640 28940 2645
rect 28970 2665 28975 2670
rect 29045 2670 29085 2675
rect 29045 2665 29050 2670
rect 28970 2645 29050 2665
rect 28970 2640 28975 2645
rect 28935 2635 28975 2640
rect 29045 2640 29050 2645
rect 29080 2640 29085 2670
rect 29045 2635 29085 2640
rect 24790 2500 24830 2505
rect 11105 2475 11145 2480
rect 11105 2445 11110 2475
rect 11140 2470 11145 2475
rect 11823 2475 11857 2480
rect 11823 2470 11826 2475
rect 11140 2450 11826 2470
rect 11140 2445 11145 2450
rect 11105 2440 11145 2445
rect 11823 2445 11826 2450
rect 11854 2445 11857 2475
rect 24790 2470 24795 2500
rect 24825 2495 24830 2500
rect 24900 2500 24940 2505
rect 24900 2495 24905 2500
rect 24825 2475 24905 2495
rect 24825 2470 24830 2475
rect 24790 2465 24830 2470
rect 24900 2470 24905 2475
rect 24935 2495 24940 2500
rect 25010 2500 25050 2505
rect 25010 2495 25015 2500
rect 24935 2475 25015 2495
rect 24935 2470 24940 2475
rect 24900 2465 24940 2470
rect 25010 2470 25015 2475
rect 25045 2495 25050 2500
rect 25120 2500 25160 2505
rect 25120 2495 25125 2500
rect 25045 2475 25125 2495
rect 25045 2470 25050 2475
rect 25010 2465 25050 2470
rect 25120 2470 25125 2475
rect 25155 2495 25160 2500
rect 25230 2500 25270 2505
rect 25230 2495 25235 2500
rect 25155 2475 25235 2495
rect 25155 2470 25160 2475
rect 25120 2465 25160 2470
rect 25230 2470 25235 2475
rect 25265 2495 25270 2500
rect 25340 2500 25380 2505
rect 25340 2495 25345 2500
rect 25265 2475 25345 2495
rect 25265 2470 25270 2475
rect 25230 2465 25270 2470
rect 25340 2470 25345 2475
rect 25375 2495 25380 2500
rect 25450 2500 25490 2505
rect 25450 2495 25455 2500
rect 25375 2475 25455 2495
rect 25375 2470 25380 2475
rect 25340 2465 25380 2470
rect 25450 2470 25455 2475
rect 25485 2495 25490 2500
rect 25560 2500 25600 2505
rect 25560 2495 25565 2500
rect 25485 2475 25565 2495
rect 25485 2470 25490 2475
rect 25450 2465 25490 2470
rect 25560 2470 25565 2475
rect 25595 2495 25600 2500
rect 25670 2500 25710 2505
rect 25670 2495 25675 2500
rect 25595 2475 25675 2495
rect 25595 2470 25600 2475
rect 25560 2465 25600 2470
rect 25670 2470 25675 2475
rect 25705 2495 25710 2500
rect 25780 2500 25820 2505
rect 25780 2495 25785 2500
rect 25705 2475 25785 2495
rect 25705 2470 25710 2475
rect 25670 2465 25710 2470
rect 25780 2470 25785 2475
rect 25815 2470 25820 2500
rect 28000 2500 28040 2505
rect 25780 2465 25820 2470
rect 25980 2475 26020 2480
rect 25980 2445 25985 2475
rect 26015 2470 26020 2475
rect 26823 2475 26857 2480
rect 26823 2470 26826 2475
rect 26015 2450 26826 2470
rect 26015 2445 26020 2450
rect 11823 2440 11857 2445
rect 25813 2440 25847 2445
rect 25980 2440 26020 2445
rect 26823 2445 26826 2450
rect 26854 2445 26857 2475
rect 28000 2470 28005 2500
rect 28035 2495 28040 2500
rect 28110 2500 28150 2505
rect 28110 2495 28115 2500
rect 28035 2475 28115 2495
rect 28035 2470 28040 2475
rect 28000 2465 28040 2470
rect 28110 2470 28115 2475
rect 28145 2495 28150 2500
rect 28220 2500 28260 2505
rect 28220 2495 28225 2500
rect 28145 2475 28225 2495
rect 28145 2470 28150 2475
rect 28110 2465 28150 2470
rect 28220 2470 28225 2475
rect 28255 2495 28260 2500
rect 28330 2500 28370 2505
rect 28330 2495 28335 2500
rect 28255 2475 28335 2495
rect 28255 2470 28260 2475
rect 28220 2465 28260 2470
rect 28330 2470 28335 2475
rect 28365 2495 28370 2500
rect 28440 2500 28480 2505
rect 28440 2495 28445 2500
rect 28365 2475 28445 2495
rect 28365 2470 28370 2475
rect 28330 2465 28370 2470
rect 28440 2470 28445 2475
rect 28475 2495 28480 2500
rect 28550 2500 28590 2505
rect 28550 2495 28555 2500
rect 28475 2475 28555 2495
rect 28475 2470 28480 2475
rect 28440 2465 28480 2470
rect 28550 2470 28555 2475
rect 28585 2495 28590 2500
rect 28660 2500 28700 2505
rect 28660 2495 28665 2500
rect 28585 2475 28665 2495
rect 28585 2470 28590 2475
rect 28550 2465 28590 2470
rect 28660 2470 28665 2475
rect 28695 2495 28700 2500
rect 28770 2500 28810 2505
rect 28770 2495 28775 2500
rect 28695 2475 28775 2495
rect 28695 2470 28700 2475
rect 28660 2465 28700 2470
rect 28770 2470 28775 2475
rect 28805 2495 28810 2500
rect 28880 2500 28920 2505
rect 28880 2495 28885 2500
rect 28805 2475 28885 2495
rect 28805 2470 28810 2475
rect 28770 2465 28810 2470
rect 28880 2470 28885 2475
rect 28915 2495 28920 2500
rect 28990 2500 29030 2505
rect 28990 2495 28995 2500
rect 28915 2475 28995 2495
rect 28915 2470 28920 2475
rect 28880 2465 28920 2470
rect 28990 2470 28995 2475
rect 29025 2470 29030 2500
rect 28990 2465 29030 2470
rect 26823 2440 26857 2445
rect 27973 2440 28007 2445
rect 10020 2435 10060 2440
rect 10020 2405 10025 2435
rect 10055 2430 10060 2435
rect 10265 2435 10305 2440
rect 10265 2430 10270 2435
rect 10055 2410 10270 2430
rect 10055 2405 10060 2410
rect 10020 2400 10060 2405
rect 10265 2405 10270 2410
rect 10300 2430 10305 2435
rect 10375 2435 10415 2440
rect 10375 2430 10380 2435
rect 10300 2410 10380 2430
rect 10300 2405 10305 2410
rect 10265 2400 10305 2405
rect 10375 2405 10380 2410
rect 10410 2430 10415 2435
rect 10485 2435 10525 2440
rect 10485 2430 10490 2435
rect 10410 2410 10490 2430
rect 10410 2405 10415 2410
rect 10375 2400 10415 2405
rect 10485 2405 10490 2410
rect 10520 2430 10525 2435
rect 10595 2435 10635 2440
rect 10595 2430 10600 2435
rect 10520 2410 10600 2430
rect 10520 2405 10525 2410
rect 10485 2400 10525 2405
rect 10595 2405 10600 2410
rect 10630 2430 10635 2435
rect 10705 2435 10745 2440
rect 10705 2430 10710 2435
rect 10630 2410 10710 2430
rect 10630 2405 10635 2410
rect 10595 2400 10635 2405
rect 10705 2405 10710 2410
rect 10740 2405 10745 2435
rect 13055 2435 13095 2440
rect 11000 2420 11040 2425
rect 11000 2415 11005 2420
rect 10705 2400 10745 2405
rect 10785 2395 11005 2415
rect 10765 2390 10805 2395
rect 3805 2380 3845 2385
rect 3355 2375 3395 2380
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2340 2660 2345
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3805 2350 3810 2380
rect 3840 2375 3845 2380
rect 4165 2380 4205 2385
rect 4165 2375 4170 2380
rect 3840 2355 4170 2375
rect 3840 2350 3845 2355
rect 3805 2345 3845 2350
rect 4165 2350 4170 2355
rect 4200 2350 4205 2380
rect 10765 2360 10770 2390
rect 10800 2360 10805 2390
rect 11000 2390 11005 2395
rect 11035 2415 11040 2420
rect 11280 2420 11320 2425
rect 11280 2415 11285 2420
rect 11035 2395 11285 2415
rect 11035 2390 11040 2395
rect 11000 2385 11040 2390
rect 11280 2390 11285 2395
rect 11315 2415 11320 2420
rect 11520 2420 11560 2425
rect 11520 2415 11525 2420
rect 11315 2395 11525 2415
rect 11315 2390 11320 2395
rect 11280 2385 11320 2390
rect 11520 2390 11525 2395
rect 11555 2415 11560 2420
rect 11760 2420 11800 2425
rect 11760 2415 11765 2420
rect 11555 2395 11765 2415
rect 11555 2390 11560 2395
rect 11520 2385 11560 2390
rect 11760 2390 11765 2395
rect 11795 2415 11800 2420
rect 12000 2420 12040 2425
rect 12000 2415 12005 2420
rect 11795 2395 12005 2415
rect 11795 2390 11800 2395
rect 11760 2385 11800 2390
rect 12000 2390 12005 2395
rect 12035 2415 12040 2420
rect 12240 2420 12280 2425
rect 12240 2415 12245 2420
rect 12035 2395 12245 2415
rect 12035 2390 12040 2395
rect 12000 2385 12040 2390
rect 12240 2390 12245 2395
rect 12275 2415 12280 2420
rect 12480 2420 12520 2425
rect 12480 2415 12485 2420
rect 12275 2395 12485 2415
rect 12275 2390 12280 2395
rect 12240 2385 12280 2390
rect 12480 2390 12485 2395
rect 12515 2390 12520 2420
rect 13055 2405 13060 2435
rect 13090 2430 13095 2435
rect 13165 2435 13205 2440
rect 13165 2430 13170 2435
rect 13090 2410 13170 2430
rect 13090 2405 13095 2410
rect 13055 2400 13095 2405
rect 13165 2405 13170 2410
rect 13200 2430 13205 2435
rect 13275 2435 13315 2440
rect 13275 2430 13280 2435
rect 13200 2410 13280 2430
rect 13200 2405 13205 2410
rect 13165 2400 13205 2405
rect 13275 2405 13280 2410
rect 13310 2430 13315 2435
rect 13385 2435 13425 2440
rect 13385 2430 13390 2435
rect 13310 2410 13390 2430
rect 13310 2405 13315 2410
rect 13275 2400 13315 2405
rect 13385 2405 13390 2410
rect 13420 2430 13425 2435
rect 13495 2435 13535 2440
rect 13495 2430 13500 2435
rect 13420 2410 13500 2430
rect 13420 2405 13425 2410
rect 13385 2400 13425 2405
rect 13495 2405 13500 2410
rect 13530 2430 13535 2435
rect 13740 2435 13780 2440
rect 13740 2430 13745 2435
rect 13530 2410 13745 2430
rect 13530 2405 13535 2410
rect 13495 2400 13535 2405
rect 13740 2405 13745 2410
rect 13775 2405 13780 2435
rect 25813 2410 25816 2440
rect 25844 2425 25847 2440
rect 25844 2420 26320 2425
rect 25844 2410 26285 2420
rect 25813 2405 26285 2410
rect 13740 2400 13780 2405
rect 12480 2385 12520 2390
rect 26280 2390 26285 2405
rect 26315 2415 26320 2420
rect 26520 2420 26560 2425
rect 26520 2415 26525 2420
rect 26315 2395 26525 2415
rect 26315 2390 26320 2395
rect 26280 2385 26320 2390
rect 26520 2390 26525 2395
rect 26555 2415 26560 2420
rect 26760 2420 26800 2425
rect 26760 2415 26765 2420
rect 26555 2395 26765 2415
rect 26555 2390 26560 2395
rect 26520 2385 26560 2390
rect 26760 2390 26765 2395
rect 26795 2415 26800 2420
rect 27000 2420 27040 2425
rect 27000 2415 27005 2420
rect 26795 2395 27005 2415
rect 26795 2390 26800 2395
rect 26760 2385 26800 2390
rect 27000 2390 27005 2395
rect 27035 2415 27040 2420
rect 27240 2420 27280 2425
rect 27240 2415 27245 2420
rect 27035 2395 27245 2415
rect 27035 2390 27040 2395
rect 27000 2385 27040 2390
rect 27240 2390 27245 2395
rect 27275 2415 27280 2420
rect 27480 2420 27520 2425
rect 27480 2415 27485 2420
rect 27275 2395 27485 2415
rect 27275 2390 27280 2395
rect 27240 2385 27280 2390
rect 27480 2390 27485 2395
rect 27515 2390 27520 2420
rect 27973 2410 27976 2440
rect 28004 2410 28007 2440
rect 27973 2405 28007 2410
rect 27480 2385 27520 2390
rect 10765 2355 10805 2360
rect 11400 2375 11440 2380
rect 4165 2345 4205 2350
rect 11400 2345 11405 2375
rect 11435 2370 11440 2375
rect 11640 2375 11680 2380
rect 11640 2370 11645 2375
rect 11435 2350 11645 2370
rect 11435 2345 11440 2350
rect 3355 2340 3395 2345
rect 11400 2340 11440 2345
rect 11640 2345 11645 2350
rect 11675 2370 11680 2375
rect 11880 2375 11920 2380
rect 11880 2370 11885 2375
rect 11675 2350 11885 2370
rect 11675 2345 11680 2350
rect 11640 2340 11680 2345
rect 11880 2345 11885 2350
rect 11915 2370 11920 2375
rect 12120 2375 12160 2380
rect 12120 2370 12125 2375
rect 11915 2350 12125 2370
rect 11915 2345 11920 2350
rect 11880 2340 11920 2345
rect 12120 2345 12125 2350
rect 12155 2370 12160 2375
rect 12360 2375 12400 2380
rect 12360 2370 12365 2375
rect 12155 2350 12365 2370
rect 12155 2345 12160 2350
rect 12120 2340 12160 2345
rect 12360 2345 12365 2350
rect 12395 2370 12400 2375
rect 12690 2375 12730 2380
rect 12690 2370 12695 2375
rect 12395 2350 12695 2370
rect 12395 2345 12400 2350
rect 12360 2340 12400 2345
rect 12690 2345 12695 2350
rect 12725 2370 12730 2375
rect 13025 2375 13065 2380
rect 13025 2370 13030 2375
rect 12725 2350 13030 2370
rect 12725 2345 12730 2350
rect 12690 2340 12730 2345
rect 13025 2345 13030 2350
rect 13060 2345 13065 2375
rect 24800 2345 24805 2380
rect 24840 2345 24845 2380
rect 25635 2345 25640 2380
rect 25675 2345 25680 2380
rect 26400 2375 26440 2380
rect 26400 2345 26405 2375
rect 26435 2370 26440 2375
rect 26640 2375 26680 2380
rect 26640 2370 26645 2375
rect 26435 2350 26645 2370
rect 26435 2345 26440 2350
rect 13025 2340 13065 2345
rect 26400 2340 26440 2345
rect 26640 2345 26645 2350
rect 26675 2370 26680 2375
rect 26880 2375 26920 2380
rect 26880 2370 26885 2375
rect 26675 2350 26885 2370
rect 26675 2345 26680 2350
rect 26640 2340 26680 2345
rect 26880 2345 26885 2350
rect 26915 2370 26920 2375
rect 27120 2375 27160 2380
rect 27120 2370 27125 2375
rect 26915 2350 27125 2370
rect 26915 2345 26920 2350
rect 26880 2340 26920 2345
rect 27120 2345 27125 2350
rect 27155 2370 27160 2375
rect 27360 2375 27400 2380
rect 27360 2370 27365 2375
rect 27155 2350 27365 2370
rect 27155 2345 27160 2350
rect 27120 2340 27160 2345
rect 27360 2345 27365 2350
rect 27395 2370 27400 2375
rect 27690 2375 27730 2380
rect 27690 2370 27695 2375
rect 27395 2350 27695 2370
rect 27395 2345 27400 2350
rect 27360 2340 27400 2345
rect 27690 2345 27695 2350
rect 27725 2370 27730 2375
rect 27970 2375 28010 2380
rect 27970 2370 27975 2375
rect 27725 2350 27975 2370
rect 27725 2345 27730 2350
rect 27690 2340 27730 2345
rect 27970 2345 27975 2350
rect 28005 2345 28010 2375
rect 28140 2345 28145 2380
rect 28180 2345 28185 2380
rect 28974 2345 28980 2380
rect 29015 2345 29020 2380
rect 27970 2340 28010 2345
rect 2655 2320 3395 2340
rect 3625 2335 3665 2340
rect 2655 2315 2660 2320
rect 2620 2310 2660 2315
rect 3625 2305 3630 2335
rect 3660 2330 3665 2335
rect 4345 2335 4385 2340
rect 4345 2330 4350 2335
rect 3660 2310 4350 2330
rect 3660 2305 3665 2310
rect 3625 2300 3665 2305
rect 4345 2305 4350 2310
rect 4380 2305 4385 2335
rect 11000 2325 11040 2330
rect 4345 2300 4385 2305
rect 10065 2315 10105 2320
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2285 2775 2290
rect 3445 2290 3485 2295
rect 3445 2285 3450 2290
rect 2770 2265 3450 2285
rect 2770 2260 2775 2265
rect 2735 2255 2775 2260
rect 3445 2260 3450 2265
rect 3480 2285 3485 2290
rect 4525 2290 4565 2295
rect 4525 2285 4530 2290
rect 3480 2265 4530 2285
rect 3480 2260 3485 2265
rect 3445 2255 3485 2260
rect 4525 2260 4530 2265
rect 4560 2285 4565 2290
rect 5270 2290 5310 2295
rect 5270 2285 5275 2290
rect 4560 2265 5275 2285
rect 4560 2260 4565 2265
rect 4525 2255 4565 2260
rect 5270 2260 5275 2265
rect 5305 2260 5310 2290
rect 10065 2285 10070 2315
rect 10100 2310 10105 2315
rect 10265 2315 10305 2320
rect 10265 2310 10270 2315
rect 10100 2290 10270 2310
rect 10100 2285 10105 2290
rect 10065 2280 10105 2285
rect 10265 2285 10270 2290
rect 10300 2310 10305 2315
rect 10375 2315 10415 2320
rect 10375 2310 10380 2315
rect 10300 2290 10380 2310
rect 10300 2285 10305 2290
rect 10265 2280 10305 2285
rect 10375 2285 10380 2290
rect 10410 2310 10415 2315
rect 10485 2315 10525 2320
rect 10485 2310 10490 2315
rect 10410 2290 10490 2310
rect 10410 2285 10415 2290
rect 10375 2280 10415 2285
rect 10485 2285 10490 2290
rect 10520 2310 10525 2315
rect 10595 2315 10635 2320
rect 10595 2310 10600 2315
rect 10520 2290 10600 2310
rect 10520 2285 10525 2290
rect 10485 2280 10525 2285
rect 10595 2285 10600 2290
rect 10630 2310 10635 2315
rect 10705 2315 10745 2320
rect 10705 2310 10710 2315
rect 10630 2290 10710 2310
rect 10630 2285 10635 2290
rect 10595 2280 10635 2285
rect 10705 2285 10710 2290
rect 10740 2285 10745 2315
rect 11000 2295 11005 2325
rect 11035 2320 11040 2325
rect 12760 2325 12800 2330
rect 12760 2320 12765 2325
rect 11035 2300 12765 2320
rect 11035 2295 11040 2300
rect 11000 2290 11040 2295
rect 12760 2295 12765 2300
rect 12795 2295 12800 2325
rect 27815 2325 27855 2330
rect 27815 2320 27820 2325
rect 12760 2290 12800 2295
rect 13055 2315 13095 2320
rect 13055 2285 13060 2315
rect 13090 2310 13095 2315
rect 13165 2315 13205 2320
rect 13165 2310 13170 2315
rect 13090 2290 13170 2310
rect 13090 2285 13095 2290
rect 10705 2280 10745 2285
rect 11440 2280 11480 2285
rect 5270 2255 5310 2260
rect 11440 2250 11445 2280
rect 11475 2275 11480 2280
rect 11660 2280 11700 2285
rect 11660 2275 11665 2280
rect 11475 2255 11665 2275
rect 11475 2250 11480 2255
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3805 2245 3845 2250
rect 11440 2245 11480 2250
rect 11660 2250 11665 2255
rect 11695 2275 11700 2280
rect 11880 2280 11920 2285
rect 11880 2275 11885 2280
rect 11695 2255 11885 2275
rect 11695 2250 11700 2255
rect 11660 2245 11700 2250
rect 11880 2250 11885 2255
rect 11915 2275 11920 2280
rect 12100 2280 12140 2285
rect 12100 2275 12105 2280
rect 11915 2255 12105 2275
rect 11915 2250 11920 2255
rect 11880 2245 11920 2250
rect 12100 2250 12105 2255
rect 12135 2275 12140 2280
rect 12320 2280 12360 2285
rect 13055 2280 13095 2285
rect 13165 2285 13170 2290
rect 13200 2310 13205 2315
rect 13275 2315 13315 2320
rect 13275 2310 13280 2315
rect 13200 2290 13280 2310
rect 13200 2285 13205 2290
rect 13165 2280 13205 2285
rect 13275 2285 13280 2290
rect 13310 2310 13315 2315
rect 13385 2315 13425 2320
rect 13385 2310 13390 2315
rect 13310 2290 13390 2310
rect 13310 2285 13315 2290
rect 13275 2280 13315 2285
rect 13385 2285 13390 2290
rect 13420 2310 13425 2315
rect 13495 2315 13535 2320
rect 13495 2310 13500 2315
rect 13420 2290 13500 2310
rect 13420 2285 13425 2290
rect 13385 2280 13425 2285
rect 13495 2285 13500 2290
rect 13530 2310 13535 2315
rect 13695 2315 13735 2320
rect 13695 2310 13700 2315
rect 13530 2290 13700 2310
rect 13530 2285 13535 2290
rect 13495 2280 13535 2285
rect 13695 2285 13700 2290
rect 13730 2285 13735 2315
rect 24800 2285 24805 2320
rect 24840 2285 24845 2320
rect 25635 2285 25640 2320
rect 25675 2300 27820 2320
rect 25675 2285 25680 2300
rect 27815 2295 27820 2300
rect 27850 2320 27855 2325
rect 27850 2300 28145 2320
rect 27850 2295 27855 2300
rect 27815 2290 27855 2295
rect 28140 2285 28145 2300
rect 28180 2285 28185 2320
rect 28975 2285 28980 2320
rect 29015 2285 29020 2320
rect 13695 2280 13735 2285
rect 25813 2280 25847 2285
rect 12320 2275 12325 2280
rect 12135 2255 12325 2275
rect 12135 2250 12140 2255
rect 12100 2245 12140 2250
rect 12320 2250 12325 2255
rect 12355 2250 12360 2280
rect 12320 2245 12360 2250
rect 25813 2250 25816 2280
rect 25844 2250 25847 2280
rect 25813 2245 25847 2250
rect 26440 2280 26480 2285
rect 26440 2250 26445 2280
rect 26475 2275 26480 2280
rect 26660 2280 26700 2285
rect 26660 2275 26665 2280
rect 26475 2255 26665 2275
rect 26475 2250 26480 2255
rect 26440 2245 26480 2250
rect 26660 2250 26665 2255
rect 26695 2275 26700 2280
rect 26880 2280 26920 2285
rect 26880 2275 26885 2280
rect 26695 2255 26885 2275
rect 26695 2250 26700 2255
rect 26660 2245 26700 2250
rect 26880 2250 26885 2255
rect 26915 2275 26920 2280
rect 27100 2280 27140 2285
rect 27100 2275 27105 2280
rect 26915 2255 27105 2275
rect 26915 2250 26920 2255
rect 26880 2245 26920 2250
rect 27100 2250 27105 2255
rect 27135 2275 27140 2280
rect 27320 2280 27360 2285
rect 27320 2275 27325 2280
rect 27135 2255 27325 2275
rect 27135 2250 27140 2255
rect 27100 2245 27140 2250
rect 27320 2250 27325 2255
rect 27355 2250 27360 2280
rect 27320 2245 27360 2250
rect 27973 2280 28007 2285
rect 27973 2250 27976 2280
rect 28004 2250 28007 2280
rect 27973 2245 28007 2250
rect 3805 2240 3810 2245
rect 2460 2220 3810 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3805 2215 3810 2220
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 11330 2235 11370 2240
rect 11330 2205 11335 2235
rect 11365 2230 11370 2235
rect 11550 2235 11590 2240
rect 11550 2230 11555 2235
rect 11365 2210 11555 2230
rect 11365 2205 11370 2210
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 3265 2200 3305 2205
rect 3265 2195 3270 2200
rect 2365 2175 3270 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 3265 2170 3270 2175
rect 3300 2195 3305 2200
rect 3985 2200 4025 2205
rect 3985 2195 3990 2200
rect 3300 2175 3990 2195
rect 3300 2170 3305 2175
rect 3265 2165 3305 2170
rect 3985 2170 3990 2175
rect 4020 2195 4025 2200
rect 4705 2200 4745 2205
rect 11330 2200 11370 2205
rect 11550 2205 11555 2210
rect 11585 2230 11590 2235
rect 11770 2235 11810 2240
rect 11770 2230 11775 2235
rect 11585 2210 11775 2230
rect 11585 2205 11590 2210
rect 11550 2200 11590 2205
rect 11770 2205 11775 2210
rect 11805 2230 11810 2235
rect 11990 2235 12030 2240
rect 11990 2230 11995 2235
rect 11805 2210 11995 2230
rect 11805 2205 11810 2210
rect 11770 2200 11810 2205
rect 11990 2205 11995 2210
rect 12025 2230 12030 2235
rect 12210 2235 12250 2240
rect 12210 2230 12215 2235
rect 12025 2210 12215 2230
rect 12025 2205 12030 2210
rect 11990 2200 12030 2205
rect 12210 2205 12215 2210
rect 12245 2230 12250 2235
rect 12430 2235 12470 2240
rect 12430 2230 12435 2235
rect 12245 2210 12435 2230
rect 12245 2205 12250 2210
rect 12210 2200 12250 2205
rect 12430 2205 12435 2210
rect 12465 2205 12470 2235
rect 26330 2235 26370 2240
rect 12430 2200 12470 2205
rect 24790 2220 24830 2225
rect 4705 2195 4710 2200
rect 4020 2175 4710 2195
rect 4020 2170 4025 2175
rect 3985 2165 4025 2170
rect 4705 2170 4710 2175
rect 4740 2170 4745 2200
rect 24790 2190 24795 2220
rect 24825 2215 24830 2220
rect 24900 2220 24940 2225
rect 24900 2215 24905 2220
rect 24825 2195 24905 2215
rect 24825 2190 24830 2195
rect 24790 2185 24830 2190
rect 24900 2190 24905 2195
rect 24935 2215 24940 2220
rect 25010 2220 25050 2225
rect 25010 2215 25015 2220
rect 24935 2195 25015 2215
rect 24935 2190 24940 2195
rect 24900 2185 24940 2190
rect 25010 2190 25015 2195
rect 25045 2215 25050 2220
rect 25120 2220 25160 2225
rect 25120 2215 25125 2220
rect 25045 2195 25125 2215
rect 25045 2190 25050 2195
rect 25010 2185 25050 2190
rect 25120 2190 25125 2195
rect 25155 2215 25160 2220
rect 25230 2220 25270 2225
rect 25230 2215 25235 2220
rect 25155 2195 25235 2215
rect 25155 2190 25160 2195
rect 25120 2185 25160 2190
rect 25230 2190 25235 2195
rect 25265 2215 25270 2220
rect 25340 2220 25380 2225
rect 25340 2215 25345 2220
rect 25265 2195 25345 2215
rect 25265 2190 25270 2195
rect 25230 2185 25270 2190
rect 25340 2190 25345 2195
rect 25375 2215 25380 2220
rect 25450 2220 25490 2225
rect 25450 2215 25455 2220
rect 25375 2195 25455 2215
rect 25375 2190 25380 2195
rect 25340 2185 25380 2190
rect 25450 2190 25455 2195
rect 25485 2215 25490 2220
rect 25560 2220 25600 2225
rect 25560 2215 25565 2220
rect 25485 2195 25565 2215
rect 25485 2190 25490 2195
rect 25450 2185 25490 2190
rect 25560 2190 25565 2195
rect 25595 2215 25600 2220
rect 25670 2220 25710 2225
rect 25670 2215 25675 2220
rect 25595 2195 25675 2215
rect 25595 2190 25600 2195
rect 25560 2185 25600 2190
rect 25670 2190 25675 2195
rect 25705 2215 25710 2220
rect 25780 2220 25820 2225
rect 25780 2215 25785 2220
rect 25705 2195 25785 2215
rect 25705 2190 25710 2195
rect 25670 2185 25710 2190
rect 25780 2190 25785 2195
rect 25815 2190 25820 2220
rect 26330 2205 26335 2235
rect 26365 2230 26370 2235
rect 26550 2235 26590 2240
rect 26550 2230 26555 2235
rect 26365 2210 26555 2230
rect 26365 2205 26370 2210
rect 26330 2200 26370 2205
rect 26550 2205 26555 2210
rect 26585 2230 26590 2235
rect 26770 2235 26810 2240
rect 26770 2230 26775 2235
rect 26585 2210 26775 2230
rect 26585 2205 26590 2210
rect 26550 2200 26590 2205
rect 26770 2205 26775 2210
rect 26805 2230 26810 2235
rect 26990 2235 27030 2240
rect 26990 2230 26995 2235
rect 26805 2210 26995 2230
rect 26805 2205 26810 2210
rect 26770 2200 26810 2205
rect 26990 2205 26995 2210
rect 27025 2230 27030 2235
rect 27210 2235 27250 2240
rect 27210 2230 27215 2235
rect 27025 2210 27215 2230
rect 27025 2205 27030 2210
rect 26990 2200 27030 2205
rect 27210 2205 27215 2210
rect 27245 2230 27250 2235
rect 27430 2235 27470 2240
rect 27430 2230 27435 2235
rect 27245 2210 27435 2230
rect 27245 2205 27250 2210
rect 27210 2200 27250 2205
rect 27430 2205 27435 2210
rect 27465 2205 27470 2235
rect 27430 2200 27470 2205
rect 28000 2220 28040 2225
rect 25780 2185 25820 2190
rect 28000 2190 28005 2220
rect 28035 2215 28040 2220
rect 28110 2220 28150 2225
rect 28110 2215 28115 2220
rect 28035 2195 28115 2215
rect 28035 2190 28040 2195
rect 28000 2185 28040 2190
rect 28110 2190 28115 2195
rect 28145 2215 28150 2220
rect 28220 2220 28260 2225
rect 28220 2215 28225 2220
rect 28145 2195 28225 2215
rect 28145 2190 28150 2195
rect 28110 2185 28150 2190
rect 28220 2190 28225 2195
rect 28255 2215 28260 2220
rect 28330 2220 28370 2225
rect 28330 2215 28335 2220
rect 28255 2195 28335 2215
rect 28255 2190 28260 2195
rect 28220 2185 28260 2190
rect 28330 2190 28335 2195
rect 28365 2215 28370 2220
rect 28440 2220 28480 2225
rect 28440 2215 28445 2220
rect 28365 2195 28445 2215
rect 28365 2190 28370 2195
rect 28330 2185 28370 2190
rect 28440 2190 28445 2195
rect 28475 2215 28480 2220
rect 28550 2220 28590 2225
rect 28550 2215 28555 2220
rect 28475 2195 28555 2215
rect 28475 2190 28480 2195
rect 28440 2185 28480 2190
rect 28550 2190 28555 2195
rect 28585 2215 28590 2220
rect 28660 2220 28700 2225
rect 28660 2215 28665 2220
rect 28585 2195 28665 2215
rect 28585 2190 28590 2195
rect 28550 2185 28590 2190
rect 28660 2190 28665 2195
rect 28695 2215 28700 2220
rect 28770 2220 28810 2225
rect 28770 2215 28775 2220
rect 28695 2195 28775 2215
rect 28695 2190 28700 2195
rect 28660 2185 28700 2190
rect 28770 2190 28775 2195
rect 28805 2215 28810 2220
rect 28880 2220 28920 2225
rect 28880 2215 28885 2220
rect 28805 2195 28885 2215
rect 28805 2190 28810 2195
rect 28770 2185 28810 2190
rect 28880 2190 28885 2195
rect 28915 2215 28920 2220
rect 28990 2220 29030 2225
rect 28990 2215 28995 2220
rect 28915 2195 28995 2215
rect 28915 2190 28920 2195
rect 28880 2185 28920 2190
rect 28990 2190 28995 2195
rect 29025 2190 29030 2220
rect 28990 2185 29030 2190
rect 4705 2165 4745 2170
rect 10950 2180 10990 2185
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3625 2150 3665 2155
rect 10950 2150 10955 2180
rect 10985 2175 10990 2180
rect 11828 2180 11862 2185
rect 11828 2175 11831 2180
rect 10985 2155 11831 2175
rect 10985 2150 10990 2155
rect 3625 2145 3630 2150
rect 2415 2125 3630 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3625 2120 3630 2125
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2140 4125 2145
rect 5315 2145 5355 2150
rect 10950 2145 10990 2150
rect 11828 2150 11831 2155
rect 11859 2150 11862 2180
rect 11828 2145 11862 2150
rect 5315 2140 5320 2145
rect 4120 2120 5320 2140
rect 4120 2115 4125 2120
rect 4085 2110 4125 2115
rect 5315 2115 5320 2120
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2090 2785 2095
rect 2865 2095 2905 2100
rect 2865 2090 2870 2095
rect 2780 2070 2870 2090
rect 2780 2065 2785 2070
rect 2745 2060 2785 2065
rect 2865 2065 2870 2070
rect 2900 2090 2905 2095
rect 2985 2095 3025 2100
rect 2985 2090 2990 2095
rect 2900 2070 2990 2090
rect 2900 2065 2905 2070
rect 2865 2060 2905 2065
rect 2985 2065 2990 2070
rect 3020 2090 3025 2095
rect 3105 2095 3145 2100
rect 3105 2090 3110 2095
rect 3020 2070 3110 2090
rect 3020 2065 3025 2070
rect 2985 2060 3025 2065
rect 3105 2065 3110 2070
rect 3140 2090 3145 2095
rect 3225 2095 3265 2100
rect 3225 2090 3230 2095
rect 3140 2070 3230 2090
rect 3140 2065 3145 2070
rect 3105 2060 3145 2065
rect 3225 2065 3230 2070
rect 3260 2090 3265 2095
rect 3345 2095 3385 2100
rect 3345 2090 3350 2095
rect 3260 2070 3350 2090
rect 3260 2065 3265 2070
rect 3225 2060 3265 2065
rect 3345 2065 3350 2070
rect 3380 2090 3385 2095
rect 3465 2095 3505 2100
rect 3465 2090 3470 2095
rect 3380 2070 3470 2090
rect 3380 2065 3385 2070
rect 3345 2060 3385 2065
rect 3465 2065 3470 2070
rect 3500 2090 3505 2095
rect 3585 2095 3625 2100
rect 3585 2090 3590 2095
rect 3500 2070 3590 2090
rect 3500 2065 3505 2070
rect 3465 2060 3505 2065
rect 3585 2065 3590 2070
rect 3620 2090 3625 2095
rect 3705 2095 3745 2100
rect 3705 2090 3710 2095
rect 3620 2070 3710 2090
rect 3620 2065 3625 2070
rect 3585 2060 3625 2065
rect 3705 2065 3710 2070
rect 3740 2090 3745 2095
rect 3825 2095 3865 2100
rect 3825 2090 3830 2095
rect 3740 2070 3830 2090
rect 3740 2065 3745 2070
rect 3705 2060 3745 2065
rect 3825 2065 3830 2070
rect 3860 2090 3865 2095
rect 3985 2095 4025 2100
rect 3985 2090 3990 2095
rect 3860 2070 3990 2090
rect 3860 2065 3865 2070
rect 3825 2060 3865 2065
rect 3985 2065 3990 2070
rect 4020 2090 4025 2095
rect 4145 2095 4185 2100
rect 4145 2090 4150 2095
rect 4020 2070 4150 2090
rect 4020 2065 4025 2070
rect 3985 2060 4025 2065
rect 4145 2065 4150 2070
rect 4180 2090 4185 2095
rect 4265 2095 4305 2100
rect 4265 2090 4270 2095
rect 4180 2070 4270 2090
rect 4180 2065 4185 2070
rect 4145 2060 4185 2065
rect 4265 2065 4270 2070
rect 4300 2090 4305 2095
rect 4385 2095 4425 2100
rect 4385 2090 4390 2095
rect 4300 2070 4390 2090
rect 4300 2065 4305 2070
rect 4265 2060 4305 2065
rect 4385 2065 4390 2070
rect 4420 2090 4425 2095
rect 4505 2095 4545 2100
rect 4505 2090 4510 2095
rect 4420 2070 4510 2090
rect 4420 2065 4425 2070
rect 4385 2060 4425 2065
rect 4505 2065 4510 2070
rect 4540 2090 4545 2095
rect 4625 2095 4665 2100
rect 4625 2090 4630 2095
rect 4540 2070 4630 2090
rect 4540 2065 4545 2070
rect 4505 2060 4545 2065
rect 4625 2065 4630 2070
rect 4660 2090 4665 2095
rect 4745 2095 4785 2100
rect 4745 2090 4750 2095
rect 4660 2070 4750 2090
rect 4660 2065 4665 2070
rect 4625 2060 4665 2065
rect 4745 2065 4750 2070
rect 4780 2090 4785 2095
rect 4865 2095 4905 2100
rect 4865 2090 4870 2095
rect 4780 2070 4870 2090
rect 4780 2065 4785 2070
rect 4745 2060 4785 2065
rect 4865 2065 4870 2070
rect 4900 2090 4905 2095
rect 4985 2095 5025 2100
rect 4985 2090 4990 2095
rect 4900 2070 4990 2090
rect 4900 2065 4905 2070
rect 4865 2060 4905 2065
rect 4985 2065 4990 2070
rect 5020 2090 5025 2095
rect 5105 2095 5145 2100
rect 5105 2090 5110 2095
rect 5020 2070 5110 2090
rect 5020 2065 5025 2070
rect 4985 2060 5025 2065
rect 5105 2065 5110 2070
rect 5140 2090 5145 2095
rect 5225 2095 5265 2100
rect 5225 2090 5230 2095
rect 5140 2070 5230 2090
rect 5140 2065 5145 2070
rect 5105 2060 5145 2065
rect 5225 2065 5230 2070
rect 5260 2090 5265 2095
rect 5550 2095 5590 2100
rect 5550 2090 5555 2095
rect 5260 2070 5555 2090
rect 5260 2065 5265 2070
rect 5225 2060 5265 2065
rect 5550 2065 5555 2070
rect 5585 2065 5590 2095
rect 5550 2060 5590 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2045 2845 2050
rect 3165 2050 3205 2055
rect 3165 2045 3170 2050
rect 2840 2025 3170 2045
rect 2840 2020 2845 2025
rect 2805 2015 2845 2020
rect 3165 2020 3170 2025
rect 3200 2045 3205 2050
rect 3525 2050 3565 2055
rect 3525 2045 3530 2050
rect 3200 2025 3530 2045
rect 3200 2020 3205 2025
rect 3165 2015 3205 2020
rect 3525 2020 3530 2025
rect 3560 2045 3565 2050
rect 3885 2050 3925 2055
rect 3885 2045 3890 2050
rect 3560 2025 3890 2045
rect 3560 2020 3565 2025
rect 3525 2015 3565 2020
rect 3885 2020 3890 2025
rect 3920 2020 3925 2050
rect 3885 2015 3925 2020
rect 4085 2050 4125 2055
rect 4085 2020 4090 2050
rect 4120 2045 4125 2050
rect 4445 2050 4485 2055
rect 4445 2045 4450 2050
rect 4120 2025 4450 2045
rect 4120 2020 4125 2025
rect 4085 2015 4125 2020
rect 4445 2020 4450 2025
rect 4480 2045 4485 2050
rect 4805 2050 4845 2055
rect 4805 2045 4810 2050
rect 4480 2025 4810 2045
rect 4480 2020 4485 2025
rect 4445 2015 4485 2020
rect 4805 2020 4810 2025
rect 4840 2045 4845 2050
rect 5165 2050 5205 2055
rect 5165 2045 5170 2050
rect 4840 2025 5170 2045
rect 4840 2020 4845 2025
rect 4805 2015 4845 2020
rect 5165 2020 5170 2025
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 9790 2010 9825 2011
rect 9790 2005 9885 2010
rect 9825 1970 9850 2005
rect 9790 1965 9885 1970
rect 9910 2005 9945 2011
rect 9910 1965 9945 1970
rect 9970 2005 10005 2010
rect 13795 2005 13830 2010
rect 10020 2000 10060 2005
rect 10020 1995 10025 2000
rect 10005 1975 10025 1995
rect 9970 1965 10005 1970
rect 10020 1970 10025 1975
rect 10055 1970 10060 2000
rect 10020 1965 10060 1970
rect 13740 2000 13780 2005
rect 13740 1970 13745 2000
rect 13775 1995 13780 2000
rect 13775 1975 13795 1995
rect 13775 1970 13780 1975
rect 13740 1965 13780 1970
rect 13795 1965 13830 1970
rect 13855 2005 13890 2011
rect 13975 2010 14010 2011
rect 13855 1965 13890 1970
rect 13915 2005 14010 2010
rect 13950 1970 13975 2005
rect 13915 1965 14010 1970
rect 24735 2000 24775 2005
rect 24735 1970 24740 2000
rect 24770 1995 24775 2000
rect 24845 2000 24885 2005
rect 24845 1995 24850 2000
rect 24770 1975 24850 1995
rect 24770 1970 24775 1975
rect 24735 1965 24775 1970
rect 24845 1970 24850 1975
rect 24880 1995 24885 2000
rect 24955 2000 24995 2005
rect 24955 1995 24960 2000
rect 24880 1975 24960 1995
rect 24880 1970 24885 1975
rect 24845 1965 24885 1970
rect 24955 1970 24960 1975
rect 24990 1995 24995 2000
rect 25065 2000 25105 2005
rect 25065 1995 25070 2000
rect 24990 1975 25070 1995
rect 24990 1970 24995 1975
rect 24955 1965 24995 1970
rect 25065 1970 25070 1975
rect 25100 1995 25105 2000
rect 25175 2000 25215 2005
rect 25175 1995 25180 2000
rect 25100 1975 25180 1995
rect 25100 1970 25105 1975
rect 25065 1965 25105 1970
rect 25175 1970 25180 1975
rect 25210 1995 25215 2000
rect 25285 2000 25325 2005
rect 25285 1995 25290 2000
rect 25210 1975 25290 1995
rect 25210 1970 25215 1975
rect 25175 1965 25215 1970
rect 25285 1970 25290 1975
rect 25320 1995 25325 2000
rect 25395 2000 25435 2005
rect 25395 1995 25400 2000
rect 25320 1975 25400 1995
rect 25320 1970 25325 1975
rect 25285 1965 25325 1970
rect 25395 1970 25400 1975
rect 25430 1995 25435 2000
rect 25505 2000 25545 2005
rect 25505 1995 25510 2000
rect 25430 1975 25510 1995
rect 25430 1970 25435 1975
rect 25395 1965 25435 1970
rect 25505 1970 25510 1975
rect 25540 1995 25545 2000
rect 25615 2000 25655 2005
rect 25615 1995 25620 2000
rect 25540 1975 25620 1995
rect 25540 1970 25545 1975
rect 25505 1965 25545 1970
rect 25615 1970 25620 1975
rect 25650 1995 25655 2000
rect 25725 2000 25765 2005
rect 25725 1995 25730 2000
rect 25650 1975 25730 1995
rect 25650 1970 25655 1975
rect 25615 1965 25655 1970
rect 25725 1970 25730 1975
rect 25760 1995 25765 2000
rect 25835 2000 25875 2005
rect 25835 1995 25840 2000
rect 25760 1975 25840 1995
rect 25760 1970 25765 1975
rect 25725 1965 25765 1970
rect 25835 1970 25840 1975
rect 25870 1970 25875 2000
rect 25835 1965 25875 1970
rect 27945 2000 27985 2005
rect 27945 1970 27950 2000
rect 27980 1995 27985 2000
rect 28055 2000 28095 2005
rect 28055 1995 28060 2000
rect 27980 1975 28060 1995
rect 27980 1970 27985 1975
rect 27945 1965 27985 1970
rect 28055 1970 28060 1975
rect 28090 1995 28095 2000
rect 28165 2000 28205 2005
rect 28165 1995 28170 2000
rect 28090 1975 28170 1995
rect 28090 1970 28095 1975
rect 28055 1965 28095 1970
rect 28165 1970 28170 1975
rect 28200 1995 28205 2000
rect 28275 2000 28315 2005
rect 28275 1995 28280 2000
rect 28200 1975 28280 1995
rect 28200 1970 28205 1975
rect 28165 1965 28205 1970
rect 28275 1970 28280 1975
rect 28310 1995 28315 2000
rect 28385 2000 28425 2005
rect 28385 1995 28390 2000
rect 28310 1975 28390 1995
rect 28310 1970 28315 1975
rect 28275 1965 28315 1970
rect 28385 1970 28390 1975
rect 28420 1995 28425 2000
rect 28495 2000 28535 2005
rect 28495 1995 28500 2000
rect 28420 1975 28500 1995
rect 28420 1970 28425 1975
rect 28385 1965 28425 1970
rect 28495 1970 28500 1975
rect 28530 1995 28535 2000
rect 28605 2000 28645 2005
rect 28605 1995 28610 2000
rect 28530 1975 28610 1995
rect 28530 1970 28535 1975
rect 28495 1965 28535 1970
rect 28605 1970 28610 1975
rect 28640 1995 28645 2000
rect 28715 2000 28755 2005
rect 28715 1995 28720 2000
rect 28640 1975 28720 1995
rect 28640 1970 28645 1975
rect 28605 1965 28645 1970
rect 28715 1970 28720 1975
rect 28750 1995 28755 2000
rect 28825 2000 28865 2005
rect 28825 1995 28830 2000
rect 28750 1975 28830 1995
rect 28750 1970 28755 1975
rect 28715 1965 28755 1970
rect 28825 1970 28830 1975
rect 28860 1995 28865 2000
rect 28935 2000 28975 2005
rect 28935 1995 28940 2000
rect 28860 1975 28940 1995
rect 28860 1970 28865 1975
rect 28825 1965 28865 1970
rect 28935 1970 28940 1975
rect 28970 1995 28975 2000
rect 29045 2000 29085 2005
rect 29045 1995 29050 2000
rect 28970 1975 29050 1995
rect 28970 1970 28975 1975
rect 28935 1965 28975 1970
rect 29045 1970 29050 1975
rect 29080 1970 29085 2000
rect 29045 1965 29085 1970
rect 11385 1960 11425 1965
rect 9910 1945 9950 1950
rect 9910 1915 9915 1945
rect 9945 1940 9950 1945
rect 10065 1945 10105 1950
rect 10065 1940 10070 1945
rect 9945 1920 10070 1940
rect 9945 1915 9950 1920
rect 9910 1910 9950 1915
rect 10065 1915 10070 1920
rect 10100 1915 10105 1945
rect 10065 1910 10105 1915
rect 10210 1945 10250 1950
rect 10210 1915 10215 1945
rect 10245 1940 10250 1945
rect 10320 1945 10360 1950
rect 10320 1940 10325 1945
rect 10245 1920 10325 1940
rect 10245 1915 10250 1920
rect 10210 1910 10250 1915
rect 10320 1915 10325 1920
rect 10355 1940 10360 1945
rect 10430 1945 10470 1950
rect 10430 1940 10435 1945
rect 10355 1920 10435 1940
rect 10355 1915 10360 1920
rect 10320 1910 10360 1915
rect 10430 1915 10435 1920
rect 10465 1940 10470 1945
rect 10540 1945 10580 1950
rect 10540 1940 10545 1945
rect 10465 1920 10545 1940
rect 10465 1915 10470 1920
rect 10430 1910 10470 1915
rect 10540 1915 10545 1920
rect 10575 1940 10580 1945
rect 10650 1945 10690 1950
rect 10650 1940 10655 1945
rect 10575 1920 10655 1940
rect 10575 1915 10580 1920
rect 10540 1910 10580 1915
rect 10650 1915 10655 1920
rect 10685 1940 10690 1945
rect 10760 1945 10800 1950
rect 10760 1940 10765 1945
rect 10685 1920 10765 1940
rect 10685 1915 10690 1920
rect 10650 1910 10690 1915
rect 10760 1915 10765 1920
rect 10795 1915 10800 1945
rect 11385 1930 11390 1960
rect 11420 1955 11425 1960
rect 11605 1960 11645 1965
rect 11605 1955 11610 1960
rect 11420 1935 11610 1955
rect 11420 1930 11425 1935
rect 11385 1925 11425 1930
rect 11605 1930 11610 1935
rect 11640 1955 11645 1960
rect 11825 1960 11865 1965
rect 11825 1955 11830 1960
rect 11640 1935 11830 1955
rect 11640 1930 11645 1935
rect 11605 1925 11645 1930
rect 11825 1930 11830 1935
rect 11860 1955 11865 1960
rect 12045 1960 12085 1965
rect 12045 1955 12050 1960
rect 11860 1935 12050 1955
rect 11860 1930 11865 1935
rect 11825 1925 11865 1930
rect 12045 1930 12050 1935
rect 12080 1955 12085 1960
rect 12265 1960 12305 1965
rect 12265 1955 12270 1960
rect 12080 1935 12270 1955
rect 12080 1930 12085 1935
rect 12045 1925 12085 1930
rect 12265 1930 12270 1935
rect 12300 1930 12305 1960
rect 26385 1960 26425 1965
rect 12265 1925 12305 1930
rect 13000 1945 13040 1950
rect 10760 1910 10800 1915
rect 13000 1915 13005 1945
rect 13035 1940 13040 1945
rect 13110 1945 13150 1950
rect 13110 1940 13115 1945
rect 13035 1920 13115 1940
rect 13035 1915 13040 1920
rect 13000 1910 13040 1915
rect 13110 1915 13115 1920
rect 13145 1940 13150 1945
rect 13220 1945 13260 1950
rect 13220 1940 13225 1945
rect 13145 1920 13225 1940
rect 13145 1915 13150 1920
rect 13110 1910 13150 1915
rect 13220 1915 13225 1920
rect 13255 1940 13260 1945
rect 13330 1945 13370 1950
rect 13330 1940 13335 1945
rect 13255 1920 13335 1940
rect 13255 1915 13260 1920
rect 13220 1910 13260 1915
rect 13330 1915 13335 1920
rect 13365 1940 13370 1945
rect 13440 1945 13480 1950
rect 13440 1940 13445 1945
rect 13365 1920 13445 1940
rect 13365 1915 13370 1920
rect 13330 1910 13370 1915
rect 13440 1915 13445 1920
rect 13475 1940 13480 1945
rect 13550 1945 13590 1950
rect 13550 1940 13555 1945
rect 13475 1920 13555 1940
rect 13475 1915 13480 1920
rect 13440 1910 13480 1915
rect 13550 1915 13555 1920
rect 13585 1915 13590 1945
rect 13550 1910 13590 1915
rect 13695 1945 13735 1950
rect 13695 1915 13700 1945
rect 13730 1940 13735 1945
rect 13850 1945 13890 1950
rect 13850 1940 13855 1945
rect 13730 1920 13855 1940
rect 13730 1915 13735 1920
rect 13695 1910 13735 1915
rect 13850 1915 13855 1920
rect 13885 1915 13890 1945
rect 26385 1930 26390 1960
rect 26420 1955 26425 1960
rect 26605 1960 26645 1965
rect 26605 1955 26610 1960
rect 26420 1935 26610 1955
rect 26420 1930 26425 1935
rect 26385 1925 26425 1930
rect 26605 1930 26610 1935
rect 26640 1955 26645 1960
rect 26825 1960 26865 1965
rect 26825 1955 26830 1960
rect 26640 1935 26830 1955
rect 26640 1930 26645 1935
rect 26605 1925 26645 1930
rect 26825 1930 26830 1935
rect 26860 1955 26865 1960
rect 27045 1960 27085 1965
rect 27045 1955 27050 1960
rect 26860 1935 27050 1955
rect 26860 1930 26865 1935
rect 26825 1925 26865 1930
rect 27045 1930 27050 1935
rect 27080 1955 27085 1960
rect 27265 1960 27305 1965
rect 27265 1955 27270 1960
rect 27080 1935 27270 1955
rect 27080 1930 27085 1935
rect 27045 1925 27085 1930
rect 27265 1930 27270 1935
rect 27300 1930 27305 1960
rect 27265 1925 27305 1930
rect 13850 1910 13890 1915
rect 11495 1905 11535 1910
rect 9790 1895 9830 1900
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1875 2965 1880
rect 3045 1875 3085 1885
rect 3285 1880 3325 1885
rect 3285 1875 3290 1880
rect 2960 1855 3290 1875
rect 2960 1850 2965 1855
rect 2925 1845 2965 1850
rect 3045 1845 3085 1855
rect 3285 1850 3290 1855
rect 3320 1875 3325 1880
rect 3405 1875 3445 1885
rect 3645 1880 3685 1885
rect 3645 1875 3650 1880
rect 3320 1855 3650 1875
rect 3320 1850 3325 1855
rect 3285 1845 3325 1850
rect 3405 1845 3445 1855
rect 3645 1850 3650 1855
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1845 3805 1885
rect 4205 1845 4245 1885
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1875 4365 1880
rect 4565 1875 4605 1885
rect 4685 1880 4725 1885
rect 4685 1875 4690 1880
rect 4360 1855 4690 1875
rect 4360 1850 4365 1855
rect 4325 1845 4365 1850
rect 4565 1845 4605 1855
rect 4685 1850 4690 1855
rect 4720 1875 4725 1880
rect 4925 1875 4965 1885
rect 5045 1880 5085 1885
rect 5045 1875 5050 1880
rect 4720 1855 5050 1875
rect 4720 1850 4725 1855
rect 4685 1845 4725 1850
rect 4925 1845 4965 1855
rect 5045 1850 5050 1855
rect 5080 1875 5085 1880
rect 5080 1855 5175 1875
rect 9790 1865 9795 1895
rect 9825 1890 9830 1895
rect 11000 1895 11040 1900
rect 11000 1890 11005 1895
rect 9825 1870 11005 1890
rect 9825 1865 9830 1870
rect 9790 1860 9830 1865
rect 11000 1865 11005 1870
rect 11035 1865 11040 1895
rect 11495 1875 11500 1905
rect 11530 1900 11535 1905
rect 11715 1905 11755 1910
rect 11715 1900 11720 1905
rect 11530 1880 11720 1900
rect 11530 1875 11535 1880
rect 11495 1870 11535 1875
rect 11715 1875 11720 1880
rect 11750 1900 11755 1905
rect 11935 1905 11975 1910
rect 11935 1900 11940 1905
rect 11750 1880 11940 1900
rect 11750 1875 11755 1880
rect 11715 1870 11755 1875
rect 11935 1875 11940 1880
rect 11970 1900 11975 1905
rect 12155 1905 12195 1910
rect 12155 1900 12160 1905
rect 11970 1880 12160 1900
rect 11970 1875 11975 1880
rect 11935 1870 11975 1875
rect 12155 1875 12160 1880
rect 12190 1900 12195 1905
rect 12375 1905 12415 1910
rect 12375 1900 12380 1905
rect 12190 1880 12380 1900
rect 12190 1875 12195 1880
rect 12155 1870 12195 1875
rect 12375 1875 12380 1880
rect 12410 1875 12415 1905
rect 26495 1905 26535 1910
rect 12375 1870 12415 1875
rect 12760 1895 12800 1900
rect 11000 1860 11040 1865
rect 12760 1865 12765 1895
rect 12795 1890 12800 1895
rect 13970 1895 14010 1900
rect 13970 1890 13975 1895
rect 12795 1870 13975 1890
rect 12795 1865 12800 1870
rect 12760 1860 12800 1865
rect 13970 1865 13975 1870
rect 14005 1865 14010 1895
rect 26495 1875 26500 1905
rect 26530 1900 26535 1905
rect 26715 1905 26755 1910
rect 26715 1900 26720 1905
rect 26530 1880 26720 1900
rect 26530 1875 26535 1880
rect 26495 1870 26535 1875
rect 26715 1875 26720 1880
rect 26750 1900 26755 1905
rect 26935 1905 26975 1910
rect 26935 1900 26940 1905
rect 26750 1880 26940 1900
rect 26750 1875 26755 1880
rect 26715 1870 26755 1875
rect 26935 1875 26940 1880
rect 26970 1900 26975 1905
rect 27155 1905 27195 1910
rect 27155 1900 27160 1905
rect 26970 1880 27160 1900
rect 26970 1875 26975 1880
rect 26935 1870 26975 1875
rect 27155 1875 27160 1880
rect 27190 1900 27195 1905
rect 27375 1905 27415 1910
rect 27375 1900 27380 1905
rect 27190 1880 27380 1900
rect 27190 1875 27195 1880
rect 27155 1870 27195 1875
rect 27375 1875 27380 1880
rect 27410 1875 27415 1905
rect 27375 1870 27415 1875
rect 28045 1905 28085 1910
rect 28045 1875 28050 1905
rect 28080 1900 28085 1905
rect 28155 1905 28195 1910
rect 28155 1900 28160 1905
rect 28080 1880 28160 1900
rect 28080 1875 28085 1880
rect 28045 1870 28085 1875
rect 28155 1875 28160 1880
rect 28190 1900 28195 1905
rect 28265 1905 28305 1910
rect 28265 1900 28270 1905
rect 28190 1880 28270 1900
rect 28190 1875 28195 1880
rect 28155 1870 28195 1875
rect 28265 1875 28270 1880
rect 28300 1875 28305 1905
rect 28265 1870 28305 1875
rect 13970 1860 14010 1865
rect 5080 1850 5085 1855
rect 5045 1845 5085 1850
rect 11190 1850 11230 1855
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2835 1820 2875 1825
rect 2835 1815 2840 1820
rect 2505 1795 2840 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2835 1790 2840 1795
rect 2870 1815 2875 1820
rect 3045 1820 3085 1825
rect 3045 1815 3050 1820
rect 2870 1795 3050 1815
rect 2870 1790 2875 1795
rect 2835 1785 2875 1790
rect 3045 1790 3050 1795
rect 3080 1815 3085 1820
rect 3165 1820 3205 1825
rect 3165 1815 3170 1820
rect 3080 1795 3170 1815
rect 3080 1790 3085 1795
rect 3045 1785 3085 1790
rect 3165 1790 3170 1795
rect 3200 1815 3205 1820
rect 3405 1820 3445 1825
rect 3405 1815 3410 1820
rect 3200 1795 3410 1815
rect 3200 1790 3205 1795
rect 3165 1785 3205 1790
rect 3405 1790 3410 1795
rect 3440 1815 3445 1820
rect 3525 1820 3565 1825
rect 3525 1815 3530 1820
rect 3440 1795 3530 1815
rect 3440 1790 3445 1795
rect 3405 1785 3445 1790
rect 3525 1790 3530 1795
rect 3560 1815 3565 1820
rect 3765 1820 3805 1825
rect 3765 1815 3770 1820
rect 3560 1795 3770 1815
rect 3560 1790 3565 1795
rect 3525 1785 3565 1790
rect 3765 1790 3770 1795
rect 3800 1815 3805 1820
rect 3855 1820 3895 1825
rect 3855 1815 3860 1820
rect 3800 1795 3860 1815
rect 3800 1790 3805 1795
rect 3765 1785 3805 1790
rect 3855 1790 3860 1795
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1815 4155 1820
rect 4205 1820 4245 1825
rect 4205 1815 4210 1820
rect 4150 1795 4210 1815
rect 4150 1790 4155 1795
rect 4115 1785 4155 1790
rect 4205 1790 4210 1795
rect 4240 1815 4245 1820
rect 4445 1820 4485 1825
rect 4445 1815 4450 1820
rect 4240 1795 4450 1815
rect 4240 1790 4245 1795
rect 4205 1785 4245 1790
rect 4445 1790 4450 1795
rect 4480 1815 4485 1820
rect 4565 1820 4605 1825
rect 4565 1815 4570 1820
rect 4480 1795 4570 1815
rect 4480 1790 4485 1795
rect 4445 1785 4485 1790
rect 4565 1790 4570 1795
rect 4600 1815 4605 1820
rect 4805 1820 4845 1825
rect 4805 1815 4810 1820
rect 4600 1795 4810 1815
rect 4600 1790 4605 1795
rect 4565 1785 4605 1790
rect 4805 1790 4810 1795
rect 4840 1815 4845 1820
rect 4925 1820 4965 1825
rect 4925 1815 4930 1820
rect 4840 1795 4930 1815
rect 4840 1790 4845 1795
rect 4805 1785 4845 1790
rect 4925 1790 4930 1795
rect 4960 1815 4965 1820
rect 5135 1820 5175 1825
rect 5135 1815 5140 1820
rect 4960 1795 5140 1815
rect 4960 1790 4965 1795
rect 4925 1785 4965 1790
rect 5135 1790 5140 1795
rect 5170 1815 5175 1820
rect 5360 1820 5400 1825
rect 5360 1815 5365 1820
rect 5170 1795 5365 1815
rect 5170 1790 5175 1795
rect 5135 1785 5175 1790
rect 5360 1790 5365 1795
rect 5395 1790 5400 1820
rect 11190 1820 11195 1850
rect 11225 1845 11230 1850
rect 11410 1850 11450 1855
rect 11410 1845 11415 1850
rect 11225 1825 11415 1845
rect 11225 1820 11230 1825
rect 11190 1815 11230 1820
rect 11410 1820 11415 1825
rect 11445 1845 11450 1850
rect 11640 1850 11680 1855
rect 11640 1845 11645 1850
rect 11445 1825 11645 1845
rect 11445 1820 11450 1825
rect 11410 1815 11450 1820
rect 11640 1820 11645 1825
rect 11675 1845 11680 1850
rect 12230 1850 12270 1855
rect 12230 1845 12235 1850
rect 11675 1825 12235 1845
rect 11675 1820 11680 1825
rect 11640 1815 11680 1820
rect 12230 1820 12235 1825
rect 12265 1845 12270 1850
rect 12450 1850 12490 1855
rect 12450 1845 12455 1850
rect 12265 1825 12455 1845
rect 12265 1820 12270 1825
rect 12230 1815 12270 1820
rect 12450 1820 12455 1825
rect 12485 1845 12490 1850
rect 12680 1850 12720 1855
rect 12680 1845 12685 1850
rect 12485 1825 12685 1845
rect 12485 1820 12490 1825
rect 12450 1815 12490 1820
rect 12680 1820 12685 1825
rect 12715 1820 12720 1850
rect 12680 1815 12720 1820
rect 26190 1850 26230 1855
rect 26190 1820 26195 1850
rect 26225 1845 26230 1850
rect 26410 1850 26450 1855
rect 26410 1845 26415 1850
rect 26225 1825 26415 1845
rect 26225 1820 26230 1825
rect 26190 1815 26230 1820
rect 26410 1820 26415 1825
rect 26445 1845 26450 1850
rect 26640 1850 26680 1855
rect 26640 1845 26645 1850
rect 26445 1825 26645 1845
rect 26445 1820 26450 1825
rect 26410 1815 26450 1820
rect 26640 1820 26645 1825
rect 26675 1845 26680 1850
rect 27230 1850 27270 1855
rect 27230 1845 27235 1850
rect 26675 1825 27235 1845
rect 26675 1820 26680 1825
rect 26640 1815 26680 1820
rect 27230 1820 27235 1825
rect 27265 1845 27270 1850
rect 27450 1850 27490 1855
rect 27450 1845 27455 1850
rect 27265 1825 27455 1845
rect 27265 1820 27270 1825
rect 27230 1815 27270 1820
rect 27450 1820 27455 1825
rect 27485 1845 27490 1850
rect 27680 1850 27720 1855
rect 27680 1845 27685 1850
rect 27485 1825 27685 1845
rect 27485 1820 27490 1825
rect 27450 1815 27490 1820
rect 27680 1820 27685 1825
rect 27715 1820 27720 1850
rect 27680 1815 27720 1820
rect 5360 1785 5400 1790
rect 11820 1805 11860 1810
rect 11820 1775 11825 1805
rect 11855 1800 11860 1805
rect 11940 1805 11980 1810
rect 11940 1800 11945 1805
rect 11855 1780 11945 1800
rect 11855 1775 11860 1780
rect 11820 1770 11860 1775
rect 11940 1775 11945 1780
rect 11975 1775 11980 1805
rect 11940 1770 11980 1775
rect 26820 1805 26860 1810
rect 26820 1775 26825 1805
rect 26855 1800 26860 1805
rect 26940 1805 26980 1810
rect 26940 1800 26945 1805
rect 26855 1780 26945 1800
rect 26855 1775 26860 1780
rect 26820 1770 26860 1775
rect 26940 1775 26945 1780
rect 26975 1775 26980 1805
rect 26940 1770 26980 1775
rect 2800 1765 2840 1770
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2565 1760 2605 1765
rect 2565 1755 2570 1760
rect 2460 1735 2570 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2565 1730 2570 1735
rect 2600 1755 2605 1760
rect 2675 1760 2715 1765
rect 2675 1755 2680 1760
rect 2600 1735 2680 1755
rect 2600 1730 2605 1735
rect 2565 1725 2605 1730
rect 2675 1730 2680 1735
rect 2710 1755 2715 1760
rect 2800 1755 2805 1765
rect 2710 1735 2805 1755
rect 2835 1755 2840 1765
rect 3225 1760 3265 1765
rect 3225 1755 3230 1760
rect 2835 1735 3230 1755
rect 2710 1730 2715 1735
rect 2800 1730 2840 1735
rect 3225 1730 3230 1735
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1755 3325 1760
rect 3525 1760 3565 1765
rect 3525 1755 3530 1760
rect 3320 1735 3530 1755
rect 3320 1730 3325 1735
rect 3285 1725 3325 1730
rect 3525 1730 3530 1735
rect 3560 1755 3565 1760
rect 3765 1760 3805 1765
rect 3765 1755 3770 1760
rect 3560 1735 3770 1755
rect 3560 1730 3565 1735
rect 3525 1725 3565 1730
rect 3765 1730 3770 1735
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1755 4245 1760
rect 4445 1760 4485 1765
rect 4445 1755 4450 1760
rect 4240 1735 4450 1755
rect 4240 1730 4245 1735
rect 4205 1725 4245 1730
rect 4445 1730 4450 1735
rect 4480 1755 4485 1760
rect 4685 1760 4725 1765
rect 4685 1755 4690 1760
rect 4480 1735 4690 1755
rect 4480 1730 4485 1735
rect 4445 1725 4485 1730
rect 4685 1730 4690 1735
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1755 4785 1760
rect 5270 1760 5310 1765
rect 5270 1755 5275 1760
rect 4780 1735 5275 1755
rect 4780 1730 4785 1735
rect 4745 1725 4785 1730
rect 5270 1730 5275 1735
rect 5305 1755 5310 1760
rect 9965 1760 10005 1765
rect 5305 1735 6100 1755
rect 5305 1730 5310 1735
rect 5270 1725 5310 1730
rect 9965 1730 9970 1760
rect 10000 1755 10005 1760
rect 10555 1760 10595 1765
rect 10555 1755 10560 1760
rect 10000 1735 10560 1755
rect 10000 1730 10005 1735
rect 9965 1725 10005 1730
rect 10555 1730 10560 1735
rect 10590 1730 10595 1760
rect 10555 1725 10595 1730
rect 11085 1760 11125 1765
rect 11085 1730 11090 1760
rect 11120 1755 11125 1760
rect 11305 1760 11345 1765
rect 11305 1755 11310 1760
rect 11120 1735 11310 1755
rect 11120 1730 11125 1735
rect 11085 1725 11125 1730
rect 11305 1730 11310 1735
rect 11340 1755 11345 1760
rect 11525 1760 11565 1765
rect 11525 1755 11530 1760
rect 11340 1735 11530 1755
rect 11340 1730 11345 1735
rect 11305 1725 11345 1730
rect 11525 1730 11530 1735
rect 11560 1755 11565 1760
rect 12125 1760 12165 1765
rect 12125 1755 12130 1760
rect 11560 1735 12130 1755
rect 11560 1730 11565 1735
rect 11525 1725 11565 1730
rect 12125 1730 12130 1735
rect 12160 1755 12165 1760
rect 12345 1760 12385 1765
rect 12345 1755 12350 1760
rect 12160 1735 12350 1755
rect 12160 1730 12165 1735
rect 12125 1725 12165 1730
rect 12345 1730 12350 1735
rect 12380 1755 12385 1760
rect 12565 1760 12605 1765
rect 12565 1755 12570 1760
rect 12380 1735 12570 1755
rect 12380 1730 12385 1735
rect 12345 1725 12385 1730
rect 12565 1730 12570 1735
rect 12600 1730 12605 1760
rect 12565 1725 12605 1730
rect 13205 1760 13245 1765
rect 13205 1730 13210 1760
rect 13240 1755 13245 1760
rect 13795 1760 13835 1765
rect 13795 1755 13800 1760
rect 13240 1735 13800 1755
rect 13240 1730 13245 1735
rect 13205 1725 13245 1730
rect 13795 1730 13800 1735
rect 13830 1730 13835 1760
rect 13795 1725 13835 1730
rect 26085 1760 26125 1765
rect 26085 1730 26090 1760
rect 26120 1755 26125 1760
rect 26305 1760 26345 1765
rect 26305 1755 26310 1760
rect 26120 1735 26310 1755
rect 26120 1730 26125 1735
rect 26085 1725 26125 1730
rect 26305 1730 26310 1735
rect 26340 1755 26345 1760
rect 26525 1760 26565 1765
rect 26525 1755 26530 1760
rect 26340 1735 26530 1755
rect 26340 1730 26345 1735
rect 26305 1725 26345 1730
rect 26525 1730 26530 1735
rect 26560 1755 26565 1760
rect 27125 1760 27165 1765
rect 27125 1755 27130 1760
rect 26560 1735 27130 1755
rect 26560 1730 26565 1735
rect 26525 1725 26565 1730
rect 27125 1730 27130 1735
rect 27160 1755 27165 1760
rect 27345 1760 27385 1765
rect 27345 1755 27350 1760
rect 27160 1735 27350 1755
rect 27160 1730 27165 1735
rect 27125 1725 27165 1730
rect 27345 1730 27350 1735
rect 27380 1755 27385 1760
rect 27565 1760 27605 1765
rect 27565 1755 27570 1760
rect 27380 1735 27570 1755
rect 27380 1730 27385 1735
rect 27345 1725 27385 1730
rect 27565 1730 27570 1735
rect 27600 1730 27605 1760
rect 27565 1725 27605 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3165 1715 3205 1720
rect -45 1685 -5 1690
rect 1262 1710 1302 1715
rect 1262 1680 1270 1710
rect 1297 1705 1302 1710
rect 2800 1710 2840 1715
rect 2800 1705 2805 1710
rect 1297 1685 2805 1705
rect 1297 1680 1302 1685
rect 1262 1675 1302 1680
rect 2800 1680 2805 1685
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1710 3205 1715
rect 3405 1715 3445 1720
rect 3405 1710 3410 1715
rect 3200 1690 3410 1710
rect 3200 1685 3205 1690
rect 3165 1680 3205 1685
rect 3405 1685 3410 1690
rect 3440 1710 3445 1715
rect 3645 1715 3685 1720
rect 3645 1710 3650 1715
rect 3440 1690 3650 1710
rect 3440 1685 3445 1690
rect 3405 1680 3445 1685
rect 3645 1685 3650 1690
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1710 4365 1715
rect 4565 1715 4605 1720
rect 4565 1710 4570 1715
rect 4360 1690 4570 1710
rect 4360 1685 4365 1690
rect 4325 1680 4365 1685
rect 4565 1685 4570 1690
rect 4600 1710 4605 1715
rect 4805 1715 4845 1720
rect 4805 1710 4810 1715
rect 4600 1690 4810 1710
rect 4600 1685 4605 1690
rect 4565 1680 4605 1685
rect 4805 1685 4810 1690
rect 4840 1685 4845 1715
rect 11237 1715 11269 1720
rect 11237 1710 11240 1715
rect 4805 1680 4845 1685
rect 9745 1705 9785 1710
rect 2800 1675 2840 1680
rect 9745 1675 9750 1705
rect 9780 1700 9785 1705
rect 10030 1705 10070 1710
rect 10030 1700 10035 1705
rect 9780 1680 10035 1700
rect 9780 1675 9785 1680
rect 9745 1670 9785 1675
rect 10030 1675 10035 1680
rect 10065 1700 10070 1705
rect 10255 1705 10295 1710
rect 10255 1700 10260 1705
rect 10065 1680 10260 1700
rect 10065 1675 10070 1680
rect 10030 1670 10070 1675
rect 10255 1675 10260 1680
rect 10290 1700 10295 1705
rect 10455 1705 10495 1710
rect 10455 1700 10460 1705
rect 10290 1680 10460 1700
rect 10290 1675 10295 1680
rect 10255 1670 10295 1675
rect 10455 1675 10460 1680
rect 10490 1700 10495 1705
rect 10655 1705 10695 1710
rect 10655 1700 10660 1705
rect 10490 1680 10660 1700
rect 10490 1675 10495 1680
rect 10455 1670 10495 1675
rect 10655 1675 10660 1680
rect 10690 1700 10695 1705
rect 10835 1705 10875 1710
rect 10835 1700 10840 1705
rect 10690 1680 10840 1700
rect 10690 1675 10695 1680
rect 10655 1670 10695 1675
rect 10835 1675 10840 1680
rect 10870 1675 10875 1705
rect 10910 1690 11240 1710
rect 11237 1685 11240 1690
rect 11266 1710 11269 1715
rect 11457 1715 11489 1720
rect 11457 1710 11460 1715
rect 11266 1690 11460 1710
rect 11266 1685 11269 1690
rect 11237 1680 11269 1685
rect 11457 1685 11460 1690
rect 11486 1710 11489 1715
rect 11601 1715 11633 1720
rect 11601 1710 11604 1715
rect 11486 1690 11604 1710
rect 11486 1685 11489 1690
rect 11457 1680 11489 1685
rect 11601 1685 11604 1690
rect 11630 1710 11633 1715
rect 11867 1715 11899 1720
rect 11867 1710 11870 1715
rect 11630 1690 11870 1710
rect 11630 1685 11633 1690
rect 11601 1680 11633 1685
rect 11867 1685 11870 1690
rect 11896 1710 11899 1715
rect 12277 1715 12309 1720
rect 12277 1710 12280 1715
rect 11896 1690 12280 1710
rect 11896 1685 11899 1690
rect 11867 1680 11899 1685
rect 12277 1685 12280 1690
rect 12306 1710 12309 1715
rect 12497 1715 12529 1720
rect 12497 1710 12500 1715
rect 12306 1690 12500 1710
rect 12306 1685 12309 1690
rect 12277 1680 12309 1685
rect 12497 1685 12500 1690
rect 12526 1710 12529 1715
rect 12641 1715 12673 1720
rect 12641 1710 12644 1715
rect 12526 1690 12644 1710
rect 12526 1685 12529 1690
rect 12497 1680 12529 1685
rect 12641 1685 12644 1690
rect 12670 1685 12673 1715
rect 26237 1715 26269 1720
rect 26237 1710 26240 1715
rect 12641 1680 12673 1685
rect 12925 1705 12965 1710
rect 10835 1670 10875 1675
rect 12925 1675 12930 1705
rect 12960 1700 12965 1705
rect 13105 1705 13145 1710
rect 13105 1700 13110 1705
rect 12960 1680 13110 1700
rect 12960 1675 12965 1680
rect 12925 1670 12965 1675
rect 13105 1675 13110 1680
rect 13140 1700 13145 1705
rect 13305 1705 13345 1710
rect 13305 1700 13310 1705
rect 13140 1680 13310 1700
rect 13140 1675 13145 1680
rect 13105 1670 13145 1675
rect 13305 1675 13310 1680
rect 13340 1700 13345 1705
rect 13505 1705 13545 1710
rect 13505 1700 13510 1705
rect 13340 1680 13510 1700
rect 13340 1675 13345 1680
rect 13305 1670 13345 1675
rect 13505 1675 13510 1680
rect 13540 1700 13545 1705
rect 13730 1705 13770 1710
rect 13730 1700 13735 1705
rect 13540 1680 13735 1700
rect 13540 1675 13545 1680
rect 13505 1670 13545 1675
rect 13730 1675 13735 1680
rect 13765 1700 13770 1705
rect 14015 1705 14055 1710
rect 14015 1700 14020 1705
rect 13765 1680 14020 1700
rect 13765 1675 13770 1680
rect 13730 1670 13770 1675
rect 14015 1675 14020 1680
rect 14050 1675 14055 1705
rect 25910 1690 26240 1710
rect 26237 1685 26240 1690
rect 26266 1710 26269 1715
rect 26457 1715 26489 1720
rect 26457 1710 26460 1715
rect 26266 1690 26460 1710
rect 26266 1685 26269 1690
rect 26237 1680 26269 1685
rect 26457 1685 26460 1690
rect 26486 1710 26489 1715
rect 26601 1715 26633 1720
rect 26601 1710 26604 1715
rect 26486 1690 26604 1710
rect 26486 1685 26489 1690
rect 26457 1680 26489 1685
rect 26601 1685 26604 1690
rect 26630 1710 26633 1715
rect 26867 1715 26899 1720
rect 26867 1710 26870 1715
rect 26630 1690 26870 1710
rect 26630 1685 26633 1690
rect 26601 1680 26633 1685
rect 26867 1685 26870 1690
rect 26896 1710 26899 1715
rect 27277 1715 27309 1720
rect 27277 1710 27280 1715
rect 26896 1690 27280 1710
rect 26896 1685 26899 1690
rect 26867 1680 26899 1685
rect 27277 1685 27280 1690
rect 27306 1710 27309 1715
rect 27497 1715 27529 1720
rect 27497 1710 27500 1715
rect 27306 1690 27500 1710
rect 27306 1685 27309 1690
rect 27277 1680 27309 1685
rect 27497 1685 27500 1690
rect 27526 1710 27529 1715
rect 27641 1715 27673 1720
rect 27641 1710 27644 1715
rect 27526 1690 27644 1710
rect 27526 1685 27529 1690
rect 27497 1680 27529 1685
rect 27641 1685 27644 1690
rect 27670 1685 27673 1715
rect 27641 1680 27673 1685
rect 28066 1680 28098 1685
rect 14015 1670 14055 1675
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2620 1665 2660 1670
rect 2620 1660 2625 1665
rect 2415 1640 2625 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2620 1635 2625 1640
rect 2655 1635 2660 1665
rect 28066 1650 28070 1680
rect 28096 1650 28098 1680
rect 2620 1630 2660 1635
rect 9970 1645 10005 1650
rect 9970 1605 10005 1610
rect 10030 1645 10065 1650
rect 10030 1605 10065 1610
rect 13735 1645 13770 1650
rect 13735 1605 13770 1610
rect 13795 1645 13830 1650
rect 28066 1645 28098 1650
rect 13795 1605 13830 1610
rect 28010 1630 28050 1635
rect 28010 1600 28015 1630
rect 28045 1625 28050 1630
rect 28116 1630 28156 1635
rect 28116 1625 28121 1630
rect 28045 1605 28121 1625
rect 28045 1600 28050 1605
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3165 1595 3205 1600
rect 3165 1590 3170 1595
rect 2365 1570 3170 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3165 1565 3170 1570
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1590 4845 1595
rect 5410 1595 5450 1600
rect 28010 1595 28050 1600
rect 28116 1600 28121 1605
rect 28151 1600 28156 1630
rect 28116 1595 28156 1600
rect 28210 1630 28250 1635
rect 28210 1600 28215 1630
rect 28245 1625 28250 1630
rect 28300 1630 28340 1635
rect 28300 1625 28305 1630
rect 28245 1605 28305 1625
rect 28245 1600 28250 1605
rect 28210 1595 28250 1600
rect 28300 1600 28305 1605
rect 28335 1600 28340 1630
rect 28300 1595 28340 1600
rect 5410 1590 5415 1595
rect 4840 1570 5415 1590
rect 4840 1565 4845 1570
rect 4805 1560 4845 1565
rect 5410 1565 5415 1570
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 27815 1570 27855 1575
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1540 2875 1545
rect 3225 1545 3265 1550
rect 3225 1540 3230 1545
rect 2870 1520 3230 1540
rect 2870 1515 2875 1520
rect 2835 1510 2875 1515
rect 3225 1515 3230 1520
rect 3260 1540 3265 1545
rect 3345 1545 3385 1550
rect 3345 1540 3350 1545
rect 3260 1520 3350 1540
rect 3260 1515 3265 1520
rect 3225 1510 3265 1515
rect 3345 1515 3350 1520
rect 3380 1540 3385 1545
rect 3465 1545 3505 1550
rect 3465 1540 3470 1545
rect 3380 1520 3470 1540
rect 3380 1515 3385 1520
rect 3345 1510 3385 1515
rect 3465 1515 3470 1520
rect 3500 1540 3505 1545
rect 3585 1545 3625 1550
rect 3585 1540 3590 1545
rect 3500 1520 3590 1540
rect 3500 1515 3505 1520
rect 3465 1510 3505 1515
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 3705 1545 3745 1550
rect 3705 1540 3710 1545
rect 3620 1520 3710 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 3705 1515 3710 1520
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1540 4305 1545
rect 4385 1545 4425 1550
rect 4385 1540 4390 1545
rect 4300 1520 4390 1540
rect 4300 1515 4305 1520
rect 4265 1510 4305 1515
rect 4385 1515 4390 1520
rect 4420 1540 4425 1545
rect 4505 1545 4545 1550
rect 4505 1540 4510 1545
rect 4420 1520 4510 1540
rect 4420 1515 4425 1520
rect 4385 1510 4425 1515
rect 4505 1515 4510 1520
rect 4540 1540 4545 1545
rect 4625 1545 4665 1550
rect 4625 1540 4630 1545
rect 4540 1520 4630 1540
rect 4540 1515 4545 1520
rect 4505 1510 4545 1515
rect 4625 1515 4630 1520
rect 4660 1540 4665 1545
rect 4745 1545 4785 1550
rect 4745 1540 4750 1545
rect 4660 1520 4750 1540
rect 4660 1515 4665 1520
rect 4625 1510 4665 1515
rect 4745 1515 4750 1520
rect 4780 1540 4785 1545
rect 5135 1545 5175 1550
rect 5135 1540 5140 1545
rect 4780 1520 5140 1540
rect 4780 1515 4785 1520
rect 4745 1510 4785 1515
rect 5135 1515 5140 1520
rect 5170 1515 5175 1545
rect 27815 1540 27820 1570
rect 27850 1565 27855 1570
rect 27971 1570 28003 1575
rect 27971 1565 27975 1570
rect 27850 1545 27975 1565
rect 27850 1540 27855 1545
rect 27815 1535 27855 1540
rect 27971 1540 27975 1545
rect 28001 1565 28003 1570
rect 28347 1570 28379 1575
rect 28347 1565 28349 1570
rect 28001 1545 28349 1565
rect 28001 1540 28003 1545
rect 27971 1535 28003 1540
rect 28347 1540 28349 1545
rect 28375 1540 28379 1570
rect 28347 1535 28379 1540
rect 5135 1510 5175 1515
rect 2925 1500 2965 1505
rect 2925 1470 2930 1500
rect 2960 1495 2965 1500
rect 3045 1500 3085 1505
rect 3045 1495 3050 1500
rect 2960 1475 3050 1495
rect 2960 1470 2965 1475
rect 2925 1465 2965 1470
rect 3045 1470 3050 1475
rect 3080 1495 3085 1500
rect 3165 1500 3205 1505
rect 3165 1495 3170 1500
rect 3080 1475 3170 1495
rect 3080 1470 3085 1475
rect 3045 1465 3085 1470
rect 3165 1470 3170 1475
rect 3200 1495 3205 1500
rect 3285 1500 3325 1505
rect 3285 1495 3290 1500
rect 3200 1475 3290 1495
rect 3200 1470 3205 1475
rect 3165 1465 3205 1470
rect 3285 1470 3290 1475
rect 3320 1495 3325 1500
rect 3525 1500 3565 1505
rect 3525 1495 3530 1500
rect 3320 1475 3530 1495
rect 3320 1470 3325 1475
rect 3285 1465 3325 1470
rect 3525 1470 3530 1475
rect 3560 1495 3565 1500
rect 3645 1500 3685 1505
rect 3645 1495 3650 1500
rect 3560 1475 3650 1495
rect 3560 1470 3565 1475
rect 3525 1465 3565 1470
rect 3645 1470 3650 1475
rect 3680 1495 3685 1500
rect 3765 1500 3805 1505
rect 3765 1495 3770 1500
rect 3680 1475 3770 1495
rect 3680 1470 3685 1475
rect 3645 1465 3685 1470
rect 3765 1470 3770 1475
rect 3800 1495 3805 1500
rect 4205 1500 4245 1505
rect 4205 1495 4210 1500
rect 3800 1475 4210 1495
rect 3800 1470 3805 1475
rect 3765 1465 3805 1470
rect 4205 1470 4210 1475
rect 4240 1495 4245 1500
rect 4325 1500 4365 1505
rect 4325 1495 4330 1500
rect 4240 1475 4330 1495
rect 4240 1470 4245 1475
rect 4205 1465 4245 1470
rect 4325 1470 4330 1475
rect 4360 1495 4365 1500
rect 4445 1500 4485 1505
rect 4445 1495 4450 1500
rect 4360 1475 4450 1495
rect 4360 1470 4365 1475
rect 4325 1465 4365 1470
rect 4445 1470 4450 1475
rect 4480 1495 4485 1500
rect 4685 1500 4725 1505
rect 4685 1495 4690 1500
rect 4480 1475 4690 1495
rect 4480 1470 4485 1475
rect 4445 1465 4485 1470
rect 4685 1470 4690 1475
rect 4720 1495 4725 1500
rect 4805 1500 4845 1505
rect 4805 1495 4810 1500
rect 4720 1475 4810 1495
rect 4720 1470 4725 1475
rect 4685 1465 4725 1470
rect 4805 1470 4810 1475
rect 4840 1495 4845 1500
rect 4925 1500 4965 1505
rect 4925 1495 4930 1500
rect 4840 1475 4930 1495
rect 4840 1470 4845 1475
rect 4805 1465 4845 1470
rect 4925 1470 4930 1475
rect 4960 1495 4965 1500
rect 5045 1500 5085 1505
rect 5045 1495 5050 1500
rect 4960 1475 5050 1495
rect 4960 1470 4965 1475
rect 4925 1465 4965 1470
rect 5045 1470 5050 1475
rect 5080 1495 5085 1500
rect 5550 1500 5590 1505
rect 5550 1495 5555 1500
rect 5080 1475 5555 1495
rect 5080 1470 5085 1475
rect 5045 1465 5085 1470
rect 5550 1470 5555 1475
rect 5585 1470 5590 1500
rect 11106 1495 11138 1500
rect 11106 1490 11109 1495
rect 10905 1470 11109 1490
rect 5550 1465 5590 1470
rect 11106 1465 11109 1470
rect 11135 1490 11138 1495
rect 11305 1495 11345 1500
rect 11305 1490 11310 1495
rect 11135 1470 11310 1490
rect 11135 1465 11138 1470
rect 11106 1460 11138 1465
rect 11305 1465 11310 1470
rect 11340 1490 11345 1495
rect 11525 1495 11565 1500
rect 11525 1490 11530 1495
rect 11340 1470 11530 1490
rect 11340 1465 11345 1470
rect 11305 1460 11345 1465
rect 11525 1465 11530 1470
rect 11560 1490 11565 1495
rect 11922 1495 11954 1500
rect 11922 1490 11925 1495
rect 11560 1470 11925 1490
rect 11560 1465 11565 1470
rect 11525 1460 11565 1465
rect 11922 1465 11925 1470
rect 11951 1490 11954 1495
rect 12146 1495 12178 1500
rect 12146 1490 12149 1495
rect 11951 1470 12149 1490
rect 11951 1465 11954 1470
rect 11922 1460 11954 1465
rect 12146 1465 12149 1470
rect 12175 1490 12178 1495
rect 12345 1495 12385 1500
rect 12345 1490 12350 1495
rect 12175 1470 12350 1490
rect 12175 1465 12178 1470
rect 12146 1460 12178 1465
rect 12345 1465 12350 1470
rect 12380 1490 12385 1495
rect 12565 1495 12605 1500
rect 12565 1490 12570 1495
rect 12380 1470 12570 1490
rect 12380 1465 12385 1470
rect 12345 1460 12385 1465
rect 12565 1465 12570 1470
rect 12600 1465 12605 1495
rect 26106 1495 26138 1500
rect 26106 1490 26109 1495
rect 25910 1470 26109 1490
rect 12565 1460 12605 1465
rect 26106 1465 26109 1470
rect 26135 1490 26138 1495
rect 26305 1495 26345 1500
rect 26305 1490 26310 1495
rect 26135 1470 26310 1490
rect 26135 1465 26138 1470
rect 26106 1460 26138 1465
rect 26305 1465 26310 1470
rect 26340 1490 26345 1495
rect 26525 1495 26565 1500
rect 26525 1490 26530 1495
rect 26340 1470 26530 1490
rect 26340 1465 26345 1470
rect 26305 1460 26345 1465
rect 26525 1465 26530 1470
rect 26560 1490 26565 1495
rect 26922 1495 26954 1500
rect 26922 1490 26925 1495
rect 26560 1470 26925 1490
rect 26560 1465 26565 1470
rect 26525 1460 26565 1465
rect 26922 1465 26925 1470
rect 26951 1490 26954 1495
rect 27146 1495 27178 1500
rect 27146 1490 27149 1495
rect 26951 1470 27149 1490
rect 26951 1465 26954 1470
rect 26922 1460 26954 1465
rect 27146 1465 27149 1470
rect 27175 1490 27178 1495
rect 27345 1495 27385 1500
rect 27345 1490 27350 1495
rect 27175 1470 27350 1490
rect 27175 1465 27178 1470
rect 27146 1460 27178 1465
rect 27345 1465 27350 1470
rect 27380 1490 27385 1495
rect 27565 1495 27605 1500
rect 27565 1490 27570 1495
rect 27380 1470 27570 1490
rect 27380 1465 27385 1470
rect 27345 1460 27385 1465
rect 27565 1465 27570 1470
rect 27600 1465 27605 1495
rect 27565 1460 27605 1465
rect 11145 1435 11185 1440
rect 11145 1405 11150 1435
rect 11180 1430 11185 1435
rect 11250 1435 11290 1440
rect 11250 1430 11255 1435
rect 11180 1410 11255 1430
rect 11180 1405 11185 1410
rect 11145 1400 11185 1405
rect 11250 1405 11255 1410
rect 11285 1430 11290 1435
rect 11360 1435 11400 1440
rect 11360 1430 11365 1435
rect 11285 1410 11365 1430
rect 11285 1405 11290 1410
rect 11250 1400 11290 1405
rect 11360 1405 11365 1410
rect 11395 1430 11400 1435
rect 11470 1435 11510 1440
rect 11470 1430 11475 1435
rect 11395 1410 11475 1430
rect 11395 1405 11400 1410
rect 11360 1400 11400 1405
rect 11470 1405 11475 1410
rect 11505 1430 11510 1435
rect 11580 1435 11620 1440
rect 11580 1430 11585 1435
rect 11505 1410 11585 1430
rect 11505 1405 11510 1410
rect 11470 1400 11510 1405
rect 11580 1405 11585 1410
rect 11615 1430 11620 1435
rect 12185 1435 12225 1440
rect 12185 1430 12190 1435
rect 11615 1410 12190 1430
rect 11615 1405 11620 1410
rect 11580 1400 11620 1405
rect 12185 1405 12190 1410
rect 12220 1430 12225 1435
rect 12290 1435 12330 1440
rect 12290 1430 12295 1435
rect 12220 1410 12295 1430
rect 12220 1405 12225 1410
rect 12185 1400 12225 1405
rect 12290 1405 12295 1410
rect 12325 1430 12330 1435
rect 12400 1435 12440 1440
rect 12400 1430 12405 1435
rect 12325 1410 12405 1430
rect 12325 1405 12330 1410
rect 12290 1400 12330 1405
rect 12400 1405 12405 1410
rect 12435 1430 12440 1435
rect 12510 1435 12550 1440
rect 12510 1430 12515 1435
rect 12435 1410 12515 1430
rect 12435 1405 12440 1410
rect 12400 1400 12440 1405
rect 12510 1405 12515 1410
rect 12545 1430 12550 1435
rect 12620 1435 12660 1440
rect 12620 1430 12625 1435
rect 12545 1410 12625 1430
rect 12545 1405 12550 1410
rect 12510 1400 12550 1405
rect 12620 1405 12625 1410
rect 12655 1405 12660 1435
rect 12620 1400 12660 1405
rect 26145 1435 26185 1440
rect 26145 1405 26150 1435
rect 26180 1430 26185 1435
rect 26250 1435 26290 1440
rect 26250 1430 26255 1435
rect 26180 1410 26255 1430
rect 26180 1405 26185 1410
rect 26145 1400 26185 1405
rect 26250 1405 26255 1410
rect 26285 1430 26290 1435
rect 26360 1435 26400 1440
rect 26360 1430 26365 1435
rect 26285 1410 26365 1430
rect 26285 1405 26290 1410
rect 26250 1400 26290 1405
rect 26360 1405 26365 1410
rect 26395 1430 26400 1435
rect 26470 1435 26510 1440
rect 26470 1430 26475 1435
rect 26395 1410 26475 1430
rect 26395 1405 26400 1410
rect 26360 1400 26400 1405
rect 26470 1405 26475 1410
rect 26505 1430 26510 1435
rect 26580 1435 26620 1440
rect 26580 1430 26585 1435
rect 26505 1410 26585 1430
rect 26505 1405 26510 1410
rect 26470 1400 26510 1405
rect 26580 1405 26585 1410
rect 26615 1430 26620 1435
rect 27185 1435 27225 1440
rect 27185 1430 27190 1435
rect 26615 1410 27190 1430
rect 26615 1405 26620 1410
rect 26580 1400 26620 1405
rect 27185 1405 27190 1410
rect 27220 1430 27225 1435
rect 27290 1435 27330 1440
rect 27290 1430 27295 1435
rect 27220 1410 27295 1430
rect 27220 1405 27225 1410
rect 27185 1400 27225 1405
rect 27290 1405 27295 1410
rect 27325 1430 27330 1435
rect 27400 1435 27440 1440
rect 27400 1430 27405 1435
rect 27325 1410 27405 1430
rect 27325 1405 27330 1410
rect 27290 1400 27330 1405
rect 27400 1405 27405 1410
rect 27435 1430 27440 1435
rect 27510 1435 27550 1440
rect 27510 1430 27515 1435
rect 27435 1410 27515 1430
rect 27435 1405 27440 1410
rect 27400 1400 27440 1405
rect 27510 1405 27515 1410
rect 27545 1430 27550 1435
rect 27620 1435 27660 1440
rect 27620 1430 27625 1435
rect 27545 1410 27625 1430
rect 27545 1405 27550 1410
rect 27510 1400 27550 1405
rect 27620 1405 27625 1410
rect 27655 1405 27660 1435
rect 27620 1400 27660 1405
rect 10835 1390 10875 1395
rect 10835 1360 10840 1390
rect 10870 1385 10875 1390
rect 12925 1390 12965 1395
rect 12925 1385 12930 1390
rect 10870 1365 12930 1385
rect 10870 1360 10875 1365
rect 10835 1355 10875 1360
rect 12925 1360 12930 1365
rect 12960 1360 12965 1390
rect 12925 1355 12965 1360
rect 26810 1385 26850 1390
rect 26810 1355 26815 1385
rect 26845 1355 26850 1385
rect 26810 1350 26850 1355
rect 28026 1350 28058 1355
rect 11005 1345 11045 1350
rect 11005 1315 11010 1345
rect 11040 1340 11045 1345
rect 11810 1345 11850 1350
rect 28026 1345 28028 1350
rect 11810 1340 11815 1345
rect 11040 1320 11815 1340
rect 11040 1315 11045 1320
rect 11005 1310 11045 1315
rect 11810 1315 11815 1320
rect 11845 1315 11850 1345
rect 11810 1310 11850 1315
rect 26315 1335 26355 1340
rect 26315 1305 26320 1335
rect 26350 1330 26355 1335
rect 26880 1335 26920 1340
rect 26880 1330 26885 1335
rect 26350 1310 26885 1330
rect 26350 1305 26355 1310
rect 26315 1300 26355 1305
rect 26880 1305 26885 1310
rect 26915 1305 26920 1335
rect 28025 1325 28028 1345
rect 28026 1320 28028 1325
rect 28054 1345 28058 1350
rect 28292 1350 28324 1355
rect 28292 1345 28296 1350
rect 28054 1325 28296 1345
rect 28054 1320 28058 1325
rect 28026 1315 28058 1320
rect 28292 1320 28296 1325
rect 28322 1345 28324 1350
rect 28322 1325 28325 1345
rect 28322 1320 28324 1325
rect 28292 1315 28324 1320
rect 26880 1300 26920 1305
rect 11315 1295 11355 1300
rect 11315 1265 11320 1295
rect 11350 1290 11355 1295
rect 11880 1295 11920 1300
rect 11880 1290 11885 1295
rect 11350 1270 11885 1290
rect 11350 1265 11355 1270
rect 11315 1260 11355 1265
rect 11880 1265 11885 1270
rect 11915 1265 11920 1295
rect 27595 1290 27635 1295
rect 11880 1260 11920 1265
rect 26425 1275 26465 1280
rect 12595 1250 12635 1255
rect 11425 1235 11465 1240
rect 11425 1205 11430 1235
rect 11460 1230 11465 1235
rect 11535 1235 11575 1240
rect 11535 1230 11540 1235
rect 11460 1210 11540 1230
rect 11460 1205 11465 1210
rect 11425 1200 11465 1205
rect 11535 1205 11540 1210
rect 11570 1230 11575 1235
rect 11645 1235 11685 1240
rect 11645 1230 11650 1235
rect 11570 1210 11650 1230
rect 11570 1205 11575 1210
rect 11535 1200 11575 1205
rect 11645 1205 11650 1210
rect 11680 1230 11685 1235
rect 11755 1235 11795 1240
rect 11755 1230 11760 1235
rect 11680 1210 11760 1230
rect 11680 1205 11685 1210
rect 11645 1200 11685 1205
rect 11755 1205 11760 1210
rect 11790 1230 11795 1235
rect 11865 1235 11905 1240
rect 11865 1230 11870 1235
rect 11790 1210 11870 1230
rect 11790 1205 11795 1210
rect 11755 1200 11795 1205
rect 11865 1205 11870 1210
rect 11900 1230 11905 1235
rect 11975 1235 12015 1240
rect 11975 1230 11980 1235
rect 11900 1210 11980 1230
rect 11900 1205 11905 1210
rect 11865 1200 11905 1205
rect 11975 1205 11980 1210
rect 12010 1230 12015 1235
rect 12085 1235 12125 1240
rect 12085 1230 12090 1235
rect 12010 1210 12090 1230
rect 12010 1205 12015 1210
rect 11975 1200 12015 1205
rect 12085 1205 12090 1210
rect 12120 1230 12125 1235
rect 12195 1235 12235 1240
rect 12195 1230 12200 1235
rect 12120 1210 12200 1230
rect 12120 1205 12125 1210
rect 12085 1200 12125 1205
rect 12195 1205 12200 1210
rect 12230 1230 12235 1235
rect 12305 1235 12345 1240
rect 12305 1230 12310 1235
rect 12230 1210 12310 1230
rect 12230 1205 12235 1210
rect 12195 1200 12235 1205
rect 12305 1205 12310 1210
rect 12340 1230 12345 1235
rect 12415 1235 12455 1240
rect 12415 1230 12420 1235
rect 12340 1210 12420 1230
rect 12340 1205 12345 1210
rect 12305 1200 12345 1205
rect 12415 1205 12420 1210
rect 12450 1230 12455 1235
rect 12525 1235 12565 1240
rect 12525 1230 12530 1235
rect 12450 1210 12530 1230
rect 12450 1205 12455 1210
rect 12415 1200 12455 1205
rect 12525 1205 12530 1210
rect 12560 1205 12565 1235
rect 12595 1220 12600 1250
rect 12630 1245 12635 1250
rect 12805 1250 12845 1255
rect 12805 1245 12810 1250
rect 12630 1225 12810 1245
rect 12630 1220 12635 1225
rect 12595 1215 12635 1220
rect 12805 1220 12810 1225
rect 12840 1220 12845 1250
rect 26425 1245 26430 1275
rect 26460 1270 26465 1275
rect 26535 1275 26575 1280
rect 26535 1270 26540 1275
rect 26460 1250 26540 1270
rect 26460 1245 26465 1250
rect 26425 1240 26465 1245
rect 26535 1245 26540 1250
rect 26570 1270 26575 1275
rect 26645 1275 26685 1280
rect 26645 1270 26650 1275
rect 26570 1250 26650 1270
rect 26570 1245 26575 1250
rect 26535 1240 26575 1245
rect 26645 1245 26650 1250
rect 26680 1270 26685 1275
rect 26755 1275 26795 1280
rect 26755 1270 26760 1275
rect 26680 1250 26760 1270
rect 26680 1245 26685 1250
rect 26645 1240 26685 1245
rect 26755 1245 26760 1250
rect 26790 1270 26795 1275
rect 26865 1275 26905 1280
rect 26865 1270 26870 1275
rect 26790 1250 26870 1270
rect 26790 1245 26795 1250
rect 26755 1240 26795 1245
rect 26865 1245 26870 1250
rect 26900 1270 26905 1275
rect 26975 1275 27015 1280
rect 26975 1270 26980 1275
rect 26900 1250 26980 1270
rect 26900 1245 26905 1250
rect 26865 1240 26905 1245
rect 26975 1245 26980 1250
rect 27010 1270 27015 1275
rect 27085 1275 27125 1280
rect 27085 1270 27090 1275
rect 27010 1250 27090 1270
rect 27010 1245 27015 1250
rect 26975 1240 27015 1245
rect 27085 1245 27090 1250
rect 27120 1270 27125 1275
rect 27195 1275 27235 1280
rect 27195 1270 27200 1275
rect 27120 1250 27200 1270
rect 27120 1245 27125 1250
rect 27085 1240 27125 1245
rect 27195 1245 27200 1250
rect 27230 1270 27235 1275
rect 27305 1275 27345 1280
rect 27305 1270 27310 1275
rect 27230 1250 27310 1270
rect 27230 1245 27235 1250
rect 27195 1240 27235 1245
rect 27305 1245 27310 1250
rect 27340 1270 27345 1275
rect 27415 1275 27455 1280
rect 27415 1270 27420 1275
rect 27340 1250 27420 1270
rect 27340 1245 27345 1250
rect 27305 1240 27345 1245
rect 27415 1245 27420 1250
rect 27450 1270 27455 1275
rect 27525 1275 27565 1280
rect 27525 1270 27530 1275
rect 27450 1250 27530 1270
rect 27450 1245 27455 1250
rect 27415 1240 27455 1245
rect 27525 1245 27530 1250
rect 27560 1245 27565 1275
rect 27595 1260 27600 1290
rect 27630 1285 27635 1290
rect 27945 1290 27985 1295
rect 27945 1285 27950 1290
rect 27630 1265 27950 1285
rect 27630 1260 27635 1265
rect 27595 1255 27635 1260
rect 27945 1260 27950 1265
rect 27980 1285 27985 1290
rect 28060 1290 28100 1295
rect 28060 1285 28065 1290
rect 27980 1265 28065 1285
rect 27980 1260 27985 1265
rect 27945 1255 27985 1260
rect 28060 1260 28065 1265
rect 28095 1260 28100 1290
rect 28060 1255 28100 1260
rect 28155 1290 28195 1295
rect 28155 1260 28160 1290
rect 28190 1285 28195 1290
rect 28250 1290 28290 1295
rect 28250 1285 28255 1290
rect 28190 1265 28255 1285
rect 28190 1260 28195 1265
rect 28155 1255 28195 1260
rect 28250 1260 28255 1265
rect 28285 1260 28290 1290
rect 28250 1255 28290 1260
rect 28365 1290 28405 1295
rect 28365 1260 28370 1290
rect 28400 1260 28405 1290
rect 28365 1255 28405 1260
rect 27525 1240 27565 1245
rect 12805 1215 12845 1220
rect 28100 1230 28140 1235
rect 12525 1200 12565 1205
rect 28100 1200 28105 1230
rect 28135 1225 28140 1230
rect 28160 1230 28190 1235
rect 28135 1205 28160 1225
rect 28135 1200 28140 1205
rect 28100 1195 28140 1200
rect 28160 1195 28190 1200
rect 28210 1230 28250 1235
rect 28210 1200 28215 1230
rect 28245 1225 28250 1230
rect 28365 1230 28405 1235
rect 28365 1225 28370 1230
rect 28245 1205 28370 1225
rect 28245 1200 28250 1205
rect 28210 1195 28250 1200
rect 28365 1200 28370 1205
rect 28400 1200 28405 1230
rect 28365 1195 28405 1200
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1180 3415 1185
rect 3985 1185 4025 1190
rect 3985 1180 3990 1185
rect 3410 1160 3990 1180
rect 3410 1155 3415 1160
rect 3375 1150 3415 1155
rect 3985 1155 3990 1160
rect 4020 1180 4025 1185
rect 4595 1185 4635 1190
rect 4595 1180 4600 1185
rect 4020 1160 4600 1180
rect 4020 1155 4025 1160
rect 3985 1150 4025 1155
rect 4595 1155 4600 1160
rect 4630 1180 4635 1185
rect 5465 1185 5505 1190
rect 5465 1180 5470 1185
rect 4630 1160 5470 1180
rect 4630 1155 4635 1160
rect 4595 1150 4635 1155
rect 5465 1155 5470 1160
rect 5500 1155 5505 1185
rect 5465 1150 5505 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1120 2985 1125
rect 3025 1125 3065 1130
rect 3025 1120 3030 1125
rect 2980 1100 3030 1120
rect 2980 1095 2985 1100
rect 2945 1090 2985 1095
rect 3025 1095 3030 1100
rect 3060 1120 3065 1125
rect 3105 1125 3145 1130
rect 3105 1120 3110 1125
rect 3060 1100 3110 1120
rect 3060 1095 3065 1100
rect 3025 1090 3065 1095
rect 3105 1095 3110 1100
rect 3140 1120 3145 1125
rect 3185 1125 3225 1130
rect 3185 1120 3190 1125
rect 3140 1100 3190 1120
rect 3140 1095 3145 1100
rect 3105 1090 3145 1095
rect 3185 1095 3190 1100
rect 3220 1120 3225 1125
rect 3265 1125 3305 1130
rect 3265 1120 3270 1125
rect 3220 1100 3270 1120
rect 3220 1095 3225 1100
rect 3185 1090 3225 1095
rect 3265 1095 3270 1100
rect 3300 1120 3305 1125
rect 3345 1125 3385 1130
rect 3345 1120 3350 1125
rect 3300 1100 3350 1120
rect 3300 1095 3305 1100
rect 3265 1090 3305 1095
rect 3345 1095 3350 1100
rect 3380 1120 3385 1125
rect 3425 1125 3465 1130
rect 3425 1120 3430 1125
rect 3380 1100 3430 1120
rect 3380 1095 3385 1100
rect 3345 1090 3385 1095
rect 3425 1095 3430 1100
rect 3460 1120 3465 1125
rect 3505 1125 3545 1130
rect 3505 1120 3510 1125
rect 3460 1100 3510 1120
rect 3460 1095 3465 1100
rect 3425 1090 3465 1095
rect 3505 1095 3510 1100
rect 3540 1120 3545 1125
rect 3585 1125 3625 1130
rect 3585 1120 3590 1125
rect 3540 1100 3590 1120
rect 3540 1095 3545 1100
rect 3505 1090 3545 1095
rect 3585 1095 3590 1100
rect 3620 1120 3625 1125
rect 3665 1125 3705 1130
rect 3665 1120 3670 1125
rect 3620 1100 3670 1120
rect 3620 1095 3625 1100
rect 3585 1090 3625 1095
rect 3665 1095 3670 1100
rect 3700 1120 3705 1125
rect 3745 1125 3785 1130
rect 3745 1120 3750 1125
rect 3700 1100 3750 1120
rect 3700 1095 3705 1100
rect 3665 1090 3705 1095
rect 3745 1095 3750 1100
rect 3780 1120 3785 1125
rect 3825 1125 3865 1130
rect 3825 1120 3830 1125
rect 3780 1100 3830 1120
rect 3780 1095 3785 1100
rect 3745 1090 3785 1095
rect 3825 1095 3830 1100
rect 3860 1120 3865 1125
rect 3905 1125 3945 1130
rect 3905 1120 3910 1125
rect 3860 1100 3910 1120
rect 3860 1095 3865 1100
rect 3825 1090 3865 1095
rect 3905 1095 3910 1100
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1120 4025 1125
rect 4065 1125 4105 1130
rect 4065 1120 4070 1125
rect 4020 1100 4070 1120
rect 4020 1095 4025 1100
rect 3985 1090 4025 1095
rect 4065 1095 4070 1100
rect 4100 1120 4105 1125
rect 4145 1125 4185 1130
rect 4145 1120 4150 1125
rect 4100 1100 4150 1120
rect 4100 1095 4105 1100
rect 4065 1090 4105 1095
rect 4145 1095 4150 1100
rect 4180 1120 4185 1125
rect 4225 1125 4265 1130
rect 4225 1120 4230 1125
rect 4180 1100 4230 1120
rect 4180 1095 4185 1100
rect 4145 1090 4185 1095
rect 4225 1095 4230 1100
rect 4260 1120 4265 1125
rect 4305 1125 4345 1130
rect 4305 1120 4310 1125
rect 4260 1100 4310 1120
rect 4260 1095 4265 1100
rect 4225 1090 4265 1095
rect 4305 1095 4310 1100
rect 4340 1120 4345 1125
rect 4385 1125 4425 1130
rect 4385 1120 4390 1125
rect 4340 1100 4390 1120
rect 4340 1095 4345 1100
rect 4305 1090 4345 1095
rect 4385 1095 4390 1100
rect 4420 1120 4425 1125
rect 4465 1125 4505 1130
rect 4465 1120 4470 1125
rect 4420 1100 4470 1120
rect 4420 1095 4425 1100
rect 4385 1090 4425 1095
rect 4465 1095 4470 1100
rect 4500 1120 4505 1125
rect 4545 1125 4585 1130
rect 4545 1120 4550 1125
rect 4500 1100 4550 1120
rect 4500 1095 4505 1100
rect 4465 1090 4505 1095
rect 4545 1095 4550 1100
rect 4580 1120 4585 1125
rect 4625 1125 4665 1130
rect 4625 1120 4630 1125
rect 4580 1100 4630 1120
rect 4580 1095 4585 1100
rect 4545 1090 4585 1095
rect 4625 1095 4630 1100
rect 4660 1120 4665 1125
rect 4705 1125 4745 1130
rect 4705 1120 4710 1125
rect 4660 1100 4710 1120
rect 4660 1095 4665 1100
rect 4625 1090 4665 1095
rect 4705 1095 4710 1100
rect 4740 1120 4745 1125
rect 4785 1125 4825 1130
rect 4785 1120 4790 1125
rect 4740 1100 4790 1120
rect 4740 1095 4745 1100
rect 4705 1090 4745 1095
rect 4785 1095 4790 1100
rect 4820 1120 4825 1125
rect 4865 1125 4905 1130
rect 4865 1120 4870 1125
rect 4820 1100 4870 1120
rect 4820 1095 4825 1100
rect 4785 1090 4825 1095
rect 4865 1095 4870 1100
rect 4900 1120 4905 1125
rect 4945 1125 4985 1130
rect 4945 1120 4950 1125
rect 4900 1100 4950 1120
rect 4900 1095 4905 1100
rect 4865 1090 4905 1095
rect 4945 1095 4950 1100
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1035 2660 1040
rect 2905 1040 2945 1045
rect 2905 1035 2910 1040
rect 2655 1015 2910 1035
rect 2655 1010 2660 1015
rect 2620 1005 2660 1010
rect 2905 1010 2910 1015
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1035 5150 1040
rect 5465 1040 5505 1045
rect 5465 1035 5470 1040
rect 5145 1015 5470 1035
rect 5145 1010 5150 1015
rect 5110 1005 5150 1010
rect 5465 1010 5470 1015
rect 5500 1010 5505 1040
rect 5465 1005 5505 1010
rect 26165 955 26205 960
rect 10355 935 10395 940
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 925 3035 930
rect 3175 930 3215 935
rect 3175 925 3180 930
rect 3030 905 3180 925
rect 3030 900 3035 905
rect 2995 895 3035 900
rect 3175 900 3180 905
rect 3210 925 3215 930
rect 3355 930 3395 935
rect 3355 925 3360 930
rect 3210 905 3360 925
rect 3210 900 3215 905
rect 3175 895 3215 900
rect 3355 900 3360 905
rect 3390 925 3395 930
rect 3535 930 3575 935
rect 3535 925 3540 930
rect 3390 905 3540 925
rect 3390 900 3395 905
rect 3355 895 3395 900
rect 3535 900 3540 905
rect 3570 925 3575 930
rect 3715 930 3755 935
rect 3715 925 3720 930
rect 3570 905 3720 925
rect 3570 900 3575 905
rect 3535 895 3575 900
rect 3715 900 3720 905
rect 3750 925 3755 930
rect 3895 930 3935 935
rect 3895 925 3900 930
rect 3750 905 3900 925
rect 3750 900 3755 905
rect 3715 895 3755 900
rect 3895 900 3900 905
rect 3930 925 3935 930
rect 4075 930 4115 935
rect 4075 925 4080 930
rect 3930 905 4080 925
rect 3930 900 3935 905
rect 3895 895 3935 900
rect 4075 900 4080 905
rect 4110 925 4115 930
rect 4255 930 4295 935
rect 4255 925 4260 930
rect 4110 905 4260 925
rect 4110 900 4115 905
rect 4075 895 4115 900
rect 4255 900 4260 905
rect 4290 925 4295 930
rect 4435 930 4475 935
rect 4435 925 4440 930
rect 4290 905 4440 925
rect 4290 900 4295 905
rect 4255 895 4295 900
rect 4435 900 4440 905
rect 4470 925 4475 930
rect 4615 930 4655 935
rect 4615 925 4620 930
rect 4470 905 4620 925
rect 4470 900 4475 905
rect 4435 895 4475 900
rect 4615 900 4620 905
rect 4650 925 4655 930
rect 4795 930 4835 935
rect 4795 925 4800 930
rect 4650 905 4800 925
rect 4650 900 4655 905
rect 4615 895 4655 900
rect 4795 900 4800 905
rect 4830 925 4835 930
rect 4975 930 5015 935
rect 4975 925 4980 930
rect 4830 905 4980 925
rect 4830 900 4835 905
rect 4795 895 4835 900
rect 4975 900 4980 905
rect 5010 925 5015 930
rect 5465 930 5505 935
rect 5465 925 5470 930
rect 5010 905 5470 925
rect 5010 900 5015 905
rect 4975 895 5015 900
rect 5465 900 5470 905
rect 5500 900 5505 930
rect 10355 905 10360 935
rect 10390 930 10395 935
rect 10555 935 10595 940
rect 10555 930 10560 935
rect 10390 910 10560 930
rect 10390 905 10395 910
rect 10355 900 10395 905
rect 10555 905 10560 910
rect 10590 905 10595 935
rect 13205 935 13245 940
rect 10555 900 10595 905
rect 11165 915 11205 920
rect 5465 895 5505 900
rect 11165 885 11170 915
rect 11200 910 11205 915
rect 11260 915 11300 920
rect 11260 910 11265 915
rect 11200 890 11265 910
rect 11200 885 11205 890
rect 11165 880 11205 885
rect 11260 885 11265 890
rect 11295 910 11300 915
rect 11370 915 11410 920
rect 11370 910 11375 915
rect 11295 890 11375 910
rect 11295 885 11300 890
rect 11260 880 11300 885
rect 11370 885 11375 890
rect 11405 910 11410 915
rect 11480 915 11520 920
rect 11480 910 11485 915
rect 11405 890 11485 910
rect 11405 885 11410 890
rect 11370 880 11410 885
rect 11480 885 11485 890
rect 11515 910 11520 915
rect 11590 915 11630 920
rect 11590 910 11595 915
rect 11515 890 11595 910
rect 11515 885 11520 890
rect 11480 880 11520 885
rect 11590 885 11595 890
rect 11625 910 11630 915
rect 11700 915 11740 920
rect 11700 910 11705 915
rect 11625 890 11705 910
rect 11625 885 11630 890
rect 11590 880 11630 885
rect 11700 885 11705 890
rect 11735 910 11740 915
rect 11810 915 11850 920
rect 11810 910 11815 915
rect 11735 890 11815 910
rect 11735 885 11740 890
rect 11700 880 11740 885
rect 11810 885 11815 890
rect 11845 910 11850 915
rect 11920 915 11960 920
rect 11920 910 11925 915
rect 11845 890 11925 910
rect 11845 885 11850 890
rect 11810 880 11850 885
rect 11920 885 11925 890
rect 11955 910 11960 915
rect 12030 915 12070 920
rect 12030 910 12035 915
rect 11955 890 12035 910
rect 11955 885 11960 890
rect 11920 880 11960 885
rect 12030 885 12035 890
rect 12065 910 12070 915
rect 12140 915 12180 920
rect 12140 910 12145 915
rect 12065 890 12145 910
rect 12065 885 12070 890
rect 12030 880 12070 885
rect 12140 885 12145 890
rect 12175 910 12180 915
rect 12250 915 12290 920
rect 12250 910 12255 915
rect 12175 890 12255 910
rect 12175 885 12180 890
rect 12140 880 12180 885
rect 12250 885 12255 890
rect 12285 910 12290 915
rect 12360 915 12400 920
rect 12360 910 12365 915
rect 12285 890 12365 910
rect 12285 885 12290 890
rect 12250 880 12290 885
rect 12360 885 12365 890
rect 12395 910 12400 915
rect 12470 915 12510 920
rect 12470 910 12475 915
rect 12395 890 12475 910
rect 12395 885 12400 890
rect 12360 880 12400 885
rect 12470 885 12475 890
rect 12505 910 12510 915
rect 12620 915 12660 920
rect 12620 910 12625 915
rect 12505 890 12625 910
rect 12505 885 12510 890
rect 12470 880 12510 885
rect 12620 885 12625 890
rect 12655 885 12660 915
rect 13205 905 13210 935
rect 13240 930 13245 935
rect 13405 935 13445 940
rect 13405 930 13410 935
rect 13240 910 13410 930
rect 13240 905 13245 910
rect 13205 900 13245 905
rect 13405 905 13410 910
rect 13440 905 13445 935
rect 26165 925 26170 955
rect 26200 950 26205 955
rect 26260 955 26300 960
rect 26260 950 26265 955
rect 26200 930 26265 950
rect 26200 925 26205 930
rect 26165 920 26205 925
rect 26260 925 26265 930
rect 26295 950 26300 955
rect 26370 955 26410 960
rect 26370 950 26375 955
rect 26295 930 26375 950
rect 26295 925 26300 930
rect 26260 920 26300 925
rect 26370 925 26375 930
rect 26405 950 26410 955
rect 26480 955 26520 960
rect 26480 950 26485 955
rect 26405 930 26485 950
rect 26405 925 26410 930
rect 26370 920 26410 925
rect 26480 925 26485 930
rect 26515 950 26520 955
rect 26590 955 26630 960
rect 26590 950 26595 955
rect 26515 930 26595 950
rect 26515 925 26520 930
rect 26480 920 26520 925
rect 26590 925 26595 930
rect 26625 950 26630 955
rect 26700 955 26740 960
rect 26700 950 26705 955
rect 26625 930 26705 950
rect 26625 925 26630 930
rect 26590 920 26630 925
rect 26700 925 26705 930
rect 26735 950 26740 955
rect 26810 955 26850 960
rect 26810 950 26815 955
rect 26735 930 26815 950
rect 26735 925 26740 930
rect 26700 920 26740 925
rect 26810 925 26815 930
rect 26845 950 26850 955
rect 26920 955 26960 960
rect 26920 950 26925 955
rect 26845 930 26925 950
rect 26845 925 26850 930
rect 26810 920 26850 925
rect 26920 925 26925 930
rect 26955 950 26960 955
rect 27030 955 27070 960
rect 27030 950 27035 955
rect 26955 930 27035 950
rect 26955 925 26960 930
rect 26920 920 26960 925
rect 27030 925 27035 930
rect 27065 950 27070 955
rect 27140 955 27180 960
rect 27140 950 27145 955
rect 27065 930 27145 950
rect 27065 925 27070 930
rect 27030 920 27070 925
rect 27140 925 27145 930
rect 27175 950 27180 955
rect 27250 955 27290 960
rect 27250 950 27255 955
rect 27175 930 27255 950
rect 27175 925 27180 930
rect 27140 920 27180 925
rect 27250 925 27255 930
rect 27285 950 27290 955
rect 27360 955 27400 960
rect 27360 950 27365 955
rect 27285 930 27365 950
rect 27285 925 27290 930
rect 27250 920 27290 925
rect 27360 925 27365 930
rect 27395 950 27400 955
rect 27470 955 27510 960
rect 27470 950 27475 955
rect 27395 930 27475 950
rect 27395 925 27400 930
rect 27360 920 27400 925
rect 27470 925 27475 930
rect 27505 950 27510 955
rect 27620 955 27660 960
rect 27620 950 27625 955
rect 27505 930 27625 950
rect 27505 925 27510 930
rect 27470 920 27510 925
rect 27620 925 27625 930
rect 27655 925 27660 955
rect 27620 920 27660 925
rect 13405 900 13445 905
rect 12620 880 12660 885
rect 11935 860 11975 865
rect 11005 855 11045 860
rect 11005 825 11010 855
rect 11040 850 11045 855
rect 11495 855 11535 860
rect 11495 850 11500 855
rect 11040 830 11500 850
rect 11040 825 11045 830
rect 11005 820 11045 825
rect 11495 825 11500 830
rect 11530 825 11535 855
rect 11935 830 11940 860
rect 11970 855 11975 860
rect 12155 860 12195 865
rect 12155 855 12160 860
rect 11970 835 12160 855
rect 11970 830 11975 835
rect 11935 825 11975 830
rect 12155 830 12160 835
rect 12190 855 12195 860
rect 12375 860 12415 865
rect 12375 855 12380 860
rect 12190 835 12380 855
rect 12190 830 12195 835
rect 12155 825 12195 830
rect 12375 830 12380 835
rect 12410 855 12415 860
rect 12860 860 12900 865
rect 12860 855 12865 860
rect 12410 835 12865 855
rect 12410 830 12415 835
rect 12375 825 12415 830
rect 12860 830 12865 835
rect 12895 830 12900 860
rect 12860 825 12900 830
rect 11495 820 11535 825
rect 12045 800 12085 805
rect 10950 795 10990 800
rect 10950 765 10955 795
rect 10985 790 10990 795
rect 11305 795 11345 800
rect 11305 790 11310 795
rect 10985 770 11310 790
rect 10985 765 10990 770
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 755 2560 760
rect 3130 760 3170 765
rect 3130 755 3135 760
rect 2555 735 3135 755
rect 2555 730 2560 735
rect 2520 725 2560 730
rect 3130 730 3135 735
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 755 3665 760
rect 3985 760 4025 765
rect 3985 755 3990 760
rect 3660 735 3990 755
rect 3660 730 3665 735
rect 3625 725 3665 730
rect 3985 730 3990 735
rect 4020 755 4025 760
rect 4345 760 4385 765
rect 4345 755 4350 760
rect 4020 735 4350 755
rect 4020 730 4025 735
rect 3985 725 4025 730
rect 4345 730 4350 735
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 755 4565 760
rect 4705 760 4745 765
rect 4705 755 4710 760
rect 4560 735 4710 755
rect 4560 730 4565 735
rect 4525 725 4565 730
rect 4705 730 4710 735
rect 4740 755 4745 760
rect 4885 760 4925 765
rect 10950 760 10990 765
rect 11305 765 11310 770
rect 11340 790 11345 795
rect 11375 795 11415 800
rect 11375 790 11380 795
rect 11340 770 11380 790
rect 11340 765 11345 770
rect 11305 760 11345 765
rect 11375 765 11380 770
rect 11410 790 11415 795
rect 11445 795 11485 800
rect 11445 790 11450 795
rect 11410 770 11450 790
rect 11410 765 11415 770
rect 11375 760 11415 765
rect 11445 765 11450 770
rect 11480 765 11485 795
rect 12045 770 12050 800
rect 12080 795 12085 800
rect 12265 800 12305 805
rect 12265 795 12270 800
rect 12080 775 12270 795
rect 12080 770 12085 775
rect 12045 765 12085 770
rect 12265 770 12270 775
rect 12300 795 12305 800
rect 12485 800 12525 805
rect 12485 795 12490 800
rect 12300 775 12490 795
rect 12300 770 12305 775
rect 12265 765 12305 770
rect 12485 770 12490 775
rect 12520 795 12525 800
rect 12805 800 12845 805
rect 12805 795 12810 800
rect 12520 775 12810 795
rect 12520 770 12525 775
rect 12485 765 12525 770
rect 12805 770 12810 775
rect 12840 770 12845 800
rect 12805 765 12845 770
rect 11445 760 11485 765
rect 4885 755 4890 760
rect 4740 735 4890 755
rect 4740 730 4745 735
rect 4705 725 4745 730
rect 4885 730 4890 735
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 700 3485 705
rect 3805 705 3845 710
rect 3805 700 3810 705
rect 3480 680 3810 700
rect 3480 675 3485 680
rect 3445 670 3485 675
rect 3805 675 3810 680
rect 3840 700 3845 705
rect 4165 705 4205 710
rect 4165 700 4170 705
rect 3840 680 4170 700
rect 3840 675 3845 680
rect 3805 670 3845 675
rect 4165 675 4170 680
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 11990 680 12030 685
rect 11990 650 11995 680
rect 12025 675 12030 680
rect 12100 680 12140 685
rect 12100 675 12105 680
rect 12025 655 12105 675
rect 12025 650 12030 655
rect 11990 645 12030 650
rect 12100 650 12105 655
rect 12135 675 12140 680
rect 12210 680 12250 685
rect 12210 675 12215 680
rect 12135 655 12215 675
rect 12135 650 12140 655
rect 12100 645 12140 650
rect 12210 650 12215 655
rect 12245 675 12250 680
rect 12320 680 12360 685
rect 12320 675 12325 680
rect 12245 655 12325 675
rect 12245 650 12250 655
rect 12210 645 12250 650
rect 12320 650 12325 655
rect 12355 675 12360 680
rect 12430 680 12470 685
rect 12430 675 12435 680
rect 12355 655 12435 675
rect 12355 650 12360 655
rect 12320 645 12360 650
rect 12430 650 12435 655
rect 12465 650 12470 680
rect 12430 645 12470 650
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 11340 -1375 11380 -1370
rect 11340 -1405 11345 -1375
rect 11375 -1380 11380 -1375
rect 11460 -1375 11500 -1370
rect 11460 -1380 11465 -1375
rect 11375 -1400 11465 -1380
rect 11375 -1405 11380 -1400
rect 11340 -1410 11380 -1405
rect 11460 -1405 11465 -1400
rect 11495 -1380 11500 -1375
rect 11580 -1375 11620 -1370
rect 11580 -1380 11585 -1375
rect 11495 -1400 11585 -1380
rect 11495 -1405 11500 -1400
rect 11460 -1410 11500 -1405
rect 11580 -1405 11585 -1400
rect 11615 -1380 11620 -1375
rect 11700 -1375 11740 -1370
rect 11700 -1380 11705 -1375
rect 11615 -1400 11705 -1380
rect 11615 -1405 11620 -1400
rect 11580 -1410 11620 -1405
rect 11700 -1405 11705 -1400
rect 11735 -1380 11740 -1375
rect 11820 -1375 11860 -1370
rect 11820 -1380 11825 -1375
rect 11735 -1400 11825 -1380
rect 11735 -1405 11740 -1400
rect 11700 -1410 11740 -1405
rect 11820 -1405 11825 -1400
rect 11855 -1380 11860 -1375
rect 11940 -1375 11980 -1370
rect 11940 -1380 11945 -1375
rect 11855 -1400 11945 -1380
rect 11855 -1405 11860 -1400
rect 11820 -1410 11860 -1405
rect 11940 -1405 11945 -1400
rect 11975 -1380 11980 -1375
rect 12060 -1375 12100 -1370
rect 12060 -1380 12065 -1375
rect 11975 -1400 12065 -1380
rect 11975 -1405 11980 -1400
rect 11940 -1410 11980 -1405
rect 12060 -1405 12065 -1400
rect 12095 -1380 12100 -1375
rect 12180 -1375 12220 -1370
rect 12180 -1380 12185 -1375
rect 12095 -1400 12185 -1380
rect 12095 -1405 12100 -1400
rect 12060 -1410 12100 -1405
rect 12180 -1405 12185 -1400
rect 12215 -1380 12220 -1375
rect 12300 -1375 12340 -1370
rect 12300 -1380 12305 -1375
rect 12215 -1400 12305 -1380
rect 12215 -1405 12220 -1400
rect 12180 -1410 12220 -1405
rect 12300 -1405 12305 -1400
rect 12335 -1380 12340 -1375
rect 12420 -1375 12460 -1370
rect 12420 -1380 12425 -1375
rect 12335 -1400 12425 -1380
rect 12335 -1405 12340 -1400
rect 12300 -1410 12340 -1405
rect 12420 -1405 12425 -1400
rect 12455 -1405 12460 -1375
rect 12420 -1410 12460 -1405
rect 10580 -1790 10620 -1785
rect 10580 -1820 10585 -1790
rect 10615 -1795 10620 -1790
rect 10980 -1790 11015 -1785
rect 10980 -1795 10985 -1790
rect 10615 -1815 10985 -1795
rect 10615 -1820 10620 -1815
rect 10580 -1825 10620 -1820
rect 10980 -1820 10985 -1815
rect 10980 -1825 11015 -1820
rect 10900 -1845 10940 -1840
rect 10900 -1875 10905 -1845
rect 10935 -1850 10940 -1845
rect 11823 -1845 11857 -1840
rect 11823 -1850 11826 -1845
rect 10935 -1870 11826 -1850
rect 10935 -1875 10940 -1870
rect 10900 -1880 10940 -1875
rect 11823 -1875 11826 -1870
rect 11854 -1875 11857 -1845
rect 11823 -1880 11857 -1875
rect 11280 -1900 11320 -1895
rect 11280 -1930 11285 -1900
rect 11315 -1905 11320 -1900
rect 11520 -1900 11560 -1895
rect 11520 -1905 11525 -1900
rect 11315 -1925 11525 -1905
rect 11315 -1930 11320 -1925
rect 11280 -1935 11320 -1930
rect 11520 -1930 11525 -1925
rect 11555 -1905 11560 -1900
rect 11760 -1900 11800 -1895
rect 11760 -1905 11765 -1900
rect 11555 -1925 11765 -1905
rect 11555 -1930 11560 -1925
rect 11520 -1935 11560 -1930
rect 11760 -1930 11765 -1925
rect 11795 -1905 11800 -1900
rect 12000 -1900 12040 -1895
rect 12000 -1905 12005 -1900
rect 11795 -1925 12005 -1905
rect 11795 -1930 11800 -1925
rect 11760 -1935 11800 -1930
rect 12000 -1930 12005 -1925
rect 12035 -1905 12040 -1900
rect 12240 -1900 12280 -1895
rect 12240 -1905 12245 -1900
rect 12035 -1925 12245 -1905
rect 12035 -1930 12040 -1925
rect 12000 -1935 12040 -1930
rect 12240 -1930 12245 -1925
rect 12275 -1905 12280 -1900
rect 12480 -1900 12520 -1895
rect 12480 -1905 12485 -1900
rect 12275 -1925 12485 -1905
rect 12275 -1930 12280 -1925
rect 12240 -1935 12280 -1930
rect 12480 -1930 12485 -1925
rect 12515 -1930 12520 -1900
rect 12480 -1935 12520 -1930
rect 11400 -1945 11440 -1940
rect 11400 -1975 11405 -1945
rect 11435 -1950 11440 -1945
rect 11640 -1945 11680 -1940
rect 11640 -1950 11645 -1945
rect 11435 -1970 11645 -1950
rect 11435 -1975 11440 -1970
rect 11400 -1980 11440 -1975
rect 11640 -1975 11645 -1970
rect 11675 -1950 11680 -1945
rect 11880 -1945 11920 -1940
rect 11880 -1950 11885 -1945
rect 11675 -1970 11885 -1950
rect 11675 -1975 11680 -1970
rect 11640 -1980 11680 -1975
rect 11880 -1975 11885 -1970
rect 11915 -1950 11920 -1945
rect 12120 -1945 12160 -1940
rect 12120 -1950 12125 -1945
rect 11915 -1970 12125 -1950
rect 11915 -1975 11920 -1970
rect 11880 -1980 11920 -1975
rect 12120 -1975 12125 -1970
rect 12155 -1950 12160 -1945
rect 12360 -1945 12400 -1940
rect 12360 -1950 12365 -1945
rect 12155 -1970 12365 -1950
rect 12155 -1975 12160 -1970
rect 12120 -1980 12160 -1975
rect 12360 -1975 12365 -1970
rect 12395 -1975 12400 -1945
rect 12360 -1980 12400 -1975
rect 12950 -1965 12990 -1960
rect 12950 -1995 12955 -1965
rect 12985 -1970 12990 -1965
rect 13060 -1965 13100 -1960
rect 13060 -1970 13065 -1965
rect 12985 -1990 13065 -1970
rect 12985 -1995 12990 -1990
rect 11340 -2000 11380 -1995
rect 11340 -2030 11345 -2000
rect 11375 -2005 11380 -2000
rect 11400 -2000 11440 -1995
rect 11400 -2005 11405 -2000
rect 11375 -2025 11405 -2005
rect 11375 -2030 11380 -2025
rect 11340 -2035 11380 -2030
rect 11400 -2030 11405 -2025
rect 11435 -2005 11440 -2000
rect 11580 -2000 11620 -1995
rect 11580 -2005 11585 -2000
rect 11435 -2025 11585 -2005
rect 11435 -2030 11440 -2025
rect 11400 -2035 11440 -2030
rect 11580 -2030 11585 -2025
rect 11615 -2005 11620 -2000
rect 11820 -2000 11860 -1995
rect 11820 -2005 11825 -2000
rect 11615 -2025 11825 -2005
rect 11615 -2030 11620 -2025
rect 11580 -2035 11620 -2030
rect 11820 -2030 11825 -2025
rect 11855 -2005 11860 -2000
rect 12060 -2000 12100 -1995
rect 12060 -2005 12065 -2000
rect 11855 -2025 12065 -2005
rect 11855 -2030 11860 -2025
rect 11820 -2035 11860 -2030
rect 12060 -2030 12065 -2025
rect 12095 -2005 12100 -2000
rect 12300 -2000 12340 -1995
rect 12950 -2000 12990 -1995
rect 13060 -1995 13065 -1990
rect 13095 -1970 13100 -1965
rect 13170 -1965 13210 -1960
rect 13170 -1970 13175 -1965
rect 13095 -1990 13175 -1970
rect 13095 -1995 13100 -1990
rect 13060 -2000 13100 -1995
rect 13170 -1995 13175 -1990
rect 13205 -1970 13210 -1965
rect 13280 -1965 13320 -1960
rect 13280 -1970 13285 -1965
rect 13205 -1990 13285 -1970
rect 13205 -1995 13210 -1990
rect 13170 -2000 13210 -1995
rect 13280 -1995 13285 -1990
rect 13315 -1970 13320 -1965
rect 13390 -1965 13430 -1960
rect 13390 -1970 13395 -1965
rect 13315 -1990 13395 -1970
rect 13315 -1995 13320 -1990
rect 13280 -2000 13320 -1995
rect 13390 -1995 13395 -1990
rect 13425 -1970 13430 -1965
rect 13500 -1965 13540 -1960
rect 13500 -1970 13505 -1965
rect 13425 -1990 13505 -1970
rect 13425 -1995 13430 -1990
rect 13390 -2000 13430 -1995
rect 13500 -1995 13505 -1990
rect 13535 -1970 13540 -1965
rect 13610 -1965 13650 -1960
rect 13610 -1970 13615 -1965
rect 13535 -1990 13615 -1970
rect 13535 -1995 13540 -1990
rect 13500 -2000 13540 -1995
rect 13610 -1995 13615 -1990
rect 13645 -1970 13650 -1965
rect 13720 -1965 13760 -1960
rect 13720 -1970 13725 -1965
rect 13645 -1990 13725 -1970
rect 13645 -1995 13650 -1990
rect 13610 -2000 13650 -1995
rect 13720 -1995 13725 -1990
rect 13755 -1970 13760 -1965
rect 13830 -1965 13870 -1960
rect 13830 -1970 13835 -1965
rect 13755 -1990 13835 -1970
rect 13755 -1995 13760 -1990
rect 13720 -2000 13760 -1995
rect 13830 -1995 13835 -1990
rect 13865 -1970 13870 -1965
rect 13940 -1965 13980 -1960
rect 13940 -1970 13945 -1965
rect 13865 -1990 13945 -1970
rect 13865 -1995 13870 -1990
rect 13830 -2000 13870 -1995
rect 13940 -1995 13945 -1990
rect 13975 -1970 13980 -1965
rect 14050 -1965 14090 -1960
rect 14050 -1970 14055 -1965
rect 13975 -1990 14055 -1970
rect 13975 -1995 13980 -1990
rect 13940 -2000 13980 -1995
rect 14050 -1995 14055 -1990
rect 14085 -1995 14090 -1965
rect 14050 -2000 14090 -1995
rect 12300 -2005 12305 -2000
rect 12095 -2025 12305 -2005
rect 12095 -2030 12100 -2025
rect 12060 -2035 12100 -2030
rect 12300 -2030 12305 -2025
rect 12335 -2030 12340 -2000
rect 12300 -2035 12340 -2030
rect 11460 -2055 11500 -2050
rect 11460 -2085 11465 -2055
rect 11495 -2060 11500 -2055
rect 11700 -2055 11740 -2050
rect 11700 -2060 11705 -2055
rect 11495 -2080 11705 -2060
rect 11495 -2085 11500 -2080
rect 11460 -2090 11500 -2085
rect 11700 -2085 11705 -2080
rect 11735 -2060 11740 -2055
rect 11940 -2055 11980 -2050
rect 11940 -2060 11945 -2055
rect 11735 -2080 11945 -2060
rect 11735 -2085 11740 -2080
rect 11700 -2090 11740 -2085
rect 11940 -2085 11945 -2080
rect 11975 -2060 11980 -2055
rect 12180 -2055 12220 -2050
rect 12180 -2060 12185 -2055
rect 11975 -2080 12185 -2060
rect 11975 -2085 11980 -2080
rect 11940 -2090 11980 -2085
rect 12180 -2085 12185 -2080
rect 12215 -2060 12220 -2055
rect 12420 -2055 12460 -2050
rect 12420 -2060 12425 -2055
rect 12215 -2080 12425 -2060
rect 12215 -2085 12220 -2080
rect 12180 -2090 12220 -2085
rect 12420 -2085 12425 -2080
rect 12455 -2060 12460 -2055
rect 12480 -2055 12520 -2050
rect 12480 -2060 12485 -2055
rect 12455 -2080 12485 -2060
rect 12455 -2085 12460 -2080
rect 12420 -2090 12460 -2085
rect 12480 -2085 12485 -2080
rect 12515 -2085 12520 -2055
rect 12480 -2090 12520 -2085
rect 12690 -2270 12730 -2265
rect 12690 -2300 12695 -2270
rect 12725 -2275 12730 -2270
rect 12725 -2295 12785 -2275
rect 12725 -2300 12730 -2295
rect 12690 -2305 12730 -2300
rect 13005 -2335 13045 -2330
rect 13005 -2365 13010 -2335
rect 13040 -2340 13045 -2335
rect 13115 -2335 13155 -2330
rect 13115 -2340 13120 -2335
rect 13040 -2360 13120 -2340
rect 13040 -2365 13045 -2360
rect 13005 -2370 13045 -2365
rect 13115 -2365 13120 -2360
rect 13150 -2340 13155 -2335
rect 13225 -2335 13265 -2330
rect 13225 -2340 13230 -2335
rect 13150 -2360 13230 -2340
rect 13150 -2365 13155 -2360
rect 13115 -2370 13155 -2365
rect 13225 -2365 13230 -2360
rect 13260 -2340 13265 -2335
rect 13335 -2335 13375 -2330
rect 13335 -2340 13340 -2335
rect 13260 -2360 13340 -2340
rect 13260 -2365 13265 -2360
rect 13225 -2370 13265 -2365
rect 13335 -2365 13340 -2360
rect 13370 -2340 13375 -2335
rect 13445 -2335 13485 -2330
rect 13445 -2340 13450 -2335
rect 13370 -2360 13450 -2340
rect 13370 -2365 13375 -2360
rect 13335 -2370 13375 -2365
rect 13445 -2365 13450 -2360
rect 13480 -2340 13485 -2335
rect 13555 -2335 13595 -2330
rect 13555 -2340 13560 -2335
rect 13480 -2360 13560 -2340
rect 13480 -2365 13485 -2360
rect 13445 -2370 13485 -2365
rect 13555 -2365 13560 -2360
rect 13590 -2340 13595 -2335
rect 13665 -2335 13705 -2330
rect 13665 -2340 13670 -2335
rect 13590 -2360 13670 -2340
rect 13590 -2365 13595 -2360
rect 13555 -2370 13595 -2365
rect 13665 -2365 13670 -2360
rect 13700 -2340 13705 -2335
rect 13775 -2335 13815 -2330
rect 13775 -2340 13780 -2335
rect 13700 -2360 13780 -2340
rect 13700 -2365 13705 -2360
rect 13665 -2370 13705 -2365
rect 13775 -2365 13780 -2360
rect 13810 -2340 13815 -2335
rect 13885 -2335 13925 -2330
rect 13885 -2340 13890 -2335
rect 13810 -2360 13890 -2340
rect 13810 -2365 13815 -2360
rect 13775 -2370 13815 -2365
rect 13885 -2365 13890 -2360
rect 13920 -2340 13925 -2335
rect 13995 -2335 14035 -2330
rect 13995 -2340 14000 -2335
rect 13920 -2360 14000 -2340
rect 13920 -2365 13925 -2360
rect 13885 -2370 13925 -2365
rect 13995 -2365 14000 -2360
rect 14030 -2365 14035 -2335
rect 13995 -2370 14035 -2365
rect 12950 -2395 12990 -2390
rect 12950 -2425 12955 -2395
rect 12985 -2400 12990 -2395
rect 13060 -2395 13100 -2390
rect 13060 -2400 13065 -2395
rect 12985 -2420 13065 -2400
rect 12985 -2425 12990 -2420
rect 12950 -2430 12990 -2425
rect 13060 -2425 13065 -2420
rect 13095 -2400 13100 -2395
rect 13170 -2395 13210 -2390
rect 13170 -2400 13175 -2395
rect 13095 -2420 13175 -2400
rect 13095 -2425 13100 -2420
rect 13060 -2430 13100 -2425
rect 13170 -2425 13175 -2420
rect 13205 -2400 13210 -2395
rect 13280 -2395 13320 -2390
rect 13280 -2400 13285 -2395
rect 13205 -2420 13285 -2400
rect 13205 -2425 13210 -2420
rect 13170 -2430 13210 -2425
rect 13280 -2425 13285 -2420
rect 13315 -2400 13320 -2395
rect 13390 -2395 13430 -2390
rect 13390 -2400 13395 -2395
rect 13315 -2420 13395 -2400
rect 13315 -2425 13320 -2420
rect 13280 -2430 13320 -2425
rect 13390 -2425 13395 -2420
rect 13425 -2400 13430 -2395
rect 13500 -2395 13540 -2390
rect 13500 -2400 13505 -2395
rect 13425 -2420 13505 -2400
rect 13425 -2425 13430 -2420
rect 13390 -2430 13430 -2425
rect 13500 -2425 13505 -2420
rect 13535 -2400 13540 -2395
rect 13610 -2395 13650 -2390
rect 13610 -2400 13615 -2395
rect 13535 -2420 13615 -2400
rect 13535 -2425 13540 -2420
rect 13500 -2430 13540 -2425
rect 13610 -2425 13615 -2420
rect 13645 -2400 13650 -2395
rect 13720 -2395 13760 -2390
rect 13720 -2400 13725 -2395
rect 13645 -2420 13725 -2400
rect 13645 -2425 13650 -2420
rect 13610 -2430 13650 -2425
rect 13720 -2425 13725 -2420
rect 13755 -2400 13760 -2395
rect 13830 -2395 13870 -2390
rect 13830 -2400 13835 -2395
rect 13755 -2420 13835 -2400
rect 13755 -2425 13760 -2420
rect 13720 -2430 13760 -2425
rect 13830 -2425 13835 -2420
rect 13865 -2400 13870 -2395
rect 13940 -2395 13980 -2390
rect 13940 -2400 13945 -2395
rect 13865 -2420 13945 -2400
rect 13865 -2425 13870 -2420
rect 13830 -2430 13870 -2425
rect 13940 -2425 13945 -2420
rect 13975 -2400 13980 -2395
rect 14050 -2395 14090 -2390
rect 14050 -2400 14055 -2395
rect 13975 -2420 14055 -2400
rect 13975 -2425 13980 -2420
rect 13940 -2430 13980 -2425
rect 14050 -2425 14055 -2420
rect 14085 -2425 14090 -2395
rect 14050 -2430 14090 -2425
rect 10980 -2525 11020 -2520
rect 10980 -2555 10985 -2525
rect 11015 -2530 11020 -2525
rect 11823 -2525 11857 -2520
rect 11823 -2530 11826 -2525
rect 11015 -2550 11826 -2530
rect 11015 -2555 11020 -2550
rect 10980 -2560 11020 -2555
rect 11823 -2555 11826 -2550
rect 11854 -2555 11857 -2525
rect 11823 -2560 11857 -2555
rect 13005 -2565 13045 -2560
rect 10970 -2580 11320 -2575
rect 10970 -2595 11285 -2580
rect 11280 -2610 11285 -2595
rect 11315 -2585 11320 -2580
rect 11520 -2580 11560 -2575
rect 11520 -2585 11525 -2580
rect 11315 -2605 11525 -2585
rect 11315 -2610 11320 -2605
rect 11280 -2615 11320 -2610
rect 11520 -2610 11525 -2605
rect 11555 -2585 11560 -2580
rect 11760 -2580 11800 -2575
rect 11760 -2585 11765 -2580
rect 11555 -2605 11765 -2585
rect 11555 -2610 11560 -2605
rect 11520 -2615 11560 -2610
rect 11760 -2610 11765 -2605
rect 11795 -2585 11800 -2580
rect 12000 -2580 12040 -2575
rect 12000 -2585 12005 -2580
rect 11795 -2605 12005 -2585
rect 11795 -2610 11800 -2605
rect 11760 -2615 11800 -2610
rect 12000 -2610 12005 -2605
rect 12035 -2585 12040 -2580
rect 12240 -2580 12280 -2575
rect 12240 -2585 12245 -2580
rect 12035 -2605 12245 -2585
rect 12035 -2610 12040 -2605
rect 12000 -2615 12040 -2610
rect 12240 -2610 12245 -2605
rect 12275 -2585 12280 -2580
rect 12480 -2580 12520 -2575
rect 12480 -2585 12485 -2580
rect 12275 -2605 12485 -2585
rect 12275 -2610 12280 -2605
rect 12240 -2615 12280 -2610
rect 12480 -2610 12485 -2605
rect 12515 -2610 12520 -2580
rect 13005 -2595 13010 -2565
rect 13040 -2570 13045 -2565
rect 13115 -2565 13155 -2560
rect 13115 -2570 13120 -2565
rect 13040 -2590 13120 -2570
rect 13040 -2595 13045 -2590
rect 13005 -2600 13045 -2595
rect 13115 -2595 13120 -2590
rect 13150 -2570 13155 -2565
rect 13225 -2565 13265 -2560
rect 13225 -2570 13230 -2565
rect 13150 -2590 13230 -2570
rect 13150 -2595 13155 -2590
rect 13115 -2600 13155 -2595
rect 13225 -2595 13230 -2590
rect 13260 -2570 13265 -2565
rect 13335 -2565 13375 -2560
rect 13335 -2570 13340 -2565
rect 13260 -2590 13340 -2570
rect 13260 -2595 13265 -2590
rect 13225 -2600 13265 -2595
rect 13335 -2595 13340 -2590
rect 13370 -2570 13375 -2565
rect 13445 -2565 13485 -2560
rect 13445 -2570 13450 -2565
rect 13370 -2590 13450 -2570
rect 13370 -2595 13375 -2590
rect 13335 -2600 13375 -2595
rect 13445 -2595 13450 -2590
rect 13480 -2570 13485 -2565
rect 13555 -2565 13595 -2560
rect 13555 -2570 13560 -2565
rect 13480 -2590 13560 -2570
rect 13480 -2595 13485 -2590
rect 13445 -2600 13485 -2595
rect 13555 -2595 13560 -2590
rect 13590 -2570 13595 -2565
rect 13665 -2565 13705 -2560
rect 13665 -2570 13670 -2565
rect 13590 -2590 13670 -2570
rect 13590 -2595 13595 -2590
rect 13555 -2600 13595 -2595
rect 13665 -2595 13670 -2590
rect 13700 -2570 13705 -2565
rect 13775 -2565 13815 -2560
rect 13775 -2570 13780 -2565
rect 13700 -2590 13780 -2570
rect 13700 -2595 13705 -2590
rect 13665 -2600 13705 -2595
rect 13775 -2595 13780 -2590
rect 13810 -2570 13815 -2565
rect 13885 -2565 13925 -2560
rect 13885 -2570 13890 -2565
rect 13810 -2590 13890 -2570
rect 13810 -2595 13815 -2590
rect 13775 -2600 13815 -2595
rect 13885 -2595 13890 -2590
rect 13920 -2570 13925 -2565
rect 13995 -2565 14035 -2560
rect 13995 -2570 14000 -2565
rect 13920 -2590 14000 -2570
rect 13920 -2595 13925 -2590
rect 13885 -2600 13925 -2595
rect 13995 -2595 14000 -2590
rect 14030 -2595 14035 -2565
rect 13995 -2600 14035 -2595
rect 12480 -2615 12520 -2610
rect 11400 -2625 11440 -2620
rect 11400 -2655 11405 -2625
rect 11435 -2630 11440 -2625
rect 11640 -2625 11680 -2620
rect 11640 -2630 11645 -2625
rect 11435 -2650 11645 -2630
rect 11435 -2655 11440 -2650
rect 11400 -2660 11440 -2655
rect 11640 -2655 11645 -2650
rect 11675 -2630 11680 -2625
rect 11880 -2625 11920 -2620
rect 11880 -2630 11885 -2625
rect 11675 -2650 11885 -2630
rect 11675 -2655 11680 -2650
rect 11640 -2660 11680 -2655
rect 11880 -2655 11885 -2650
rect 11915 -2630 11920 -2625
rect 12120 -2625 12160 -2620
rect 12120 -2630 12125 -2625
rect 11915 -2650 12125 -2630
rect 11915 -2655 11920 -2650
rect 11880 -2660 11920 -2655
rect 12120 -2655 12125 -2650
rect 12155 -2630 12160 -2625
rect 12360 -2625 12400 -2620
rect 12360 -2630 12365 -2625
rect 12155 -2650 12365 -2630
rect 12155 -2655 12160 -2650
rect 12120 -2660 12160 -2655
rect 12360 -2655 12365 -2650
rect 12395 -2630 12400 -2625
rect 12690 -2625 12730 -2620
rect 12690 -2630 12695 -2625
rect 12395 -2650 12695 -2630
rect 12395 -2655 12400 -2650
rect 12360 -2660 12400 -2655
rect 12690 -2655 12695 -2650
rect 12725 -2630 12730 -2625
rect 12975 -2625 13015 -2620
rect 12975 -2630 12980 -2625
rect 12725 -2650 12980 -2630
rect 12725 -2655 12730 -2650
rect 12690 -2660 12730 -2655
rect 12975 -2655 12980 -2650
rect 13010 -2655 13015 -2625
rect 12975 -2660 13015 -2655
rect 13005 -2685 13045 -2680
rect 13005 -2715 13010 -2685
rect 13040 -2690 13045 -2685
rect 13115 -2685 13155 -2680
rect 13115 -2690 13120 -2685
rect 13040 -2710 13120 -2690
rect 13040 -2715 13045 -2710
rect 11440 -2720 11480 -2715
rect 11440 -2750 11445 -2720
rect 11475 -2725 11480 -2720
rect 11660 -2720 11700 -2715
rect 11660 -2725 11665 -2720
rect 11475 -2745 11665 -2725
rect 11475 -2750 11480 -2745
rect 11440 -2755 11480 -2750
rect 11660 -2750 11665 -2745
rect 11695 -2725 11700 -2720
rect 11880 -2720 11920 -2715
rect 11880 -2725 11885 -2720
rect 11695 -2745 11885 -2725
rect 11695 -2750 11700 -2745
rect 11660 -2755 11700 -2750
rect 11880 -2750 11885 -2745
rect 11915 -2725 11920 -2720
rect 12100 -2720 12140 -2715
rect 12100 -2725 12105 -2720
rect 11915 -2745 12105 -2725
rect 11915 -2750 11920 -2745
rect 11880 -2755 11920 -2750
rect 12100 -2750 12105 -2745
rect 12135 -2725 12140 -2720
rect 12320 -2720 12360 -2715
rect 13005 -2720 13045 -2715
rect 13115 -2715 13120 -2710
rect 13150 -2690 13155 -2685
rect 13225 -2685 13265 -2680
rect 13225 -2690 13230 -2685
rect 13150 -2710 13230 -2690
rect 13150 -2715 13155 -2710
rect 13115 -2720 13155 -2715
rect 13225 -2715 13230 -2710
rect 13260 -2690 13265 -2685
rect 13335 -2685 13375 -2680
rect 13335 -2690 13340 -2685
rect 13260 -2710 13340 -2690
rect 13260 -2715 13265 -2710
rect 13225 -2720 13265 -2715
rect 13335 -2715 13340 -2710
rect 13370 -2690 13375 -2685
rect 13445 -2685 13485 -2680
rect 13445 -2690 13450 -2685
rect 13370 -2710 13450 -2690
rect 13370 -2715 13375 -2710
rect 13335 -2720 13375 -2715
rect 13445 -2715 13450 -2710
rect 13480 -2690 13485 -2685
rect 13555 -2685 13595 -2680
rect 13555 -2690 13560 -2685
rect 13480 -2710 13560 -2690
rect 13480 -2715 13485 -2710
rect 13445 -2720 13485 -2715
rect 13555 -2715 13560 -2710
rect 13590 -2690 13595 -2685
rect 13665 -2685 13705 -2680
rect 13665 -2690 13670 -2685
rect 13590 -2710 13670 -2690
rect 13590 -2715 13595 -2710
rect 13555 -2720 13595 -2715
rect 13665 -2715 13670 -2710
rect 13700 -2690 13705 -2685
rect 13775 -2685 13815 -2680
rect 13775 -2690 13780 -2685
rect 13700 -2710 13780 -2690
rect 13700 -2715 13705 -2710
rect 13665 -2720 13705 -2715
rect 13775 -2715 13780 -2710
rect 13810 -2690 13815 -2685
rect 13885 -2685 13925 -2680
rect 13885 -2690 13890 -2685
rect 13810 -2710 13890 -2690
rect 13810 -2715 13815 -2710
rect 13775 -2720 13815 -2715
rect 13885 -2715 13890 -2710
rect 13920 -2690 13925 -2685
rect 13995 -2685 14035 -2680
rect 13995 -2690 14000 -2685
rect 13920 -2710 14000 -2690
rect 13920 -2715 13925 -2710
rect 13885 -2720 13925 -2715
rect 13995 -2715 14000 -2710
rect 14030 -2715 14035 -2685
rect 13995 -2720 14035 -2715
rect 12320 -2725 12325 -2720
rect 12135 -2745 12325 -2725
rect 12135 -2750 12140 -2745
rect 12100 -2755 12140 -2750
rect 12320 -2750 12325 -2745
rect 12355 -2750 12360 -2720
rect 12320 -2755 12360 -2750
rect 11330 -2765 11370 -2760
rect 11330 -2795 11335 -2765
rect 11365 -2770 11370 -2765
rect 11550 -2765 11590 -2760
rect 11550 -2770 11555 -2765
rect 11365 -2790 11555 -2770
rect 11365 -2795 11370 -2790
rect 11330 -2800 11370 -2795
rect 11550 -2795 11555 -2790
rect 11585 -2770 11590 -2765
rect 11770 -2765 11810 -2760
rect 11770 -2770 11775 -2765
rect 11585 -2790 11775 -2770
rect 11585 -2795 11590 -2790
rect 11550 -2800 11590 -2795
rect 11770 -2795 11775 -2790
rect 11805 -2770 11810 -2765
rect 11990 -2765 12030 -2760
rect 11990 -2770 11995 -2765
rect 11805 -2790 11995 -2770
rect 11805 -2795 11810 -2790
rect 11770 -2800 11810 -2795
rect 11990 -2795 11995 -2790
rect 12025 -2770 12030 -2765
rect 12210 -2765 12250 -2760
rect 12210 -2770 12215 -2765
rect 12025 -2790 12215 -2770
rect 12025 -2795 12030 -2790
rect 11990 -2800 12030 -2795
rect 12210 -2795 12215 -2790
rect 12245 -2770 12250 -2765
rect 12430 -2765 12470 -2760
rect 12430 -2770 12435 -2765
rect 12245 -2790 12435 -2770
rect 12245 -2795 12250 -2790
rect 12210 -2800 12250 -2795
rect 12430 -2795 12435 -2790
rect 12465 -2795 12470 -2765
rect 12430 -2800 12470 -2795
rect 12950 -2905 12990 -2900
rect 12950 -2935 12955 -2905
rect 12985 -2910 12990 -2905
rect 13060 -2905 13100 -2900
rect 13060 -2910 13065 -2905
rect 12985 -2930 13065 -2910
rect 12985 -2935 12990 -2930
rect 12950 -2940 12990 -2935
rect 13060 -2935 13065 -2930
rect 13095 -2910 13100 -2905
rect 13170 -2905 13210 -2900
rect 13170 -2910 13175 -2905
rect 13095 -2930 13175 -2910
rect 13095 -2935 13100 -2930
rect 13060 -2940 13100 -2935
rect 13170 -2935 13175 -2930
rect 13205 -2910 13210 -2905
rect 13280 -2905 13320 -2900
rect 13280 -2910 13285 -2905
rect 13205 -2930 13285 -2910
rect 13205 -2935 13210 -2930
rect 13170 -2940 13210 -2935
rect 13280 -2935 13285 -2930
rect 13315 -2910 13320 -2905
rect 13390 -2905 13430 -2900
rect 13390 -2910 13395 -2905
rect 13315 -2930 13395 -2910
rect 13315 -2935 13320 -2930
rect 13280 -2940 13320 -2935
rect 13390 -2935 13395 -2930
rect 13425 -2910 13430 -2905
rect 13500 -2905 13540 -2900
rect 13500 -2910 13505 -2905
rect 13425 -2930 13505 -2910
rect 13425 -2935 13430 -2930
rect 13390 -2940 13430 -2935
rect 13500 -2935 13505 -2930
rect 13535 -2910 13540 -2905
rect 13610 -2905 13650 -2900
rect 13610 -2910 13615 -2905
rect 13535 -2930 13615 -2910
rect 13535 -2935 13540 -2930
rect 13500 -2940 13540 -2935
rect 13610 -2935 13615 -2930
rect 13645 -2910 13650 -2905
rect 13720 -2905 13760 -2900
rect 13720 -2910 13725 -2905
rect 13645 -2930 13725 -2910
rect 13645 -2935 13650 -2930
rect 13610 -2940 13650 -2935
rect 13720 -2935 13725 -2930
rect 13755 -2910 13760 -2905
rect 13830 -2905 13870 -2900
rect 13830 -2910 13835 -2905
rect 13755 -2930 13835 -2910
rect 13755 -2935 13760 -2930
rect 13720 -2940 13760 -2935
rect 13830 -2935 13835 -2930
rect 13865 -2910 13870 -2905
rect 13940 -2905 13980 -2900
rect 13940 -2910 13945 -2905
rect 13865 -2930 13945 -2910
rect 13865 -2935 13870 -2930
rect 13830 -2940 13870 -2935
rect 13940 -2935 13945 -2930
rect 13975 -2910 13980 -2905
rect 14050 -2905 14090 -2900
rect 14050 -2910 14055 -2905
rect 13975 -2930 14055 -2910
rect 13975 -2935 13980 -2930
rect 13940 -2940 13980 -2935
rect 14050 -2935 14055 -2930
rect 14085 -2935 14090 -2905
rect 14050 -2940 14090 -2935
rect 12995 -2965 13035 -2960
rect 12995 -2995 13000 -2965
rect 13030 -2970 13035 -2965
rect 13195 -2965 13235 -2960
rect 13195 -2970 13200 -2965
rect 13030 -2990 13200 -2970
rect 13030 -2995 13035 -2990
rect 12995 -3000 13035 -2995
rect 13195 -2995 13200 -2990
rect 13230 -2970 13235 -2965
rect 13395 -2965 13435 -2960
rect 13395 -2970 13400 -2965
rect 13230 -2990 13400 -2970
rect 13230 -2995 13235 -2990
rect 13195 -3000 13235 -2995
rect 13395 -2995 13400 -2990
rect 13430 -2970 13435 -2965
rect 13595 -2965 13635 -2960
rect 13595 -2970 13600 -2965
rect 13430 -2990 13600 -2970
rect 13430 -2995 13435 -2990
rect 13395 -3000 13435 -2995
rect 13595 -2995 13600 -2990
rect 13630 -2970 13635 -2965
rect 13795 -2965 13835 -2960
rect 13795 -2970 13800 -2965
rect 13630 -2990 13800 -2970
rect 13630 -2995 13635 -2990
rect 13595 -3000 13635 -2995
rect 13795 -2995 13800 -2990
rect 13830 -2970 13835 -2965
rect 13995 -2965 14035 -2960
rect 13995 -2970 14000 -2965
rect 13830 -2990 14000 -2970
rect 13830 -2995 13835 -2990
rect 13795 -3000 13835 -2995
rect 13995 -2995 14000 -2990
rect 14030 -2995 14035 -2965
rect 13995 -3000 14035 -2995
rect 11385 -3040 11425 -3035
rect 11385 -3070 11390 -3040
rect 11420 -3045 11425 -3040
rect 11605 -3040 11645 -3035
rect 11605 -3045 11610 -3040
rect 11420 -3065 11610 -3045
rect 11420 -3070 11425 -3065
rect 11385 -3075 11425 -3070
rect 11605 -3070 11610 -3065
rect 11640 -3045 11645 -3040
rect 11825 -3040 11865 -3035
rect 11825 -3045 11830 -3040
rect 11640 -3065 11830 -3045
rect 11640 -3070 11645 -3065
rect 11605 -3075 11645 -3070
rect 11825 -3070 11830 -3065
rect 11860 -3045 11865 -3040
rect 12045 -3040 12085 -3035
rect 12045 -3045 12050 -3040
rect 11860 -3065 12050 -3045
rect 11860 -3070 11865 -3065
rect 11825 -3075 11865 -3070
rect 12045 -3070 12050 -3065
rect 12080 -3045 12085 -3040
rect 12265 -3040 12305 -3035
rect 12265 -3045 12270 -3040
rect 12080 -3065 12270 -3045
rect 12080 -3070 12085 -3065
rect 12045 -3075 12085 -3070
rect 12265 -3070 12270 -3065
rect 12300 -3070 12305 -3040
rect 12265 -3075 12305 -3070
rect 11495 -3095 11535 -3090
rect 11495 -3125 11500 -3095
rect 11530 -3100 11535 -3095
rect 11715 -3095 11755 -3090
rect 11715 -3100 11720 -3095
rect 11530 -3120 11720 -3100
rect 11530 -3125 11535 -3120
rect 11495 -3130 11535 -3125
rect 11715 -3125 11720 -3120
rect 11750 -3100 11755 -3095
rect 11935 -3095 11975 -3090
rect 11935 -3100 11940 -3095
rect 11750 -3120 11940 -3100
rect 11750 -3125 11755 -3120
rect 11715 -3130 11755 -3125
rect 11935 -3125 11940 -3120
rect 11970 -3100 11975 -3095
rect 12155 -3095 12195 -3090
rect 12155 -3100 12160 -3095
rect 11970 -3120 12160 -3100
rect 11970 -3125 11975 -3120
rect 11935 -3130 11975 -3125
rect 12155 -3125 12160 -3120
rect 12190 -3100 12195 -3095
rect 12375 -3095 12415 -3090
rect 12375 -3100 12380 -3095
rect 12190 -3120 12380 -3100
rect 12190 -3125 12195 -3120
rect 12155 -3130 12195 -3125
rect 12375 -3125 12380 -3120
rect 12410 -3125 12415 -3095
rect 12375 -3130 12415 -3125
rect 11190 -3150 11230 -3145
rect 11190 -3180 11195 -3150
rect 11225 -3155 11230 -3150
rect 11410 -3150 11450 -3145
rect 11410 -3155 11415 -3150
rect 11225 -3175 11415 -3155
rect 11225 -3180 11230 -3175
rect 11190 -3185 11230 -3180
rect 11410 -3180 11415 -3175
rect 11445 -3155 11450 -3150
rect 11640 -3150 11680 -3145
rect 11640 -3155 11645 -3150
rect 11445 -3175 11645 -3155
rect 11445 -3180 11450 -3175
rect 11410 -3185 11450 -3180
rect 11640 -3180 11645 -3175
rect 11675 -3155 11680 -3150
rect 12230 -3150 12270 -3145
rect 12230 -3155 12235 -3150
rect 11675 -3175 12235 -3155
rect 11675 -3180 11680 -3175
rect 11640 -3185 11680 -3180
rect 12230 -3180 12235 -3175
rect 12265 -3155 12270 -3150
rect 12450 -3150 12490 -3145
rect 12450 -3155 12455 -3150
rect 12265 -3175 12455 -3155
rect 12265 -3180 12270 -3175
rect 12230 -3185 12270 -3180
rect 12450 -3180 12455 -3175
rect 12485 -3155 12490 -3150
rect 12680 -3150 12720 -3145
rect 12680 -3155 12685 -3150
rect 12485 -3175 12685 -3155
rect 12485 -3180 12490 -3175
rect 12450 -3185 12490 -3180
rect 12680 -3180 12685 -3175
rect 12715 -3180 12720 -3150
rect 12680 -3185 12720 -3180
rect 11820 -3195 11860 -3190
rect 11820 -3225 11825 -3195
rect 11855 -3200 11860 -3195
rect 11940 -3195 11980 -3190
rect 11940 -3200 11945 -3195
rect 11855 -3220 11945 -3200
rect 11855 -3225 11860 -3220
rect 11820 -3230 11860 -3225
rect 11940 -3225 11945 -3220
rect 11975 -3225 11980 -3195
rect 11940 -3230 11980 -3225
rect 11085 -3240 11125 -3235
rect 11085 -3270 11090 -3240
rect 11120 -3245 11125 -3240
rect 11305 -3240 11345 -3235
rect 11305 -3245 11310 -3240
rect 11120 -3265 11310 -3245
rect 11120 -3270 11125 -3265
rect 11085 -3275 11125 -3270
rect 11305 -3270 11310 -3265
rect 11340 -3245 11345 -3240
rect 11525 -3240 11565 -3235
rect 11525 -3245 11530 -3240
rect 11340 -3265 11530 -3245
rect 11340 -3270 11345 -3265
rect 11305 -3275 11345 -3270
rect 11525 -3270 11530 -3265
rect 11560 -3245 11565 -3240
rect 12125 -3240 12165 -3235
rect 12125 -3245 12130 -3240
rect 11560 -3265 12130 -3245
rect 11560 -3270 11565 -3265
rect 11525 -3275 11565 -3270
rect 12125 -3270 12130 -3265
rect 12160 -3245 12165 -3240
rect 12345 -3240 12385 -3235
rect 12345 -3245 12350 -3240
rect 12160 -3265 12350 -3245
rect 12160 -3270 12165 -3265
rect 12125 -3275 12165 -3270
rect 12345 -3270 12350 -3265
rect 12380 -3245 12385 -3240
rect 12565 -3240 12605 -3235
rect 12565 -3245 12570 -3240
rect 12380 -3265 12570 -3245
rect 12380 -3270 12385 -3265
rect 12345 -3275 12385 -3270
rect 12565 -3270 12570 -3265
rect 12600 -3270 12605 -3240
rect 12565 -3275 12605 -3270
rect 11237 -3285 11269 -3280
rect 11237 -3290 11240 -3285
rect 10970 -3310 11240 -3290
rect 11237 -3315 11240 -3310
rect 11266 -3290 11269 -3285
rect 11457 -3285 11489 -3280
rect 11457 -3290 11460 -3285
rect 11266 -3310 11460 -3290
rect 11266 -3315 11269 -3310
rect 11237 -3320 11269 -3315
rect 11457 -3315 11460 -3310
rect 11486 -3290 11489 -3285
rect 11601 -3285 11633 -3280
rect 11601 -3290 11604 -3285
rect 11486 -3310 11604 -3290
rect 11486 -3315 11489 -3310
rect 11457 -3320 11489 -3315
rect 11601 -3315 11604 -3310
rect 11630 -3290 11633 -3285
rect 11867 -3285 11899 -3280
rect 11867 -3290 11870 -3285
rect 11630 -3310 11870 -3290
rect 11630 -3315 11633 -3310
rect 11601 -3320 11633 -3315
rect 11867 -3315 11870 -3310
rect 11896 -3290 11899 -3285
rect 12277 -3285 12309 -3280
rect 12277 -3290 12280 -3285
rect 11896 -3310 12280 -3290
rect 11896 -3315 11899 -3310
rect 11867 -3320 11899 -3315
rect 12277 -3315 12280 -3310
rect 12306 -3290 12309 -3285
rect 12497 -3285 12529 -3280
rect 12497 -3290 12500 -3285
rect 12306 -3310 12500 -3290
rect 12306 -3315 12309 -3310
rect 12277 -3320 12309 -3315
rect 12497 -3315 12500 -3310
rect 12526 -3290 12529 -3285
rect 12641 -3285 12673 -3280
rect 12641 -3290 12644 -3285
rect 12526 -3310 12644 -3290
rect 12526 -3315 12529 -3310
rect 12497 -3320 12529 -3315
rect 12641 -3315 12644 -3310
rect 12670 -3315 12673 -3285
rect 12641 -3320 12673 -3315
rect 13095 -3315 13135 -3310
rect 13095 -3345 13100 -3315
rect 13130 -3320 13135 -3315
rect 13295 -3315 13335 -3310
rect 13295 -3320 13300 -3315
rect 13130 -3340 13300 -3320
rect 13130 -3345 13135 -3340
rect 13095 -3350 13135 -3345
rect 13295 -3345 13300 -3340
rect 13330 -3320 13335 -3315
rect 13495 -3315 13535 -3310
rect 13495 -3320 13500 -3315
rect 13330 -3340 13500 -3320
rect 13330 -3345 13335 -3340
rect 13295 -3350 13335 -3345
rect 13495 -3345 13500 -3340
rect 13530 -3320 13535 -3315
rect 13695 -3315 13735 -3310
rect 13695 -3320 13700 -3315
rect 13530 -3340 13700 -3320
rect 13530 -3345 13535 -3340
rect 13495 -3350 13535 -3345
rect 13695 -3345 13700 -3340
rect 13730 -3320 13735 -3315
rect 13895 -3315 13935 -3310
rect 13895 -3320 13900 -3315
rect 13730 -3340 13900 -3320
rect 13730 -3345 13735 -3340
rect 13695 -3350 13735 -3345
rect 13895 -3345 13900 -3340
rect 13930 -3345 13935 -3315
rect 13895 -3350 13935 -3345
rect 11106 -3505 11138 -3500
rect 11106 -3510 11109 -3505
rect 10970 -3530 11109 -3510
rect 11106 -3535 11109 -3530
rect 11135 -3510 11138 -3505
rect 11305 -3505 11345 -3500
rect 11305 -3510 11310 -3505
rect 11135 -3530 11310 -3510
rect 11135 -3535 11138 -3530
rect 11106 -3540 11138 -3535
rect 11305 -3535 11310 -3530
rect 11340 -3510 11345 -3505
rect 11525 -3505 11565 -3500
rect 11525 -3510 11530 -3505
rect 11340 -3530 11530 -3510
rect 11340 -3535 11345 -3530
rect 11305 -3540 11345 -3535
rect 11525 -3535 11530 -3530
rect 11560 -3510 11565 -3505
rect 11922 -3505 11954 -3500
rect 11922 -3510 11925 -3505
rect 11560 -3530 11925 -3510
rect 11560 -3535 11565 -3530
rect 11525 -3540 11565 -3535
rect 11922 -3535 11925 -3530
rect 11951 -3510 11954 -3505
rect 12146 -3505 12178 -3500
rect 12146 -3510 12149 -3505
rect 11951 -3530 12149 -3510
rect 11951 -3535 11954 -3530
rect 11922 -3540 11954 -3535
rect 12146 -3535 12149 -3530
rect 12175 -3510 12178 -3505
rect 12345 -3505 12385 -3500
rect 12345 -3510 12350 -3505
rect 12175 -3530 12350 -3510
rect 12175 -3535 12178 -3530
rect 12146 -3540 12178 -3535
rect 12345 -3535 12350 -3530
rect 12380 -3510 12385 -3505
rect 12565 -3505 12605 -3500
rect 12565 -3510 12570 -3505
rect 12380 -3530 12570 -3510
rect 12380 -3535 12385 -3530
rect 12345 -3540 12385 -3535
rect 12565 -3535 12570 -3530
rect 12600 -3535 12605 -3505
rect 12565 -3540 12605 -3535
rect 11145 -3565 11185 -3560
rect 11145 -3595 11150 -3565
rect 11180 -3570 11185 -3565
rect 11250 -3565 11290 -3560
rect 11250 -3570 11255 -3565
rect 11180 -3590 11255 -3570
rect 11180 -3595 11185 -3590
rect 11145 -3600 11185 -3595
rect 11250 -3595 11255 -3590
rect 11285 -3570 11290 -3565
rect 11360 -3565 11400 -3560
rect 11360 -3570 11365 -3565
rect 11285 -3590 11365 -3570
rect 11285 -3595 11290 -3590
rect 11250 -3600 11290 -3595
rect 11360 -3595 11365 -3590
rect 11395 -3570 11400 -3565
rect 11470 -3565 11510 -3560
rect 11470 -3570 11475 -3565
rect 11395 -3590 11475 -3570
rect 11395 -3595 11400 -3590
rect 11360 -3600 11400 -3595
rect 11470 -3595 11475 -3590
rect 11505 -3570 11510 -3565
rect 11580 -3565 11620 -3560
rect 11580 -3570 11585 -3565
rect 11505 -3590 11585 -3570
rect 11505 -3595 11510 -3590
rect 11470 -3600 11510 -3595
rect 11580 -3595 11585 -3590
rect 11615 -3570 11620 -3565
rect 12185 -3565 12225 -3560
rect 12185 -3570 12190 -3565
rect 11615 -3590 12190 -3570
rect 11615 -3595 11620 -3590
rect 11580 -3600 11620 -3595
rect 12185 -3595 12190 -3590
rect 12220 -3570 12225 -3565
rect 12290 -3565 12330 -3560
rect 12290 -3570 12295 -3565
rect 12220 -3590 12295 -3570
rect 12220 -3595 12225 -3590
rect 12185 -3600 12225 -3595
rect 12290 -3595 12295 -3590
rect 12325 -3570 12330 -3565
rect 12400 -3565 12440 -3560
rect 12400 -3570 12405 -3565
rect 12325 -3590 12405 -3570
rect 12325 -3595 12330 -3590
rect 12290 -3600 12330 -3595
rect 12400 -3595 12405 -3590
rect 12435 -3570 12440 -3565
rect 12510 -3565 12550 -3560
rect 12510 -3570 12515 -3565
rect 12435 -3590 12515 -3570
rect 12435 -3595 12440 -3590
rect 12400 -3600 12440 -3595
rect 12510 -3595 12515 -3590
rect 12545 -3570 12550 -3565
rect 12620 -3565 12660 -3560
rect 12620 -3570 12625 -3565
rect 12545 -3590 12625 -3570
rect 12545 -3595 12550 -3590
rect 12510 -3600 12550 -3595
rect 12620 -3595 12625 -3590
rect 12655 -3595 12660 -3565
rect 12620 -3600 12660 -3595
rect 10970 -3635 12805 -3615
rect 11810 -3655 11850 -3650
rect 11810 -3685 11815 -3655
rect 11845 -3685 11850 -3655
rect 11810 -3690 11850 -3685
rect 11315 -3705 11355 -3700
rect 11315 -3735 11320 -3705
rect 11350 -3710 11355 -3705
rect 11880 -3705 11920 -3700
rect 11880 -3710 11885 -3705
rect 11350 -3730 11885 -3710
rect 11350 -3735 11355 -3730
rect 11315 -3740 11355 -3735
rect 11880 -3735 11885 -3730
rect 11915 -3735 11920 -3705
rect 11880 -3740 11920 -3735
rect 12595 -3750 12635 -3745
rect 11425 -3765 11465 -3760
rect 11425 -3795 11430 -3765
rect 11460 -3770 11465 -3765
rect 11535 -3765 11575 -3760
rect 11535 -3770 11540 -3765
rect 11460 -3790 11540 -3770
rect 11460 -3795 11465 -3790
rect 11425 -3800 11465 -3795
rect 11535 -3795 11540 -3790
rect 11570 -3770 11575 -3765
rect 11645 -3765 11685 -3760
rect 11645 -3770 11650 -3765
rect 11570 -3790 11650 -3770
rect 11570 -3795 11575 -3790
rect 11535 -3800 11575 -3795
rect 11645 -3795 11650 -3790
rect 11680 -3770 11685 -3765
rect 11755 -3765 11795 -3760
rect 11755 -3770 11760 -3765
rect 11680 -3790 11760 -3770
rect 11680 -3795 11685 -3790
rect 11645 -3800 11685 -3795
rect 11755 -3795 11760 -3790
rect 11790 -3770 11795 -3765
rect 11865 -3765 11905 -3760
rect 11865 -3770 11870 -3765
rect 11790 -3790 11870 -3770
rect 11790 -3795 11795 -3790
rect 11755 -3800 11795 -3795
rect 11865 -3795 11870 -3790
rect 11900 -3770 11905 -3765
rect 11975 -3765 12015 -3760
rect 11975 -3770 11980 -3765
rect 11900 -3790 11980 -3770
rect 11900 -3795 11905 -3790
rect 11865 -3800 11905 -3795
rect 11975 -3795 11980 -3790
rect 12010 -3770 12015 -3765
rect 12085 -3765 12125 -3760
rect 12085 -3770 12090 -3765
rect 12010 -3790 12090 -3770
rect 12010 -3795 12015 -3790
rect 11975 -3800 12015 -3795
rect 12085 -3795 12090 -3790
rect 12120 -3770 12125 -3765
rect 12195 -3765 12235 -3760
rect 12195 -3770 12200 -3765
rect 12120 -3790 12200 -3770
rect 12120 -3795 12125 -3790
rect 12085 -3800 12125 -3795
rect 12195 -3795 12200 -3790
rect 12230 -3770 12235 -3765
rect 12305 -3765 12345 -3760
rect 12305 -3770 12310 -3765
rect 12230 -3790 12310 -3770
rect 12230 -3795 12235 -3790
rect 12195 -3800 12235 -3795
rect 12305 -3795 12310 -3790
rect 12340 -3770 12345 -3765
rect 12415 -3765 12455 -3760
rect 12415 -3770 12420 -3765
rect 12340 -3790 12420 -3770
rect 12340 -3795 12345 -3790
rect 12305 -3800 12345 -3795
rect 12415 -3795 12420 -3790
rect 12450 -3770 12455 -3765
rect 12525 -3765 12565 -3760
rect 12525 -3770 12530 -3765
rect 12450 -3790 12530 -3770
rect 12450 -3795 12455 -3790
rect 12415 -3800 12455 -3795
rect 12525 -3795 12530 -3790
rect 12560 -3795 12565 -3765
rect 12595 -3780 12600 -3750
rect 12630 -3755 12635 -3750
rect 12630 -3775 12695 -3755
rect 12630 -3780 12635 -3775
rect 12595 -3785 12635 -3780
rect 12525 -3800 12565 -3795
rect 11165 -4085 11205 -4080
rect 11165 -4115 11170 -4085
rect 11200 -4090 11205 -4085
rect 11260 -4085 11300 -4080
rect 11260 -4090 11265 -4085
rect 11200 -4110 11265 -4090
rect 11200 -4115 11205 -4110
rect 11165 -4120 11205 -4115
rect 11260 -4115 11265 -4110
rect 11295 -4090 11300 -4085
rect 11370 -4085 11410 -4080
rect 11370 -4090 11375 -4085
rect 11295 -4110 11375 -4090
rect 11295 -4115 11300 -4110
rect 11260 -4120 11300 -4115
rect 11370 -4115 11375 -4110
rect 11405 -4090 11410 -4085
rect 11480 -4085 11520 -4080
rect 11480 -4090 11485 -4085
rect 11405 -4110 11485 -4090
rect 11405 -4115 11410 -4110
rect 11370 -4120 11410 -4115
rect 11480 -4115 11485 -4110
rect 11515 -4090 11520 -4085
rect 11590 -4085 11630 -4080
rect 11590 -4090 11595 -4085
rect 11515 -4110 11595 -4090
rect 11515 -4115 11520 -4110
rect 11480 -4120 11520 -4115
rect 11590 -4115 11595 -4110
rect 11625 -4090 11630 -4085
rect 11700 -4085 11740 -4080
rect 11700 -4090 11705 -4085
rect 11625 -4110 11705 -4090
rect 11625 -4115 11630 -4110
rect 11590 -4120 11630 -4115
rect 11700 -4115 11705 -4110
rect 11735 -4090 11740 -4085
rect 11810 -4085 11850 -4080
rect 11810 -4090 11815 -4085
rect 11735 -4110 11815 -4090
rect 11735 -4115 11740 -4110
rect 11700 -4120 11740 -4115
rect 11810 -4115 11815 -4110
rect 11845 -4090 11850 -4085
rect 11920 -4085 11960 -4080
rect 11920 -4090 11925 -4085
rect 11845 -4110 11925 -4090
rect 11845 -4115 11850 -4110
rect 11810 -4120 11850 -4115
rect 11920 -4115 11925 -4110
rect 11955 -4090 11960 -4085
rect 12030 -4085 12070 -4080
rect 12030 -4090 12035 -4085
rect 11955 -4110 12035 -4090
rect 11955 -4115 11960 -4110
rect 11920 -4120 11960 -4115
rect 12030 -4115 12035 -4110
rect 12065 -4090 12070 -4085
rect 12140 -4085 12180 -4080
rect 12140 -4090 12145 -4085
rect 12065 -4110 12145 -4090
rect 12065 -4115 12070 -4110
rect 12030 -4120 12070 -4115
rect 12140 -4115 12145 -4110
rect 12175 -4090 12180 -4085
rect 12250 -4085 12290 -4080
rect 12250 -4090 12255 -4085
rect 12175 -4110 12255 -4090
rect 12175 -4115 12180 -4110
rect 12140 -4120 12180 -4115
rect 12250 -4115 12255 -4110
rect 12285 -4090 12290 -4085
rect 12360 -4085 12400 -4080
rect 12360 -4090 12365 -4085
rect 12285 -4110 12365 -4090
rect 12285 -4115 12290 -4110
rect 12250 -4120 12290 -4115
rect 12360 -4115 12365 -4110
rect 12395 -4090 12400 -4085
rect 12470 -4085 12510 -4080
rect 12470 -4090 12475 -4085
rect 12395 -4110 12475 -4090
rect 12395 -4115 12400 -4110
rect 12360 -4120 12400 -4115
rect 12470 -4115 12475 -4110
rect 12505 -4090 12510 -4085
rect 12620 -4085 12660 -4080
rect 12620 -4090 12625 -4085
rect 12505 -4110 12625 -4090
rect 12505 -4115 12510 -4110
rect 12470 -4120 12510 -4115
rect 12620 -4115 12625 -4110
rect 12655 -4115 12660 -4085
rect 12620 -4120 12660 -4115
<< via2 >>
rect -190 4960 -160 4990
rect 5555 4960 5585 4990
rect -105 3495 -75 3525
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 5555 3415 5585 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 3110 -75 3140
rect -105 2970 -75 3000
rect -105 2880 -75 2910
rect 5555 2780 5585 2810
rect 5555 2065 5585 2095
rect -105 1690 -75 1720
rect 5555 1470 5585 1500
rect 5470 1155 5500 1185
rect 5470 1010 5500 1040
rect 5470 900 5500 930
rect -190 545 -160 575
<< metal3 >>
rect -200 4995 -150 5000
rect -200 4955 -195 4995
rect -155 4955 -150 4995
rect -200 4950 -150 4955
rect 5545 4995 5595 5000
rect 5545 4955 5550 4995
rect 5590 4955 5595 4995
rect 5545 4950 5595 4955
rect -195 585 -155 4950
rect -115 4910 -65 4915
rect -115 4870 -110 4910
rect -70 4870 -65 4910
rect -115 4865 -65 4870
rect 5460 4910 5510 4915
rect 5460 4870 5465 4910
rect 5505 4870 5510 4910
rect 5460 4865 5510 4870
rect -110 3525 -70 4865
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3140 -70 3495
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 3110 -105 3140
rect -75 3110 -70 3140
rect -110 3000 -70 3110
rect -110 2970 -105 3000
rect -75 2970 -70 3000
rect -110 2910 -70 2970
rect -110 2880 -105 2910
rect -75 2880 -70 2910
rect -110 1720 -70 2880
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5465 1185 5505 4865
rect 5465 1155 5470 1185
rect 5500 1155 5505 1185
rect 5465 1040 5505 1155
rect 5465 1010 5470 1040
rect 5500 1010 5505 1040
rect 5465 930 5505 1010
rect 5465 900 5470 930
rect 5500 900 5505 930
rect 5465 665 5505 900
rect 5550 3445 5590 4950
rect 12965 4375 13195 4605
rect 13315 4375 13545 4605
rect 13665 4375 13895 4605
rect 14015 4375 14245 4605
rect 14365 4375 14595 4605
rect 14715 4375 14945 4605
rect 15065 4375 15295 4605
rect 15415 4375 15645 4605
rect 12965 4025 13195 4255
rect 13315 4025 13545 4255
rect 13665 4025 13895 4255
rect 14015 4025 14245 4255
rect 14365 4025 14595 4255
rect 14715 4025 14945 4255
rect 15065 4025 15295 4255
rect 15415 4025 15645 4255
rect 12965 3675 13195 3905
rect 13315 3675 13545 3905
rect 13665 3675 13895 3905
rect 14015 3675 14245 3905
rect 14365 3675 14595 3905
rect 14715 3675 14945 3905
rect 15065 3675 15295 3905
rect 15415 3675 15645 3905
rect 5550 3415 5555 3445
rect 5585 3415 5590 3445
rect 5550 2810 5590 3415
rect 14365 3325 14595 3555
rect 14715 3325 14945 3555
rect 15065 3325 15295 3555
rect 15415 3325 15645 3555
rect 14365 2975 14595 3205
rect 14715 2975 14945 3205
rect 15065 2975 15295 3205
rect 15415 2975 15645 3205
rect 5550 2780 5555 2810
rect 5585 2780 5590 2810
rect 5550 2095 5590 2780
rect 14365 2625 14595 2855
rect 14715 2625 14945 2855
rect 15065 2625 15295 2855
rect 15415 2625 15645 2855
rect 14365 2275 14595 2505
rect 14715 2275 14945 2505
rect 15065 2275 15295 2505
rect 15415 2275 15645 2505
rect 5550 2065 5555 2095
rect 5585 2065 5590 2095
rect 5550 1500 5590 2065
rect 14365 1925 14595 2155
rect 14715 1925 14945 2155
rect 15065 1925 15295 2155
rect 15415 1925 15645 2155
rect 14365 1575 14595 1805
rect 14715 1575 14945 1805
rect 15065 1575 15295 1805
rect 15415 1575 15645 1805
rect 5550 1470 5555 1500
rect 5585 1470 5590 1500
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5460 660 5510 665
rect 5460 620 5465 660
rect 5505 620 5510 660
rect 5460 615 5510 620
rect 5550 585 5590 1470
rect 14365 1225 14595 1455
rect 14715 1225 14945 1455
rect 15065 1225 15295 1455
rect 15415 1225 15645 1455
rect 14365 875 14595 1105
rect 14715 875 14945 1105
rect 15065 875 15295 1105
rect 15415 875 15645 1105
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5545 580 5595 585
rect 5545 540 5550 580
rect 5590 540 5595 580
rect 5545 535 5595 540
rect 14365 525 14595 755
rect 14715 525 14945 755
rect 15065 525 15295 755
rect 15415 525 15645 755
rect 11915 175 12145 405
rect 12265 175 12495 405
rect 12615 175 12845 405
rect 12965 175 13195 405
rect 13315 175 13545 405
rect 13665 175 13895 405
rect 14015 175 14245 405
rect 14365 175 14595 405
rect 14715 175 14945 405
rect 15065 175 15295 405
rect 15415 175 15645 405
rect 11915 -175 12145 55
rect 12265 -175 12495 55
rect 12615 -175 12845 55
rect 12965 -175 13195 55
rect 13315 -175 13545 55
rect 13665 -175 13895 55
rect 14015 -175 14245 55
rect 14365 -175 14595 55
rect 14715 -175 14945 55
rect 15065 -175 15295 55
rect 15415 -175 15645 55
rect 11915 -525 12145 -295
rect 12265 -525 12495 -295
rect 12615 -525 12845 -295
rect 12965 -525 13195 -295
rect 13315 -525 13545 -295
rect 13665 -525 13895 -295
rect 14015 -525 14245 -295
rect 14365 -525 14595 -295
rect 14715 -525 14945 -295
rect 15065 -525 15295 -295
rect 15415 -525 15645 -295
<< via3 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -190 4960 -160 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5555 4960 5585 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect -110 4870 -70 4910
rect 5465 4870 5505 4910
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect -110 620 -70 660
rect 5465 620 5505 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5550 540 5590 580
<< mimcap >>
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 12980 4515 13180 4590
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 12980 4475 13060 4515
rect 13100 4475 13180 4515
rect 12980 4390 13180 4475
rect 13330 4515 13530 4590
rect 13330 4475 13410 4515
rect 13450 4475 13530 4515
rect 13330 4390 13530 4475
rect 13680 4515 13880 4590
rect 13680 4475 13760 4515
rect 13800 4475 13880 4515
rect 13680 4390 13880 4475
rect 14030 4515 14230 4590
rect 14030 4475 14110 4515
rect 14150 4475 14230 4515
rect 14030 4390 14230 4475
rect 14380 4515 14580 4590
rect 14380 4475 14460 4515
rect 14500 4475 14580 4515
rect 14380 4390 14580 4475
rect 14730 4515 14930 4590
rect 14730 4475 14810 4515
rect 14850 4475 14930 4515
rect 14730 4390 14930 4475
rect 15080 4515 15280 4590
rect 15080 4475 15160 4515
rect 15200 4475 15280 4515
rect 15080 4390 15280 4475
rect 15430 4515 15630 4590
rect 15430 4475 15510 4515
rect 15550 4475 15630 4515
rect 15430 4390 15630 4475
rect 5060 4290 5260 4375
rect 12980 4165 13180 4240
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 12980 4125 13060 4165
rect 13100 4125 13180 4165
rect 12980 4040 13180 4125
rect 13330 4165 13530 4240
rect 13330 4125 13410 4165
rect 13450 4125 13530 4165
rect 13330 4040 13530 4125
rect 13680 4165 13880 4240
rect 13680 4125 13760 4165
rect 13800 4125 13880 4165
rect 13680 4040 13880 4125
rect 14030 4165 14230 4240
rect 14030 4125 14110 4165
rect 14150 4125 14230 4165
rect 14030 4040 14230 4125
rect 14380 4165 14580 4240
rect 14380 4125 14460 4165
rect 14500 4125 14580 4165
rect 14380 4040 14580 4125
rect 14730 4165 14930 4240
rect 14730 4125 14810 4165
rect 14850 4125 14930 4165
rect 14730 4040 14930 4125
rect 15080 4165 15280 4240
rect 15080 4125 15160 4165
rect 15200 4125 15280 4165
rect 15080 4040 15280 4125
rect 15430 4165 15630 4240
rect 15430 4125 15510 4165
rect 15550 4125 15630 4165
rect 15430 4040 15630 4125
rect 5060 3940 5260 4025
rect 12980 3815 13180 3890
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 12980 3775 13060 3815
rect 13100 3775 13180 3815
rect 12980 3690 13180 3775
rect 13330 3815 13530 3890
rect 13330 3775 13410 3815
rect 13450 3775 13530 3815
rect 13330 3690 13530 3775
rect 13680 3815 13880 3890
rect 13680 3775 13760 3815
rect 13800 3775 13880 3815
rect 13680 3690 13880 3775
rect 14030 3815 14230 3890
rect 14030 3775 14110 3815
rect 14150 3775 14230 3815
rect 14030 3690 14230 3775
rect 14380 3815 14580 3890
rect 14380 3775 14460 3815
rect 14500 3775 14580 3815
rect 14380 3690 14580 3775
rect 14730 3815 14930 3890
rect 14730 3775 14810 3815
rect 14850 3775 14930 3815
rect 14730 3690 14930 3775
rect 15080 3815 15280 3890
rect 15080 3775 15160 3815
rect 15200 3775 15280 3815
rect 15080 3690 15280 3775
rect 15430 3815 15630 3890
rect 15430 3775 15510 3815
rect 15550 3775 15630 3815
rect 15430 3690 15630 3775
rect 5060 3590 5260 3675
rect 14380 3465 14580 3540
rect 14380 3425 14460 3465
rect 14500 3425 14580 3465
rect 14380 3340 14580 3425
rect 14730 3465 14930 3540
rect 14730 3425 14810 3465
rect 14850 3425 14930 3465
rect 14730 3340 14930 3425
rect 15080 3465 15280 3540
rect 15080 3425 15160 3465
rect 15200 3425 15280 3465
rect 15080 3340 15280 3425
rect 15430 3465 15630 3540
rect 15430 3425 15510 3465
rect 15550 3425 15630 3465
rect 15430 3340 15630 3425
rect 14380 3115 14580 3190
rect 14380 3075 14460 3115
rect 14500 3075 14580 3115
rect 14380 2990 14580 3075
rect 14730 3115 14930 3190
rect 14730 3075 14810 3115
rect 14850 3075 14930 3115
rect 14730 2990 14930 3075
rect 15080 3115 15280 3190
rect 15080 3075 15160 3115
rect 15200 3075 15280 3115
rect 15080 2990 15280 3075
rect 15430 3115 15630 3190
rect 15430 3075 15510 3115
rect 15550 3075 15630 3115
rect 15430 2990 15630 3075
rect 14380 2765 14580 2840
rect 14380 2725 14460 2765
rect 14500 2725 14580 2765
rect 14380 2640 14580 2725
rect 14730 2765 14930 2840
rect 14730 2725 14810 2765
rect 14850 2725 14930 2765
rect 14730 2640 14930 2725
rect 15080 2765 15280 2840
rect 15080 2725 15160 2765
rect 15200 2725 15280 2765
rect 15080 2640 15280 2725
rect 15430 2765 15630 2840
rect 15430 2725 15510 2765
rect 15550 2725 15630 2765
rect 15430 2640 15630 2725
rect 14380 2415 14580 2490
rect 14380 2375 14460 2415
rect 14500 2375 14580 2415
rect 14380 2290 14580 2375
rect 14730 2415 14930 2490
rect 14730 2375 14810 2415
rect 14850 2375 14930 2415
rect 14730 2290 14930 2375
rect 15080 2415 15280 2490
rect 15080 2375 15160 2415
rect 15200 2375 15280 2415
rect 15080 2290 15280 2375
rect 15430 2415 15630 2490
rect 15430 2375 15510 2415
rect 15550 2375 15630 2415
rect 15430 2290 15630 2375
rect 14380 2065 14580 2140
rect 14380 2025 14460 2065
rect 14500 2025 14580 2065
rect 14380 1940 14580 2025
rect 14730 2065 14930 2140
rect 14730 2025 14810 2065
rect 14850 2025 14930 2065
rect 14730 1940 14930 2025
rect 15080 2065 15280 2140
rect 15080 2025 15160 2065
rect 15200 2025 15280 2065
rect 15080 1940 15280 2025
rect 15430 2065 15630 2140
rect 15430 2025 15510 2065
rect 15550 2025 15630 2065
rect 15430 1940 15630 2025
rect 14380 1715 14580 1790
rect 14380 1675 14460 1715
rect 14500 1675 14580 1715
rect 14380 1590 14580 1675
rect 14730 1715 14930 1790
rect 14730 1675 14810 1715
rect 14850 1675 14930 1715
rect 14730 1590 14930 1675
rect 15080 1715 15280 1790
rect 15080 1675 15160 1715
rect 15200 1675 15280 1715
rect 15080 1590 15280 1675
rect 15430 1715 15630 1790
rect 15430 1675 15510 1715
rect 15550 1675 15630 1715
rect 15430 1590 15630 1675
rect 14380 1365 14580 1440
rect 14380 1325 14460 1365
rect 14500 1325 14580 1365
rect 14380 1240 14580 1325
rect 14730 1365 14930 1440
rect 14730 1325 14810 1365
rect 14850 1325 14930 1365
rect 14730 1240 14930 1325
rect 15080 1365 15280 1440
rect 15080 1325 15160 1365
rect 15200 1325 15280 1365
rect 15080 1240 15280 1325
rect 15430 1365 15630 1440
rect 15430 1325 15510 1365
rect 15550 1325 15630 1365
rect 15430 1240 15630 1325
rect 14380 1015 14580 1090
rect 14380 975 14460 1015
rect 14500 975 14580 1015
rect 14380 890 14580 975
rect 14730 1015 14930 1090
rect 14730 975 14810 1015
rect 14850 975 14930 1015
rect 14730 890 14930 975
rect 15080 1015 15280 1090
rect 15080 975 15160 1015
rect 15200 975 15280 1015
rect 15080 890 15280 975
rect 15430 1015 15630 1090
rect 15430 975 15510 1015
rect 15550 975 15630 1015
rect 15430 890 15630 975
rect 14380 665 14580 740
rect 14380 625 14460 665
rect 14500 625 14580 665
rect 14380 540 14580 625
rect 14730 665 14930 740
rect 14730 625 14810 665
rect 14850 625 14930 665
rect 14730 540 14930 625
rect 15080 665 15280 740
rect 15080 625 15160 665
rect 15200 625 15280 665
rect 15080 540 15280 625
rect 15430 665 15630 740
rect 15430 625 15510 665
rect 15550 625 15630 665
rect 15430 540 15630 625
rect 11930 315 12130 390
rect 11930 275 12010 315
rect 12050 275 12130 315
rect 11930 190 12130 275
rect 12280 315 12480 390
rect 12280 275 12360 315
rect 12400 275 12480 315
rect 12280 190 12480 275
rect 12630 315 12830 390
rect 12630 275 12710 315
rect 12750 275 12830 315
rect 12630 190 12830 275
rect 12980 315 13180 390
rect 12980 275 13060 315
rect 13100 275 13180 315
rect 12980 190 13180 275
rect 13330 315 13530 390
rect 13330 275 13410 315
rect 13450 275 13530 315
rect 13330 190 13530 275
rect 13680 315 13880 390
rect 13680 275 13760 315
rect 13800 275 13880 315
rect 13680 190 13880 275
rect 14030 315 14230 390
rect 14030 275 14110 315
rect 14150 275 14230 315
rect 14030 190 14230 275
rect 14380 315 14580 390
rect 14380 275 14460 315
rect 14500 275 14580 315
rect 14380 190 14580 275
rect 14730 315 14930 390
rect 14730 275 14810 315
rect 14850 275 14930 315
rect 14730 190 14930 275
rect 15080 315 15280 390
rect 15080 275 15160 315
rect 15200 275 15280 315
rect 15080 190 15280 275
rect 15430 315 15630 390
rect 15430 275 15510 315
rect 15550 275 15630 315
rect 15430 190 15630 275
rect 11930 -35 12130 40
rect 11930 -75 12010 -35
rect 12050 -75 12130 -35
rect 11930 -160 12130 -75
rect 12280 -35 12480 40
rect 12280 -75 12360 -35
rect 12400 -75 12480 -35
rect 12280 -160 12480 -75
rect 12630 -35 12830 40
rect 12630 -75 12710 -35
rect 12750 -75 12830 -35
rect 12630 -160 12830 -75
rect 12980 -35 13180 40
rect 12980 -75 13060 -35
rect 13100 -75 13180 -35
rect 12980 -160 13180 -75
rect 13330 -35 13530 40
rect 13330 -75 13410 -35
rect 13450 -75 13530 -35
rect 13330 -160 13530 -75
rect 13680 -35 13880 40
rect 13680 -75 13760 -35
rect 13800 -75 13880 -35
rect 13680 -160 13880 -75
rect 14030 -35 14230 40
rect 14030 -75 14110 -35
rect 14150 -75 14230 -35
rect 14030 -160 14230 -75
rect 14380 -35 14580 40
rect 14380 -75 14460 -35
rect 14500 -75 14580 -35
rect 14380 -160 14580 -75
rect 14730 -35 14930 40
rect 14730 -75 14810 -35
rect 14850 -75 14930 -35
rect 14730 -160 14930 -75
rect 15080 -35 15280 40
rect 15080 -75 15160 -35
rect 15200 -75 15280 -35
rect 15080 -160 15280 -75
rect 15430 -35 15630 40
rect 15430 -75 15510 -35
rect 15550 -75 15630 -35
rect 15430 -160 15630 -75
rect 11930 -385 12130 -310
rect 11930 -425 12010 -385
rect 12050 -425 12130 -385
rect 11930 -510 12130 -425
rect 12280 -385 12480 -310
rect 12280 -425 12360 -385
rect 12400 -425 12480 -385
rect 12280 -510 12480 -425
rect 12630 -385 12830 -310
rect 12630 -425 12710 -385
rect 12750 -425 12830 -385
rect 12630 -510 12830 -425
rect 12980 -385 13180 -310
rect 12980 -425 13060 -385
rect 13100 -425 13180 -385
rect 12980 -510 13180 -425
rect 13330 -385 13530 -310
rect 13330 -425 13410 -385
rect 13450 -425 13530 -385
rect 13330 -510 13530 -425
rect 13680 -385 13880 -310
rect 13680 -425 13760 -385
rect 13800 -425 13880 -385
rect 13680 -510 13880 -425
rect 14030 -385 14230 -310
rect 14030 -425 14110 -385
rect 14150 -425 14230 -385
rect 14030 -510 14230 -425
rect 14380 -385 14580 -310
rect 14380 -425 14460 -385
rect 14500 -425 14580 -385
rect 14380 -510 14580 -425
rect 14730 -385 14930 -310
rect 14730 -425 14810 -385
rect 14850 -425 14930 -385
rect 14730 -510 14930 -425
rect 15080 -385 15280 -310
rect 15080 -425 15160 -385
rect 15200 -425 15280 -385
rect 15080 -510 15280 -425
rect 15430 -385 15630 -310
rect 15430 -425 15510 -385
rect 15550 -425 15630 -385
rect 15430 -510 15630 -425
<< mimcapcontact >>
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 5140 4725 5180 4765
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 5140 4375 5180 4415
rect 13060 4475 13100 4515
rect 13410 4475 13450 4515
rect 13760 4475 13800 4515
rect 14110 4475 14150 4515
rect 14460 4475 14500 4515
rect 14810 4475 14850 4515
rect 15160 4475 15200 4515
rect 15510 4475 15550 4515
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 5140 4025 5180 4065
rect 13060 4125 13100 4165
rect 13410 4125 13450 4165
rect 13760 4125 13800 4165
rect 14110 4125 14150 4165
rect 14460 4125 14500 4165
rect 14810 4125 14850 4165
rect 15160 4125 15200 4165
rect 15510 4125 15550 4165
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 5140 3675 5180 3715
rect 13060 3775 13100 3815
rect 13410 3775 13450 3815
rect 13760 3775 13800 3815
rect 14110 3775 14150 3815
rect 14460 3775 14500 3815
rect 14810 3775 14850 3815
rect 15160 3775 15200 3815
rect 15510 3775 15550 3815
rect 14460 3425 14500 3465
rect 14810 3425 14850 3465
rect 15160 3425 15200 3465
rect 15510 3425 15550 3465
rect 14460 3075 14500 3115
rect 14810 3075 14850 3115
rect 15160 3075 15200 3115
rect 15510 3075 15550 3115
rect 14460 2725 14500 2765
rect 14810 2725 14850 2765
rect 15160 2725 15200 2765
rect 15510 2725 15550 2765
rect 14460 2375 14500 2415
rect 14810 2375 14850 2415
rect 15160 2375 15200 2415
rect 15510 2375 15550 2415
rect 14460 2025 14500 2065
rect 14810 2025 14850 2065
rect 15160 2025 15200 2065
rect 15510 2025 15550 2065
rect 14460 1675 14500 1715
rect 14810 1675 14850 1715
rect 15160 1675 15200 1715
rect 15510 1675 15550 1715
rect 14460 1325 14500 1365
rect 14810 1325 14850 1365
rect 15160 1325 15200 1365
rect 15510 1325 15550 1365
rect 14460 975 14500 1015
rect 14810 975 14850 1015
rect 15160 975 15200 1015
rect 15510 975 15550 1015
rect 14460 625 14500 665
rect 14810 625 14850 665
rect 15160 625 15200 665
rect 15510 625 15550 665
rect 12010 275 12050 315
rect 12360 275 12400 315
rect 12710 275 12750 315
rect 13060 275 13100 315
rect 13410 275 13450 315
rect 13760 275 13800 315
rect 14110 275 14150 315
rect 14460 275 14500 315
rect 14810 275 14850 315
rect 15160 275 15200 315
rect 15510 275 15550 315
rect 12010 -75 12050 -35
rect 12360 -75 12400 -35
rect 12710 -75 12750 -35
rect 13060 -75 13100 -35
rect 13410 -75 13450 -35
rect 13760 -75 13800 -35
rect 14110 -75 14150 -35
rect 14460 -75 14500 -35
rect 14810 -75 14850 -35
rect 15160 -75 15200 -35
rect 15510 -75 15550 -35
rect 12010 -425 12050 -385
rect 12360 -425 12400 -385
rect 12710 -425 12750 -385
rect 13060 -425 13100 -385
rect 13410 -425 13450 -385
rect 13760 -425 13800 -385
rect 14110 -425 14150 -385
rect 14460 -425 14500 -385
rect 14810 -425 14850 -385
rect 15160 -425 15200 -385
rect 15510 -425 15550 -385
<< metal4 >>
rect -200 4995 5595 5000
rect -200 4955 -195 4995
rect -155 4955 5550 4995
rect 5590 4955 5595 4995
rect -200 4950 5595 4955
rect -115 4910 5510 4915
rect -115 4870 -110 4910
rect -70 4870 5465 4910
rect 5505 4870 5510 4910
rect -115 4865 5510 4870
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 13055 4515 13105 4520
rect 13055 4475 13060 4515
rect 13100 4475 13105 4515
rect 13055 4470 13105 4475
rect 13405 4515 13455 4520
rect 13405 4475 13410 4515
rect 13450 4475 13455 4515
rect 13405 4470 13455 4475
rect 13755 4515 13805 4520
rect 13755 4475 13760 4515
rect 13800 4475 13805 4515
rect 13755 4470 13805 4475
rect 14105 4515 14155 4520
rect 14105 4475 14110 4515
rect 14150 4475 14155 4515
rect 14105 4470 14155 4475
rect 14455 4515 14505 4520
rect 14455 4475 14460 4515
rect 14500 4475 14505 4515
rect 14455 4470 14505 4475
rect 14805 4515 14855 4520
rect 14805 4475 14810 4515
rect 14850 4475 14855 4515
rect 14805 4470 14855 4475
rect 15155 4515 15205 4520
rect 15155 4475 15160 4515
rect 15200 4475 15205 4515
rect 15155 4470 15205 4475
rect 15505 4515 15555 4520
rect 15505 4475 15510 4515
rect 15550 4475 15555 4515
rect 15505 4470 15555 4475
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 13055 4165 13105 4170
rect 13055 4125 13060 4165
rect 13100 4125 13105 4165
rect 13055 4120 13105 4125
rect 13405 4165 13455 4170
rect 13405 4125 13410 4165
rect 13450 4125 13455 4165
rect 13405 4120 13455 4125
rect 13755 4165 13805 4170
rect 13755 4125 13760 4165
rect 13800 4125 13805 4165
rect 13755 4120 13805 4125
rect 14105 4165 14155 4170
rect 14105 4125 14110 4165
rect 14150 4125 14155 4165
rect 14105 4120 14155 4125
rect 14455 4165 14505 4170
rect 14455 4125 14460 4165
rect 14500 4125 14505 4165
rect 14455 4120 14505 4125
rect 14805 4165 14855 4170
rect 14805 4125 14810 4165
rect 14850 4125 14855 4165
rect 14805 4120 14855 4125
rect 15155 4165 15205 4170
rect 15155 4125 15160 4165
rect 15200 4125 15205 4165
rect 15155 4120 15205 4125
rect 15505 4165 15555 4170
rect 15505 4125 15510 4165
rect 15550 4125 15555 4165
rect 15505 4120 15555 4125
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 13055 3815 13105 3820
rect 13055 3775 13060 3815
rect 13100 3775 13105 3815
rect 13055 3770 13105 3775
rect 13405 3815 13455 3820
rect 13405 3775 13410 3815
rect 13450 3775 13455 3815
rect 13405 3770 13455 3775
rect 13755 3815 13805 3820
rect 13755 3775 13760 3815
rect 13800 3775 13805 3815
rect 13755 3770 13805 3775
rect 14105 3815 14155 3820
rect 14105 3775 14110 3815
rect 14150 3775 14155 3815
rect 14105 3770 14155 3775
rect 14455 3815 14505 3820
rect 14455 3775 14460 3815
rect 14500 3775 14505 3815
rect 14455 3770 14505 3775
rect 14805 3815 14855 3820
rect 14805 3775 14810 3815
rect 14850 3775 14855 3815
rect 14805 3770 14855 3775
rect 15155 3815 15205 3820
rect 15155 3775 15160 3815
rect 15200 3775 15205 3815
rect 15155 3770 15205 3775
rect 15505 3815 15555 3820
rect 15505 3775 15510 3815
rect 15550 3775 15555 3815
rect 15505 3770 15555 3775
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 14455 3465 14505 3470
rect 14455 3425 14460 3465
rect 14500 3425 14505 3465
rect 14455 3420 14505 3425
rect 14805 3465 14855 3470
rect 14805 3425 14810 3465
rect 14850 3425 14855 3465
rect 14805 3420 14855 3425
rect 15155 3465 15205 3470
rect 15155 3425 15160 3465
rect 15200 3425 15205 3465
rect 15155 3420 15205 3425
rect 15505 3465 15555 3470
rect 15505 3425 15510 3465
rect 15550 3425 15555 3465
rect 15505 3420 15555 3425
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect 14455 3115 14505 3120
rect 14455 3075 14460 3115
rect 14500 3075 14505 3115
rect 14455 3070 14505 3075
rect 14805 3115 14855 3120
rect 14805 3075 14810 3115
rect 14850 3075 14855 3115
rect 14805 3070 14855 3075
rect 15155 3115 15205 3120
rect 15155 3075 15160 3115
rect 15200 3075 15205 3115
rect 15155 3070 15205 3075
rect 15505 3115 15555 3120
rect 15505 3075 15510 3115
rect 15550 3075 15555 3115
rect 15505 3070 15555 3075
rect 14455 2765 14505 2770
rect 14455 2725 14460 2765
rect 14500 2725 14505 2765
rect 14455 2720 14505 2725
rect 14805 2765 14855 2770
rect 14805 2725 14810 2765
rect 14850 2725 14855 2765
rect 14805 2720 14855 2725
rect 15155 2765 15205 2770
rect 15155 2725 15160 2765
rect 15200 2725 15205 2765
rect 15155 2720 15205 2725
rect 15505 2765 15555 2770
rect 15505 2725 15510 2765
rect 15550 2725 15555 2765
rect 15505 2720 15555 2725
rect 14455 2415 14505 2420
rect 14455 2375 14460 2415
rect 14500 2375 14505 2415
rect 14455 2370 14505 2375
rect 14805 2415 14855 2420
rect 14805 2375 14810 2415
rect 14850 2375 14855 2415
rect 14805 2370 14855 2375
rect 15155 2415 15205 2420
rect 15155 2375 15160 2415
rect 15200 2375 15205 2415
rect 15155 2370 15205 2375
rect 15505 2415 15555 2420
rect 15505 2375 15510 2415
rect 15550 2375 15555 2415
rect 15505 2370 15555 2375
rect 14455 2065 14505 2070
rect 14455 2025 14460 2065
rect 14500 2025 14505 2065
rect 14455 2020 14505 2025
rect 14805 2065 14855 2070
rect 14805 2025 14810 2065
rect 14850 2025 14855 2065
rect 14805 2020 14855 2025
rect 15155 2065 15205 2070
rect 15155 2025 15160 2065
rect 15200 2025 15205 2065
rect 15155 2020 15205 2025
rect 15505 2065 15555 2070
rect 15505 2025 15510 2065
rect 15550 2025 15555 2065
rect 15505 2020 15555 2025
rect 14455 1715 14505 1720
rect 14455 1675 14460 1715
rect 14500 1675 14505 1715
rect 14455 1670 14505 1675
rect 14805 1715 14855 1720
rect 14805 1675 14810 1715
rect 14850 1675 14855 1715
rect 14805 1670 14855 1675
rect 15155 1715 15205 1720
rect 15155 1675 15160 1715
rect 15200 1675 15205 1715
rect 15155 1670 15205 1675
rect 15505 1715 15555 1720
rect 15505 1675 15510 1715
rect 15550 1675 15555 1715
rect 15505 1670 15555 1675
rect 14455 1365 14505 1370
rect 14455 1325 14460 1365
rect 14500 1325 14505 1365
rect 14455 1320 14505 1325
rect 14805 1365 14855 1370
rect 14805 1325 14810 1365
rect 14850 1325 14855 1365
rect 14805 1320 14855 1325
rect 15155 1365 15205 1370
rect 15155 1325 15160 1365
rect 15200 1325 15205 1365
rect 15155 1320 15205 1325
rect 15505 1365 15555 1370
rect 15505 1325 15510 1365
rect 15550 1325 15555 1365
rect 15505 1320 15555 1325
rect 14455 1015 14505 1020
rect 14455 975 14460 1015
rect 14500 975 14505 1015
rect 14455 970 14505 975
rect 14805 1015 14855 1020
rect 14805 975 14810 1015
rect 14850 975 14855 1015
rect 14805 970 14855 975
rect 15155 1015 15205 1020
rect 15155 975 15160 1015
rect 15200 975 15205 1015
rect 15155 970 15205 975
rect 15505 1015 15555 1020
rect 15505 975 15510 1015
rect 15550 975 15555 1015
rect 15505 970 15555 975
rect 14455 665 14505 670
rect -115 660 5510 665
rect -115 620 -110 660
rect -70 620 5465 660
rect 5505 620 5510 660
rect 14455 625 14460 665
rect 14500 625 14505 665
rect 14455 620 14505 625
rect 14805 665 14855 670
rect 14805 625 14810 665
rect 14850 625 14855 665
rect 14805 620 14855 625
rect 15155 665 15205 670
rect 15155 625 15160 665
rect 15200 625 15205 665
rect 15155 620 15205 625
rect 15505 665 15555 670
rect 15505 625 15510 665
rect 15550 625 15555 665
rect 15505 620 15555 625
rect -115 615 5510 620
rect -200 580 5595 585
rect -200 540 -195 580
rect -155 540 5550 580
rect 5590 540 5595 580
rect -200 535 5595 540
rect 12005 315 12055 320
rect 12005 275 12010 315
rect 12050 275 12055 315
rect 12005 270 12055 275
rect 12355 315 12405 320
rect 12355 275 12360 315
rect 12400 275 12405 315
rect 12355 270 12405 275
rect 12705 315 12755 320
rect 12705 275 12710 315
rect 12750 275 12755 315
rect 12705 270 12755 275
rect 13055 315 13105 320
rect 13055 275 13060 315
rect 13100 275 13105 315
rect 13055 270 13105 275
rect 13405 315 13455 320
rect 13405 275 13410 315
rect 13450 275 13455 315
rect 13405 270 13455 275
rect 13755 315 13805 320
rect 13755 275 13760 315
rect 13800 275 13805 315
rect 13755 270 13805 275
rect 14105 315 14155 320
rect 14105 275 14110 315
rect 14150 275 14155 315
rect 14105 270 14155 275
rect 14455 315 14505 320
rect 14455 275 14460 315
rect 14500 275 14505 315
rect 14455 270 14505 275
rect 14805 315 14855 320
rect 14805 275 14810 315
rect 14850 275 14855 315
rect 14805 270 14855 275
rect 15155 315 15205 320
rect 15155 275 15160 315
rect 15200 275 15205 315
rect 15155 270 15205 275
rect 15505 315 15555 320
rect 15505 275 15510 315
rect 15550 275 15555 315
rect 15505 270 15555 275
rect 12005 -35 12055 -30
rect 12005 -75 12010 -35
rect 12050 -75 12055 -35
rect 12005 -80 12055 -75
rect 12355 -35 12405 -30
rect 12355 -75 12360 -35
rect 12400 -75 12405 -35
rect 12355 -80 12405 -75
rect 12705 -35 12755 -30
rect 12705 -75 12710 -35
rect 12750 -75 12755 -35
rect 12705 -80 12755 -75
rect 13055 -35 13105 -30
rect 13055 -75 13060 -35
rect 13100 -75 13105 -35
rect 13055 -80 13105 -75
rect 13405 -35 13455 -30
rect 13405 -75 13410 -35
rect 13450 -75 13455 -35
rect 13405 -80 13455 -75
rect 13755 -35 13805 -30
rect 13755 -75 13760 -35
rect 13800 -75 13805 -35
rect 13755 -80 13805 -75
rect 14105 -35 14155 -30
rect 14105 -75 14110 -35
rect 14150 -75 14155 -35
rect 14105 -80 14155 -75
rect 14455 -35 14505 -30
rect 14455 -75 14460 -35
rect 14500 -75 14505 -35
rect 14455 -80 14505 -75
rect 14805 -35 14855 -30
rect 14805 -75 14810 -35
rect 14850 -75 14855 -35
rect 14805 -80 14855 -75
rect 15155 -35 15205 -30
rect 15155 -75 15160 -35
rect 15200 -75 15205 -35
rect 15155 -80 15205 -75
rect 15505 -35 15555 -30
rect 15505 -75 15510 -35
rect 15550 -75 15555 -35
rect 15505 -80 15555 -75
rect 12005 -385 12055 -380
rect 12005 -425 12010 -385
rect 12050 -425 12055 -385
rect 12005 -430 12055 -425
rect 12355 -385 12405 -380
rect 12355 -425 12360 -385
rect 12400 -425 12405 -385
rect 12355 -430 12405 -425
rect 12705 -385 12755 -380
rect 12705 -425 12710 -385
rect 12750 -425 12755 -385
rect 12705 -430 12755 -425
rect 13055 -385 13105 -380
rect 13055 -425 13060 -385
rect 13100 -425 13105 -385
rect 13055 -430 13105 -425
rect 13405 -385 13455 -380
rect 13405 -425 13410 -385
rect 13450 -425 13455 -385
rect 13405 -430 13455 -425
rect 13755 -385 13805 -380
rect 13755 -425 13760 -385
rect 13800 -425 13805 -385
rect 13755 -430 13805 -425
rect 14105 -385 14155 -380
rect 14105 -425 14110 -385
rect 14150 -425 14155 -385
rect 14105 -430 14155 -425
rect 14455 -385 14505 -380
rect 14455 -425 14460 -385
rect 14500 -425 14505 -385
rect 14455 -430 14505 -425
rect 14805 -385 14855 -380
rect 14805 -425 14810 -385
rect 14850 -425 14855 -385
rect 14805 -430 14855 -425
rect 15155 -385 15205 -380
rect 15155 -425 15160 -385
rect 15200 -425 15205 -385
rect 15155 -430 15205 -425
rect 15505 -385 15555 -380
rect 15505 -425 15510 -385
rect 15550 -425 15555 -385
rect 15505 -430 15555 -425
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal2 2950 1735 2950 1735 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2955 1590 2955 1590 1 FreeSans 400 0 0 80 Vin+
flabel metal2 2945 1845 2945 1845 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 3745 1530 3745 1530 3 FreeSans 400 0 40 0 V_p1
flabel metal1 2650 1155 2650 1155 3 FreeSans 400 0 200 0 START_UP
flabel metal2 3785 1785 3785 1785 5 FreeSans 400 0 0 -40 1st_Vout1
flabel metal2 455 3440 455 3440 1 FreeSans 400 0 0 40 cap_res1
flabel metal3 2730 3375 2730 3375 3 FreeSans 400 0 40 0 cap_res2
flabel metal1 2550 845 2550 845 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal2 5120 1590 5120 1590 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 4225 1785 4225 1785 5 FreeSans 400 0 0 -40 1st_Vout2
flabel metal2 5065 1845 5065 1845 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 4265 1530 4265 1530 7 FreeSans 400 0 -40 0 V_p2
flabel metal1 3275 350 3275 350 7 FreeSans 400 0 -400 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 3825 295 3825 295 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal1 4015 350 4015 350 3 FreeSans 400 0 200 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 4725 295 4725 295 5 FreeSans 400 0 0 -200 VB3_CUR_BIAS
port 6 s
flabel metal1 4985 1110 4985 1110 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 4115 3135 4115 3135 1 FreeSans 400 0 0 40 PFET_GATE_10uA
flabel metal2 6080 3075 6080 3075 1 FreeSans 400 0 0 200 VB1_CUR_BIAS
port 1 n
flabel metal2 6100 3020 6100 3020 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6080 2955 6080 2955 5 FreeSans 400 0 0 -200 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal2 6100 1745 6100 1745 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
flabel metal3 5590 4400 5590 4400 3 FreeSans 800 0 80 0 VDDA
port 4 e
flabel metal3 5505 4175 5505 4175 3 FreeSans 800 0 80 0 GNDA
port 2 e
flabel metal1 2180 1010 2180 1010 3 FreeSans 400 0 40 0 Vbe2
flabel poly 4635 2375 4635 2375 5 FreeSans 400 0 0 -40 V_TOP
<< end >>
