* PEX produced on Mon Feb 17 04:29:33 AM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_7.ext - technology: sky130A

.subckt phase_frequency_detector_magic F_REF F_VCO VDDA QA QB GNDA
X0 GNDA.t29 E.t3 QA.t2 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X1 a_4210_n7910.t1 before_Reset.t3 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X2 F.t2 QB_b.t3 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X3 GNDA.t32 QA.t3 QA_b.t0 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X4 GNDA.t25 Reset.t2 E_b.t2 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X5 VDDA.t14 E.t4 a_2350_n7910.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X6 a_4210_n7910.t0 before_Reset.t4 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X7 GNDA.t1 E_b.t3 E.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X8 before_Reset.t0 QA.t4 a_3770_n7290.t1 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X9 VDDA.t24 F.t3 a_2350_n8670.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X10 GNDA.t42 a_4060_n9120.t2 a_3730_n9120.t0 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X11 GNDA.t36 a_4390_n9120.t2 a_4060_n9120.t1 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X12 QA_b.t1 QA.t5 a_1830_n7910.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X13 VDDA.t23 Reset.t3 a_3250_n7910.t1 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X14 QB_b.t0 QB.t3 a_1830_n8670.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X15 E.t1 E_b.t4 a_2730_n7910.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X16 VDDA.t16 QA.t6 before_Reset.t1 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X17 VDDA.t22 Reset.t4 a_3250_n8670.t0 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X18 F.t0 F_b.t3 a_2730_n8670.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X19 GNDA.t3 a_3730_n9120.t2 Reset.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X20 QA.t0 QA_b.t3 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X21 a_4390_n9120.t0 a_4210_n7910.t2 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X22 QA_b.t2 F_REF.t0 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X23 E_b.t1 E.t5 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X24 E.t2 QA_b.t4 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X25 a_3770_n7290.t0 QB.t4 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X26 a_2350_n7910.t1 QA_b.t5 QA.t1 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X27 a_4390_n9120.t1 a_4210_n7910.t3 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X28 a_1830_n7910.t0 F_REF.t1 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X29 a_2350_n8670.t0 QB_b.t4 QB.t1 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X30 a_3250_n7910.t0 E.t6 E_b.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X31 a_2730_n7910.t1 QA_b.t6 VDDA.t25 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X32 a_1830_n8670.t1 F_VCO.t0 VDDA.t6 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X33 a_3250_n8670.t1 F.t4 F_b.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X34 GNDA.t17 F.t5 QB.t2 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X35 before_Reset.t2 QB.t5 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X36 a_2730_n8670.t1 QB_b.t5 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X37 GNDA.t38 QB.t6 QB_b.t2 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X38 GNDA.t21 Reset.t5 F_b.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X39 GNDA.t15 F_b.t4 F.t1 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X40 VDDA.t27 a_4060_n9120.t3 a_3730_n9120.t1 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X41 VDDA.t8 a_4390_n9120.t3 a_4060_n9120.t0 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X42 VDDA.t2 a_3730_n9120.t3 Reset.t1 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X43 QB.t0 QB_b.t6 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X44 QB_b.t1 F_VCO.t1 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X45 F_b.t2 F.t6 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
R0 E.n4 E.n0 1319.38
R1 E.n0 E.t6 562.333
R2 E.n2 E.t4 388.813
R3 E.n2 E.t3 356.68
R4 E.n3 E.n2 232
R5 E.n0 E.t5 224.934
R6 E.t1 E.n4 221.411
R7 E.n3 E.n1 157.278
R8 E.n4 E.n3 90.64
R9 E.n1 E.t0 24.0005
R10 E.n1 E.t2 24.0005
R11 QA.t4 QA.t6 835.467
R12 QA.n2 QA.t5 517.347
R13 QA QA.t4 450.418
R14 QA.n1 QA.n0 244.715
R15 QA.n2 QA.t3 228.148
R16 QA.n1 QA.t1 221.411
R17 QA.n3 QA.n2 216
R18 QA.n3 QA.n1 201.573
R19 QA QA.n3 60.8005
R20 QA.n0 QA.t2 24.0005
R21 QA.n0 QA.t0 24.0005
R22 GNDA.n89 GNDA.n88 21560
R23 GNDA.t26 GNDA.t0 3006.67
R24 GNDA.t4 GNDA.t31 3006.67
R25 GNDA.t6 GNDA.t14 3006.67
R26 GNDA.t39 GNDA.t37 3006.67
R27 GNDA.t2 GNDA.n92 1943.33
R28 GNDA.t35 GNDA.n19 1575
R29 GNDA.n37 GNDA.t18 1430
R30 GNDA.n36 GNDA.t30 1430
R31 GNDA.n94 GNDA.t35 1430
R32 GNDA.t41 GNDA.n93 1430
R33 GNDA.n54 GNDA.n50 1026.67
R34 GNDA.n37 GNDA.t8 990
R35 GNDA.t18 GNDA.n36 990
R36 GNDA.n50 GNDA.t22 990
R37 GNDA.n54 GNDA.t24 990
R38 GNDA.t12 GNDA.n53 990
R39 GNDA.n53 GNDA.t28 990
R40 GNDA.n88 GNDA.t43 990
R41 GNDA.n94 GNDA.t41 990
R42 GNDA.n93 GNDA.t2 990
R43 GNDA.n92 GNDA.t20 990
R44 GNDA.t33 GNDA.n91 990
R45 GNDA.n91 GNDA.t16 990
R46 GNDA.t10 GNDA.n89 990
R47 GNDA.t30 GNDA.t22 806.668
R48 GNDA.t24 GNDA.t26 806.668
R49 GNDA.t0 GNDA.t12 806.668
R50 GNDA.t28 GNDA.t4 806.668
R51 GNDA.t31 GNDA.t43 806.668
R52 GNDA.t20 GNDA.t6 806.668
R53 GNDA.t14 GNDA.t33 806.668
R54 GNDA.t16 GNDA.t39 806.668
R55 GNDA.t37 GNDA.t10 806.668
R56 GNDA.n91 GNDA.n90 585.003
R57 GNDA.n53 GNDA.n52 585.003
R58 GNDA.n38 GNDA.n37 585.001
R59 GNDA.n55 GNDA.n54 585.001
R60 GNDA.n50 GNDA.n49 585.001
R61 GNDA.n36 GNDA.n35 585.001
R62 GNDA.n88 GNDA.n87 585.001
R63 GNDA.n95 GNDA.n94 585.001
R64 GNDA.n93 GNDA.n16 585.001
R65 GNDA.n92 GNDA.n13 585.001
R66 GNDA.n89 GNDA.n2 585.001
R67 GNDA.n3 GNDA.t38 198.058
R68 GNDA.n129 GNDA.t40 198.058
R69 GNDA.n117 GNDA.t15 198.058
R70 GNDA.n11 GNDA.t7 198.058
R71 GNDA.n81 GNDA.t32 198.058
R72 GNDA.n22 GNDA.t5 198.058
R73 GNDA.n67 GNDA.t1 198.058
R74 GNDA.n62 GNDA.t27 198.058
R75 GNDA.n7 GNDA.t17 130.713
R76 GNDA.n13 GNDA.t21 130.001
R77 GNDA.n16 GNDA.t3 130.001
R78 GNDA.n95 GNDA.t42 130.001
R79 GNDA.n19 GNDA.t36 130.001
R80 GNDA.n87 GNDA.t44 130.001
R81 GNDA.n55 GNDA.t25 130.001
R82 GNDA.n49 GNDA.t23 130.001
R83 GNDA.n35 GNDA.t19 130.001
R84 GNDA.n38 GNDA.t9 130.001
R85 GNDA.n2 GNDA.t11 130.001
R86 GNDA.n8 GNDA.t34 130.001
R87 GNDA.n51 GNDA.t13 130.001
R88 GNDA.n24 GNDA.t29 130.001
R89 GNDA.n19 GNDA.n18 70.3675
R90 GNDA.n39 GNDA.n38 68.9179
R91 GNDA.n109 GNDA.n13 60.29
R92 GNDA.n102 GNDA.n16 60.29
R93 GNDA.n96 GNDA.n95 60.29
R94 GNDA.n87 GNDA.n86 60.29
R95 GNDA.n56 GNDA.n55 60.29
R96 GNDA.n49 GNDA.n48 60.29
R97 GNDA.n35 GNDA.n34 60.29
R98 GNDA.n137 GNDA.n2 60.29
R99 GNDA.n122 GNDA.n8 54.4005
R100 GNDA.n124 GNDA.n7 54.4005
R101 GNDA.n73 GNDA.n24 54.4005
R102 GNDA.n51 GNDA.n25 54.4005
R103 GNDA.n86 GNDA.n0 33.0991
R104 GNDA.n138 GNDA.n137 33.0991
R105 GNDA.n42 GNDA.n41 32.0005
R106 GNDA.n43 GNDA.n42 32.0005
R107 GNDA.n43 GNDA.n32 32.0005
R108 GNDA.n57 GNDA.n31 32.0005
R109 GNDA.n61 GNDA.n29 32.0005
R110 GNDA.n62 GNDA.n61 32.0005
R111 GNDA.n63 GNDA.n62 32.0005
R112 GNDA.n63 GNDA.n27 32.0005
R113 GNDA.n67 GNDA.n27 32.0005
R114 GNDA.n68 GNDA.n67 32.0005
R115 GNDA.n69 GNDA.n68 32.0005
R116 GNDA.n75 GNDA.n74 32.0005
R117 GNDA.n75 GNDA.n22 32.0005
R118 GNDA.n79 GNDA.n22 32.0005
R119 GNDA.n80 GNDA.n79 32.0005
R120 GNDA.n81 GNDA.n80 32.0005
R121 GNDA.n81 GNDA.n20 32.0005
R122 GNDA.n85 GNDA.n20 32.0005
R123 GNDA.n97 GNDA.n17 32.0005
R124 GNDA.n101 GNDA.n17 32.0005
R125 GNDA.n104 GNDA.n103 32.0005
R126 GNDA.n104 GNDA.n14 32.0005
R127 GNDA.n108 GNDA.n14 32.0005
R128 GNDA.n111 GNDA.n110 32.0005
R129 GNDA.n111 GNDA.n11 32.0005
R130 GNDA.n115 GNDA.n11 32.0005
R131 GNDA.n116 GNDA.n115 32.0005
R132 GNDA.n117 GNDA.n116 32.0005
R133 GNDA.n117 GNDA.n9 32.0005
R134 GNDA.n121 GNDA.n9 32.0005
R135 GNDA.n125 GNDA.n5 32.0005
R136 GNDA.n129 GNDA.n5 32.0005
R137 GNDA.n130 GNDA.n129 32.0005
R138 GNDA.n131 GNDA.n130 32.0005
R139 GNDA.n131 GNDA.n3 32.0005
R140 GNDA.n135 GNDA.n3 32.0005
R141 GNDA.n136 GNDA.n135 32.0005
R142 GNDA.n47 GNDA.n31 28.8005
R143 GNDA.n41 GNDA.n34 25.6005
R144 GNDA.n57 GNDA.n56 25.6005
R145 GNDA.n72 GNDA.n25 25.6005
R146 GNDA.n73 GNDA.n72 25.6005
R147 GNDA.n102 GNDA.n101 25.6005
R148 GNDA.n109 GNDA.n108 25.6005
R149 GNDA.n123 GNDA.n122 25.6005
R150 GNDA.n96 GNDA.n18 23.4035
R151 GNDA.n124 GNDA.n123 22.4005
R152 GNDA.n48 GNDA.n32 19.2005
R153 GNDA.n97 GNDA.n96 16.0005
R154 GNDA.n39 GNDA.n34 13.8517
R155 GNDA GNDA.n0 12.7806
R156 GNDA GNDA.n138 11.8876
R157 GNDA.n48 GNDA.n47 9.6005
R158 GNDA.n125 GNDA.n124 9.6005
R159 GNDA.n41 GNDA.n40 9.3005
R160 GNDA.n42 GNDA.n33 9.3005
R161 GNDA.n44 GNDA.n43 9.3005
R162 GNDA.n45 GNDA.n32 9.3005
R163 GNDA.n47 GNDA.n46 9.3005
R164 GNDA.n31 GNDA.n30 9.3005
R165 GNDA.n58 GNDA.n57 9.3005
R166 GNDA.n59 GNDA.n29 9.3005
R167 GNDA.n61 GNDA.n60 9.3005
R168 GNDA.n62 GNDA.n28 9.3005
R169 GNDA.n64 GNDA.n63 9.3005
R170 GNDA.n65 GNDA.n27 9.3005
R171 GNDA.n67 GNDA.n66 9.3005
R172 GNDA.n68 GNDA.n26 9.3005
R173 GNDA.n70 GNDA.n69 9.3005
R174 GNDA.n72 GNDA.n71 9.3005
R175 GNDA.n74 GNDA.n23 9.3005
R176 GNDA.n76 GNDA.n75 9.3005
R177 GNDA.n77 GNDA.n22 9.3005
R178 GNDA.n79 GNDA.n78 9.3005
R179 GNDA.n80 GNDA.n21 9.3005
R180 GNDA.n82 GNDA.n81 9.3005
R181 GNDA.n83 GNDA.n20 9.3005
R182 GNDA.n85 GNDA.n84 9.3005
R183 GNDA.n98 GNDA.n97 9.3005
R184 GNDA.n99 GNDA.n17 9.3005
R185 GNDA.n101 GNDA.n100 9.3005
R186 GNDA.n103 GNDA.n15 9.3005
R187 GNDA.n105 GNDA.n104 9.3005
R188 GNDA.n106 GNDA.n14 9.3005
R189 GNDA.n108 GNDA.n107 9.3005
R190 GNDA.n110 GNDA.n12 9.3005
R191 GNDA.n112 GNDA.n111 9.3005
R192 GNDA.n113 GNDA.n11 9.3005
R193 GNDA.n115 GNDA.n114 9.3005
R194 GNDA.n116 GNDA.n10 9.3005
R195 GNDA.n118 GNDA.n117 9.3005
R196 GNDA.n119 GNDA.n9 9.3005
R197 GNDA.n121 GNDA.n120 9.3005
R198 GNDA.n123 GNDA.n6 9.3005
R199 GNDA.n126 GNDA.n125 9.3005
R200 GNDA.n127 GNDA.n5 9.3005
R201 GNDA.n129 GNDA.n128 9.3005
R202 GNDA.n130 GNDA.n4 9.3005
R203 GNDA.n132 GNDA.n131 9.3005
R204 GNDA.n133 GNDA.n3 9.3005
R205 GNDA.n135 GNDA.n134 9.3005
R206 GNDA.n136 GNDA.n1 9.3005
R207 GNDA.n56 GNDA.n29 6.4005
R208 GNDA.n69 GNDA.n25 6.4005
R209 GNDA.n74 GNDA.n73 6.4005
R210 GNDA.n86 GNDA.n85 6.4005
R211 GNDA.n103 GNDA.n102 6.4005
R212 GNDA.n110 GNDA.n109 6.4005
R213 GNDA.n122 GNDA.n121 6.4005
R214 GNDA.n137 GNDA.n136 6.4005
R215 GNDA.n90 GNDA.n8 5.68939
R216 GNDA.n52 GNDA.n51 5.68939
R217 GNDA.n52 GNDA.n24 5.68939
R218 GNDA.n90 GNDA.n7 4.97828
R219 GNDA.n98 GNDA.n18 0.289336
R220 GNDA.n40 GNDA.n39 0.241128
R221 GNDA.n84 GNDA.n0 0.193881
R222 GNDA.n138 GNDA.n1 0.193881
R223 GNDA.n40 GNDA.n33 0.15675
R224 GNDA.n44 GNDA.n33 0.15675
R225 GNDA.n45 GNDA.n44 0.15675
R226 GNDA.n58 GNDA.n30 0.15675
R227 GNDA.n59 GNDA.n58 0.15675
R228 GNDA.n60 GNDA.n59 0.15675
R229 GNDA.n60 GNDA.n28 0.15675
R230 GNDA.n64 GNDA.n28 0.15675
R231 GNDA.n65 GNDA.n64 0.15675
R232 GNDA.n66 GNDA.n65 0.15675
R233 GNDA.n66 GNDA.n26 0.15675
R234 GNDA.n70 GNDA.n26 0.15675
R235 GNDA.n71 GNDA.n70 0.15675
R236 GNDA.n71 GNDA.n23 0.15675
R237 GNDA.n76 GNDA.n23 0.15675
R238 GNDA.n77 GNDA.n76 0.15675
R239 GNDA.n78 GNDA.n77 0.15675
R240 GNDA.n78 GNDA.n21 0.15675
R241 GNDA.n82 GNDA.n21 0.15675
R242 GNDA.n83 GNDA.n82 0.15675
R243 GNDA.n84 GNDA.n83 0.15675
R244 GNDA.n99 GNDA.n98 0.15675
R245 GNDA.n100 GNDA.n99 0.15675
R246 GNDA.n100 GNDA.n15 0.15675
R247 GNDA.n105 GNDA.n15 0.15675
R248 GNDA.n106 GNDA.n105 0.15675
R249 GNDA.n107 GNDA.n106 0.15675
R250 GNDA.n107 GNDA.n12 0.15675
R251 GNDA.n112 GNDA.n12 0.15675
R252 GNDA.n113 GNDA.n112 0.15675
R253 GNDA.n114 GNDA.n113 0.15675
R254 GNDA.n114 GNDA.n10 0.15675
R255 GNDA.n118 GNDA.n10 0.15675
R256 GNDA.n119 GNDA.n118 0.15675
R257 GNDA.n120 GNDA.n119 0.15675
R258 GNDA.n120 GNDA.n6 0.15675
R259 GNDA.n126 GNDA.n6 0.15675
R260 GNDA.n127 GNDA.n126 0.15675
R261 GNDA.n128 GNDA.n127 0.15675
R262 GNDA.n128 GNDA.n4 0.15675
R263 GNDA.n132 GNDA.n4 0.15675
R264 GNDA.n133 GNDA.n132 0.15675
R265 GNDA.n134 GNDA.n133 0.15675
R266 GNDA.n134 GNDA.n1 0.15675
R267 GNDA.n46 GNDA.n45 0.141125
R268 GNDA.n46 GNDA.n30 0.141125
R269 before_Reset.n1 before_Reset.n0 481.334
R270 before_Reset.n0 before_Reset.t4 465.933
R271 before_Reset.n0 before_Reset.t3 321.334
R272 before_Reset.n2 before_Reset.n1 226.889
R273 before_Reset.n1 before_Reset.t0 172.458
R274 before_Reset.t1 before_Reset.n2 19.7005
R275 before_Reset.n2 before_Reset.t2 19.7005
R276 a_4210_n7910.t0 a_4210_n7910.n2 500.086
R277 a_4210_n7910.n1 a_4210_n7910.n0 473.334
R278 a_4210_n7910.n0 a_4210_n7910.t3 465.933
R279 a_4210_n7910.t0 a_4210_n7910.n2 461.389
R280 a_4210_n7910.n0 a_4210_n7910.t2 321.334
R281 a_4210_n7910.n1 a_4210_n7910.t1 177.577
R282 a_4210_n7910.n2 a_4210_n7910.n1 48.3899
R283 QB_b.t6 QB_b.t3 1188.93
R284 QB_b QB_b.n2 899.734
R285 QB_b.t3 QB_b.t5 835.467
R286 QB_b.n2 QB_b.t4 562.333
R287 QB_b QB_b.n1 419.647
R288 QB_b.n1 QB_b.n0 247.917
R289 QB_b.n2 QB_b.t6 224.934
R290 QB_b.n1 QB_b.t0 221.411
R291 QB_b.n0 QB_b.t2 24.0005
R292 QB_b.n0 QB_b.t1 24.0005
R293 F.n4 F.n0 1319.38
R294 F.n0 F.t4 562.333
R295 F.n2 F.t3 388.813
R296 F.n2 F.t5 356.68
R297 F.n3 F.n2 232
R298 F.n0 F.t6 224.934
R299 F.t0 F.n4 221.411
R300 F.n3 F.n1 157.278
R301 F.n4 F.n3 90.64
R302 F.n1 F.t1 24.0005
R303 F.n1 F.t2 24.0005
R304 QA_b.t3 QA_b.t4 1188.93
R305 QA_b QA_b.n2 837.38
R306 QA_b.t4 QA_b.t6 835.467
R307 QA_b.n0 QA_b.t5 562.333
R308 QA_b QA_b.n0 482
R309 QA_b.n2 QA_b.n1 247.917
R310 QA_b.n0 QA_b.t3 224.934
R311 QA_b.n2 QA_b.t1 221.411
R312 QA_b.n1 QA_b.t0 24.0005
R313 QA_b.n1 QA_b.t2 24.0005
R314 Reset.n1 Reset.t3 562.333
R315 Reset.n2 Reset.n1 480.45
R316 Reset.n0 Reset.t4 417.733
R317 Reset.n0 Reset.t5 369.534
R318 Reset.n3 Reset.n2 328.733
R319 Reset.t1 Reset.n3 288.37
R320 Reset.n1 Reset.t2 224.934
R321 Reset.n3 Reset.t0 177.577
R322 Reset.n2 Reset.n0 176.733
R323 E_b.n0 E_b.t4 517.347
R324 E_b.n2 E_b.n0 417.574
R325 E_b.n2 E_b.n1 244.716
R326 E_b.n0 E_b.t3 228.148
R327 E_b.t0 E_b.n2 221.411
R328 E_b.n1 E_b.t2 24.0005
R329 E_b.n1 E_b.t1 24.0005
R330 a_2350_n7910.t0 a_2350_n7910.t1 39.4005
R331 VDDA.n129 VDDA.n121 831.25
R332 VDDA.n124 VDDA.n123 831.25
R333 VDDA.n118 VDDA.n110 831.25
R334 VDDA.n113 VDDA.n112 831.25
R335 VDDA.n122 VDDA.n121 585
R336 VDDA.n126 VDDA.n124 585
R337 VDDA.n111 VDDA.n110 585
R338 VDDA.n115 VDDA.n113 585
R339 VDDA.n128 VDDA.t25 465.079
R340 VDDA.t25 VDDA.n127 465.079
R341 VDDA.n117 VDDA.t10 465.079
R342 VDDA.t10 VDDA.n116 465.079
R343 VDDA.t27 VDDA.n47 464.281
R344 VDDA.n49 VDDA.t27 464.281
R345 VDDA.t4 VDDA.n102 464.281
R346 VDDA.n103 VDDA.t4 464.281
R347 VDDA.n145 VDDA.t23 464.281
R348 VDDA.t23 VDDA.n144 464.281
R349 VDDA.n151 VDDA.t20 464.281
R350 VDDA.t20 VDDA.n18 464.281
R351 VDDA.n29 VDDA.t18 464.281
R352 VDDA.t18 VDDA.n26 464.281
R353 VDDA.n61 VDDA.t29 464.281
R354 VDDA.t29 VDDA.n60 464.281
R355 VDDA.t6 VDDA.n94 464.281
R356 VDDA.n95 VDDA.t6 464.281
R357 VDDA.t22 VDDA.n134 464.281
R358 VDDA.n135 VDDA.t22 464.281
R359 VDDA.n85 VDDA.t2 464.281
R360 VDDA.t2 VDDA.n84 464.281
R361 VDDA.t8 VDDA.n37 464.281
R362 VDDA.n39 VDDA.t8 464.281
R363 VDDA.n23 VDDA.t16 315.25
R364 VDDA.t12 VDDA.t5 314.113
R365 VDDA.t11 VDDA.t0 314.113
R366 VDDA.n102 VDDA.n91 243.698
R367 VDDA.n146 VDDA.n145 243.698
R368 VDDA.n152 VDDA.n151 243.698
R369 VDDA.n29 VDDA.n28 243.698
R370 VDDA.n62 VDDA.n61 243.698
R371 VDDA.n95 VDDA.n92 243.698
R372 VDDA.n135 VDDA.n132 243.698
R373 VDDA.n84 VDDA.n21 243.698
R374 VDDA.n43 VDDA.n39 243.698
R375 VDDA.n130 VDDA.n129 238.367
R376 VDDA.n123 VDDA.n90 238.367
R377 VDDA.n89 VDDA.n13 238.367
R378 VDDA.n155 VDDA.n154 238.367
R379 VDDA.n34 VDDA.n33 238.367
R380 VDDA.n57 VDDA.n44 238.367
R381 VDDA.n99 VDDA.n2 238.367
R382 VDDA.n119 VDDA.n118 238.367
R383 VDDA.n139 VDDA.n14 238.367
R384 VDDA.n87 VDDA.n86 238.367
R385 VDDA.n66 VDDA.n65 238.367
R386 VDDA.n112 VDDA.n108 238.367
R387 VDDA.n106 VDDA.n1 238.367
R388 VDDA.n49 VDDA.n46 190.333
R389 VDDA.n40 VDDA.n38 185
R390 VDDA.n42 VDDA.n41 185
R391 VDDA.n81 VDDA.n22 185
R392 VDDA.n83 VDDA.n82 185
R393 VDDA.n138 VDDA.n137 185
R394 VDDA.n136 VDDA.n133 185
R395 VDDA.n111 VDDA.n109 185
R396 VDDA.n115 VDDA.n114 185
R397 VDDA.n98 VDDA.n97 185
R398 VDDA.n96 VDDA.n93 185
R399 VDDA.n56 VDDA.n55 185
R400 VDDA.n59 VDDA.n58 185
R401 VDDA.n30 VDDA.n27 185
R402 VDDA.n32 VDDA.n31 185
R403 VDDA.n150 VDDA.n148 185
R404 VDDA.n149 VDDA.n19 185
R405 VDDA.n141 VDDA.n140 185
R406 VDDA.n143 VDDA.n142 185
R407 VDDA.n122 VDDA.n120 185
R408 VDDA.n126 VDDA.n125 185
R409 VDDA.n101 VDDA.n100 185
R410 VDDA.n105 VDDA.n104 185
R411 VDDA.n53 VDDA.n25 185
R412 VDDA.n54 VDDA.n53 185
R413 VDDA.n52 VDDA.n51 185
R414 VDDA.n50 VDDA.n48 185
R415 VDDA.n54 VDDA.n46 185
R416 VDDA.n105 VDDA.n100 150
R417 VDDA.n125 VDDA.n120 150
R418 VDDA.n142 VDDA.n140 150
R419 VDDA.n148 VDDA.n19 150
R420 VDDA.n32 VDDA.n27 150
R421 VDDA.n58 VDDA.n55 150
R422 VDDA.n98 VDDA.n93 150
R423 VDDA.n114 VDDA.n109 150
R424 VDDA.n138 VDDA.n133 150
R425 VDDA.n82 VDDA.n22 150
R426 VDDA.n42 VDDA.n38 150
R427 VDDA.n53 VDDA.n52 150
R428 VDDA.n48 VDDA.n46 150
R429 VDDA.n63 VDDA.n54 137.904
R430 VDDA.n88 VDDA.n20 137.904
R431 VDDA.t14 VDDA.n121 123.126
R432 VDDA.n124 VDDA.t14 123.126
R433 VDDA.t24 VDDA.n110 123.126
R434 VDDA.n113 VDDA.t24 123.126
R435 VDDA.n153 VDDA.n147 107.258
R436 VDDA.n147 VDDA.t21 103.427
R437 VDDA.t9 VDDA.n131 103.427
R438 VDDA.n131 VDDA.t13 103.427
R439 VDDA.t3 VDDA.n107 103.427
R440 VDDA.n153 VDDA.t1 95.7666
R441 VDDA.t28 VDDA.t7 91.936
R442 VDDA.t17 VDDA.t26 91.936
R443 VDDA.t19 VDDA.t15 84.2747
R444 VDDA.t21 VDDA.t12 84.2747
R445 VDDA.t5 VDDA.t9 84.2747
R446 VDDA.t13 VDDA.t11 84.2747
R447 VDDA.t0 VDDA.t3 84.2747
R448 VDDA.n65 VDDA.n64 65.8183
R449 VDDA.n64 VDDA.n43 65.8183
R450 VDDA.n88 VDDA.n87 65.8183
R451 VDDA.n88 VDDA.n21 65.8183
R452 VDDA.n147 VDDA.n139 65.8183
R453 VDDA.n147 VDDA.n132 65.8183
R454 VDDA.n131 VDDA.n119 65.8183
R455 VDDA.n131 VDDA.n108 65.8183
R456 VDDA.n107 VDDA.n99 65.8183
R457 VDDA.n107 VDDA.n92 65.8183
R458 VDDA.n63 VDDA.n62 65.8183
R459 VDDA.n63 VDDA.n44 65.8183
R460 VDDA.n28 VDDA.n20 65.8183
R461 VDDA.n33 VDDA.n20 65.8183
R462 VDDA.n153 VDDA.n152 65.8183
R463 VDDA.n154 VDDA.n153 65.8183
R464 VDDA.n147 VDDA.n146 65.8183
R465 VDDA.n147 VDDA.n89 65.8183
R466 VDDA.n131 VDDA.n130 65.8183
R467 VDDA.n131 VDDA.n90 65.8183
R468 VDDA.n107 VDDA.n91 65.8183
R469 VDDA.n107 VDDA.n106 65.8183
R470 VDDA.n54 VDDA.n45 65.8183
R471 VDDA.n57 VDDA.n36 60.4427
R472 VDDA.n190 VDDA.n1 58.0576
R473 VDDA.n162 VDDA.n13 58.0576
R474 VDDA.n156 VDDA.n155 58.0576
R475 VDDA.n73 VDDA.n34 58.0576
R476 VDDA.n190 VDDA.n2 58.0576
R477 VDDA.n162 VDDA.n14 58.0576
R478 VDDA.n86 VDDA.n80 58.0576
R479 VDDA.n67 VDDA.n66 58.0576
R480 VDDA.n74 VDDA.n25 58.0576
R481 VDDA.n177 VDDA.n7 54.4005
R482 VDDA.n175 VDDA.n7 54.4005
R483 VDDA.n175 VDDA.n8 54.4005
R484 VDDA.n177 VDDA.n8 54.4005
R485 VDDA.n100 VDDA.n91 53.3664
R486 VDDA.n106 VDDA.n105 53.3664
R487 VDDA.n93 VDDA.n92 53.3664
R488 VDDA.n114 VDDA.n108 53.3664
R489 VDDA.n133 VDDA.n132 53.3664
R490 VDDA.n65 VDDA.n38 53.3664
R491 VDDA.n43 VDDA.n42 53.3664
R492 VDDA.n87 VDDA.n22 53.3664
R493 VDDA.n82 VDDA.n21 53.3664
R494 VDDA.n139 VDDA.n138 53.3664
R495 VDDA.n119 VDDA.n109 53.3664
R496 VDDA.n99 VDDA.n98 53.3664
R497 VDDA.n62 VDDA.n55 53.3664
R498 VDDA.n58 VDDA.n44 53.3664
R499 VDDA.n28 VDDA.n27 53.3664
R500 VDDA.n33 VDDA.n32 53.3664
R501 VDDA.n152 VDDA.n148 53.3664
R502 VDDA.n154 VDDA.n19 53.3664
R503 VDDA.n146 VDDA.n140 53.3664
R504 VDDA.n142 VDDA.n89 53.3664
R505 VDDA.n130 VDDA.n120 53.3664
R506 VDDA.n125 VDDA.n90 53.3664
R507 VDDA.n52 VDDA.n45 53.3664
R508 VDDA.n48 VDDA.n45 53.3664
R509 VDDA.n191 VDDA.n190 34.9005
R510 VDDA.n68 VDDA.n67 32.0005
R511 VDDA.n68 VDDA.n35 32.0005
R512 VDDA.n72 VDDA.n35 32.0005
R513 VDDA.n76 VDDA.n75 32.0005
R514 VDDA.n161 VDDA.n15 32.0005
R515 VDDA.n164 VDDA.n163 32.0005
R516 VDDA.n164 VDDA.n11 32.0005
R517 VDDA.n168 VDDA.n11 32.0005
R518 VDDA.n169 VDDA.n168 32.0005
R519 VDDA.n170 VDDA.n169 32.0005
R520 VDDA.n170 VDDA.n9 32.0005
R521 VDDA.n174 VDDA.n9 32.0005
R522 VDDA.n178 VDDA.n5 32.0005
R523 VDDA.n182 VDDA.n5 32.0005
R524 VDDA.n183 VDDA.n182 32.0005
R525 VDDA.n184 VDDA.n183 32.0005
R526 VDDA.n184 VDDA.n3 32.0005
R527 VDDA.n188 VDDA.n3 32.0005
R528 VDDA.n189 VDDA.n188 32.0005
R529 VDDA.n157 VDDA.n17 28.8005
R530 VDDA.n156 VDDA.n15 25.6005
R531 VDDA.n162 VDDA.n161 25.6005
R532 VDDA.n176 VDDA.n175 25.6005
R533 VDDA.n177 VDDA.n176 25.6005
R534 VDDA.n75 VDDA.n74 22.4005
R535 VDDA.n79 VDDA.n23 19.2005
R536 VDDA.n80 VDDA.n79 19.2005
R537 VDDA.n76 VDDA.n23 12.8005
R538 VDDA.n80 VDDA.n17 12.8005
R539 VDDA.n64 VDDA.t28 11.4924
R540 VDDA.t7 VDDA.n63 11.4924
R541 VDDA.n54 VDDA.t17 11.4924
R542 VDDA.t26 VDDA.n20 11.4924
R543 VDDA.t15 VDDA.n88 11.4924
R544 VDDA.n69 VDDA.n68 9.3005
R545 VDDA.n70 VDDA.n35 9.3005
R546 VDDA.n72 VDDA.n71 9.3005
R547 VDDA.n75 VDDA.n24 9.3005
R548 VDDA.n77 VDDA.n76 9.3005
R549 VDDA.n79 VDDA.n78 9.3005
R550 VDDA.n17 VDDA.n16 9.3005
R551 VDDA.n158 VDDA.n157 9.3005
R552 VDDA.n159 VDDA.n15 9.3005
R553 VDDA.n161 VDDA.n160 9.3005
R554 VDDA.n163 VDDA.n12 9.3005
R555 VDDA.n165 VDDA.n164 9.3005
R556 VDDA.n166 VDDA.n11 9.3005
R557 VDDA.n168 VDDA.n167 9.3005
R558 VDDA.n169 VDDA.n10 9.3005
R559 VDDA.n171 VDDA.n170 9.3005
R560 VDDA.n172 VDDA.n9 9.3005
R561 VDDA.n174 VDDA.n173 9.3005
R562 VDDA.n176 VDDA.n6 9.3005
R563 VDDA.n179 VDDA.n178 9.3005
R564 VDDA.n180 VDDA.n5 9.3005
R565 VDDA.n182 VDDA.n181 9.3005
R566 VDDA.n183 VDDA.n4 9.3005
R567 VDDA.n185 VDDA.n184 9.3005
R568 VDDA.n186 VDDA.n3 9.3005
R569 VDDA.n188 VDDA.n187 9.3005
R570 VDDA.n189 VDDA.n0 9.3005
R571 VDDA.n104 VDDA.n101 9.14336
R572 VDDA.n143 VDDA.n141 9.14336
R573 VDDA.n150 VDDA.n149 9.14336
R574 VDDA.n31 VDDA.n30 9.14336
R575 VDDA.n59 VDDA.n56 9.14336
R576 VDDA.n97 VDDA.n96 9.14336
R577 VDDA.n137 VDDA.n136 9.14336
R578 VDDA.n83 VDDA.n81 9.14336
R579 VDDA.n41 VDDA.n40 9.14336
R580 VDDA.n51 VDDA.n50 9.14336
R581 VDDA.t1 VDDA.t19 7.66179
R582 VDDA.n69 VDDA.n36 7.08733
R583 VDDA.n73 VDDA.n72 6.4005
R584 VDDA.n163 VDDA.n162 6.4005
R585 VDDA.n175 VDDA.n174 6.4005
R586 VDDA.n178 VDDA.n177 6.4005
R587 VDDA.n190 VDDA.n189 6.4005
R588 VDDA.n126 VDDA.n122 5.81868
R589 VDDA.n115 VDDA.n111 5.81868
R590 VDDA.n47 VDDA.n25 5.33286
R591 VDDA.n103 VDDA.n1 5.33286
R592 VDDA.n144 VDDA.n13 5.33286
R593 VDDA.n155 VDDA.n18 5.33286
R594 VDDA.n34 VDDA.n26 5.33286
R595 VDDA.n60 VDDA.n57 5.33286
R596 VDDA.n94 VDDA.n2 5.33286
R597 VDDA.n134 VDDA.n14 5.33286
R598 VDDA.n86 VDDA.n85 5.33286
R599 VDDA.n66 VDDA.n37 5.33286
R600 VDDA.n102 VDDA.n101 3.75335
R601 VDDA.n104 VDDA.n103 3.75335
R602 VDDA.n145 VDDA.n141 3.75335
R603 VDDA.n144 VDDA.n143 3.75335
R604 VDDA.n151 VDDA.n150 3.75335
R605 VDDA.n149 VDDA.n18 3.75335
R606 VDDA.n30 VDDA.n29 3.75335
R607 VDDA.n31 VDDA.n26 3.75335
R608 VDDA.n61 VDDA.n56 3.75335
R609 VDDA.n60 VDDA.n59 3.75335
R610 VDDA.n97 VDDA.n94 3.75335
R611 VDDA.n96 VDDA.n95 3.75335
R612 VDDA.n137 VDDA.n134 3.75335
R613 VDDA.n136 VDDA.n135 3.75335
R614 VDDA.n85 VDDA.n81 3.75335
R615 VDDA.n84 VDDA.n83 3.75335
R616 VDDA.n40 VDDA.n37 3.75335
R617 VDDA.n41 VDDA.n39 3.75335
R618 VDDA.n51 VDDA.n47 3.75335
R619 VDDA.n50 VDDA.n49 3.75335
R620 VDDA.n129 VDDA.n128 3.40194
R621 VDDA.n127 VDDA.n123 3.40194
R622 VDDA.n118 VDDA.n117 3.40194
R623 VDDA.n116 VDDA.n112 3.40194
R624 VDDA.n74 VDDA.n73 3.2005
R625 VDDA.n157 VDDA.n156 3.2005
R626 VDDA.n128 VDDA.n122 2.39444
R627 VDDA.n127 VDDA.n126 2.39444
R628 VDDA.n117 VDDA.n111 2.39444
R629 VDDA.n116 VDDA.n115 2.39444
R630 VDDA.n123 VDDA.n7 2.32777
R631 VDDA.n118 VDDA.n8 2.32777
R632 VDDA.n67 VDDA.n36 0.6077
R633 VDDA.n70 VDDA.n69 0.15675
R634 VDDA.n71 VDDA.n70 0.15675
R635 VDDA.n71 VDDA.n24 0.15675
R636 VDDA.n77 VDDA.n24 0.15675
R637 VDDA.n78 VDDA.n77 0.15675
R638 VDDA.n78 VDDA.n16 0.15675
R639 VDDA.n160 VDDA.n159 0.15675
R640 VDDA.n160 VDDA.n12 0.15675
R641 VDDA.n165 VDDA.n12 0.15675
R642 VDDA.n166 VDDA.n165 0.15675
R643 VDDA.n167 VDDA.n166 0.15675
R644 VDDA.n167 VDDA.n10 0.15675
R645 VDDA.n171 VDDA.n10 0.15675
R646 VDDA.n172 VDDA.n171 0.15675
R647 VDDA.n173 VDDA.n172 0.15675
R648 VDDA.n173 VDDA.n6 0.15675
R649 VDDA.n179 VDDA.n6 0.15675
R650 VDDA.n180 VDDA.n179 0.15675
R651 VDDA.n181 VDDA.n180 0.15675
R652 VDDA.n181 VDDA.n4 0.15675
R653 VDDA.n185 VDDA.n4 0.15675
R654 VDDA.n186 VDDA.n185 0.15675
R655 VDDA.n187 VDDA.n186 0.15675
R656 VDDA.n187 VDDA.n0 0.15675
R657 VDDA.n191 VDDA.n0 0.15675
R658 VDDA.n158 VDDA.n16 0.141125
R659 VDDA.n159 VDDA.n158 0.141125
R660 VDDA VDDA.n191 0.1255
R661 a_3770_n7290.t0 a_3770_n7290.t1 48.0005
R662 a_2350_n8670.t0 a_2350_n8670.t1 39.4005
R663 a_4060_n9120.t0 a_4060_n9120.n2 500.086
R664 a_4060_n9120.n1 a_4060_n9120.n0 473.334
R665 a_4060_n9120.n0 a_4060_n9120.t3 465.933
R666 a_4060_n9120.t0 a_4060_n9120.n2 461.389
R667 a_4060_n9120.n0 a_4060_n9120.t2 321.334
R668 a_4060_n9120.n1 a_4060_n9120.t1 177.577
R669 a_4060_n9120.n2 a_4060_n9120.n1 48.3898
R670 a_3730_n9120.t1 a_3730_n9120.n2 500.086
R671 a_3730_n9120.n1 a_3730_n9120.n0 473.334
R672 a_3730_n9120.n0 a_3730_n9120.t3 465.933
R673 a_3730_n9120.t1 a_3730_n9120.n2 461.389
R674 a_3730_n9120.n0 a_3730_n9120.t2 321.334
R675 a_3730_n9120.n1 a_3730_n9120.t0 177.577
R676 a_3730_n9120.n2 a_3730_n9120.n1 48.3898
R677 a_4390_n9120.t1 a_4390_n9120.n2 500.086
R678 a_4390_n9120.n0 a_4390_n9120.t3 465.933
R679 a_4390_n9120.t1 a_4390_n9120.n2 461.389
R680 a_4390_n9120.n1 a_4390_n9120.n0 392.623
R681 a_4390_n9120.n0 a_4390_n9120.t2 321.334
R682 a_4390_n9120.n1 a_4390_n9120.t0 177.577
R683 a_4390_n9120.n2 a_4390_n9120.n1 48.3899
R684 a_1830_n7910.t0 a_1830_n7910.t1 39.4005
R685 a_3250_n7910.t0 a_3250_n7910.t1 39.4005
R686 QB.t5 QB.t4 835.467
R687 QB QB.t5 581.653
R688 QB.n0 QB.t3 517.347
R689 QB.n3 QB.n0 363.2
R690 QB.n2 QB.n1 244.716
R691 QB.n0 QB.t6 228.148
R692 QB.n2 QB.t1 221.411
R693 QB.n3 QB.n2 54.3734
R694 QB.n1 QB.t2 24.0005
R695 QB.n1 QB.t0 24.0005
R696 QB QB.n3 12.8005
R697 a_1830_n8670.t0 a_1830_n8670.t1 39.4005
R698 a_2730_n7910.t0 a_2730_n7910.t1 39.4005
R699 a_3250_n8670.t0 a_3250_n8670.t1 39.4005
R700 F_b.n0 F_b.t3 517.347
R701 F_b.n2 F_b.n0 417.574
R702 F_b.n2 F_b.n1 244.716
R703 F_b.n0 F_b.t4 228.148
R704 F_b.t1 F_b.n2 221.411
R705 F_b.n1 F_b.t0 24.0005
R706 F_b.n1 F_b.t2 24.0005
R707 a_2730_n8670.t0 a_2730_n8670.t1 39.4005
R708 F_REF.n0 F_REF.t1 514.134
R709 F_REF.n0 F_REF.t0 273.134
R710 F_REF F_REF.n0 216.9
R711 F_VCO.n0 F_VCO.t0 514.134
R712 F_VCO.n0 F_VCO.t1 273.134
R713 F_VCO F_VCO.n0 216.9
C0 QB F_VCO 0.056153f
C1 QB QA 0.068636f
C2 VDDA QB 2.25074f
C3 F_REF QA 0.056f
C4 QB_b F_VCO 0.026369f
C5 VDDA F_REF 0.085173f
C6 VDDA QB_b 0.513239f
C7 VDDA F_VCO 0.085127f
C8 VDDA QA 0.393128f
C9 F_REF QA_b 0.026369f
C10 QA_b QA 0.422694f
C11 VDDA QA_b 0.521329f
C12 QB_b QB 0.386189f
C13 F_VCO GNDA 0.236218f
C14 QB GNDA 1.49618f
C15 QA GNDA 2.60115f
C16 F_REF GNDA 0.236218f
C17 VDDA GNDA 11.876046f
C18 QB_b GNDA 1.06416f
C19 QA_b GNDA 1.05219f
C20 QB.t3 GNDA 0.087036f
C21 QB.t6 GNDA 0.038163f
C22 QB.n0 GNDA 0.219846f
C23 QB.t1 GNDA 0.183277f
C24 QB.t2 GNDA 0.034822f
C25 QB.t0 GNDA 0.034822f
C26 QB.n1 GNDA 0.185934f
C27 QB.n2 GNDA 0.330337f
C28 QB.n3 GNDA 0.285611f
C29 QB.t4 GNDA 0.086185f
C30 QB.t5 GNDA 0.145983f
C31 VDDA.n20 GNDA 0.047111f
C32 VDDA.t16 GNDA 0.011828f
C33 VDDA.n23 GNDA 0.012955f
C34 VDDA.t26 GNDA 0.032616f
C35 VDDA.t17 GNDA 0.032616f
C36 VDDA.n54 GNDA 0.047111f
C37 VDDA.n63 GNDA 0.047111f
C38 VDDA.t7 GNDA 0.032616f
C39 VDDA.t28 GNDA 0.032616f
C40 VDDA.n64 GNDA 0.080935f
C41 VDDA.n69 GNDA 0.014374f
C42 VDDA.n88 GNDA 0.047111f
C43 VDDA.t15 GNDA 0.0302f
C44 VDDA.t19 GNDA 0.028992f
C45 VDDA.t1 GNDA 0.032616f
C46 VDDA.n107 GNDA 0.071271f
C47 VDDA.t3 GNDA 0.059191f
C48 VDDA.t0 GNDA 0.12563f
C49 VDDA.t11 GNDA 0.12563f
C50 VDDA.t13 GNDA 0.059191f
C51 VDDA.n112 GNDA 0.01026f
C52 VDDA.n129 GNDA 0.01026f
C53 VDDA.n131 GNDA 0.065231f
C54 VDDA.t9 GNDA 0.059191f
C55 VDDA.t5 GNDA 0.12563f
C56 VDDA.t12 GNDA 0.12563f
C57 VDDA.t21 GNDA 0.059191f
C58 VDDA.n147 GNDA 0.066439f
C59 VDDA.n153 GNDA 0.064023f
.ends

