magic
tech sky130A
timestamp 1737822713
<< nmos >>
rect -850 350 -800 600
rect -750 350 -700 600
rect -650 350 -600 600
rect -550 350 -500 600
rect -450 350 -400 600
rect -350 350 -300 600
rect -250 350 -200 600
rect -150 350 -100 600
rect -450 0 -400 250
rect -350 0 -300 250
rect -250 0 -200 250
rect -150 0 -100 250
rect 300 190 315 240
rect 365 190 380 240
rect 430 190 445 240
rect 495 190 510 240
rect 560 190 575 240
rect 625 190 640 240
rect 690 190 705 240
rect 755 190 770 240
rect 900 190 915 240
rect 965 190 980 240
rect 1030 190 1045 240
rect 1095 190 1110 240
rect 1160 190 1175 240
rect 1225 190 1240 240
rect 1290 190 1305 240
rect 1355 190 1370 240
rect 1500 190 1515 240
rect 1565 190 1580 240
rect 1630 190 1645 240
rect 1695 190 1710 240
rect 1760 190 1775 240
rect 1825 190 1840 240
rect 1890 190 1905 240
rect 1955 190 1970 240
rect 300 -5 315 45
rect 365 -5 380 45
rect 430 -5 445 45
rect 495 -5 510 45
rect 640 -5 655 45
rect 705 -5 720 45
rect 770 -5 785 45
rect 835 -5 850 45
rect 980 -5 995 45
rect 1045 -5 1060 45
rect 1110 -5 1125 45
rect 1175 -5 1190 45
<< ndiff >>
rect -900 585 -850 600
rect -900 365 -885 585
rect -865 365 -850 585
rect -900 350 -850 365
rect -800 585 -750 600
rect -800 365 -785 585
rect -765 365 -750 585
rect -800 350 -750 365
rect -700 585 -650 600
rect -700 365 -685 585
rect -665 365 -650 585
rect -700 350 -650 365
rect -600 585 -550 600
rect -600 365 -585 585
rect -565 365 -550 585
rect -600 350 -550 365
rect -500 585 -450 600
rect -500 365 -485 585
rect -465 365 -450 585
rect -500 350 -450 365
rect -400 585 -350 600
rect -400 365 -385 585
rect -365 365 -350 585
rect -400 350 -350 365
rect -300 585 -250 600
rect -300 365 -285 585
rect -265 365 -250 585
rect -300 350 -250 365
rect -200 585 -150 600
rect -200 365 -185 585
rect -165 365 -150 585
rect -200 350 -150 365
rect -100 585 -50 600
rect -100 365 -85 585
rect -65 365 -50 585
rect -100 350 -50 365
rect -500 235 -450 250
rect -500 15 -485 235
rect -465 15 -450 235
rect -500 0 -450 15
rect -400 235 -350 250
rect -400 15 -385 235
rect -365 15 -350 235
rect -400 0 -350 15
rect -300 235 -250 250
rect -300 15 -285 235
rect -265 15 -250 235
rect -300 0 -250 15
rect -200 235 -150 250
rect -200 15 -185 235
rect -165 15 -150 235
rect -200 0 -150 15
rect -100 235 -50 250
rect -100 15 -85 235
rect -65 15 -50 235
rect 250 225 300 240
rect 250 205 265 225
rect 285 205 300 225
rect 250 190 300 205
rect 315 225 365 240
rect 315 205 330 225
rect 350 205 365 225
rect 315 190 365 205
rect 380 225 430 240
rect 380 205 395 225
rect 415 205 430 225
rect 380 190 430 205
rect 445 225 495 240
rect 445 205 460 225
rect 480 205 495 225
rect 445 190 495 205
rect 510 225 560 240
rect 510 205 525 225
rect 545 205 560 225
rect 510 190 560 205
rect 575 225 625 240
rect 575 205 590 225
rect 610 205 625 225
rect 575 190 625 205
rect 640 225 690 240
rect 640 205 655 225
rect 675 205 690 225
rect 640 190 690 205
rect 705 225 755 240
rect 705 205 720 225
rect 740 205 755 225
rect 705 190 755 205
rect 770 225 820 240
rect 770 205 785 225
rect 805 205 820 225
rect 770 190 820 205
rect 850 225 900 240
rect 850 205 865 225
rect 885 205 900 225
rect 850 190 900 205
rect 915 225 965 240
rect 915 205 930 225
rect 950 205 965 225
rect 915 190 965 205
rect 980 225 1030 240
rect 980 205 995 225
rect 1015 205 1030 225
rect 980 190 1030 205
rect 1045 225 1095 240
rect 1045 205 1060 225
rect 1080 205 1095 225
rect 1045 190 1095 205
rect 1110 225 1160 240
rect 1110 205 1125 225
rect 1145 205 1160 225
rect 1110 190 1160 205
rect 1175 225 1225 240
rect 1175 205 1190 225
rect 1210 205 1225 225
rect 1175 190 1225 205
rect 1240 225 1290 240
rect 1240 205 1255 225
rect 1275 205 1290 225
rect 1240 190 1290 205
rect 1305 225 1355 240
rect 1305 205 1320 225
rect 1340 205 1355 225
rect 1305 190 1355 205
rect 1370 225 1420 240
rect 1370 205 1385 225
rect 1405 205 1420 225
rect 1370 190 1420 205
rect 1450 225 1500 240
rect 1450 205 1465 225
rect 1485 205 1500 225
rect 1450 190 1500 205
rect 1515 225 1565 240
rect 1515 205 1530 225
rect 1550 205 1565 225
rect 1515 190 1565 205
rect 1580 225 1630 240
rect 1580 205 1595 225
rect 1615 205 1630 225
rect 1580 190 1630 205
rect 1645 225 1695 240
rect 1645 205 1660 225
rect 1680 205 1695 225
rect 1645 190 1695 205
rect 1710 225 1760 240
rect 1710 205 1725 225
rect 1745 205 1760 225
rect 1710 190 1760 205
rect 1775 225 1825 240
rect 1775 205 1790 225
rect 1810 205 1825 225
rect 1775 190 1825 205
rect 1840 225 1890 240
rect 1840 205 1855 225
rect 1875 205 1890 225
rect 1840 190 1890 205
rect 1905 225 1955 240
rect 1905 205 1920 225
rect 1940 205 1955 225
rect 1905 190 1955 205
rect 1970 225 2020 240
rect 1970 205 1985 225
rect 2005 205 2020 225
rect 1970 190 2020 205
rect -100 0 -50 15
rect 250 30 300 45
rect 250 10 265 30
rect 285 10 300 30
rect 250 -5 300 10
rect 315 30 365 45
rect 315 10 330 30
rect 350 10 365 30
rect 315 -5 365 10
rect 380 30 430 45
rect 380 10 395 30
rect 415 10 430 30
rect 380 -5 430 10
rect 445 30 495 45
rect 445 10 460 30
rect 480 10 495 30
rect 445 -5 495 10
rect 510 30 560 45
rect 510 10 525 30
rect 545 10 560 30
rect 510 -5 560 10
rect 590 30 640 45
rect 590 10 605 30
rect 625 10 640 30
rect 590 -5 640 10
rect 655 30 705 45
rect 655 10 670 30
rect 690 10 705 30
rect 655 -5 705 10
rect 720 30 770 45
rect 720 10 735 30
rect 755 10 770 30
rect 720 -5 770 10
rect 785 30 835 45
rect 785 10 800 30
rect 820 10 835 30
rect 785 -5 835 10
rect 850 30 900 45
rect 850 10 865 30
rect 885 10 900 30
rect 850 -5 900 10
rect 930 30 980 45
rect 930 10 945 30
rect 965 10 980 30
rect 930 -5 980 10
rect 995 30 1045 45
rect 995 10 1010 30
rect 1030 10 1045 30
rect 995 -5 1045 10
rect 1060 30 1110 45
rect 1060 10 1075 30
rect 1095 10 1110 30
rect 1060 -5 1110 10
rect 1125 30 1175 45
rect 1125 10 1140 30
rect 1160 10 1175 30
rect 1125 -5 1175 10
rect 1190 30 1240 45
rect 1190 10 1205 30
rect 1225 10 1240 30
rect 1190 -5 1240 10
<< ndiffc >>
rect -885 365 -865 585
rect -785 365 -765 585
rect -685 365 -665 585
rect -585 365 -565 585
rect -485 365 -465 585
rect -385 365 -365 585
rect -285 365 -265 585
rect -185 365 -165 585
rect -85 365 -65 585
rect -485 15 -465 235
rect -385 15 -365 235
rect -285 15 -265 235
rect -185 15 -165 235
rect -85 15 -65 235
rect 265 205 285 225
rect 330 205 350 225
rect 395 205 415 225
rect 460 205 480 225
rect 525 205 545 225
rect 590 205 610 225
rect 655 205 675 225
rect 720 205 740 225
rect 785 205 805 225
rect 865 205 885 225
rect 930 205 950 225
rect 995 205 1015 225
rect 1060 205 1080 225
rect 1125 205 1145 225
rect 1190 205 1210 225
rect 1255 205 1275 225
rect 1320 205 1340 225
rect 1385 205 1405 225
rect 1465 205 1485 225
rect 1530 205 1550 225
rect 1595 205 1615 225
rect 1660 205 1680 225
rect 1725 205 1745 225
rect 1790 205 1810 225
rect 1855 205 1875 225
rect 1920 205 1940 225
rect 1985 205 2005 225
rect 265 10 285 30
rect 330 10 350 30
rect 395 10 415 30
rect 460 10 480 30
rect 525 10 545 30
rect 605 10 625 30
rect 670 10 690 30
rect 735 10 755 30
rect 800 10 820 30
rect 865 10 885 30
rect 945 10 965 30
rect 1010 10 1030 30
rect 1075 10 1095 30
rect 1140 10 1160 30
rect 1205 10 1225 30
<< poly >>
rect -850 600 -800 615
rect -750 600 -700 615
rect -650 600 -600 615
rect -550 600 -500 615
rect -450 600 -400 615
rect -350 600 -300 615
rect -250 600 -200 615
rect -150 600 -100 615
rect -850 335 -800 350
rect -750 335 -700 350
rect -650 335 -600 350
rect -550 335 -500 350
rect -450 335 -400 350
rect -350 335 -300 350
rect -250 335 -200 350
rect -150 335 -100 350
rect -450 250 -400 265
rect -350 250 -300 265
rect -250 250 -200 265
rect -150 250 -100 265
rect 300 240 315 255
rect 365 240 380 255
rect 430 240 445 255
rect 495 240 510 255
rect 560 240 575 255
rect 625 240 640 255
rect 690 240 705 255
rect 755 240 770 255
rect 900 240 915 255
rect 965 240 980 255
rect 1030 240 1045 255
rect 1095 240 1110 255
rect 1160 240 1175 255
rect 1225 240 1240 255
rect 1290 240 1305 255
rect 1355 240 1370 255
rect 1500 240 1515 255
rect 1565 240 1580 255
rect 1630 240 1645 255
rect 1695 240 1710 255
rect 1760 240 1775 255
rect 1825 240 1840 255
rect 1890 240 1905 255
rect 1955 240 1970 255
rect 300 175 315 190
rect 365 175 380 190
rect 430 175 445 190
rect 495 175 510 190
rect 560 175 575 190
rect 625 175 640 190
rect 690 175 705 190
rect 755 175 770 190
rect 300 165 770 175
rect 300 160 330 165
rect 320 145 330 160
rect 350 160 460 165
rect 350 145 360 160
rect 320 135 360 145
rect 450 145 460 160
rect 480 160 590 165
rect 480 145 490 160
rect 450 135 490 145
rect 580 145 590 160
rect 610 160 720 165
rect 610 145 620 160
rect 580 135 620 145
rect 710 145 720 160
rect 740 160 770 165
rect 900 175 915 190
rect 965 175 980 190
rect 1030 175 1045 190
rect 1095 175 1110 190
rect 1160 175 1175 190
rect 1225 175 1240 190
rect 1290 175 1305 190
rect 1355 175 1370 190
rect 900 165 1370 175
rect 1500 180 1515 190
rect 1565 180 1580 190
rect 1630 180 1645 190
rect 1695 180 1710 190
rect 1760 180 1775 190
rect 1825 180 1840 190
rect 1890 180 1905 190
rect 1955 180 1970 190
rect 1500 165 1970 180
rect 900 160 930 165
rect 740 145 750 160
rect 710 135 750 145
rect 920 145 930 160
rect 950 160 1060 165
rect 950 145 960 160
rect 920 135 960 145
rect 1050 145 1060 160
rect 1080 160 1190 165
rect 1080 145 1090 160
rect 1050 135 1090 145
rect 1180 145 1190 160
rect 1210 160 1320 165
rect 1210 145 1220 160
rect 1180 135 1220 145
rect 1310 145 1320 160
rect 1340 160 1370 165
rect 1340 145 1350 160
rect 1310 135 1350 145
rect 320 90 360 100
rect 320 75 330 90
rect 300 70 330 75
rect 350 75 360 90
rect 450 90 490 100
rect 450 75 460 90
rect 350 70 460 75
rect 480 75 490 90
rect 660 90 700 100
rect 660 75 670 90
rect 480 70 510 75
rect 300 60 510 70
rect 300 45 315 60
rect 365 45 380 60
rect 430 45 445 60
rect 495 45 510 60
rect 640 70 670 75
rect 690 75 700 90
rect 790 90 830 100
rect 790 75 800 90
rect 690 70 800 75
rect 820 75 830 90
rect 820 70 850 75
rect 640 60 850 70
rect 640 45 655 60
rect 705 45 720 60
rect 770 45 785 60
rect 835 45 850 60
rect 980 55 1190 70
rect 980 45 995 55
rect 1045 45 1060 55
rect 1110 45 1125 55
rect 1175 45 1190 55
rect -450 -15 -400 0
rect -350 -15 -300 0
rect -250 -15 -200 0
rect -150 -15 -100 0
rect 300 -20 315 -5
rect 365 -20 380 -5
rect 430 -20 445 -5
rect 495 -20 510 -5
rect 640 -20 655 -5
rect 705 -20 720 -5
rect 770 -20 785 -5
rect 835 -20 850 -5
rect 980 -20 995 -5
rect 1045 -20 1060 -5
rect 1110 -20 1125 -5
rect 1175 -20 1190 -5
<< polycont >>
rect 330 145 350 165
rect 460 145 480 165
rect 590 145 610 165
rect 720 145 740 165
rect 930 145 950 165
rect 1060 145 1080 165
rect 1190 145 1210 165
rect 1320 145 1340 165
rect 330 70 350 90
rect 460 70 480 90
rect 670 70 690 90
rect 800 70 820 90
<< locali >>
rect -895 585 -855 595
rect -895 365 -885 585
rect -865 365 -855 585
rect -895 355 -855 365
rect -795 585 -755 595
rect -795 365 -785 585
rect -765 365 -755 585
rect -795 355 -755 365
rect -695 585 -655 595
rect -695 365 -685 585
rect -665 365 -655 585
rect -695 355 -655 365
rect -595 585 -555 595
rect -595 365 -585 585
rect -565 365 -555 585
rect -595 355 -555 365
rect -495 585 -455 595
rect -495 365 -485 585
rect -465 365 -455 585
rect -495 355 -455 365
rect -395 585 -355 595
rect -395 365 -385 585
rect -365 365 -355 585
rect -395 355 -355 365
rect -295 585 -255 595
rect -295 365 -285 585
rect -265 365 -255 585
rect -295 355 -255 365
rect -195 585 -155 595
rect -195 365 -185 585
rect -165 365 -155 585
rect -195 355 -155 365
rect -95 585 -55 595
rect -95 365 -85 585
rect -65 365 -55 585
rect -95 355 -55 365
rect -495 235 -455 245
rect -495 15 -485 235
rect -465 15 -455 235
rect -495 5 -455 15
rect -395 235 -355 245
rect -395 15 -385 235
rect -365 15 -355 235
rect -395 5 -355 15
rect -295 235 -255 245
rect -295 15 -285 235
rect -265 15 -255 235
rect -295 5 -255 15
rect -195 235 -155 245
rect -195 15 -185 235
rect -165 15 -155 235
rect -195 5 -155 15
rect -95 235 -55 245
rect 265 235 285 275
rect 395 235 415 275
rect 525 235 545 275
rect 655 235 675 275
rect 785 235 805 270
rect 865 235 885 275
rect 995 235 1015 275
rect 1125 235 1145 275
rect 1255 235 1275 275
rect 1385 235 1405 270
rect 1465 235 1485 275
rect 1595 235 1615 275
rect 1725 235 1745 275
rect 1855 235 1875 275
rect 1985 235 2005 270
rect -95 15 -85 235
rect -65 15 -55 235
rect 255 225 295 235
rect 255 205 265 225
rect 285 205 295 225
rect 255 195 295 205
rect 320 225 360 235
rect 320 205 330 225
rect 350 205 360 225
rect 320 195 360 205
rect 385 225 425 235
rect 385 205 395 225
rect 415 205 425 225
rect 385 195 425 205
rect 450 225 490 235
rect 450 205 460 225
rect 480 205 490 225
rect 450 195 490 205
rect 515 225 555 235
rect 515 205 525 225
rect 545 205 555 225
rect 515 195 555 205
rect 580 225 620 235
rect 580 205 590 225
rect 610 205 620 225
rect 580 195 620 205
rect 645 225 685 235
rect 645 205 655 225
rect 675 205 685 225
rect 645 195 685 205
rect 710 225 750 235
rect 710 205 720 225
rect 740 205 750 225
rect 710 195 750 205
rect 775 225 815 235
rect 775 205 785 225
rect 805 205 815 225
rect 775 195 815 205
rect 855 225 895 235
rect 855 205 865 225
rect 885 205 895 225
rect 855 195 895 205
rect 920 225 960 235
rect 920 205 930 225
rect 950 205 960 225
rect 920 195 960 205
rect 985 225 1025 235
rect 985 205 995 225
rect 1015 205 1025 225
rect 985 195 1025 205
rect 1050 225 1090 235
rect 1050 205 1060 225
rect 1080 205 1090 225
rect 1050 195 1090 205
rect 1115 225 1155 235
rect 1115 205 1125 225
rect 1145 205 1155 225
rect 1115 195 1155 205
rect 1180 225 1220 235
rect 1180 205 1190 225
rect 1210 205 1220 225
rect 1180 195 1220 205
rect 1245 225 1285 235
rect 1245 205 1255 225
rect 1275 205 1285 225
rect 1245 195 1285 205
rect 1310 225 1350 235
rect 1310 205 1320 225
rect 1340 205 1350 225
rect 1310 195 1350 205
rect 1375 225 1415 235
rect 1375 205 1385 225
rect 1405 205 1415 225
rect 1375 195 1415 205
rect 1455 225 1495 235
rect 1455 205 1465 225
rect 1485 205 1495 225
rect 1455 195 1495 205
rect 1520 225 1560 235
rect 1520 205 1530 225
rect 1550 205 1560 225
rect 1520 195 1560 205
rect 1585 225 1625 235
rect 1585 205 1595 225
rect 1615 205 1625 225
rect 1585 195 1625 205
rect 1650 225 1690 235
rect 1650 205 1660 225
rect 1680 205 1690 225
rect 1650 195 1690 205
rect 1715 225 1755 235
rect 1715 205 1725 225
rect 1745 205 1755 225
rect 1715 195 1755 205
rect 1780 225 1820 235
rect 1780 205 1790 225
rect 1810 205 1820 225
rect 1780 195 1820 205
rect 1845 225 1885 235
rect 1845 205 1855 225
rect 1875 205 1885 225
rect 1845 195 1885 205
rect 1910 225 1950 235
rect 1910 205 1920 225
rect 1940 205 1950 225
rect 1910 195 1950 205
rect 1975 225 2015 235
rect 1975 205 1985 225
rect 2005 205 2015 225
rect 1975 195 2015 205
rect 330 175 350 195
rect 460 175 480 195
rect 590 175 610 195
rect 720 175 740 195
rect 930 175 950 195
rect 1060 175 1080 195
rect 1190 175 1210 195
rect 1320 175 1340 195
rect 320 165 360 175
rect 320 145 330 165
rect 350 145 360 165
rect 320 135 360 145
rect 450 165 490 175
rect 450 145 460 165
rect 480 145 490 165
rect 450 135 490 145
rect 580 165 620 175
rect 580 145 590 165
rect 610 145 620 165
rect 580 135 620 145
rect 710 165 750 175
rect 710 145 720 165
rect 740 145 750 165
rect 710 135 750 145
rect 920 165 960 175
rect 920 145 930 165
rect 950 145 960 165
rect 920 135 960 145
rect 1050 165 1090 175
rect 1050 145 1060 165
rect 1080 145 1090 165
rect 1050 135 1090 145
rect 1180 165 1220 175
rect 1180 145 1190 165
rect 1210 145 1220 165
rect 1180 135 1220 145
rect 1310 165 1350 175
rect 1310 145 1320 165
rect 1340 145 1350 165
rect 1310 135 1350 145
rect 320 90 360 100
rect 320 70 330 90
rect 350 70 360 90
rect 320 60 360 70
rect 450 90 490 100
rect 450 70 460 90
rect 480 70 490 90
rect 450 60 490 70
rect 660 90 700 100
rect 660 70 670 90
rect 690 70 700 90
rect 660 60 700 70
rect 790 90 830 100
rect 790 70 800 90
rect 820 70 830 90
rect 790 60 830 70
rect 330 40 350 60
rect 460 40 480 60
rect 670 40 690 60
rect 800 40 820 60
rect -95 5 -55 15
rect 255 30 295 40
rect 255 10 265 30
rect 285 10 295 30
rect 255 0 295 10
rect 320 30 360 40
rect 320 10 330 30
rect 350 10 360 30
rect 320 0 360 10
rect 385 30 425 40
rect 385 10 395 30
rect 415 10 425 30
rect 385 0 425 10
rect 450 30 490 40
rect 450 10 460 30
rect 480 10 490 30
rect 450 0 490 10
rect 515 30 555 40
rect 515 10 525 30
rect 545 10 555 30
rect 515 0 555 10
rect 595 30 635 40
rect 595 10 605 30
rect 625 10 635 30
rect 595 0 635 10
rect 660 30 700 40
rect 660 10 670 30
rect 690 10 700 30
rect 660 0 700 10
rect 725 30 765 40
rect 725 10 735 30
rect 755 10 765 30
rect 725 0 765 10
rect 790 30 830 40
rect 790 10 800 30
rect 820 10 830 30
rect 790 0 830 10
rect 855 30 895 40
rect 855 10 865 30
rect 885 10 895 30
rect 855 0 895 10
rect 935 30 975 40
rect 935 10 945 30
rect 965 10 975 30
rect 935 0 975 10
rect 1000 30 1040 40
rect 1000 10 1010 30
rect 1030 10 1040 30
rect 1000 0 1040 10
rect 1065 30 1105 40
rect 1065 10 1075 30
rect 1095 10 1105 30
rect 1065 0 1105 10
rect 1130 30 1170 40
rect 1130 10 1140 30
rect 1160 10 1170 30
rect 1130 0 1170 10
rect 1195 30 1235 40
rect 1195 10 1205 30
rect 1225 10 1235 30
rect 1195 0 1235 10
rect 265 -35 285 0
rect 395 -40 415 0
rect 525 -40 545 0
rect 605 -35 625 0
rect 735 -40 755 0
rect 865 -40 885 0
rect 945 -35 965 0
rect 1075 -40 1095 0
rect 1205 -40 1225 0
<< end >>
