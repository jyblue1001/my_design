** sch_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/phase_frequency_detector_5.sch
**.subckt phase_frequency_detector_5 F_REF F_VCO VDDA QA QB GNDA
*.ipin F_REF
*.opin QA
*.ipin F_VCO
*.opin QB
*.ipin VDDA
*.ipin GNDA
x1 VDDA GNDA QA F_REF QA_b nor_pfd
x2 VDDA GNDA QB F_VCO QB_b nor_pfd
x3 VDDA GNDA QA_b E QA nor_pfd
x4 VDDA GNDA QB_b F QB nor_pfd
x5 VDDA GNDA E_b QA_b E nor_pfd
x6 VDDA GNDA F_b QB_b F nor_pfd
x7 VDDA GNDA E Reset E_b nor_pfd
x12 VDDA GNDA F Reset F_b nor_pfd
x8 VDDA GNDA QB QA before_Reset nand_pfd
x9 VDDA GNDA before_Reset net1 inv_pfd
x10 VDDA GNDA net1 net2 inv_pfd
x11 VDDA GNDA net2 net3 inv_pfd
x13 VDDA GNDA net3 net4 inv_pfd
x14 VDDA GNDA net4 Reset inv_pfd
**.ends

* expanding   symbol:  /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/nor_pfd.sym # of pins=5
** sym_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/nor_pfd.sym
** sch_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/nor_pfd.sch
.subckt nor_pfd VDDA GNDA A B Y
*.ipin A
*.opin Y
*.ipin VDDA
*.ipin GNDA
*.ipin B
XM4 net1 B VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 GNDA B Y GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 GNDA A Y GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A net1 VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/nand_pfd.sym # of pins=5
** sym_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/nand_pfd.sym
** sch_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/nand_pfd.sch
.subckt nand_pfd VDDA GNDA A B Y
*.ipin A
*.opin Y
*.ipin VDDA
*.ipin GNDA
*.ipin B
XM4 Y B VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 B Y GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 GNDA A net1 GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/inv_pfd.sym # of pins=4
** sym_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/inv_pfd.sym
** sch_path: /foss/designs/my_design/projects/pll/pfd/xschem_ngspice/inv_pfd.sch
.subckt inv_pfd VDDA GNDA A Y
*.ipin A
*.opin Y
*.ipin VDDA
*.ipin GNDA
XM2 Y A VDDA VDDA sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 GNDA A Y GNDA sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
