magic
tech sky130A
magscale 1 2
timestamp 1746289854
<< pwell >>
rect 1350 1187 2690 1340
rect 1350 153 1503 1187
rect 2537 153 2690 1187
rect 1350 0 2690 153
rect 2700 1187 4040 1340
rect 2700 153 2853 1187
rect 3887 153 4040 1187
rect 2700 0 4040 153
rect 4050 1187 5390 1340
rect 4050 153 4203 1187
rect 5237 153 5390 1187
rect 4050 0 5390 153
rect 5400 1187 6740 1340
rect 5400 153 5553 1187
rect 6587 153 6740 1187
rect 5400 0 6740 153
rect 6750 1187 8090 1340
rect 6750 153 6903 1187
rect 7937 153 8090 1187
rect 6750 0 8090 153
rect 8100 1187 9440 1340
rect 8100 153 8253 1187
rect 9287 153 9440 1187
rect 8100 0 9440 153
<< nbase >>
rect 1503 153 2537 1187
rect 2853 153 3887 1187
rect 4203 153 5237 1187
rect 5553 153 6587 1187
rect 6903 153 7937 1187
rect 8253 153 9287 1187
<< nmos >>
rect -1610 3960 -1580 4360
rect -1310 3960 -1280 4360
rect 1970 3960 2090 4760
rect 2190 3960 2310 4760
rect 2410 3960 2530 4760
rect 2630 3960 2750 4760
rect 2850 3960 2970 4760
rect 3070 3960 3190 4760
rect 3290 3960 3410 4760
rect 3510 3960 3630 4760
rect 3730 3960 3850 4760
rect 3950 3960 4070 4760
rect 4170 3960 4290 4760
rect 4390 3960 4510 4760
rect 5390 4460 5510 4860
rect 5610 4460 5730 4860
rect 5830 4460 5950 4860
rect 6050 4460 6170 4860
rect 6270 4460 6390 4860
rect 6490 4460 6610 4860
rect 6710 4460 6830 4860
rect 6930 4460 7050 4860
rect 7150 4460 7270 4860
rect 7370 4460 7490 4860
rect 7590 4460 7710 4860
rect 7810 4460 7930 4860
rect 5830 3710 5950 3910
rect 6050 3710 6170 3910
rect 6270 3710 6390 3910
rect 6490 3710 6610 3910
rect 6710 3710 6830 3910
rect 6930 3710 7050 3910
rect 7150 3710 7270 3910
rect 7370 3710 7490 3910
rect -2710 3460 -710 3660
rect 5810 2560 6610 3360
rect 6710 2560 7510 3360
<< ndiff >>
rect 5290 4830 5390 4860
rect 5290 4790 5320 4830
rect 5360 4790 5390 4830
rect 1870 4730 1970 4760
rect -1710 4330 -1610 4360
rect -1710 3990 -1680 4330
rect -1640 3990 -1610 4330
rect -1710 3960 -1610 3990
rect -1580 4330 -1480 4360
rect -1580 3990 -1550 4330
rect -1510 3990 -1480 4330
rect -1580 3960 -1480 3990
rect -1410 4330 -1310 4360
rect -1410 3990 -1380 4330
rect -1340 3990 -1310 4330
rect -1410 3960 -1310 3990
rect -1280 4330 -1180 4360
rect -1280 3990 -1250 4330
rect -1210 3990 -1180 4330
rect -1280 3960 -1180 3990
rect 1870 3990 1900 4730
rect 1940 3990 1970 4730
rect 1870 3960 1970 3990
rect 2090 4730 2190 4760
rect 2090 3990 2120 4730
rect 2160 3990 2190 4730
rect 2090 3960 2190 3990
rect 2310 4730 2410 4760
rect 2310 3990 2340 4730
rect 2380 3990 2410 4730
rect 2310 3960 2410 3990
rect 2530 4730 2630 4760
rect 2530 3990 2560 4730
rect 2600 3990 2630 4730
rect 2530 3960 2630 3990
rect 2750 4730 2850 4760
rect 2750 3990 2780 4730
rect 2820 3990 2850 4730
rect 2750 3960 2850 3990
rect 2970 4730 3070 4760
rect 2970 3990 3000 4730
rect 3040 3990 3070 4730
rect 2970 3960 3070 3990
rect 3190 4730 3290 4760
rect 3190 3990 3220 4730
rect 3260 3990 3290 4730
rect 3190 3960 3290 3990
rect 3410 4730 3510 4760
rect 3410 3990 3440 4730
rect 3480 3990 3510 4730
rect 3410 3960 3510 3990
rect 3630 4730 3730 4760
rect 3630 3990 3660 4730
rect 3700 3990 3730 4730
rect 3630 3960 3730 3990
rect 3850 4730 3950 4760
rect 3850 3990 3880 4730
rect 3920 3990 3950 4730
rect 3850 3960 3950 3990
rect 4070 4730 4170 4760
rect 4070 3990 4100 4730
rect 4140 3990 4170 4730
rect 4070 3960 4170 3990
rect 4290 4730 4390 4760
rect 4290 3990 4320 4730
rect 4360 3990 4390 4730
rect 4290 3960 4390 3990
rect 4510 4730 4610 4760
rect 4510 3990 4540 4730
rect 4580 3990 4610 4730
rect 5290 4730 5390 4790
rect 5290 4690 5320 4730
rect 5360 4690 5390 4730
rect 5290 4630 5390 4690
rect 5290 4590 5320 4630
rect 5360 4590 5390 4630
rect 5290 4530 5390 4590
rect 5290 4490 5320 4530
rect 5360 4490 5390 4530
rect 5290 4460 5390 4490
rect 5510 4830 5610 4860
rect 5510 4790 5540 4830
rect 5580 4790 5610 4830
rect 5510 4730 5610 4790
rect 5510 4690 5540 4730
rect 5580 4690 5610 4730
rect 5510 4630 5610 4690
rect 5510 4590 5540 4630
rect 5580 4590 5610 4630
rect 5510 4530 5610 4590
rect 5510 4490 5540 4530
rect 5580 4490 5610 4530
rect 5510 4460 5610 4490
rect 5730 4830 5830 4860
rect 5730 4790 5760 4830
rect 5800 4790 5830 4830
rect 5730 4730 5830 4790
rect 5730 4690 5760 4730
rect 5800 4690 5830 4730
rect 5730 4630 5830 4690
rect 5730 4590 5760 4630
rect 5800 4590 5830 4630
rect 5730 4530 5830 4590
rect 5730 4490 5760 4530
rect 5800 4490 5830 4530
rect 5730 4460 5830 4490
rect 5950 4830 6050 4860
rect 5950 4790 5980 4830
rect 6020 4790 6050 4830
rect 5950 4730 6050 4790
rect 5950 4690 5980 4730
rect 6020 4690 6050 4730
rect 5950 4630 6050 4690
rect 5950 4590 5980 4630
rect 6020 4590 6050 4630
rect 5950 4530 6050 4590
rect 5950 4490 5980 4530
rect 6020 4490 6050 4530
rect 5950 4460 6050 4490
rect 6170 4830 6270 4860
rect 6170 4790 6200 4830
rect 6240 4790 6270 4830
rect 6170 4730 6270 4790
rect 6170 4690 6200 4730
rect 6240 4690 6270 4730
rect 6170 4630 6270 4690
rect 6170 4590 6200 4630
rect 6240 4590 6270 4630
rect 6170 4530 6270 4590
rect 6170 4490 6200 4530
rect 6240 4490 6270 4530
rect 6170 4460 6270 4490
rect 6390 4830 6490 4860
rect 6390 4790 6420 4830
rect 6460 4790 6490 4830
rect 6390 4730 6490 4790
rect 6390 4690 6420 4730
rect 6460 4690 6490 4730
rect 6390 4630 6490 4690
rect 6390 4590 6420 4630
rect 6460 4590 6490 4630
rect 6390 4530 6490 4590
rect 6390 4490 6420 4530
rect 6460 4490 6490 4530
rect 6390 4460 6490 4490
rect 6610 4830 6710 4860
rect 6610 4790 6640 4830
rect 6680 4790 6710 4830
rect 6610 4730 6710 4790
rect 6610 4690 6640 4730
rect 6680 4690 6710 4730
rect 6610 4630 6710 4690
rect 6610 4590 6640 4630
rect 6680 4590 6710 4630
rect 6610 4530 6710 4590
rect 6610 4490 6640 4530
rect 6680 4490 6710 4530
rect 6610 4460 6710 4490
rect 6830 4830 6930 4860
rect 6830 4790 6860 4830
rect 6900 4790 6930 4830
rect 6830 4730 6930 4790
rect 6830 4690 6860 4730
rect 6900 4690 6930 4730
rect 6830 4630 6930 4690
rect 6830 4590 6860 4630
rect 6900 4590 6930 4630
rect 6830 4530 6930 4590
rect 6830 4490 6860 4530
rect 6900 4490 6930 4530
rect 6830 4460 6930 4490
rect 7050 4830 7150 4860
rect 7050 4790 7080 4830
rect 7120 4790 7150 4830
rect 7050 4730 7150 4790
rect 7050 4690 7080 4730
rect 7120 4690 7150 4730
rect 7050 4630 7150 4690
rect 7050 4590 7080 4630
rect 7120 4590 7150 4630
rect 7050 4530 7150 4590
rect 7050 4490 7080 4530
rect 7120 4490 7150 4530
rect 7050 4460 7150 4490
rect 7270 4830 7370 4860
rect 7270 4790 7300 4830
rect 7340 4790 7370 4830
rect 7270 4730 7370 4790
rect 7270 4690 7300 4730
rect 7340 4690 7370 4730
rect 7270 4630 7370 4690
rect 7270 4590 7300 4630
rect 7340 4590 7370 4630
rect 7270 4530 7370 4590
rect 7270 4490 7300 4530
rect 7340 4490 7370 4530
rect 7270 4460 7370 4490
rect 7490 4830 7590 4860
rect 7490 4790 7520 4830
rect 7560 4790 7590 4830
rect 7490 4730 7590 4790
rect 7490 4690 7520 4730
rect 7560 4690 7590 4730
rect 7490 4630 7590 4690
rect 7490 4590 7520 4630
rect 7560 4590 7590 4630
rect 7490 4530 7590 4590
rect 7490 4490 7520 4530
rect 7560 4490 7590 4530
rect 7490 4460 7590 4490
rect 7710 4830 7810 4860
rect 7710 4790 7740 4830
rect 7780 4790 7810 4830
rect 7710 4730 7810 4790
rect 7710 4690 7740 4730
rect 7780 4690 7810 4730
rect 7710 4630 7810 4690
rect 7710 4590 7740 4630
rect 7780 4590 7810 4630
rect 7710 4530 7810 4590
rect 7710 4490 7740 4530
rect 7780 4490 7810 4530
rect 7710 4460 7810 4490
rect 7930 4830 8030 4860
rect 7930 4790 7960 4830
rect 8000 4790 8030 4830
rect 7930 4730 8030 4790
rect 7930 4690 7960 4730
rect 8000 4690 8030 4730
rect 7930 4630 8030 4690
rect 7930 4590 7960 4630
rect 8000 4590 8030 4630
rect 7930 4530 8030 4590
rect 7930 4490 7960 4530
rect 8000 4490 8030 4530
rect 7930 4460 8030 4490
rect 4510 3960 4610 3990
rect 5730 3880 5830 3910
rect 5730 3840 5760 3880
rect 5800 3840 5830 3880
rect 5730 3780 5830 3840
rect 5730 3740 5760 3780
rect 5800 3740 5830 3780
rect 5730 3710 5830 3740
rect 5950 3880 6050 3910
rect 5950 3840 5980 3880
rect 6020 3840 6050 3880
rect 5950 3780 6050 3840
rect 5950 3740 5980 3780
rect 6020 3740 6050 3780
rect 5950 3710 6050 3740
rect 6170 3880 6270 3910
rect 6170 3840 6200 3880
rect 6240 3840 6270 3880
rect 6170 3780 6270 3840
rect 6170 3740 6200 3780
rect 6240 3740 6270 3780
rect 6170 3710 6270 3740
rect 6390 3880 6490 3910
rect 6390 3840 6420 3880
rect 6460 3840 6490 3880
rect 6390 3780 6490 3840
rect 6390 3740 6420 3780
rect 6460 3740 6490 3780
rect 6390 3710 6490 3740
rect 6610 3880 6710 3910
rect 6610 3840 6640 3880
rect 6680 3840 6710 3880
rect 6610 3780 6710 3840
rect 6610 3740 6640 3780
rect 6680 3740 6710 3780
rect 6610 3710 6710 3740
rect 6830 3880 6930 3910
rect 6830 3840 6860 3880
rect 6900 3840 6930 3880
rect 6830 3780 6930 3840
rect 6830 3740 6860 3780
rect 6900 3740 6930 3780
rect 6830 3710 6930 3740
rect 7050 3880 7150 3910
rect 7050 3840 7080 3880
rect 7120 3840 7150 3880
rect 7050 3780 7150 3840
rect 7050 3740 7080 3780
rect 7120 3740 7150 3780
rect 7050 3710 7150 3740
rect 7270 3880 7370 3910
rect 7270 3840 7300 3880
rect 7340 3840 7370 3880
rect 7270 3780 7370 3840
rect 7270 3740 7300 3780
rect 7340 3740 7370 3780
rect 7270 3710 7370 3740
rect 7490 3880 7590 3910
rect 7490 3840 7520 3880
rect 7560 3840 7590 3880
rect 7490 3780 7590 3840
rect 7490 3740 7520 3780
rect 7560 3740 7590 3780
rect 7490 3710 7590 3740
rect -2810 3630 -2710 3660
rect -2810 3490 -2780 3630
rect -2740 3490 -2710 3630
rect -2810 3460 -2710 3490
rect -710 3630 -610 3660
rect -710 3490 -680 3630
rect -640 3490 -610 3630
rect -710 3460 -610 3490
rect 5710 3330 5810 3360
rect 5710 3290 5740 3330
rect 5780 3290 5810 3330
rect 5710 3230 5810 3290
rect 5710 3190 5740 3230
rect 5780 3190 5810 3230
rect 5710 3130 5810 3190
rect 5710 3090 5740 3130
rect 5780 3090 5810 3130
rect 5710 3030 5810 3090
rect 5710 2990 5740 3030
rect 5780 2990 5810 3030
rect 5710 2930 5810 2990
rect 5710 2890 5740 2930
rect 5780 2890 5810 2930
rect 5710 2830 5810 2890
rect 5710 2790 5740 2830
rect 5780 2790 5810 2830
rect 5710 2730 5810 2790
rect 5710 2690 5740 2730
rect 5780 2690 5810 2730
rect 5710 2630 5810 2690
rect 5710 2590 5740 2630
rect 5780 2590 5810 2630
rect 5710 2560 5810 2590
rect 6610 3330 6710 3360
rect 6610 3290 6640 3330
rect 6680 3290 6710 3330
rect 6610 3230 6710 3290
rect 6610 3190 6640 3230
rect 6680 3190 6710 3230
rect 6610 3130 6710 3190
rect 6610 3090 6640 3130
rect 6680 3090 6710 3130
rect 6610 3030 6710 3090
rect 6610 2990 6640 3030
rect 6680 2990 6710 3030
rect 6610 2930 6710 2990
rect 6610 2890 6640 2930
rect 6680 2890 6710 2930
rect 6610 2830 6710 2890
rect 6610 2790 6640 2830
rect 6680 2790 6710 2830
rect 6610 2730 6710 2790
rect 6610 2690 6640 2730
rect 6680 2690 6710 2730
rect 6610 2630 6710 2690
rect 6610 2590 6640 2630
rect 6680 2590 6710 2630
rect 6610 2560 6710 2590
rect 7510 3330 7610 3360
rect 7510 3290 7540 3330
rect 7580 3290 7610 3330
rect 7510 3230 7610 3290
rect 7510 3190 7540 3230
rect 7580 3190 7610 3230
rect 7510 3130 7610 3190
rect 7510 3090 7540 3130
rect 7580 3090 7610 3130
rect 7510 3030 7610 3090
rect 7510 2990 7540 3030
rect 7580 2990 7610 3030
rect 7510 2930 7610 2990
rect 7510 2890 7540 2930
rect 7580 2890 7610 2930
rect 7510 2830 7610 2890
rect 7510 2790 7540 2830
rect 7580 2790 7610 2830
rect 7510 2730 7610 2790
rect 7510 2690 7540 2730
rect 7580 2690 7610 2730
rect 7510 2630 7610 2690
rect 7510 2590 7540 2630
rect 7580 2590 7610 2630
rect 7510 2560 7610 2590
<< pdiff >>
rect 1680 958 2360 1010
rect 1680 924 1734 958
rect 1768 924 1824 958
rect 1858 924 1914 958
rect 1948 924 2004 958
rect 2038 924 2094 958
rect 2128 924 2184 958
rect 2218 924 2274 958
rect 2308 924 2360 958
rect 1680 868 2360 924
rect 1680 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2360 868
rect 1680 778 2360 834
rect 1680 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2360 778
rect 1680 688 2360 744
rect 1680 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2360 688
rect 1680 598 2360 654
rect 1680 564 1734 598
rect 1768 564 1824 598
rect 1858 564 1914 598
rect 1948 564 2004 598
rect 2038 564 2094 598
rect 2128 564 2184 598
rect 2218 564 2274 598
rect 2308 564 2360 598
rect 1680 508 2360 564
rect 1680 474 1734 508
rect 1768 474 1824 508
rect 1858 474 1914 508
rect 1948 474 2004 508
rect 2038 474 2094 508
rect 2128 474 2184 508
rect 2218 474 2274 508
rect 2308 474 2360 508
rect 1680 418 2360 474
rect 1680 384 1734 418
rect 1768 384 1824 418
rect 1858 384 1914 418
rect 1948 384 2004 418
rect 2038 384 2094 418
rect 2128 384 2184 418
rect 2218 384 2274 418
rect 2308 384 2360 418
rect 1680 330 2360 384
rect 3030 958 3710 1010
rect 3030 924 3084 958
rect 3118 924 3174 958
rect 3208 924 3264 958
rect 3298 924 3354 958
rect 3388 924 3444 958
rect 3478 924 3534 958
rect 3568 924 3624 958
rect 3658 924 3710 958
rect 3030 868 3710 924
rect 3030 834 3084 868
rect 3118 834 3174 868
rect 3208 834 3264 868
rect 3298 834 3354 868
rect 3388 834 3444 868
rect 3478 834 3534 868
rect 3568 834 3624 868
rect 3658 834 3710 868
rect 3030 778 3710 834
rect 3030 744 3084 778
rect 3118 744 3174 778
rect 3208 744 3264 778
rect 3298 744 3354 778
rect 3388 744 3444 778
rect 3478 744 3534 778
rect 3568 744 3624 778
rect 3658 744 3710 778
rect 3030 688 3710 744
rect 3030 654 3084 688
rect 3118 654 3174 688
rect 3208 654 3264 688
rect 3298 654 3354 688
rect 3388 654 3444 688
rect 3478 654 3534 688
rect 3568 654 3624 688
rect 3658 654 3710 688
rect 3030 598 3710 654
rect 3030 564 3084 598
rect 3118 564 3174 598
rect 3208 564 3264 598
rect 3298 564 3354 598
rect 3388 564 3444 598
rect 3478 564 3534 598
rect 3568 564 3624 598
rect 3658 564 3710 598
rect 3030 508 3710 564
rect 3030 474 3084 508
rect 3118 474 3174 508
rect 3208 474 3264 508
rect 3298 474 3354 508
rect 3388 474 3444 508
rect 3478 474 3534 508
rect 3568 474 3624 508
rect 3658 474 3710 508
rect 3030 418 3710 474
rect 3030 384 3084 418
rect 3118 384 3174 418
rect 3208 384 3264 418
rect 3298 384 3354 418
rect 3388 384 3444 418
rect 3478 384 3534 418
rect 3568 384 3624 418
rect 3658 384 3710 418
rect 3030 330 3710 384
rect 4380 958 5060 1010
rect 4380 924 4434 958
rect 4468 924 4524 958
rect 4558 924 4614 958
rect 4648 924 4704 958
rect 4738 924 4794 958
rect 4828 924 4884 958
rect 4918 924 4974 958
rect 5008 924 5060 958
rect 4380 868 5060 924
rect 4380 834 4434 868
rect 4468 834 4524 868
rect 4558 834 4614 868
rect 4648 834 4704 868
rect 4738 834 4794 868
rect 4828 834 4884 868
rect 4918 834 4974 868
rect 5008 834 5060 868
rect 4380 778 5060 834
rect 4380 744 4434 778
rect 4468 744 4524 778
rect 4558 744 4614 778
rect 4648 744 4704 778
rect 4738 744 4794 778
rect 4828 744 4884 778
rect 4918 744 4974 778
rect 5008 744 5060 778
rect 4380 688 5060 744
rect 4380 654 4434 688
rect 4468 654 4524 688
rect 4558 654 4614 688
rect 4648 654 4704 688
rect 4738 654 4794 688
rect 4828 654 4884 688
rect 4918 654 4974 688
rect 5008 654 5060 688
rect 4380 598 5060 654
rect 4380 564 4434 598
rect 4468 564 4524 598
rect 4558 564 4614 598
rect 4648 564 4704 598
rect 4738 564 4794 598
rect 4828 564 4884 598
rect 4918 564 4974 598
rect 5008 564 5060 598
rect 4380 508 5060 564
rect 4380 474 4434 508
rect 4468 474 4524 508
rect 4558 474 4614 508
rect 4648 474 4704 508
rect 4738 474 4794 508
rect 4828 474 4884 508
rect 4918 474 4974 508
rect 5008 474 5060 508
rect 4380 418 5060 474
rect 4380 384 4434 418
rect 4468 384 4524 418
rect 4558 384 4614 418
rect 4648 384 4704 418
rect 4738 384 4794 418
rect 4828 384 4884 418
rect 4918 384 4974 418
rect 5008 384 5060 418
rect 4380 330 5060 384
rect 5730 958 6410 1010
rect 5730 924 5784 958
rect 5818 924 5874 958
rect 5908 924 5964 958
rect 5998 924 6054 958
rect 6088 924 6144 958
rect 6178 924 6234 958
rect 6268 924 6324 958
rect 6358 924 6410 958
rect 5730 868 6410 924
rect 5730 834 5784 868
rect 5818 834 5874 868
rect 5908 834 5964 868
rect 5998 834 6054 868
rect 6088 834 6144 868
rect 6178 834 6234 868
rect 6268 834 6324 868
rect 6358 834 6410 868
rect 5730 778 6410 834
rect 5730 744 5784 778
rect 5818 744 5874 778
rect 5908 744 5964 778
rect 5998 744 6054 778
rect 6088 744 6144 778
rect 6178 744 6234 778
rect 6268 744 6324 778
rect 6358 744 6410 778
rect 5730 688 6410 744
rect 5730 654 5784 688
rect 5818 654 5874 688
rect 5908 654 5964 688
rect 5998 654 6054 688
rect 6088 654 6144 688
rect 6178 654 6234 688
rect 6268 654 6324 688
rect 6358 654 6410 688
rect 5730 598 6410 654
rect 5730 564 5784 598
rect 5818 564 5874 598
rect 5908 564 5964 598
rect 5998 564 6054 598
rect 6088 564 6144 598
rect 6178 564 6234 598
rect 6268 564 6324 598
rect 6358 564 6410 598
rect 5730 508 6410 564
rect 5730 474 5784 508
rect 5818 474 5874 508
rect 5908 474 5964 508
rect 5998 474 6054 508
rect 6088 474 6144 508
rect 6178 474 6234 508
rect 6268 474 6324 508
rect 6358 474 6410 508
rect 5730 418 6410 474
rect 5730 384 5784 418
rect 5818 384 5874 418
rect 5908 384 5964 418
rect 5998 384 6054 418
rect 6088 384 6144 418
rect 6178 384 6234 418
rect 6268 384 6324 418
rect 6358 384 6410 418
rect 5730 330 6410 384
rect 7080 958 7760 1010
rect 7080 924 7134 958
rect 7168 924 7224 958
rect 7258 924 7314 958
rect 7348 924 7404 958
rect 7438 924 7494 958
rect 7528 924 7584 958
rect 7618 924 7674 958
rect 7708 924 7760 958
rect 7080 868 7760 924
rect 7080 834 7134 868
rect 7168 834 7224 868
rect 7258 834 7314 868
rect 7348 834 7404 868
rect 7438 834 7494 868
rect 7528 834 7584 868
rect 7618 834 7674 868
rect 7708 834 7760 868
rect 7080 778 7760 834
rect 7080 744 7134 778
rect 7168 744 7224 778
rect 7258 744 7314 778
rect 7348 744 7404 778
rect 7438 744 7494 778
rect 7528 744 7584 778
rect 7618 744 7674 778
rect 7708 744 7760 778
rect 7080 688 7760 744
rect 7080 654 7134 688
rect 7168 654 7224 688
rect 7258 654 7314 688
rect 7348 654 7404 688
rect 7438 654 7494 688
rect 7528 654 7584 688
rect 7618 654 7674 688
rect 7708 654 7760 688
rect 7080 598 7760 654
rect 7080 564 7134 598
rect 7168 564 7224 598
rect 7258 564 7314 598
rect 7348 564 7404 598
rect 7438 564 7494 598
rect 7528 564 7584 598
rect 7618 564 7674 598
rect 7708 564 7760 598
rect 7080 508 7760 564
rect 7080 474 7134 508
rect 7168 474 7224 508
rect 7258 474 7314 508
rect 7348 474 7404 508
rect 7438 474 7494 508
rect 7528 474 7584 508
rect 7618 474 7674 508
rect 7708 474 7760 508
rect 7080 418 7760 474
rect 7080 384 7134 418
rect 7168 384 7224 418
rect 7258 384 7314 418
rect 7348 384 7404 418
rect 7438 384 7494 418
rect 7528 384 7584 418
rect 7618 384 7674 418
rect 7708 384 7760 418
rect 7080 330 7760 384
rect 8430 958 9110 1010
rect 8430 924 8484 958
rect 8518 924 8574 958
rect 8608 924 8664 958
rect 8698 924 8754 958
rect 8788 924 8844 958
rect 8878 924 8934 958
rect 8968 924 9024 958
rect 9058 924 9110 958
rect 8430 868 9110 924
rect 8430 834 8484 868
rect 8518 834 8574 868
rect 8608 834 8664 868
rect 8698 834 8754 868
rect 8788 834 8844 868
rect 8878 834 8934 868
rect 8968 834 9024 868
rect 9058 834 9110 868
rect 8430 778 9110 834
rect 8430 744 8484 778
rect 8518 744 8574 778
rect 8608 744 8664 778
rect 8698 744 8754 778
rect 8788 744 8844 778
rect 8878 744 8934 778
rect 8968 744 9024 778
rect 9058 744 9110 778
rect 8430 688 9110 744
rect 8430 654 8484 688
rect 8518 654 8574 688
rect 8608 654 8664 688
rect 8698 654 8754 688
rect 8788 654 8844 688
rect 8878 654 8934 688
rect 8968 654 9024 688
rect 9058 654 9110 688
rect 8430 598 9110 654
rect 8430 564 8484 598
rect 8518 564 8574 598
rect 8608 564 8664 598
rect 8698 564 8754 598
rect 8788 564 8844 598
rect 8878 564 8934 598
rect 8968 564 9024 598
rect 9058 564 9110 598
rect 8430 508 9110 564
rect 8430 474 8484 508
rect 8518 474 8574 508
rect 8608 474 8664 508
rect 8698 474 8754 508
rect 8788 474 8844 508
rect 8878 474 8934 508
rect 8968 474 9024 508
rect 9058 474 9110 508
rect 8430 418 9110 474
rect 8430 384 8484 418
rect 8518 384 8574 418
rect 8608 384 8664 418
rect 8698 384 8754 418
rect 8788 384 8844 418
rect 8878 384 8934 418
rect 8968 384 9024 418
rect 9058 384 9110 418
rect 8430 330 9110 384
<< ndiffc >>
rect 5320 4790 5360 4830
rect -1680 3990 -1640 4330
rect -1550 3990 -1510 4330
rect -1380 3990 -1340 4330
rect -1250 3990 -1210 4330
rect 1900 3990 1940 4730
rect 2120 3990 2160 4730
rect 2340 3990 2380 4730
rect 2560 3990 2600 4730
rect 2780 3990 2820 4730
rect 3000 3990 3040 4730
rect 3220 3990 3260 4730
rect 3440 3990 3480 4730
rect 3660 3990 3700 4730
rect 3880 3990 3920 4730
rect 4100 3990 4140 4730
rect 4320 3990 4360 4730
rect 4540 3990 4580 4730
rect 5320 4690 5360 4730
rect 5320 4590 5360 4630
rect 5320 4490 5360 4530
rect 5540 4790 5580 4830
rect 5540 4690 5580 4730
rect 5540 4590 5580 4630
rect 5540 4490 5580 4530
rect 5760 4790 5800 4830
rect 5760 4690 5800 4730
rect 5760 4590 5800 4630
rect 5760 4490 5800 4530
rect 5980 4790 6020 4830
rect 5980 4690 6020 4730
rect 5980 4590 6020 4630
rect 5980 4490 6020 4530
rect 6200 4790 6240 4830
rect 6200 4690 6240 4730
rect 6200 4590 6240 4630
rect 6200 4490 6240 4530
rect 6420 4790 6460 4830
rect 6420 4690 6460 4730
rect 6420 4590 6460 4630
rect 6420 4490 6460 4530
rect 6640 4790 6680 4830
rect 6640 4690 6680 4730
rect 6640 4590 6680 4630
rect 6640 4490 6680 4530
rect 6860 4790 6900 4830
rect 6860 4690 6900 4730
rect 6860 4590 6900 4630
rect 6860 4490 6900 4530
rect 7080 4790 7120 4830
rect 7080 4690 7120 4730
rect 7080 4590 7120 4630
rect 7080 4490 7120 4530
rect 7300 4790 7340 4830
rect 7300 4690 7340 4730
rect 7300 4590 7340 4630
rect 7300 4490 7340 4530
rect 7520 4790 7560 4830
rect 7520 4690 7560 4730
rect 7520 4590 7560 4630
rect 7520 4490 7560 4530
rect 7740 4790 7780 4830
rect 7740 4690 7780 4730
rect 7740 4590 7780 4630
rect 7740 4490 7780 4530
rect 7960 4790 8000 4830
rect 7960 4690 8000 4730
rect 7960 4590 8000 4630
rect 7960 4490 8000 4530
rect 5760 3840 5800 3880
rect 5760 3740 5800 3780
rect 5980 3840 6020 3880
rect 5980 3740 6020 3780
rect 6200 3840 6240 3880
rect 6200 3740 6240 3780
rect 6420 3840 6460 3880
rect 6420 3740 6460 3780
rect 6640 3840 6680 3880
rect 6640 3740 6680 3780
rect 6860 3840 6900 3880
rect 6860 3740 6900 3780
rect 7080 3840 7120 3880
rect 7080 3740 7120 3780
rect 7300 3840 7340 3880
rect 7300 3740 7340 3780
rect 7520 3840 7560 3880
rect 7520 3740 7560 3780
rect -2780 3490 -2740 3630
rect -680 3490 -640 3630
rect 5740 3290 5780 3330
rect 5740 3190 5780 3230
rect 5740 3090 5780 3130
rect 5740 2990 5780 3030
rect 5740 2890 5780 2930
rect 5740 2790 5780 2830
rect 5740 2690 5780 2730
rect 5740 2590 5780 2630
rect 6640 3290 6680 3330
rect 6640 3190 6680 3230
rect 6640 3090 6680 3130
rect 6640 2990 6680 3030
rect 6640 2890 6680 2930
rect 6640 2790 6680 2830
rect 6640 2690 6680 2730
rect 6640 2590 6680 2630
rect 7540 3290 7580 3330
rect 7540 3190 7580 3230
rect 7540 3090 7580 3130
rect 7540 2990 7580 3030
rect 7540 2890 7580 2930
rect 7540 2790 7580 2830
rect 7540 2690 7580 2730
rect 7540 2590 7580 2630
<< pdiffc >>
rect 1734 924 1768 958
rect 1824 924 1858 958
rect 1914 924 1948 958
rect 2004 924 2038 958
rect 2094 924 2128 958
rect 2184 924 2218 958
rect 2274 924 2308 958
rect 1734 834 1768 868
rect 1824 834 1858 868
rect 1914 834 1948 868
rect 2004 834 2038 868
rect 2094 834 2128 868
rect 2184 834 2218 868
rect 2274 834 2308 868
rect 1734 744 1768 778
rect 1824 744 1858 778
rect 1914 744 1948 778
rect 2004 744 2038 778
rect 2094 744 2128 778
rect 2184 744 2218 778
rect 2274 744 2308 778
rect 1734 654 1768 688
rect 1824 654 1858 688
rect 1914 654 1948 688
rect 2004 654 2038 688
rect 2094 654 2128 688
rect 2184 654 2218 688
rect 2274 654 2308 688
rect 1734 564 1768 598
rect 1824 564 1858 598
rect 1914 564 1948 598
rect 2004 564 2038 598
rect 2094 564 2128 598
rect 2184 564 2218 598
rect 2274 564 2308 598
rect 1734 474 1768 508
rect 1824 474 1858 508
rect 1914 474 1948 508
rect 2004 474 2038 508
rect 2094 474 2128 508
rect 2184 474 2218 508
rect 2274 474 2308 508
rect 1734 384 1768 418
rect 1824 384 1858 418
rect 1914 384 1948 418
rect 2004 384 2038 418
rect 2094 384 2128 418
rect 2184 384 2218 418
rect 2274 384 2308 418
rect 3084 924 3118 958
rect 3174 924 3208 958
rect 3264 924 3298 958
rect 3354 924 3388 958
rect 3444 924 3478 958
rect 3534 924 3568 958
rect 3624 924 3658 958
rect 3084 834 3118 868
rect 3174 834 3208 868
rect 3264 834 3298 868
rect 3354 834 3388 868
rect 3444 834 3478 868
rect 3534 834 3568 868
rect 3624 834 3658 868
rect 3084 744 3118 778
rect 3174 744 3208 778
rect 3264 744 3298 778
rect 3354 744 3388 778
rect 3444 744 3478 778
rect 3534 744 3568 778
rect 3624 744 3658 778
rect 3084 654 3118 688
rect 3174 654 3208 688
rect 3264 654 3298 688
rect 3354 654 3388 688
rect 3444 654 3478 688
rect 3534 654 3568 688
rect 3624 654 3658 688
rect 3084 564 3118 598
rect 3174 564 3208 598
rect 3264 564 3298 598
rect 3354 564 3388 598
rect 3444 564 3478 598
rect 3534 564 3568 598
rect 3624 564 3658 598
rect 3084 474 3118 508
rect 3174 474 3208 508
rect 3264 474 3298 508
rect 3354 474 3388 508
rect 3444 474 3478 508
rect 3534 474 3568 508
rect 3624 474 3658 508
rect 3084 384 3118 418
rect 3174 384 3208 418
rect 3264 384 3298 418
rect 3354 384 3388 418
rect 3444 384 3478 418
rect 3534 384 3568 418
rect 3624 384 3658 418
rect 4434 924 4468 958
rect 4524 924 4558 958
rect 4614 924 4648 958
rect 4704 924 4738 958
rect 4794 924 4828 958
rect 4884 924 4918 958
rect 4974 924 5008 958
rect 4434 834 4468 868
rect 4524 834 4558 868
rect 4614 834 4648 868
rect 4704 834 4738 868
rect 4794 834 4828 868
rect 4884 834 4918 868
rect 4974 834 5008 868
rect 4434 744 4468 778
rect 4524 744 4558 778
rect 4614 744 4648 778
rect 4704 744 4738 778
rect 4794 744 4828 778
rect 4884 744 4918 778
rect 4974 744 5008 778
rect 4434 654 4468 688
rect 4524 654 4558 688
rect 4614 654 4648 688
rect 4704 654 4738 688
rect 4794 654 4828 688
rect 4884 654 4918 688
rect 4974 654 5008 688
rect 4434 564 4468 598
rect 4524 564 4558 598
rect 4614 564 4648 598
rect 4704 564 4738 598
rect 4794 564 4828 598
rect 4884 564 4918 598
rect 4974 564 5008 598
rect 4434 474 4468 508
rect 4524 474 4558 508
rect 4614 474 4648 508
rect 4704 474 4738 508
rect 4794 474 4828 508
rect 4884 474 4918 508
rect 4974 474 5008 508
rect 4434 384 4468 418
rect 4524 384 4558 418
rect 4614 384 4648 418
rect 4704 384 4738 418
rect 4794 384 4828 418
rect 4884 384 4918 418
rect 4974 384 5008 418
rect 5784 924 5818 958
rect 5874 924 5908 958
rect 5964 924 5998 958
rect 6054 924 6088 958
rect 6144 924 6178 958
rect 6234 924 6268 958
rect 6324 924 6358 958
rect 5784 834 5818 868
rect 5874 834 5908 868
rect 5964 834 5998 868
rect 6054 834 6088 868
rect 6144 834 6178 868
rect 6234 834 6268 868
rect 6324 834 6358 868
rect 5784 744 5818 778
rect 5874 744 5908 778
rect 5964 744 5998 778
rect 6054 744 6088 778
rect 6144 744 6178 778
rect 6234 744 6268 778
rect 6324 744 6358 778
rect 5784 654 5818 688
rect 5874 654 5908 688
rect 5964 654 5998 688
rect 6054 654 6088 688
rect 6144 654 6178 688
rect 6234 654 6268 688
rect 6324 654 6358 688
rect 5784 564 5818 598
rect 5874 564 5908 598
rect 5964 564 5998 598
rect 6054 564 6088 598
rect 6144 564 6178 598
rect 6234 564 6268 598
rect 6324 564 6358 598
rect 5784 474 5818 508
rect 5874 474 5908 508
rect 5964 474 5998 508
rect 6054 474 6088 508
rect 6144 474 6178 508
rect 6234 474 6268 508
rect 6324 474 6358 508
rect 5784 384 5818 418
rect 5874 384 5908 418
rect 5964 384 5998 418
rect 6054 384 6088 418
rect 6144 384 6178 418
rect 6234 384 6268 418
rect 6324 384 6358 418
rect 7134 924 7168 958
rect 7224 924 7258 958
rect 7314 924 7348 958
rect 7404 924 7438 958
rect 7494 924 7528 958
rect 7584 924 7618 958
rect 7674 924 7708 958
rect 7134 834 7168 868
rect 7224 834 7258 868
rect 7314 834 7348 868
rect 7404 834 7438 868
rect 7494 834 7528 868
rect 7584 834 7618 868
rect 7674 834 7708 868
rect 7134 744 7168 778
rect 7224 744 7258 778
rect 7314 744 7348 778
rect 7404 744 7438 778
rect 7494 744 7528 778
rect 7584 744 7618 778
rect 7674 744 7708 778
rect 7134 654 7168 688
rect 7224 654 7258 688
rect 7314 654 7348 688
rect 7404 654 7438 688
rect 7494 654 7528 688
rect 7584 654 7618 688
rect 7674 654 7708 688
rect 7134 564 7168 598
rect 7224 564 7258 598
rect 7314 564 7348 598
rect 7404 564 7438 598
rect 7494 564 7528 598
rect 7584 564 7618 598
rect 7674 564 7708 598
rect 7134 474 7168 508
rect 7224 474 7258 508
rect 7314 474 7348 508
rect 7404 474 7438 508
rect 7494 474 7528 508
rect 7584 474 7618 508
rect 7674 474 7708 508
rect 7134 384 7168 418
rect 7224 384 7258 418
rect 7314 384 7348 418
rect 7404 384 7438 418
rect 7494 384 7528 418
rect 7584 384 7618 418
rect 7674 384 7708 418
rect 8484 924 8518 958
rect 8574 924 8608 958
rect 8664 924 8698 958
rect 8754 924 8788 958
rect 8844 924 8878 958
rect 8934 924 8968 958
rect 9024 924 9058 958
rect 8484 834 8518 868
rect 8574 834 8608 868
rect 8664 834 8698 868
rect 8754 834 8788 868
rect 8844 834 8878 868
rect 8934 834 8968 868
rect 9024 834 9058 868
rect 8484 744 8518 778
rect 8574 744 8608 778
rect 8664 744 8698 778
rect 8754 744 8788 778
rect 8844 744 8878 778
rect 8934 744 8968 778
rect 9024 744 9058 778
rect 8484 654 8518 688
rect 8574 654 8608 688
rect 8664 654 8698 688
rect 8754 654 8788 688
rect 8844 654 8878 688
rect 8934 654 8968 688
rect 9024 654 9058 688
rect 8484 564 8518 598
rect 8574 564 8608 598
rect 8664 564 8698 598
rect 8754 564 8788 598
rect 8844 564 8878 598
rect 8934 564 8968 598
rect 9024 564 9058 598
rect 8484 474 8518 508
rect 8574 474 8608 508
rect 8664 474 8698 508
rect 8754 474 8788 508
rect 8844 474 8878 508
rect 8934 474 8968 508
rect 9024 474 9058 508
rect 8484 384 8518 418
rect 8574 384 8608 418
rect 8664 384 8698 418
rect 8754 384 8788 418
rect 8844 384 8878 418
rect 8934 384 8968 418
rect 9024 384 9058 418
<< psubdiff >>
rect 1376 1279 2664 1314
rect 1376 1256 1506 1279
rect 1376 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2664 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2664 1256
rect 1376 1213 2664 1222
rect 1376 1166 1477 1213
rect 1376 1132 1410 1166
rect 1444 1132 1477 1166
rect 2563 1166 2664 1213
rect 1376 1076 1477 1132
rect 1376 1042 1410 1076
rect 1444 1042 1477 1076
rect 1376 986 1477 1042
rect 1376 952 1410 986
rect 1444 952 1477 986
rect 1376 896 1477 952
rect 1376 862 1410 896
rect 1444 862 1477 896
rect 1376 806 1477 862
rect 1376 772 1410 806
rect 1444 772 1477 806
rect 1376 716 1477 772
rect 1376 682 1410 716
rect 1444 682 1477 716
rect 1376 626 1477 682
rect 1376 592 1410 626
rect 1444 592 1477 626
rect 1376 536 1477 592
rect 1376 502 1410 536
rect 1444 502 1477 536
rect 1376 446 1477 502
rect 1376 412 1410 446
rect 1444 412 1477 446
rect 1376 356 1477 412
rect 1376 322 1410 356
rect 1444 322 1477 356
rect 1376 266 1477 322
rect 1376 232 1410 266
rect 1444 232 1477 266
rect 1376 176 1477 232
rect 2563 1132 2597 1166
rect 2631 1132 2664 1166
rect 2563 1076 2664 1132
rect 2563 1042 2597 1076
rect 2631 1042 2664 1076
rect 2563 986 2664 1042
rect 2563 952 2597 986
rect 2631 952 2664 986
rect 2563 896 2664 952
rect 2563 862 2597 896
rect 2631 862 2664 896
rect 2563 806 2664 862
rect 2563 772 2597 806
rect 2631 772 2664 806
rect 2563 716 2664 772
rect 2563 682 2597 716
rect 2631 682 2664 716
rect 2563 626 2664 682
rect 2563 592 2597 626
rect 2631 592 2664 626
rect 2563 536 2664 592
rect 2563 502 2597 536
rect 2631 502 2664 536
rect 2563 446 2664 502
rect 2563 412 2597 446
rect 2631 412 2664 446
rect 2563 356 2664 412
rect 2563 322 2597 356
rect 2631 322 2664 356
rect 2563 266 2664 322
rect 2563 232 2597 266
rect 2631 232 2664 266
rect 1376 142 1410 176
rect 1444 142 1477 176
rect 1376 127 1477 142
rect 2563 176 2664 232
rect 2563 142 2597 176
rect 2631 142 2664 176
rect 2563 127 2664 142
rect 1376 92 2664 127
rect 1376 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 58 2664 92
rect 1376 26 2664 58
rect 2726 1279 4014 1314
rect 2726 1256 2856 1279
rect 2726 1222 2760 1256
rect 2794 1245 2856 1256
rect 2890 1245 2946 1279
rect 2980 1245 3036 1279
rect 3070 1245 3126 1279
rect 3160 1245 3216 1279
rect 3250 1245 3306 1279
rect 3340 1245 3396 1279
rect 3430 1245 3486 1279
rect 3520 1245 3576 1279
rect 3610 1245 3666 1279
rect 3700 1245 3756 1279
rect 3790 1245 3846 1279
rect 3880 1256 4014 1279
rect 3880 1245 3947 1256
rect 2794 1222 3947 1245
rect 3981 1222 4014 1256
rect 2726 1213 4014 1222
rect 2726 1166 2827 1213
rect 2726 1132 2760 1166
rect 2794 1132 2827 1166
rect 3913 1166 4014 1213
rect 2726 1076 2827 1132
rect 2726 1042 2760 1076
rect 2794 1042 2827 1076
rect 2726 986 2827 1042
rect 2726 952 2760 986
rect 2794 952 2827 986
rect 2726 896 2827 952
rect 2726 862 2760 896
rect 2794 862 2827 896
rect 2726 806 2827 862
rect 2726 772 2760 806
rect 2794 772 2827 806
rect 2726 716 2827 772
rect 2726 682 2760 716
rect 2794 682 2827 716
rect 2726 626 2827 682
rect 2726 592 2760 626
rect 2794 592 2827 626
rect 2726 536 2827 592
rect 2726 502 2760 536
rect 2794 502 2827 536
rect 2726 446 2827 502
rect 2726 412 2760 446
rect 2794 412 2827 446
rect 2726 356 2827 412
rect 2726 322 2760 356
rect 2794 322 2827 356
rect 2726 266 2827 322
rect 2726 232 2760 266
rect 2794 232 2827 266
rect 2726 176 2827 232
rect 3913 1132 3947 1166
rect 3981 1132 4014 1166
rect 3913 1076 4014 1132
rect 3913 1042 3947 1076
rect 3981 1042 4014 1076
rect 3913 986 4014 1042
rect 3913 952 3947 986
rect 3981 952 4014 986
rect 3913 896 4014 952
rect 3913 862 3947 896
rect 3981 862 4014 896
rect 3913 806 4014 862
rect 3913 772 3947 806
rect 3981 772 4014 806
rect 3913 716 4014 772
rect 3913 682 3947 716
rect 3981 682 4014 716
rect 3913 626 4014 682
rect 3913 592 3947 626
rect 3981 592 4014 626
rect 3913 536 4014 592
rect 3913 502 3947 536
rect 3981 502 4014 536
rect 3913 446 4014 502
rect 3913 412 3947 446
rect 3981 412 4014 446
rect 3913 356 4014 412
rect 3913 322 3947 356
rect 3981 322 4014 356
rect 3913 266 4014 322
rect 3913 232 3947 266
rect 3981 232 4014 266
rect 2726 142 2760 176
rect 2794 142 2827 176
rect 2726 127 2827 142
rect 3913 176 4014 232
rect 3913 142 3947 176
rect 3981 142 4014 176
rect 3913 127 4014 142
rect 2726 92 4014 127
rect 2726 58 2856 92
rect 2890 58 2946 92
rect 2980 58 3036 92
rect 3070 58 3126 92
rect 3160 58 3216 92
rect 3250 58 3306 92
rect 3340 58 3396 92
rect 3430 58 3486 92
rect 3520 58 3576 92
rect 3610 58 3666 92
rect 3700 58 3756 92
rect 3790 58 3846 92
rect 3880 58 4014 92
rect 2726 26 4014 58
rect 4076 1279 5364 1314
rect 4076 1256 4206 1279
rect 4076 1222 4110 1256
rect 4144 1245 4206 1256
rect 4240 1245 4296 1279
rect 4330 1245 4386 1279
rect 4420 1245 4476 1279
rect 4510 1245 4566 1279
rect 4600 1245 4656 1279
rect 4690 1245 4746 1279
rect 4780 1245 4836 1279
rect 4870 1245 4926 1279
rect 4960 1245 5016 1279
rect 5050 1245 5106 1279
rect 5140 1245 5196 1279
rect 5230 1256 5364 1279
rect 5230 1245 5297 1256
rect 4144 1222 5297 1245
rect 5331 1222 5364 1256
rect 4076 1213 5364 1222
rect 4076 1166 4177 1213
rect 4076 1132 4110 1166
rect 4144 1132 4177 1166
rect 5263 1166 5364 1213
rect 4076 1076 4177 1132
rect 4076 1042 4110 1076
rect 4144 1042 4177 1076
rect 4076 986 4177 1042
rect 4076 952 4110 986
rect 4144 952 4177 986
rect 4076 896 4177 952
rect 4076 862 4110 896
rect 4144 862 4177 896
rect 4076 806 4177 862
rect 4076 772 4110 806
rect 4144 772 4177 806
rect 4076 716 4177 772
rect 4076 682 4110 716
rect 4144 682 4177 716
rect 4076 626 4177 682
rect 4076 592 4110 626
rect 4144 592 4177 626
rect 4076 536 4177 592
rect 4076 502 4110 536
rect 4144 502 4177 536
rect 4076 446 4177 502
rect 4076 412 4110 446
rect 4144 412 4177 446
rect 4076 356 4177 412
rect 4076 322 4110 356
rect 4144 322 4177 356
rect 4076 266 4177 322
rect 4076 232 4110 266
rect 4144 232 4177 266
rect 4076 176 4177 232
rect 5263 1132 5297 1166
rect 5331 1132 5364 1166
rect 5263 1076 5364 1132
rect 5263 1042 5297 1076
rect 5331 1042 5364 1076
rect 5263 986 5364 1042
rect 5263 952 5297 986
rect 5331 952 5364 986
rect 5263 896 5364 952
rect 5263 862 5297 896
rect 5331 862 5364 896
rect 5263 806 5364 862
rect 5263 772 5297 806
rect 5331 772 5364 806
rect 5263 716 5364 772
rect 5263 682 5297 716
rect 5331 682 5364 716
rect 5263 626 5364 682
rect 5263 592 5297 626
rect 5331 592 5364 626
rect 5263 536 5364 592
rect 5263 502 5297 536
rect 5331 502 5364 536
rect 5263 446 5364 502
rect 5263 412 5297 446
rect 5331 412 5364 446
rect 5263 356 5364 412
rect 5263 322 5297 356
rect 5331 322 5364 356
rect 5263 266 5364 322
rect 5263 232 5297 266
rect 5331 232 5364 266
rect 4076 142 4110 176
rect 4144 142 4177 176
rect 4076 127 4177 142
rect 5263 176 5364 232
rect 5263 142 5297 176
rect 5331 142 5364 176
rect 5263 127 5364 142
rect 4076 92 5364 127
rect 4076 58 4206 92
rect 4240 58 4296 92
rect 4330 58 4386 92
rect 4420 58 4476 92
rect 4510 58 4566 92
rect 4600 58 4656 92
rect 4690 58 4746 92
rect 4780 58 4836 92
rect 4870 58 4926 92
rect 4960 58 5016 92
rect 5050 58 5106 92
rect 5140 58 5196 92
rect 5230 58 5364 92
rect 4076 26 5364 58
rect 5426 1279 6714 1314
rect 5426 1256 5556 1279
rect 5426 1222 5460 1256
rect 5494 1245 5556 1256
rect 5590 1245 5646 1279
rect 5680 1245 5736 1279
rect 5770 1245 5826 1279
rect 5860 1245 5916 1279
rect 5950 1245 6006 1279
rect 6040 1245 6096 1279
rect 6130 1245 6186 1279
rect 6220 1245 6276 1279
rect 6310 1245 6366 1279
rect 6400 1245 6456 1279
rect 6490 1245 6546 1279
rect 6580 1256 6714 1279
rect 6580 1245 6647 1256
rect 5494 1222 6647 1245
rect 6681 1222 6714 1256
rect 5426 1213 6714 1222
rect 5426 1166 5527 1213
rect 5426 1132 5460 1166
rect 5494 1132 5527 1166
rect 6613 1166 6714 1213
rect 5426 1076 5527 1132
rect 5426 1042 5460 1076
rect 5494 1042 5527 1076
rect 5426 986 5527 1042
rect 5426 952 5460 986
rect 5494 952 5527 986
rect 5426 896 5527 952
rect 5426 862 5460 896
rect 5494 862 5527 896
rect 5426 806 5527 862
rect 5426 772 5460 806
rect 5494 772 5527 806
rect 5426 716 5527 772
rect 5426 682 5460 716
rect 5494 682 5527 716
rect 5426 626 5527 682
rect 5426 592 5460 626
rect 5494 592 5527 626
rect 5426 536 5527 592
rect 5426 502 5460 536
rect 5494 502 5527 536
rect 5426 446 5527 502
rect 5426 412 5460 446
rect 5494 412 5527 446
rect 5426 356 5527 412
rect 5426 322 5460 356
rect 5494 322 5527 356
rect 5426 266 5527 322
rect 5426 232 5460 266
rect 5494 232 5527 266
rect 5426 176 5527 232
rect 6613 1132 6647 1166
rect 6681 1132 6714 1166
rect 6613 1076 6714 1132
rect 6613 1042 6647 1076
rect 6681 1042 6714 1076
rect 6613 986 6714 1042
rect 6613 952 6647 986
rect 6681 952 6714 986
rect 6613 896 6714 952
rect 6613 862 6647 896
rect 6681 862 6714 896
rect 6613 806 6714 862
rect 6613 772 6647 806
rect 6681 772 6714 806
rect 6613 716 6714 772
rect 6613 682 6647 716
rect 6681 682 6714 716
rect 6613 626 6714 682
rect 6613 592 6647 626
rect 6681 592 6714 626
rect 6613 536 6714 592
rect 6613 502 6647 536
rect 6681 502 6714 536
rect 6613 446 6714 502
rect 6613 412 6647 446
rect 6681 412 6714 446
rect 6613 356 6714 412
rect 6613 322 6647 356
rect 6681 322 6714 356
rect 6613 266 6714 322
rect 6613 232 6647 266
rect 6681 232 6714 266
rect 5426 142 5460 176
rect 5494 142 5527 176
rect 5426 127 5527 142
rect 6613 176 6714 232
rect 6613 142 6647 176
rect 6681 142 6714 176
rect 6613 127 6714 142
rect 5426 92 6714 127
rect 5426 58 5556 92
rect 5590 58 5646 92
rect 5680 58 5736 92
rect 5770 58 5826 92
rect 5860 58 5916 92
rect 5950 58 6006 92
rect 6040 58 6096 92
rect 6130 58 6186 92
rect 6220 58 6276 92
rect 6310 58 6366 92
rect 6400 58 6456 92
rect 6490 58 6546 92
rect 6580 58 6714 92
rect 5426 26 6714 58
rect 6776 1279 8064 1314
rect 6776 1256 6906 1279
rect 6776 1222 6810 1256
rect 6844 1245 6906 1256
rect 6940 1245 6996 1279
rect 7030 1245 7086 1279
rect 7120 1245 7176 1279
rect 7210 1245 7266 1279
rect 7300 1245 7356 1279
rect 7390 1245 7446 1279
rect 7480 1245 7536 1279
rect 7570 1245 7626 1279
rect 7660 1245 7716 1279
rect 7750 1245 7806 1279
rect 7840 1245 7896 1279
rect 7930 1256 8064 1279
rect 7930 1245 7997 1256
rect 6844 1222 7997 1245
rect 8031 1222 8064 1256
rect 6776 1213 8064 1222
rect 6776 1166 6877 1213
rect 6776 1132 6810 1166
rect 6844 1132 6877 1166
rect 7963 1166 8064 1213
rect 6776 1076 6877 1132
rect 6776 1042 6810 1076
rect 6844 1042 6877 1076
rect 6776 986 6877 1042
rect 6776 952 6810 986
rect 6844 952 6877 986
rect 6776 896 6877 952
rect 6776 862 6810 896
rect 6844 862 6877 896
rect 6776 806 6877 862
rect 6776 772 6810 806
rect 6844 772 6877 806
rect 6776 716 6877 772
rect 6776 682 6810 716
rect 6844 682 6877 716
rect 6776 626 6877 682
rect 6776 592 6810 626
rect 6844 592 6877 626
rect 6776 536 6877 592
rect 6776 502 6810 536
rect 6844 502 6877 536
rect 6776 446 6877 502
rect 6776 412 6810 446
rect 6844 412 6877 446
rect 6776 356 6877 412
rect 6776 322 6810 356
rect 6844 322 6877 356
rect 6776 266 6877 322
rect 6776 232 6810 266
rect 6844 232 6877 266
rect 6776 176 6877 232
rect 7963 1132 7997 1166
rect 8031 1132 8064 1166
rect 7963 1076 8064 1132
rect 7963 1042 7997 1076
rect 8031 1042 8064 1076
rect 7963 986 8064 1042
rect 7963 952 7997 986
rect 8031 952 8064 986
rect 7963 896 8064 952
rect 7963 862 7997 896
rect 8031 862 8064 896
rect 7963 806 8064 862
rect 7963 772 7997 806
rect 8031 772 8064 806
rect 7963 716 8064 772
rect 7963 682 7997 716
rect 8031 682 8064 716
rect 7963 626 8064 682
rect 7963 592 7997 626
rect 8031 592 8064 626
rect 7963 536 8064 592
rect 7963 502 7997 536
rect 8031 502 8064 536
rect 7963 446 8064 502
rect 7963 412 7997 446
rect 8031 412 8064 446
rect 7963 356 8064 412
rect 7963 322 7997 356
rect 8031 322 8064 356
rect 7963 266 8064 322
rect 7963 232 7997 266
rect 8031 232 8064 266
rect 6776 142 6810 176
rect 6844 142 6877 176
rect 6776 127 6877 142
rect 7963 176 8064 232
rect 7963 142 7997 176
rect 8031 142 8064 176
rect 7963 127 8064 142
rect 6776 92 8064 127
rect 6776 58 6906 92
rect 6940 58 6996 92
rect 7030 58 7086 92
rect 7120 58 7176 92
rect 7210 58 7266 92
rect 7300 58 7356 92
rect 7390 58 7446 92
rect 7480 58 7536 92
rect 7570 58 7626 92
rect 7660 58 7716 92
rect 7750 58 7806 92
rect 7840 58 7896 92
rect 7930 58 8064 92
rect 6776 26 8064 58
rect 8126 1279 9414 1314
rect 8126 1256 8256 1279
rect 8126 1222 8160 1256
rect 8194 1245 8256 1256
rect 8290 1245 8346 1279
rect 8380 1245 8436 1279
rect 8470 1245 8526 1279
rect 8560 1245 8616 1279
rect 8650 1245 8706 1279
rect 8740 1245 8796 1279
rect 8830 1245 8886 1279
rect 8920 1245 8976 1279
rect 9010 1245 9066 1279
rect 9100 1245 9156 1279
rect 9190 1245 9246 1279
rect 9280 1256 9414 1279
rect 9280 1245 9347 1256
rect 8194 1222 9347 1245
rect 9381 1222 9414 1256
rect 8126 1213 9414 1222
rect 8126 1166 8227 1213
rect 8126 1132 8160 1166
rect 8194 1132 8227 1166
rect 9313 1166 9414 1213
rect 8126 1076 8227 1132
rect 8126 1042 8160 1076
rect 8194 1042 8227 1076
rect 8126 986 8227 1042
rect 8126 952 8160 986
rect 8194 952 8227 986
rect 8126 896 8227 952
rect 8126 862 8160 896
rect 8194 862 8227 896
rect 8126 806 8227 862
rect 8126 772 8160 806
rect 8194 772 8227 806
rect 8126 716 8227 772
rect 8126 682 8160 716
rect 8194 682 8227 716
rect 8126 626 8227 682
rect 8126 592 8160 626
rect 8194 592 8227 626
rect 8126 536 8227 592
rect 8126 502 8160 536
rect 8194 502 8227 536
rect 8126 446 8227 502
rect 8126 412 8160 446
rect 8194 412 8227 446
rect 8126 356 8227 412
rect 8126 322 8160 356
rect 8194 322 8227 356
rect 8126 266 8227 322
rect 8126 232 8160 266
rect 8194 232 8227 266
rect 8126 176 8227 232
rect 9313 1132 9347 1166
rect 9381 1132 9414 1166
rect 9313 1076 9414 1132
rect 9313 1042 9347 1076
rect 9381 1042 9414 1076
rect 9313 986 9414 1042
rect 9313 952 9347 986
rect 9381 952 9414 986
rect 9313 896 9414 952
rect 9313 862 9347 896
rect 9381 862 9414 896
rect 9313 806 9414 862
rect 9313 772 9347 806
rect 9381 772 9414 806
rect 9313 716 9414 772
rect 9313 682 9347 716
rect 9381 682 9414 716
rect 9313 626 9414 682
rect 9313 592 9347 626
rect 9381 592 9414 626
rect 9313 536 9414 592
rect 9313 502 9347 536
rect 9381 502 9414 536
rect 9313 446 9414 502
rect 9313 412 9347 446
rect 9381 412 9414 446
rect 9313 356 9414 412
rect 9313 322 9347 356
rect 9381 322 9414 356
rect 9313 266 9414 322
rect 9313 232 9347 266
rect 9381 232 9414 266
rect 8126 142 8160 176
rect 8194 142 8227 176
rect 8126 127 8227 142
rect 9313 176 9414 232
rect 9313 142 9347 176
rect 9381 142 9414 176
rect 9313 127 9414 142
rect 8126 92 9414 127
rect 8126 58 8256 92
rect 8290 58 8346 92
rect 8380 58 8436 92
rect 8470 58 8526 92
rect 8560 58 8616 92
rect 8650 58 8706 92
rect 8740 58 8796 92
rect 8830 58 8886 92
rect 8920 58 8976 92
rect 9010 58 9066 92
rect 9100 58 9156 92
rect 9190 58 9246 92
rect 9280 58 9414 92
rect 8126 26 9414 58
<< nsubdiff >>
rect 1539 1132 2501 1151
rect 1539 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 2501 1132
rect 1539 1079 2501 1098
rect 1539 1075 1611 1079
rect 1539 1041 1558 1075
rect 1592 1041 1611 1075
rect 1539 985 1611 1041
rect 2429 1056 2501 1079
rect 2429 1022 2448 1056
rect 2482 1022 2501 1056
rect 1539 951 1558 985
rect 1592 951 1611 985
rect 1539 895 1611 951
rect 1539 861 1558 895
rect 1592 861 1611 895
rect 1539 805 1611 861
rect 1539 771 1558 805
rect 1592 771 1611 805
rect 1539 715 1611 771
rect 1539 681 1558 715
rect 1592 681 1611 715
rect 1539 625 1611 681
rect 1539 591 1558 625
rect 1592 591 1611 625
rect 1539 535 1611 591
rect 1539 501 1558 535
rect 1592 501 1611 535
rect 1539 445 1611 501
rect 1539 411 1558 445
rect 1592 411 1611 445
rect 1539 355 1611 411
rect 1539 321 1558 355
rect 1592 321 1611 355
rect 2429 966 2501 1022
rect 2429 932 2448 966
rect 2482 932 2501 966
rect 2429 876 2501 932
rect 2429 842 2448 876
rect 2482 842 2501 876
rect 2429 786 2501 842
rect 2429 752 2448 786
rect 2482 752 2501 786
rect 2429 696 2501 752
rect 2429 662 2448 696
rect 2482 662 2501 696
rect 2429 606 2501 662
rect 2429 572 2448 606
rect 2482 572 2501 606
rect 2429 516 2501 572
rect 2429 482 2448 516
rect 2482 482 2501 516
rect 2429 426 2501 482
rect 2429 392 2448 426
rect 2482 392 2501 426
rect 2429 336 2501 392
rect 1539 261 1611 321
rect 2429 302 2448 336
rect 2482 302 2501 336
rect 2429 261 2501 302
rect 1539 242 2501 261
rect 1539 208 1636 242
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 208 2501 242
rect 1539 189 2501 208
rect 2889 1132 3851 1151
rect 2889 1098 3020 1132
rect 3054 1098 3110 1132
rect 3144 1098 3200 1132
rect 3234 1098 3290 1132
rect 3324 1098 3380 1132
rect 3414 1098 3470 1132
rect 3504 1098 3560 1132
rect 3594 1098 3650 1132
rect 3684 1098 3740 1132
rect 3774 1098 3851 1132
rect 2889 1079 3851 1098
rect 2889 1075 2961 1079
rect 2889 1041 2908 1075
rect 2942 1041 2961 1075
rect 2889 985 2961 1041
rect 3779 1056 3851 1079
rect 3779 1022 3798 1056
rect 3832 1022 3851 1056
rect 2889 951 2908 985
rect 2942 951 2961 985
rect 2889 895 2961 951
rect 2889 861 2908 895
rect 2942 861 2961 895
rect 2889 805 2961 861
rect 2889 771 2908 805
rect 2942 771 2961 805
rect 2889 715 2961 771
rect 2889 681 2908 715
rect 2942 681 2961 715
rect 2889 625 2961 681
rect 2889 591 2908 625
rect 2942 591 2961 625
rect 2889 535 2961 591
rect 2889 501 2908 535
rect 2942 501 2961 535
rect 2889 445 2961 501
rect 2889 411 2908 445
rect 2942 411 2961 445
rect 2889 355 2961 411
rect 2889 321 2908 355
rect 2942 321 2961 355
rect 3779 966 3851 1022
rect 3779 932 3798 966
rect 3832 932 3851 966
rect 3779 876 3851 932
rect 3779 842 3798 876
rect 3832 842 3851 876
rect 3779 786 3851 842
rect 3779 752 3798 786
rect 3832 752 3851 786
rect 3779 696 3851 752
rect 3779 662 3798 696
rect 3832 662 3851 696
rect 3779 606 3851 662
rect 3779 572 3798 606
rect 3832 572 3851 606
rect 3779 516 3851 572
rect 3779 482 3798 516
rect 3832 482 3851 516
rect 3779 426 3851 482
rect 3779 392 3798 426
rect 3832 392 3851 426
rect 3779 336 3851 392
rect 2889 261 2961 321
rect 3779 302 3798 336
rect 3832 302 3851 336
rect 3779 261 3851 302
rect 2889 242 3851 261
rect 2889 208 2986 242
rect 3020 208 3076 242
rect 3110 208 3166 242
rect 3200 208 3256 242
rect 3290 208 3346 242
rect 3380 208 3436 242
rect 3470 208 3526 242
rect 3560 208 3616 242
rect 3650 208 3706 242
rect 3740 208 3851 242
rect 2889 189 3851 208
rect 4239 1132 5201 1151
rect 4239 1098 4370 1132
rect 4404 1098 4460 1132
rect 4494 1098 4550 1132
rect 4584 1098 4640 1132
rect 4674 1098 4730 1132
rect 4764 1098 4820 1132
rect 4854 1098 4910 1132
rect 4944 1098 5000 1132
rect 5034 1098 5090 1132
rect 5124 1098 5201 1132
rect 4239 1079 5201 1098
rect 4239 1075 4311 1079
rect 4239 1041 4258 1075
rect 4292 1041 4311 1075
rect 4239 985 4311 1041
rect 5129 1056 5201 1079
rect 5129 1022 5148 1056
rect 5182 1022 5201 1056
rect 4239 951 4258 985
rect 4292 951 4311 985
rect 4239 895 4311 951
rect 4239 861 4258 895
rect 4292 861 4311 895
rect 4239 805 4311 861
rect 4239 771 4258 805
rect 4292 771 4311 805
rect 4239 715 4311 771
rect 4239 681 4258 715
rect 4292 681 4311 715
rect 4239 625 4311 681
rect 4239 591 4258 625
rect 4292 591 4311 625
rect 4239 535 4311 591
rect 4239 501 4258 535
rect 4292 501 4311 535
rect 4239 445 4311 501
rect 4239 411 4258 445
rect 4292 411 4311 445
rect 4239 355 4311 411
rect 4239 321 4258 355
rect 4292 321 4311 355
rect 5129 966 5201 1022
rect 5129 932 5148 966
rect 5182 932 5201 966
rect 5129 876 5201 932
rect 5129 842 5148 876
rect 5182 842 5201 876
rect 5129 786 5201 842
rect 5129 752 5148 786
rect 5182 752 5201 786
rect 5129 696 5201 752
rect 5129 662 5148 696
rect 5182 662 5201 696
rect 5129 606 5201 662
rect 5129 572 5148 606
rect 5182 572 5201 606
rect 5129 516 5201 572
rect 5129 482 5148 516
rect 5182 482 5201 516
rect 5129 426 5201 482
rect 5129 392 5148 426
rect 5182 392 5201 426
rect 5129 336 5201 392
rect 4239 261 4311 321
rect 5129 302 5148 336
rect 5182 302 5201 336
rect 5129 261 5201 302
rect 4239 242 5201 261
rect 4239 208 4336 242
rect 4370 208 4426 242
rect 4460 208 4516 242
rect 4550 208 4606 242
rect 4640 208 4696 242
rect 4730 208 4786 242
rect 4820 208 4876 242
rect 4910 208 4966 242
rect 5000 208 5056 242
rect 5090 208 5201 242
rect 4239 189 5201 208
rect 5589 1132 6551 1151
rect 5589 1098 5720 1132
rect 5754 1098 5810 1132
rect 5844 1098 5900 1132
rect 5934 1098 5990 1132
rect 6024 1098 6080 1132
rect 6114 1098 6170 1132
rect 6204 1098 6260 1132
rect 6294 1098 6350 1132
rect 6384 1098 6440 1132
rect 6474 1098 6551 1132
rect 5589 1079 6551 1098
rect 5589 1075 5661 1079
rect 5589 1041 5608 1075
rect 5642 1041 5661 1075
rect 5589 985 5661 1041
rect 6479 1056 6551 1079
rect 6479 1022 6498 1056
rect 6532 1022 6551 1056
rect 5589 951 5608 985
rect 5642 951 5661 985
rect 5589 895 5661 951
rect 5589 861 5608 895
rect 5642 861 5661 895
rect 5589 805 5661 861
rect 5589 771 5608 805
rect 5642 771 5661 805
rect 5589 715 5661 771
rect 5589 681 5608 715
rect 5642 681 5661 715
rect 5589 625 5661 681
rect 5589 591 5608 625
rect 5642 591 5661 625
rect 5589 535 5661 591
rect 5589 501 5608 535
rect 5642 501 5661 535
rect 5589 445 5661 501
rect 5589 411 5608 445
rect 5642 411 5661 445
rect 5589 355 5661 411
rect 5589 321 5608 355
rect 5642 321 5661 355
rect 6479 966 6551 1022
rect 6479 932 6498 966
rect 6532 932 6551 966
rect 6479 876 6551 932
rect 6479 842 6498 876
rect 6532 842 6551 876
rect 6479 786 6551 842
rect 6479 752 6498 786
rect 6532 752 6551 786
rect 6479 696 6551 752
rect 6479 662 6498 696
rect 6532 662 6551 696
rect 6479 606 6551 662
rect 6479 572 6498 606
rect 6532 572 6551 606
rect 6479 516 6551 572
rect 6479 482 6498 516
rect 6532 482 6551 516
rect 6479 426 6551 482
rect 6479 392 6498 426
rect 6532 392 6551 426
rect 6479 336 6551 392
rect 5589 261 5661 321
rect 6479 302 6498 336
rect 6532 302 6551 336
rect 6479 261 6551 302
rect 5589 242 6551 261
rect 5589 208 5686 242
rect 5720 208 5776 242
rect 5810 208 5866 242
rect 5900 208 5956 242
rect 5990 208 6046 242
rect 6080 208 6136 242
rect 6170 208 6226 242
rect 6260 208 6316 242
rect 6350 208 6406 242
rect 6440 208 6551 242
rect 5589 189 6551 208
rect 6939 1132 7901 1151
rect 6939 1098 7070 1132
rect 7104 1098 7160 1132
rect 7194 1098 7250 1132
rect 7284 1098 7340 1132
rect 7374 1098 7430 1132
rect 7464 1098 7520 1132
rect 7554 1098 7610 1132
rect 7644 1098 7700 1132
rect 7734 1098 7790 1132
rect 7824 1098 7901 1132
rect 6939 1079 7901 1098
rect 6939 1075 7011 1079
rect 6939 1041 6958 1075
rect 6992 1041 7011 1075
rect 6939 985 7011 1041
rect 7829 1056 7901 1079
rect 7829 1022 7848 1056
rect 7882 1022 7901 1056
rect 6939 951 6958 985
rect 6992 951 7011 985
rect 6939 895 7011 951
rect 6939 861 6958 895
rect 6992 861 7011 895
rect 6939 805 7011 861
rect 6939 771 6958 805
rect 6992 771 7011 805
rect 6939 715 7011 771
rect 6939 681 6958 715
rect 6992 681 7011 715
rect 6939 625 7011 681
rect 6939 591 6958 625
rect 6992 591 7011 625
rect 6939 535 7011 591
rect 6939 501 6958 535
rect 6992 501 7011 535
rect 6939 445 7011 501
rect 6939 411 6958 445
rect 6992 411 7011 445
rect 6939 355 7011 411
rect 6939 321 6958 355
rect 6992 321 7011 355
rect 7829 966 7901 1022
rect 7829 932 7848 966
rect 7882 932 7901 966
rect 7829 876 7901 932
rect 7829 842 7848 876
rect 7882 842 7901 876
rect 7829 786 7901 842
rect 7829 752 7848 786
rect 7882 752 7901 786
rect 7829 696 7901 752
rect 7829 662 7848 696
rect 7882 662 7901 696
rect 7829 606 7901 662
rect 7829 572 7848 606
rect 7882 572 7901 606
rect 7829 516 7901 572
rect 7829 482 7848 516
rect 7882 482 7901 516
rect 7829 426 7901 482
rect 7829 392 7848 426
rect 7882 392 7901 426
rect 7829 336 7901 392
rect 6939 261 7011 321
rect 7829 302 7848 336
rect 7882 302 7901 336
rect 7829 261 7901 302
rect 6939 242 7901 261
rect 6939 208 7036 242
rect 7070 208 7126 242
rect 7160 208 7216 242
rect 7250 208 7306 242
rect 7340 208 7396 242
rect 7430 208 7486 242
rect 7520 208 7576 242
rect 7610 208 7666 242
rect 7700 208 7756 242
rect 7790 208 7901 242
rect 6939 189 7901 208
rect 8289 1132 9251 1151
rect 8289 1098 8420 1132
rect 8454 1098 8510 1132
rect 8544 1098 8600 1132
rect 8634 1098 8690 1132
rect 8724 1098 8780 1132
rect 8814 1098 8870 1132
rect 8904 1098 8960 1132
rect 8994 1098 9050 1132
rect 9084 1098 9140 1132
rect 9174 1098 9251 1132
rect 8289 1079 9251 1098
rect 8289 1075 8361 1079
rect 8289 1041 8308 1075
rect 8342 1041 8361 1075
rect 8289 985 8361 1041
rect 9179 1056 9251 1079
rect 9179 1022 9198 1056
rect 9232 1022 9251 1056
rect 8289 951 8308 985
rect 8342 951 8361 985
rect 8289 895 8361 951
rect 8289 861 8308 895
rect 8342 861 8361 895
rect 8289 805 8361 861
rect 8289 771 8308 805
rect 8342 771 8361 805
rect 8289 715 8361 771
rect 8289 681 8308 715
rect 8342 681 8361 715
rect 8289 625 8361 681
rect 8289 591 8308 625
rect 8342 591 8361 625
rect 8289 535 8361 591
rect 8289 501 8308 535
rect 8342 501 8361 535
rect 8289 445 8361 501
rect 8289 411 8308 445
rect 8342 411 8361 445
rect 8289 355 8361 411
rect 8289 321 8308 355
rect 8342 321 8361 355
rect 9179 966 9251 1022
rect 9179 932 9198 966
rect 9232 932 9251 966
rect 9179 876 9251 932
rect 9179 842 9198 876
rect 9232 842 9251 876
rect 9179 786 9251 842
rect 9179 752 9198 786
rect 9232 752 9251 786
rect 9179 696 9251 752
rect 9179 662 9198 696
rect 9232 662 9251 696
rect 9179 606 9251 662
rect 9179 572 9198 606
rect 9232 572 9251 606
rect 9179 516 9251 572
rect 9179 482 9198 516
rect 9232 482 9251 516
rect 9179 426 9251 482
rect 9179 392 9198 426
rect 9232 392 9251 426
rect 9179 336 9251 392
rect 8289 261 8361 321
rect 9179 302 9198 336
rect 9232 302 9251 336
rect 9179 261 9251 302
rect 8289 242 9251 261
rect 8289 208 8386 242
rect 8420 208 8476 242
rect 8510 208 8566 242
rect 8600 208 8656 242
rect 8690 208 8746 242
rect 8780 208 8836 242
rect 8870 208 8926 242
rect 8960 208 9016 242
rect 9050 208 9106 242
rect 9140 208 9251 242
rect 8289 189 9251 208
<< psubdiffcont >>
rect 1410 1222 1444 1256
rect 1506 1245 1540 1279
rect 1596 1245 1630 1279
rect 1686 1245 1720 1279
rect 1776 1245 1810 1279
rect 1866 1245 1900 1279
rect 1956 1245 1990 1279
rect 2046 1245 2080 1279
rect 2136 1245 2170 1279
rect 2226 1245 2260 1279
rect 2316 1245 2350 1279
rect 2406 1245 2440 1279
rect 2496 1245 2530 1279
rect 2597 1222 2631 1256
rect 1410 1132 1444 1166
rect 1410 1042 1444 1076
rect 1410 952 1444 986
rect 1410 862 1444 896
rect 1410 772 1444 806
rect 1410 682 1444 716
rect 1410 592 1444 626
rect 1410 502 1444 536
rect 1410 412 1444 446
rect 1410 322 1444 356
rect 1410 232 1444 266
rect 2597 1132 2631 1166
rect 2597 1042 2631 1076
rect 2597 952 2631 986
rect 2597 862 2631 896
rect 2597 772 2631 806
rect 2597 682 2631 716
rect 2597 592 2631 626
rect 2597 502 2631 536
rect 2597 412 2631 446
rect 2597 322 2631 356
rect 2597 232 2631 266
rect 1410 142 1444 176
rect 2597 142 2631 176
rect 1506 58 1540 92
rect 1596 58 1630 92
rect 1686 58 1720 92
rect 1776 58 1810 92
rect 1866 58 1900 92
rect 1956 58 1990 92
rect 2046 58 2080 92
rect 2136 58 2170 92
rect 2226 58 2260 92
rect 2316 58 2350 92
rect 2406 58 2440 92
rect 2496 58 2530 92
rect 2760 1222 2794 1256
rect 2856 1245 2890 1279
rect 2946 1245 2980 1279
rect 3036 1245 3070 1279
rect 3126 1245 3160 1279
rect 3216 1245 3250 1279
rect 3306 1245 3340 1279
rect 3396 1245 3430 1279
rect 3486 1245 3520 1279
rect 3576 1245 3610 1279
rect 3666 1245 3700 1279
rect 3756 1245 3790 1279
rect 3846 1245 3880 1279
rect 3947 1222 3981 1256
rect 2760 1132 2794 1166
rect 2760 1042 2794 1076
rect 2760 952 2794 986
rect 2760 862 2794 896
rect 2760 772 2794 806
rect 2760 682 2794 716
rect 2760 592 2794 626
rect 2760 502 2794 536
rect 2760 412 2794 446
rect 2760 322 2794 356
rect 2760 232 2794 266
rect 3947 1132 3981 1166
rect 3947 1042 3981 1076
rect 3947 952 3981 986
rect 3947 862 3981 896
rect 3947 772 3981 806
rect 3947 682 3981 716
rect 3947 592 3981 626
rect 3947 502 3981 536
rect 3947 412 3981 446
rect 3947 322 3981 356
rect 3947 232 3981 266
rect 2760 142 2794 176
rect 3947 142 3981 176
rect 2856 58 2890 92
rect 2946 58 2980 92
rect 3036 58 3070 92
rect 3126 58 3160 92
rect 3216 58 3250 92
rect 3306 58 3340 92
rect 3396 58 3430 92
rect 3486 58 3520 92
rect 3576 58 3610 92
rect 3666 58 3700 92
rect 3756 58 3790 92
rect 3846 58 3880 92
rect 4110 1222 4144 1256
rect 4206 1245 4240 1279
rect 4296 1245 4330 1279
rect 4386 1245 4420 1279
rect 4476 1245 4510 1279
rect 4566 1245 4600 1279
rect 4656 1245 4690 1279
rect 4746 1245 4780 1279
rect 4836 1245 4870 1279
rect 4926 1245 4960 1279
rect 5016 1245 5050 1279
rect 5106 1245 5140 1279
rect 5196 1245 5230 1279
rect 5297 1222 5331 1256
rect 4110 1132 4144 1166
rect 4110 1042 4144 1076
rect 4110 952 4144 986
rect 4110 862 4144 896
rect 4110 772 4144 806
rect 4110 682 4144 716
rect 4110 592 4144 626
rect 4110 502 4144 536
rect 4110 412 4144 446
rect 4110 322 4144 356
rect 4110 232 4144 266
rect 5297 1132 5331 1166
rect 5297 1042 5331 1076
rect 5297 952 5331 986
rect 5297 862 5331 896
rect 5297 772 5331 806
rect 5297 682 5331 716
rect 5297 592 5331 626
rect 5297 502 5331 536
rect 5297 412 5331 446
rect 5297 322 5331 356
rect 5297 232 5331 266
rect 4110 142 4144 176
rect 5297 142 5331 176
rect 4206 58 4240 92
rect 4296 58 4330 92
rect 4386 58 4420 92
rect 4476 58 4510 92
rect 4566 58 4600 92
rect 4656 58 4690 92
rect 4746 58 4780 92
rect 4836 58 4870 92
rect 4926 58 4960 92
rect 5016 58 5050 92
rect 5106 58 5140 92
rect 5196 58 5230 92
rect 5460 1222 5494 1256
rect 5556 1245 5590 1279
rect 5646 1245 5680 1279
rect 5736 1245 5770 1279
rect 5826 1245 5860 1279
rect 5916 1245 5950 1279
rect 6006 1245 6040 1279
rect 6096 1245 6130 1279
rect 6186 1245 6220 1279
rect 6276 1245 6310 1279
rect 6366 1245 6400 1279
rect 6456 1245 6490 1279
rect 6546 1245 6580 1279
rect 6647 1222 6681 1256
rect 5460 1132 5494 1166
rect 5460 1042 5494 1076
rect 5460 952 5494 986
rect 5460 862 5494 896
rect 5460 772 5494 806
rect 5460 682 5494 716
rect 5460 592 5494 626
rect 5460 502 5494 536
rect 5460 412 5494 446
rect 5460 322 5494 356
rect 5460 232 5494 266
rect 6647 1132 6681 1166
rect 6647 1042 6681 1076
rect 6647 952 6681 986
rect 6647 862 6681 896
rect 6647 772 6681 806
rect 6647 682 6681 716
rect 6647 592 6681 626
rect 6647 502 6681 536
rect 6647 412 6681 446
rect 6647 322 6681 356
rect 6647 232 6681 266
rect 5460 142 5494 176
rect 6647 142 6681 176
rect 5556 58 5590 92
rect 5646 58 5680 92
rect 5736 58 5770 92
rect 5826 58 5860 92
rect 5916 58 5950 92
rect 6006 58 6040 92
rect 6096 58 6130 92
rect 6186 58 6220 92
rect 6276 58 6310 92
rect 6366 58 6400 92
rect 6456 58 6490 92
rect 6546 58 6580 92
rect 6810 1222 6844 1256
rect 6906 1245 6940 1279
rect 6996 1245 7030 1279
rect 7086 1245 7120 1279
rect 7176 1245 7210 1279
rect 7266 1245 7300 1279
rect 7356 1245 7390 1279
rect 7446 1245 7480 1279
rect 7536 1245 7570 1279
rect 7626 1245 7660 1279
rect 7716 1245 7750 1279
rect 7806 1245 7840 1279
rect 7896 1245 7930 1279
rect 7997 1222 8031 1256
rect 6810 1132 6844 1166
rect 6810 1042 6844 1076
rect 6810 952 6844 986
rect 6810 862 6844 896
rect 6810 772 6844 806
rect 6810 682 6844 716
rect 6810 592 6844 626
rect 6810 502 6844 536
rect 6810 412 6844 446
rect 6810 322 6844 356
rect 6810 232 6844 266
rect 7997 1132 8031 1166
rect 7997 1042 8031 1076
rect 7997 952 8031 986
rect 7997 862 8031 896
rect 7997 772 8031 806
rect 7997 682 8031 716
rect 7997 592 8031 626
rect 7997 502 8031 536
rect 7997 412 8031 446
rect 7997 322 8031 356
rect 7997 232 8031 266
rect 6810 142 6844 176
rect 7997 142 8031 176
rect 6906 58 6940 92
rect 6996 58 7030 92
rect 7086 58 7120 92
rect 7176 58 7210 92
rect 7266 58 7300 92
rect 7356 58 7390 92
rect 7446 58 7480 92
rect 7536 58 7570 92
rect 7626 58 7660 92
rect 7716 58 7750 92
rect 7806 58 7840 92
rect 7896 58 7930 92
rect 8160 1222 8194 1256
rect 8256 1245 8290 1279
rect 8346 1245 8380 1279
rect 8436 1245 8470 1279
rect 8526 1245 8560 1279
rect 8616 1245 8650 1279
rect 8706 1245 8740 1279
rect 8796 1245 8830 1279
rect 8886 1245 8920 1279
rect 8976 1245 9010 1279
rect 9066 1245 9100 1279
rect 9156 1245 9190 1279
rect 9246 1245 9280 1279
rect 9347 1222 9381 1256
rect 8160 1132 8194 1166
rect 8160 1042 8194 1076
rect 8160 952 8194 986
rect 8160 862 8194 896
rect 8160 772 8194 806
rect 8160 682 8194 716
rect 8160 592 8194 626
rect 8160 502 8194 536
rect 8160 412 8194 446
rect 8160 322 8194 356
rect 8160 232 8194 266
rect 9347 1132 9381 1166
rect 9347 1042 9381 1076
rect 9347 952 9381 986
rect 9347 862 9381 896
rect 9347 772 9381 806
rect 9347 682 9381 716
rect 9347 592 9381 626
rect 9347 502 9381 536
rect 9347 412 9381 446
rect 9347 322 9381 356
rect 9347 232 9381 266
rect 8160 142 8194 176
rect 9347 142 9381 176
rect 8256 58 8290 92
rect 8346 58 8380 92
rect 8436 58 8470 92
rect 8526 58 8560 92
rect 8616 58 8650 92
rect 8706 58 8740 92
rect 8796 58 8830 92
rect 8886 58 8920 92
rect 8976 58 9010 92
rect 9066 58 9100 92
rect 9156 58 9190 92
rect 9246 58 9280 92
<< nsubdiffcont >>
rect 1670 1098 1704 1132
rect 1760 1098 1794 1132
rect 1850 1098 1884 1132
rect 1940 1098 1974 1132
rect 2030 1098 2064 1132
rect 2120 1098 2154 1132
rect 2210 1098 2244 1132
rect 2300 1098 2334 1132
rect 2390 1098 2424 1132
rect 1558 1041 1592 1075
rect 2448 1022 2482 1056
rect 1558 951 1592 985
rect 1558 861 1592 895
rect 1558 771 1592 805
rect 1558 681 1592 715
rect 1558 591 1592 625
rect 1558 501 1592 535
rect 1558 411 1592 445
rect 1558 321 1592 355
rect 2448 932 2482 966
rect 2448 842 2482 876
rect 2448 752 2482 786
rect 2448 662 2482 696
rect 2448 572 2482 606
rect 2448 482 2482 516
rect 2448 392 2482 426
rect 2448 302 2482 336
rect 1636 208 1670 242
rect 1726 208 1760 242
rect 1816 208 1850 242
rect 1906 208 1940 242
rect 1996 208 2030 242
rect 2086 208 2120 242
rect 2176 208 2210 242
rect 2266 208 2300 242
rect 2356 208 2390 242
rect 3020 1098 3054 1132
rect 3110 1098 3144 1132
rect 3200 1098 3234 1132
rect 3290 1098 3324 1132
rect 3380 1098 3414 1132
rect 3470 1098 3504 1132
rect 3560 1098 3594 1132
rect 3650 1098 3684 1132
rect 3740 1098 3774 1132
rect 2908 1041 2942 1075
rect 3798 1022 3832 1056
rect 2908 951 2942 985
rect 2908 861 2942 895
rect 2908 771 2942 805
rect 2908 681 2942 715
rect 2908 591 2942 625
rect 2908 501 2942 535
rect 2908 411 2942 445
rect 2908 321 2942 355
rect 3798 932 3832 966
rect 3798 842 3832 876
rect 3798 752 3832 786
rect 3798 662 3832 696
rect 3798 572 3832 606
rect 3798 482 3832 516
rect 3798 392 3832 426
rect 3798 302 3832 336
rect 2986 208 3020 242
rect 3076 208 3110 242
rect 3166 208 3200 242
rect 3256 208 3290 242
rect 3346 208 3380 242
rect 3436 208 3470 242
rect 3526 208 3560 242
rect 3616 208 3650 242
rect 3706 208 3740 242
rect 4370 1098 4404 1132
rect 4460 1098 4494 1132
rect 4550 1098 4584 1132
rect 4640 1098 4674 1132
rect 4730 1098 4764 1132
rect 4820 1098 4854 1132
rect 4910 1098 4944 1132
rect 5000 1098 5034 1132
rect 5090 1098 5124 1132
rect 4258 1041 4292 1075
rect 5148 1022 5182 1056
rect 4258 951 4292 985
rect 4258 861 4292 895
rect 4258 771 4292 805
rect 4258 681 4292 715
rect 4258 591 4292 625
rect 4258 501 4292 535
rect 4258 411 4292 445
rect 4258 321 4292 355
rect 5148 932 5182 966
rect 5148 842 5182 876
rect 5148 752 5182 786
rect 5148 662 5182 696
rect 5148 572 5182 606
rect 5148 482 5182 516
rect 5148 392 5182 426
rect 5148 302 5182 336
rect 4336 208 4370 242
rect 4426 208 4460 242
rect 4516 208 4550 242
rect 4606 208 4640 242
rect 4696 208 4730 242
rect 4786 208 4820 242
rect 4876 208 4910 242
rect 4966 208 5000 242
rect 5056 208 5090 242
rect 5720 1098 5754 1132
rect 5810 1098 5844 1132
rect 5900 1098 5934 1132
rect 5990 1098 6024 1132
rect 6080 1098 6114 1132
rect 6170 1098 6204 1132
rect 6260 1098 6294 1132
rect 6350 1098 6384 1132
rect 6440 1098 6474 1132
rect 5608 1041 5642 1075
rect 6498 1022 6532 1056
rect 5608 951 5642 985
rect 5608 861 5642 895
rect 5608 771 5642 805
rect 5608 681 5642 715
rect 5608 591 5642 625
rect 5608 501 5642 535
rect 5608 411 5642 445
rect 5608 321 5642 355
rect 6498 932 6532 966
rect 6498 842 6532 876
rect 6498 752 6532 786
rect 6498 662 6532 696
rect 6498 572 6532 606
rect 6498 482 6532 516
rect 6498 392 6532 426
rect 6498 302 6532 336
rect 5686 208 5720 242
rect 5776 208 5810 242
rect 5866 208 5900 242
rect 5956 208 5990 242
rect 6046 208 6080 242
rect 6136 208 6170 242
rect 6226 208 6260 242
rect 6316 208 6350 242
rect 6406 208 6440 242
rect 7070 1098 7104 1132
rect 7160 1098 7194 1132
rect 7250 1098 7284 1132
rect 7340 1098 7374 1132
rect 7430 1098 7464 1132
rect 7520 1098 7554 1132
rect 7610 1098 7644 1132
rect 7700 1098 7734 1132
rect 7790 1098 7824 1132
rect 6958 1041 6992 1075
rect 7848 1022 7882 1056
rect 6958 951 6992 985
rect 6958 861 6992 895
rect 6958 771 6992 805
rect 6958 681 6992 715
rect 6958 591 6992 625
rect 6958 501 6992 535
rect 6958 411 6992 445
rect 6958 321 6992 355
rect 7848 932 7882 966
rect 7848 842 7882 876
rect 7848 752 7882 786
rect 7848 662 7882 696
rect 7848 572 7882 606
rect 7848 482 7882 516
rect 7848 392 7882 426
rect 7848 302 7882 336
rect 7036 208 7070 242
rect 7126 208 7160 242
rect 7216 208 7250 242
rect 7306 208 7340 242
rect 7396 208 7430 242
rect 7486 208 7520 242
rect 7576 208 7610 242
rect 7666 208 7700 242
rect 7756 208 7790 242
rect 8420 1098 8454 1132
rect 8510 1098 8544 1132
rect 8600 1098 8634 1132
rect 8690 1098 8724 1132
rect 8780 1098 8814 1132
rect 8870 1098 8904 1132
rect 8960 1098 8994 1132
rect 9050 1098 9084 1132
rect 9140 1098 9174 1132
rect 8308 1041 8342 1075
rect 9198 1022 9232 1056
rect 8308 951 8342 985
rect 8308 861 8342 895
rect 8308 771 8342 805
rect 8308 681 8342 715
rect 8308 591 8342 625
rect 8308 501 8342 535
rect 8308 411 8342 445
rect 8308 321 8342 355
rect 9198 932 9232 966
rect 9198 842 9232 876
rect 9198 752 9232 786
rect 9198 662 9232 696
rect 9198 572 9232 606
rect 9198 482 9232 516
rect 9198 392 9232 426
rect 9198 302 9232 336
rect 8386 208 8420 242
rect 8476 208 8510 242
rect 8566 208 8600 242
rect 8656 208 8690 242
rect 8746 208 8780 242
rect 8836 208 8870 242
rect 8926 208 8960 242
rect 9016 208 9050 242
rect 9106 208 9140 242
<< poly >>
rect 5390 4860 5510 4890
rect 5610 4860 5730 4890
rect 5830 4860 5950 4890
rect 6050 4860 6170 4890
rect 6270 4860 6390 4890
rect 6490 4880 6830 4910
rect 6490 4860 6610 4880
rect 6710 4860 6830 4880
rect 6930 4860 7050 4890
rect 7150 4860 7270 4890
rect 7370 4860 7490 4890
rect 7590 4860 7710 4890
rect 7810 4860 7930 4890
rect 1970 4760 2090 4790
rect 2190 4760 2310 4790
rect 2410 4760 2530 4790
rect 2630 4760 2750 4790
rect 2850 4760 2970 4790
rect 3070 4760 3190 4790
rect 3290 4760 3410 4790
rect 3510 4760 3630 4790
rect 3730 4760 3850 4790
rect 3950 4760 4070 4790
rect 4170 4760 4290 4790
rect 4390 4760 4510 4790
rect -1610 4360 -1580 4390
rect -1310 4360 -1280 4390
rect 5390 4440 5510 4460
rect 5610 4440 5730 4460
rect 5830 4440 5950 4460
rect 6050 4440 6170 4460
rect 6270 4440 6390 4460
rect 5390 4410 6390 4440
rect 6490 4430 6610 4460
rect 6710 4430 6830 4460
rect 6930 4440 7050 4460
rect 7150 4440 7270 4460
rect 7370 4440 7490 4460
rect 7590 4440 7710 4460
rect 7810 4440 7930 4460
rect 6930 4410 7930 4440
rect 5960 4370 5980 4410
rect 6020 4370 6040 4410
rect 5960 4350 6040 4370
rect 7280 4370 7300 4410
rect 7340 4370 7360 4410
rect 7280 4350 7360 4370
rect 6290 4000 6370 4020
rect 6290 3960 6310 4000
rect 6350 3960 6370 4000
rect 6950 4000 7030 4020
rect 6950 3960 6970 4000
rect 7010 3960 7030 4000
rect -1610 3930 -1580 3960
rect -1310 3930 -1280 3960
rect 1970 3930 2090 3960
rect 2190 3930 2310 3960
rect 2410 3930 2530 3960
rect 2630 3930 2750 3960
rect 2850 3930 2970 3960
rect 3070 3930 3190 3960
rect 3290 3930 3410 3960
rect 3510 3930 3630 3960
rect 3730 3930 3850 3960
rect 3950 3930 4070 3960
rect 4170 3930 4290 3960
rect 4390 3930 4510 3960
rect 5830 3910 5950 3940
rect 6050 3910 6170 3940
rect 6270 3930 7050 3960
rect 6270 3910 6390 3930
rect 6490 3910 6610 3930
rect 6710 3910 6830 3930
rect 6930 3910 7050 3930
rect 7150 3910 7270 3940
rect 7370 3910 7490 3940
rect 5830 3690 5950 3710
rect 6050 3690 6170 3710
rect -2710 3660 -710 3690
rect 5830 3660 6170 3690
rect 6270 3680 6390 3710
rect 6490 3680 6610 3710
rect 6710 3680 6830 3710
rect 6930 3680 7050 3710
rect 7150 3690 7270 3710
rect 7370 3690 7490 3710
rect 7150 3660 7490 3690
rect -2710 3430 -710 3460
rect 5810 3450 6610 3470
rect 5810 3410 5830 3450
rect 5870 3410 5910 3450
rect 5950 3410 5990 3450
rect 6030 3410 6070 3450
rect 6110 3410 6150 3450
rect 6190 3410 6230 3450
rect 6270 3410 6310 3450
rect 6350 3410 6390 3450
rect 6430 3410 6470 3450
rect 6510 3410 6550 3450
rect 6590 3410 6610 3450
rect 5810 3360 6610 3410
rect 6710 3450 7510 3470
rect 6710 3410 6730 3450
rect 6770 3410 6810 3450
rect 6850 3410 6890 3450
rect 6930 3410 6970 3450
rect 7010 3410 7050 3450
rect 7090 3410 7130 3450
rect 7170 3410 7210 3450
rect 7250 3410 7290 3450
rect 7330 3410 7370 3450
rect 7410 3410 7450 3450
rect 7490 3410 7510 3450
rect 6710 3360 7510 3410
rect 5810 2530 6610 2560
rect 6710 2530 7510 2560
<< polycont >>
rect 5980 4370 6020 4410
rect 7300 4370 7340 4410
rect 6310 3960 6350 4000
rect 6970 3960 7010 4000
rect 5830 3410 5870 3450
rect 5910 3410 5950 3450
rect 5990 3410 6030 3450
rect 6070 3410 6110 3450
rect 6150 3410 6190 3450
rect 6230 3410 6270 3450
rect 6310 3410 6350 3450
rect 6390 3410 6430 3450
rect 6470 3410 6510 3450
rect 6550 3410 6590 3450
rect 6730 3410 6770 3450
rect 6810 3410 6850 3450
rect 6890 3410 6930 3450
rect 6970 3410 7010 3450
rect 7050 3410 7090 3450
rect 7130 3410 7170 3450
rect 7210 3410 7250 3450
rect 7290 3410 7330 3450
rect 7370 3410 7410 3450
rect 7450 3410 7490 3450
<< xpolycontact >>
rect 40 3170 110 3610
rect 40 1890 110 2330
rect 160 3170 230 3610
rect 160 1890 230 2330
rect 280 3170 350 3610
rect 280 1890 350 2330
rect 400 3170 470 3610
rect 400 1890 470 2330
rect 520 3170 590 3610
rect 520 1890 590 2330
rect 640 3170 710 3610
rect 640 1890 710 2330
rect 760 3170 830 3610
rect 760 1890 830 2330
rect 880 3170 950 3610
rect 880 1890 950 2330
rect 1240 3170 1310 3610
rect 1240 1890 1310 2330
rect 1360 3170 1430 3610
rect 1360 1890 1430 2330
rect 1480 3170 1550 3610
rect 1480 1890 1550 2330
rect 1600 3170 1670 3610
rect 1600 1890 1670 2330
rect 1720 3170 1790 3610
rect 1720 1890 1790 2330
rect 1840 3170 1910 3610
rect 1840 1890 1910 2330
rect 1960 3170 2030 3610
rect 1960 1890 2030 2330
rect 2080 3170 2150 3610
rect 2080 1890 2150 2330
rect 2440 3170 2510 3610
rect 2440 1890 2510 2330
rect 2560 3170 2630 3610
rect 2560 1890 2630 2330
rect 2680 3170 2750 3610
rect 2680 1890 2750 2330
rect 2800 3170 2870 3610
rect 2800 1890 2870 2330
rect 2920 3170 2990 3610
rect 2920 1890 2990 2330
rect 3040 3170 3110 3610
rect 3040 1890 3110 2330
rect 3160 3170 3230 3610
rect 3160 1890 3230 2330
rect 3280 3170 3350 3610
rect 3280 1890 3350 2330
rect 4280 3030 4350 3470
rect 4280 1890 4350 2330
<< xpolyres >>
rect 40 2330 110 3170
rect 160 2330 230 3170
rect 280 2330 350 3170
rect 400 2330 470 3170
rect 520 2330 590 3170
rect 640 2330 710 3170
rect 760 2330 830 3170
rect 880 2330 950 3170
rect 1240 2330 1310 3170
rect 1360 2330 1430 3170
rect 1480 2330 1550 3170
rect 1600 2330 1670 3170
rect 1720 2330 1790 3170
rect 1840 2330 1910 3170
rect 1960 2330 2030 3170
rect 2080 2330 2150 3170
rect 2440 2330 2510 3170
rect 2560 2330 2630 3170
rect 2680 2330 2750 3170
rect 2800 2330 2870 3170
rect 2920 2330 2990 3170
rect 3040 2330 3110 3170
rect 3160 2330 3230 3170
rect 3280 2330 3350 3170
rect 4280 2330 4350 3030
<< locali >>
rect 5300 4950 5380 4970
rect 5300 4910 5320 4950
rect 5360 4910 5380 4950
rect 5300 4890 5380 4910
rect 5740 4950 5820 4970
rect 5740 4910 5760 4950
rect 5800 4910 5820 4950
rect 5740 4890 5820 4910
rect 6180 4950 6260 4970
rect 6180 4910 6200 4950
rect 6240 4910 6260 4950
rect 6180 4890 6260 4910
rect 6620 4950 6700 4970
rect 6620 4910 6640 4950
rect 6680 4910 6700 4950
rect 6620 4890 6700 4910
rect 7060 4950 7140 4970
rect 7060 4910 7080 4950
rect 7120 4910 7140 4950
rect 7060 4890 7140 4910
rect 7500 4950 7580 4970
rect 7500 4910 7520 4950
rect 7560 4910 7580 4950
rect 7500 4890 7580 4910
rect 7940 4950 8020 4970
rect 7940 4910 7960 4950
rect 8000 4910 8020 4950
rect 7940 4890 8020 4910
rect 5320 4850 5360 4890
rect 5760 4850 5800 4890
rect 6200 4850 6240 4890
rect 6640 4850 6680 4890
rect 7080 4850 7120 4890
rect 7520 4850 7560 4890
rect 7960 4850 8000 4890
rect 5300 4830 5380 4850
rect 1900 4790 4580 4830
rect 1900 4750 1940 4790
rect 4540 4750 4580 4790
rect 5300 4790 5320 4830
rect 5360 4790 5380 4830
rect 1880 4730 1960 4750
rect -1700 4330 -1620 4350
rect -1700 3990 -1680 4330
rect -1640 3990 -1620 4330
rect -1700 3970 -1620 3990
rect -1570 4330 -1490 4350
rect -1570 3990 -1550 4330
rect -1510 3990 -1490 4330
rect -1570 3970 -1490 3990
rect -1400 4330 -1320 4350
rect -1400 3990 -1380 4330
rect -1340 3990 -1320 4330
rect -1400 3970 -1320 3990
rect -1270 4330 -1190 4350
rect -1270 3990 -1250 4330
rect -1210 3990 -1190 4330
rect -1270 3970 -1190 3990
rect 1880 3990 1900 4730
rect 1940 3990 1960 4730
rect 1880 3970 1960 3990
rect 2100 4730 2180 4750
rect 2100 3990 2120 4730
rect 2160 3990 2180 4730
rect 2100 3970 2180 3990
rect 2320 4730 2400 4750
rect 2320 3990 2340 4730
rect 2380 3990 2400 4730
rect 2320 3970 2400 3990
rect 2540 4730 2620 4750
rect 2540 3990 2560 4730
rect 2600 3990 2620 4730
rect 2540 3970 2620 3990
rect 2760 4730 2840 4750
rect 2760 3990 2780 4730
rect 2820 3990 2840 4730
rect 2760 3970 2840 3990
rect 2980 4730 3060 4750
rect 2980 3990 3000 4730
rect 3040 3990 3060 4730
rect 2980 3970 3060 3990
rect 3200 4730 3280 4750
rect 3200 3990 3220 4730
rect 3260 3990 3280 4730
rect 3200 3970 3280 3990
rect 3420 4730 3500 4750
rect 3420 3990 3440 4730
rect 3480 3990 3500 4730
rect 3420 3970 3500 3990
rect 3640 4730 3720 4750
rect 3640 3990 3660 4730
rect 3700 3990 3720 4730
rect 3640 3970 3720 3990
rect 3860 4730 3940 4750
rect 3860 3990 3880 4730
rect 3920 3990 3940 4730
rect 3860 3970 3940 3990
rect 4080 4730 4160 4750
rect 4080 3990 4100 4730
rect 4140 3990 4160 4730
rect 4080 3970 4160 3990
rect 4300 4730 4380 4750
rect 4300 3990 4320 4730
rect 4360 3990 4380 4730
rect 4300 3970 4380 3990
rect 4520 4730 4600 4750
rect 4520 3990 4540 4730
rect 4580 3990 4600 4730
rect 5300 4730 5380 4790
rect 5300 4690 5320 4730
rect 5360 4690 5380 4730
rect 5300 4630 5380 4690
rect 5300 4590 5320 4630
rect 5360 4590 5380 4630
rect 5300 4530 5380 4590
rect 5300 4490 5320 4530
rect 5360 4490 5380 4530
rect 5300 4470 5380 4490
rect 5520 4830 5600 4850
rect 5520 4790 5540 4830
rect 5580 4790 5600 4830
rect 5520 4730 5600 4790
rect 5520 4690 5540 4730
rect 5580 4690 5600 4730
rect 5520 4630 5600 4690
rect 5520 4590 5540 4630
rect 5580 4590 5600 4630
rect 5520 4530 5600 4590
rect 5520 4490 5540 4530
rect 5580 4490 5600 4530
rect 5520 4470 5600 4490
rect 5740 4830 5820 4850
rect 5740 4790 5760 4830
rect 5800 4790 5820 4830
rect 5740 4730 5820 4790
rect 5740 4690 5760 4730
rect 5800 4690 5820 4730
rect 5740 4630 5820 4690
rect 5740 4590 5760 4630
rect 5800 4590 5820 4630
rect 5740 4530 5820 4590
rect 5740 4490 5760 4530
rect 5800 4490 5820 4530
rect 5740 4470 5820 4490
rect 5960 4830 6040 4850
rect 5960 4790 5980 4830
rect 6020 4790 6040 4830
rect 5960 4730 6040 4790
rect 5960 4690 5980 4730
rect 6020 4690 6040 4730
rect 5960 4630 6040 4690
rect 5960 4590 5980 4630
rect 6020 4590 6040 4630
rect 5960 4530 6040 4590
rect 5960 4490 5980 4530
rect 6020 4490 6040 4530
rect 5960 4470 6040 4490
rect 6180 4830 6260 4850
rect 6180 4790 6200 4830
rect 6240 4790 6260 4830
rect 6180 4730 6260 4790
rect 6180 4690 6200 4730
rect 6240 4690 6260 4730
rect 6180 4630 6260 4690
rect 6180 4590 6200 4630
rect 6240 4590 6260 4630
rect 6180 4530 6260 4590
rect 6180 4490 6200 4530
rect 6240 4490 6260 4530
rect 6180 4470 6260 4490
rect 6400 4830 6480 4850
rect 6400 4790 6420 4830
rect 6460 4790 6480 4830
rect 6400 4730 6480 4790
rect 6400 4690 6420 4730
rect 6460 4690 6480 4730
rect 6400 4630 6480 4690
rect 6400 4590 6420 4630
rect 6460 4590 6480 4630
rect 6400 4530 6480 4590
rect 6400 4490 6420 4530
rect 6460 4490 6480 4530
rect 6400 4470 6480 4490
rect 6620 4830 6700 4850
rect 6620 4790 6640 4830
rect 6680 4790 6700 4830
rect 6620 4730 6700 4790
rect 6620 4690 6640 4730
rect 6680 4690 6700 4730
rect 6620 4630 6700 4690
rect 6620 4590 6640 4630
rect 6680 4590 6700 4630
rect 6620 4530 6700 4590
rect 6620 4490 6640 4530
rect 6680 4490 6700 4530
rect 6620 4470 6700 4490
rect 6840 4830 6920 4850
rect 6840 4790 6860 4830
rect 6900 4790 6920 4830
rect 6840 4730 6920 4790
rect 6840 4690 6860 4730
rect 6900 4690 6920 4730
rect 6840 4630 6920 4690
rect 6840 4590 6860 4630
rect 6900 4590 6920 4630
rect 6840 4530 6920 4590
rect 6840 4490 6860 4530
rect 6900 4490 6920 4530
rect 6840 4470 6920 4490
rect 7060 4830 7140 4850
rect 7060 4790 7080 4830
rect 7120 4790 7140 4830
rect 7060 4730 7140 4790
rect 7060 4690 7080 4730
rect 7120 4690 7140 4730
rect 7060 4630 7140 4690
rect 7060 4590 7080 4630
rect 7120 4590 7140 4630
rect 7060 4530 7140 4590
rect 7060 4490 7080 4530
rect 7120 4490 7140 4530
rect 7060 4470 7140 4490
rect 7280 4830 7360 4850
rect 7280 4790 7300 4830
rect 7340 4790 7360 4830
rect 7280 4730 7360 4790
rect 7280 4690 7300 4730
rect 7340 4690 7360 4730
rect 7280 4630 7360 4690
rect 7280 4590 7300 4630
rect 7340 4590 7360 4630
rect 7280 4530 7360 4590
rect 7280 4490 7300 4530
rect 7340 4490 7360 4530
rect 7280 4470 7360 4490
rect 7500 4830 7580 4850
rect 7500 4790 7520 4830
rect 7560 4790 7580 4830
rect 7500 4730 7580 4790
rect 7500 4690 7520 4730
rect 7560 4690 7580 4730
rect 7500 4630 7580 4690
rect 7500 4590 7520 4630
rect 7560 4590 7580 4630
rect 7500 4530 7580 4590
rect 7500 4490 7520 4530
rect 7560 4490 7580 4530
rect 7500 4470 7580 4490
rect 7720 4830 7800 4850
rect 7720 4790 7740 4830
rect 7780 4790 7800 4830
rect 7720 4730 7800 4790
rect 7720 4690 7740 4730
rect 7780 4690 7800 4730
rect 7720 4630 7800 4690
rect 7720 4590 7740 4630
rect 7780 4590 7800 4630
rect 7720 4530 7800 4590
rect 7720 4490 7740 4530
rect 7780 4490 7800 4530
rect 7720 4470 7800 4490
rect 7940 4830 8020 4850
rect 7940 4790 7960 4830
rect 8000 4790 8020 4830
rect 7940 4730 8020 4790
rect 7940 4690 7960 4730
rect 8000 4690 8020 4730
rect 7940 4630 8020 4690
rect 7940 4590 7960 4630
rect 8000 4590 8020 4630
rect 7940 4530 8020 4590
rect 7940 4490 7960 4530
rect 8000 4490 8020 4530
rect 7940 4470 8020 4490
rect 5540 4230 5580 4470
rect 5980 4430 6020 4470
rect 6420 4430 6460 4470
rect 6860 4430 6900 4470
rect 7300 4430 7340 4470
rect 5960 4410 6040 4430
rect 5960 4370 5980 4410
rect 6020 4370 6040 4410
rect 6420 4390 6900 4430
rect 7280 4410 7360 4430
rect 5960 4350 6040 4370
rect 6640 4340 6680 4390
rect 7280 4370 7300 4410
rect 7340 4370 7360 4410
rect 7280 4350 7360 4370
rect 6620 4320 6700 4340
rect 6620 4280 6640 4320
rect 6680 4280 6700 4320
rect 6620 4260 6700 4280
rect 7620 4320 7700 4340
rect 7620 4280 7640 4320
rect 7680 4280 7700 4320
rect 7620 4260 7700 4280
rect 7740 4230 7780 4470
rect 5520 4210 5600 4230
rect 5520 4170 5540 4210
rect 5580 4170 5600 4210
rect 5520 4150 5600 4170
rect 6620 4200 6700 4220
rect 6620 4160 6640 4200
rect 6680 4160 6700 4200
rect 6620 4140 6700 4160
rect 7720 4210 7800 4230
rect 7720 4170 7740 4210
rect 7780 4170 7800 4210
rect 7720 4150 7800 4170
rect 5960 4100 6040 4120
rect 5960 4060 5980 4100
rect 6020 4060 6040 4100
rect 5960 4040 6040 4060
rect 7280 4100 7360 4120
rect 7280 4060 7300 4100
rect 7340 4060 7360 4100
rect 7280 4040 7360 4060
rect 4520 3970 4600 3990
rect 5980 3900 6020 4040
rect 6290 4000 6370 4020
rect 6290 3960 6310 4000
rect 6350 3960 6370 4000
rect 6620 4000 6700 4020
rect 6620 3980 6640 4000
rect 6290 3940 6370 3960
rect 6420 3960 6640 3980
rect 6680 3980 6700 4000
rect 6950 4000 7030 4020
rect 6680 3960 6900 3980
rect 6420 3940 6900 3960
rect 6950 3960 6970 4000
rect 7010 3960 7030 4000
rect 6950 3940 7030 3960
rect 6420 3900 6460 3940
rect 6860 3900 6900 3940
rect 7300 3900 7340 4040
rect 5740 3880 5820 3900
rect 5740 3840 5760 3880
rect 5800 3840 5820 3880
rect 5740 3780 5820 3840
rect 5740 3740 5760 3780
rect 5800 3740 5820 3780
rect 5740 3720 5820 3740
rect 5960 3880 6040 3900
rect 5960 3840 5980 3880
rect 6020 3840 6040 3880
rect 5960 3780 6040 3840
rect 5960 3740 5980 3780
rect 6020 3740 6040 3780
rect 5960 3720 6040 3740
rect 6180 3880 6260 3900
rect 6180 3840 6200 3880
rect 6240 3840 6260 3880
rect 6180 3780 6260 3840
rect 6180 3740 6200 3780
rect 6240 3740 6260 3780
rect 6180 3720 6260 3740
rect 6400 3880 6480 3900
rect 6400 3840 6420 3880
rect 6460 3840 6480 3880
rect 6400 3780 6480 3840
rect 6400 3740 6420 3780
rect 6460 3740 6480 3780
rect 6400 3720 6480 3740
rect 6620 3880 6700 3900
rect 6620 3840 6640 3880
rect 6680 3840 6700 3880
rect 6620 3780 6700 3840
rect 6620 3740 6640 3780
rect 6680 3740 6700 3780
rect 6620 3720 6700 3740
rect 6840 3880 6920 3900
rect 6840 3840 6860 3880
rect 6900 3840 6920 3880
rect 6840 3780 6920 3840
rect 6840 3740 6860 3780
rect 6900 3740 6920 3780
rect 6840 3720 6920 3740
rect 7060 3880 7140 3900
rect 7060 3840 7080 3880
rect 7120 3840 7140 3880
rect 7060 3780 7140 3840
rect 7060 3740 7080 3780
rect 7120 3740 7140 3780
rect 7060 3720 7140 3740
rect 7280 3880 7360 3900
rect 7280 3840 7300 3880
rect 7340 3840 7360 3880
rect 7280 3780 7360 3840
rect 7280 3740 7300 3780
rect 7340 3740 7360 3780
rect 7280 3720 7360 3740
rect 7500 3880 7580 3900
rect 7500 3840 7520 3880
rect 7560 3840 7580 3880
rect 7500 3780 7580 3840
rect 7500 3740 7520 3780
rect 7560 3740 7580 3780
rect 7500 3720 7580 3740
rect -2800 3630 -2720 3650
rect -2800 3490 -2780 3630
rect -2740 3490 -2720 3630
rect -2800 3470 -2720 3490
rect -700 3630 -620 3650
rect -700 3490 -680 3630
rect -640 3490 -620 3630
rect -700 3470 -620 3490
rect 110 3170 160 3610
rect 350 3170 400 3610
rect 590 3170 640 3610
rect 830 3170 880 3610
rect 1310 3170 1360 3610
rect 1550 3170 1600 3610
rect 1790 3170 1840 3610
rect 2030 3170 2080 3610
rect 2510 3170 2560 3610
rect 2750 3170 2800 3610
rect 2990 3170 3040 3610
rect 3230 3170 3280 3610
rect 5760 3590 5800 3720
rect 5960 3660 6040 3680
rect 5960 3620 5980 3660
rect 6020 3620 6040 3660
rect 5960 3600 6040 3620
rect 6200 3590 6240 3720
rect 6640 3590 6680 3720
rect 7080 3590 7120 3720
rect 7280 3660 7360 3680
rect 7280 3620 7300 3660
rect 7340 3620 7360 3660
rect 7280 3600 7360 3620
rect 7520 3590 7560 3720
rect 5740 3570 5820 3590
rect 5740 3530 5760 3570
rect 5800 3530 5820 3570
rect 5740 3510 5820 3530
rect 6180 3570 6260 3590
rect 6180 3530 6200 3570
rect 6240 3530 6260 3570
rect 6180 3510 6260 3530
rect 6620 3570 6700 3590
rect 6620 3530 6640 3570
rect 6680 3530 6700 3570
rect 6620 3510 6700 3530
rect 7060 3570 7140 3590
rect 7060 3530 7080 3570
rect 7120 3530 7140 3570
rect 7060 3510 7140 3530
rect 7500 3570 7580 3590
rect 7500 3530 7520 3570
rect 7560 3530 7580 3570
rect 7500 3510 7580 3530
rect 5740 3470 5780 3510
rect 5740 3450 6610 3470
rect 5740 3410 5830 3450
rect 5870 3410 5910 3450
rect 5950 3410 5990 3450
rect 6030 3410 6070 3450
rect 6110 3410 6150 3450
rect 6190 3410 6230 3450
rect 6270 3410 6310 3450
rect 6350 3410 6390 3450
rect 6430 3410 6470 3450
rect 6510 3410 6550 3450
rect 6590 3410 6610 3450
rect 5740 3390 6610 3410
rect 6710 3450 7580 3470
rect 6710 3410 6730 3450
rect 6770 3410 6810 3450
rect 6850 3410 6890 3450
rect 6930 3410 6970 3450
rect 7010 3410 7050 3450
rect 7090 3410 7130 3450
rect 7170 3410 7210 3450
rect 7250 3410 7290 3450
rect 7330 3410 7370 3450
rect 7410 3410 7450 3450
rect 7490 3410 7580 3450
rect 6710 3390 7580 3410
rect 5740 3350 5780 3390
rect 7540 3350 7580 3390
rect 5720 3330 5800 3350
rect 5720 3290 5740 3330
rect 5780 3290 5800 3330
rect 5720 3230 5800 3290
rect 5720 3190 5740 3230
rect 5780 3190 5800 3230
rect 5720 3130 5800 3190
rect 5720 3090 5740 3130
rect 5780 3090 5800 3130
rect 5720 3030 5800 3090
rect 5720 2990 5740 3030
rect 5780 2990 5800 3030
rect 5720 2930 5800 2990
rect 5720 2890 5740 2930
rect 5780 2890 5800 2930
rect 5720 2830 5800 2890
rect 5720 2790 5740 2830
rect 5780 2790 5800 2830
rect 5720 2730 5800 2790
rect 5720 2690 5740 2730
rect 5780 2690 5800 2730
rect 5720 2630 5800 2690
rect 5720 2590 5740 2630
rect 5780 2590 5800 2630
rect 5720 2570 5800 2590
rect 6620 3330 6700 3350
rect 6620 3290 6640 3330
rect 6680 3290 6700 3330
rect 6620 3230 6700 3290
rect 6620 3190 6640 3230
rect 6680 3190 6700 3230
rect 6620 3130 6700 3190
rect 6620 3090 6640 3130
rect 6680 3090 6700 3130
rect 6620 3030 6700 3090
rect 6620 2990 6640 3030
rect 6680 2990 6700 3030
rect 6620 2930 6700 2990
rect 6620 2890 6640 2930
rect 6680 2890 6700 2930
rect 6620 2830 6700 2890
rect 6620 2790 6640 2830
rect 6680 2790 6700 2830
rect 6620 2730 6700 2790
rect 6620 2690 6640 2730
rect 6680 2690 6700 2730
rect 6620 2630 6700 2690
rect 6620 2590 6640 2630
rect 6680 2590 6700 2630
rect 6620 2570 6700 2590
rect 7520 3330 7720 3350
rect 7520 3290 7540 3330
rect 7580 3310 7660 3330
rect 7580 3290 7600 3310
rect 7520 3230 7600 3290
rect 7640 3290 7660 3310
rect 7700 3290 7720 3330
rect 7640 3270 7720 3290
rect 7520 3190 7540 3230
rect 7580 3190 7600 3230
rect 7520 3130 7600 3190
rect 7520 3090 7540 3130
rect 7580 3090 7600 3130
rect 7520 3030 7600 3090
rect 7520 2990 7540 3030
rect 7580 2990 7600 3030
rect 7520 2930 7600 2990
rect 7520 2890 7540 2930
rect 7580 2890 7600 2930
rect 7520 2830 7600 2890
rect 7520 2790 7540 2830
rect 7580 2790 7600 2830
rect 7520 2730 7600 2790
rect 7520 2690 7540 2730
rect 7580 2690 7600 2730
rect 7520 2630 7600 2690
rect 7520 2590 7540 2630
rect 7580 2590 7600 2630
rect 7520 2570 7600 2590
rect 230 1890 280 2330
rect 470 1890 520 2330
rect 710 1890 760 2330
rect 1430 1890 1480 2330
rect 1670 1890 1720 2330
rect 1910 1890 1960 2330
rect 2630 1890 2680 2330
rect 2870 1890 2920 2330
rect 3110 1890 3160 2330
rect 20 1080 1320 1320
rect 20 270 270 1080
rect 1070 270 1320 1080
rect 20 20 1320 270
rect 1370 1279 9420 1320
rect 1370 1256 1506 1279
rect 1370 1222 1410 1256
rect 1444 1245 1506 1256
rect 1540 1245 1596 1279
rect 1630 1245 1686 1279
rect 1720 1245 1776 1279
rect 1810 1245 1866 1279
rect 1900 1245 1956 1279
rect 1990 1245 2046 1279
rect 2080 1245 2136 1279
rect 2170 1245 2226 1279
rect 2260 1245 2316 1279
rect 2350 1245 2406 1279
rect 2440 1245 2496 1279
rect 2530 1256 2856 1279
rect 2530 1245 2597 1256
rect 1444 1222 2597 1245
rect 2631 1222 2760 1256
rect 2794 1245 2856 1256
rect 2890 1245 2946 1279
rect 2980 1245 3036 1279
rect 3070 1245 3126 1279
rect 3160 1245 3216 1279
rect 3250 1245 3306 1279
rect 3340 1245 3396 1279
rect 3430 1245 3486 1279
rect 3520 1245 3576 1279
rect 3610 1245 3666 1279
rect 3700 1245 3756 1279
rect 3790 1245 3846 1279
rect 3880 1256 4206 1279
rect 3880 1245 3947 1256
rect 2794 1222 3947 1245
rect 3981 1222 4110 1256
rect 4144 1245 4206 1256
rect 4240 1245 4296 1279
rect 4330 1245 4386 1279
rect 4420 1245 4476 1279
rect 4510 1245 4566 1279
rect 4600 1245 4656 1279
rect 4690 1245 4746 1279
rect 4780 1245 4836 1279
rect 4870 1245 4926 1279
rect 4960 1245 5016 1279
rect 5050 1245 5106 1279
rect 5140 1245 5196 1279
rect 5230 1256 5556 1279
rect 5230 1245 5297 1256
rect 4144 1222 5297 1245
rect 5331 1222 5460 1256
rect 5494 1245 5556 1256
rect 5590 1245 5646 1279
rect 5680 1245 5736 1279
rect 5770 1245 5826 1279
rect 5860 1245 5916 1279
rect 5950 1245 6006 1279
rect 6040 1245 6096 1279
rect 6130 1245 6186 1279
rect 6220 1245 6276 1279
rect 6310 1245 6366 1279
rect 6400 1245 6456 1279
rect 6490 1245 6546 1279
rect 6580 1256 6906 1279
rect 6580 1245 6647 1256
rect 5494 1222 6647 1245
rect 6681 1222 6810 1256
rect 6844 1245 6906 1256
rect 6940 1245 6996 1279
rect 7030 1245 7086 1279
rect 7120 1245 7176 1279
rect 7210 1245 7266 1279
rect 7300 1245 7356 1279
rect 7390 1245 7446 1279
rect 7480 1245 7536 1279
rect 7570 1245 7626 1279
rect 7660 1245 7716 1279
rect 7750 1245 7806 1279
rect 7840 1245 7896 1279
rect 7930 1256 8256 1279
rect 7930 1245 7997 1256
rect 6844 1222 7997 1245
rect 8031 1222 8160 1256
rect 8194 1245 8256 1256
rect 8290 1245 8346 1279
rect 8380 1245 8436 1279
rect 8470 1245 8526 1279
rect 8560 1245 8616 1279
rect 8650 1245 8706 1279
rect 8740 1245 8796 1279
rect 8830 1245 8886 1279
rect 8920 1245 8976 1279
rect 9010 1245 9066 1279
rect 9100 1245 9156 1279
rect 9190 1245 9246 1279
rect 9280 1256 9420 1279
rect 9280 1245 9347 1256
rect 8194 1222 9347 1245
rect 9381 1222 9420 1256
rect 1370 1166 9420 1222
rect 1370 1132 1410 1166
rect 1444 1132 2597 1166
rect 2631 1132 2760 1166
rect 2794 1132 3947 1166
rect 3981 1132 4110 1166
rect 4144 1132 5297 1166
rect 5331 1132 5460 1166
rect 5494 1132 6647 1166
rect 6681 1132 6810 1166
rect 6844 1132 7997 1166
rect 8031 1132 8160 1166
rect 8194 1132 9347 1166
rect 9381 1132 9420 1166
rect 1370 1098 1670 1132
rect 1704 1098 1760 1132
rect 1794 1098 1850 1132
rect 1884 1098 1940 1132
rect 1974 1098 2030 1132
rect 2064 1098 2120 1132
rect 2154 1098 2210 1132
rect 2244 1098 2300 1132
rect 2334 1098 2390 1132
rect 2424 1098 3020 1132
rect 3054 1098 3110 1132
rect 3144 1098 3200 1132
rect 3234 1098 3290 1132
rect 3324 1098 3380 1132
rect 3414 1098 3470 1132
rect 3504 1098 3560 1132
rect 3594 1098 3650 1132
rect 3684 1098 3740 1132
rect 3774 1098 4370 1132
rect 4404 1098 4460 1132
rect 4494 1098 4550 1132
rect 4584 1098 4640 1132
rect 4674 1098 4730 1132
rect 4764 1098 4820 1132
rect 4854 1098 4910 1132
rect 4944 1098 5000 1132
rect 5034 1098 5090 1132
rect 5124 1098 5720 1132
rect 5754 1098 5810 1132
rect 5844 1098 5900 1132
rect 5934 1098 5990 1132
rect 6024 1098 6080 1132
rect 6114 1098 6170 1132
rect 6204 1098 6260 1132
rect 6294 1098 6350 1132
rect 6384 1098 6440 1132
rect 6474 1098 7070 1132
rect 7104 1098 7160 1132
rect 7194 1098 7250 1132
rect 7284 1098 7340 1132
rect 7374 1098 7430 1132
rect 7464 1098 7520 1132
rect 7554 1098 7610 1132
rect 7644 1098 7700 1132
rect 7734 1098 7790 1132
rect 7824 1098 8420 1132
rect 8454 1098 8510 1132
rect 8544 1098 8600 1132
rect 8634 1098 8690 1132
rect 8724 1098 8780 1132
rect 8814 1098 8870 1132
rect 8904 1098 8960 1132
rect 8994 1098 9050 1132
rect 9084 1098 9140 1132
rect 9174 1098 9420 1132
rect 1370 1079 9420 1098
rect 1370 1076 1620 1079
rect 1370 1042 1410 1076
rect 1444 1075 1620 1076
rect 1444 1042 1558 1075
rect 1370 1041 1558 1042
rect 1592 1041 1620 1075
rect 1370 986 1620 1041
rect 2420 1076 2970 1079
rect 2420 1056 2597 1076
rect 2420 1022 2448 1056
rect 2482 1042 2597 1056
rect 2631 1042 2760 1076
rect 2794 1075 2970 1076
rect 2794 1042 2908 1075
rect 2482 1041 2908 1042
rect 2942 1041 2970 1075
rect 2482 1022 2970 1041
rect 1370 952 1410 986
rect 1444 985 1620 986
rect 1444 952 1558 985
rect 1370 951 1558 952
rect 1592 951 1620 985
rect 1370 896 1620 951
rect 1370 862 1410 896
rect 1444 895 1620 896
rect 1444 862 1558 895
rect 1370 861 1558 862
rect 1592 861 1620 895
rect 1370 806 1620 861
rect 1370 772 1410 806
rect 1444 805 1620 806
rect 1444 772 1558 805
rect 1370 771 1558 772
rect 1592 771 1620 805
rect 1370 716 1620 771
rect 1370 682 1410 716
rect 1444 715 1620 716
rect 1444 682 1558 715
rect 1370 681 1558 682
rect 1592 681 1620 715
rect 1370 626 1620 681
rect 1370 592 1410 626
rect 1444 625 1620 626
rect 1444 592 1558 625
rect 1370 591 1558 592
rect 1592 591 1620 625
rect 1370 536 1620 591
rect 1370 502 1410 536
rect 1444 535 1620 536
rect 1444 502 1558 535
rect 1370 501 1558 502
rect 1592 501 1620 535
rect 1370 446 1620 501
rect 1370 412 1410 446
rect 1444 445 1620 446
rect 1444 412 1558 445
rect 1370 411 1558 412
rect 1592 411 1620 445
rect 1370 356 1620 411
rect 1370 322 1410 356
rect 1444 355 1620 356
rect 1444 322 1558 355
rect 1370 321 1558 322
rect 1592 321 1620 355
rect 1673 958 2367 1017
rect 1673 924 1734 958
rect 1768 930 1824 958
rect 1858 930 1914 958
rect 1948 930 2004 958
rect 1780 924 1824 930
rect 1880 924 1914 930
rect 1980 924 2004 930
rect 2038 930 2094 958
rect 2038 924 2046 930
rect 1673 896 1746 924
rect 1780 896 1846 924
rect 1880 896 1946 924
rect 1980 896 2046 924
rect 2080 924 2094 930
rect 2128 930 2184 958
rect 2128 924 2146 930
rect 2080 896 2146 924
rect 2180 924 2184 930
rect 2218 930 2274 958
rect 2218 924 2246 930
rect 2308 924 2367 958
rect 2180 896 2246 924
rect 2280 896 2367 924
rect 1673 868 2367 896
rect 1673 834 1734 868
rect 1768 834 1824 868
rect 1858 834 1914 868
rect 1948 834 2004 868
rect 2038 834 2094 868
rect 2128 834 2184 868
rect 2218 834 2274 868
rect 2308 834 2367 868
rect 1673 830 2367 834
rect 1673 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2367 830
rect 1673 778 2367 796
rect 1673 744 1734 778
rect 1768 744 1824 778
rect 1858 744 1914 778
rect 1948 744 2004 778
rect 2038 744 2094 778
rect 2128 744 2184 778
rect 2218 744 2274 778
rect 2308 744 2367 778
rect 1673 730 2367 744
rect 1673 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2367 730
rect 1673 688 2367 696
rect 1673 654 1734 688
rect 1768 654 1824 688
rect 1858 654 1914 688
rect 1948 654 2004 688
rect 2038 654 2094 688
rect 2128 654 2184 688
rect 2218 654 2274 688
rect 2308 654 2367 688
rect 1673 630 2367 654
rect 1673 598 1746 630
rect 1780 598 1846 630
rect 1880 598 1946 630
rect 1980 598 2046 630
rect 1673 564 1734 598
rect 1780 596 1824 598
rect 1880 596 1914 598
rect 1980 596 2004 598
rect 1768 564 1824 596
rect 1858 564 1914 596
rect 1948 564 2004 596
rect 2038 596 2046 598
rect 2080 598 2146 630
rect 2080 596 2094 598
rect 2038 564 2094 596
rect 2128 596 2146 598
rect 2180 598 2246 630
rect 2280 598 2367 630
rect 2180 596 2184 598
rect 2128 564 2184 596
rect 2218 596 2246 598
rect 2218 564 2274 596
rect 2308 564 2367 598
rect 1673 530 2367 564
rect 1673 508 1746 530
rect 1780 508 1846 530
rect 1880 508 1946 530
rect 1980 508 2046 530
rect 1673 474 1734 508
rect 1780 496 1824 508
rect 1880 496 1914 508
rect 1980 496 2004 508
rect 1768 474 1824 496
rect 1858 474 1914 496
rect 1948 474 2004 496
rect 2038 496 2046 508
rect 2080 508 2146 530
rect 2080 496 2094 508
rect 2038 474 2094 496
rect 2128 496 2146 508
rect 2180 508 2246 530
rect 2280 508 2367 530
rect 2180 496 2184 508
rect 2128 474 2184 496
rect 2218 496 2246 508
rect 2218 474 2274 496
rect 2308 474 2367 508
rect 1673 430 2367 474
rect 1673 418 1746 430
rect 1780 418 1846 430
rect 1880 418 1946 430
rect 1980 418 2046 430
rect 1673 384 1734 418
rect 1780 396 1824 418
rect 1880 396 1914 418
rect 1980 396 2004 418
rect 1768 384 1824 396
rect 1858 384 1914 396
rect 1948 384 2004 396
rect 2038 396 2046 418
rect 2080 418 2146 430
rect 2080 396 2094 418
rect 2038 384 2094 396
rect 2128 396 2146 418
rect 2180 418 2246 430
rect 2280 418 2367 430
rect 2180 396 2184 418
rect 2128 384 2184 396
rect 2218 396 2246 418
rect 2218 384 2274 396
rect 2308 384 2367 418
rect 1673 323 2367 384
rect 2420 986 2970 1022
rect 3770 1076 4320 1079
rect 3770 1056 3947 1076
rect 3770 1022 3798 1056
rect 3832 1042 3947 1056
rect 3981 1042 4110 1076
rect 4144 1075 4320 1076
rect 4144 1042 4258 1075
rect 3832 1041 4258 1042
rect 4292 1041 4320 1075
rect 3832 1022 4320 1041
rect 2420 966 2597 986
rect 2420 932 2448 966
rect 2482 952 2597 966
rect 2631 952 2760 986
rect 2794 985 2970 986
rect 2794 952 2908 985
rect 2482 951 2908 952
rect 2942 951 2970 985
rect 2482 932 2970 951
rect 2420 896 2970 932
rect 2420 876 2597 896
rect 2420 842 2448 876
rect 2482 862 2597 876
rect 2631 862 2760 896
rect 2794 895 2970 896
rect 2794 862 2908 895
rect 2482 861 2908 862
rect 2942 861 2970 895
rect 2482 842 2970 861
rect 2420 806 2970 842
rect 2420 786 2597 806
rect 2420 752 2448 786
rect 2482 772 2597 786
rect 2631 772 2760 806
rect 2794 805 2970 806
rect 2794 772 2908 805
rect 2482 771 2908 772
rect 2942 771 2970 805
rect 2482 752 2970 771
rect 2420 716 2970 752
rect 2420 696 2597 716
rect 2420 662 2448 696
rect 2482 682 2597 696
rect 2631 682 2760 716
rect 2794 715 2970 716
rect 2794 682 2908 715
rect 2482 681 2908 682
rect 2942 681 2970 715
rect 2482 662 2970 681
rect 2420 626 2970 662
rect 2420 606 2597 626
rect 2420 572 2448 606
rect 2482 592 2597 606
rect 2631 592 2760 626
rect 2794 625 2970 626
rect 2794 592 2908 625
rect 2482 591 2908 592
rect 2942 591 2970 625
rect 2482 572 2970 591
rect 2420 536 2970 572
rect 2420 516 2597 536
rect 2420 482 2448 516
rect 2482 502 2597 516
rect 2631 502 2760 536
rect 2794 535 2970 536
rect 2794 502 2908 535
rect 2482 501 2908 502
rect 2942 501 2970 535
rect 2482 482 2970 501
rect 2420 446 2970 482
rect 2420 426 2597 446
rect 2420 392 2448 426
rect 2482 412 2597 426
rect 2631 412 2760 446
rect 2794 445 2970 446
rect 2794 412 2908 445
rect 2482 411 2908 412
rect 2942 411 2970 445
rect 2482 392 2970 411
rect 2420 356 2970 392
rect 2420 336 2597 356
rect 1370 270 1620 321
rect 2420 302 2448 336
rect 2482 322 2597 336
rect 2631 322 2760 356
rect 2794 355 2970 356
rect 2794 322 2908 355
rect 2482 321 2908 322
rect 2942 321 2970 355
rect 3023 958 3717 1017
rect 3023 924 3084 958
rect 3118 930 3174 958
rect 3208 930 3264 958
rect 3298 930 3354 958
rect 3130 924 3174 930
rect 3230 924 3264 930
rect 3330 924 3354 930
rect 3388 930 3444 958
rect 3388 924 3396 930
rect 3023 896 3096 924
rect 3130 896 3196 924
rect 3230 896 3296 924
rect 3330 896 3396 924
rect 3430 924 3444 930
rect 3478 930 3534 958
rect 3478 924 3496 930
rect 3430 896 3496 924
rect 3530 924 3534 930
rect 3568 930 3624 958
rect 3568 924 3596 930
rect 3658 924 3717 958
rect 3530 896 3596 924
rect 3630 896 3717 924
rect 3023 868 3717 896
rect 3023 834 3084 868
rect 3118 834 3174 868
rect 3208 834 3264 868
rect 3298 834 3354 868
rect 3388 834 3444 868
rect 3478 834 3534 868
rect 3568 834 3624 868
rect 3658 834 3717 868
rect 3023 830 3717 834
rect 3023 796 3096 830
rect 3130 796 3196 830
rect 3230 796 3296 830
rect 3330 796 3396 830
rect 3430 796 3496 830
rect 3530 796 3596 830
rect 3630 796 3717 830
rect 3023 778 3717 796
rect 3023 744 3084 778
rect 3118 744 3174 778
rect 3208 744 3264 778
rect 3298 744 3354 778
rect 3388 744 3444 778
rect 3478 744 3534 778
rect 3568 744 3624 778
rect 3658 744 3717 778
rect 3023 730 3717 744
rect 3023 696 3096 730
rect 3130 696 3196 730
rect 3230 696 3296 730
rect 3330 696 3396 730
rect 3430 696 3496 730
rect 3530 696 3596 730
rect 3630 696 3717 730
rect 3023 688 3717 696
rect 3023 654 3084 688
rect 3118 654 3174 688
rect 3208 654 3264 688
rect 3298 654 3354 688
rect 3388 654 3444 688
rect 3478 654 3534 688
rect 3568 654 3624 688
rect 3658 654 3717 688
rect 3023 630 3717 654
rect 3023 598 3096 630
rect 3130 598 3196 630
rect 3230 598 3296 630
rect 3330 598 3396 630
rect 3023 564 3084 598
rect 3130 596 3174 598
rect 3230 596 3264 598
rect 3330 596 3354 598
rect 3118 564 3174 596
rect 3208 564 3264 596
rect 3298 564 3354 596
rect 3388 596 3396 598
rect 3430 598 3496 630
rect 3430 596 3444 598
rect 3388 564 3444 596
rect 3478 596 3496 598
rect 3530 598 3596 630
rect 3630 598 3717 630
rect 3530 596 3534 598
rect 3478 564 3534 596
rect 3568 596 3596 598
rect 3568 564 3624 596
rect 3658 564 3717 598
rect 3023 530 3717 564
rect 3023 508 3096 530
rect 3130 508 3196 530
rect 3230 508 3296 530
rect 3330 508 3396 530
rect 3023 474 3084 508
rect 3130 496 3174 508
rect 3230 496 3264 508
rect 3330 496 3354 508
rect 3118 474 3174 496
rect 3208 474 3264 496
rect 3298 474 3354 496
rect 3388 496 3396 508
rect 3430 508 3496 530
rect 3430 496 3444 508
rect 3388 474 3444 496
rect 3478 496 3496 508
rect 3530 508 3596 530
rect 3630 508 3717 530
rect 3530 496 3534 508
rect 3478 474 3534 496
rect 3568 496 3596 508
rect 3568 474 3624 496
rect 3658 474 3717 508
rect 3023 430 3717 474
rect 3023 418 3096 430
rect 3130 418 3196 430
rect 3230 418 3296 430
rect 3330 418 3396 430
rect 3023 384 3084 418
rect 3130 396 3174 418
rect 3230 396 3264 418
rect 3330 396 3354 418
rect 3118 384 3174 396
rect 3208 384 3264 396
rect 3298 384 3354 396
rect 3388 396 3396 418
rect 3430 418 3496 430
rect 3430 396 3444 418
rect 3388 384 3444 396
rect 3478 396 3496 418
rect 3530 418 3596 430
rect 3630 418 3717 430
rect 3530 396 3534 418
rect 3478 384 3534 396
rect 3568 396 3596 418
rect 3568 384 3624 396
rect 3658 384 3717 418
rect 3023 323 3717 384
rect 3770 986 4320 1022
rect 5120 1076 5670 1079
rect 5120 1056 5297 1076
rect 5120 1022 5148 1056
rect 5182 1042 5297 1056
rect 5331 1042 5460 1076
rect 5494 1075 5670 1076
rect 5494 1042 5608 1075
rect 5182 1041 5608 1042
rect 5642 1041 5670 1075
rect 5182 1022 5670 1041
rect 3770 966 3947 986
rect 3770 932 3798 966
rect 3832 952 3947 966
rect 3981 952 4110 986
rect 4144 985 4320 986
rect 4144 952 4258 985
rect 3832 951 4258 952
rect 4292 951 4320 985
rect 3832 932 4320 951
rect 3770 896 4320 932
rect 3770 876 3947 896
rect 3770 842 3798 876
rect 3832 862 3947 876
rect 3981 862 4110 896
rect 4144 895 4320 896
rect 4144 862 4258 895
rect 3832 861 4258 862
rect 4292 861 4320 895
rect 3832 842 4320 861
rect 3770 806 4320 842
rect 3770 786 3947 806
rect 3770 752 3798 786
rect 3832 772 3947 786
rect 3981 772 4110 806
rect 4144 805 4320 806
rect 4144 772 4258 805
rect 3832 771 4258 772
rect 4292 771 4320 805
rect 3832 752 4320 771
rect 3770 716 4320 752
rect 3770 696 3947 716
rect 3770 662 3798 696
rect 3832 682 3947 696
rect 3981 682 4110 716
rect 4144 715 4320 716
rect 4144 682 4258 715
rect 3832 681 4258 682
rect 4292 681 4320 715
rect 3832 662 4320 681
rect 3770 626 4320 662
rect 3770 606 3947 626
rect 3770 572 3798 606
rect 3832 592 3947 606
rect 3981 592 4110 626
rect 4144 625 4320 626
rect 4144 592 4258 625
rect 3832 591 4258 592
rect 4292 591 4320 625
rect 3832 572 4320 591
rect 3770 536 4320 572
rect 3770 516 3947 536
rect 3770 482 3798 516
rect 3832 502 3947 516
rect 3981 502 4110 536
rect 4144 535 4320 536
rect 4144 502 4258 535
rect 3832 501 4258 502
rect 4292 501 4320 535
rect 3832 482 4320 501
rect 3770 446 4320 482
rect 3770 426 3947 446
rect 3770 392 3798 426
rect 3832 412 3947 426
rect 3981 412 4110 446
rect 4144 445 4320 446
rect 4144 412 4258 445
rect 3832 411 4258 412
rect 4292 411 4320 445
rect 3832 392 4320 411
rect 3770 356 4320 392
rect 3770 336 3947 356
rect 2482 302 2970 321
rect 2420 270 2970 302
rect 3770 302 3798 336
rect 3832 322 3947 336
rect 3981 322 4110 356
rect 4144 355 4320 356
rect 4144 322 4258 355
rect 3832 321 4258 322
rect 4292 321 4320 355
rect 4373 958 5067 1017
rect 4373 924 4434 958
rect 4468 930 4524 958
rect 4558 930 4614 958
rect 4648 930 4704 958
rect 4480 924 4524 930
rect 4580 924 4614 930
rect 4680 924 4704 930
rect 4738 930 4794 958
rect 4738 924 4746 930
rect 4373 896 4446 924
rect 4480 896 4546 924
rect 4580 896 4646 924
rect 4680 896 4746 924
rect 4780 924 4794 930
rect 4828 930 4884 958
rect 4828 924 4846 930
rect 4780 896 4846 924
rect 4880 924 4884 930
rect 4918 930 4974 958
rect 4918 924 4946 930
rect 5008 924 5067 958
rect 4880 896 4946 924
rect 4980 896 5067 924
rect 4373 868 5067 896
rect 4373 834 4434 868
rect 4468 834 4524 868
rect 4558 834 4614 868
rect 4648 834 4704 868
rect 4738 834 4794 868
rect 4828 834 4884 868
rect 4918 834 4974 868
rect 5008 834 5067 868
rect 4373 830 5067 834
rect 4373 796 4446 830
rect 4480 796 4546 830
rect 4580 796 4646 830
rect 4680 796 4746 830
rect 4780 796 4846 830
rect 4880 796 4946 830
rect 4980 796 5067 830
rect 4373 778 5067 796
rect 4373 744 4434 778
rect 4468 744 4524 778
rect 4558 744 4614 778
rect 4648 744 4704 778
rect 4738 744 4794 778
rect 4828 744 4884 778
rect 4918 744 4974 778
rect 5008 744 5067 778
rect 4373 730 5067 744
rect 4373 696 4446 730
rect 4480 696 4546 730
rect 4580 696 4646 730
rect 4680 696 4746 730
rect 4780 696 4846 730
rect 4880 696 4946 730
rect 4980 696 5067 730
rect 4373 688 5067 696
rect 4373 654 4434 688
rect 4468 654 4524 688
rect 4558 654 4614 688
rect 4648 654 4704 688
rect 4738 654 4794 688
rect 4828 654 4884 688
rect 4918 654 4974 688
rect 5008 654 5067 688
rect 4373 630 5067 654
rect 4373 598 4446 630
rect 4480 598 4546 630
rect 4580 598 4646 630
rect 4680 598 4746 630
rect 4373 564 4434 598
rect 4480 596 4524 598
rect 4580 596 4614 598
rect 4680 596 4704 598
rect 4468 564 4524 596
rect 4558 564 4614 596
rect 4648 564 4704 596
rect 4738 596 4746 598
rect 4780 598 4846 630
rect 4780 596 4794 598
rect 4738 564 4794 596
rect 4828 596 4846 598
rect 4880 598 4946 630
rect 4980 598 5067 630
rect 4880 596 4884 598
rect 4828 564 4884 596
rect 4918 596 4946 598
rect 4918 564 4974 596
rect 5008 564 5067 598
rect 4373 530 5067 564
rect 4373 508 4446 530
rect 4480 508 4546 530
rect 4580 508 4646 530
rect 4680 508 4746 530
rect 4373 474 4434 508
rect 4480 496 4524 508
rect 4580 496 4614 508
rect 4680 496 4704 508
rect 4468 474 4524 496
rect 4558 474 4614 496
rect 4648 474 4704 496
rect 4738 496 4746 508
rect 4780 508 4846 530
rect 4780 496 4794 508
rect 4738 474 4794 496
rect 4828 496 4846 508
rect 4880 508 4946 530
rect 4980 508 5067 530
rect 4880 496 4884 508
rect 4828 474 4884 496
rect 4918 496 4946 508
rect 4918 474 4974 496
rect 5008 474 5067 508
rect 4373 430 5067 474
rect 4373 418 4446 430
rect 4480 418 4546 430
rect 4580 418 4646 430
rect 4680 418 4746 430
rect 4373 384 4434 418
rect 4480 396 4524 418
rect 4580 396 4614 418
rect 4680 396 4704 418
rect 4468 384 4524 396
rect 4558 384 4614 396
rect 4648 384 4704 396
rect 4738 396 4746 418
rect 4780 418 4846 430
rect 4780 396 4794 418
rect 4738 384 4794 396
rect 4828 396 4846 418
rect 4880 418 4946 430
rect 4980 418 5067 430
rect 4880 396 4884 418
rect 4828 384 4884 396
rect 4918 396 4946 418
rect 4918 384 4974 396
rect 5008 384 5067 418
rect 4373 323 5067 384
rect 5120 986 5670 1022
rect 6470 1076 7020 1079
rect 6470 1056 6647 1076
rect 6470 1022 6498 1056
rect 6532 1042 6647 1056
rect 6681 1042 6810 1076
rect 6844 1075 7020 1076
rect 6844 1042 6958 1075
rect 6532 1041 6958 1042
rect 6992 1041 7020 1075
rect 6532 1022 7020 1041
rect 5120 966 5297 986
rect 5120 932 5148 966
rect 5182 952 5297 966
rect 5331 952 5460 986
rect 5494 985 5670 986
rect 5494 952 5608 985
rect 5182 951 5608 952
rect 5642 951 5670 985
rect 5182 932 5670 951
rect 5120 896 5670 932
rect 5120 876 5297 896
rect 5120 842 5148 876
rect 5182 862 5297 876
rect 5331 862 5460 896
rect 5494 895 5670 896
rect 5494 862 5608 895
rect 5182 861 5608 862
rect 5642 861 5670 895
rect 5182 842 5670 861
rect 5120 806 5670 842
rect 5120 786 5297 806
rect 5120 752 5148 786
rect 5182 772 5297 786
rect 5331 772 5460 806
rect 5494 805 5670 806
rect 5494 772 5608 805
rect 5182 771 5608 772
rect 5642 771 5670 805
rect 5182 752 5670 771
rect 5120 716 5670 752
rect 5120 696 5297 716
rect 5120 662 5148 696
rect 5182 682 5297 696
rect 5331 682 5460 716
rect 5494 715 5670 716
rect 5494 682 5608 715
rect 5182 681 5608 682
rect 5642 681 5670 715
rect 5182 662 5670 681
rect 5120 626 5670 662
rect 5120 606 5297 626
rect 5120 572 5148 606
rect 5182 592 5297 606
rect 5331 592 5460 626
rect 5494 625 5670 626
rect 5494 592 5608 625
rect 5182 591 5608 592
rect 5642 591 5670 625
rect 5182 572 5670 591
rect 5120 536 5670 572
rect 5120 516 5297 536
rect 5120 482 5148 516
rect 5182 502 5297 516
rect 5331 502 5460 536
rect 5494 535 5670 536
rect 5494 502 5608 535
rect 5182 501 5608 502
rect 5642 501 5670 535
rect 5182 482 5670 501
rect 5120 446 5670 482
rect 5120 426 5297 446
rect 5120 392 5148 426
rect 5182 412 5297 426
rect 5331 412 5460 446
rect 5494 445 5670 446
rect 5494 412 5608 445
rect 5182 411 5608 412
rect 5642 411 5670 445
rect 5182 392 5670 411
rect 5120 356 5670 392
rect 5120 336 5297 356
rect 3832 302 4320 321
rect 3770 270 4320 302
rect 5120 302 5148 336
rect 5182 322 5297 336
rect 5331 322 5460 356
rect 5494 355 5670 356
rect 5494 322 5608 355
rect 5182 321 5608 322
rect 5642 321 5670 355
rect 5723 958 6417 1017
rect 5723 924 5784 958
rect 5818 930 5874 958
rect 5908 930 5964 958
rect 5998 930 6054 958
rect 5830 924 5874 930
rect 5930 924 5964 930
rect 6030 924 6054 930
rect 6088 930 6144 958
rect 6088 924 6096 930
rect 5723 896 5796 924
rect 5830 896 5896 924
rect 5930 896 5996 924
rect 6030 896 6096 924
rect 6130 924 6144 930
rect 6178 930 6234 958
rect 6178 924 6196 930
rect 6130 896 6196 924
rect 6230 924 6234 930
rect 6268 930 6324 958
rect 6268 924 6296 930
rect 6358 924 6417 958
rect 6230 896 6296 924
rect 6330 896 6417 924
rect 5723 868 6417 896
rect 5723 834 5784 868
rect 5818 834 5874 868
rect 5908 834 5964 868
rect 5998 834 6054 868
rect 6088 834 6144 868
rect 6178 834 6234 868
rect 6268 834 6324 868
rect 6358 834 6417 868
rect 5723 830 6417 834
rect 5723 796 5796 830
rect 5830 796 5896 830
rect 5930 796 5996 830
rect 6030 796 6096 830
rect 6130 796 6196 830
rect 6230 796 6296 830
rect 6330 796 6417 830
rect 5723 778 6417 796
rect 5723 744 5784 778
rect 5818 744 5874 778
rect 5908 744 5964 778
rect 5998 744 6054 778
rect 6088 744 6144 778
rect 6178 744 6234 778
rect 6268 744 6324 778
rect 6358 744 6417 778
rect 5723 730 6417 744
rect 5723 696 5796 730
rect 5830 696 5896 730
rect 5930 696 5996 730
rect 6030 696 6096 730
rect 6130 696 6196 730
rect 6230 696 6296 730
rect 6330 696 6417 730
rect 5723 688 6417 696
rect 5723 654 5784 688
rect 5818 654 5874 688
rect 5908 654 5964 688
rect 5998 654 6054 688
rect 6088 654 6144 688
rect 6178 654 6234 688
rect 6268 654 6324 688
rect 6358 654 6417 688
rect 5723 630 6417 654
rect 5723 598 5796 630
rect 5830 598 5896 630
rect 5930 598 5996 630
rect 6030 598 6096 630
rect 5723 564 5784 598
rect 5830 596 5874 598
rect 5930 596 5964 598
rect 6030 596 6054 598
rect 5818 564 5874 596
rect 5908 564 5964 596
rect 5998 564 6054 596
rect 6088 596 6096 598
rect 6130 598 6196 630
rect 6130 596 6144 598
rect 6088 564 6144 596
rect 6178 596 6196 598
rect 6230 598 6296 630
rect 6330 598 6417 630
rect 6230 596 6234 598
rect 6178 564 6234 596
rect 6268 596 6296 598
rect 6268 564 6324 596
rect 6358 564 6417 598
rect 5723 530 6417 564
rect 5723 508 5796 530
rect 5830 508 5896 530
rect 5930 508 5996 530
rect 6030 508 6096 530
rect 5723 474 5784 508
rect 5830 496 5874 508
rect 5930 496 5964 508
rect 6030 496 6054 508
rect 5818 474 5874 496
rect 5908 474 5964 496
rect 5998 474 6054 496
rect 6088 496 6096 508
rect 6130 508 6196 530
rect 6130 496 6144 508
rect 6088 474 6144 496
rect 6178 496 6196 508
rect 6230 508 6296 530
rect 6330 508 6417 530
rect 6230 496 6234 508
rect 6178 474 6234 496
rect 6268 496 6296 508
rect 6268 474 6324 496
rect 6358 474 6417 508
rect 5723 430 6417 474
rect 5723 418 5796 430
rect 5830 418 5896 430
rect 5930 418 5996 430
rect 6030 418 6096 430
rect 5723 384 5784 418
rect 5830 396 5874 418
rect 5930 396 5964 418
rect 6030 396 6054 418
rect 5818 384 5874 396
rect 5908 384 5964 396
rect 5998 384 6054 396
rect 6088 396 6096 418
rect 6130 418 6196 430
rect 6130 396 6144 418
rect 6088 384 6144 396
rect 6178 396 6196 418
rect 6230 418 6296 430
rect 6330 418 6417 430
rect 6230 396 6234 418
rect 6178 384 6234 396
rect 6268 396 6296 418
rect 6268 384 6324 396
rect 6358 384 6417 418
rect 5723 323 6417 384
rect 6470 986 7020 1022
rect 7820 1076 8370 1079
rect 7820 1056 7997 1076
rect 7820 1022 7848 1056
rect 7882 1042 7997 1056
rect 8031 1042 8160 1076
rect 8194 1075 8370 1076
rect 8194 1042 8308 1075
rect 7882 1041 8308 1042
rect 8342 1041 8370 1075
rect 7882 1022 8370 1041
rect 6470 966 6647 986
rect 6470 932 6498 966
rect 6532 952 6647 966
rect 6681 952 6810 986
rect 6844 985 7020 986
rect 6844 952 6958 985
rect 6532 951 6958 952
rect 6992 951 7020 985
rect 6532 932 7020 951
rect 6470 896 7020 932
rect 6470 876 6647 896
rect 6470 842 6498 876
rect 6532 862 6647 876
rect 6681 862 6810 896
rect 6844 895 7020 896
rect 6844 862 6958 895
rect 6532 861 6958 862
rect 6992 861 7020 895
rect 6532 842 7020 861
rect 6470 806 7020 842
rect 6470 786 6647 806
rect 6470 752 6498 786
rect 6532 772 6647 786
rect 6681 772 6810 806
rect 6844 805 7020 806
rect 6844 772 6958 805
rect 6532 771 6958 772
rect 6992 771 7020 805
rect 6532 752 7020 771
rect 6470 716 7020 752
rect 6470 696 6647 716
rect 6470 662 6498 696
rect 6532 682 6647 696
rect 6681 682 6810 716
rect 6844 715 7020 716
rect 6844 682 6958 715
rect 6532 681 6958 682
rect 6992 681 7020 715
rect 6532 662 7020 681
rect 6470 626 7020 662
rect 6470 606 6647 626
rect 6470 572 6498 606
rect 6532 592 6647 606
rect 6681 592 6810 626
rect 6844 625 7020 626
rect 6844 592 6958 625
rect 6532 591 6958 592
rect 6992 591 7020 625
rect 6532 572 7020 591
rect 6470 536 7020 572
rect 6470 516 6647 536
rect 6470 482 6498 516
rect 6532 502 6647 516
rect 6681 502 6810 536
rect 6844 535 7020 536
rect 6844 502 6958 535
rect 6532 501 6958 502
rect 6992 501 7020 535
rect 6532 482 7020 501
rect 6470 446 7020 482
rect 6470 426 6647 446
rect 6470 392 6498 426
rect 6532 412 6647 426
rect 6681 412 6810 446
rect 6844 445 7020 446
rect 6844 412 6958 445
rect 6532 411 6958 412
rect 6992 411 7020 445
rect 6532 392 7020 411
rect 6470 356 7020 392
rect 6470 336 6647 356
rect 5182 302 5670 321
rect 5120 270 5670 302
rect 6470 302 6498 336
rect 6532 322 6647 336
rect 6681 322 6810 356
rect 6844 355 7020 356
rect 6844 322 6958 355
rect 6532 321 6958 322
rect 6992 321 7020 355
rect 7073 958 7767 1017
rect 7073 924 7134 958
rect 7168 930 7224 958
rect 7258 930 7314 958
rect 7348 930 7404 958
rect 7180 924 7224 930
rect 7280 924 7314 930
rect 7380 924 7404 930
rect 7438 930 7494 958
rect 7438 924 7446 930
rect 7073 896 7146 924
rect 7180 896 7246 924
rect 7280 896 7346 924
rect 7380 896 7446 924
rect 7480 924 7494 930
rect 7528 930 7584 958
rect 7528 924 7546 930
rect 7480 896 7546 924
rect 7580 924 7584 930
rect 7618 930 7674 958
rect 7618 924 7646 930
rect 7708 924 7767 958
rect 7580 896 7646 924
rect 7680 896 7767 924
rect 7073 868 7767 896
rect 7073 834 7134 868
rect 7168 834 7224 868
rect 7258 834 7314 868
rect 7348 834 7404 868
rect 7438 834 7494 868
rect 7528 834 7584 868
rect 7618 834 7674 868
rect 7708 834 7767 868
rect 7073 830 7767 834
rect 7073 796 7146 830
rect 7180 796 7246 830
rect 7280 796 7346 830
rect 7380 796 7446 830
rect 7480 796 7546 830
rect 7580 796 7646 830
rect 7680 796 7767 830
rect 7073 778 7767 796
rect 7073 744 7134 778
rect 7168 744 7224 778
rect 7258 744 7314 778
rect 7348 744 7404 778
rect 7438 744 7494 778
rect 7528 744 7584 778
rect 7618 744 7674 778
rect 7708 744 7767 778
rect 7073 730 7767 744
rect 7073 696 7146 730
rect 7180 696 7246 730
rect 7280 696 7346 730
rect 7380 696 7446 730
rect 7480 696 7546 730
rect 7580 696 7646 730
rect 7680 696 7767 730
rect 7073 688 7767 696
rect 7073 654 7134 688
rect 7168 654 7224 688
rect 7258 654 7314 688
rect 7348 654 7404 688
rect 7438 654 7494 688
rect 7528 654 7584 688
rect 7618 654 7674 688
rect 7708 654 7767 688
rect 7073 630 7767 654
rect 7073 598 7146 630
rect 7180 598 7246 630
rect 7280 598 7346 630
rect 7380 598 7446 630
rect 7073 564 7134 598
rect 7180 596 7224 598
rect 7280 596 7314 598
rect 7380 596 7404 598
rect 7168 564 7224 596
rect 7258 564 7314 596
rect 7348 564 7404 596
rect 7438 596 7446 598
rect 7480 598 7546 630
rect 7480 596 7494 598
rect 7438 564 7494 596
rect 7528 596 7546 598
rect 7580 598 7646 630
rect 7680 598 7767 630
rect 7580 596 7584 598
rect 7528 564 7584 596
rect 7618 596 7646 598
rect 7618 564 7674 596
rect 7708 564 7767 598
rect 7073 530 7767 564
rect 7073 508 7146 530
rect 7180 508 7246 530
rect 7280 508 7346 530
rect 7380 508 7446 530
rect 7073 474 7134 508
rect 7180 496 7224 508
rect 7280 496 7314 508
rect 7380 496 7404 508
rect 7168 474 7224 496
rect 7258 474 7314 496
rect 7348 474 7404 496
rect 7438 496 7446 508
rect 7480 508 7546 530
rect 7480 496 7494 508
rect 7438 474 7494 496
rect 7528 496 7546 508
rect 7580 508 7646 530
rect 7680 508 7767 530
rect 7580 496 7584 508
rect 7528 474 7584 496
rect 7618 496 7646 508
rect 7618 474 7674 496
rect 7708 474 7767 508
rect 7073 430 7767 474
rect 7073 418 7146 430
rect 7180 418 7246 430
rect 7280 418 7346 430
rect 7380 418 7446 430
rect 7073 384 7134 418
rect 7180 396 7224 418
rect 7280 396 7314 418
rect 7380 396 7404 418
rect 7168 384 7224 396
rect 7258 384 7314 396
rect 7348 384 7404 396
rect 7438 396 7446 418
rect 7480 418 7546 430
rect 7480 396 7494 418
rect 7438 384 7494 396
rect 7528 396 7546 418
rect 7580 418 7646 430
rect 7680 418 7767 430
rect 7580 396 7584 418
rect 7528 384 7584 396
rect 7618 396 7646 418
rect 7618 384 7674 396
rect 7708 384 7767 418
rect 7073 323 7767 384
rect 7820 986 8370 1022
rect 9170 1076 9420 1079
rect 9170 1056 9347 1076
rect 9170 1022 9198 1056
rect 9232 1042 9347 1056
rect 9381 1042 9420 1076
rect 9232 1022 9420 1042
rect 7820 966 7997 986
rect 7820 932 7848 966
rect 7882 952 7997 966
rect 8031 952 8160 986
rect 8194 985 8370 986
rect 8194 952 8308 985
rect 7882 951 8308 952
rect 8342 951 8370 985
rect 7882 932 8370 951
rect 7820 896 8370 932
rect 7820 876 7997 896
rect 7820 842 7848 876
rect 7882 862 7997 876
rect 8031 862 8160 896
rect 8194 895 8370 896
rect 8194 862 8308 895
rect 7882 861 8308 862
rect 8342 861 8370 895
rect 7882 842 8370 861
rect 7820 806 8370 842
rect 7820 786 7997 806
rect 7820 752 7848 786
rect 7882 772 7997 786
rect 8031 772 8160 806
rect 8194 805 8370 806
rect 8194 772 8308 805
rect 7882 771 8308 772
rect 8342 771 8370 805
rect 7882 752 8370 771
rect 7820 716 8370 752
rect 7820 696 7997 716
rect 7820 662 7848 696
rect 7882 682 7997 696
rect 8031 682 8160 716
rect 8194 715 8370 716
rect 8194 682 8308 715
rect 7882 681 8308 682
rect 8342 681 8370 715
rect 7882 662 8370 681
rect 7820 626 8370 662
rect 7820 606 7997 626
rect 7820 572 7848 606
rect 7882 592 7997 606
rect 8031 592 8160 626
rect 8194 625 8370 626
rect 8194 592 8308 625
rect 7882 591 8308 592
rect 8342 591 8370 625
rect 7882 572 8370 591
rect 7820 536 8370 572
rect 7820 516 7997 536
rect 7820 482 7848 516
rect 7882 502 7997 516
rect 8031 502 8160 536
rect 8194 535 8370 536
rect 8194 502 8308 535
rect 7882 501 8308 502
rect 8342 501 8370 535
rect 7882 482 8370 501
rect 7820 446 8370 482
rect 7820 426 7997 446
rect 7820 392 7848 426
rect 7882 412 7997 426
rect 8031 412 8160 446
rect 8194 445 8370 446
rect 8194 412 8308 445
rect 7882 411 8308 412
rect 8342 411 8370 445
rect 7882 392 8370 411
rect 7820 356 8370 392
rect 7820 336 7997 356
rect 6532 302 7020 321
rect 6470 270 7020 302
rect 7820 302 7848 336
rect 7882 322 7997 336
rect 8031 322 8160 356
rect 8194 355 8370 356
rect 8194 322 8308 355
rect 7882 321 8308 322
rect 8342 321 8370 355
rect 8423 958 9117 1017
rect 8423 924 8484 958
rect 8518 930 8574 958
rect 8608 930 8664 958
rect 8698 930 8754 958
rect 8530 924 8574 930
rect 8630 924 8664 930
rect 8730 924 8754 930
rect 8788 930 8844 958
rect 8788 924 8796 930
rect 8423 896 8496 924
rect 8530 896 8596 924
rect 8630 896 8696 924
rect 8730 896 8796 924
rect 8830 924 8844 930
rect 8878 930 8934 958
rect 8878 924 8896 930
rect 8830 896 8896 924
rect 8930 924 8934 930
rect 8968 930 9024 958
rect 8968 924 8996 930
rect 9058 924 9117 958
rect 8930 896 8996 924
rect 9030 896 9117 924
rect 8423 868 9117 896
rect 8423 834 8484 868
rect 8518 834 8574 868
rect 8608 834 8664 868
rect 8698 834 8754 868
rect 8788 834 8844 868
rect 8878 834 8934 868
rect 8968 834 9024 868
rect 9058 834 9117 868
rect 8423 830 9117 834
rect 8423 796 8496 830
rect 8530 796 8596 830
rect 8630 796 8696 830
rect 8730 796 8796 830
rect 8830 796 8896 830
rect 8930 796 8996 830
rect 9030 796 9117 830
rect 8423 778 9117 796
rect 8423 744 8484 778
rect 8518 744 8574 778
rect 8608 744 8664 778
rect 8698 744 8754 778
rect 8788 744 8844 778
rect 8878 744 8934 778
rect 8968 744 9024 778
rect 9058 744 9117 778
rect 8423 730 9117 744
rect 8423 696 8496 730
rect 8530 696 8596 730
rect 8630 696 8696 730
rect 8730 696 8796 730
rect 8830 696 8896 730
rect 8930 696 8996 730
rect 9030 696 9117 730
rect 8423 688 9117 696
rect 8423 654 8484 688
rect 8518 654 8574 688
rect 8608 654 8664 688
rect 8698 654 8754 688
rect 8788 654 8844 688
rect 8878 654 8934 688
rect 8968 654 9024 688
rect 9058 654 9117 688
rect 8423 630 9117 654
rect 8423 598 8496 630
rect 8530 598 8596 630
rect 8630 598 8696 630
rect 8730 598 8796 630
rect 8423 564 8484 598
rect 8530 596 8574 598
rect 8630 596 8664 598
rect 8730 596 8754 598
rect 8518 564 8574 596
rect 8608 564 8664 596
rect 8698 564 8754 596
rect 8788 596 8796 598
rect 8830 598 8896 630
rect 8830 596 8844 598
rect 8788 564 8844 596
rect 8878 596 8896 598
rect 8930 598 8996 630
rect 9030 598 9117 630
rect 8930 596 8934 598
rect 8878 564 8934 596
rect 8968 596 8996 598
rect 8968 564 9024 596
rect 9058 564 9117 598
rect 8423 530 9117 564
rect 8423 508 8496 530
rect 8530 508 8596 530
rect 8630 508 8696 530
rect 8730 508 8796 530
rect 8423 474 8484 508
rect 8530 496 8574 508
rect 8630 496 8664 508
rect 8730 496 8754 508
rect 8518 474 8574 496
rect 8608 474 8664 496
rect 8698 474 8754 496
rect 8788 496 8796 508
rect 8830 508 8896 530
rect 8830 496 8844 508
rect 8788 474 8844 496
rect 8878 496 8896 508
rect 8930 508 8996 530
rect 9030 508 9117 530
rect 8930 496 8934 508
rect 8878 474 8934 496
rect 8968 496 8996 508
rect 8968 474 9024 496
rect 9058 474 9117 508
rect 8423 430 9117 474
rect 8423 418 8496 430
rect 8530 418 8596 430
rect 8630 418 8696 430
rect 8730 418 8796 430
rect 8423 384 8484 418
rect 8530 396 8574 418
rect 8630 396 8664 418
rect 8730 396 8754 418
rect 8518 384 8574 396
rect 8608 384 8664 396
rect 8698 384 8754 396
rect 8788 396 8796 418
rect 8830 418 8896 430
rect 8830 396 8844 418
rect 8788 384 8844 396
rect 8878 396 8896 418
rect 8930 418 8996 430
rect 9030 418 9117 430
rect 8930 396 8934 418
rect 8878 384 8934 396
rect 8968 396 8996 418
rect 8968 384 9024 396
rect 9058 384 9117 418
rect 8423 323 9117 384
rect 9170 986 9420 1022
rect 9170 966 9347 986
rect 9170 932 9198 966
rect 9232 952 9347 966
rect 9381 952 9420 986
rect 9232 932 9420 952
rect 9170 896 9420 932
rect 9170 876 9347 896
rect 9170 842 9198 876
rect 9232 862 9347 876
rect 9381 862 9420 896
rect 9232 842 9420 862
rect 9170 806 9420 842
rect 9170 786 9347 806
rect 9170 752 9198 786
rect 9232 772 9347 786
rect 9381 772 9420 806
rect 9232 752 9420 772
rect 9170 716 9420 752
rect 9170 696 9347 716
rect 9170 662 9198 696
rect 9232 682 9347 696
rect 9381 682 9420 716
rect 9232 662 9420 682
rect 9170 626 9420 662
rect 9170 606 9347 626
rect 9170 572 9198 606
rect 9232 592 9347 606
rect 9381 592 9420 626
rect 9232 572 9420 592
rect 9170 536 9420 572
rect 9170 516 9347 536
rect 9170 482 9198 516
rect 9232 502 9347 516
rect 9381 502 9420 536
rect 9232 482 9420 502
rect 9170 446 9420 482
rect 9170 426 9347 446
rect 9170 392 9198 426
rect 9232 412 9347 426
rect 9381 412 9420 446
rect 9232 392 9420 412
rect 9170 356 9420 392
rect 9170 336 9347 356
rect 7882 302 8370 321
rect 7820 270 8370 302
rect 9170 302 9198 336
rect 9232 322 9347 336
rect 9381 322 9420 356
rect 9232 302 9420 322
rect 9170 270 9420 302
rect 1370 266 9420 270
rect 1370 232 1410 266
rect 1444 242 2597 266
rect 1444 232 1636 242
rect 1370 208 1636 232
rect 1670 208 1726 242
rect 1760 208 1816 242
rect 1850 208 1906 242
rect 1940 208 1996 242
rect 2030 208 2086 242
rect 2120 208 2176 242
rect 2210 208 2266 242
rect 2300 208 2356 242
rect 2390 232 2597 242
rect 2631 232 2760 266
rect 2794 242 3947 266
rect 2794 232 2986 242
rect 2390 208 2986 232
rect 3020 208 3076 242
rect 3110 208 3166 242
rect 3200 208 3256 242
rect 3290 208 3346 242
rect 3380 208 3436 242
rect 3470 208 3526 242
rect 3560 208 3616 242
rect 3650 208 3706 242
rect 3740 232 3947 242
rect 3981 232 4110 266
rect 4144 242 5297 266
rect 4144 232 4336 242
rect 3740 208 4336 232
rect 4370 208 4426 242
rect 4460 208 4516 242
rect 4550 208 4606 242
rect 4640 208 4696 242
rect 4730 208 4786 242
rect 4820 208 4876 242
rect 4910 208 4966 242
rect 5000 208 5056 242
rect 5090 232 5297 242
rect 5331 232 5460 266
rect 5494 242 6647 266
rect 5494 232 5686 242
rect 5090 208 5686 232
rect 5720 208 5776 242
rect 5810 208 5866 242
rect 5900 208 5956 242
rect 5990 208 6046 242
rect 6080 208 6136 242
rect 6170 208 6226 242
rect 6260 208 6316 242
rect 6350 208 6406 242
rect 6440 232 6647 242
rect 6681 232 6810 266
rect 6844 242 7997 266
rect 6844 232 7036 242
rect 6440 208 7036 232
rect 7070 208 7126 242
rect 7160 208 7216 242
rect 7250 208 7306 242
rect 7340 208 7396 242
rect 7430 208 7486 242
rect 7520 208 7576 242
rect 7610 208 7666 242
rect 7700 208 7756 242
rect 7790 232 7997 242
rect 8031 232 8160 266
rect 8194 242 9347 266
rect 8194 232 8386 242
rect 7790 208 8386 232
rect 8420 208 8476 242
rect 8510 208 8566 242
rect 8600 208 8656 242
rect 8690 208 8746 242
rect 8780 208 8836 242
rect 8870 208 8926 242
rect 8960 208 9016 242
rect 9050 208 9106 242
rect 9140 232 9347 242
rect 9381 232 9420 266
rect 9140 208 9420 232
rect 1370 176 9420 208
rect 1370 142 1410 176
rect 1444 142 2597 176
rect 2631 142 2760 176
rect 2794 142 3947 176
rect 3981 142 4110 176
rect 4144 142 5297 176
rect 5331 142 5460 176
rect 5494 142 6647 176
rect 6681 142 6810 176
rect 6844 142 7997 176
rect 8031 142 8160 176
rect 8194 142 9347 176
rect 9381 142 9420 176
rect 1370 92 9420 142
rect 1370 58 1506 92
rect 1540 58 1596 92
rect 1630 58 1686 92
rect 1720 58 1776 92
rect 1810 58 1866 92
rect 1900 58 1956 92
rect 1990 58 2046 92
rect 2080 58 2136 92
rect 2170 58 2226 92
rect 2260 58 2316 92
rect 2350 58 2406 92
rect 2440 58 2496 92
rect 2530 58 2856 92
rect 2890 58 2946 92
rect 2980 58 3036 92
rect 3070 58 3126 92
rect 3160 58 3216 92
rect 3250 58 3306 92
rect 3340 58 3396 92
rect 3430 58 3486 92
rect 3520 58 3576 92
rect 3610 58 3666 92
rect 3700 58 3756 92
rect 3790 58 3846 92
rect 3880 58 4206 92
rect 4240 58 4296 92
rect 4330 58 4386 92
rect 4420 58 4476 92
rect 4510 58 4566 92
rect 4600 58 4656 92
rect 4690 58 4746 92
rect 4780 58 4836 92
rect 4870 58 4926 92
rect 4960 58 5016 92
rect 5050 58 5106 92
rect 5140 58 5196 92
rect 5230 58 5556 92
rect 5590 58 5646 92
rect 5680 58 5736 92
rect 5770 58 5826 92
rect 5860 58 5916 92
rect 5950 58 6006 92
rect 6040 58 6096 92
rect 6130 58 6186 92
rect 6220 58 6276 92
rect 6310 58 6366 92
rect 6400 58 6456 92
rect 6490 58 6546 92
rect 6580 58 6906 92
rect 6940 58 6996 92
rect 7030 58 7086 92
rect 7120 58 7176 92
rect 7210 58 7266 92
rect 7300 58 7356 92
rect 7390 58 7446 92
rect 7480 58 7536 92
rect 7570 58 7626 92
rect 7660 58 7716 92
rect 7750 58 7806 92
rect 7840 58 7896 92
rect 7930 58 8256 92
rect 8290 58 8346 92
rect 8380 58 8436 92
rect 8470 58 8526 92
rect 8560 58 8616 92
rect 8650 58 8706 92
rect 8740 58 8796 92
rect 8830 58 8886 92
rect 8920 58 8976 92
rect 9010 58 9066 92
rect 9100 58 9156 92
rect 9190 58 9246 92
rect 9280 58 9420 92
rect 1370 20 9420 58
<< viali >>
rect 5320 4910 5360 4950
rect 5760 4910 5800 4950
rect 6200 4910 6240 4950
rect 6640 4910 6680 4950
rect 7080 4910 7120 4950
rect 7520 4910 7560 4950
rect 7960 4910 8000 4950
rect 7300 4370 7340 4410
rect 6640 4280 6680 4320
rect 7640 4280 7680 4320
rect 5540 4170 5580 4210
rect 6640 4160 6680 4200
rect 7740 4170 7780 4210
rect 5980 4060 6020 4100
rect 7300 4060 7340 4100
rect 6310 3960 6350 4000
rect 6640 3960 6680 4000
rect 6970 3960 7010 4000
rect 5980 3620 6020 3660
rect 7300 3620 7340 3660
rect 5760 3530 5800 3570
rect 6200 3530 6240 3570
rect 6640 3530 6680 3570
rect 7080 3530 7120 3570
rect 7520 3530 7560 3570
rect 7660 3290 7700 3330
rect 1746 924 1768 930
rect 1768 924 1780 930
rect 1846 924 1858 930
rect 1858 924 1880 930
rect 1946 924 1948 930
rect 1948 924 1980 930
rect 1746 896 1780 924
rect 1846 896 1880 924
rect 1946 896 1980 924
rect 2046 896 2080 930
rect 2146 896 2180 930
rect 2246 924 2274 930
rect 2274 924 2280 930
rect 2246 896 2280 924
rect 1746 796 1780 830
rect 1846 796 1880 830
rect 1946 796 1980 830
rect 2046 796 2080 830
rect 2146 796 2180 830
rect 2246 796 2280 830
rect 1746 696 1780 730
rect 1846 696 1880 730
rect 1946 696 1980 730
rect 2046 696 2080 730
rect 2146 696 2180 730
rect 2246 696 2280 730
rect 1746 598 1780 630
rect 1846 598 1880 630
rect 1946 598 1980 630
rect 1746 596 1768 598
rect 1768 596 1780 598
rect 1846 596 1858 598
rect 1858 596 1880 598
rect 1946 596 1948 598
rect 1948 596 1980 598
rect 2046 596 2080 630
rect 2146 596 2180 630
rect 2246 598 2280 630
rect 2246 596 2274 598
rect 2274 596 2280 598
rect 1746 508 1780 530
rect 1846 508 1880 530
rect 1946 508 1980 530
rect 1746 496 1768 508
rect 1768 496 1780 508
rect 1846 496 1858 508
rect 1858 496 1880 508
rect 1946 496 1948 508
rect 1948 496 1980 508
rect 2046 496 2080 530
rect 2146 496 2180 530
rect 2246 508 2280 530
rect 2246 496 2274 508
rect 2274 496 2280 508
rect 1746 418 1780 430
rect 1846 418 1880 430
rect 1946 418 1980 430
rect 1746 396 1768 418
rect 1768 396 1780 418
rect 1846 396 1858 418
rect 1858 396 1880 418
rect 1946 396 1948 418
rect 1948 396 1980 418
rect 2046 396 2080 430
rect 2146 396 2180 430
rect 2246 418 2280 430
rect 2246 396 2274 418
rect 2274 396 2280 418
rect 3096 924 3118 930
rect 3118 924 3130 930
rect 3196 924 3208 930
rect 3208 924 3230 930
rect 3296 924 3298 930
rect 3298 924 3330 930
rect 3096 896 3130 924
rect 3196 896 3230 924
rect 3296 896 3330 924
rect 3396 896 3430 930
rect 3496 896 3530 930
rect 3596 924 3624 930
rect 3624 924 3630 930
rect 3596 896 3630 924
rect 3096 796 3130 830
rect 3196 796 3230 830
rect 3296 796 3330 830
rect 3396 796 3430 830
rect 3496 796 3530 830
rect 3596 796 3630 830
rect 3096 696 3130 730
rect 3196 696 3230 730
rect 3296 696 3330 730
rect 3396 696 3430 730
rect 3496 696 3530 730
rect 3596 696 3630 730
rect 3096 598 3130 630
rect 3196 598 3230 630
rect 3296 598 3330 630
rect 3096 596 3118 598
rect 3118 596 3130 598
rect 3196 596 3208 598
rect 3208 596 3230 598
rect 3296 596 3298 598
rect 3298 596 3330 598
rect 3396 596 3430 630
rect 3496 596 3530 630
rect 3596 598 3630 630
rect 3596 596 3624 598
rect 3624 596 3630 598
rect 3096 508 3130 530
rect 3196 508 3230 530
rect 3296 508 3330 530
rect 3096 496 3118 508
rect 3118 496 3130 508
rect 3196 496 3208 508
rect 3208 496 3230 508
rect 3296 496 3298 508
rect 3298 496 3330 508
rect 3396 496 3430 530
rect 3496 496 3530 530
rect 3596 508 3630 530
rect 3596 496 3624 508
rect 3624 496 3630 508
rect 3096 418 3130 430
rect 3196 418 3230 430
rect 3296 418 3330 430
rect 3096 396 3118 418
rect 3118 396 3130 418
rect 3196 396 3208 418
rect 3208 396 3230 418
rect 3296 396 3298 418
rect 3298 396 3330 418
rect 3396 396 3430 430
rect 3496 396 3530 430
rect 3596 418 3630 430
rect 3596 396 3624 418
rect 3624 396 3630 418
rect 4446 924 4468 930
rect 4468 924 4480 930
rect 4546 924 4558 930
rect 4558 924 4580 930
rect 4646 924 4648 930
rect 4648 924 4680 930
rect 4446 896 4480 924
rect 4546 896 4580 924
rect 4646 896 4680 924
rect 4746 896 4780 930
rect 4846 896 4880 930
rect 4946 924 4974 930
rect 4974 924 4980 930
rect 4946 896 4980 924
rect 4446 796 4480 830
rect 4546 796 4580 830
rect 4646 796 4680 830
rect 4746 796 4780 830
rect 4846 796 4880 830
rect 4946 796 4980 830
rect 4446 696 4480 730
rect 4546 696 4580 730
rect 4646 696 4680 730
rect 4746 696 4780 730
rect 4846 696 4880 730
rect 4946 696 4980 730
rect 4446 598 4480 630
rect 4546 598 4580 630
rect 4646 598 4680 630
rect 4446 596 4468 598
rect 4468 596 4480 598
rect 4546 596 4558 598
rect 4558 596 4580 598
rect 4646 596 4648 598
rect 4648 596 4680 598
rect 4746 596 4780 630
rect 4846 596 4880 630
rect 4946 598 4980 630
rect 4946 596 4974 598
rect 4974 596 4980 598
rect 4446 508 4480 530
rect 4546 508 4580 530
rect 4646 508 4680 530
rect 4446 496 4468 508
rect 4468 496 4480 508
rect 4546 496 4558 508
rect 4558 496 4580 508
rect 4646 496 4648 508
rect 4648 496 4680 508
rect 4746 496 4780 530
rect 4846 496 4880 530
rect 4946 508 4980 530
rect 4946 496 4974 508
rect 4974 496 4980 508
rect 4446 418 4480 430
rect 4546 418 4580 430
rect 4646 418 4680 430
rect 4446 396 4468 418
rect 4468 396 4480 418
rect 4546 396 4558 418
rect 4558 396 4580 418
rect 4646 396 4648 418
rect 4648 396 4680 418
rect 4746 396 4780 430
rect 4846 396 4880 430
rect 4946 418 4980 430
rect 4946 396 4974 418
rect 4974 396 4980 418
rect 5796 924 5818 930
rect 5818 924 5830 930
rect 5896 924 5908 930
rect 5908 924 5930 930
rect 5996 924 5998 930
rect 5998 924 6030 930
rect 5796 896 5830 924
rect 5896 896 5930 924
rect 5996 896 6030 924
rect 6096 896 6130 930
rect 6196 896 6230 930
rect 6296 924 6324 930
rect 6324 924 6330 930
rect 6296 896 6330 924
rect 5796 796 5830 830
rect 5896 796 5930 830
rect 5996 796 6030 830
rect 6096 796 6130 830
rect 6196 796 6230 830
rect 6296 796 6330 830
rect 5796 696 5830 730
rect 5896 696 5930 730
rect 5996 696 6030 730
rect 6096 696 6130 730
rect 6196 696 6230 730
rect 6296 696 6330 730
rect 5796 598 5830 630
rect 5896 598 5930 630
rect 5996 598 6030 630
rect 5796 596 5818 598
rect 5818 596 5830 598
rect 5896 596 5908 598
rect 5908 596 5930 598
rect 5996 596 5998 598
rect 5998 596 6030 598
rect 6096 596 6130 630
rect 6196 596 6230 630
rect 6296 598 6330 630
rect 6296 596 6324 598
rect 6324 596 6330 598
rect 5796 508 5830 530
rect 5896 508 5930 530
rect 5996 508 6030 530
rect 5796 496 5818 508
rect 5818 496 5830 508
rect 5896 496 5908 508
rect 5908 496 5930 508
rect 5996 496 5998 508
rect 5998 496 6030 508
rect 6096 496 6130 530
rect 6196 496 6230 530
rect 6296 508 6330 530
rect 6296 496 6324 508
rect 6324 496 6330 508
rect 5796 418 5830 430
rect 5896 418 5930 430
rect 5996 418 6030 430
rect 5796 396 5818 418
rect 5818 396 5830 418
rect 5896 396 5908 418
rect 5908 396 5930 418
rect 5996 396 5998 418
rect 5998 396 6030 418
rect 6096 396 6130 430
rect 6196 396 6230 430
rect 6296 418 6330 430
rect 6296 396 6324 418
rect 6324 396 6330 418
rect 7146 924 7168 930
rect 7168 924 7180 930
rect 7246 924 7258 930
rect 7258 924 7280 930
rect 7346 924 7348 930
rect 7348 924 7380 930
rect 7146 896 7180 924
rect 7246 896 7280 924
rect 7346 896 7380 924
rect 7446 896 7480 930
rect 7546 896 7580 930
rect 7646 924 7674 930
rect 7674 924 7680 930
rect 7646 896 7680 924
rect 7146 796 7180 830
rect 7246 796 7280 830
rect 7346 796 7380 830
rect 7446 796 7480 830
rect 7546 796 7580 830
rect 7646 796 7680 830
rect 7146 696 7180 730
rect 7246 696 7280 730
rect 7346 696 7380 730
rect 7446 696 7480 730
rect 7546 696 7580 730
rect 7646 696 7680 730
rect 7146 598 7180 630
rect 7246 598 7280 630
rect 7346 598 7380 630
rect 7146 596 7168 598
rect 7168 596 7180 598
rect 7246 596 7258 598
rect 7258 596 7280 598
rect 7346 596 7348 598
rect 7348 596 7380 598
rect 7446 596 7480 630
rect 7546 596 7580 630
rect 7646 598 7680 630
rect 7646 596 7674 598
rect 7674 596 7680 598
rect 7146 508 7180 530
rect 7246 508 7280 530
rect 7346 508 7380 530
rect 7146 496 7168 508
rect 7168 496 7180 508
rect 7246 496 7258 508
rect 7258 496 7280 508
rect 7346 496 7348 508
rect 7348 496 7380 508
rect 7446 496 7480 530
rect 7546 496 7580 530
rect 7646 508 7680 530
rect 7646 496 7674 508
rect 7674 496 7680 508
rect 7146 418 7180 430
rect 7246 418 7280 430
rect 7346 418 7380 430
rect 7146 396 7168 418
rect 7168 396 7180 418
rect 7246 396 7258 418
rect 7258 396 7280 418
rect 7346 396 7348 418
rect 7348 396 7380 418
rect 7446 396 7480 430
rect 7546 396 7580 430
rect 7646 418 7680 430
rect 7646 396 7674 418
rect 7674 396 7680 418
rect 8496 924 8518 930
rect 8518 924 8530 930
rect 8596 924 8608 930
rect 8608 924 8630 930
rect 8696 924 8698 930
rect 8698 924 8730 930
rect 8496 896 8530 924
rect 8596 896 8630 924
rect 8696 896 8730 924
rect 8796 896 8830 930
rect 8896 896 8930 930
rect 8996 924 9024 930
rect 9024 924 9030 930
rect 8996 896 9030 924
rect 8496 796 8530 830
rect 8596 796 8630 830
rect 8696 796 8730 830
rect 8796 796 8830 830
rect 8896 796 8930 830
rect 8996 796 9030 830
rect 8496 696 8530 730
rect 8596 696 8630 730
rect 8696 696 8730 730
rect 8796 696 8830 730
rect 8896 696 8930 730
rect 8996 696 9030 730
rect 8496 598 8530 630
rect 8596 598 8630 630
rect 8696 598 8730 630
rect 8496 596 8518 598
rect 8518 596 8530 598
rect 8596 596 8608 598
rect 8608 596 8630 598
rect 8696 596 8698 598
rect 8698 596 8730 598
rect 8796 596 8830 630
rect 8896 596 8930 630
rect 8996 598 9030 630
rect 8996 596 9024 598
rect 9024 596 9030 598
rect 8496 508 8530 530
rect 8596 508 8630 530
rect 8696 508 8730 530
rect 8496 496 8518 508
rect 8518 496 8530 508
rect 8596 496 8608 508
rect 8608 496 8630 508
rect 8696 496 8698 508
rect 8698 496 8730 508
rect 8796 496 8830 530
rect 8896 496 8930 530
rect 8996 508 9030 530
rect 8996 496 9024 508
rect 9024 496 9030 508
rect 8496 418 8530 430
rect 8596 418 8630 430
rect 8696 418 8730 430
rect 8496 396 8518 418
rect 8518 396 8530 418
rect 8596 396 8608 418
rect 8608 396 8630 418
rect 8696 396 8698 418
rect 8698 396 8730 418
rect 8796 396 8830 430
rect 8896 396 8930 430
rect 8996 418 9030 430
rect 8996 396 9024 418
rect 9024 396 9030 418
<< metal1 >>
rect 5300 4960 5380 4970
rect 5300 4900 5310 4960
rect 5370 4900 5380 4960
rect 5300 4890 5380 4900
rect 5740 4960 5820 4970
rect 5740 4900 5750 4960
rect 5810 4900 5820 4960
rect 5740 4890 5820 4900
rect 6180 4960 6260 4970
rect 6180 4900 6190 4960
rect 6250 4900 6260 4960
rect 6180 4890 6260 4900
rect 6620 4960 6700 4970
rect 6620 4900 6630 4960
rect 6690 4900 6700 4960
rect 6620 4890 6700 4900
rect 7060 4960 7140 4970
rect 7060 4900 7070 4960
rect 7130 4900 7140 4960
rect 7060 4890 7140 4900
rect 7500 4960 7580 4970
rect 7500 4900 7510 4960
rect 7570 4900 7580 4960
rect 7500 4890 7580 4900
rect 7940 4960 8020 4970
rect 7940 4900 7950 4960
rect 8010 4900 8020 4960
rect 7940 4890 8020 4900
rect 5960 4420 6040 4430
rect 5960 4360 5970 4420
rect 6030 4360 6040 4420
rect 5960 4350 6040 4360
rect 7280 4420 7360 4430
rect 7280 4360 7290 4420
rect 7350 4360 7360 4420
rect 7280 4350 7360 4360
rect 5520 4220 5600 4230
rect 5520 4160 5530 4220
rect 5590 4160 5600 4220
rect 5520 4150 5600 4160
rect 5980 4120 6020 4350
rect 6620 4330 6700 4340
rect 6620 4270 6630 4330
rect 6690 4270 6700 4330
rect 6620 4260 6700 4270
rect 6620 4210 6700 4220
rect 6620 4150 6630 4210
rect 6690 4150 6700 4210
rect 6620 4140 6700 4150
rect 5960 4110 6040 4120
rect 5960 4050 5970 4110
rect 6030 4050 6040 4110
rect 5960 4040 6040 4050
rect 6640 4020 6680 4140
rect 7300 4120 7340 4350
rect 7620 4330 7700 4340
rect 7620 4270 7630 4330
rect 7690 4270 7700 4330
rect 7620 4260 7700 4270
rect 7280 4110 7360 4120
rect 7280 4050 7290 4110
rect 7350 4050 7360 4110
rect 7280 4040 7360 4050
rect 6290 4010 6370 4020
rect 6290 3950 6300 4010
rect 6360 3950 6370 4010
rect 6290 3940 6370 3950
rect 6620 4000 6700 4020
rect 6620 3960 6640 4000
rect 6680 3960 6700 4000
rect 6620 3940 6700 3960
rect 6950 4010 7030 4020
rect 6950 3950 6960 4010
rect 7020 3950 7030 4010
rect 6950 3940 7030 3950
rect 5960 3670 6040 3680
rect 5960 3610 5970 3670
rect 6030 3610 6040 3670
rect 7280 3670 7360 3680
rect 7280 3610 7290 3670
rect 7350 3610 7360 3670
rect 7280 3600 7360 3610
rect 5740 3580 5820 3590
rect 5740 3520 5750 3580
rect 5810 3520 5820 3580
rect 5740 3510 5820 3520
rect 6180 3580 6260 3590
rect 6180 3520 6190 3580
rect 6250 3520 6260 3580
rect 6180 3510 6260 3520
rect 6620 3580 6700 3590
rect 6620 3520 6630 3580
rect 6690 3520 6700 3580
rect 6620 3510 6700 3520
rect 7060 3580 7140 3590
rect 7060 3520 7070 3580
rect 7130 3520 7140 3580
rect 7060 3510 7140 3520
rect 7500 3580 7580 3590
rect 7500 3520 7510 3580
rect 7570 3520 7580 3580
rect 7500 3510 7580 3520
rect 7640 3350 7680 4260
rect 7720 4220 7800 4230
rect 7720 4160 7730 4220
rect 7790 4160 7800 4220
rect 7720 4150 7800 4160
rect 7640 3330 7720 3350
rect 7640 3290 7660 3330
rect 7700 3290 7720 3330
rect 7640 3270 7720 3290
rect 370 370 970 1460
rect 1720 1420 9070 1460
rect 1720 975 2320 1420
rect 3070 975 3670 1420
rect 4420 975 5020 1420
rect 5770 975 6370 1420
rect 7120 975 7720 1420
rect 8470 975 9070 1420
rect 1715 930 2325 975
rect 1715 896 1746 930
rect 1780 896 1846 930
rect 1880 896 1946 930
rect 1980 896 2046 930
rect 2080 896 2146 930
rect 2180 896 2246 930
rect 2280 896 2325 930
rect 1715 830 2325 896
rect 1715 796 1746 830
rect 1780 796 1846 830
rect 1880 796 1946 830
rect 1980 796 2046 830
rect 2080 796 2146 830
rect 2180 796 2246 830
rect 2280 796 2325 830
rect 1715 730 2325 796
rect 1715 696 1746 730
rect 1780 696 1846 730
rect 1880 696 1946 730
rect 1980 696 2046 730
rect 2080 696 2146 730
rect 2180 696 2246 730
rect 2280 696 2325 730
rect 1715 630 2325 696
rect 1715 596 1746 630
rect 1780 596 1846 630
rect 1880 596 1946 630
rect 1980 596 2046 630
rect 2080 596 2146 630
rect 2180 596 2246 630
rect 2280 596 2325 630
rect 1715 530 2325 596
rect 1715 496 1746 530
rect 1780 496 1846 530
rect 1880 496 1946 530
rect 1980 496 2046 530
rect 2080 496 2146 530
rect 2180 496 2246 530
rect 2280 496 2325 530
rect 1715 430 2325 496
rect 1715 396 1746 430
rect 1780 396 1846 430
rect 1880 396 1946 430
rect 1980 396 2046 430
rect 2080 396 2146 430
rect 2180 396 2246 430
rect 2280 396 2325 430
rect 1715 365 2325 396
rect 3065 930 3675 975
rect 3065 896 3096 930
rect 3130 896 3196 930
rect 3230 896 3296 930
rect 3330 896 3396 930
rect 3430 896 3496 930
rect 3530 896 3596 930
rect 3630 896 3675 930
rect 3065 830 3675 896
rect 3065 796 3096 830
rect 3130 796 3196 830
rect 3230 796 3296 830
rect 3330 796 3396 830
rect 3430 796 3496 830
rect 3530 796 3596 830
rect 3630 796 3675 830
rect 3065 730 3675 796
rect 3065 696 3096 730
rect 3130 696 3196 730
rect 3230 696 3296 730
rect 3330 696 3396 730
rect 3430 696 3496 730
rect 3530 696 3596 730
rect 3630 696 3675 730
rect 3065 630 3675 696
rect 3065 596 3096 630
rect 3130 596 3196 630
rect 3230 596 3296 630
rect 3330 596 3396 630
rect 3430 596 3496 630
rect 3530 596 3596 630
rect 3630 596 3675 630
rect 3065 530 3675 596
rect 3065 496 3096 530
rect 3130 496 3196 530
rect 3230 496 3296 530
rect 3330 496 3396 530
rect 3430 496 3496 530
rect 3530 496 3596 530
rect 3630 496 3675 530
rect 3065 430 3675 496
rect 3065 396 3096 430
rect 3130 396 3196 430
rect 3230 396 3296 430
rect 3330 396 3396 430
rect 3430 396 3496 430
rect 3530 396 3596 430
rect 3630 396 3675 430
rect 3065 365 3675 396
rect 4415 930 5025 975
rect 4415 896 4446 930
rect 4480 896 4546 930
rect 4580 896 4646 930
rect 4680 896 4746 930
rect 4780 896 4846 930
rect 4880 896 4946 930
rect 4980 896 5025 930
rect 4415 830 5025 896
rect 4415 796 4446 830
rect 4480 796 4546 830
rect 4580 796 4646 830
rect 4680 796 4746 830
rect 4780 796 4846 830
rect 4880 796 4946 830
rect 4980 796 5025 830
rect 4415 730 5025 796
rect 4415 696 4446 730
rect 4480 696 4546 730
rect 4580 696 4646 730
rect 4680 696 4746 730
rect 4780 696 4846 730
rect 4880 696 4946 730
rect 4980 696 5025 730
rect 4415 630 5025 696
rect 4415 596 4446 630
rect 4480 596 4546 630
rect 4580 596 4646 630
rect 4680 596 4746 630
rect 4780 596 4846 630
rect 4880 596 4946 630
rect 4980 596 5025 630
rect 4415 530 5025 596
rect 4415 496 4446 530
rect 4480 496 4546 530
rect 4580 496 4646 530
rect 4680 496 4746 530
rect 4780 496 4846 530
rect 4880 496 4946 530
rect 4980 496 5025 530
rect 4415 430 5025 496
rect 4415 396 4446 430
rect 4480 396 4546 430
rect 4580 396 4646 430
rect 4680 396 4746 430
rect 4780 396 4846 430
rect 4880 396 4946 430
rect 4980 396 5025 430
rect 4415 365 5025 396
rect 5765 930 6375 975
rect 5765 896 5796 930
rect 5830 896 5896 930
rect 5930 896 5996 930
rect 6030 896 6096 930
rect 6130 896 6196 930
rect 6230 896 6296 930
rect 6330 896 6375 930
rect 5765 830 6375 896
rect 5765 796 5796 830
rect 5830 796 5896 830
rect 5930 796 5996 830
rect 6030 796 6096 830
rect 6130 796 6196 830
rect 6230 796 6296 830
rect 6330 796 6375 830
rect 5765 730 6375 796
rect 5765 696 5796 730
rect 5830 696 5896 730
rect 5930 696 5996 730
rect 6030 696 6096 730
rect 6130 696 6196 730
rect 6230 696 6296 730
rect 6330 696 6375 730
rect 5765 630 6375 696
rect 5765 596 5796 630
rect 5830 596 5896 630
rect 5930 596 5996 630
rect 6030 596 6096 630
rect 6130 596 6196 630
rect 6230 596 6296 630
rect 6330 596 6375 630
rect 5765 530 6375 596
rect 5765 496 5796 530
rect 5830 496 5896 530
rect 5930 496 5996 530
rect 6030 496 6096 530
rect 6130 496 6196 530
rect 6230 496 6296 530
rect 6330 496 6375 530
rect 5765 430 6375 496
rect 5765 396 5796 430
rect 5830 396 5896 430
rect 5930 396 5996 430
rect 6030 396 6096 430
rect 6130 396 6196 430
rect 6230 396 6296 430
rect 6330 396 6375 430
rect 5765 365 6375 396
rect 7115 930 7725 975
rect 7115 896 7146 930
rect 7180 896 7246 930
rect 7280 896 7346 930
rect 7380 896 7446 930
rect 7480 896 7546 930
rect 7580 896 7646 930
rect 7680 896 7725 930
rect 7115 830 7725 896
rect 7115 796 7146 830
rect 7180 796 7246 830
rect 7280 796 7346 830
rect 7380 796 7446 830
rect 7480 796 7546 830
rect 7580 796 7646 830
rect 7680 796 7725 830
rect 7115 730 7725 796
rect 7115 696 7146 730
rect 7180 696 7246 730
rect 7280 696 7346 730
rect 7380 696 7446 730
rect 7480 696 7546 730
rect 7580 696 7646 730
rect 7680 696 7725 730
rect 7115 630 7725 696
rect 7115 596 7146 630
rect 7180 596 7246 630
rect 7280 596 7346 630
rect 7380 596 7446 630
rect 7480 596 7546 630
rect 7580 596 7646 630
rect 7680 596 7725 630
rect 7115 530 7725 596
rect 7115 496 7146 530
rect 7180 496 7246 530
rect 7280 496 7346 530
rect 7380 496 7446 530
rect 7480 496 7546 530
rect 7580 496 7646 530
rect 7680 496 7725 530
rect 7115 430 7725 496
rect 7115 396 7146 430
rect 7180 396 7246 430
rect 7280 396 7346 430
rect 7380 396 7446 430
rect 7480 396 7546 430
rect 7580 396 7646 430
rect 7680 396 7725 430
rect 7115 365 7725 396
rect 8465 930 9075 975
rect 8465 896 8496 930
rect 8530 896 8596 930
rect 8630 896 8696 930
rect 8730 896 8796 930
rect 8830 896 8896 930
rect 8930 896 8996 930
rect 9030 896 9075 930
rect 8465 830 9075 896
rect 8465 796 8496 830
rect 8530 796 8596 830
rect 8630 796 8696 830
rect 8730 796 8796 830
rect 8830 796 8896 830
rect 8930 796 8996 830
rect 9030 796 9075 830
rect 8465 730 9075 796
rect 8465 696 8496 730
rect 8530 696 8596 730
rect 8630 696 8696 730
rect 8730 696 8796 730
rect 8830 696 8896 730
rect 8930 696 8996 730
rect 9030 696 9075 730
rect 8465 630 9075 696
rect 8465 596 8496 630
rect 8530 596 8596 630
rect 8630 596 8696 630
rect 8730 596 8796 630
rect 8830 596 8896 630
rect 8930 596 8996 630
rect 9030 596 9075 630
rect 8465 530 9075 596
rect 8465 496 8496 530
rect 8530 496 8596 530
rect 8630 496 8696 530
rect 8730 496 8796 530
rect 8830 496 8896 530
rect 8930 496 8996 530
rect 9030 496 9075 530
rect 8465 430 9075 496
rect 8465 396 8496 430
rect 8530 396 8596 430
rect 8630 396 8696 430
rect 8730 396 8796 430
rect 8830 396 8896 430
rect 8930 396 8996 430
rect 9030 396 9075 430
rect 8465 365 9075 396
<< via1 >>
rect 5310 4950 5370 4960
rect 5310 4910 5320 4950
rect 5320 4910 5360 4950
rect 5360 4910 5370 4950
rect 5310 4900 5370 4910
rect 5750 4950 5810 4960
rect 5750 4910 5760 4950
rect 5760 4910 5800 4950
rect 5800 4910 5810 4950
rect 5750 4900 5810 4910
rect 6190 4950 6250 4960
rect 6190 4910 6200 4950
rect 6200 4910 6240 4950
rect 6240 4910 6250 4950
rect 6190 4900 6250 4910
rect 6630 4950 6690 4960
rect 6630 4910 6640 4950
rect 6640 4910 6680 4950
rect 6680 4910 6690 4950
rect 6630 4900 6690 4910
rect 7070 4950 7130 4960
rect 7070 4910 7080 4950
rect 7080 4910 7120 4950
rect 7120 4910 7130 4950
rect 7070 4900 7130 4910
rect 7510 4950 7570 4960
rect 7510 4910 7520 4950
rect 7520 4910 7560 4950
rect 7560 4910 7570 4950
rect 7510 4900 7570 4910
rect 7950 4950 8010 4960
rect 7950 4910 7960 4950
rect 7960 4910 8000 4950
rect 8000 4910 8010 4950
rect 7950 4900 8010 4910
rect 5970 4360 6030 4420
rect 7290 4410 7350 4420
rect 7290 4370 7300 4410
rect 7300 4370 7340 4410
rect 7340 4370 7350 4410
rect 7290 4360 7350 4370
rect 5530 4210 5590 4220
rect 5530 4170 5540 4210
rect 5540 4170 5580 4210
rect 5580 4170 5590 4210
rect 5530 4160 5590 4170
rect 6630 4320 6690 4330
rect 6630 4280 6640 4320
rect 6640 4280 6680 4320
rect 6680 4280 6690 4320
rect 6630 4270 6690 4280
rect 6630 4200 6690 4210
rect 6630 4160 6640 4200
rect 6640 4160 6680 4200
rect 6680 4160 6690 4200
rect 6630 4150 6690 4160
rect 5970 4100 6030 4110
rect 5970 4060 5980 4100
rect 5980 4060 6020 4100
rect 6020 4060 6030 4100
rect 5970 4050 6030 4060
rect 7630 4320 7690 4330
rect 7630 4280 7640 4320
rect 7640 4280 7680 4320
rect 7680 4280 7690 4320
rect 7630 4270 7690 4280
rect 7290 4100 7350 4110
rect 7290 4060 7300 4100
rect 7300 4060 7340 4100
rect 7340 4060 7350 4100
rect 7290 4050 7350 4060
rect 6300 4000 6360 4010
rect 6300 3960 6310 4000
rect 6310 3960 6350 4000
rect 6350 3960 6360 4000
rect 6300 3950 6360 3960
rect 6960 4000 7020 4010
rect 6960 3960 6970 4000
rect 6970 3960 7010 4000
rect 7010 3960 7020 4000
rect 6960 3950 7020 3960
rect 5970 3660 6030 3670
rect 5970 3620 5980 3660
rect 5980 3620 6020 3660
rect 6020 3620 6030 3660
rect 5970 3610 6030 3620
rect 7290 3660 7350 3670
rect 7290 3620 7300 3660
rect 7300 3620 7340 3660
rect 7340 3620 7350 3660
rect 7290 3610 7350 3620
rect 5750 3570 5810 3580
rect 5750 3530 5760 3570
rect 5760 3530 5800 3570
rect 5800 3530 5810 3570
rect 5750 3520 5810 3530
rect 6190 3570 6250 3580
rect 6190 3530 6200 3570
rect 6200 3530 6240 3570
rect 6240 3530 6250 3570
rect 6190 3520 6250 3530
rect 6630 3570 6690 3580
rect 6630 3530 6640 3570
rect 6640 3530 6680 3570
rect 6680 3530 6690 3570
rect 6630 3520 6690 3530
rect 7070 3570 7130 3580
rect 7070 3530 7080 3570
rect 7080 3530 7120 3570
rect 7120 3530 7130 3570
rect 7070 3520 7130 3530
rect 7510 3570 7570 3580
rect 7510 3530 7520 3570
rect 7520 3530 7560 3570
rect 7560 3530 7570 3570
rect 7510 3520 7570 3530
rect 7730 4210 7790 4220
rect 7730 4170 7740 4210
rect 7740 4170 7780 4210
rect 7780 4170 7790 4210
rect 7730 4160 7790 4170
<< metal2 >>
rect 5300 4960 5380 4970
rect 5300 4900 5310 4960
rect 5370 4950 5380 4960
rect 5740 4960 5820 4970
rect 5740 4950 5750 4960
rect 5370 4910 5750 4950
rect 5370 4900 5380 4910
rect 5300 4890 5380 4900
rect 5740 4900 5750 4910
rect 5810 4950 5820 4960
rect 6180 4960 6260 4970
rect 6180 4950 6190 4960
rect 5810 4910 6190 4950
rect 5810 4900 5820 4910
rect 5740 4890 5820 4900
rect 6180 4900 6190 4910
rect 6250 4950 6260 4960
rect 6620 4960 6700 4970
rect 6620 4950 6630 4960
rect 6250 4910 6630 4950
rect 6250 4900 6260 4910
rect 6180 4890 6260 4900
rect 6620 4900 6630 4910
rect 6690 4950 6700 4960
rect 7060 4960 7140 4970
rect 7060 4950 7070 4960
rect 6690 4910 7070 4950
rect 6690 4900 6700 4910
rect 6620 4890 6700 4900
rect 7060 4900 7070 4910
rect 7130 4950 7140 4960
rect 7500 4960 7580 4970
rect 7500 4950 7510 4960
rect 7130 4910 7510 4950
rect 7130 4900 7140 4910
rect 7060 4890 7140 4900
rect 7500 4900 7510 4910
rect 7570 4950 7580 4960
rect 7940 4960 8020 4970
rect 7940 4950 7950 4960
rect 7570 4910 7950 4950
rect 7570 4900 7580 4910
rect 7500 4890 7580 4900
rect 7940 4900 7950 4910
rect 8010 4900 8020 4960
rect 7940 4890 8020 4900
rect 5960 4420 6040 4430
rect 5960 4360 5970 4420
rect 6030 4410 6040 4420
rect 7280 4420 7360 4430
rect 7280 4410 7290 4420
rect 6030 4370 7290 4410
rect 6030 4360 6040 4370
rect 5960 4350 6040 4360
rect 7280 4360 7290 4370
rect 7350 4360 7360 4420
rect 7280 4350 7360 4360
rect 6620 4330 6700 4340
rect 6620 4270 6630 4330
rect 6690 4320 6700 4330
rect 7620 4330 7700 4340
rect 7620 4320 7630 4330
rect 6690 4280 7630 4320
rect 6690 4270 6700 4280
rect 6620 4260 6700 4270
rect 7620 4270 7630 4280
rect 7690 4270 7700 4330
rect 7620 4260 7700 4270
rect 5520 4220 5600 4230
rect 7720 4220 7800 4230
rect 5520 4160 5530 4220
rect 5590 4200 5600 4220
rect 6620 4210 6700 4220
rect 6620 4200 6630 4210
rect 5590 4160 6630 4200
rect 5520 4150 5600 4160
rect 6620 4150 6630 4160
rect 6690 4200 6700 4210
rect 7720 4200 7730 4220
rect 6690 4160 7730 4200
rect 7790 4160 7800 4220
rect 6690 4150 6700 4160
rect 7720 4150 7800 4160
rect 6620 4140 6700 4150
rect 5960 4110 6040 4120
rect 5960 4050 5970 4110
rect 6030 4100 6040 4110
rect 7280 4110 7360 4120
rect 7280 4100 7290 4110
rect 6030 4060 7290 4100
rect 6030 4050 6040 4060
rect 5960 4040 6040 4050
rect 7280 4050 7290 4060
rect 7350 4050 7360 4110
rect 7280 4040 7360 4050
rect 6290 4010 6370 4020
rect 6290 4000 6300 4010
rect 5510 3960 6300 4000
rect 6290 3950 6300 3960
rect 6360 4000 6370 4010
rect 6950 4010 7030 4020
rect 6950 4000 6960 4010
rect 6360 3960 6960 4000
rect 6360 3950 6370 3960
rect 6290 3940 6370 3950
rect 6950 3950 6960 3960
rect 7020 3950 7030 4010
rect 6950 3940 7030 3950
rect 5960 3670 6040 3680
rect 5960 3660 5970 3670
rect 5510 3620 5970 3660
rect 5960 3610 5970 3620
rect 6030 3660 6040 3670
rect 7280 3670 7360 3680
rect 7280 3660 7290 3670
rect 6030 3620 7290 3660
rect 6030 3610 6040 3620
rect 5960 3600 6040 3610
rect 7280 3610 7290 3620
rect 7350 3610 7360 3670
rect 7280 3600 7360 3610
rect 5740 3580 5820 3590
rect 5740 3520 5750 3580
rect 5810 3570 5820 3580
rect 6180 3580 6260 3590
rect 6180 3570 6190 3580
rect 5810 3530 6190 3570
rect 5810 3520 5820 3530
rect 5740 3510 5820 3520
rect 6180 3520 6190 3530
rect 6250 3570 6260 3580
rect 6620 3580 6700 3590
rect 6620 3570 6630 3580
rect 6250 3530 6630 3570
rect 6250 3520 6260 3530
rect 6180 3510 6260 3520
rect 6620 3520 6630 3530
rect 6690 3570 6700 3580
rect 7060 3580 7140 3590
rect 7060 3570 7070 3580
rect 6690 3530 7070 3570
rect 6690 3520 6700 3530
rect 6620 3510 6700 3520
rect 7060 3520 7070 3530
rect 7130 3570 7140 3580
rect 7500 3580 7580 3590
rect 7500 3570 7510 3580
rect 7130 3530 7510 3570
rect 7130 3520 7140 3530
rect 7060 3510 7140 3520
rect 7500 3520 7510 3530
rect 7570 3520 7580 3580
rect 7500 3510 7580 3520
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 0 0 1 0
box 0 0 1340 1340
<< labels >>
flabel locali s 1940 1102 2058 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 1963 1252 2064 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 1904 626 2152 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 3290 1102 3408 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 3313 1252 3414 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 3254 626 3502 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 4640 1102 4758 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 4663 1252 4764 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 4604 626 4852 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 5990 1102 6108 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 6013 1252 6114 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 5954 626 6202 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 7340 1102 7458 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 7363 1252 7464 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 7304 626 7552 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 8690 1102 8808 1142 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 8713 1252 8814 1301 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 8654 626 8902 730 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
<< end >>
