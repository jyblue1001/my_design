magic
tech sky130A
magscale 1 2
timestamp 1755890037
<< nwell >>
rect 109180 9060 110940 9840
rect 111850 8760 112530 9540
rect 112790 8760 113470 9200
rect 114130 8760 114810 9540
rect 115070 8760 115750 9540
rect 116660 9060 118420 9840
rect 109060 7540 110820 8320
rect 112900 7530 114700 8110
rect 116780 7540 118540 8320
rect 109120 5690 110760 6970
rect 116840 5690 118480 6970
rect 117830 5680 118110 5690
rect 109120 3940 110760 4420
rect 116840 3940 118480 4420
<< nmos >>
rect 113620 6360 113650 6860
rect 113730 6360 113760 6860
rect 113840 6360 113870 6860
rect 113950 6360 113980 6860
rect 112140 5430 112170 5730
rect 112250 5430 112280 5730
rect 112360 5430 112390 5730
rect 112470 5430 112500 5730
rect 112580 5430 112610 5730
rect 112690 5430 112720 5730
rect 112800 5430 112830 5730
rect 112910 5430 112940 5730
rect 113020 5430 113050 5730
rect 113130 5430 113160 5730
rect 113240 5430 113270 5730
rect 113350 5430 113380 5730
rect 114220 5430 114250 5730
rect 114330 5430 114360 5730
rect 114440 5430 114470 5730
rect 114550 5430 114580 5730
rect 114660 5430 114690 5730
rect 114770 5430 114800 5730
rect 114880 5430 114910 5730
rect 114990 5430 115020 5730
rect 115100 5430 115130 5730
rect 115210 5430 115240 5730
rect 115320 5430 115350 5730
rect 115430 5430 115460 5730
rect 112140 3560 112170 3860
rect 112250 3560 112280 3860
rect 112360 3560 112390 3860
rect 112470 3560 112500 3860
rect 112580 3560 112610 3860
rect 112690 3560 112720 3860
rect 112800 3560 112830 3860
rect 112910 3560 112940 3860
rect 113020 3560 113050 3860
rect 113130 3560 113160 3860
rect 113240 3560 113270 3860
rect 113350 3560 113380 3860
rect 113620 3560 113650 3860
rect 113730 3560 113760 3860
rect 113840 3560 113870 3860
rect 113950 3560 113980 3860
rect 114220 3560 114250 3860
rect 114330 3560 114360 3860
rect 114440 3560 114470 3860
rect 114550 3560 114580 3860
rect 114660 3560 114690 3860
rect 114770 3560 114800 3860
rect 114880 3560 114910 3860
rect 114990 3560 115020 3860
rect 115100 3560 115130 3860
rect 115210 3560 115240 3860
rect 115320 3560 115350 3860
rect 115430 3560 115460 3860
rect 109320 2900 109350 3500
rect 109430 2900 109460 3500
rect 109540 2900 109570 3500
rect 109650 2900 109680 3500
rect 109760 2900 109790 3500
rect 109870 2900 109900 3500
rect 109980 2900 110010 3500
rect 110090 2900 110120 3500
rect 110200 2900 110230 3500
rect 110310 2900 110340 3500
rect 110420 2900 110450 3500
rect 110530 2900 110560 3500
rect 117040 2900 117070 3500
rect 117150 2900 117180 3500
rect 117260 2900 117290 3500
rect 117370 2900 117400 3500
rect 117480 2900 117510 3500
rect 117590 2900 117620 3500
rect 117700 2900 117730 3500
rect 117810 2900 117840 3500
rect 117920 2900 117950 3500
rect 118030 2900 118060 3500
rect 118140 2900 118170 3500
rect 118250 2900 118280 3500
rect 109380 -20 109500 1380
rect 109580 -20 109700 1380
rect 109780 -20 109900 1380
rect 109980 -20 110100 1380
rect 110180 -20 110300 1380
rect 110380 -20 110500 1380
rect 112520 1110 112550 1610
rect 112630 1110 112660 1610
rect 112740 1110 112770 1610
rect 112850 1110 112880 1610
rect 112960 1110 112990 1610
rect 113070 1110 113100 1610
rect 113180 1110 113210 1610
rect 113290 1110 113320 1610
rect 113400 1110 113430 1610
rect 113510 1110 113540 1610
rect 113620 1110 113650 1610
rect 113730 1110 113760 1610
rect 113840 1110 113870 1610
rect 113950 1110 113980 1610
rect 114060 1110 114090 1610
rect 114170 1110 114200 1610
rect 114280 1110 114310 1610
rect 114390 1110 114420 1610
rect 114500 1110 114530 1610
rect 114610 1110 114640 1610
rect 114720 1110 114750 1610
rect 114830 1110 114860 1610
rect 114940 1110 114970 1610
rect 113510 -200 113540 100
rect 113620 -200 113650 100
rect 113730 -200 113760 100
rect 113840 -200 113870 100
rect 113950 -200 113980 100
rect 114060 -200 114090 100
rect 117100 -20 117220 1380
rect 117300 -20 117420 1380
rect 117500 -20 117620 1380
rect 117700 -20 117820 1380
rect 117900 -20 118020 1380
rect 118100 -20 118220 1380
rect 113500 -720 114100 -420
<< pmos >>
rect 109380 9100 109420 9800
rect 109500 9100 109540 9800
rect 109620 9100 109660 9800
rect 109740 9100 109780 9800
rect 109860 9100 109900 9800
rect 109980 9100 110020 9800
rect 110100 9100 110140 9800
rect 110220 9100 110260 9800
rect 110340 9100 110380 9800
rect 110460 9100 110500 9800
rect 110580 9100 110620 9800
rect 110700 9100 110740 9800
rect 112050 8800 112090 9500
rect 112170 8800 112210 9500
rect 112290 8800 112330 9500
rect 112990 8800 113030 9160
rect 113110 8800 113150 9160
rect 113230 8800 113270 9160
rect 114330 8800 114370 9500
rect 114450 8800 114490 9500
rect 114570 8800 114610 9500
rect 115270 8800 115310 9500
rect 115390 8800 115430 9500
rect 115510 8800 115550 9500
rect 116860 9100 116900 9800
rect 116980 9100 117020 9800
rect 117100 9100 117140 9800
rect 117220 9100 117260 9800
rect 117340 9100 117380 9800
rect 117460 9100 117500 9800
rect 117580 9100 117620 9800
rect 117700 9100 117740 9800
rect 117820 9100 117860 9800
rect 117940 9100 117980 9800
rect 118060 9100 118100 9800
rect 118180 9100 118220 9800
rect 109260 7580 109300 8280
rect 109380 7580 109420 8280
rect 109500 7580 109540 8280
rect 109620 7580 109660 8280
rect 109740 7580 109780 8280
rect 109860 7580 109900 8280
rect 109980 7580 110020 8280
rect 110100 7580 110140 8280
rect 110220 7580 110260 8280
rect 110340 7580 110380 8280
rect 110460 7580 110500 8280
rect 110580 7580 110620 8280
rect 113100 7570 113130 8070
rect 113210 7570 113240 8070
rect 113320 7570 113350 8070
rect 113430 7570 113460 8070
rect 113540 7570 113570 8070
rect 113650 7570 113680 8070
rect 113920 7570 113950 8070
rect 114030 7570 114060 8070
rect 114140 7570 114170 8070
rect 114250 7570 114280 8070
rect 114360 7570 114390 8070
rect 114470 7570 114500 8070
rect 116980 7580 117020 8280
rect 117100 7580 117140 8280
rect 117220 7580 117260 8280
rect 117340 7580 117380 8280
rect 117460 7580 117500 8280
rect 117580 7580 117620 8280
rect 117700 7580 117740 8280
rect 117820 7580 117860 8280
rect 117940 7580 117980 8280
rect 118060 7580 118100 8280
rect 118180 7580 118220 8280
rect 118300 7580 118340 8280
rect 109320 5730 109350 6930
rect 109430 5730 109460 6930
rect 109540 5730 109570 6930
rect 109650 5730 109680 6930
rect 109760 5730 109790 6930
rect 109870 5730 109900 6930
rect 109980 5730 110010 6930
rect 110090 5730 110120 6930
rect 110200 5730 110230 6930
rect 110310 5730 110340 6930
rect 110420 5730 110450 6930
rect 110530 5730 110560 6930
rect 117040 5730 117070 6930
rect 117150 5730 117180 6930
rect 117260 5730 117290 6930
rect 117370 5730 117400 6930
rect 117480 5730 117510 6930
rect 117590 5730 117620 6930
rect 117700 5730 117730 6930
rect 117810 5730 117840 6930
rect 117920 5730 117950 6930
rect 118030 5730 118060 6930
rect 118140 5730 118170 6930
rect 118250 5730 118280 6930
rect 109320 3980 109350 4380
rect 109430 3980 109460 4380
rect 109540 3980 109570 4380
rect 109650 3980 109680 4380
rect 109760 3980 109790 4380
rect 109870 3980 109900 4380
rect 109980 3980 110010 4380
rect 110090 3980 110120 4380
rect 110200 3980 110230 4380
rect 110310 3980 110340 4380
rect 110420 3980 110450 4380
rect 110530 3980 110560 4380
rect 117040 3980 117070 4380
rect 117150 3980 117180 4380
rect 117260 3980 117290 4380
rect 117370 3980 117400 4380
rect 117480 3980 117510 4380
rect 117590 3980 117620 4380
rect 117700 3980 117730 4380
rect 117810 3980 117840 4380
rect 117920 3980 117950 4380
rect 118030 3980 118060 4380
rect 118140 3980 118170 4380
rect 118250 3980 118280 4380
<< ndiff >>
rect 113540 6830 113620 6860
rect 113540 6390 113560 6830
rect 113600 6390 113620 6830
rect 113540 6360 113620 6390
rect 113650 6830 113730 6860
rect 113650 6390 113670 6830
rect 113710 6390 113730 6830
rect 113650 6360 113730 6390
rect 113760 6830 113840 6860
rect 113760 6390 113780 6830
rect 113820 6390 113840 6830
rect 113760 6360 113840 6390
rect 113870 6830 113950 6860
rect 113870 6390 113890 6830
rect 113930 6390 113950 6830
rect 113870 6360 113950 6390
rect 113980 6830 114060 6860
rect 113980 6390 114000 6830
rect 114040 6390 114060 6830
rect 113980 6360 114060 6390
rect 112060 5700 112140 5730
rect 112060 5460 112080 5700
rect 112120 5460 112140 5700
rect 112060 5430 112140 5460
rect 112170 5700 112250 5730
rect 112170 5460 112190 5700
rect 112230 5460 112250 5700
rect 112170 5430 112250 5460
rect 112280 5700 112360 5730
rect 112280 5460 112300 5700
rect 112340 5460 112360 5700
rect 112280 5430 112360 5460
rect 112390 5700 112470 5730
rect 112390 5460 112410 5700
rect 112450 5460 112470 5700
rect 112390 5430 112470 5460
rect 112500 5700 112580 5730
rect 112500 5460 112520 5700
rect 112560 5460 112580 5700
rect 112500 5430 112580 5460
rect 112610 5700 112690 5730
rect 112610 5460 112630 5700
rect 112670 5460 112690 5700
rect 112610 5430 112690 5460
rect 112720 5700 112800 5730
rect 112720 5460 112740 5700
rect 112780 5460 112800 5700
rect 112720 5430 112800 5460
rect 112830 5700 112910 5730
rect 112830 5460 112850 5700
rect 112890 5460 112910 5700
rect 112830 5430 112910 5460
rect 112940 5700 113020 5730
rect 112940 5460 112960 5700
rect 113000 5460 113020 5700
rect 112940 5430 113020 5460
rect 113050 5700 113130 5730
rect 113050 5460 113070 5700
rect 113110 5460 113130 5700
rect 113050 5430 113130 5460
rect 113160 5700 113240 5730
rect 113160 5460 113180 5700
rect 113220 5460 113240 5700
rect 113160 5430 113240 5460
rect 113270 5700 113350 5730
rect 113270 5460 113290 5700
rect 113330 5460 113350 5700
rect 113270 5430 113350 5460
rect 113380 5700 113460 5730
rect 113380 5460 113400 5700
rect 113440 5460 113460 5700
rect 113380 5430 113460 5460
rect 114140 5700 114220 5730
rect 114140 5460 114160 5700
rect 114200 5460 114220 5700
rect 114140 5430 114220 5460
rect 114250 5700 114330 5730
rect 114250 5460 114270 5700
rect 114310 5460 114330 5700
rect 114250 5430 114330 5460
rect 114360 5700 114440 5730
rect 114360 5460 114380 5700
rect 114420 5460 114440 5700
rect 114360 5430 114440 5460
rect 114470 5700 114550 5730
rect 114470 5460 114490 5700
rect 114530 5460 114550 5700
rect 114470 5430 114550 5460
rect 114580 5700 114660 5730
rect 114580 5460 114600 5700
rect 114640 5460 114660 5700
rect 114580 5430 114660 5460
rect 114690 5700 114770 5730
rect 114690 5460 114710 5700
rect 114750 5460 114770 5700
rect 114690 5430 114770 5460
rect 114800 5700 114880 5730
rect 114800 5460 114820 5700
rect 114860 5460 114880 5700
rect 114800 5430 114880 5460
rect 114910 5700 114990 5730
rect 114910 5460 114930 5700
rect 114970 5460 114990 5700
rect 114910 5430 114990 5460
rect 115020 5700 115100 5730
rect 115020 5460 115040 5700
rect 115080 5460 115100 5700
rect 115020 5430 115100 5460
rect 115130 5700 115210 5730
rect 115130 5460 115150 5700
rect 115190 5460 115210 5700
rect 115130 5430 115210 5460
rect 115240 5700 115320 5730
rect 115240 5460 115260 5700
rect 115300 5460 115320 5700
rect 115240 5430 115320 5460
rect 115350 5700 115430 5730
rect 115350 5460 115370 5700
rect 115410 5460 115430 5700
rect 115350 5430 115430 5460
rect 115460 5700 115540 5730
rect 115460 5460 115480 5700
rect 115520 5460 115540 5700
rect 115460 5430 115540 5460
rect 112060 3830 112140 3860
rect 112060 3590 112080 3830
rect 112120 3590 112140 3830
rect 112060 3560 112140 3590
rect 112170 3830 112250 3860
rect 112170 3590 112190 3830
rect 112230 3590 112250 3830
rect 112170 3560 112250 3590
rect 112280 3830 112360 3860
rect 112280 3590 112300 3830
rect 112340 3590 112360 3830
rect 112280 3560 112360 3590
rect 112390 3830 112470 3860
rect 112390 3590 112410 3830
rect 112450 3590 112470 3830
rect 112390 3560 112470 3590
rect 112500 3830 112580 3860
rect 112500 3590 112520 3830
rect 112560 3590 112580 3830
rect 112500 3560 112580 3590
rect 112610 3830 112690 3860
rect 112610 3590 112630 3830
rect 112670 3590 112690 3830
rect 112610 3560 112690 3590
rect 112720 3830 112800 3860
rect 112720 3590 112740 3830
rect 112780 3590 112800 3830
rect 112720 3560 112800 3590
rect 112830 3830 112910 3860
rect 112830 3590 112850 3830
rect 112890 3590 112910 3830
rect 112830 3560 112910 3590
rect 112940 3830 113020 3860
rect 112940 3590 112960 3830
rect 113000 3590 113020 3830
rect 112940 3560 113020 3590
rect 113050 3830 113130 3860
rect 113050 3590 113070 3830
rect 113110 3590 113130 3830
rect 113050 3560 113130 3590
rect 113160 3830 113240 3860
rect 113160 3590 113180 3830
rect 113220 3590 113240 3830
rect 113160 3560 113240 3590
rect 113270 3830 113350 3860
rect 113270 3590 113290 3830
rect 113330 3590 113350 3830
rect 113270 3560 113350 3590
rect 113380 3830 113460 3860
rect 113540 3830 113620 3860
rect 113380 3590 113400 3830
rect 113440 3590 113460 3830
rect 113540 3590 113560 3830
rect 113600 3590 113620 3830
rect 113380 3560 113460 3590
rect 113540 3560 113620 3590
rect 113650 3830 113730 3860
rect 113650 3590 113670 3830
rect 113710 3590 113730 3830
rect 113650 3560 113730 3590
rect 113760 3830 113840 3860
rect 113760 3590 113780 3830
rect 113820 3590 113840 3830
rect 113760 3560 113840 3590
rect 113870 3830 113950 3860
rect 113870 3590 113890 3830
rect 113930 3590 113950 3830
rect 113870 3560 113950 3590
rect 113980 3830 114060 3860
rect 114140 3830 114220 3860
rect 113980 3590 114000 3830
rect 114040 3590 114060 3830
rect 114140 3590 114160 3830
rect 114200 3590 114220 3830
rect 113980 3560 114060 3590
rect 114140 3560 114220 3590
rect 114250 3830 114330 3860
rect 114250 3590 114270 3830
rect 114310 3590 114330 3830
rect 114250 3560 114330 3590
rect 114360 3830 114440 3860
rect 114360 3590 114380 3830
rect 114420 3590 114440 3830
rect 114360 3560 114440 3590
rect 114470 3830 114550 3860
rect 114470 3590 114490 3830
rect 114530 3590 114550 3830
rect 114470 3560 114550 3590
rect 114580 3830 114660 3860
rect 114580 3590 114600 3830
rect 114640 3590 114660 3830
rect 114580 3560 114660 3590
rect 114690 3830 114770 3860
rect 114690 3590 114710 3830
rect 114750 3590 114770 3830
rect 114690 3560 114770 3590
rect 114800 3830 114880 3860
rect 114800 3590 114820 3830
rect 114860 3590 114880 3830
rect 114800 3560 114880 3590
rect 114910 3830 114990 3860
rect 114910 3590 114930 3830
rect 114970 3590 114990 3830
rect 114910 3560 114990 3590
rect 115020 3830 115100 3860
rect 115020 3590 115040 3830
rect 115080 3590 115100 3830
rect 115020 3560 115100 3590
rect 115130 3830 115210 3860
rect 115130 3590 115150 3830
rect 115190 3590 115210 3830
rect 115130 3560 115210 3590
rect 115240 3830 115320 3860
rect 115240 3590 115260 3830
rect 115300 3590 115320 3830
rect 115240 3560 115320 3590
rect 115350 3830 115430 3860
rect 115350 3590 115370 3830
rect 115410 3590 115430 3830
rect 115350 3560 115430 3590
rect 115460 3830 115540 3860
rect 115460 3590 115480 3830
rect 115520 3590 115540 3830
rect 115460 3560 115540 3590
rect 109240 3470 109320 3500
rect 109240 2930 109260 3470
rect 109300 2930 109320 3470
rect 109240 2900 109320 2930
rect 109350 3470 109430 3500
rect 109350 2930 109370 3470
rect 109410 2930 109430 3470
rect 109350 2900 109430 2930
rect 109460 3470 109540 3500
rect 109460 2930 109480 3470
rect 109520 2930 109540 3470
rect 109460 2900 109540 2930
rect 109570 3470 109650 3500
rect 109570 2930 109590 3470
rect 109630 2930 109650 3470
rect 109570 2900 109650 2930
rect 109680 3470 109760 3500
rect 109680 2930 109700 3470
rect 109740 2930 109760 3470
rect 109680 2900 109760 2930
rect 109790 3470 109870 3500
rect 109790 2930 109810 3470
rect 109850 2930 109870 3470
rect 109790 2900 109870 2930
rect 109900 3470 109980 3500
rect 109900 2930 109920 3470
rect 109960 2930 109980 3470
rect 109900 2900 109980 2930
rect 110010 3470 110090 3500
rect 110010 2930 110030 3470
rect 110070 2930 110090 3470
rect 110010 2900 110090 2930
rect 110120 3470 110200 3500
rect 110120 2930 110140 3470
rect 110180 2930 110200 3470
rect 110120 2900 110200 2930
rect 110230 3470 110310 3500
rect 110230 2930 110250 3470
rect 110290 2930 110310 3470
rect 110230 2900 110310 2930
rect 110340 3470 110420 3500
rect 110340 2930 110360 3470
rect 110400 2930 110420 3470
rect 110340 2900 110420 2930
rect 110450 3470 110530 3500
rect 110450 2930 110470 3470
rect 110510 2930 110530 3470
rect 110450 2900 110530 2930
rect 110560 3470 110640 3500
rect 110560 2930 110580 3470
rect 110620 2930 110640 3470
rect 116960 3470 117040 3500
rect 110560 2900 110640 2930
rect 116960 2930 116980 3470
rect 117020 2930 117040 3470
rect 116960 2900 117040 2930
rect 117070 3470 117150 3500
rect 117070 2930 117090 3470
rect 117130 2930 117150 3470
rect 117070 2900 117150 2930
rect 117180 3470 117260 3500
rect 117180 2930 117200 3470
rect 117240 2930 117260 3470
rect 117180 2900 117260 2930
rect 117290 3470 117370 3500
rect 117290 2930 117310 3470
rect 117350 2930 117370 3470
rect 117290 2900 117370 2930
rect 117400 3470 117480 3500
rect 117400 2930 117420 3470
rect 117460 2930 117480 3470
rect 117400 2900 117480 2930
rect 117510 3470 117590 3500
rect 117510 2930 117530 3470
rect 117570 2930 117590 3470
rect 117510 2900 117590 2930
rect 117620 3470 117700 3500
rect 117620 2930 117640 3470
rect 117680 2930 117700 3470
rect 117620 2900 117700 2930
rect 117730 3470 117810 3500
rect 117730 2930 117750 3470
rect 117790 2930 117810 3470
rect 117730 2900 117810 2930
rect 117840 3470 117920 3500
rect 117840 2930 117860 3470
rect 117900 2930 117920 3470
rect 117840 2900 117920 2930
rect 117950 3470 118030 3500
rect 117950 2930 117970 3470
rect 118010 2930 118030 3470
rect 117950 2900 118030 2930
rect 118060 3470 118140 3500
rect 118060 2930 118080 3470
rect 118120 2930 118140 3470
rect 118060 2900 118140 2930
rect 118170 3470 118250 3500
rect 118170 2930 118190 3470
rect 118230 2930 118250 3470
rect 118170 2900 118250 2930
rect 118280 3470 118360 3500
rect 118280 2930 118300 3470
rect 118340 2930 118360 3470
rect 118280 2900 118360 2930
rect 112440 1580 112520 1610
rect 109300 1350 109380 1380
rect 109300 10 109320 1350
rect 109360 10 109380 1350
rect 109300 -20 109380 10
rect 109500 1350 109580 1380
rect 109500 10 109520 1350
rect 109560 10 109580 1350
rect 109500 -20 109580 10
rect 109700 1350 109780 1380
rect 109700 10 109720 1350
rect 109760 10 109780 1350
rect 109700 -20 109780 10
rect 109900 1350 109980 1380
rect 109900 10 109920 1350
rect 109960 10 109980 1350
rect 109900 -20 109980 10
rect 110100 1350 110180 1380
rect 110100 10 110120 1350
rect 110160 10 110180 1350
rect 110100 -20 110180 10
rect 110300 1350 110380 1380
rect 110300 10 110320 1350
rect 110360 10 110380 1350
rect 110300 -20 110380 10
rect 110500 1350 110580 1380
rect 110500 10 110520 1350
rect 110560 10 110580 1350
rect 112440 1140 112460 1580
rect 112500 1140 112520 1580
rect 112440 1110 112520 1140
rect 112550 1580 112630 1610
rect 112550 1140 112570 1580
rect 112610 1140 112630 1580
rect 112550 1110 112630 1140
rect 112660 1580 112740 1610
rect 112660 1140 112680 1580
rect 112720 1140 112740 1580
rect 112660 1110 112740 1140
rect 112770 1580 112850 1610
rect 112770 1140 112790 1580
rect 112830 1140 112850 1580
rect 112770 1110 112850 1140
rect 112880 1580 112960 1610
rect 112880 1140 112900 1580
rect 112940 1140 112960 1580
rect 112880 1110 112960 1140
rect 112990 1580 113070 1610
rect 112990 1140 113010 1580
rect 113050 1140 113070 1580
rect 112990 1110 113070 1140
rect 113100 1580 113180 1610
rect 113100 1140 113120 1580
rect 113160 1140 113180 1580
rect 113100 1110 113180 1140
rect 113210 1580 113290 1610
rect 113210 1140 113230 1580
rect 113270 1140 113290 1580
rect 113210 1110 113290 1140
rect 113320 1580 113400 1610
rect 113320 1140 113340 1580
rect 113380 1140 113400 1580
rect 113320 1110 113400 1140
rect 113430 1580 113510 1610
rect 113430 1140 113450 1580
rect 113490 1140 113510 1580
rect 113430 1110 113510 1140
rect 113540 1580 113620 1610
rect 113540 1140 113560 1580
rect 113600 1140 113620 1580
rect 113540 1110 113620 1140
rect 113650 1580 113730 1610
rect 113650 1140 113670 1580
rect 113710 1140 113730 1580
rect 113650 1110 113730 1140
rect 113760 1580 113840 1610
rect 113760 1140 113780 1580
rect 113820 1140 113840 1580
rect 113760 1110 113840 1140
rect 113870 1580 113950 1610
rect 113870 1140 113890 1580
rect 113930 1140 113950 1580
rect 113870 1110 113950 1140
rect 113980 1580 114060 1610
rect 113980 1140 114000 1580
rect 114040 1140 114060 1580
rect 113980 1110 114060 1140
rect 114090 1580 114170 1610
rect 114090 1140 114110 1580
rect 114150 1140 114170 1580
rect 114090 1110 114170 1140
rect 114200 1580 114280 1610
rect 114200 1140 114220 1580
rect 114260 1140 114280 1580
rect 114200 1110 114280 1140
rect 114310 1580 114390 1610
rect 114310 1140 114330 1580
rect 114370 1140 114390 1580
rect 114310 1110 114390 1140
rect 114420 1580 114500 1610
rect 114420 1140 114440 1580
rect 114480 1140 114500 1580
rect 114420 1110 114500 1140
rect 114530 1580 114610 1610
rect 114530 1140 114550 1580
rect 114590 1140 114610 1580
rect 114530 1110 114610 1140
rect 114640 1580 114720 1610
rect 114640 1140 114660 1580
rect 114700 1140 114720 1580
rect 114640 1110 114720 1140
rect 114750 1580 114830 1610
rect 114750 1140 114770 1580
rect 114810 1140 114830 1580
rect 114750 1110 114830 1140
rect 114860 1580 114940 1610
rect 114860 1140 114880 1580
rect 114920 1140 114940 1580
rect 114860 1110 114940 1140
rect 114970 1580 115050 1610
rect 114970 1140 114990 1580
rect 115030 1140 115050 1580
rect 114970 1110 115050 1140
rect 117020 1350 117100 1380
rect 110500 -20 110580 10
rect 113430 70 113510 100
rect 113430 -170 113450 70
rect 113490 -170 113510 70
rect 113430 -200 113510 -170
rect 113540 70 113620 100
rect 113540 -170 113560 70
rect 113600 -170 113620 70
rect 113540 -200 113620 -170
rect 113650 70 113730 100
rect 113650 -170 113670 70
rect 113710 -170 113730 70
rect 113650 -200 113730 -170
rect 113760 70 113840 100
rect 113760 -170 113780 70
rect 113820 -170 113840 70
rect 113760 -200 113840 -170
rect 113870 70 113950 100
rect 113870 -170 113890 70
rect 113930 -170 113950 70
rect 113870 -200 113950 -170
rect 113980 70 114060 100
rect 113980 -170 114000 70
rect 114040 -170 114060 70
rect 113980 -200 114060 -170
rect 114090 70 114170 100
rect 114090 -170 114110 70
rect 114150 -170 114170 70
rect 117020 10 117040 1350
rect 117080 10 117100 1350
rect 117020 -20 117100 10
rect 117220 1350 117300 1380
rect 117220 10 117240 1350
rect 117280 10 117300 1350
rect 117220 -20 117300 10
rect 117420 1350 117500 1380
rect 117420 10 117440 1350
rect 117480 10 117500 1350
rect 117420 -20 117500 10
rect 117620 1350 117700 1380
rect 117620 10 117640 1350
rect 117680 10 117700 1350
rect 117620 -20 117700 10
rect 117820 1350 117900 1380
rect 117820 10 117840 1350
rect 117880 10 117900 1350
rect 117820 -20 117900 10
rect 118020 1350 118100 1380
rect 118020 10 118040 1350
rect 118080 10 118100 1350
rect 118020 -20 118100 10
rect 118220 1350 118300 1380
rect 118220 10 118240 1350
rect 118280 10 118300 1350
rect 118220 -20 118300 10
rect 114090 -200 114170 -170
rect 113420 -450 113500 -420
rect 113420 -690 113440 -450
rect 113480 -690 113500 -450
rect 113420 -720 113500 -690
rect 114100 -450 114180 -420
rect 114100 -690 114120 -450
rect 114160 -690 114180 -450
rect 114100 -720 114180 -690
<< pdiff >>
rect 109300 9770 109380 9800
rect 109300 9130 109320 9770
rect 109360 9130 109380 9770
rect 109300 9100 109380 9130
rect 109420 9770 109500 9800
rect 109420 9130 109440 9770
rect 109480 9130 109500 9770
rect 109420 9100 109500 9130
rect 109540 9770 109620 9800
rect 109540 9130 109560 9770
rect 109600 9130 109620 9770
rect 109540 9100 109620 9130
rect 109660 9770 109740 9800
rect 109660 9130 109680 9770
rect 109720 9130 109740 9770
rect 109660 9100 109740 9130
rect 109780 9770 109860 9800
rect 109780 9130 109800 9770
rect 109840 9130 109860 9770
rect 109780 9100 109860 9130
rect 109900 9770 109980 9800
rect 109900 9130 109920 9770
rect 109960 9130 109980 9770
rect 109900 9100 109980 9130
rect 110020 9770 110100 9800
rect 110020 9130 110040 9770
rect 110080 9130 110100 9770
rect 110020 9100 110100 9130
rect 110140 9770 110220 9800
rect 110140 9130 110160 9770
rect 110200 9130 110220 9770
rect 110140 9100 110220 9130
rect 110260 9770 110340 9800
rect 110260 9130 110280 9770
rect 110320 9130 110340 9770
rect 110260 9100 110340 9130
rect 110380 9770 110460 9800
rect 110380 9130 110400 9770
rect 110440 9130 110460 9770
rect 110380 9100 110460 9130
rect 110500 9770 110580 9800
rect 110500 9130 110520 9770
rect 110560 9130 110580 9770
rect 110500 9100 110580 9130
rect 110620 9770 110700 9800
rect 110620 9130 110640 9770
rect 110680 9130 110700 9770
rect 110620 9100 110700 9130
rect 110740 9770 110820 9800
rect 110740 9130 110760 9770
rect 110800 9130 110820 9770
rect 116780 9770 116860 9800
rect 110740 9100 110820 9130
rect 111970 9470 112050 9500
rect 111970 8830 111990 9470
rect 112030 8830 112050 9470
rect 111970 8800 112050 8830
rect 112090 9470 112170 9500
rect 112090 8830 112110 9470
rect 112150 8830 112170 9470
rect 112090 8800 112170 8830
rect 112210 9470 112290 9500
rect 112210 8830 112230 9470
rect 112270 8830 112290 9470
rect 112210 8800 112290 8830
rect 112330 9470 112410 9500
rect 112330 8830 112350 9470
rect 112390 8830 112410 9470
rect 114250 9470 114330 9500
rect 112330 8800 112410 8830
rect 112910 9130 112990 9160
rect 112910 8830 112930 9130
rect 112970 8830 112990 9130
rect 112910 8800 112990 8830
rect 113030 9130 113110 9160
rect 113030 8830 113050 9130
rect 113090 8830 113110 9130
rect 113030 8800 113110 8830
rect 113150 9130 113230 9160
rect 113150 8830 113170 9130
rect 113210 8830 113230 9130
rect 113150 8800 113230 8830
rect 113270 9130 113350 9160
rect 113270 8830 113290 9130
rect 113330 8830 113350 9130
rect 113270 8800 113350 8830
rect 114250 8830 114270 9470
rect 114310 8830 114330 9470
rect 114250 8800 114330 8830
rect 114370 9470 114450 9500
rect 114370 8830 114390 9470
rect 114430 8830 114450 9470
rect 114370 8800 114450 8830
rect 114490 9470 114570 9500
rect 114490 8830 114510 9470
rect 114550 8830 114570 9470
rect 114490 8800 114570 8830
rect 114610 9470 114690 9500
rect 114610 8830 114630 9470
rect 114670 8830 114690 9470
rect 114610 8800 114690 8830
rect 115190 9470 115270 9500
rect 115190 8830 115210 9470
rect 115250 8830 115270 9470
rect 115190 8800 115270 8830
rect 115310 9470 115390 9500
rect 115310 8830 115330 9470
rect 115370 8830 115390 9470
rect 115310 8800 115390 8830
rect 115430 9470 115510 9500
rect 115430 8830 115450 9470
rect 115490 8830 115510 9470
rect 115430 8800 115510 8830
rect 115550 9470 115630 9500
rect 115550 8830 115570 9470
rect 115610 8830 115630 9470
rect 116780 9130 116800 9770
rect 116840 9130 116860 9770
rect 116780 9100 116860 9130
rect 116900 9770 116980 9800
rect 116900 9130 116920 9770
rect 116960 9130 116980 9770
rect 116900 9100 116980 9130
rect 117020 9770 117100 9800
rect 117020 9130 117040 9770
rect 117080 9130 117100 9770
rect 117020 9100 117100 9130
rect 117140 9770 117220 9800
rect 117140 9130 117160 9770
rect 117200 9130 117220 9770
rect 117140 9100 117220 9130
rect 117260 9770 117340 9800
rect 117260 9130 117280 9770
rect 117320 9130 117340 9770
rect 117260 9100 117340 9130
rect 117380 9770 117460 9800
rect 117380 9130 117400 9770
rect 117440 9130 117460 9770
rect 117380 9100 117460 9130
rect 117500 9770 117580 9800
rect 117500 9130 117520 9770
rect 117560 9130 117580 9770
rect 117500 9100 117580 9130
rect 117620 9770 117700 9800
rect 117620 9130 117640 9770
rect 117680 9130 117700 9770
rect 117620 9100 117700 9130
rect 117740 9770 117820 9800
rect 117740 9130 117760 9770
rect 117800 9130 117820 9770
rect 117740 9100 117820 9130
rect 117860 9770 117940 9800
rect 117860 9130 117880 9770
rect 117920 9130 117940 9770
rect 117860 9100 117940 9130
rect 117980 9770 118060 9800
rect 117980 9130 118000 9770
rect 118040 9130 118060 9770
rect 117980 9100 118060 9130
rect 118100 9770 118180 9800
rect 118100 9130 118120 9770
rect 118160 9130 118180 9770
rect 118100 9100 118180 9130
rect 118220 9770 118300 9800
rect 118220 9130 118240 9770
rect 118280 9130 118300 9770
rect 118220 9100 118300 9130
rect 115550 8800 115630 8830
rect 109180 8250 109260 8280
rect 109180 7610 109200 8250
rect 109240 7610 109260 8250
rect 109180 7580 109260 7610
rect 109300 8250 109380 8280
rect 109300 7610 109320 8250
rect 109360 7610 109380 8250
rect 109300 7580 109380 7610
rect 109420 8250 109500 8280
rect 109420 7610 109440 8250
rect 109480 7610 109500 8250
rect 109420 7580 109500 7610
rect 109540 8250 109620 8280
rect 109540 7610 109560 8250
rect 109600 7610 109620 8250
rect 109540 7580 109620 7610
rect 109660 8250 109740 8280
rect 109660 7610 109680 8250
rect 109720 7610 109740 8250
rect 109660 7580 109740 7610
rect 109780 8250 109860 8280
rect 109780 7610 109800 8250
rect 109840 7610 109860 8250
rect 109780 7580 109860 7610
rect 109900 8250 109980 8280
rect 109900 7610 109920 8250
rect 109960 7610 109980 8250
rect 109900 7580 109980 7610
rect 110020 8250 110100 8280
rect 110020 7610 110040 8250
rect 110080 7610 110100 8250
rect 110020 7580 110100 7610
rect 110140 8250 110220 8280
rect 110140 7610 110160 8250
rect 110200 7610 110220 8250
rect 110140 7580 110220 7610
rect 110260 8250 110340 8280
rect 110260 7610 110280 8250
rect 110320 7610 110340 8250
rect 110260 7580 110340 7610
rect 110380 8250 110460 8280
rect 110380 7610 110400 8250
rect 110440 7610 110460 8250
rect 110380 7580 110460 7610
rect 110500 8250 110580 8280
rect 110500 7610 110520 8250
rect 110560 7610 110580 8250
rect 110500 7580 110580 7610
rect 110620 8250 110700 8280
rect 110620 7610 110640 8250
rect 110680 7610 110700 8250
rect 116900 8250 116980 8280
rect 110620 7580 110700 7610
rect 113020 8040 113100 8070
rect 113020 7600 113040 8040
rect 113080 7600 113100 8040
rect 113020 7570 113100 7600
rect 113130 8040 113210 8070
rect 113130 7600 113150 8040
rect 113190 7600 113210 8040
rect 113130 7570 113210 7600
rect 113240 8040 113320 8070
rect 113240 7600 113260 8040
rect 113300 7600 113320 8040
rect 113240 7570 113320 7600
rect 113350 8040 113430 8070
rect 113350 7600 113370 8040
rect 113410 7600 113430 8040
rect 113350 7570 113430 7600
rect 113460 8040 113540 8070
rect 113460 7600 113480 8040
rect 113520 7600 113540 8040
rect 113460 7570 113540 7600
rect 113570 8040 113650 8070
rect 113570 7600 113590 8040
rect 113630 7600 113650 8040
rect 113570 7570 113650 7600
rect 113680 8040 113760 8070
rect 113840 8040 113920 8070
rect 113680 7600 113700 8040
rect 113740 7600 113760 8040
rect 113840 7600 113860 8040
rect 113900 7600 113920 8040
rect 113680 7570 113760 7600
rect 113840 7570 113920 7600
rect 113950 8040 114030 8070
rect 113950 7600 113970 8040
rect 114010 7600 114030 8040
rect 113950 7570 114030 7600
rect 114060 8040 114140 8070
rect 114060 7600 114080 8040
rect 114120 7600 114140 8040
rect 114060 7570 114140 7600
rect 114170 8040 114250 8070
rect 114170 7600 114190 8040
rect 114230 7600 114250 8040
rect 114170 7570 114250 7600
rect 114280 8040 114360 8070
rect 114280 7600 114300 8040
rect 114340 7600 114360 8040
rect 114280 7570 114360 7600
rect 114390 8040 114470 8070
rect 114390 7600 114410 8040
rect 114450 7600 114470 8040
rect 114390 7570 114470 7600
rect 114500 8040 114580 8070
rect 114500 7600 114520 8040
rect 114560 7600 114580 8040
rect 114500 7570 114580 7600
rect 116900 7610 116920 8250
rect 116960 7610 116980 8250
rect 116900 7580 116980 7610
rect 117020 8250 117100 8280
rect 117020 7610 117040 8250
rect 117080 7610 117100 8250
rect 117020 7580 117100 7610
rect 117140 8250 117220 8280
rect 117140 7610 117160 8250
rect 117200 7610 117220 8250
rect 117140 7580 117220 7610
rect 117260 8250 117340 8280
rect 117260 7610 117280 8250
rect 117320 7610 117340 8250
rect 117260 7580 117340 7610
rect 117380 8250 117460 8280
rect 117380 7610 117400 8250
rect 117440 7610 117460 8250
rect 117380 7580 117460 7610
rect 117500 8250 117580 8280
rect 117500 7610 117520 8250
rect 117560 7610 117580 8250
rect 117500 7580 117580 7610
rect 117620 8250 117700 8280
rect 117620 7610 117640 8250
rect 117680 7610 117700 8250
rect 117620 7580 117700 7610
rect 117740 8250 117820 8280
rect 117740 7610 117760 8250
rect 117800 7610 117820 8250
rect 117740 7580 117820 7610
rect 117860 8250 117940 8280
rect 117860 7610 117880 8250
rect 117920 7610 117940 8250
rect 117860 7580 117940 7610
rect 117980 8250 118060 8280
rect 117980 7610 118000 8250
rect 118040 7610 118060 8250
rect 117980 7580 118060 7610
rect 118100 8250 118180 8280
rect 118100 7610 118120 8250
rect 118160 7610 118180 8250
rect 118100 7580 118180 7610
rect 118220 8250 118300 8280
rect 118220 7610 118240 8250
rect 118280 7610 118300 8250
rect 118220 7580 118300 7610
rect 118340 8250 118420 8280
rect 118340 7610 118360 8250
rect 118400 7610 118420 8250
rect 118340 7580 118420 7610
rect 109240 6900 109320 6930
rect 109240 5760 109260 6900
rect 109300 5760 109320 6900
rect 109240 5730 109320 5760
rect 109350 6900 109430 6930
rect 109350 5760 109370 6900
rect 109410 5760 109430 6900
rect 109350 5730 109430 5760
rect 109460 6900 109540 6930
rect 109460 5760 109480 6900
rect 109520 5760 109540 6900
rect 109460 5730 109540 5760
rect 109570 6900 109650 6930
rect 109570 5760 109590 6900
rect 109630 5760 109650 6900
rect 109570 5730 109650 5760
rect 109680 6900 109760 6930
rect 109680 5760 109700 6900
rect 109740 5760 109760 6900
rect 109680 5730 109760 5760
rect 109790 6900 109870 6930
rect 109790 5760 109810 6900
rect 109850 5760 109870 6900
rect 109790 5730 109870 5760
rect 109900 6900 109980 6930
rect 109900 5760 109920 6900
rect 109960 5760 109980 6900
rect 109900 5730 109980 5760
rect 110010 6900 110090 6930
rect 110010 5760 110030 6900
rect 110070 5760 110090 6900
rect 110010 5730 110090 5760
rect 110120 6900 110200 6930
rect 110120 5760 110140 6900
rect 110180 5760 110200 6900
rect 110120 5730 110200 5760
rect 110230 6900 110310 6930
rect 110230 5760 110250 6900
rect 110290 5760 110310 6900
rect 110230 5730 110310 5760
rect 110340 6900 110420 6930
rect 110340 5760 110360 6900
rect 110400 5760 110420 6900
rect 110340 5730 110420 5760
rect 110450 6900 110530 6930
rect 110450 5760 110470 6900
rect 110510 5760 110530 6900
rect 110450 5730 110530 5760
rect 110560 6900 110640 6930
rect 110560 5760 110580 6900
rect 110620 5760 110640 6900
rect 116960 6900 117040 6930
rect 116960 5760 116980 6900
rect 117020 5760 117040 6900
rect 110560 5730 110640 5760
rect 116960 5730 117040 5760
rect 117070 6900 117150 6930
rect 117070 5760 117090 6900
rect 117130 5760 117150 6900
rect 117070 5730 117150 5760
rect 117180 6900 117260 6930
rect 117180 5760 117200 6900
rect 117240 5760 117260 6900
rect 117180 5730 117260 5760
rect 117290 6900 117370 6930
rect 117290 5760 117310 6900
rect 117350 5760 117370 6900
rect 117290 5730 117370 5760
rect 117400 6900 117480 6930
rect 117400 5760 117420 6900
rect 117460 5760 117480 6900
rect 117400 5730 117480 5760
rect 117510 6900 117590 6930
rect 117510 5760 117530 6900
rect 117570 5760 117590 6900
rect 117510 5730 117590 5760
rect 117620 6900 117700 6930
rect 117620 5760 117640 6900
rect 117680 5760 117700 6900
rect 117620 5730 117700 5760
rect 117730 6900 117810 6930
rect 117730 5760 117750 6900
rect 117790 5760 117810 6900
rect 117730 5730 117810 5760
rect 117840 6900 117920 6930
rect 117840 5760 117860 6900
rect 117900 5760 117920 6900
rect 117840 5730 117920 5760
rect 117950 6900 118030 6930
rect 117950 5760 117970 6900
rect 118010 5760 118030 6900
rect 117950 5730 118030 5760
rect 118060 6900 118140 6930
rect 118060 5760 118080 6900
rect 118120 5760 118140 6900
rect 118060 5730 118140 5760
rect 118170 6900 118250 6930
rect 118170 5760 118190 6900
rect 118230 5760 118250 6900
rect 118170 5730 118250 5760
rect 118280 6900 118360 6930
rect 118280 5760 118300 6900
rect 118340 5760 118360 6900
rect 118280 5730 118360 5760
rect 109240 4350 109320 4380
rect 109240 4010 109260 4350
rect 109300 4010 109320 4350
rect 109240 3980 109320 4010
rect 109350 4350 109430 4380
rect 109350 4010 109370 4350
rect 109410 4010 109430 4350
rect 109350 3980 109430 4010
rect 109460 4350 109540 4380
rect 109460 4010 109480 4350
rect 109520 4010 109540 4350
rect 109460 3980 109540 4010
rect 109570 4350 109650 4380
rect 109570 4010 109590 4350
rect 109630 4010 109650 4350
rect 109570 3980 109650 4010
rect 109680 4350 109760 4380
rect 109680 4010 109700 4350
rect 109740 4010 109760 4350
rect 109680 3980 109760 4010
rect 109790 4350 109870 4380
rect 109790 4010 109810 4350
rect 109850 4010 109870 4350
rect 109790 3980 109870 4010
rect 109900 4350 109980 4380
rect 109900 4010 109920 4350
rect 109960 4010 109980 4350
rect 109900 3980 109980 4010
rect 110010 4350 110090 4380
rect 110010 4010 110030 4350
rect 110070 4010 110090 4350
rect 110010 3980 110090 4010
rect 110120 4350 110200 4380
rect 110120 4010 110140 4350
rect 110180 4010 110200 4350
rect 110120 3980 110200 4010
rect 110230 4350 110310 4380
rect 110230 4010 110250 4350
rect 110290 4010 110310 4350
rect 110230 3980 110310 4010
rect 110340 4350 110420 4380
rect 110340 4010 110360 4350
rect 110400 4010 110420 4350
rect 110340 3980 110420 4010
rect 110450 4350 110530 4380
rect 110450 4010 110470 4350
rect 110510 4010 110530 4350
rect 110450 3980 110530 4010
rect 110560 4350 110640 4380
rect 110560 4010 110580 4350
rect 110620 4010 110640 4350
rect 116960 4350 117040 4380
rect 110560 3980 110640 4010
rect 116960 4010 116980 4350
rect 117020 4010 117040 4350
rect 116960 3980 117040 4010
rect 117070 4350 117150 4380
rect 117070 4010 117090 4350
rect 117130 4010 117150 4350
rect 117070 3980 117150 4010
rect 117180 4350 117260 4380
rect 117180 4010 117200 4350
rect 117240 4010 117260 4350
rect 117180 3980 117260 4010
rect 117290 4350 117370 4380
rect 117290 4010 117310 4350
rect 117350 4010 117370 4350
rect 117290 3980 117370 4010
rect 117400 4350 117480 4380
rect 117400 4010 117420 4350
rect 117460 4010 117480 4350
rect 117400 3980 117480 4010
rect 117510 4350 117590 4380
rect 117510 4010 117530 4350
rect 117570 4010 117590 4350
rect 117510 3980 117590 4010
rect 117620 4350 117700 4380
rect 117620 4010 117640 4350
rect 117680 4010 117700 4350
rect 117620 3980 117700 4010
rect 117730 4350 117810 4380
rect 117730 4010 117750 4350
rect 117790 4010 117810 4350
rect 117730 3980 117810 4010
rect 117840 4350 117920 4380
rect 117840 4010 117860 4350
rect 117900 4010 117920 4350
rect 117840 3980 117920 4010
rect 117950 4350 118030 4380
rect 117950 4010 117970 4350
rect 118010 4010 118030 4350
rect 117950 3980 118030 4010
rect 118060 4350 118140 4380
rect 118060 4010 118080 4350
rect 118120 4010 118140 4350
rect 118060 3980 118140 4010
rect 118170 4350 118250 4380
rect 118170 4010 118190 4350
rect 118230 4010 118250 4350
rect 118170 3980 118250 4010
rect 118280 4350 118360 4380
rect 118280 4010 118300 4350
rect 118340 4010 118360 4350
rect 118280 3980 118360 4010
<< ndiffc >>
rect 113560 6390 113600 6830
rect 113670 6390 113710 6830
rect 113780 6390 113820 6830
rect 113890 6390 113930 6830
rect 114000 6390 114040 6830
rect 112080 5460 112120 5700
rect 112190 5460 112230 5700
rect 112300 5460 112340 5700
rect 112410 5460 112450 5700
rect 112520 5460 112560 5700
rect 112630 5460 112670 5700
rect 112740 5460 112780 5700
rect 112850 5460 112890 5700
rect 112960 5460 113000 5700
rect 113070 5460 113110 5700
rect 113180 5460 113220 5700
rect 113290 5460 113330 5700
rect 113400 5460 113440 5700
rect 114160 5460 114200 5700
rect 114270 5460 114310 5700
rect 114380 5460 114420 5700
rect 114490 5460 114530 5700
rect 114600 5460 114640 5700
rect 114710 5460 114750 5700
rect 114820 5460 114860 5700
rect 114930 5460 114970 5700
rect 115040 5460 115080 5700
rect 115150 5460 115190 5700
rect 115260 5460 115300 5700
rect 115370 5460 115410 5700
rect 115480 5460 115520 5700
rect 112080 3590 112120 3830
rect 112190 3590 112230 3830
rect 112300 3590 112340 3830
rect 112410 3590 112450 3830
rect 112520 3590 112560 3830
rect 112630 3590 112670 3830
rect 112740 3590 112780 3830
rect 112850 3590 112890 3830
rect 112960 3590 113000 3830
rect 113070 3590 113110 3830
rect 113180 3590 113220 3830
rect 113290 3590 113330 3830
rect 113400 3590 113440 3830
rect 113560 3590 113600 3830
rect 113670 3590 113710 3830
rect 113780 3590 113820 3830
rect 113890 3590 113930 3830
rect 114000 3590 114040 3830
rect 114160 3590 114200 3830
rect 114270 3590 114310 3830
rect 114380 3590 114420 3830
rect 114490 3590 114530 3830
rect 114600 3590 114640 3830
rect 114710 3590 114750 3830
rect 114820 3590 114860 3830
rect 114930 3590 114970 3830
rect 115040 3590 115080 3830
rect 115150 3590 115190 3830
rect 115260 3590 115300 3830
rect 115370 3590 115410 3830
rect 115480 3590 115520 3830
rect 109260 2930 109300 3470
rect 109370 2930 109410 3470
rect 109480 2930 109520 3470
rect 109590 2930 109630 3470
rect 109700 2930 109740 3470
rect 109810 2930 109850 3470
rect 109920 2930 109960 3470
rect 110030 2930 110070 3470
rect 110140 2930 110180 3470
rect 110250 2930 110290 3470
rect 110360 2930 110400 3470
rect 110470 2930 110510 3470
rect 110580 2930 110620 3470
rect 116980 2930 117020 3470
rect 117090 2930 117130 3470
rect 117200 2930 117240 3470
rect 117310 2930 117350 3470
rect 117420 2930 117460 3470
rect 117530 2930 117570 3470
rect 117640 2930 117680 3470
rect 117750 2930 117790 3470
rect 117860 2930 117900 3470
rect 117970 2930 118010 3470
rect 118080 2930 118120 3470
rect 118190 2930 118230 3470
rect 118300 2930 118340 3470
rect 109320 10 109360 1350
rect 109520 10 109560 1350
rect 109720 10 109760 1350
rect 109920 10 109960 1350
rect 110120 10 110160 1350
rect 110320 10 110360 1350
rect 110520 10 110560 1350
rect 112460 1140 112500 1580
rect 112570 1140 112610 1580
rect 112680 1140 112720 1580
rect 112790 1140 112830 1580
rect 112900 1140 112940 1580
rect 113010 1140 113050 1580
rect 113120 1140 113160 1580
rect 113230 1140 113270 1580
rect 113340 1140 113380 1580
rect 113450 1140 113490 1580
rect 113560 1140 113600 1580
rect 113670 1140 113710 1580
rect 113780 1140 113820 1580
rect 113890 1140 113930 1580
rect 114000 1140 114040 1580
rect 114110 1140 114150 1580
rect 114220 1140 114260 1580
rect 114330 1140 114370 1580
rect 114440 1140 114480 1580
rect 114550 1140 114590 1580
rect 114660 1140 114700 1580
rect 114770 1140 114810 1580
rect 114880 1140 114920 1580
rect 114990 1140 115030 1580
rect 113450 -170 113490 70
rect 113560 -170 113600 70
rect 113670 -170 113710 70
rect 113780 -170 113820 70
rect 113890 -170 113930 70
rect 114000 -170 114040 70
rect 114110 -170 114150 70
rect 117040 10 117080 1350
rect 117240 10 117280 1350
rect 117440 10 117480 1350
rect 117640 10 117680 1350
rect 117840 10 117880 1350
rect 118040 10 118080 1350
rect 118240 10 118280 1350
rect 113440 -690 113480 -450
rect 114120 -690 114160 -450
<< pdiffc >>
rect 109320 9130 109360 9770
rect 109440 9130 109480 9770
rect 109560 9130 109600 9770
rect 109680 9130 109720 9770
rect 109800 9130 109840 9770
rect 109920 9130 109960 9770
rect 110040 9130 110080 9770
rect 110160 9130 110200 9770
rect 110280 9130 110320 9770
rect 110400 9130 110440 9770
rect 110520 9130 110560 9770
rect 110640 9130 110680 9770
rect 110760 9130 110800 9770
rect 111990 8830 112030 9470
rect 112110 8830 112150 9470
rect 112230 8830 112270 9470
rect 112350 8830 112390 9470
rect 112930 8830 112970 9130
rect 113050 8830 113090 9130
rect 113170 8830 113210 9130
rect 113290 8830 113330 9130
rect 114270 8830 114310 9470
rect 114390 8830 114430 9470
rect 114510 8830 114550 9470
rect 114630 8830 114670 9470
rect 115210 8830 115250 9470
rect 115330 8830 115370 9470
rect 115450 8830 115490 9470
rect 115570 8830 115610 9470
rect 116800 9130 116840 9770
rect 116920 9130 116960 9770
rect 117040 9130 117080 9770
rect 117160 9130 117200 9770
rect 117280 9130 117320 9770
rect 117400 9130 117440 9770
rect 117520 9130 117560 9770
rect 117640 9130 117680 9770
rect 117760 9130 117800 9770
rect 117880 9130 117920 9770
rect 118000 9130 118040 9770
rect 118120 9130 118160 9770
rect 118240 9130 118280 9770
rect 109200 7610 109240 8250
rect 109320 7610 109360 8250
rect 109440 7610 109480 8250
rect 109560 7610 109600 8250
rect 109680 7610 109720 8250
rect 109800 7610 109840 8250
rect 109920 7610 109960 8250
rect 110040 7610 110080 8250
rect 110160 7610 110200 8250
rect 110280 7610 110320 8250
rect 110400 7610 110440 8250
rect 110520 7610 110560 8250
rect 110640 7610 110680 8250
rect 113040 7600 113080 8040
rect 113150 7600 113190 8040
rect 113260 7600 113300 8040
rect 113370 7600 113410 8040
rect 113480 7600 113520 8040
rect 113590 7600 113630 8040
rect 113700 7600 113740 8040
rect 113860 7600 113900 8040
rect 113970 7600 114010 8040
rect 114080 7600 114120 8040
rect 114190 7600 114230 8040
rect 114300 7600 114340 8040
rect 114410 7600 114450 8040
rect 114520 7600 114560 8040
rect 116920 7610 116960 8250
rect 117040 7610 117080 8250
rect 117160 7610 117200 8250
rect 117280 7610 117320 8250
rect 117400 7610 117440 8250
rect 117520 7610 117560 8250
rect 117640 7610 117680 8250
rect 117760 7610 117800 8250
rect 117880 7610 117920 8250
rect 118000 7610 118040 8250
rect 118120 7610 118160 8250
rect 118240 7610 118280 8250
rect 118360 7610 118400 8250
rect 109260 5760 109300 6900
rect 109370 5760 109410 6900
rect 109480 5760 109520 6900
rect 109590 5760 109630 6900
rect 109700 5760 109740 6900
rect 109810 5760 109850 6900
rect 109920 5760 109960 6900
rect 110030 5760 110070 6900
rect 110140 5760 110180 6900
rect 110250 5760 110290 6900
rect 110360 5760 110400 6900
rect 110470 5760 110510 6900
rect 110580 5760 110620 6900
rect 116980 5760 117020 6900
rect 117090 5760 117130 6900
rect 117200 5760 117240 6900
rect 117310 5760 117350 6900
rect 117420 5760 117460 6900
rect 117530 5760 117570 6900
rect 117640 5760 117680 6900
rect 117750 5760 117790 6900
rect 117860 5760 117900 6900
rect 117970 5760 118010 6900
rect 118080 5760 118120 6900
rect 118190 5760 118230 6900
rect 118300 5760 118340 6900
rect 109260 4010 109300 4350
rect 109370 4010 109410 4350
rect 109480 4010 109520 4350
rect 109590 4010 109630 4350
rect 109700 4010 109740 4350
rect 109810 4010 109850 4350
rect 109920 4010 109960 4350
rect 110030 4010 110070 4350
rect 110140 4010 110180 4350
rect 110250 4010 110290 4350
rect 110360 4010 110400 4350
rect 110470 4010 110510 4350
rect 110580 4010 110620 4350
rect 116980 4010 117020 4350
rect 117090 4010 117130 4350
rect 117200 4010 117240 4350
rect 117310 4010 117350 4350
rect 117420 4010 117460 4350
rect 117530 4010 117570 4350
rect 117640 4010 117680 4350
rect 117750 4010 117790 4350
rect 117860 4010 117900 4350
rect 117970 4010 118010 4350
rect 118080 4010 118120 4350
rect 118190 4010 118230 4350
rect 118300 4010 118340 4350
<< psubdiff >>
rect 113460 6830 113540 6860
rect 113460 6390 113480 6830
rect 113520 6390 113540 6830
rect 113460 6360 113540 6390
rect 114060 6830 114140 6860
rect 114060 6390 114080 6830
rect 114120 6390 114140 6830
rect 114060 6360 114140 6390
rect 111980 5700 112060 5730
rect 111980 5460 112000 5700
rect 112040 5460 112060 5700
rect 111980 5430 112060 5460
rect 113460 5700 113540 5730
rect 113460 5460 113480 5700
rect 113520 5460 113540 5700
rect 113460 5430 113540 5460
rect 114060 5700 114140 5730
rect 114060 5460 114080 5700
rect 114120 5460 114140 5700
rect 114060 5430 114140 5460
rect 115540 5700 115620 5730
rect 115540 5460 115560 5700
rect 115600 5460 115620 5700
rect 115540 5430 115620 5460
rect 111980 3830 112060 3860
rect 111980 3590 112000 3830
rect 112040 3590 112060 3830
rect 111980 3560 112060 3590
rect 113460 3830 113540 3860
rect 113460 3590 113480 3830
rect 113520 3590 113540 3830
rect 113460 3560 113540 3590
rect 114060 3830 114140 3860
rect 114060 3590 114080 3830
rect 114120 3590 114140 3830
rect 114060 3560 114140 3590
rect 115540 3830 115620 3860
rect 115540 3590 115560 3830
rect 115600 3590 115620 3830
rect 115540 3560 115620 3590
rect 109160 3470 109240 3500
rect 109160 2930 109180 3470
rect 109220 2930 109240 3470
rect 109160 2900 109240 2930
rect 110640 3470 110720 3500
rect 110640 2930 110660 3470
rect 110700 2930 110720 3470
rect 116880 3470 116960 3500
rect 110640 2900 110720 2930
rect 116880 2930 116900 3470
rect 116940 2930 116960 3470
rect 116880 2900 116960 2930
rect 118360 3470 118440 3500
rect 118360 2930 118380 3470
rect 118420 2930 118440 3470
rect 118360 2900 118440 2930
rect 112360 1580 112440 1610
rect 109220 1350 109300 1380
rect 109220 10 109240 1350
rect 109280 10 109300 1350
rect 109220 -20 109300 10
rect 110580 1350 110660 1380
rect 110580 10 110600 1350
rect 110640 10 110660 1350
rect 112360 1140 112380 1580
rect 112420 1140 112440 1580
rect 112360 1110 112440 1140
rect 115050 1580 115130 1610
rect 115050 1140 115070 1580
rect 115110 1140 115130 1580
rect 115050 1110 115130 1140
rect 116940 1350 117020 1380
rect 110580 -20 110660 10
rect 113350 70 113430 100
rect 113350 -170 113370 70
rect 113410 -170 113430 70
rect 113350 -200 113430 -170
rect 114170 70 114250 100
rect 114170 -170 114190 70
rect 114230 -170 114250 70
rect 116940 10 116960 1350
rect 117000 10 117020 1350
rect 116940 -20 117020 10
rect 118300 1350 118380 1380
rect 118300 10 118320 1350
rect 118360 10 118380 1350
rect 118300 -20 118380 10
rect 114170 -200 114250 -170
<< nsubdiff >>
rect 109220 9770 109300 9800
rect 109220 9130 109240 9770
rect 109280 9130 109300 9770
rect 109220 9100 109300 9130
rect 110820 9770 110900 9800
rect 110820 9130 110840 9770
rect 110880 9130 110900 9770
rect 116700 9770 116780 9800
rect 110820 9100 110900 9130
rect 111890 9470 111970 9500
rect 111890 8830 111910 9470
rect 111950 8830 111970 9470
rect 111890 8800 111970 8830
rect 112410 9470 112490 9500
rect 112410 8830 112430 9470
rect 112470 8830 112490 9470
rect 114170 9470 114250 9500
rect 112410 8800 112490 8830
rect 112830 9130 112910 9160
rect 112830 8830 112850 9130
rect 112890 8830 112910 9130
rect 112830 8800 112910 8830
rect 113350 9130 113430 9160
rect 113350 8830 113370 9130
rect 113410 8830 113430 9130
rect 113350 8800 113430 8830
rect 114170 8830 114190 9470
rect 114230 8830 114250 9470
rect 114170 8800 114250 8830
rect 114690 9470 114770 9500
rect 114690 8830 114710 9470
rect 114750 8830 114770 9470
rect 114690 8800 114770 8830
rect 115110 9470 115190 9500
rect 115110 8830 115130 9470
rect 115170 8830 115190 9470
rect 115110 8800 115190 8830
rect 115630 9470 115710 9500
rect 115630 8830 115650 9470
rect 115690 8830 115710 9470
rect 116700 9130 116720 9770
rect 116760 9130 116780 9770
rect 116700 9100 116780 9130
rect 118300 9770 118380 9800
rect 118300 9130 118320 9770
rect 118360 9130 118380 9770
rect 118300 9100 118380 9130
rect 115630 8800 115710 8830
rect 109100 8250 109180 8280
rect 109100 7610 109120 8250
rect 109160 7610 109180 8250
rect 109100 7580 109180 7610
rect 110700 8250 110780 8280
rect 110700 7610 110720 8250
rect 110760 7610 110780 8250
rect 116820 8250 116900 8280
rect 110700 7580 110780 7610
rect 112940 8040 113020 8070
rect 112940 7600 112960 8040
rect 113000 7600 113020 8040
rect 112940 7570 113020 7600
rect 113760 8040 113840 8070
rect 113760 7600 113780 8040
rect 113820 7600 113840 8040
rect 113760 7570 113840 7600
rect 114580 8040 114660 8070
rect 114580 7600 114600 8040
rect 114640 7600 114660 8040
rect 114580 7570 114660 7600
rect 116820 7610 116840 8250
rect 116880 7610 116900 8250
rect 116820 7580 116900 7610
rect 118420 8250 118500 8280
rect 118420 7610 118440 8250
rect 118480 7610 118500 8250
rect 118420 7580 118500 7610
rect 109160 6900 109240 6930
rect 109160 5760 109180 6900
rect 109220 5760 109240 6900
rect 109160 5730 109240 5760
rect 110640 6900 110720 6930
rect 110640 5760 110660 6900
rect 110700 5760 110720 6900
rect 116880 6900 116960 6930
rect 116880 5760 116900 6900
rect 116940 5760 116960 6900
rect 110640 5730 110720 5760
rect 116880 5730 116960 5760
rect 118360 6900 118440 6930
rect 118360 5760 118380 6900
rect 118420 5760 118440 6900
rect 118360 5730 118440 5760
rect 109160 4350 109240 4380
rect 109160 4010 109180 4350
rect 109220 4010 109240 4350
rect 109160 3980 109240 4010
rect 110640 4350 110720 4380
rect 110640 4010 110660 4350
rect 110700 4010 110720 4350
rect 116880 4350 116960 4380
rect 110640 3980 110720 4010
rect 116880 4010 116900 4350
rect 116940 4010 116960 4350
rect 116880 3980 116960 4010
rect 118360 4350 118440 4380
rect 118360 4010 118380 4350
rect 118420 4010 118440 4350
rect 118360 3980 118440 4010
<< psubdiffcont >>
rect 113480 6390 113520 6830
rect 114080 6390 114120 6830
rect 112000 5460 112040 5700
rect 113480 5460 113520 5700
rect 114080 5460 114120 5700
rect 115560 5460 115600 5700
rect 112000 3590 112040 3830
rect 113480 3590 113520 3830
rect 114080 3590 114120 3830
rect 115560 3590 115600 3830
rect 109180 2930 109220 3470
rect 110660 2930 110700 3470
rect 116900 2930 116940 3470
rect 118380 2930 118420 3470
rect 109240 10 109280 1350
rect 110600 10 110640 1350
rect 112380 1140 112420 1580
rect 115070 1140 115110 1580
rect 113370 -170 113410 70
rect 114190 -170 114230 70
rect 116960 10 117000 1350
rect 118320 10 118360 1350
<< nsubdiffcont >>
rect 109240 9130 109280 9770
rect 110840 9130 110880 9770
rect 111910 8830 111950 9470
rect 112430 8830 112470 9470
rect 112850 8830 112890 9130
rect 113370 8830 113410 9130
rect 114190 8830 114230 9470
rect 114710 8830 114750 9470
rect 115130 8830 115170 9470
rect 115650 8830 115690 9470
rect 116720 9130 116760 9770
rect 118320 9130 118360 9770
rect 109120 7610 109160 8250
rect 110720 7610 110760 8250
rect 112960 7600 113000 8040
rect 113780 7600 113820 8040
rect 114600 7600 114640 8040
rect 116840 7610 116880 8250
rect 118440 7610 118480 8250
rect 109180 5760 109220 6900
rect 110660 5760 110700 6900
rect 116900 5760 116940 6900
rect 118380 5760 118420 6900
rect 109180 4010 109220 4350
rect 110660 4010 110700 4350
rect 116900 4010 116940 4350
rect 118380 4010 118420 4350
<< poly >>
rect 109490 9970 109550 9990
rect 109490 9930 109500 9970
rect 109540 9930 109550 9970
rect 109490 9910 109550 9930
rect 109610 9970 109670 9990
rect 109610 9930 109620 9970
rect 109660 9930 109670 9970
rect 109610 9910 109670 9930
rect 109730 9970 109790 9990
rect 109730 9930 109740 9970
rect 109780 9930 109790 9970
rect 109730 9910 109790 9930
rect 109850 9970 109910 9990
rect 109850 9930 109860 9970
rect 109900 9930 109910 9970
rect 109850 9910 109910 9930
rect 109970 9970 110030 9990
rect 109970 9930 109980 9970
rect 110020 9930 110030 9970
rect 109970 9910 110030 9930
rect 110090 9970 110150 9990
rect 110090 9930 110100 9970
rect 110140 9930 110150 9970
rect 110090 9910 110150 9930
rect 110210 9970 110270 9990
rect 110210 9930 110220 9970
rect 110260 9930 110270 9970
rect 110210 9910 110270 9930
rect 110330 9970 110390 9990
rect 110330 9930 110340 9970
rect 110380 9930 110390 9970
rect 110330 9910 110390 9930
rect 110450 9970 110510 9990
rect 110450 9930 110460 9970
rect 110500 9930 110510 9970
rect 110450 9910 110510 9930
rect 110570 9970 110630 9990
rect 110570 9930 110580 9970
rect 110620 9930 110630 9970
rect 110570 9910 110630 9930
rect 116970 9970 117030 9990
rect 116970 9930 116980 9970
rect 117020 9930 117030 9970
rect 116970 9910 117030 9930
rect 117090 9970 117150 9990
rect 117090 9930 117100 9970
rect 117140 9930 117150 9970
rect 117090 9910 117150 9930
rect 117210 9970 117270 9990
rect 117210 9930 117220 9970
rect 117260 9930 117270 9970
rect 117210 9910 117270 9930
rect 117330 9970 117390 9990
rect 117330 9930 117340 9970
rect 117380 9930 117390 9970
rect 117330 9910 117390 9930
rect 117450 9970 117510 9990
rect 117450 9930 117460 9970
rect 117500 9930 117510 9970
rect 117450 9910 117510 9930
rect 117570 9970 117630 9990
rect 117570 9930 117580 9970
rect 117620 9930 117630 9970
rect 117570 9910 117630 9930
rect 117690 9970 117750 9990
rect 117690 9930 117700 9970
rect 117740 9930 117750 9970
rect 117690 9910 117750 9930
rect 117810 9970 117870 9990
rect 117810 9930 117820 9970
rect 117860 9930 117870 9970
rect 117810 9910 117870 9930
rect 117930 9970 117990 9990
rect 117930 9930 117940 9970
rect 117980 9930 117990 9970
rect 117930 9910 117990 9930
rect 118050 9970 118110 9990
rect 118050 9930 118060 9970
rect 118100 9930 118110 9970
rect 118050 9910 118110 9930
rect 109380 9800 109420 9830
rect 109500 9800 109540 9910
rect 109620 9800 109660 9910
rect 109740 9800 109780 9910
rect 109860 9800 109900 9910
rect 109980 9800 110020 9910
rect 110100 9800 110140 9910
rect 110220 9800 110260 9910
rect 110340 9800 110380 9910
rect 110460 9800 110500 9910
rect 110580 9800 110620 9910
rect 110700 9800 110740 9830
rect 116860 9800 116900 9830
rect 116980 9800 117020 9910
rect 117100 9800 117140 9910
rect 117220 9800 117260 9910
rect 117340 9800 117380 9910
rect 117460 9800 117500 9910
rect 117580 9800 117620 9910
rect 117700 9800 117740 9910
rect 117820 9800 117860 9910
rect 117940 9800 117980 9910
rect 118060 9800 118100 9910
rect 118180 9800 118220 9830
rect 111970 9590 112050 9610
rect 111970 9550 111990 9590
rect 112030 9560 112050 9590
rect 112330 9590 112410 9610
rect 112330 9560 112350 9590
rect 112030 9550 112090 9560
rect 111970 9530 112090 9550
rect 112290 9550 112350 9560
rect 112390 9550 112410 9590
rect 112290 9530 112410 9550
rect 114250 9590 114330 9610
rect 114250 9550 114270 9590
rect 114310 9560 114330 9590
rect 114610 9590 114690 9610
rect 114610 9560 114630 9590
rect 114310 9550 114370 9560
rect 114250 9530 114370 9550
rect 114570 9550 114630 9560
rect 114670 9550 114690 9590
rect 114570 9530 114690 9550
rect 115190 9590 115270 9610
rect 115190 9550 115210 9590
rect 115250 9560 115270 9590
rect 115550 9590 115630 9610
rect 115550 9560 115570 9590
rect 115250 9550 115310 9560
rect 115190 9530 115310 9550
rect 115510 9550 115570 9560
rect 115610 9550 115630 9590
rect 115510 9530 115630 9550
rect 112050 9500 112090 9530
rect 112170 9500 112210 9530
rect 112290 9500 112330 9530
rect 114330 9500 114370 9530
rect 114450 9500 114490 9530
rect 114570 9500 114610 9530
rect 115270 9500 115310 9530
rect 115390 9500 115430 9530
rect 115510 9500 115550 9530
rect 109380 9070 109420 9100
rect 109500 9070 109540 9100
rect 109620 9070 109660 9100
rect 109740 9070 109780 9100
rect 109860 9070 109900 9100
rect 109980 9070 110020 9100
rect 110100 9070 110140 9100
rect 110220 9070 110260 9100
rect 110340 9070 110380 9100
rect 110460 9070 110500 9100
rect 110580 9070 110620 9100
rect 110700 9070 110740 9100
rect 109300 9050 109420 9070
rect 109300 9010 109320 9050
rect 109360 9040 109420 9050
rect 110700 9050 110820 9070
rect 110700 9040 110760 9050
rect 109360 9010 109380 9040
rect 109300 8990 109380 9010
rect 110740 9010 110760 9040
rect 110800 9010 110820 9050
rect 110740 8990 110820 9010
rect 112910 9250 112990 9270
rect 112910 9210 112930 9250
rect 112970 9220 112990 9250
rect 113270 9250 113350 9270
rect 113270 9220 113290 9250
rect 112970 9210 113030 9220
rect 112910 9190 113030 9210
rect 113230 9210 113290 9220
rect 113330 9210 113350 9250
rect 113230 9190 113350 9210
rect 112990 9160 113030 9190
rect 113110 9160 113150 9190
rect 113230 9160 113270 9190
rect 116860 9070 116900 9100
rect 116980 9070 117020 9100
rect 117100 9070 117140 9100
rect 117220 9070 117260 9100
rect 117340 9070 117380 9100
rect 117460 9070 117500 9100
rect 117580 9070 117620 9100
rect 117700 9070 117740 9100
rect 117820 9070 117860 9100
rect 117940 9070 117980 9100
rect 118060 9070 118100 9100
rect 118180 9070 118220 9100
rect 116780 9050 116900 9070
rect 116780 9010 116800 9050
rect 116840 9040 116900 9050
rect 118180 9050 118300 9070
rect 118180 9040 118240 9050
rect 116840 9010 116860 9040
rect 116780 8990 116860 9010
rect 118220 9010 118240 9040
rect 118280 9010 118300 9050
rect 118220 8990 118300 9010
rect 112050 8770 112090 8800
rect 112170 8690 112210 8800
rect 112290 8770 112330 8800
rect 112990 8770 113030 8800
rect 113110 8690 113150 8800
rect 113230 8770 113270 8800
rect 114330 8770 114370 8800
rect 112100 8670 112210 8690
rect 112100 8630 112120 8670
rect 112160 8630 112210 8670
rect 112100 8610 112210 8630
rect 113060 8670 113150 8690
rect 113060 8630 113070 8670
rect 113110 8660 113150 8670
rect 114450 8690 114490 8800
rect 114570 8770 114610 8800
rect 115270 8770 115310 8800
rect 115390 8690 115430 8800
rect 115510 8770 115550 8800
rect 114450 8670 114540 8690
rect 114450 8660 114490 8670
rect 113110 8630 113120 8660
rect 113060 8610 113120 8630
rect 114480 8630 114490 8660
rect 114530 8630 114540 8670
rect 114480 8610 114540 8630
rect 115352 8670 115430 8690
rect 115352 8630 115362 8670
rect 115402 8660 115430 8670
rect 115402 8630 115412 8660
rect 115352 8610 115412 8630
rect 109190 8370 109250 8390
rect 109190 8330 109200 8370
rect 109240 8340 109250 8370
rect 110630 8370 110690 8390
rect 110630 8340 110640 8370
rect 109240 8330 109300 8340
rect 109190 8310 109300 8330
rect 110580 8330 110640 8340
rect 110680 8330 110690 8370
rect 110580 8310 110690 8330
rect 116910 8370 116970 8390
rect 116910 8330 116920 8370
rect 116960 8340 116970 8370
rect 118350 8370 118410 8390
rect 118350 8340 118360 8370
rect 116960 8330 117020 8340
rect 116910 8310 117020 8330
rect 118300 8330 118360 8340
rect 118400 8330 118410 8370
rect 118300 8310 118410 8330
rect 109260 8280 109300 8310
rect 109380 8280 109420 8310
rect 109500 8280 109540 8310
rect 109620 8280 109660 8310
rect 109740 8280 109780 8310
rect 109860 8280 109900 8310
rect 109980 8280 110020 8310
rect 110100 8280 110140 8310
rect 110220 8280 110260 8310
rect 110340 8280 110380 8310
rect 110460 8280 110500 8310
rect 110580 8280 110620 8310
rect 113020 8290 113100 8310
rect 113020 8250 113040 8290
rect 113080 8260 113100 8290
rect 113680 8290 113760 8310
rect 113680 8260 113700 8290
rect 113080 8250 113130 8260
rect 113020 8230 113130 8250
rect 113100 8070 113130 8230
rect 113650 8250 113700 8260
rect 113740 8250 113760 8290
rect 113650 8230 113760 8250
rect 113840 8290 113920 8310
rect 113840 8250 113860 8290
rect 113900 8260 113920 8290
rect 114500 8290 114580 8310
rect 114500 8260 114520 8290
rect 113900 8250 113950 8260
rect 113840 8230 113950 8250
rect 113210 8070 113240 8100
rect 113320 8070 113350 8100
rect 113430 8070 113460 8100
rect 113540 8070 113570 8100
rect 113650 8070 113680 8230
rect 113920 8070 113950 8230
rect 114470 8250 114520 8260
rect 114560 8250 114580 8290
rect 116980 8280 117020 8310
rect 117100 8280 117140 8310
rect 117220 8280 117260 8310
rect 117340 8280 117380 8310
rect 117460 8280 117500 8310
rect 117580 8280 117620 8310
rect 117700 8280 117740 8310
rect 117820 8280 117860 8310
rect 117940 8280 117980 8310
rect 118060 8280 118100 8310
rect 118180 8280 118220 8310
rect 118300 8280 118340 8310
rect 114470 8230 114580 8250
rect 114030 8070 114060 8100
rect 114140 8070 114170 8100
rect 114250 8070 114280 8100
rect 114360 8070 114390 8100
rect 114470 8070 114500 8230
rect 109260 7550 109300 7580
rect 109380 7470 109420 7580
rect 109500 7470 109540 7580
rect 109620 7470 109660 7580
rect 109740 7470 109780 7580
rect 109860 7470 109900 7580
rect 109980 7470 110020 7580
rect 110100 7470 110140 7580
rect 110220 7470 110260 7580
rect 110340 7470 110380 7580
rect 110460 7470 110500 7580
rect 110580 7550 110620 7580
rect 113100 7540 113130 7570
rect 113210 7540 113240 7570
rect 113320 7550 113350 7570
rect 113430 7550 113460 7570
rect 113210 7520 113274 7540
rect 113320 7520 113460 7550
rect 113540 7540 113570 7570
rect 113650 7540 113680 7570
rect 113920 7540 113950 7570
rect 114030 7540 114060 7570
rect 114140 7550 114170 7570
rect 114250 7550 114280 7570
rect 113506 7520 113570 7540
rect 114030 7520 114094 7540
rect 114140 7520 114280 7550
rect 114360 7540 114390 7570
rect 114470 7540 114500 7570
rect 116980 7550 117020 7580
rect 114326 7520 114390 7540
rect 113214 7480 113224 7520
rect 113264 7480 113274 7520
rect 109370 7450 109430 7470
rect 109370 7410 109380 7450
rect 109420 7410 109430 7450
rect 109370 7390 109430 7410
rect 109490 7450 109550 7470
rect 109490 7410 109500 7450
rect 109540 7410 109550 7450
rect 109490 7390 109550 7410
rect 109610 7450 109670 7470
rect 109610 7410 109620 7450
rect 109660 7410 109670 7450
rect 109610 7390 109670 7410
rect 109730 7450 109790 7470
rect 109730 7410 109740 7450
rect 109780 7410 109790 7450
rect 109730 7390 109790 7410
rect 109850 7450 109910 7470
rect 109850 7410 109860 7450
rect 109900 7410 109910 7450
rect 109850 7390 109910 7410
rect 109970 7450 110030 7470
rect 109970 7410 109980 7450
rect 110020 7410 110030 7450
rect 109970 7390 110030 7410
rect 110090 7450 110150 7470
rect 110090 7410 110100 7450
rect 110140 7410 110150 7450
rect 110090 7390 110150 7410
rect 110210 7450 110270 7470
rect 110210 7410 110220 7450
rect 110260 7410 110270 7450
rect 110210 7390 110270 7410
rect 110330 7450 110390 7470
rect 110330 7410 110340 7450
rect 110380 7410 110390 7450
rect 110330 7390 110390 7410
rect 110450 7450 110510 7470
rect 113214 7460 113274 7480
rect 113350 7480 113370 7520
rect 113410 7480 113430 7520
rect 113350 7460 113430 7480
rect 113506 7480 113516 7520
rect 113556 7480 113566 7520
rect 113506 7460 113566 7480
rect 114034 7480 114044 7520
rect 114084 7480 114094 7520
rect 114034 7460 114094 7480
rect 114170 7480 114190 7520
rect 114230 7480 114250 7520
rect 114170 7460 114250 7480
rect 114326 7480 114336 7520
rect 114376 7480 114386 7520
rect 114326 7460 114386 7480
rect 117100 7470 117140 7580
rect 117220 7470 117260 7580
rect 117340 7470 117380 7580
rect 117460 7470 117500 7580
rect 117580 7470 117620 7580
rect 117700 7470 117740 7580
rect 117820 7470 117860 7580
rect 117940 7470 117980 7580
rect 118060 7470 118100 7580
rect 118180 7470 118220 7580
rect 118300 7550 118340 7580
rect 110450 7410 110460 7450
rect 110500 7410 110510 7450
rect 110450 7390 110510 7410
rect 117090 7450 117150 7470
rect 117090 7410 117100 7450
rect 117140 7410 117150 7450
rect 117090 7390 117150 7410
rect 117210 7450 117270 7470
rect 117210 7410 117220 7450
rect 117260 7410 117270 7450
rect 117210 7390 117270 7410
rect 117330 7450 117390 7470
rect 117330 7410 117340 7450
rect 117380 7410 117390 7450
rect 117330 7390 117390 7410
rect 117450 7450 117510 7470
rect 117450 7410 117460 7450
rect 117500 7410 117510 7450
rect 117450 7390 117510 7410
rect 117570 7450 117630 7470
rect 117570 7410 117580 7450
rect 117620 7410 117630 7450
rect 117570 7390 117630 7410
rect 117690 7450 117750 7470
rect 117690 7410 117700 7450
rect 117740 7410 117750 7450
rect 117690 7390 117750 7410
rect 117810 7450 117870 7470
rect 117810 7410 117820 7450
rect 117860 7410 117870 7450
rect 117810 7390 117870 7410
rect 117930 7450 117990 7470
rect 117930 7410 117940 7450
rect 117980 7410 117990 7450
rect 117930 7390 117990 7410
rect 118050 7450 118110 7470
rect 118050 7410 118060 7450
rect 118100 7410 118110 7450
rect 118050 7390 118110 7410
rect 118170 7450 118230 7470
rect 118170 7410 118180 7450
rect 118220 7410 118230 7450
rect 118170 7390 118230 7410
rect 109250 7020 109310 7040
rect 109250 6980 109260 7020
rect 109300 6990 109310 7020
rect 110570 7020 110630 7040
rect 110570 6990 110580 7020
rect 109300 6980 109350 6990
rect 109250 6960 109350 6980
rect 110530 6980 110580 6990
rect 110620 6980 110630 7020
rect 110530 6960 110630 6980
rect 116970 7020 117030 7040
rect 116970 6980 116980 7020
rect 117020 6990 117030 7020
rect 118290 7020 118350 7040
rect 118290 6990 118300 7020
rect 117020 6980 117070 6990
rect 109320 6930 109350 6960
rect 109430 6930 109460 6960
rect 109540 6930 109570 6960
rect 109650 6930 109680 6960
rect 109760 6930 109790 6960
rect 109870 6930 109900 6960
rect 109980 6930 110010 6960
rect 110090 6930 110120 6960
rect 110200 6930 110230 6960
rect 110310 6930 110340 6960
rect 110420 6930 110450 6960
rect 110530 6930 110560 6960
rect 113700 6950 113780 6970
rect 116970 6960 117070 6980
rect 118250 6980 118300 6990
rect 118340 6980 118350 7020
rect 118250 6960 118350 6980
rect 113700 6910 113720 6950
rect 113760 6910 113780 6950
rect 117040 6930 117070 6960
rect 117150 6930 117180 6960
rect 117260 6930 117290 6960
rect 117370 6930 117400 6960
rect 117480 6930 117510 6960
rect 117590 6930 117620 6960
rect 117700 6930 117730 6960
rect 117810 6930 117840 6960
rect 117920 6930 117950 6960
rect 118030 6930 118060 6960
rect 118140 6930 118170 6960
rect 118250 6930 118280 6960
rect 113700 6890 113870 6910
rect 113620 6860 113650 6890
rect 113730 6880 113870 6890
rect 113730 6860 113760 6880
rect 113840 6860 113870 6880
rect 113950 6860 113980 6890
rect 113620 6330 113650 6360
rect 113730 6330 113760 6360
rect 113840 6330 113870 6360
rect 113950 6330 113980 6360
rect 113540 6310 113650 6330
rect 113540 6270 113560 6310
rect 113600 6300 113650 6310
rect 113950 6310 114060 6330
rect 113950 6300 114000 6310
rect 113600 6270 113620 6300
rect 113540 6250 113620 6270
rect 113980 6270 114000 6300
rect 114040 6270 114060 6310
rect 113980 6250 114060 6270
rect 112232 5820 112298 5840
rect 112232 5780 112245 5820
rect 112285 5780 112298 5820
rect 112232 5760 112298 5780
rect 112342 5820 112408 5840
rect 112342 5780 112355 5820
rect 112395 5780 112408 5820
rect 112342 5760 112408 5780
rect 112452 5820 112518 5840
rect 112452 5780 112465 5820
rect 112505 5780 112518 5820
rect 112452 5760 112518 5780
rect 112562 5820 112628 5840
rect 112562 5780 112575 5820
rect 112615 5780 112628 5820
rect 112562 5760 112628 5780
rect 112672 5820 112738 5840
rect 112672 5780 112685 5820
rect 112725 5780 112738 5820
rect 112672 5760 112738 5780
rect 112782 5820 112848 5840
rect 112782 5780 112795 5820
rect 112835 5780 112848 5820
rect 112782 5760 112848 5780
rect 112892 5820 112958 5840
rect 112892 5780 112905 5820
rect 112945 5780 112958 5820
rect 112892 5760 112958 5780
rect 113002 5820 113068 5840
rect 113002 5780 113015 5820
rect 113055 5780 113068 5820
rect 113002 5760 113068 5780
rect 113112 5820 113178 5840
rect 113112 5780 113125 5820
rect 113165 5780 113178 5820
rect 113112 5760 113178 5780
rect 113222 5820 113288 5840
rect 113222 5780 113235 5820
rect 113275 5780 113288 5820
rect 113222 5760 113288 5780
rect 114312 5820 114378 5840
rect 114312 5780 114325 5820
rect 114365 5780 114378 5820
rect 114312 5760 114378 5780
rect 114422 5820 114488 5840
rect 114422 5780 114435 5820
rect 114475 5780 114488 5820
rect 114422 5760 114488 5780
rect 114532 5820 114598 5840
rect 114532 5780 114545 5820
rect 114585 5780 114598 5820
rect 114532 5760 114598 5780
rect 114642 5820 114708 5840
rect 114642 5780 114655 5820
rect 114695 5780 114708 5820
rect 114642 5760 114708 5780
rect 114752 5820 114818 5840
rect 114752 5780 114765 5820
rect 114805 5780 114818 5820
rect 114752 5760 114818 5780
rect 114862 5820 114928 5840
rect 114862 5780 114875 5820
rect 114915 5780 114928 5820
rect 114862 5760 114928 5780
rect 114972 5820 115038 5840
rect 114972 5780 114985 5820
rect 115025 5780 115038 5820
rect 114972 5760 115038 5780
rect 115082 5820 115148 5840
rect 115082 5780 115095 5820
rect 115135 5780 115148 5820
rect 115082 5760 115148 5780
rect 115192 5820 115258 5840
rect 115192 5780 115205 5820
rect 115245 5780 115258 5820
rect 115192 5760 115258 5780
rect 115302 5820 115368 5840
rect 115302 5780 115315 5820
rect 115355 5780 115368 5820
rect 115302 5760 115368 5780
rect 112140 5730 112170 5760
rect 112250 5730 112280 5760
rect 112360 5730 112390 5760
rect 112470 5730 112500 5760
rect 112580 5730 112610 5760
rect 112690 5730 112720 5760
rect 112800 5730 112830 5760
rect 112910 5730 112940 5760
rect 113020 5730 113050 5760
rect 113130 5730 113160 5760
rect 113240 5730 113270 5760
rect 113350 5730 113380 5760
rect 114220 5730 114250 5760
rect 114330 5730 114360 5760
rect 114440 5730 114470 5760
rect 114550 5730 114580 5760
rect 114660 5730 114690 5760
rect 114770 5730 114800 5760
rect 114880 5730 114910 5760
rect 114990 5730 115020 5760
rect 115100 5730 115130 5760
rect 115210 5730 115240 5760
rect 115320 5730 115350 5760
rect 115430 5730 115460 5760
rect 109320 5700 109350 5730
rect 109430 5710 109460 5730
rect 109540 5710 109570 5730
rect 109650 5710 109680 5730
rect 109760 5710 109790 5730
rect 109870 5710 109900 5730
rect 109980 5710 110010 5730
rect 110090 5710 110120 5730
rect 110200 5710 110230 5730
rect 110310 5710 110340 5730
rect 110420 5710 110450 5730
rect 109430 5680 110450 5710
rect 110530 5700 110560 5730
rect 109910 5640 109920 5680
rect 109960 5640 109970 5680
rect 109910 5570 109970 5640
rect 109900 5550 109980 5570
rect 109900 5510 109920 5550
rect 109960 5510 109980 5550
rect 109900 5470 109980 5510
rect 109900 5430 109920 5470
rect 109960 5430 109980 5470
rect 117040 5700 117070 5730
rect 117150 5710 117180 5730
rect 117260 5710 117290 5730
rect 117370 5710 117400 5730
rect 117480 5710 117510 5730
rect 117590 5710 117620 5730
rect 117700 5710 117730 5730
rect 117810 5710 117840 5730
rect 117920 5710 117950 5730
rect 118030 5710 118060 5730
rect 118140 5710 118170 5730
rect 117150 5680 118170 5710
rect 118250 5700 118280 5730
rect 117630 5640 117640 5680
rect 117680 5640 117690 5680
rect 117630 5570 117690 5640
rect 117620 5550 117700 5570
rect 117620 5510 117640 5550
rect 117680 5510 117700 5550
rect 117620 5470 117700 5510
rect 117620 5430 117640 5470
rect 117680 5430 117700 5470
rect 109900 5390 109980 5430
rect 112140 5400 112170 5430
rect 112250 5400 112280 5430
rect 112360 5400 112390 5430
rect 112470 5400 112500 5430
rect 112580 5400 112610 5430
rect 112690 5400 112720 5430
rect 112800 5400 112830 5430
rect 112910 5400 112940 5430
rect 113020 5400 113050 5430
rect 113130 5400 113160 5430
rect 113240 5400 113270 5430
rect 113350 5400 113380 5430
rect 114220 5400 114250 5430
rect 114330 5400 114360 5430
rect 114440 5400 114470 5430
rect 114550 5400 114580 5430
rect 114660 5400 114690 5430
rect 114770 5400 114800 5430
rect 114880 5400 114910 5430
rect 114990 5400 115020 5430
rect 115100 5400 115130 5430
rect 115210 5400 115240 5430
rect 115320 5400 115350 5430
rect 115430 5400 115460 5430
rect 109900 5350 109920 5390
rect 109960 5350 109980 5390
rect 109900 5330 109980 5350
rect 112070 5380 112170 5400
rect 112070 5340 112080 5380
rect 112120 5370 112170 5380
rect 113350 5380 113450 5400
rect 113350 5370 113400 5380
rect 112120 5340 112130 5370
rect 112070 5320 112130 5340
rect 113390 5340 113400 5370
rect 113440 5340 113450 5380
rect 113390 5320 113450 5340
rect 114150 5380 114250 5400
rect 114150 5340 114160 5380
rect 114200 5370 114250 5380
rect 115430 5380 115530 5400
rect 115430 5370 115480 5380
rect 114200 5340 114210 5370
rect 114150 5320 114210 5340
rect 115470 5340 115480 5370
rect 115520 5340 115530 5380
rect 115470 5320 115530 5340
rect 117620 5390 117700 5430
rect 117620 5350 117640 5390
rect 117680 5350 117700 5390
rect 117620 5330 117700 5350
rect 109250 4470 109310 4490
rect 109250 4430 109260 4470
rect 109300 4440 109310 4470
rect 110570 4470 110630 4490
rect 110570 4440 110580 4470
rect 109300 4430 109350 4440
rect 109250 4410 109350 4430
rect 110530 4430 110580 4440
rect 110620 4430 110630 4470
rect 110530 4410 110630 4430
rect 116970 4470 117030 4490
rect 116970 4430 116980 4470
rect 117020 4440 117030 4470
rect 118290 4470 118350 4490
rect 118290 4440 118300 4470
rect 117020 4430 117070 4440
rect 116970 4410 117070 4430
rect 118250 4430 118300 4440
rect 118340 4430 118350 4470
rect 118250 4410 118350 4430
rect 109320 4380 109350 4410
rect 109430 4380 109460 4410
rect 109540 4380 109570 4410
rect 109650 4380 109680 4410
rect 109760 4380 109790 4410
rect 109870 4380 109900 4410
rect 109980 4380 110010 4410
rect 110090 4380 110120 4410
rect 110200 4380 110230 4410
rect 110310 4380 110340 4410
rect 110420 4380 110450 4410
rect 110530 4380 110560 4410
rect 117040 4380 117070 4410
rect 117150 4380 117180 4410
rect 117260 4380 117290 4410
rect 117370 4380 117400 4410
rect 117480 4380 117510 4410
rect 117590 4380 117620 4410
rect 117700 4380 117730 4410
rect 117810 4380 117840 4410
rect 117920 4380 117950 4410
rect 118030 4380 118060 4410
rect 118140 4380 118170 4410
rect 118250 4380 118280 4410
rect 113380 4020 113440 4040
rect 112080 4000 112140 4020
rect 109320 3950 109350 3980
rect 109430 3960 109460 3980
rect 109540 3960 109570 3980
rect 109650 3960 109680 3980
rect 109760 3960 109790 3980
rect 109870 3960 109900 3980
rect 109980 3960 110010 3980
rect 110090 3960 110120 3980
rect 110200 3960 110230 3980
rect 110310 3960 110340 3980
rect 110420 3960 110450 3980
rect 109430 3930 110450 3960
rect 110530 3950 110560 3980
rect 112080 3960 112090 4000
rect 112130 3970 112140 4000
rect 113380 3990 113390 4020
rect 113240 3980 113390 3990
rect 113430 3980 113440 4020
rect 112130 3960 112280 3970
rect 112080 3940 112280 3960
rect 110240 3890 110250 3930
rect 110290 3890 110300 3930
rect 112250 3910 112280 3940
rect 113240 3960 113440 3980
rect 113680 4020 113740 4040
rect 113680 3980 113690 4020
rect 113730 3990 113740 4020
rect 113860 4020 113920 4040
rect 113860 3990 113870 4020
rect 113730 3980 113760 3990
rect 113680 3960 113760 3980
rect 113240 3910 113270 3960
rect 110240 3870 110300 3890
rect 110250 3820 110290 3870
rect 112140 3860 112170 3890
rect 112250 3880 113270 3910
rect 112250 3860 112280 3880
rect 112360 3860 112390 3880
rect 112470 3860 112500 3880
rect 112580 3860 112610 3880
rect 112690 3860 112720 3880
rect 112800 3860 112830 3880
rect 112910 3860 112940 3880
rect 113020 3860 113050 3880
rect 113130 3860 113160 3880
rect 113240 3860 113270 3880
rect 113350 3860 113380 3890
rect 113620 3860 113650 3890
rect 113730 3860 113760 3960
rect 113840 3980 113870 3990
rect 113910 3980 113920 4020
rect 113840 3960 113920 3980
rect 114160 4020 114220 4040
rect 114160 3980 114170 4020
rect 114210 3990 114220 4020
rect 115460 4000 115520 4020
rect 114210 3980 114360 3990
rect 114160 3960 114360 3980
rect 115460 3970 115470 4000
rect 113840 3860 113870 3960
rect 114330 3910 114360 3960
rect 115320 3960 115470 3970
rect 115510 3960 115520 4000
rect 115320 3940 115520 3960
rect 117040 3950 117070 3980
rect 117150 3960 117180 3980
rect 117260 3960 117290 3980
rect 117370 3960 117400 3980
rect 117480 3960 117510 3980
rect 117590 3960 117620 3980
rect 117700 3960 117730 3980
rect 117810 3960 117840 3980
rect 117920 3960 117950 3980
rect 118030 3960 118060 3980
rect 118140 3960 118170 3980
rect 115320 3910 115350 3940
rect 117150 3930 118170 3960
rect 118250 3950 118280 3980
rect 113950 3860 113980 3890
rect 114220 3860 114250 3890
rect 114330 3880 115350 3910
rect 117300 3890 117310 3930
rect 117350 3890 117360 3930
rect 114330 3860 114360 3880
rect 114440 3860 114470 3880
rect 114550 3860 114580 3880
rect 114660 3860 114690 3880
rect 114770 3860 114800 3880
rect 114880 3860 114910 3880
rect 114990 3860 115020 3880
rect 115100 3860 115130 3880
rect 115210 3860 115240 3880
rect 115320 3860 115350 3880
rect 115430 3860 115460 3890
rect 117300 3870 117360 3890
rect 110230 3800 110310 3820
rect 110230 3760 110250 3800
rect 110290 3760 110310 3800
rect 110230 3720 110310 3760
rect 110230 3680 110250 3720
rect 110290 3680 110310 3720
rect 110230 3660 110310 3680
rect 110250 3610 110290 3660
rect 110240 3590 110300 3610
rect 110240 3550 110250 3590
rect 110290 3550 110300 3590
rect 117310 3820 117350 3870
rect 117290 3800 117370 3820
rect 117290 3760 117310 3800
rect 117350 3760 117370 3800
rect 117290 3720 117370 3760
rect 117290 3680 117310 3720
rect 117350 3680 117370 3720
rect 117290 3660 117370 3680
rect 117310 3610 117350 3660
rect 117300 3590 117360 3610
rect 109320 3500 109350 3530
rect 109430 3520 110450 3550
rect 112140 3530 112170 3560
rect 112250 3530 112280 3560
rect 112360 3530 112390 3560
rect 112470 3530 112500 3560
rect 112580 3530 112610 3560
rect 112690 3530 112720 3560
rect 112800 3530 112830 3560
rect 112910 3530 112940 3560
rect 113020 3530 113050 3560
rect 113130 3530 113160 3560
rect 113240 3530 113270 3560
rect 113350 3530 113380 3560
rect 113620 3530 113650 3560
rect 113730 3530 113760 3560
rect 113840 3530 113870 3560
rect 113950 3530 113980 3560
rect 114220 3530 114250 3560
rect 114330 3530 114360 3560
rect 114440 3530 114470 3560
rect 114550 3530 114580 3560
rect 114660 3530 114690 3560
rect 114770 3530 114800 3560
rect 114880 3530 114910 3560
rect 114990 3530 115020 3560
rect 115100 3530 115130 3560
rect 115210 3530 115240 3560
rect 115320 3530 115350 3560
rect 115430 3530 115460 3560
rect 117300 3550 117310 3590
rect 117350 3550 117360 3590
rect 109430 3500 109460 3520
rect 109540 3500 109570 3520
rect 109650 3500 109680 3520
rect 109760 3500 109790 3520
rect 109870 3500 109900 3520
rect 109980 3500 110010 3520
rect 110090 3500 110120 3520
rect 110200 3500 110230 3520
rect 110310 3500 110340 3520
rect 110420 3500 110450 3520
rect 110530 3500 110560 3530
rect 112070 3510 112170 3530
rect 112070 3470 112080 3510
rect 112120 3500 112170 3510
rect 113350 3510 113650 3530
rect 113350 3500 113480 3510
rect 112120 3470 112130 3500
rect 112070 3450 112130 3470
rect 113470 3470 113480 3500
rect 113520 3500 113650 3510
rect 113950 3510 114250 3530
rect 113950 3500 114080 3510
rect 113520 3470 113530 3500
rect 113470 3450 113530 3470
rect 114070 3470 114080 3500
rect 114120 3500 114250 3510
rect 115430 3510 115530 3530
rect 115430 3500 115480 3510
rect 114120 3470 114130 3500
rect 114070 3450 114130 3470
rect 115470 3470 115480 3500
rect 115520 3470 115530 3510
rect 117040 3500 117070 3530
rect 117150 3520 118170 3550
rect 117150 3500 117180 3520
rect 117260 3500 117290 3520
rect 117370 3500 117400 3520
rect 117480 3500 117510 3520
rect 117590 3500 117620 3520
rect 117700 3500 117730 3520
rect 117810 3500 117840 3520
rect 117920 3500 117950 3520
rect 118030 3500 118060 3520
rect 118140 3500 118170 3520
rect 118250 3500 118280 3530
rect 115470 3450 115530 3470
rect 109320 2870 109350 2900
rect 109430 2870 109460 2900
rect 109540 2870 109570 2900
rect 109650 2870 109680 2900
rect 109760 2870 109790 2900
rect 109870 2870 109900 2900
rect 109980 2870 110010 2900
rect 110090 2870 110120 2900
rect 110200 2870 110230 2900
rect 110310 2870 110340 2900
rect 110420 2870 110450 2900
rect 110530 2870 110560 2900
rect 117040 2870 117070 2900
rect 117150 2870 117180 2900
rect 117260 2870 117290 2900
rect 117370 2870 117400 2900
rect 117480 2870 117510 2900
rect 117590 2870 117620 2900
rect 117700 2870 117730 2900
rect 117810 2870 117840 2900
rect 117920 2870 117950 2900
rect 118030 2870 118060 2900
rect 118140 2870 118170 2900
rect 118250 2870 118280 2900
rect 109250 2850 109350 2870
rect 109250 2810 109260 2850
rect 109300 2840 109350 2850
rect 110530 2850 110630 2870
rect 110530 2840 110580 2850
rect 109300 2810 109310 2840
rect 109250 2790 109310 2810
rect 110570 2810 110580 2840
rect 110620 2810 110630 2850
rect 110570 2790 110630 2810
rect 116970 2850 117070 2870
rect 116970 2810 116980 2850
rect 117020 2840 117070 2850
rect 118250 2850 118350 2870
rect 118250 2840 118300 2850
rect 117020 2810 117030 2840
rect 116970 2780 117030 2810
rect 118290 2810 118300 2840
rect 118340 2810 118350 2850
rect 118290 2790 118350 2810
rect 113650 1700 113730 1720
rect 113650 1660 113670 1700
rect 113710 1660 113730 1700
rect 113870 1700 113950 1720
rect 113870 1660 113890 1700
rect 113930 1660 113950 1700
rect 112520 1610 112550 1640
rect 112630 1630 114750 1660
rect 112630 1610 112660 1630
rect 112740 1610 112770 1630
rect 112850 1610 112880 1630
rect 112960 1610 112990 1630
rect 113070 1610 113100 1630
rect 113180 1610 113210 1630
rect 113290 1610 113320 1630
rect 113400 1610 113430 1630
rect 113510 1610 113540 1630
rect 113620 1610 113650 1630
rect 113730 1610 113760 1630
rect 113840 1610 113870 1630
rect 113950 1610 113980 1630
rect 114060 1610 114090 1630
rect 114170 1610 114200 1630
rect 114280 1610 114310 1630
rect 114390 1610 114420 1630
rect 114500 1610 114530 1630
rect 114610 1610 114640 1630
rect 114720 1610 114750 1630
rect 114830 1610 114860 1640
rect 114940 1610 114970 1640
rect 109600 1460 109680 1480
rect 109600 1430 109620 1460
rect 109580 1420 109620 1430
rect 109660 1430 109680 1460
rect 109800 1460 109880 1480
rect 109800 1430 109820 1460
rect 109660 1420 109820 1430
rect 109860 1430 109880 1460
rect 110000 1460 110080 1480
rect 110000 1430 110020 1460
rect 109860 1420 110020 1430
rect 110060 1430 110080 1460
rect 110200 1460 110280 1480
rect 110200 1430 110220 1460
rect 110060 1420 110220 1430
rect 110260 1430 110280 1460
rect 110260 1420 110300 1430
rect 109380 1380 109500 1410
rect 109580 1400 110300 1420
rect 109580 1380 109700 1400
rect 109780 1380 109900 1400
rect 109980 1380 110100 1400
rect 110180 1380 110300 1400
rect 110380 1380 110500 1410
rect 117320 1460 117400 1480
rect 117320 1420 117340 1460
rect 117380 1420 117400 1460
rect 117320 1410 117400 1420
rect 117520 1460 117600 1480
rect 117520 1420 117540 1460
rect 117580 1420 117600 1460
rect 117520 1410 117600 1420
rect 117720 1460 117800 1480
rect 117720 1420 117740 1460
rect 117780 1420 117800 1460
rect 117720 1410 117800 1420
rect 117920 1460 118000 1480
rect 117920 1420 117940 1460
rect 117980 1420 118000 1460
rect 117920 1410 118000 1420
rect 117100 1380 117220 1410
rect 117300 1380 117420 1410
rect 117500 1380 117620 1410
rect 117700 1380 117820 1410
rect 117900 1380 118020 1410
rect 118100 1380 118220 1410
rect 112520 1080 112550 1110
rect 112630 1080 112660 1110
rect 112740 1080 112770 1110
rect 112850 1080 112880 1110
rect 112960 1080 112990 1110
rect 113070 1080 113100 1110
rect 113180 1080 113210 1110
rect 113290 1080 113320 1110
rect 113400 1080 113430 1110
rect 113510 1080 113540 1110
rect 113620 1080 113650 1110
rect 113730 1080 113760 1110
rect 113840 1080 113870 1110
rect 113950 1080 113980 1110
rect 114060 1080 114090 1110
rect 114170 1080 114200 1110
rect 114280 1080 114310 1110
rect 114390 1080 114420 1110
rect 114500 1080 114530 1110
rect 114610 1080 114640 1110
rect 114720 1080 114750 1110
rect 112440 1060 112550 1080
rect 112440 1020 112460 1060
rect 112500 1050 112550 1060
rect 112500 1020 112520 1050
rect 112440 1000 112520 1020
rect 114830 700 114860 1110
rect 114940 1080 114970 1110
rect 114940 1060 115050 1080
rect 114940 1050 114990 1060
rect 114970 1020 114990 1050
rect 115030 1020 115050 1060
rect 114970 1000 115050 1020
rect 114830 680 114910 700
rect 114830 640 114850 680
rect 114890 640 114910 680
rect 114830 620 114910 640
rect 113760 190 113840 210
rect 113760 150 113780 190
rect 113820 150 113840 190
rect 113510 100 113540 130
rect 113620 120 113980 150
rect 113620 100 113650 120
rect 113730 100 113760 120
rect 113840 100 113870 120
rect 113950 100 113980 120
rect 114060 100 114090 130
rect 109380 -50 109500 -20
rect 109580 -50 109700 -20
rect 109780 -50 109900 -20
rect 109980 -50 110100 -20
rect 110180 -50 110300 -20
rect 110380 -50 110500 -20
rect 109310 -70 109500 -50
rect 109310 -110 109320 -70
rect 109360 -80 109500 -70
rect 110380 -70 110570 -50
rect 110380 -80 110520 -70
rect 109360 -110 109370 -80
rect 109310 -130 109370 -110
rect 110510 -110 110520 -80
rect 110560 -110 110570 -70
rect 110510 -130 110570 -110
rect 117100 -50 117220 -20
rect 117300 -50 117420 -20
rect 117500 -50 117620 -20
rect 117700 -50 117820 -20
rect 117900 -50 118020 -20
rect 118100 -50 118220 -20
rect 117030 -70 117220 -50
rect 117030 -110 117040 -70
rect 117080 -80 117220 -70
rect 118100 -70 118290 -50
rect 118100 -80 118240 -70
rect 117080 -110 117090 -80
rect 117030 -130 117090 -110
rect 118230 -110 118240 -80
rect 118280 -110 118290 -70
rect 118230 -130 118290 -110
rect 113510 -230 113540 -200
rect 113620 -230 113650 -200
rect 113730 -230 113760 -200
rect 113840 -230 113870 -200
rect 113950 -230 113980 -200
rect 114060 -230 114090 -200
rect 113440 -250 113540 -230
rect 113440 -290 113450 -250
rect 113490 -260 113540 -250
rect 114060 -250 114160 -230
rect 114060 -260 114110 -250
rect 113490 -290 113500 -260
rect 113440 -310 113500 -290
rect 114100 -290 114110 -260
rect 114150 -290 114160 -250
rect 114100 -310 114160 -290
rect 113760 -330 113840 -310
rect 113760 -370 113780 -330
rect 113820 -370 113840 -330
rect 113760 -390 113840 -370
rect 113500 -420 114100 -390
rect 113500 -750 114100 -720
<< polycont >>
rect 109500 9930 109540 9970
rect 109620 9930 109660 9970
rect 109740 9930 109780 9970
rect 109860 9930 109900 9970
rect 109980 9930 110020 9970
rect 110100 9930 110140 9970
rect 110220 9930 110260 9970
rect 110340 9930 110380 9970
rect 110460 9930 110500 9970
rect 110580 9930 110620 9970
rect 116980 9930 117020 9970
rect 117100 9930 117140 9970
rect 117220 9930 117260 9970
rect 117340 9930 117380 9970
rect 117460 9930 117500 9970
rect 117580 9930 117620 9970
rect 117700 9930 117740 9970
rect 117820 9930 117860 9970
rect 117940 9930 117980 9970
rect 118060 9930 118100 9970
rect 111990 9550 112030 9590
rect 112350 9550 112390 9590
rect 114270 9550 114310 9590
rect 114630 9550 114670 9590
rect 115210 9550 115250 9590
rect 115570 9550 115610 9590
rect 109320 9010 109360 9050
rect 110760 9010 110800 9050
rect 112930 9210 112970 9250
rect 113290 9210 113330 9250
rect 116800 9010 116840 9050
rect 118240 9010 118280 9050
rect 112120 8630 112160 8670
rect 113070 8630 113110 8670
rect 114490 8630 114530 8670
rect 115362 8630 115402 8670
rect 109200 8330 109240 8370
rect 110640 8330 110680 8370
rect 116920 8330 116960 8370
rect 118360 8330 118400 8370
rect 113040 8250 113080 8290
rect 113700 8250 113740 8290
rect 113860 8250 113900 8290
rect 114520 8250 114560 8290
rect 113224 7480 113264 7520
rect 109380 7410 109420 7450
rect 109500 7410 109540 7450
rect 109620 7410 109660 7450
rect 109740 7410 109780 7450
rect 109860 7410 109900 7450
rect 109980 7410 110020 7450
rect 110100 7410 110140 7450
rect 110220 7410 110260 7450
rect 110340 7410 110380 7450
rect 113370 7480 113410 7520
rect 113516 7480 113556 7520
rect 114044 7480 114084 7520
rect 114190 7480 114230 7520
rect 114336 7480 114376 7520
rect 110460 7410 110500 7450
rect 117100 7410 117140 7450
rect 117220 7410 117260 7450
rect 117340 7410 117380 7450
rect 117460 7410 117500 7450
rect 117580 7410 117620 7450
rect 117700 7410 117740 7450
rect 117820 7410 117860 7450
rect 117940 7410 117980 7450
rect 118060 7410 118100 7450
rect 118180 7410 118220 7450
rect 109260 6980 109300 7020
rect 110580 6980 110620 7020
rect 116980 6980 117020 7020
rect 118300 6980 118340 7020
rect 113720 6910 113760 6950
rect 113560 6270 113600 6310
rect 114000 6270 114040 6310
rect 112245 5780 112285 5820
rect 112355 5780 112395 5820
rect 112465 5780 112505 5820
rect 112575 5780 112615 5820
rect 112685 5780 112725 5820
rect 112795 5780 112835 5820
rect 112905 5780 112945 5820
rect 113015 5780 113055 5820
rect 113125 5780 113165 5820
rect 113235 5780 113275 5820
rect 114325 5780 114365 5820
rect 114435 5780 114475 5820
rect 114545 5780 114585 5820
rect 114655 5780 114695 5820
rect 114765 5780 114805 5820
rect 114875 5780 114915 5820
rect 114985 5780 115025 5820
rect 115095 5780 115135 5820
rect 115205 5780 115245 5820
rect 115315 5780 115355 5820
rect 109920 5640 109960 5680
rect 109920 5510 109960 5550
rect 109920 5430 109960 5470
rect 117640 5640 117680 5680
rect 117640 5510 117680 5550
rect 117640 5430 117680 5470
rect 109920 5350 109960 5390
rect 112080 5340 112120 5380
rect 113400 5340 113440 5380
rect 114160 5340 114200 5380
rect 115480 5340 115520 5380
rect 117640 5350 117680 5390
rect 109260 4430 109300 4470
rect 110580 4430 110620 4470
rect 116980 4430 117020 4470
rect 118300 4430 118340 4470
rect 112090 3960 112130 4000
rect 113390 3980 113430 4020
rect 110250 3890 110290 3930
rect 113690 3980 113730 4020
rect 113870 3980 113910 4020
rect 114170 3980 114210 4020
rect 115470 3960 115510 4000
rect 117310 3890 117350 3930
rect 110250 3760 110290 3800
rect 110250 3680 110290 3720
rect 110250 3550 110290 3590
rect 117310 3760 117350 3800
rect 117310 3680 117350 3720
rect 117310 3550 117350 3590
rect 112080 3470 112120 3510
rect 113480 3470 113520 3510
rect 114080 3470 114120 3510
rect 115480 3470 115520 3510
rect 109260 2810 109300 2850
rect 110580 2810 110620 2850
rect 116980 2810 117020 2850
rect 118300 2810 118340 2850
rect 113670 1660 113710 1700
rect 113890 1660 113930 1700
rect 109620 1420 109660 1460
rect 109820 1420 109860 1460
rect 110020 1420 110060 1460
rect 110220 1420 110260 1460
rect 117340 1420 117380 1460
rect 117540 1420 117580 1460
rect 117740 1420 117780 1460
rect 117940 1420 117980 1460
rect 112460 1020 112500 1060
rect 114990 1020 115030 1060
rect 114850 640 114890 680
rect 113780 150 113820 190
rect 109320 -110 109360 -70
rect 110520 -110 110560 -70
rect 117040 -110 117080 -70
rect 118240 -110 118280 -70
rect 113450 -290 113490 -250
rect 114110 -290 114150 -250
rect 113780 -370 113820 -330
<< xpolycontact >>
rect 108408 6500 108690 6940
rect 108408 5810 108690 6250
rect 118910 6500 119192 6940
rect 118910 5810 119192 6250
rect 108510 3708 108580 4148
rect 108510 2950 108580 3390
rect 108630 3708 108700 4148
rect 108630 2950 108700 3390
rect 108750 3708 108820 4148
rect 108750 2950 108820 3390
rect 108870 3708 108940 4148
rect 118660 3708 118730 4148
rect 108870 2950 108940 3390
rect 118660 2950 118730 3390
rect 118780 3708 118850 4148
rect 118780 2950 118850 3390
rect 118900 3708 118970 4148
rect 118900 2950 118970 3390
rect 119020 3708 119090 4148
rect 119020 2950 119090 3390
rect 108650 840 108720 1280
rect 108650 -94 108720 346
rect 108770 840 108840 1280
rect 108770 -94 108840 346
rect 118760 840 118830 1280
rect 118760 -94 118830 346
rect 118880 840 118950 1280
rect 118880 -94 118950 346
<< ppolyres >>
rect 108408 6250 108690 6500
rect 118910 6250 119192 6500
<< xpolyres >>
rect 108510 3390 108580 3708
rect 108630 3390 108700 3708
rect 108750 3390 108820 3708
rect 108870 3390 108940 3708
rect 118660 3390 118730 3708
rect 118780 3390 118850 3708
rect 118900 3390 118970 3708
rect 119020 3390 119090 3708
rect 108650 346 108720 840
rect 108770 346 108840 840
rect 118760 346 118830 840
rect 118880 346 118950 840
<< locali >>
rect 109490 9970 109550 9990
rect 109490 9930 109500 9970
rect 109540 9930 109550 9970
rect 109490 9910 109550 9930
rect 109610 9970 109670 9990
rect 109610 9930 109620 9970
rect 109660 9930 109670 9970
rect 109610 9910 109670 9930
rect 109730 9970 109790 9990
rect 109730 9930 109740 9970
rect 109780 9930 109790 9970
rect 109730 9910 109790 9930
rect 109850 9970 109910 9990
rect 109850 9930 109860 9970
rect 109900 9930 109910 9970
rect 109850 9910 109910 9930
rect 109970 9970 110030 9990
rect 109970 9930 109980 9970
rect 110020 9930 110030 9970
rect 109970 9910 110030 9930
rect 110090 9970 110150 9990
rect 110090 9930 110100 9970
rect 110140 9930 110150 9970
rect 110090 9910 110150 9930
rect 110210 9970 110270 9990
rect 110210 9930 110220 9970
rect 110260 9930 110270 9970
rect 110210 9910 110270 9930
rect 110330 9970 110390 9990
rect 110330 9930 110340 9970
rect 110380 9930 110390 9970
rect 110330 9910 110390 9930
rect 110450 9970 110510 9990
rect 110450 9930 110460 9970
rect 110500 9930 110510 9970
rect 110450 9910 110510 9930
rect 110570 9970 110630 9990
rect 110570 9930 110580 9970
rect 110620 9930 110630 9970
rect 110570 9910 110630 9930
rect 116970 9970 117030 9990
rect 116970 9930 116980 9970
rect 117020 9930 117030 9970
rect 116970 9910 117030 9930
rect 117090 9970 117150 9990
rect 117090 9930 117100 9970
rect 117140 9930 117150 9970
rect 117090 9910 117150 9930
rect 117210 9970 117270 9990
rect 117210 9930 117220 9970
rect 117260 9930 117270 9970
rect 117210 9910 117270 9930
rect 117330 9970 117390 9990
rect 117330 9930 117340 9970
rect 117380 9930 117390 9970
rect 117330 9910 117390 9930
rect 117450 9970 117510 9990
rect 117450 9930 117460 9970
rect 117500 9930 117510 9970
rect 117450 9910 117510 9930
rect 117570 9970 117630 9990
rect 117570 9930 117580 9970
rect 117620 9930 117630 9970
rect 117570 9910 117630 9930
rect 117690 9970 117750 9990
rect 117690 9930 117700 9970
rect 117740 9930 117750 9970
rect 117690 9910 117750 9930
rect 117810 9970 117870 9990
rect 117810 9930 117820 9970
rect 117860 9930 117870 9970
rect 117810 9910 117870 9930
rect 117930 9970 117990 9990
rect 117930 9930 117940 9970
rect 117980 9930 117990 9970
rect 117930 9910 117990 9930
rect 118050 9970 118110 9990
rect 118050 9930 118060 9970
rect 118100 9930 118110 9970
rect 118050 9910 118110 9930
rect 109230 9770 109370 9790
rect 109230 9130 109240 9770
rect 109280 9130 109320 9770
rect 109360 9130 109370 9770
rect 109230 9110 109370 9130
rect 109430 9770 109490 9790
rect 109430 9130 109440 9770
rect 109480 9130 109490 9770
rect 109430 9110 109490 9130
rect 109550 9770 109610 9790
rect 109550 9130 109560 9770
rect 109600 9130 109610 9770
rect 109550 9110 109610 9130
rect 109670 9770 109730 9790
rect 109670 9130 109680 9770
rect 109720 9130 109730 9770
rect 109670 9110 109730 9130
rect 109790 9770 109850 9790
rect 109790 9130 109800 9770
rect 109840 9130 109850 9770
rect 109790 9110 109850 9130
rect 109910 9770 109970 9790
rect 109910 9130 109920 9770
rect 109960 9130 109970 9770
rect 109910 9110 109970 9130
rect 110030 9770 110090 9790
rect 110030 9130 110040 9770
rect 110080 9130 110090 9770
rect 110030 9110 110090 9130
rect 110150 9770 110210 9790
rect 110150 9130 110160 9770
rect 110200 9130 110210 9770
rect 110150 9110 110210 9130
rect 110270 9770 110330 9790
rect 110270 9130 110280 9770
rect 110320 9130 110330 9770
rect 110270 9110 110330 9130
rect 110390 9770 110450 9790
rect 110390 9130 110400 9770
rect 110440 9130 110450 9770
rect 110390 9110 110450 9130
rect 110510 9770 110570 9790
rect 110510 9130 110520 9770
rect 110560 9130 110570 9770
rect 110510 9110 110570 9130
rect 110630 9770 110690 9790
rect 110630 9130 110640 9770
rect 110680 9130 110690 9770
rect 110630 9110 110690 9130
rect 110750 9770 110890 9790
rect 110750 9130 110760 9770
rect 110800 9130 110840 9770
rect 110880 9130 110890 9770
rect 116710 9770 116850 9790
rect 111970 9590 112050 9610
rect 111970 9550 111990 9590
rect 112030 9550 112050 9590
rect 111970 9530 112050 9550
rect 112330 9590 112410 9610
rect 112330 9550 112350 9590
rect 112390 9550 112410 9590
rect 112330 9530 112410 9550
rect 114250 9590 114330 9610
rect 114250 9550 114270 9590
rect 114310 9550 114330 9590
rect 114250 9530 114330 9550
rect 114610 9590 114690 9610
rect 114610 9550 114630 9590
rect 114670 9550 114690 9590
rect 114610 9530 114690 9550
rect 115190 9590 115270 9610
rect 115190 9550 115210 9590
rect 115250 9550 115270 9590
rect 115190 9530 115270 9550
rect 115550 9590 115630 9610
rect 115550 9550 115570 9590
rect 115610 9550 115630 9590
rect 115550 9530 115630 9550
rect 110750 9110 110890 9130
rect 111900 9470 112040 9490
rect 109300 9050 109380 9070
rect 109300 9010 109320 9050
rect 109360 9010 109380 9050
rect 109300 8990 109380 9010
rect 110740 9050 110820 9070
rect 110740 9010 110760 9050
rect 110800 9010 110820 9050
rect 110740 8990 110820 9010
rect 111900 8830 111910 9470
rect 111950 8830 111990 9470
rect 112030 8830 112040 9470
rect 111900 8810 112040 8830
rect 112100 9470 112160 9490
rect 112100 8830 112110 9470
rect 112150 8830 112160 9470
rect 112100 8810 112160 8830
rect 112220 9470 112280 9490
rect 112220 8830 112230 9470
rect 112270 8830 112280 9470
rect 112220 8810 112280 8830
rect 112340 9470 112480 9490
rect 112340 8830 112350 9470
rect 112390 8830 112430 9470
rect 112470 8830 112480 9470
rect 114180 9470 114320 9490
rect 112910 9250 112990 9270
rect 112910 9210 112930 9250
rect 112970 9210 112990 9250
rect 112910 9190 112990 9210
rect 113270 9250 113350 9270
rect 113270 9210 113290 9250
rect 113330 9210 113350 9250
rect 113270 9190 113350 9210
rect 112340 8810 112480 8830
rect 112840 9130 112980 9150
rect 112840 8830 112850 9130
rect 112890 8830 112930 9130
rect 112970 8830 112980 9130
rect 112840 8810 112980 8830
rect 113040 9130 113100 9150
rect 113040 8830 113050 9130
rect 113090 8830 113100 9130
rect 113040 8810 113100 8830
rect 113160 9130 113220 9150
rect 113160 8830 113170 9130
rect 113210 8830 113220 9130
rect 113160 8810 113220 8830
rect 113280 9130 113420 9150
rect 113280 8830 113290 9130
rect 113330 8830 113370 9130
rect 113410 8830 113420 9130
rect 113280 8810 113420 8830
rect 114180 8830 114190 9470
rect 114230 8830 114270 9470
rect 114310 8830 114320 9470
rect 114180 8810 114320 8830
rect 114380 9470 114440 9490
rect 114380 8830 114390 9470
rect 114430 8830 114440 9470
rect 114380 8810 114440 8830
rect 114500 9470 114560 9490
rect 114500 8830 114510 9470
rect 114550 8830 114560 9470
rect 114500 8810 114560 8830
rect 114620 9470 114760 9490
rect 114620 8830 114630 9470
rect 114670 8830 114710 9470
rect 114750 8830 114760 9470
rect 114620 8810 114760 8830
rect 115120 9470 115260 9490
rect 115120 8830 115130 9470
rect 115170 8830 115210 9470
rect 115250 8830 115260 9470
rect 115120 8810 115260 8830
rect 115320 9470 115380 9490
rect 115320 8830 115330 9470
rect 115370 8830 115380 9470
rect 115320 8810 115380 8830
rect 115440 9470 115500 9490
rect 115440 8830 115450 9470
rect 115490 8830 115500 9470
rect 115440 8810 115500 8830
rect 115560 9470 115700 9490
rect 115560 8830 115570 9470
rect 115610 8830 115650 9470
rect 115690 8830 115700 9470
rect 116710 9130 116720 9770
rect 116760 9130 116800 9770
rect 116840 9130 116850 9770
rect 116710 9110 116850 9130
rect 116910 9770 116970 9790
rect 116910 9130 116920 9770
rect 116960 9130 116970 9770
rect 116910 9110 116970 9130
rect 117030 9770 117090 9790
rect 117030 9130 117040 9770
rect 117080 9130 117090 9770
rect 117030 9110 117090 9130
rect 117150 9770 117210 9790
rect 117150 9130 117160 9770
rect 117200 9130 117210 9770
rect 117150 9110 117210 9130
rect 117270 9770 117330 9790
rect 117270 9130 117280 9770
rect 117320 9130 117330 9770
rect 117270 9110 117330 9130
rect 117390 9770 117450 9790
rect 117390 9130 117400 9770
rect 117440 9130 117450 9770
rect 117390 9110 117450 9130
rect 117510 9770 117570 9790
rect 117510 9130 117520 9770
rect 117560 9130 117570 9770
rect 117510 9110 117570 9130
rect 117630 9770 117690 9790
rect 117630 9130 117640 9770
rect 117680 9130 117690 9770
rect 117630 9110 117690 9130
rect 117750 9770 117810 9790
rect 117750 9130 117760 9770
rect 117800 9130 117810 9770
rect 117750 9110 117810 9130
rect 117870 9770 117930 9790
rect 117870 9130 117880 9770
rect 117920 9130 117930 9770
rect 117870 9110 117930 9130
rect 117990 9770 118050 9790
rect 117990 9130 118000 9770
rect 118040 9130 118050 9770
rect 117990 9110 118050 9130
rect 118110 9770 118170 9790
rect 118110 9130 118120 9770
rect 118160 9130 118170 9770
rect 118110 9110 118170 9130
rect 118230 9770 118370 9790
rect 118230 9130 118240 9770
rect 118280 9130 118320 9770
rect 118360 9130 118370 9770
rect 118230 9110 118370 9130
rect 116780 9050 116860 9070
rect 116780 9010 116800 9050
rect 116840 9010 116860 9050
rect 116780 8990 116860 9010
rect 118220 9050 118300 9070
rect 118220 9010 118240 9050
rect 118280 9010 118300 9050
rect 118220 8990 118300 9010
rect 115560 8810 115700 8830
rect 112100 8670 112180 8690
rect 112100 8630 112120 8670
rect 112160 8630 112180 8670
rect 112100 8610 112180 8630
rect 113060 8670 113120 8690
rect 113060 8630 113070 8670
rect 113110 8630 113120 8670
rect 113060 8610 113120 8630
rect 114480 8670 114540 8690
rect 114480 8630 114490 8670
rect 114530 8630 114540 8670
rect 114480 8610 114540 8630
rect 115352 8670 115412 8690
rect 115352 8630 115362 8670
rect 115402 8630 115412 8670
rect 115352 8610 115412 8630
rect 109190 8370 109250 8390
rect 109190 8330 109200 8370
rect 109240 8330 109250 8370
rect 109190 8310 109250 8330
rect 110630 8370 110690 8390
rect 110630 8330 110640 8370
rect 110680 8330 110690 8370
rect 110630 8310 110690 8330
rect 116910 8370 116970 8390
rect 116910 8330 116920 8370
rect 116960 8330 116970 8370
rect 116910 8310 116970 8330
rect 118350 8370 118410 8390
rect 118350 8330 118360 8370
rect 118400 8330 118410 8370
rect 118350 8310 118410 8330
rect 113020 8290 113100 8310
rect 109110 8250 109250 8270
rect 109110 7610 109120 8250
rect 109160 7610 109200 8250
rect 109240 7610 109250 8250
rect 109110 7590 109250 7610
rect 109310 8250 109370 8270
rect 109310 7610 109320 8250
rect 109360 7610 109370 8250
rect 109310 7590 109370 7610
rect 109430 8250 109490 8270
rect 109430 7610 109440 8250
rect 109480 7610 109490 8250
rect 109430 7590 109490 7610
rect 109550 8250 109610 8270
rect 109550 7610 109560 8250
rect 109600 7610 109610 8250
rect 109550 7590 109610 7610
rect 109670 8250 109730 8270
rect 109670 7610 109680 8250
rect 109720 7610 109730 8250
rect 109670 7590 109730 7610
rect 109790 8250 109850 8270
rect 109790 7610 109800 8250
rect 109840 7610 109850 8250
rect 109790 7590 109850 7610
rect 109910 8250 109970 8270
rect 109910 7610 109920 8250
rect 109960 7610 109970 8250
rect 109910 7590 109970 7610
rect 110030 8250 110090 8270
rect 110030 7610 110040 8250
rect 110080 7610 110090 8250
rect 110030 7590 110090 7610
rect 110150 8250 110210 8270
rect 110150 7610 110160 8250
rect 110200 7610 110210 8250
rect 110150 7590 110210 7610
rect 110270 8250 110330 8270
rect 110270 7610 110280 8250
rect 110320 7610 110330 8250
rect 110270 7590 110330 7610
rect 110390 8250 110450 8270
rect 110390 7610 110400 8250
rect 110440 7610 110450 8250
rect 110390 7590 110450 7610
rect 110510 8250 110570 8270
rect 110510 7610 110520 8250
rect 110560 7610 110570 8250
rect 110510 7590 110570 7610
rect 110630 8250 110770 8270
rect 110630 7610 110640 8250
rect 110680 7610 110720 8250
rect 110760 7610 110770 8250
rect 113020 8250 113040 8290
rect 113080 8250 113100 8290
rect 113020 8230 113100 8250
rect 113360 8290 113420 8310
rect 113360 8250 113370 8290
rect 113410 8250 113420 8290
rect 113360 8230 113420 8250
rect 113680 8290 113760 8310
rect 113680 8250 113700 8290
rect 113740 8250 113760 8290
rect 113680 8230 113760 8250
rect 113840 8290 113920 8310
rect 113840 8250 113860 8290
rect 113900 8250 113920 8290
rect 113840 8230 113920 8250
rect 114180 8290 114240 8310
rect 114180 8250 114190 8290
rect 114230 8250 114240 8290
rect 114180 8230 114240 8250
rect 114500 8290 114580 8310
rect 114500 8250 114520 8290
rect 114560 8250 114580 8290
rect 114500 8230 114580 8250
rect 116830 8250 116970 8270
rect 113040 8060 113080 8230
rect 113240 8160 113320 8180
rect 113240 8120 113260 8160
rect 113300 8120 113320 8160
rect 113240 8100 113320 8120
rect 113260 8060 113300 8100
rect 113370 8060 113410 8230
rect 113460 8160 113540 8180
rect 113460 8120 113480 8160
rect 113520 8120 113540 8160
rect 113460 8100 113540 8120
rect 113480 8060 113520 8100
rect 113700 8060 113740 8230
rect 113860 8060 113900 8230
rect 114060 8160 114140 8180
rect 114060 8120 114080 8160
rect 114120 8120 114140 8160
rect 114060 8100 114140 8120
rect 114080 8060 114120 8100
rect 114190 8060 114230 8230
rect 114280 8160 114360 8180
rect 114280 8120 114300 8160
rect 114340 8120 114360 8160
rect 114280 8100 114360 8120
rect 114300 8060 114340 8100
rect 114520 8060 114560 8230
rect 110630 7590 110770 7610
rect 112950 8040 113090 8060
rect 112950 7600 112960 8040
rect 113000 7600 113040 8040
rect 113080 7600 113090 8040
rect 112950 7580 113090 7600
rect 113140 8040 113200 8060
rect 113140 7600 113150 8040
rect 113190 7600 113200 8040
rect 113140 7580 113200 7600
rect 113250 8040 113310 8060
rect 113250 7600 113260 8040
rect 113300 7600 113310 8040
rect 113250 7580 113310 7600
rect 113360 8040 113420 8060
rect 113360 7600 113370 8040
rect 113410 7600 113420 8040
rect 113360 7580 113420 7600
rect 113470 8040 113530 8060
rect 113470 7600 113480 8040
rect 113520 7600 113530 8040
rect 113470 7580 113530 7600
rect 113580 8040 113640 8060
rect 113580 7600 113590 8040
rect 113630 7600 113640 8040
rect 113580 7580 113640 7600
rect 113690 8040 113910 8060
rect 113690 7600 113700 8040
rect 113740 7600 113780 8040
rect 113820 7600 113860 8040
rect 113900 7600 113910 8040
rect 113690 7580 113910 7600
rect 113960 8040 114020 8060
rect 113960 7600 113970 8040
rect 114010 7600 114020 8040
rect 113960 7580 114020 7600
rect 114070 8040 114130 8060
rect 114070 7600 114080 8040
rect 114120 7600 114130 8040
rect 114070 7580 114130 7600
rect 114180 8040 114240 8060
rect 114180 7600 114190 8040
rect 114230 7600 114240 8040
rect 114180 7580 114240 7600
rect 114290 8040 114350 8060
rect 114290 7600 114300 8040
rect 114340 7600 114350 8040
rect 114290 7580 114350 7600
rect 114400 8040 114460 8060
rect 114400 7600 114410 8040
rect 114450 7600 114460 8040
rect 114400 7580 114460 7600
rect 114510 8040 114650 8060
rect 114510 7600 114520 8040
rect 114560 7600 114600 8040
rect 114640 7600 114650 8040
rect 114510 7580 114650 7600
rect 116830 7610 116840 8250
rect 116880 7610 116920 8250
rect 116960 7610 116970 8250
rect 116830 7590 116970 7610
rect 117030 8250 117090 8270
rect 117030 7610 117040 8250
rect 117080 7610 117090 8250
rect 117030 7590 117090 7610
rect 117150 8250 117210 8270
rect 117150 7610 117160 8250
rect 117200 7610 117210 8250
rect 117150 7590 117210 7610
rect 117270 8250 117330 8270
rect 117270 7610 117280 8250
rect 117320 7610 117330 8250
rect 117270 7590 117330 7610
rect 117390 8250 117450 8270
rect 117390 7610 117400 8250
rect 117440 7610 117450 8250
rect 117390 7590 117450 7610
rect 117510 8250 117570 8270
rect 117510 7610 117520 8250
rect 117560 7610 117570 8250
rect 117510 7590 117570 7610
rect 117630 8250 117690 8270
rect 117630 7610 117640 8250
rect 117680 7610 117690 8250
rect 117630 7590 117690 7610
rect 117750 8250 117810 8270
rect 117750 7610 117760 8250
rect 117800 7610 117810 8250
rect 117750 7590 117810 7610
rect 117870 8250 117930 8270
rect 117870 7610 117880 8250
rect 117920 7610 117930 8250
rect 117870 7590 117930 7610
rect 117990 8250 118050 8270
rect 117990 7610 118000 8250
rect 118040 7610 118050 8250
rect 117990 7590 118050 7610
rect 118110 8250 118170 8270
rect 118110 7610 118120 8250
rect 118160 7610 118170 8250
rect 118110 7590 118170 7610
rect 118230 8250 118290 8270
rect 118230 7610 118240 8250
rect 118280 7610 118290 8250
rect 118230 7590 118290 7610
rect 118350 8250 118490 8270
rect 118350 7610 118360 8250
rect 118400 7610 118440 8250
rect 118480 7610 118490 8250
rect 118350 7590 118490 7610
rect 113140 7560 113180 7580
rect 113120 7540 113180 7560
rect 113600 7560 113640 7580
rect 113960 7560 114000 7580
rect 113600 7540 113660 7560
rect 113120 7500 113130 7540
rect 113170 7500 113180 7540
rect 113120 7480 113180 7500
rect 113214 7520 113274 7540
rect 113214 7480 113224 7520
rect 113264 7480 113274 7520
rect 109370 7450 109430 7470
rect 109370 7410 109380 7450
rect 109420 7410 109430 7450
rect 109370 7390 109430 7410
rect 109490 7450 109550 7470
rect 109490 7410 109500 7450
rect 109540 7410 109550 7450
rect 109490 7390 109550 7410
rect 109610 7450 109670 7470
rect 109610 7410 109620 7450
rect 109660 7410 109670 7450
rect 109610 7390 109670 7410
rect 109730 7450 109790 7470
rect 109730 7410 109740 7450
rect 109780 7410 109790 7450
rect 109730 7390 109790 7410
rect 109850 7450 109910 7470
rect 109850 7410 109860 7450
rect 109900 7410 109910 7450
rect 109850 7390 109910 7410
rect 109970 7450 110030 7470
rect 109970 7410 109980 7450
rect 110020 7410 110030 7450
rect 109970 7390 110030 7410
rect 110090 7450 110150 7470
rect 110090 7410 110100 7450
rect 110140 7410 110150 7450
rect 110090 7390 110150 7410
rect 110210 7450 110270 7470
rect 110210 7410 110220 7450
rect 110260 7410 110270 7450
rect 110210 7390 110270 7410
rect 110330 7450 110390 7470
rect 110330 7410 110340 7450
rect 110380 7410 110390 7450
rect 110330 7390 110390 7410
rect 110450 7450 110510 7470
rect 113214 7460 113274 7480
rect 113350 7520 113430 7540
rect 113350 7480 113370 7520
rect 113410 7480 113430 7520
rect 113350 7460 113430 7480
rect 113506 7520 113566 7540
rect 113506 7480 113516 7520
rect 113556 7480 113566 7520
rect 113600 7500 113610 7540
rect 113650 7500 113660 7540
rect 113600 7480 113660 7500
rect 113940 7540 114000 7560
rect 114420 7560 114460 7580
rect 114420 7540 114480 7560
rect 113940 7500 113950 7540
rect 113990 7500 114000 7540
rect 113940 7480 114000 7500
rect 114034 7520 114094 7540
rect 114034 7480 114044 7520
rect 114084 7480 114094 7520
rect 113506 7460 113566 7480
rect 114034 7460 114094 7480
rect 114170 7520 114250 7540
rect 114170 7480 114190 7520
rect 114230 7480 114250 7520
rect 114170 7460 114250 7480
rect 114326 7520 114386 7540
rect 114326 7480 114336 7520
rect 114376 7480 114386 7520
rect 114420 7500 114430 7540
rect 114470 7500 114480 7540
rect 114420 7480 114480 7500
rect 114326 7460 114386 7480
rect 110450 7410 110460 7450
rect 110500 7410 110510 7450
rect 117090 7450 117150 7470
rect 110450 7390 110510 7410
rect 113200 7400 113280 7420
rect 113200 7360 113220 7400
rect 113260 7360 113280 7400
rect 113200 7340 113280 7360
rect 114320 7400 114400 7420
rect 114320 7360 114340 7400
rect 114380 7360 114400 7400
rect 117090 7410 117100 7450
rect 117140 7410 117150 7450
rect 117090 7390 117150 7410
rect 117210 7450 117270 7470
rect 117210 7410 117220 7450
rect 117260 7410 117270 7450
rect 117210 7390 117270 7410
rect 117330 7450 117390 7470
rect 117330 7410 117340 7450
rect 117380 7410 117390 7450
rect 117330 7390 117390 7410
rect 117450 7450 117510 7470
rect 117450 7410 117460 7450
rect 117500 7410 117510 7450
rect 117450 7390 117510 7410
rect 117570 7450 117630 7470
rect 117570 7410 117580 7450
rect 117620 7410 117630 7450
rect 117570 7390 117630 7410
rect 117690 7450 117750 7470
rect 117690 7410 117700 7450
rect 117740 7410 117750 7450
rect 117690 7390 117750 7410
rect 117810 7450 117870 7470
rect 117810 7410 117820 7450
rect 117860 7410 117870 7450
rect 117810 7390 117870 7410
rect 117930 7450 117990 7470
rect 117930 7410 117940 7450
rect 117980 7410 117990 7450
rect 117930 7390 117990 7410
rect 118050 7450 118110 7470
rect 118050 7410 118060 7450
rect 118100 7410 118110 7450
rect 118050 7390 118110 7410
rect 118170 7450 118230 7470
rect 118170 7410 118180 7450
rect 118220 7410 118230 7450
rect 118170 7390 118230 7410
rect 114320 7340 114400 7360
rect 109250 7020 109310 7040
rect 108408 7000 108690 7020
rect 108408 6960 108420 7000
rect 108460 6960 108530 7000
rect 108570 6960 108640 7000
rect 108680 6960 108690 7000
rect 109250 6980 109260 7020
rect 109300 6980 109310 7020
rect 109250 6960 109310 6980
rect 110570 7020 110630 7040
rect 110570 6980 110580 7020
rect 110620 6980 110630 7020
rect 110570 6960 110630 6980
rect 116970 7020 117030 7040
rect 116970 6980 116980 7020
rect 117020 6980 117030 7020
rect 108408 6940 108690 6960
rect 113700 6950 113780 6970
rect 109170 6900 109310 6920
rect 108408 5790 108690 5810
rect 108408 5750 108420 5790
rect 108460 5750 108530 5790
rect 108570 5750 108640 5790
rect 108680 5750 108690 5790
rect 108408 5730 108690 5750
rect 109170 5760 109180 6900
rect 109220 5760 109260 6900
rect 109300 5760 109310 6900
rect 109170 5740 109310 5760
rect 109360 6900 109420 6920
rect 109360 5760 109370 6900
rect 109410 5760 109420 6900
rect 109360 5740 109420 5760
rect 109470 6900 109530 6920
rect 109470 5760 109480 6900
rect 109520 5760 109530 6900
rect 109470 5740 109530 5760
rect 109580 6900 109640 6920
rect 109580 5760 109590 6900
rect 109630 5760 109640 6900
rect 109580 5740 109640 5760
rect 109690 6900 109750 6920
rect 109690 5760 109700 6900
rect 109740 5760 109750 6900
rect 109690 5740 109750 5760
rect 109800 6900 109860 6920
rect 109800 5760 109810 6900
rect 109850 5760 109860 6900
rect 109800 5740 109860 5760
rect 109910 6900 109970 6920
rect 109910 5760 109920 6900
rect 109960 5760 109970 6900
rect 109910 5740 109970 5760
rect 110020 6900 110080 6920
rect 110020 5760 110030 6900
rect 110070 5760 110080 6900
rect 110020 5740 110080 5760
rect 110130 6900 110190 6920
rect 110130 5760 110140 6900
rect 110180 5760 110190 6900
rect 110130 5740 110190 5760
rect 110240 6900 110300 6920
rect 110240 5760 110250 6900
rect 110290 5760 110300 6900
rect 110240 5740 110300 5760
rect 110350 6900 110410 6920
rect 110350 5760 110360 6900
rect 110400 5760 110410 6900
rect 110350 5740 110410 5760
rect 110460 6900 110520 6920
rect 110460 5760 110470 6900
rect 110510 5760 110520 6900
rect 110460 5740 110520 5760
rect 110570 6900 110710 6920
rect 110570 5760 110580 6900
rect 110620 5760 110660 6900
rect 110700 5760 110710 6900
rect 113700 6910 113720 6950
rect 113760 6910 113780 6950
rect 113700 6890 113780 6910
rect 113870 6950 113950 6970
rect 116970 6960 117030 6980
rect 118290 7020 118350 7040
rect 118290 6980 118300 7020
rect 118340 6980 118350 7020
rect 118290 6960 118350 6980
rect 118910 7000 119192 7020
rect 118910 6960 118920 7000
rect 118960 6960 119030 7000
rect 119070 6960 119140 7000
rect 119180 6960 119192 7000
rect 113870 6910 113890 6950
rect 113930 6910 113950 6950
rect 118910 6940 119192 6960
rect 113870 6890 113950 6910
rect 116890 6900 117030 6920
rect 113470 6830 113610 6850
rect 113470 6390 113480 6830
rect 113520 6390 113560 6830
rect 113600 6390 113610 6830
rect 113470 6370 113610 6390
rect 113660 6830 113720 6850
rect 113660 6390 113670 6830
rect 113710 6390 113720 6830
rect 113660 6370 113720 6390
rect 113770 6830 113830 6850
rect 113770 6390 113780 6830
rect 113820 6390 113830 6830
rect 113770 6370 113830 6390
rect 113880 6830 113940 6850
rect 113880 6390 113890 6830
rect 113930 6390 113940 6830
rect 113880 6370 113940 6390
rect 113990 6830 114130 6850
rect 113990 6390 114000 6830
rect 114040 6390 114080 6830
rect 114120 6390 114130 6830
rect 113990 6370 114130 6390
rect 113540 6310 113620 6330
rect 113540 6270 113560 6310
rect 113600 6270 113620 6310
rect 113540 6250 113620 6270
rect 113980 6310 114060 6330
rect 113980 6270 114000 6310
rect 114040 6270 114060 6310
rect 113980 6250 114060 6270
rect 112232 5820 112298 5840
rect 112232 5780 112245 5820
rect 112285 5780 112298 5820
rect 112232 5760 112298 5780
rect 112342 5820 112408 5840
rect 112342 5780 112355 5820
rect 112395 5780 112408 5820
rect 112342 5760 112408 5780
rect 112452 5820 112518 5840
rect 112452 5780 112465 5820
rect 112505 5780 112518 5820
rect 112452 5760 112518 5780
rect 112562 5820 112628 5840
rect 112562 5780 112575 5820
rect 112615 5780 112628 5820
rect 112562 5760 112628 5780
rect 112672 5820 112738 5840
rect 112672 5780 112685 5820
rect 112725 5780 112738 5820
rect 112672 5760 112738 5780
rect 112782 5820 112848 5840
rect 112782 5780 112795 5820
rect 112835 5780 112848 5820
rect 112782 5760 112848 5780
rect 112892 5820 112958 5840
rect 112892 5780 112905 5820
rect 112945 5780 112958 5820
rect 112892 5760 112958 5780
rect 113002 5820 113068 5840
rect 113002 5780 113015 5820
rect 113055 5780 113068 5820
rect 113002 5760 113068 5780
rect 113112 5820 113178 5840
rect 113112 5780 113125 5820
rect 113165 5780 113178 5820
rect 113112 5760 113178 5780
rect 113222 5820 113288 5840
rect 113222 5780 113235 5820
rect 113275 5780 113288 5820
rect 113222 5760 113288 5780
rect 114312 5820 114378 5840
rect 114312 5780 114325 5820
rect 114365 5780 114378 5820
rect 114312 5760 114378 5780
rect 114422 5820 114488 5840
rect 114422 5780 114435 5820
rect 114475 5780 114488 5820
rect 114422 5760 114488 5780
rect 114532 5820 114598 5840
rect 114532 5780 114545 5820
rect 114585 5780 114598 5820
rect 114532 5760 114598 5780
rect 114642 5820 114708 5840
rect 114642 5780 114655 5820
rect 114695 5780 114708 5820
rect 114642 5760 114708 5780
rect 114752 5820 114818 5840
rect 114752 5780 114765 5820
rect 114805 5780 114818 5820
rect 114752 5760 114818 5780
rect 114862 5820 114928 5840
rect 114862 5780 114875 5820
rect 114915 5780 114928 5820
rect 114862 5760 114928 5780
rect 114972 5820 115038 5840
rect 114972 5780 114985 5820
rect 115025 5780 115038 5820
rect 114972 5760 115038 5780
rect 115082 5820 115148 5840
rect 115082 5780 115095 5820
rect 115135 5780 115148 5820
rect 115082 5760 115148 5780
rect 115192 5820 115258 5840
rect 115192 5780 115205 5820
rect 115245 5780 115258 5820
rect 115192 5760 115258 5780
rect 115302 5820 115368 5840
rect 115302 5780 115315 5820
rect 115355 5780 115368 5820
rect 115302 5760 115368 5780
rect 116890 5760 116900 6900
rect 116940 5760 116980 6900
rect 117020 5760 117030 6900
rect 110570 5740 110710 5760
rect 116890 5740 117030 5760
rect 117080 6900 117140 6920
rect 117080 5760 117090 6900
rect 117130 5760 117140 6900
rect 117080 5740 117140 5760
rect 117190 6900 117250 6920
rect 117190 5760 117200 6900
rect 117240 5760 117250 6900
rect 117190 5740 117250 5760
rect 117300 6900 117360 6920
rect 117300 5760 117310 6900
rect 117350 5760 117360 6900
rect 117300 5740 117360 5760
rect 117410 6900 117470 6920
rect 117410 5760 117420 6900
rect 117460 5760 117470 6900
rect 117410 5740 117470 5760
rect 117520 6900 117580 6920
rect 117520 5760 117530 6900
rect 117570 5760 117580 6900
rect 117520 5740 117580 5760
rect 117630 6900 117690 6920
rect 117630 5760 117640 6900
rect 117680 5760 117690 6900
rect 117630 5740 117690 5760
rect 117740 6900 117800 6920
rect 117740 5760 117750 6900
rect 117790 5760 117800 6900
rect 117740 5740 117800 5760
rect 117850 6900 117910 6920
rect 117850 5760 117860 6900
rect 117900 5760 117910 6900
rect 117850 5740 117910 5760
rect 117960 6900 118020 6920
rect 117960 5760 117970 6900
rect 118010 5760 118020 6900
rect 117960 5740 118020 5760
rect 118070 6900 118130 6920
rect 118070 5760 118080 6900
rect 118120 5760 118130 6900
rect 118070 5740 118130 5760
rect 118180 6900 118240 6920
rect 118180 5760 118190 6900
rect 118230 5760 118240 6900
rect 118180 5740 118240 5760
rect 118290 6900 118430 6920
rect 118290 5760 118300 6900
rect 118340 5760 118380 6900
rect 118420 5760 118430 6900
rect 118290 5740 118430 5760
rect 118910 5790 119192 5810
rect 118910 5750 118920 5790
rect 118960 5750 119030 5790
rect 119070 5750 119140 5790
rect 119180 5750 119192 5790
rect 118910 5730 119192 5750
rect 111990 5700 112130 5720
rect 109910 5680 109970 5700
rect 109910 5640 109920 5680
rect 109960 5640 109970 5680
rect 109910 5620 109970 5640
rect 109900 5550 109980 5570
rect 109900 5510 109920 5550
rect 109960 5510 109980 5550
rect 109900 5470 109980 5510
rect 109900 5430 109920 5470
rect 109960 5430 109980 5470
rect 111990 5460 112000 5700
rect 112040 5460 112080 5700
rect 112120 5460 112130 5700
rect 111990 5440 112130 5460
rect 112180 5700 112240 5720
rect 112180 5460 112190 5700
rect 112230 5460 112240 5700
rect 112180 5440 112240 5460
rect 112290 5700 112350 5720
rect 112290 5460 112300 5700
rect 112340 5460 112350 5700
rect 112290 5440 112350 5460
rect 112400 5700 112460 5720
rect 112400 5460 112410 5700
rect 112450 5460 112460 5700
rect 112400 5440 112460 5460
rect 112510 5700 112570 5720
rect 112510 5460 112520 5700
rect 112560 5460 112570 5700
rect 112510 5440 112570 5460
rect 112620 5700 112680 5720
rect 112620 5460 112630 5700
rect 112670 5460 112680 5700
rect 112620 5440 112680 5460
rect 112730 5700 112790 5720
rect 112730 5460 112740 5700
rect 112780 5460 112790 5700
rect 112730 5440 112790 5460
rect 112840 5700 112900 5720
rect 112840 5460 112850 5700
rect 112890 5460 112900 5700
rect 112840 5440 112900 5460
rect 112950 5700 113010 5720
rect 112950 5460 112960 5700
rect 113000 5460 113010 5700
rect 112950 5440 113010 5460
rect 113060 5700 113120 5720
rect 113060 5460 113070 5700
rect 113110 5460 113120 5700
rect 113060 5440 113120 5460
rect 113170 5700 113230 5720
rect 113170 5460 113180 5700
rect 113220 5460 113230 5700
rect 113170 5440 113230 5460
rect 113280 5700 113340 5720
rect 113280 5460 113290 5700
rect 113330 5460 113340 5700
rect 113280 5440 113340 5460
rect 113390 5700 113530 5720
rect 113390 5460 113400 5700
rect 113440 5460 113480 5700
rect 113520 5460 113530 5700
rect 113390 5440 113530 5460
rect 114070 5700 114210 5720
rect 114070 5460 114080 5700
rect 114120 5460 114160 5700
rect 114200 5460 114210 5700
rect 114070 5440 114210 5460
rect 114260 5700 114320 5720
rect 114260 5460 114270 5700
rect 114310 5460 114320 5700
rect 114260 5440 114320 5460
rect 114370 5700 114430 5720
rect 114370 5460 114380 5700
rect 114420 5460 114430 5700
rect 114370 5440 114430 5460
rect 114480 5700 114540 5720
rect 114480 5460 114490 5700
rect 114530 5460 114540 5700
rect 114480 5440 114540 5460
rect 114590 5700 114650 5720
rect 114590 5460 114600 5700
rect 114640 5460 114650 5700
rect 114590 5440 114650 5460
rect 114700 5700 114760 5720
rect 114700 5460 114710 5700
rect 114750 5460 114760 5700
rect 114700 5440 114760 5460
rect 114810 5700 114870 5720
rect 114810 5460 114820 5700
rect 114860 5460 114870 5700
rect 114810 5440 114870 5460
rect 114920 5700 114980 5720
rect 114920 5460 114930 5700
rect 114970 5460 114980 5700
rect 114920 5440 114980 5460
rect 115030 5700 115090 5720
rect 115030 5460 115040 5700
rect 115080 5460 115090 5700
rect 115030 5440 115090 5460
rect 115140 5700 115200 5720
rect 115140 5460 115150 5700
rect 115190 5460 115200 5700
rect 115140 5440 115200 5460
rect 115250 5700 115310 5720
rect 115250 5460 115260 5700
rect 115300 5460 115310 5700
rect 115250 5440 115310 5460
rect 115360 5700 115420 5720
rect 115360 5460 115370 5700
rect 115410 5460 115420 5700
rect 115360 5440 115420 5460
rect 115470 5700 115610 5720
rect 115470 5460 115480 5700
rect 115520 5460 115560 5700
rect 115600 5460 115610 5700
rect 117630 5680 117690 5700
rect 117630 5640 117640 5680
rect 117680 5640 117690 5680
rect 117630 5620 117690 5640
rect 115470 5440 115610 5460
rect 117620 5550 117700 5570
rect 117620 5510 117640 5550
rect 117680 5510 117700 5550
rect 117620 5470 117700 5510
rect 109900 5390 109980 5430
rect 109900 5350 109920 5390
rect 109960 5350 109980 5390
rect 109900 5330 109980 5350
rect 112070 5380 112130 5440
rect 112070 5340 112080 5380
rect 112120 5340 112130 5380
rect 112070 5320 112130 5340
rect 113390 5380 113450 5400
rect 113390 5340 113400 5380
rect 113440 5340 113450 5380
rect 113390 5320 113450 5340
rect 114150 5380 114210 5400
rect 114150 5340 114160 5380
rect 114200 5340 114210 5380
rect 114150 5320 114210 5340
rect 115470 5380 115530 5440
rect 115470 5340 115480 5380
rect 115520 5340 115530 5380
rect 115470 5320 115530 5340
rect 117620 5430 117640 5470
rect 117680 5430 117700 5470
rect 117620 5390 117700 5430
rect 117620 5350 117640 5390
rect 117680 5350 117700 5390
rect 117620 5330 117700 5350
rect 109250 4470 109310 4490
rect 109250 4430 109260 4470
rect 109300 4430 109310 4470
rect 109250 4410 109310 4430
rect 110570 4470 110630 4490
rect 110570 4430 110580 4470
rect 110620 4430 110630 4470
rect 110570 4410 110630 4430
rect 116970 4470 117030 4490
rect 116970 4430 116980 4470
rect 117020 4430 117030 4470
rect 116970 4410 117030 4430
rect 118290 4470 118350 4490
rect 118290 4430 118300 4470
rect 118340 4430 118350 4470
rect 118290 4410 118350 4430
rect 109170 4350 109310 4370
rect 108510 4182 108940 4222
rect 108510 4148 108580 4182
rect 108870 4148 108940 4182
rect 108700 4048 108750 4148
rect 109170 4010 109180 4350
rect 109220 4010 109260 4350
rect 109300 4010 109310 4350
rect 109170 3990 109310 4010
rect 109360 4350 109420 4370
rect 109360 4010 109370 4350
rect 109410 4010 109420 4350
rect 109360 3990 109420 4010
rect 109470 4350 109530 4370
rect 109470 4010 109480 4350
rect 109520 4010 109530 4350
rect 109470 3990 109530 4010
rect 109580 4350 109640 4370
rect 109580 4010 109590 4350
rect 109630 4010 109640 4350
rect 109580 3990 109640 4010
rect 109690 4350 109750 4370
rect 109690 4010 109700 4350
rect 109740 4010 109750 4350
rect 109690 3990 109750 4010
rect 109800 4350 109860 4370
rect 109800 4010 109810 4350
rect 109850 4010 109860 4350
rect 109800 3990 109860 4010
rect 109910 4350 109970 4370
rect 109910 4010 109920 4350
rect 109960 4010 109970 4350
rect 109910 3990 109970 4010
rect 110020 4350 110080 4370
rect 110020 4010 110030 4350
rect 110070 4010 110080 4350
rect 110020 3990 110080 4010
rect 110130 4350 110190 4370
rect 110130 4010 110140 4350
rect 110180 4010 110190 4350
rect 110130 3990 110190 4010
rect 110240 4350 110300 4370
rect 110240 4010 110250 4350
rect 110290 4010 110300 4350
rect 110240 3990 110300 4010
rect 110350 4350 110410 4370
rect 110350 4010 110360 4350
rect 110400 4010 110410 4350
rect 110350 3990 110410 4010
rect 110460 4350 110520 4370
rect 110460 4010 110470 4350
rect 110510 4010 110520 4350
rect 110460 3990 110520 4010
rect 110570 4350 110710 4370
rect 110570 4010 110580 4350
rect 110620 4010 110660 4350
rect 110700 4010 110710 4350
rect 116890 4350 117030 4370
rect 113380 4020 113440 4040
rect 110570 3990 110710 4010
rect 112080 4000 112140 4020
rect 112080 3960 112090 4000
rect 112130 3960 112140 4000
rect 113380 3980 113390 4020
rect 113430 3980 113440 4020
rect 113380 3960 113440 3980
rect 113680 4020 113740 4040
rect 113680 3980 113690 4020
rect 113730 3980 113740 4020
rect 113680 3960 113740 3980
rect 113860 4020 113920 4040
rect 113860 3980 113870 4020
rect 113910 3980 113920 4020
rect 113860 3960 113920 3980
rect 114160 4020 114220 4040
rect 114160 3980 114170 4020
rect 114210 3980 114220 4020
rect 114160 3960 114220 3980
rect 115460 4000 115520 4020
rect 115460 3960 115470 4000
rect 115510 3960 115520 4000
rect 116890 4010 116900 4350
rect 116940 4010 116980 4350
rect 117020 4010 117030 4350
rect 116890 3990 117030 4010
rect 117080 4350 117140 4370
rect 117080 4010 117090 4350
rect 117130 4010 117140 4350
rect 117080 3990 117140 4010
rect 117190 4350 117250 4370
rect 117190 4010 117200 4350
rect 117240 4010 117250 4350
rect 117190 3990 117250 4010
rect 117300 4350 117360 4370
rect 117300 4010 117310 4350
rect 117350 4010 117360 4350
rect 117300 3990 117360 4010
rect 117410 4350 117470 4370
rect 117410 4010 117420 4350
rect 117460 4010 117470 4350
rect 117410 3990 117470 4010
rect 117520 4350 117580 4370
rect 117520 4010 117530 4350
rect 117570 4010 117580 4350
rect 117520 3990 117580 4010
rect 117630 4350 117690 4370
rect 117630 4010 117640 4350
rect 117680 4010 117690 4350
rect 117630 3990 117690 4010
rect 117740 4350 117800 4370
rect 117740 4010 117750 4350
rect 117790 4010 117800 4350
rect 117740 3990 117800 4010
rect 117850 4350 117910 4370
rect 117850 4010 117860 4350
rect 117900 4010 117910 4350
rect 117850 3990 117910 4010
rect 117960 4350 118020 4370
rect 117960 4010 117970 4350
rect 118010 4010 118020 4350
rect 117960 3990 118020 4010
rect 118070 4350 118130 4370
rect 118070 4010 118080 4350
rect 118120 4010 118130 4350
rect 118070 3990 118130 4010
rect 118180 4350 118240 4370
rect 118180 4010 118190 4350
rect 118230 4010 118240 4350
rect 118180 3990 118240 4010
rect 118290 4350 118430 4370
rect 118290 4010 118300 4350
rect 118340 4010 118380 4350
rect 118420 4010 118430 4350
rect 118290 3990 118430 4010
rect 118660 4182 119090 4222
rect 118660 4148 118730 4182
rect 119020 4148 119090 4182
rect 109460 3930 109540 3950
rect 109460 3890 109480 3930
rect 109520 3890 109540 3930
rect 109460 3870 109540 3890
rect 109680 3930 109760 3950
rect 109680 3890 109700 3930
rect 109740 3890 109760 3930
rect 109680 3870 109760 3890
rect 109900 3930 109980 3950
rect 109900 3890 109920 3930
rect 109960 3890 109980 3930
rect 109900 3870 109980 3890
rect 110120 3930 110200 3950
rect 110120 3890 110140 3930
rect 110180 3890 110200 3930
rect 110120 3870 110200 3890
rect 110240 3930 110300 3950
rect 110240 3890 110250 3930
rect 110290 3890 110300 3930
rect 110240 3870 110300 3890
rect 110340 3930 110420 3950
rect 112080 3940 112140 3960
rect 115460 3940 115520 3960
rect 110340 3890 110360 3930
rect 110400 3890 110420 3930
rect 110340 3870 110420 3890
rect 117180 3930 117260 3950
rect 117180 3890 117200 3930
rect 117240 3890 117260 3930
rect 117180 3870 117260 3890
rect 117300 3930 117360 3950
rect 117300 3890 117310 3930
rect 117350 3890 117360 3930
rect 117300 3870 117360 3890
rect 117400 3930 117480 3950
rect 117400 3890 117420 3930
rect 117460 3890 117480 3930
rect 117400 3870 117480 3890
rect 117620 3930 117700 3950
rect 117620 3890 117640 3930
rect 117680 3890 117700 3930
rect 117620 3870 117700 3890
rect 117840 3930 117920 3950
rect 117840 3890 117860 3930
rect 117900 3890 117920 3930
rect 117840 3870 117920 3890
rect 118060 3930 118140 3950
rect 118060 3890 118080 3930
rect 118120 3890 118140 3930
rect 118060 3870 118140 3890
rect 111990 3830 112130 3850
rect 110230 3800 110310 3820
rect 110230 3760 110250 3800
rect 110290 3760 110310 3800
rect 110230 3720 110310 3760
rect 110230 3680 110250 3720
rect 110290 3680 110310 3720
rect 110230 3660 110310 3680
rect 110240 3590 110300 3610
rect 110240 3550 110250 3590
rect 110290 3550 110300 3590
rect 111990 3590 112000 3830
rect 112040 3590 112080 3830
rect 112120 3590 112130 3830
rect 111990 3570 112130 3590
rect 112180 3830 112240 3850
rect 112180 3590 112190 3830
rect 112230 3590 112240 3830
rect 112180 3570 112240 3590
rect 112290 3830 112350 3850
rect 112290 3590 112300 3830
rect 112340 3590 112350 3830
rect 112290 3570 112350 3590
rect 112400 3830 112460 3850
rect 112400 3590 112410 3830
rect 112450 3590 112460 3830
rect 112400 3570 112460 3590
rect 112510 3830 112570 3850
rect 112510 3590 112520 3830
rect 112560 3590 112570 3830
rect 112510 3570 112570 3590
rect 112620 3830 112680 3850
rect 112620 3590 112630 3830
rect 112670 3590 112680 3830
rect 112620 3570 112680 3590
rect 112730 3830 112790 3850
rect 112730 3590 112740 3830
rect 112780 3590 112790 3830
rect 112730 3570 112790 3590
rect 112840 3830 112900 3850
rect 112840 3590 112850 3830
rect 112890 3590 112900 3830
rect 112840 3570 112900 3590
rect 112950 3830 113010 3850
rect 112950 3590 112960 3830
rect 113000 3590 113010 3830
rect 112950 3570 113010 3590
rect 113060 3830 113120 3850
rect 113060 3590 113070 3830
rect 113110 3590 113120 3830
rect 113060 3570 113120 3590
rect 113170 3830 113230 3850
rect 113170 3590 113180 3830
rect 113220 3590 113230 3830
rect 113170 3570 113230 3590
rect 113280 3830 113340 3850
rect 113280 3590 113290 3830
rect 113330 3590 113340 3830
rect 113280 3570 113340 3590
rect 113390 3830 113610 3850
rect 113390 3590 113400 3830
rect 113440 3590 113480 3830
rect 113520 3590 113560 3830
rect 113600 3590 113610 3830
rect 113390 3570 113610 3590
rect 113660 3830 113720 3850
rect 113660 3590 113670 3830
rect 113710 3590 113720 3830
rect 113660 3570 113720 3590
rect 113770 3830 113830 3850
rect 113770 3590 113780 3830
rect 113820 3590 113830 3830
rect 113770 3570 113830 3590
rect 113880 3830 113940 3850
rect 113880 3590 113890 3830
rect 113930 3590 113940 3830
rect 113880 3570 113940 3590
rect 113990 3830 114210 3850
rect 113990 3590 114000 3830
rect 114040 3590 114080 3830
rect 114120 3590 114160 3830
rect 114200 3590 114210 3830
rect 113990 3570 114210 3590
rect 114260 3830 114320 3850
rect 114260 3590 114270 3830
rect 114310 3590 114320 3830
rect 114260 3570 114320 3590
rect 114370 3830 114430 3850
rect 114370 3590 114380 3830
rect 114420 3590 114430 3830
rect 114370 3570 114430 3590
rect 114480 3830 114540 3850
rect 114480 3590 114490 3830
rect 114530 3590 114540 3830
rect 114480 3570 114540 3590
rect 114590 3830 114650 3850
rect 114590 3590 114600 3830
rect 114640 3590 114650 3830
rect 114590 3570 114650 3590
rect 114700 3830 114760 3850
rect 114700 3590 114710 3830
rect 114750 3590 114760 3830
rect 114700 3570 114760 3590
rect 114810 3830 114870 3850
rect 114810 3590 114820 3830
rect 114860 3590 114870 3830
rect 114810 3570 114870 3590
rect 114920 3830 114980 3850
rect 114920 3590 114930 3830
rect 114970 3590 114980 3830
rect 114920 3570 114980 3590
rect 115030 3830 115090 3850
rect 115030 3590 115040 3830
rect 115080 3590 115090 3830
rect 115030 3570 115090 3590
rect 115140 3830 115200 3850
rect 115140 3590 115150 3830
rect 115190 3590 115200 3830
rect 115140 3570 115200 3590
rect 115250 3830 115310 3850
rect 115250 3590 115260 3830
rect 115300 3590 115310 3830
rect 115250 3570 115310 3590
rect 115360 3830 115420 3850
rect 115360 3590 115370 3830
rect 115410 3590 115420 3830
rect 115360 3570 115420 3590
rect 115470 3830 115610 3850
rect 115470 3590 115480 3830
rect 115520 3590 115560 3830
rect 115600 3590 115610 3830
rect 117290 3800 117370 3820
rect 117290 3760 117310 3800
rect 117350 3760 117370 3800
rect 117290 3720 117370 3760
rect 117290 3680 117310 3720
rect 117350 3680 117370 3720
rect 118850 4048 118900 4148
rect 117290 3660 117370 3680
rect 115470 3570 115610 3590
rect 117300 3590 117360 3610
rect 110240 3530 110300 3550
rect 112080 3530 112130 3570
rect 112070 3510 112130 3530
rect 109170 3470 109310 3490
rect 108510 2930 108580 2950
rect 108510 2880 108520 2930
rect 108570 2880 108580 2930
rect 108510 2860 108580 2880
rect 108630 2930 108700 2950
rect 108630 2880 108640 2930
rect 108690 2880 108700 2930
rect 108630 2860 108700 2880
rect 108750 2930 108820 2950
rect 108750 2880 108760 2930
rect 108810 2880 108820 2930
rect 108750 2860 108820 2880
rect 108870 2930 108940 2950
rect 108870 2880 108880 2930
rect 108930 2880 108940 2930
rect 109170 2930 109180 3470
rect 109220 2930 109260 3470
rect 109300 2930 109310 3470
rect 109170 2910 109310 2930
rect 109360 3470 109420 3490
rect 109360 2930 109370 3470
rect 109410 2930 109420 3470
rect 109360 2910 109420 2930
rect 109470 3470 109530 3490
rect 109470 2930 109480 3470
rect 109520 2930 109530 3470
rect 109470 2910 109530 2930
rect 109580 3470 109640 3490
rect 109580 2930 109590 3470
rect 109630 2930 109640 3470
rect 109580 2910 109640 2930
rect 109690 3470 109750 3490
rect 109690 2930 109700 3470
rect 109740 2930 109750 3470
rect 109690 2910 109750 2930
rect 109800 3470 109860 3490
rect 109800 2930 109810 3470
rect 109850 2930 109860 3470
rect 109800 2910 109860 2930
rect 109910 3470 109970 3490
rect 109910 2930 109920 3470
rect 109960 2930 109970 3470
rect 109910 2910 109970 2930
rect 110020 3470 110080 3490
rect 110020 2930 110030 3470
rect 110070 2930 110080 3470
rect 110020 2910 110080 2930
rect 110130 3470 110190 3490
rect 110130 2930 110140 3470
rect 110180 2930 110190 3470
rect 110130 2910 110190 2930
rect 110240 3470 110300 3490
rect 110240 2930 110250 3470
rect 110290 2930 110300 3470
rect 110240 2910 110300 2930
rect 110350 3470 110410 3490
rect 110350 2930 110360 3470
rect 110400 2930 110410 3470
rect 110350 2910 110410 2930
rect 110460 3470 110520 3490
rect 110460 2930 110470 3470
rect 110510 2930 110520 3470
rect 110460 2910 110520 2930
rect 110570 3470 110710 3490
rect 110570 2930 110580 3470
rect 110620 2930 110660 3470
rect 110700 2930 110710 3470
rect 112070 3470 112080 3510
rect 112120 3470 112130 3510
rect 112070 3450 112130 3470
rect 113470 3510 113530 3530
rect 113470 3470 113480 3510
rect 113520 3470 113530 3510
rect 113470 3450 113530 3470
rect 114070 3510 114130 3530
rect 114070 3470 114080 3510
rect 114120 3470 114130 3510
rect 114070 3450 114130 3470
rect 115470 3510 115530 3570
rect 117300 3550 117310 3590
rect 117350 3550 117360 3590
rect 117300 3530 117360 3550
rect 115470 3470 115480 3510
rect 115520 3470 115530 3510
rect 115470 3450 115530 3470
rect 116890 3470 117030 3490
rect 110570 2910 110710 2930
rect 116890 2930 116900 3470
rect 116940 2930 116980 3470
rect 117020 2930 117030 3470
rect 116890 2910 117030 2930
rect 117080 3470 117140 3490
rect 117080 2930 117090 3470
rect 117130 2930 117140 3470
rect 117080 2910 117140 2930
rect 117190 3470 117250 3490
rect 117190 2930 117200 3470
rect 117240 2930 117250 3470
rect 117190 2910 117250 2930
rect 117300 3470 117360 3490
rect 117300 2930 117310 3470
rect 117350 2930 117360 3470
rect 117300 2910 117360 2930
rect 117410 3470 117470 3490
rect 117410 2930 117420 3470
rect 117460 2930 117470 3470
rect 117410 2910 117470 2930
rect 117520 3470 117580 3490
rect 117520 2930 117530 3470
rect 117570 2930 117580 3470
rect 117520 2910 117580 2930
rect 117630 3470 117690 3490
rect 117630 2930 117640 3470
rect 117680 2930 117690 3470
rect 117630 2910 117690 2930
rect 117740 3470 117800 3490
rect 117740 2930 117750 3470
rect 117790 2930 117800 3470
rect 117740 2910 117800 2930
rect 117850 3470 117910 3490
rect 117850 2930 117860 3470
rect 117900 2930 117910 3470
rect 117850 2910 117910 2930
rect 117960 3470 118020 3490
rect 117960 2930 117970 3470
rect 118010 2930 118020 3470
rect 117960 2910 118020 2930
rect 118070 3470 118130 3490
rect 118070 2930 118080 3470
rect 118120 2930 118130 3470
rect 118070 2910 118130 2930
rect 118180 3470 118240 3490
rect 118180 2930 118190 3470
rect 118230 2930 118240 3470
rect 118180 2910 118240 2930
rect 118290 3470 118430 3490
rect 118290 2930 118300 3470
rect 118340 2930 118380 3470
rect 118420 2930 118430 3470
rect 118290 2910 118430 2930
rect 118660 2930 118730 2950
rect 108870 2860 108940 2880
rect 118660 2880 118670 2930
rect 118720 2880 118730 2930
rect 109250 2850 109310 2870
rect 109250 2810 109260 2850
rect 109300 2810 109310 2850
rect 109250 2790 109310 2810
rect 110570 2850 110630 2870
rect 110570 2810 110580 2850
rect 110620 2810 110630 2850
rect 110570 2790 110630 2810
rect 116970 2850 117030 2870
rect 116970 2810 116980 2850
rect 117020 2810 117030 2850
rect 116970 2780 117030 2810
rect 118290 2850 118350 2870
rect 118660 2860 118730 2880
rect 118780 2930 118850 2950
rect 118780 2880 118790 2930
rect 118840 2880 118850 2930
rect 118780 2860 118850 2880
rect 118900 2930 118970 2950
rect 118900 2880 118910 2930
rect 118960 2880 118970 2930
rect 118900 2860 118970 2880
rect 119020 2930 119090 2950
rect 119020 2880 119030 2930
rect 119080 2880 119090 2930
rect 119020 2860 119090 2880
rect 118290 2810 118300 2850
rect 118340 2810 118350 2850
rect 118290 2790 118350 2810
rect 113650 1700 113730 1720
rect 113650 1660 113670 1700
rect 113710 1660 113730 1700
rect 113650 1640 113730 1660
rect 113870 1700 113950 1720
rect 113870 1660 113890 1700
rect 113930 1660 113950 1700
rect 113870 1640 113950 1660
rect 112370 1580 112510 1600
rect 109600 1460 109680 1480
rect 109600 1420 109620 1460
rect 109660 1420 109680 1460
rect 109600 1400 109680 1420
rect 109800 1460 109880 1480
rect 109800 1420 109820 1460
rect 109860 1420 109880 1460
rect 109800 1400 109880 1420
rect 110000 1460 110080 1480
rect 110000 1420 110020 1460
rect 110060 1420 110080 1460
rect 110000 1400 110080 1420
rect 110200 1460 110280 1480
rect 110200 1420 110220 1460
rect 110260 1420 110280 1460
rect 110200 1400 110280 1420
rect 108650 1350 108720 1370
rect 108650 1300 108660 1350
rect 108710 1300 108720 1350
rect 108650 1280 108720 1300
rect 108770 1350 108840 1370
rect 108770 1300 108780 1350
rect 108830 1300 108840 1350
rect 108770 1280 108840 1300
rect 109230 1350 109370 1370
rect 108720 -94 108770 6
rect 109230 10 109240 1350
rect 109280 10 109320 1350
rect 109360 10 109370 1350
rect 109230 -10 109370 10
rect 109510 1350 109570 1370
rect 109510 10 109520 1350
rect 109560 10 109570 1350
rect 109510 -10 109570 10
rect 109710 1350 109770 1370
rect 109710 10 109720 1350
rect 109760 10 109770 1350
rect 109710 -10 109770 10
rect 109910 1350 109970 1370
rect 109910 10 109920 1350
rect 109960 10 109970 1350
rect 109910 -10 109970 10
rect 110110 1350 110170 1370
rect 110110 10 110120 1350
rect 110160 10 110170 1350
rect 110110 -10 110170 10
rect 110310 1350 110370 1370
rect 110310 10 110320 1350
rect 110360 10 110370 1350
rect 110310 -10 110370 10
rect 110510 1350 110650 1370
rect 110510 10 110520 1350
rect 110560 10 110600 1350
rect 110640 10 110650 1350
rect 112370 1140 112380 1580
rect 112420 1140 112460 1580
rect 112500 1140 112510 1580
rect 112370 1120 112510 1140
rect 112560 1580 112620 1600
rect 112560 1140 112570 1580
rect 112610 1140 112620 1580
rect 112560 1120 112620 1140
rect 112670 1580 112730 1600
rect 112670 1140 112680 1580
rect 112720 1140 112730 1580
rect 112670 1120 112730 1140
rect 112780 1580 112840 1600
rect 112780 1140 112790 1580
rect 112830 1140 112840 1580
rect 112780 1120 112840 1140
rect 112890 1580 112950 1600
rect 112890 1140 112900 1580
rect 112940 1140 112950 1580
rect 112890 1120 112950 1140
rect 113000 1580 113060 1600
rect 113000 1140 113010 1580
rect 113050 1140 113060 1580
rect 113000 1120 113060 1140
rect 113110 1580 113170 1600
rect 113110 1140 113120 1580
rect 113160 1140 113170 1580
rect 113110 1120 113170 1140
rect 113220 1580 113280 1600
rect 113220 1140 113230 1580
rect 113270 1140 113280 1580
rect 113220 1120 113280 1140
rect 113330 1580 113390 1600
rect 113330 1140 113340 1580
rect 113380 1140 113390 1580
rect 113330 1120 113390 1140
rect 113440 1580 113500 1600
rect 113440 1140 113450 1580
rect 113490 1140 113500 1580
rect 113440 1120 113500 1140
rect 113550 1580 113610 1600
rect 113550 1140 113560 1580
rect 113600 1140 113610 1580
rect 113550 1120 113610 1140
rect 113660 1580 113720 1600
rect 113660 1140 113670 1580
rect 113710 1140 113720 1580
rect 113660 1120 113720 1140
rect 113770 1580 113830 1600
rect 113770 1140 113780 1580
rect 113820 1140 113830 1580
rect 113770 1120 113830 1140
rect 113880 1580 113940 1600
rect 113880 1140 113890 1580
rect 113930 1140 113940 1580
rect 113880 1120 113940 1140
rect 113990 1580 114050 1600
rect 113990 1140 114000 1580
rect 114040 1140 114050 1580
rect 113990 1120 114050 1140
rect 114100 1580 114160 1600
rect 114100 1140 114110 1580
rect 114150 1140 114160 1580
rect 114100 1120 114160 1140
rect 114210 1580 114270 1600
rect 114210 1140 114220 1580
rect 114260 1140 114270 1580
rect 114210 1120 114270 1140
rect 114320 1580 114380 1600
rect 114320 1140 114330 1580
rect 114370 1140 114380 1580
rect 114320 1120 114380 1140
rect 114430 1580 114490 1600
rect 114430 1140 114440 1580
rect 114480 1140 114490 1580
rect 114430 1120 114490 1140
rect 114540 1580 114600 1600
rect 114540 1140 114550 1580
rect 114590 1140 114600 1580
rect 114540 1120 114600 1140
rect 114650 1580 114710 1600
rect 114650 1140 114660 1580
rect 114700 1140 114710 1580
rect 114650 1120 114710 1140
rect 114760 1580 114820 1600
rect 114760 1140 114770 1580
rect 114810 1140 114820 1580
rect 114760 1120 114820 1140
rect 114870 1580 114930 1600
rect 114870 1140 114880 1580
rect 114920 1140 114930 1580
rect 114870 1120 114930 1140
rect 114980 1580 115120 1600
rect 114980 1140 114990 1580
rect 115030 1140 115070 1580
rect 115110 1140 115120 1580
rect 117320 1460 117400 1480
rect 117320 1420 117340 1460
rect 117380 1420 117400 1460
rect 117320 1400 117400 1420
rect 117520 1460 117600 1480
rect 117520 1420 117540 1460
rect 117580 1420 117600 1460
rect 117520 1400 117600 1420
rect 117720 1460 117800 1480
rect 117720 1420 117740 1460
rect 117780 1420 117800 1460
rect 117720 1400 117800 1420
rect 117920 1460 118000 1480
rect 117920 1420 117940 1460
rect 117980 1420 118000 1460
rect 117920 1400 118000 1420
rect 114980 1120 115120 1140
rect 116950 1350 117090 1370
rect 112440 1060 112520 1080
rect 112440 1020 112460 1060
rect 112500 1020 112520 1060
rect 112440 1000 112520 1020
rect 114970 1060 115050 1080
rect 114970 1020 114990 1060
rect 115030 1020 115050 1060
rect 114970 1000 115050 1020
rect 114830 680 114910 700
rect 114830 640 114850 680
rect 114890 640 114910 680
rect 114830 620 114910 640
rect 113760 190 113840 210
rect 113760 150 113780 190
rect 113820 150 113840 190
rect 113760 130 113840 150
rect 110510 -10 110650 10
rect 113360 70 113500 90
rect 109310 -70 109370 -50
rect 109310 -110 109320 -70
rect 109360 -110 109370 -70
rect 109310 -130 109370 -110
rect 110510 -70 110570 -50
rect 110510 -110 110520 -70
rect 110560 -110 110570 -70
rect 110510 -130 110570 -110
rect 113360 -170 113370 70
rect 113410 -170 113450 70
rect 113490 -170 113500 70
rect 113360 -190 113500 -170
rect 113550 70 113610 90
rect 113550 -170 113560 70
rect 113600 -170 113610 70
rect 113550 -190 113610 -170
rect 113660 70 113720 90
rect 113660 -170 113670 70
rect 113710 -170 113720 70
rect 113660 -190 113720 -170
rect 113770 70 113830 90
rect 113770 -170 113780 70
rect 113820 -170 113830 70
rect 113770 -190 113830 -170
rect 113880 70 113940 90
rect 113880 -170 113890 70
rect 113930 -170 113940 70
rect 113880 -190 113940 -170
rect 113990 70 114050 90
rect 113990 -170 114000 70
rect 114040 -170 114050 70
rect 113990 -190 114050 -170
rect 114100 70 114240 90
rect 114100 -170 114110 70
rect 114150 -170 114190 70
rect 114230 -170 114240 70
rect 116950 10 116960 1350
rect 117000 10 117040 1350
rect 117080 10 117090 1350
rect 116950 -10 117090 10
rect 117230 1350 117290 1370
rect 117230 10 117240 1350
rect 117280 10 117290 1350
rect 117230 -10 117290 10
rect 117430 1350 117490 1370
rect 117430 10 117440 1350
rect 117480 10 117490 1350
rect 117430 -10 117490 10
rect 117630 1350 117690 1370
rect 117630 10 117640 1350
rect 117680 10 117690 1350
rect 117630 -10 117690 10
rect 117830 1350 117890 1370
rect 117830 10 117840 1350
rect 117880 10 117890 1350
rect 117830 -10 117890 10
rect 118030 1350 118090 1370
rect 118030 10 118040 1350
rect 118080 10 118090 1350
rect 118030 -10 118090 10
rect 118230 1350 118370 1370
rect 118230 10 118240 1350
rect 118280 10 118320 1350
rect 118360 10 118370 1350
rect 118760 1350 118830 1370
rect 118760 1300 118770 1350
rect 118820 1300 118830 1350
rect 118760 1280 118830 1300
rect 118880 1350 118950 1370
rect 118880 1300 118890 1350
rect 118940 1300 118950 1350
rect 118880 1280 118950 1300
rect 118230 -10 118370 10
rect 117030 -70 117090 -50
rect 117030 -110 117040 -70
rect 117080 -110 117090 -70
rect 117030 -130 117090 -110
rect 118230 -70 118290 -50
rect 118230 -110 118240 -70
rect 118280 -110 118290 -70
rect 118830 -94 118880 6
rect 118230 -130 118290 -110
rect 114100 -190 114240 -170
rect 113440 -250 113500 -230
rect 113440 -290 113450 -250
rect 113490 -290 113500 -250
rect 113440 -310 113500 -290
rect 114100 -250 114160 -230
rect 114100 -290 114110 -250
rect 114150 -290 114160 -250
rect 114100 -310 114160 -290
rect 113760 -330 113840 -310
rect 113760 -370 113780 -330
rect 113820 -370 113840 -330
rect 113760 -390 113840 -370
rect 113430 -450 113490 -430
rect 113430 -690 113440 -450
rect 113480 -690 113490 -450
rect 113430 -710 113490 -690
rect 114110 -450 114170 -430
rect 114110 -690 114120 -450
rect 114160 -690 114170 -450
rect 114110 -710 114170 -690
<< viali >>
rect 109500 9930 109540 9970
rect 109620 9930 109660 9970
rect 109740 9930 109780 9970
rect 109860 9930 109900 9970
rect 109980 9930 110020 9970
rect 110100 9930 110140 9970
rect 110220 9930 110260 9970
rect 110340 9930 110380 9970
rect 110460 9930 110500 9970
rect 110580 9930 110620 9970
rect 116980 9930 117020 9970
rect 117100 9930 117140 9970
rect 117220 9930 117260 9970
rect 117340 9930 117380 9970
rect 117460 9930 117500 9970
rect 117580 9930 117620 9970
rect 117700 9930 117740 9970
rect 117820 9930 117860 9970
rect 117940 9930 117980 9970
rect 118060 9930 118100 9970
rect 109320 9130 109360 9770
rect 109440 9130 109480 9770
rect 109560 9130 109600 9770
rect 109680 9130 109720 9770
rect 109800 9130 109840 9770
rect 109920 9130 109960 9770
rect 110040 9130 110080 9770
rect 110160 9130 110200 9770
rect 110280 9130 110320 9770
rect 110400 9130 110440 9770
rect 110520 9130 110560 9770
rect 110640 9130 110680 9770
rect 110760 9130 110800 9770
rect 111990 9550 112030 9590
rect 112350 9550 112390 9590
rect 114270 9550 114310 9590
rect 114630 9550 114670 9590
rect 115210 9550 115250 9590
rect 115570 9550 115610 9590
rect 109320 9010 109360 9050
rect 110760 9010 110800 9050
rect 111990 8830 112030 9470
rect 112110 8830 112150 9470
rect 112230 8830 112270 9470
rect 112350 8830 112390 9470
rect 112930 9210 112970 9250
rect 113290 9210 113330 9250
rect 112930 8830 112970 9130
rect 113050 8830 113090 9130
rect 113170 8830 113210 9130
rect 113290 8830 113330 9130
rect 114270 8830 114310 9470
rect 114390 8830 114430 9470
rect 114510 8830 114550 9470
rect 114630 8830 114670 9470
rect 115210 8830 115250 9470
rect 115330 8830 115370 9470
rect 115450 8830 115490 9470
rect 115570 8830 115610 9470
rect 116800 9130 116840 9770
rect 116920 9130 116960 9770
rect 117040 9130 117080 9770
rect 117160 9130 117200 9770
rect 117280 9130 117320 9770
rect 117400 9130 117440 9770
rect 117520 9130 117560 9770
rect 117640 9130 117680 9770
rect 117760 9130 117800 9770
rect 117880 9130 117920 9770
rect 118000 9130 118040 9770
rect 118120 9130 118160 9770
rect 118240 9130 118280 9770
rect 116800 9010 116840 9050
rect 118240 9010 118280 9050
rect 112120 8630 112160 8670
rect 113070 8630 113110 8670
rect 114490 8630 114530 8670
rect 115362 8630 115402 8670
rect 109200 8330 109240 8370
rect 110640 8330 110680 8370
rect 116920 8330 116960 8370
rect 118360 8330 118400 8370
rect 109200 7610 109240 8250
rect 109320 7610 109360 8250
rect 109440 7610 109480 8250
rect 109560 7610 109600 8250
rect 109680 7610 109720 8250
rect 109800 7610 109840 8250
rect 109920 7610 109960 8250
rect 110040 7610 110080 8250
rect 110160 7610 110200 8250
rect 110280 7610 110320 8250
rect 110400 7610 110440 8250
rect 110520 7610 110560 8250
rect 110640 7610 110680 8250
rect 113040 8250 113080 8290
rect 113370 8250 113410 8290
rect 113700 8250 113740 8290
rect 113860 8250 113900 8290
rect 114190 8250 114230 8290
rect 114520 8250 114560 8290
rect 113260 8120 113300 8160
rect 113480 8120 113520 8160
rect 114080 8120 114120 8160
rect 114300 8120 114340 8160
rect 116920 7610 116960 8250
rect 117040 7610 117080 8250
rect 117160 7610 117200 8250
rect 117280 7610 117320 8250
rect 117400 7610 117440 8250
rect 117520 7610 117560 8250
rect 117640 7610 117680 8250
rect 117760 7610 117800 8250
rect 117880 7610 117920 8250
rect 118000 7610 118040 8250
rect 118120 7610 118160 8250
rect 118240 7610 118280 8250
rect 118360 7610 118400 8250
rect 113130 7500 113170 7540
rect 113224 7480 113264 7520
rect 109380 7410 109420 7450
rect 109500 7410 109540 7450
rect 109620 7410 109660 7450
rect 109740 7410 109780 7450
rect 109860 7410 109900 7450
rect 109980 7410 110020 7450
rect 110100 7410 110140 7450
rect 110220 7410 110260 7450
rect 110340 7410 110380 7450
rect 113370 7480 113410 7520
rect 113516 7480 113556 7520
rect 113610 7500 113650 7540
rect 113950 7500 113990 7540
rect 114044 7480 114084 7520
rect 114190 7480 114230 7520
rect 114336 7480 114376 7520
rect 114430 7500 114470 7540
rect 110460 7410 110500 7450
rect 113220 7360 113260 7400
rect 114340 7360 114380 7400
rect 117100 7410 117140 7450
rect 117220 7410 117260 7450
rect 117340 7410 117380 7450
rect 117460 7410 117500 7450
rect 117580 7410 117620 7450
rect 117700 7410 117740 7450
rect 117820 7410 117860 7450
rect 117940 7410 117980 7450
rect 118060 7410 118100 7450
rect 118180 7410 118220 7450
rect 108420 6960 108460 7000
rect 108530 6960 108570 7000
rect 108640 6960 108680 7000
rect 109260 6980 109300 7020
rect 110580 6980 110620 7020
rect 116980 6980 117020 7020
rect 108420 5750 108460 5790
rect 108530 5750 108570 5790
rect 108640 5750 108680 5790
rect 109260 5760 109300 6900
rect 109370 5760 109410 6900
rect 109480 5760 109520 6900
rect 109590 5760 109630 6900
rect 109700 5760 109740 6900
rect 109810 5760 109850 6900
rect 109920 5760 109960 6900
rect 110030 5760 110070 6900
rect 110140 5760 110180 6900
rect 110250 5760 110290 6900
rect 110360 5760 110400 6900
rect 110470 5760 110510 6900
rect 110580 5760 110620 6900
rect 113720 6910 113760 6950
rect 118300 6980 118340 7020
rect 118920 6960 118960 7000
rect 119030 6960 119070 7000
rect 119140 6960 119180 7000
rect 113890 6910 113930 6950
rect 113560 6390 113600 6830
rect 113670 6390 113710 6830
rect 113780 6390 113820 6830
rect 113890 6390 113930 6830
rect 114000 6390 114040 6830
rect 113560 6270 113600 6310
rect 114000 6270 114040 6310
rect 112245 5780 112285 5820
rect 112355 5780 112395 5820
rect 112465 5780 112505 5820
rect 112575 5780 112615 5820
rect 112685 5780 112725 5820
rect 112795 5780 112835 5820
rect 112905 5780 112945 5820
rect 113015 5780 113055 5820
rect 113125 5780 113165 5820
rect 113235 5780 113275 5820
rect 114325 5780 114365 5820
rect 114435 5780 114475 5820
rect 114545 5780 114585 5820
rect 114655 5780 114695 5820
rect 114765 5780 114805 5820
rect 114875 5780 114915 5820
rect 114985 5780 115025 5820
rect 115095 5780 115135 5820
rect 115205 5780 115245 5820
rect 115315 5780 115355 5820
rect 116980 5760 117020 6900
rect 117090 5760 117130 6900
rect 117200 5760 117240 6900
rect 117310 5760 117350 6900
rect 117420 5760 117460 6900
rect 117530 5760 117570 6900
rect 117640 5760 117680 6900
rect 117750 5760 117790 6900
rect 117860 5760 117900 6900
rect 117970 5760 118010 6900
rect 118080 5760 118120 6900
rect 118190 5760 118230 6900
rect 118300 5760 118340 6900
rect 118920 5750 118960 5790
rect 119030 5750 119070 5790
rect 119140 5750 119180 5790
rect 109920 5510 109960 5550
rect 109920 5430 109960 5470
rect 112080 5460 112120 5700
rect 112190 5460 112230 5700
rect 112300 5460 112340 5700
rect 112410 5460 112450 5700
rect 112520 5460 112560 5700
rect 112630 5460 112670 5700
rect 112740 5460 112780 5700
rect 112850 5460 112890 5700
rect 112960 5460 113000 5700
rect 113070 5460 113110 5700
rect 113180 5460 113220 5700
rect 113290 5460 113330 5700
rect 113400 5460 113440 5700
rect 114160 5460 114200 5700
rect 114270 5460 114310 5700
rect 114380 5460 114420 5700
rect 114490 5460 114530 5700
rect 114600 5460 114640 5700
rect 114710 5460 114750 5700
rect 114820 5460 114860 5700
rect 114930 5460 114970 5700
rect 115040 5460 115080 5700
rect 115150 5460 115190 5700
rect 115260 5460 115300 5700
rect 115370 5460 115410 5700
rect 115480 5460 115520 5700
rect 117640 5510 117680 5550
rect 109920 5350 109960 5390
rect 112080 5340 112120 5380
rect 113400 5340 113440 5380
rect 114160 5340 114200 5380
rect 115480 5340 115520 5380
rect 117640 5430 117680 5470
rect 117640 5350 117680 5390
rect 109260 4430 109300 4470
rect 110580 4430 110620 4470
rect 116980 4430 117020 4470
rect 118300 4430 118340 4470
rect 109260 4010 109300 4350
rect 109370 4010 109410 4350
rect 109480 4010 109520 4350
rect 109590 4010 109630 4350
rect 109700 4010 109740 4350
rect 109810 4010 109850 4350
rect 109920 4010 109960 4350
rect 110030 4010 110070 4350
rect 110140 4010 110180 4350
rect 110250 4010 110290 4350
rect 110360 4010 110400 4350
rect 110470 4010 110510 4350
rect 110580 4010 110620 4350
rect 112090 3960 112130 4000
rect 113390 3980 113430 4020
rect 113690 3980 113730 4020
rect 113870 3980 113910 4020
rect 114170 3980 114210 4020
rect 115470 3960 115510 4000
rect 116980 4010 117020 4350
rect 117090 4010 117130 4350
rect 117200 4010 117240 4350
rect 117310 4010 117350 4350
rect 117420 4010 117460 4350
rect 117530 4010 117570 4350
rect 117640 4010 117680 4350
rect 117750 4010 117790 4350
rect 117860 4010 117900 4350
rect 117970 4010 118010 4350
rect 118080 4010 118120 4350
rect 118190 4010 118230 4350
rect 118300 4010 118340 4350
rect 109480 3890 109520 3930
rect 109700 3890 109740 3930
rect 109920 3890 109960 3930
rect 110140 3890 110180 3930
rect 110360 3890 110400 3930
rect 117200 3890 117240 3930
rect 117420 3890 117460 3930
rect 117640 3890 117680 3930
rect 117860 3890 117900 3930
rect 118080 3890 118120 3930
rect 110250 3760 110290 3800
rect 110250 3680 110290 3720
rect 112080 3590 112120 3830
rect 112190 3590 112230 3830
rect 112300 3590 112340 3830
rect 112410 3590 112450 3830
rect 112520 3590 112560 3830
rect 112630 3590 112670 3830
rect 112740 3590 112780 3830
rect 112850 3590 112890 3830
rect 112960 3590 113000 3830
rect 113070 3590 113110 3830
rect 113180 3590 113220 3830
rect 113290 3590 113330 3830
rect 113400 3590 113440 3830
rect 113560 3590 113600 3830
rect 113670 3590 113710 3830
rect 113780 3590 113820 3830
rect 113890 3590 113930 3830
rect 114000 3590 114040 3830
rect 114160 3590 114200 3830
rect 114270 3590 114310 3830
rect 114380 3590 114420 3830
rect 114490 3590 114530 3830
rect 114600 3590 114640 3830
rect 114710 3590 114750 3830
rect 114820 3590 114860 3830
rect 114930 3590 114970 3830
rect 115040 3590 115080 3830
rect 115150 3590 115190 3830
rect 115260 3590 115300 3830
rect 115370 3590 115410 3830
rect 115480 3590 115520 3830
rect 117310 3760 117350 3800
rect 117310 3680 117350 3720
rect 108520 2880 108570 2930
rect 108640 2880 108690 2930
rect 108760 2880 108810 2930
rect 108880 2880 108930 2930
rect 109260 2930 109300 3470
rect 109370 2930 109410 3470
rect 109480 2930 109520 3470
rect 109590 2930 109630 3470
rect 109700 2930 109740 3470
rect 109810 2930 109850 3470
rect 109920 2930 109960 3470
rect 110030 2930 110070 3470
rect 110140 2930 110180 3470
rect 110250 2930 110290 3470
rect 110360 2930 110400 3470
rect 110470 2930 110510 3470
rect 110580 2930 110620 3470
rect 112080 3470 112120 3510
rect 113480 3470 113520 3510
rect 114080 3470 114120 3510
rect 115480 3470 115520 3510
rect 116980 2930 117020 3470
rect 117090 2930 117130 3470
rect 117200 2930 117240 3470
rect 117310 2930 117350 3470
rect 117420 2930 117460 3470
rect 117530 2930 117570 3470
rect 117640 2930 117680 3470
rect 117750 2930 117790 3470
rect 117860 2930 117900 3470
rect 117970 2930 118010 3470
rect 118080 2930 118120 3470
rect 118190 2930 118230 3470
rect 118300 2930 118340 3470
rect 118670 2880 118720 2930
rect 109260 2810 109300 2850
rect 110580 2810 110620 2850
rect 116980 2810 117020 2850
rect 118790 2880 118840 2930
rect 118910 2880 118960 2930
rect 119030 2880 119080 2930
rect 118300 2810 118340 2850
rect 113670 1660 113710 1700
rect 113890 1660 113930 1700
rect 109620 1420 109660 1460
rect 109820 1420 109860 1460
rect 110020 1420 110060 1460
rect 110220 1420 110260 1460
rect 108660 1300 108710 1350
rect 108780 1300 108830 1350
rect 109320 10 109360 1350
rect 109520 10 109560 1350
rect 109720 10 109760 1350
rect 109920 10 109960 1350
rect 110120 10 110160 1350
rect 110320 10 110360 1350
rect 110520 10 110560 1350
rect 112460 1140 112500 1580
rect 112570 1140 112610 1580
rect 112680 1140 112720 1580
rect 112790 1140 112830 1580
rect 112900 1140 112940 1580
rect 113010 1140 113050 1580
rect 113120 1140 113160 1580
rect 113230 1140 113270 1580
rect 113340 1140 113380 1580
rect 113450 1140 113490 1580
rect 113560 1140 113600 1580
rect 113670 1140 113710 1580
rect 113780 1140 113820 1580
rect 113890 1140 113930 1580
rect 114000 1140 114040 1580
rect 114110 1140 114150 1580
rect 114220 1140 114260 1580
rect 114330 1140 114370 1580
rect 114440 1140 114480 1580
rect 114550 1140 114590 1580
rect 114660 1140 114700 1580
rect 114770 1140 114810 1580
rect 114880 1140 114920 1580
rect 114990 1140 115030 1580
rect 117340 1420 117380 1460
rect 117540 1420 117580 1460
rect 117740 1420 117780 1460
rect 117940 1420 117980 1460
rect 112460 1020 112500 1060
rect 114990 1020 115030 1060
rect 114850 640 114890 680
rect 113780 150 113820 190
rect 109320 -110 109360 -70
rect 110520 -110 110560 -70
rect 113450 -170 113490 70
rect 113560 -170 113600 70
rect 113670 -170 113710 70
rect 113780 -170 113820 70
rect 113890 -170 113930 70
rect 114000 -170 114040 70
rect 114110 -170 114150 70
rect 117040 10 117080 1350
rect 117240 10 117280 1350
rect 117440 10 117480 1350
rect 117640 10 117680 1350
rect 117840 10 117880 1350
rect 118040 10 118080 1350
rect 118240 10 118280 1350
rect 118770 1300 118820 1350
rect 118890 1300 118940 1350
rect 117040 -110 117080 -70
rect 118240 -110 118280 -70
rect 113450 -290 113490 -250
rect 114110 -290 114150 -250
rect 113780 -370 113820 -330
rect 113440 -690 113480 -450
rect 114120 -690 114160 -450
<< metal1 >>
rect 104580 9340 104820 12220
rect 104580 9280 104590 9340
rect 104650 9280 104670 9340
rect 104730 9280 104750 9340
rect 104810 9280 104820 9340
rect 104580 9260 104820 9280
rect 104580 9200 104590 9260
rect 104650 9200 104670 9260
rect 104730 9200 104750 9260
rect 104810 9200 104820 9260
rect 104580 9180 104820 9200
rect 104580 9120 104590 9180
rect 104650 9120 104670 9180
rect 104730 9120 104750 9180
rect 104810 9120 104820 9180
rect 104580 9110 104820 9120
rect 105280 9340 105520 12220
rect 105280 9280 105290 9340
rect 105350 9280 105370 9340
rect 105430 9280 105450 9340
rect 105510 9280 105520 9340
rect 105280 9260 105520 9280
rect 105280 9200 105290 9260
rect 105350 9200 105370 9260
rect 105430 9200 105450 9260
rect 105510 9200 105520 9260
rect 105280 9180 105520 9200
rect 105280 9120 105290 9180
rect 105350 9120 105370 9180
rect 105430 9120 105450 9180
rect 105510 9120 105520 9180
rect 105280 9110 105520 9120
rect 105980 9340 106220 12220
rect 105980 9280 105990 9340
rect 106050 9280 106070 9340
rect 106130 9280 106150 9340
rect 106210 9280 106220 9340
rect 105980 9260 106220 9280
rect 105980 9200 105990 9260
rect 106050 9200 106070 9260
rect 106130 9200 106150 9260
rect 106210 9200 106220 9260
rect 105980 9180 106220 9200
rect 105980 9120 105990 9180
rect 106050 9120 106070 9180
rect 106130 9120 106150 9180
rect 106210 9120 106220 9180
rect 105980 9110 106220 9120
rect 106680 9340 106920 12220
rect 106680 9280 106690 9340
rect 106750 9280 106770 9340
rect 106830 9280 106850 9340
rect 106910 9280 106920 9340
rect 106680 9260 106920 9280
rect 106680 9200 106690 9260
rect 106750 9200 106770 9260
rect 106830 9200 106850 9260
rect 106910 9200 106920 9260
rect 106680 9180 106920 9200
rect 106680 9120 106690 9180
rect 106750 9120 106770 9180
rect 106830 9120 106850 9180
rect 106910 9120 106920 9180
rect 106680 9110 106920 9120
rect 108080 9340 108320 12220
rect 109490 9980 109550 9990
rect 109490 9910 109550 9920
rect 109610 9980 109670 9990
rect 109610 9910 109670 9920
rect 109730 9980 109790 9990
rect 109730 9910 109790 9920
rect 109850 9980 109910 9990
rect 109850 9910 109910 9920
rect 109970 9980 110150 9990
rect 110030 9920 110090 9980
rect 109970 9910 110150 9920
rect 110210 9980 110270 9990
rect 110210 9910 110270 9920
rect 110330 9980 110390 9990
rect 110330 9910 110390 9920
rect 110450 9980 110510 9990
rect 110450 9910 110510 9920
rect 110570 9980 110630 9990
rect 110570 9910 110630 9920
rect 114900 9980 114980 9990
rect 114900 9920 114910 9980
rect 114970 9920 114980 9980
rect 109420 9870 109500 9880
rect 109420 9810 109430 9870
rect 109490 9810 109500 9870
rect 109420 9800 109500 9810
rect 109660 9870 109740 9880
rect 109660 9810 109670 9870
rect 109730 9810 109740 9870
rect 109660 9800 109740 9810
rect 109900 9870 109980 9880
rect 109900 9810 109910 9870
rect 109970 9810 109980 9870
rect 109900 9800 109980 9810
rect 110140 9870 110220 9880
rect 110140 9810 110150 9870
rect 110210 9810 110220 9870
rect 110140 9800 110220 9810
rect 110380 9870 110460 9880
rect 110380 9810 110390 9870
rect 110450 9810 110460 9870
rect 110380 9800 110460 9810
rect 110620 9870 110700 9880
rect 110620 9810 110630 9870
rect 110690 9810 110700 9870
rect 110620 9800 110700 9810
rect 112210 9870 112290 9880
rect 112210 9810 112220 9870
rect 112280 9810 112290 9870
rect 108080 9280 108090 9340
rect 108150 9280 108170 9340
rect 108230 9280 108250 9340
rect 108310 9280 108320 9340
rect 108080 9260 108320 9280
rect 108080 9200 108090 9260
rect 108150 9200 108170 9260
rect 108230 9200 108250 9260
rect 108310 9200 108320 9260
rect 108080 9180 108320 9200
rect 108080 9120 108090 9180
rect 108150 9120 108170 9180
rect 108230 9120 108250 9180
rect 108310 9120 108320 9180
rect 108080 7350 108320 9120
rect 109310 9770 109370 9790
rect 109310 9130 109320 9770
rect 109360 9130 109370 9770
rect 109310 9070 109370 9130
rect 109430 9770 109490 9800
rect 109430 9130 109440 9770
rect 109480 9130 109490 9770
rect 109300 9060 109380 9070
rect 109300 9000 109310 9060
rect 109370 9000 109380 9060
rect 109300 8990 109380 9000
rect 109430 8960 109490 9130
rect 109550 9770 109610 9790
rect 109550 9130 109560 9770
rect 109600 9130 109610 9770
rect 109550 9070 109610 9130
rect 109670 9770 109730 9800
rect 109670 9130 109680 9770
rect 109720 9130 109730 9770
rect 109540 9060 109620 9070
rect 109540 9000 109550 9060
rect 109610 9000 109620 9060
rect 109540 8990 109620 9000
rect 109670 8960 109730 9130
rect 109790 9770 109850 9790
rect 109790 9130 109800 9770
rect 109840 9130 109850 9770
rect 109790 9070 109850 9130
rect 109910 9770 109970 9800
rect 109910 9130 109920 9770
rect 109960 9130 109970 9770
rect 109780 9060 109860 9070
rect 109780 9000 109790 9060
rect 109850 9000 109860 9060
rect 109780 8990 109860 9000
rect 109910 8960 109970 9130
rect 110030 9770 110090 9790
rect 110030 9130 110040 9770
rect 110080 9130 110090 9770
rect 110030 9070 110090 9130
rect 110150 9770 110210 9800
rect 110150 9130 110160 9770
rect 110200 9130 110210 9770
rect 110020 9060 110100 9070
rect 110020 9000 110030 9060
rect 110090 9000 110100 9060
rect 110020 8990 110100 9000
rect 110150 8960 110210 9130
rect 110270 9770 110330 9790
rect 110270 9130 110280 9770
rect 110320 9130 110330 9770
rect 110270 9070 110330 9130
rect 110390 9770 110450 9800
rect 110390 9130 110400 9770
rect 110440 9130 110450 9770
rect 110260 9060 110340 9070
rect 110260 9000 110270 9060
rect 110330 9000 110340 9060
rect 110260 8990 110340 9000
rect 110390 8960 110450 9130
rect 110510 9770 110570 9790
rect 110510 9130 110520 9770
rect 110560 9130 110570 9770
rect 110510 9070 110570 9130
rect 110630 9770 110690 9800
rect 110630 9130 110640 9770
rect 110680 9130 110690 9770
rect 110500 9060 110580 9070
rect 110500 9000 110510 9060
rect 110570 9000 110580 9060
rect 110500 8990 110580 9000
rect 110630 8960 110690 9130
rect 110750 9770 110810 9790
rect 110750 9130 110760 9770
rect 110800 9130 110810 9770
rect 111970 9600 112050 9610
rect 111970 9540 111980 9600
rect 112040 9540 112050 9600
rect 111970 9530 112050 9540
rect 112210 9600 112290 9810
rect 113150 9870 113230 9880
rect 113150 9810 113160 9870
rect 113220 9810 113230 9870
rect 113150 9800 113230 9810
rect 114370 9870 114450 9880
rect 114370 9810 114380 9870
rect 114440 9810 114450 9870
rect 114370 9800 114450 9810
rect 112210 9540 112220 9600
rect 112280 9540 112290 9600
rect 112210 9530 112290 9540
rect 112330 9600 112410 9610
rect 112330 9540 112340 9600
rect 112400 9540 112410 9600
rect 112330 9530 112410 9540
rect 110750 9070 110810 9130
rect 111980 9470 112040 9530
rect 110740 9060 110820 9070
rect 110740 9000 110750 9060
rect 110810 9000 110820 9060
rect 110740 8990 110820 9000
rect 111070 9060 111310 9070
rect 111070 9000 111080 9060
rect 111140 9000 111160 9060
rect 111220 9000 111240 9060
rect 111300 9000 111310 9060
rect 109180 8950 110700 8960
rect 109180 8890 109190 8950
rect 109250 8890 109430 8950
rect 109490 8890 109670 8950
rect 109730 8890 109910 8950
rect 109970 8890 110150 8950
rect 110210 8890 110390 8950
rect 110450 8890 110630 8950
rect 110690 8890 110700 8950
rect 109180 8870 110700 8890
rect 109180 8810 109190 8870
rect 109250 8810 109430 8870
rect 109490 8810 109670 8870
rect 109730 8810 109910 8870
rect 109970 8810 110150 8870
rect 110210 8810 110390 8870
rect 110450 8810 110630 8870
rect 110690 8810 110700 8870
rect 109180 8790 110700 8810
rect 109180 8730 109190 8790
rect 109250 8730 109430 8790
rect 109490 8730 109670 8790
rect 109730 8730 109910 8790
rect 109970 8730 110150 8790
rect 110210 8730 110390 8790
rect 110450 8730 110630 8790
rect 110690 8730 110700 8790
rect 109180 8710 110700 8730
rect 109180 8650 109190 8710
rect 109250 8650 109430 8710
rect 109490 8650 109670 8710
rect 109730 8650 109910 8710
rect 109970 8650 110150 8710
rect 110210 8650 110390 8710
rect 110450 8650 110630 8710
rect 110690 8650 110700 8710
rect 109180 8630 110700 8650
rect 109180 8570 109190 8630
rect 109250 8570 109430 8630
rect 109490 8570 109670 8630
rect 109730 8570 109910 8630
rect 109970 8570 110150 8630
rect 110210 8570 110390 8630
rect 110450 8570 110630 8630
rect 110690 8570 110700 8630
rect 109180 8550 110700 8570
rect 109180 8490 109190 8550
rect 109250 8490 109430 8550
rect 109490 8490 109670 8550
rect 109730 8490 109910 8550
rect 109970 8490 110150 8550
rect 110210 8490 110390 8550
rect 110450 8490 110630 8550
rect 110690 8490 110700 8550
rect 109180 8470 110700 8490
rect 109180 8410 109190 8470
rect 109250 8410 109430 8470
rect 109490 8410 109670 8470
rect 109730 8410 109910 8470
rect 109970 8410 110150 8470
rect 110210 8410 110390 8470
rect 110450 8410 110630 8470
rect 110690 8410 110700 8470
rect 109180 8400 110700 8410
rect 111070 8460 111310 9000
rect 111980 8830 111990 9470
rect 112030 8830 112040 9470
rect 111980 8810 112040 8830
rect 112100 9470 112160 9490
rect 112100 8830 112110 9470
rect 112150 8830 112160 9470
rect 112100 8690 112160 8830
rect 112220 9470 112280 9530
rect 112220 8830 112230 9470
rect 112270 8830 112280 9470
rect 112220 8800 112280 8830
rect 112340 9470 112400 9530
rect 112340 8830 112350 9470
rect 112390 8830 112400 9470
rect 112910 9420 112990 9430
rect 112910 9360 112920 9420
rect 112980 9360 112990 9420
rect 112910 9340 112990 9360
rect 112910 9280 112920 9340
rect 112980 9280 112990 9340
rect 112910 9260 112990 9280
rect 112910 9200 112920 9260
rect 112980 9200 112990 9260
rect 112910 9190 112990 9200
rect 113030 9420 113110 9430
rect 113030 9360 113040 9420
rect 113100 9360 113110 9420
rect 113030 9340 113110 9360
rect 113030 9280 113040 9340
rect 113100 9280 113110 9340
rect 113030 9260 113110 9280
rect 113030 9200 113040 9260
rect 113100 9200 113110 9260
rect 113030 9190 113110 9200
rect 112340 8810 112400 8830
rect 112920 9130 112980 9190
rect 112920 8830 112930 9130
rect 112970 8830 112980 9130
rect 112920 8810 112980 8830
rect 113040 9130 113100 9190
rect 113040 8830 113050 9130
rect 113090 8830 113100 9130
rect 113040 8810 113100 8830
rect 113160 9130 113220 9800
rect 113680 9760 113920 9770
rect 113680 9700 113690 9760
rect 113750 9700 113770 9760
rect 113830 9700 113850 9760
rect 113910 9700 113920 9760
rect 113680 9680 113920 9700
rect 113680 9620 113690 9680
rect 113750 9620 113770 9680
rect 113830 9620 113850 9680
rect 113910 9620 113920 9680
rect 113680 9600 113920 9620
rect 113680 9540 113690 9600
rect 113750 9540 113770 9600
rect 113830 9540 113850 9600
rect 113910 9540 113920 9600
rect 113270 9420 113350 9430
rect 113270 9360 113280 9420
rect 113340 9360 113350 9420
rect 113270 9340 113350 9360
rect 113270 9280 113280 9340
rect 113340 9280 113350 9340
rect 113270 9260 113350 9280
rect 113270 9200 113280 9260
rect 113340 9200 113350 9260
rect 113270 9190 113350 9200
rect 113680 9420 113920 9540
rect 114250 9760 114330 9770
rect 114250 9700 114260 9760
rect 114320 9700 114330 9760
rect 114250 9680 114330 9700
rect 114250 9620 114260 9680
rect 114320 9620 114330 9680
rect 114250 9600 114330 9620
rect 114250 9540 114260 9600
rect 114320 9540 114330 9600
rect 114250 9530 114330 9540
rect 113680 9360 113690 9420
rect 113750 9360 113770 9420
rect 113830 9360 113850 9420
rect 113910 9360 113920 9420
rect 113680 9340 113920 9360
rect 113680 9280 113690 9340
rect 113750 9280 113770 9340
rect 113830 9280 113850 9340
rect 113910 9280 113920 9340
rect 113680 9260 113920 9280
rect 113680 9200 113690 9260
rect 113750 9200 113770 9260
rect 113830 9200 113850 9260
rect 113910 9200 113920 9260
rect 113160 8830 113170 9130
rect 113210 8830 113220 9130
rect 113160 8800 113220 8830
rect 113280 9130 113340 9190
rect 113280 8830 113290 9130
rect 113330 8830 113340 9130
rect 113280 8810 113340 8830
rect 112210 8790 112290 8800
rect 112210 8730 112220 8790
rect 112280 8730 112290 8790
rect 112210 8720 112290 8730
rect 113150 8790 113230 8800
rect 113150 8730 113160 8790
rect 113220 8730 113230 8790
rect 113150 8720 113230 8730
rect 111340 8680 111420 8690
rect 111340 8620 111350 8680
rect 111410 8620 111420 8680
rect 111340 8610 111420 8620
rect 112100 8680 112180 8690
rect 112100 8620 112110 8680
rect 112170 8620 112180 8680
rect 112100 8610 112180 8620
rect 113060 8680 113120 8690
rect 113060 8610 113120 8620
rect 111070 8400 111080 8460
rect 111140 8400 111160 8460
rect 111220 8400 111240 8460
rect 111300 8400 111310 8460
rect 109190 8370 109250 8400
rect 109190 8330 109200 8370
rect 109240 8330 109250 8370
rect 109190 8250 109250 8330
rect 109300 8350 109380 8360
rect 109300 8290 109310 8350
rect 109370 8290 109380 8350
rect 109300 8280 109380 8290
rect 108080 7290 108090 7350
rect 108150 7290 108170 7350
rect 108230 7290 108250 7350
rect 108310 7290 108320 7350
rect 108080 7270 108320 7290
rect 108080 7210 108090 7270
rect 108150 7210 108170 7270
rect 108230 7210 108250 7270
rect 108310 7210 108320 7270
rect 108080 7190 108320 7210
rect 108080 7130 108090 7190
rect 108150 7130 108170 7190
rect 108230 7130 108250 7190
rect 108310 7130 108320 7190
rect 108080 7120 108320 7130
rect 108510 7670 108590 7680
rect 108510 7610 108520 7670
rect 108580 7610 108590 7670
rect 108510 7020 108590 7610
rect 109190 7610 109200 8250
rect 109240 7610 109250 8250
rect 109190 7590 109250 7610
rect 109310 8250 109370 8280
rect 109310 7610 109320 8250
rect 109360 7610 109370 8250
rect 109310 7580 109370 7610
rect 109430 8250 109490 8400
rect 109540 8350 109620 8360
rect 109540 8290 109550 8350
rect 109610 8290 109620 8350
rect 109540 8280 109620 8290
rect 109430 7610 109440 8250
rect 109480 7610 109490 8250
rect 109430 7590 109490 7610
rect 109550 8250 109610 8280
rect 109550 7610 109560 8250
rect 109600 7610 109610 8250
rect 109550 7580 109610 7610
rect 109670 8250 109730 8400
rect 109780 8350 109860 8360
rect 109780 8290 109790 8350
rect 109850 8290 109860 8350
rect 109780 8280 109860 8290
rect 109670 7610 109680 8250
rect 109720 7610 109730 8250
rect 109670 7590 109730 7610
rect 109790 8250 109850 8280
rect 109790 7610 109800 8250
rect 109840 7610 109850 8250
rect 109790 7580 109850 7610
rect 109910 8250 109970 8400
rect 110020 8350 110100 8360
rect 110020 8290 110030 8350
rect 110090 8290 110100 8350
rect 110020 8280 110100 8290
rect 109910 7610 109920 8250
rect 109960 7610 109970 8250
rect 109910 7590 109970 7610
rect 110030 8250 110090 8280
rect 110030 7610 110040 8250
rect 110080 7610 110090 8250
rect 110030 7580 110090 7610
rect 110150 8250 110210 8400
rect 110260 8350 110340 8360
rect 110260 8290 110270 8350
rect 110330 8290 110340 8350
rect 110260 8280 110340 8290
rect 110150 7610 110160 8250
rect 110200 7610 110210 8250
rect 110150 7590 110210 7610
rect 110270 8250 110330 8280
rect 110270 7610 110280 8250
rect 110320 7610 110330 8250
rect 110270 7580 110330 7610
rect 110390 8250 110450 8400
rect 110630 8370 110690 8400
rect 110500 8350 110580 8360
rect 110500 8290 110510 8350
rect 110570 8290 110580 8350
rect 110500 8280 110580 8290
rect 110630 8330 110640 8370
rect 110680 8330 110690 8370
rect 110390 7610 110400 8250
rect 110440 7610 110450 8250
rect 110390 7590 110450 7610
rect 110510 8250 110570 8280
rect 110510 7610 110520 8250
rect 110560 7610 110570 8250
rect 110510 7580 110570 7610
rect 110630 8250 110690 8330
rect 110630 7610 110640 8250
rect 110680 7610 110690 8250
rect 110630 7590 110690 7610
rect 111070 8380 111310 8400
rect 111070 8320 111080 8380
rect 111140 8320 111160 8380
rect 111220 8320 111240 8380
rect 111300 8320 111310 8380
rect 111070 8300 111310 8320
rect 111070 8240 111080 8300
rect 111140 8240 111160 8300
rect 111220 8240 111240 8300
rect 111300 8240 111310 8300
rect 109300 7570 109380 7580
rect 109300 7510 109310 7570
rect 109370 7510 109380 7570
rect 109300 7500 109380 7510
rect 109540 7570 109620 7580
rect 109540 7510 109550 7570
rect 109610 7510 109620 7570
rect 109540 7500 109620 7510
rect 109780 7570 109860 7580
rect 109780 7510 109790 7570
rect 109850 7510 109860 7570
rect 109780 7500 109860 7510
rect 110020 7570 110100 7580
rect 110020 7510 110030 7570
rect 110090 7510 110100 7570
rect 110020 7500 110100 7510
rect 110260 7570 110340 7580
rect 110260 7510 110270 7570
rect 110330 7510 110340 7570
rect 110260 7500 110340 7510
rect 110500 7570 110580 7580
rect 110500 7510 110510 7570
rect 110570 7510 110580 7570
rect 110500 7500 110580 7510
rect 110800 7570 111040 7580
rect 110800 7510 110810 7570
rect 110870 7510 110890 7570
rect 110950 7510 110970 7570
rect 111030 7510 111040 7570
rect 109370 7460 109430 7470
rect 109370 7390 109430 7400
rect 109490 7460 109550 7470
rect 109490 7390 109550 7400
rect 109610 7460 109670 7470
rect 109610 7390 109670 7400
rect 109730 7460 109790 7470
rect 109730 7390 109790 7400
rect 109850 7460 109910 7470
rect 109850 7390 109910 7400
rect 109970 7460 110030 7470
rect 109970 7390 110030 7400
rect 110090 7460 110150 7470
rect 110090 7390 110150 7400
rect 110210 7460 110270 7470
rect 110210 7390 110270 7400
rect 110330 7460 110390 7470
rect 110330 7390 110390 7400
rect 110450 7460 110510 7470
rect 110450 7390 110510 7400
rect 109240 7350 109320 7360
rect 109240 7290 109250 7350
rect 109310 7290 109320 7350
rect 109240 7270 109320 7290
rect 109240 7210 109250 7270
rect 109310 7210 109320 7270
rect 109240 7190 109320 7210
rect 109240 7130 109250 7190
rect 109310 7130 109320 7190
rect 109240 7120 109320 7130
rect 109460 7350 109540 7360
rect 109460 7290 109470 7350
rect 109530 7290 109540 7350
rect 109460 7270 109540 7290
rect 109460 7210 109470 7270
rect 109530 7210 109540 7270
rect 109460 7190 109540 7210
rect 109460 7130 109470 7190
rect 109530 7130 109540 7190
rect 109460 7120 109540 7130
rect 109680 7350 109760 7360
rect 109680 7290 109690 7350
rect 109750 7290 109760 7350
rect 109680 7270 109760 7290
rect 109680 7210 109690 7270
rect 109750 7210 109760 7270
rect 109680 7190 109760 7210
rect 109680 7130 109690 7190
rect 109750 7130 109760 7190
rect 109680 7120 109760 7130
rect 109900 7350 109980 7360
rect 109900 7290 109910 7350
rect 109970 7290 109980 7350
rect 109900 7270 109980 7290
rect 109900 7210 109910 7270
rect 109970 7210 109980 7270
rect 109900 7190 109980 7210
rect 109900 7130 109910 7190
rect 109970 7130 109980 7190
rect 109900 7120 109980 7130
rect 110120 7350 110200 7360
rect 110120 7290 110130 7350
rect 110190 7290 110200 7350
rect 110120 7270 110200 7290
rect 110120 7210 110130 7270
rect 110190 7210 110200 7270
rect 110120 7190 110200 7210
rect 110120 7130 110130 7190
rect 110190 7130 110200 7190
rect 110120 7120 110200 7130
rect 110340 7350 110420 7360
rect 110340 7290 110350 7350
rect 110410 7290 110420 7350
rect 110340 7270 110420 7290
rect 110340 7210 110350 7270
rect 110410 7210 110420 7270
rect 110340 7190 110420 7210
rect 110340 7130 110350 7190
rect 110410 7130 110420 7190
rect 110340 7120 110420 7130
rect 110560 7350 110640 7360
rect 110560 7290 110570 7350
rect 110630 7290 110640 7350
rect 110560 7270 110640 7290
rect 110560 7210 110570 7270
rect 110630 7210 110640 7270
rect 110560 7190 110640 7210
rect 110560 7130 110570 7190
rect 110630 7130 110640 7190
rect 110560 7120 110640 7130
rect 109250 7020 109310 7120
rect 108408 7000 108690 7020
rect 108408 6960 108420 7000
rect 108460 6960 108530 7000
rect 108570 6960 108640 7000
rect 108680 6960 108690 7000
rect 108408 6940 108690 6960
rect 109250 6980 109260 7020
rect 109300 6980 109310 7020
rect 109250 6900 109310 6980
rect 109350 7000 109430 7010
rect 109350 6940 109360 7000
rect 109420 6940 109430 7000
rect 109350 6930 109430 6940
rect 108408 5790 108690 5810
rect 108408 5750 108420 5790
rect 108460 5750 108530 5790
rect 108570 5750 108640 5790
rect 108680 5750 108690 5790
rect 108408 5730 108690 5750
rect 109250 5760 109260 6900
rect 109300 5760 109310 6900
rect 109250 5740 109310 5760
rect 109360 6900 109420 6930
rect 109360 5760 109370 6900
rect 109410 5760 109420 6900
rect 109360 5730 109420 5760
rect 109470 6900 109530 7120
rect 109570 7000 109650 7010
rect 109570 6940 109580 7000
rect 109640 6940 109650 7000
rect 109570 6930 109650 6940
rect 109470 5760 109480 6900
rect 109520 5760 109530 6900
rect 109470 5740 109530 5760
rect 109580 6900 109640 6930
rect 109580 5760 109590 6900
rect 109630 5760 109640 6900
rect 109580 5730 109640 5760
rect 109690 6900 109750 7120
rect 109790 7000 109870 7010
rect 109790 6940 109800 7000
rect 109860 6940 109870 7000
rect 109790 6930 109870 6940
rect 109690 5760 109700 6900
rect 109740 5760 109750 6900
rect 109690 5740 109750 5760
rect 109800 6900 109860 6930
rect 109800 5760 109810 6900
rect 109850 5760 109860 6900
rect 109800 5730 109860 5760
rect 109910 6900 109970 7120
rect 110010 7000 110090 7010
rect 110010 6940 110020 7000
rect 110080 6940 110090 7000
rect 110010 6930 110090 6940
rect 109910 5760 109920 6900
rect 109960 5760 109970 6900
rect 109910 5740 109970 5760
rect 110020 6900 110080 6930
rect 110020 5760 110030 6900
rect 110070 5760 110080 6900
rect 110020 5730 110080 5760
rect 110130 6900 110190 7120
rect 110230 7000 110310 7010
rect 110230 6940 110240 7000
rect 110300 6940 110310 7000
rect 110230 6930 110310 6940
rect 110130 5760 110140 6900
rect 110180 5760 110190 6900
rect 110130 5740 110190 5760
rect 110240 6900 110300 6930
rect 110240 5760 110250 6900
rect 110290 5760 110300 6900
rect 110240 5730 110300 5760
rect 110350 6900 110410 7120
rect 110570 7020 110630 7120
rect 110450 7000 110530 7010
rect 110450 6940 110460 7000
rect 110520 6940 110530 7000
rect 110450 6930 110530 6940
rect 110570 6980 110580 7020
rect 110620 6980 110630 7020
rect 110350 5760 110360 6900
rect 110400 5760 110410 6900
rect 110350 5740 110410 5760
rect 110460 6900 110520 6930
rect 110460 5760 110470 6900
rect 110510 5760 110520 6900
rect 110460 5730 110520 5760
rect 110570 6900 110630 6980
rect 110570 5760 110580 6900
rect 110620 5760 110630 6900
rect 110570 5740 110630 5760
rect 110800 6960 111040 7510
rect 110800 6900 110810 6960
rect 110870 6900 110890 6960
rect 110950 6900 110970 6960
rect 111030 6900 111040 6960
rect 110800 6880 111040 6900
rect 110800 6820 110810 6880
rect 110870 6820 110890 6880
rect 110950 6820 110970 6880
rect 111030 6820 111040 6880
rect 110800 6800 111040 6820
rect 110800 6740 110810 6800
rect 110870 6740 110890 6800
rect 110950 6740 110970 6800
rect 111030 6740 111040 6800
rect 108430 5560 108670 5730
rect 108430 5500 108440 5560
rect 108500 5500 108520 5560
rect 108580 5500 108600 5560
rect 108660 5500 108670 5560
rect 108430 5480 108670 5500
rect 108430 5420 108440 5480
rect 108500 5420 108520 5480
rect 108580 5420 108600 5480
rect 108660 5420 108670 5480
rect 108430 5400 108670 5420
rect 108430 5340 108440 5400
rect 108500 5340 108520 5400
rect 108580 5340 108600 5400
rect 108660 5340 108670 5400
rect 108430 5330 108670 5340
rect 109350 5720 109430 5730
rect 109350 5660 109360 5720
rect 109420 5660 109430 5720
rect 109350 5270 109430 5660
rect 109570 5720 109650 5730
rect 109570 5660 109580 5720
rect 109640 5660 109650 5720
rect 109570 5270 109650 5660
rect 109790 5720 109870 5730
rect 109790 5660 109800 5720
rect 109860 5660 109870 5720
rect 109790 5270 109870 5660
rect 110010 5720 110090 5730
rect 110010 5660 110020 5720
rect 110080 5660 110090 5720
rect 109900 5560 109980 5570
rect 109900 5500 109910 5560
rect 109970 5500 109980 5560
rect 109900 5480 109980 5500
rect 109900 5420 109910 5480
rect 109970 5420 109980 5480
rect 109900 5400 109980 5420
rect 109900 5340 109910 5400
rect 109970 5340 109980 5400
rect 109900 5330 109980 5340
rect 110010 5270 110090 5660
rect 110230 5720 110310 5730
rect 110230 5660 110240 5720
rect 110300 5660 110310 5720
rect 110230 5270 110310 5660
rect 110450 5720 110530 5730
rect 110450 5660 110460 5720
rect 110520 5660 110530 5720
rect 110450 5270 110530 5660
rect 107980 5260 108480 5270
rect 107980 5200 107990 5260
rect 108050 5200 108070 5260
rect 108130 5200 108160 5260
rect 108220 5200 108240 5260
rect 108300 5200 108330 5260
rect 108390 5200 108410 5260
rect 108470 5200 108480 5260
rect 107980 5180 108480 5200
rect 107980 5120 107990 5180
rect 108050 5120 108070 5180
rect 108130 5120 108160 5180
rect 108220 5120 108240 5180
rect 108300 5120 108330 5180
rect 108390 5120 108410 5180
rect 108470 5120 108480 5180
rect 107980 5100 108480 5120
rect 107980 5040 107990 5100
rect 108050 5040 108070 5100
rect 108130 5040 108160 5100
rect 108220 5040 108240 5100
rect 108300 5040 108330 5100
rect 108390 5040 108410 5100
rect 108470 5040 108480 5100
rect 107680 4720 107920 4730
rect 107680 4660 107690 4720
rect 107750 4660 107770 4720
rect 107830 4660 107850 4720
rect 107910 4660 107920 4720
rect 107680 4640 107920 4660
rect 107680 4580 107690 4640
rect 107750 4580 107770 4640
rect 107830 4580 107850 4640
rect 107910 4580 107920 4640
rect 107680 4560 107920 4580
rect 107680 4500 107690 4560
rect 107750 4500 107770 4560
rect 107830 4500 107850 4560
rect 107910 4500 107920 4560
rect 107680 2500 107920 4500
rect 107680 2440 107690 2500
rect 107750 2440 107770 2500
rect 107830 2440 107850 2500
rect 107910 2440 107920 2500
rect 107680 2420 107920 2440
rect 107680 2360 107690 2420
rect 107750 2360 107770 2420
rect 107830 2360 107850 2420
rect 107910 2360 107920 2420
rect 107680 2340 107920 2360
rect 107680 2280 107690 2340
rect 107750 2280 107770 2340
rect 107830 2280 107850 2340
rect 107910 2280 107920 2340
rect 104580 -1160 104820 -1150
rect 104580 -1220 104590 -1160
rect 104650 -1220 104670 -1160
rect 104730 -1220 104750 -1160
rect 104810 -1220 104820 -1160
rect 104580 -1240 104820 -1220
rect 104580 -1300 104590 -1240
rect 104650 -1300 104670 -1240
rect 104730 -1300 104750 -1240
rect 104810 -1300 104820 -1240
rect 104580 -1320 104820 -1300
rect 104580 -1380 104590 -1320
rect 104650 -1380 104670 -1320
rect 104730 -1380 104750 -1320
rect 104810 -1380 104820 -1320
rect 104580 -3000 104820 -1380
rect 105280 -1160 105520 -1150
rect 105280 -1220 105290 -1160
rect 105350 -1220 105370 -1160
rect 105430 -1220 105450 -1160
rect 105510 -1220 105520 -1160
rect 105280 -1240 105520 -1220
rect 105280 -1300 105290 -1240
rect 105350 -1300 105370 -1240
rect 105430 -1300 105450 -1240
rect 105510 -1300 105520 -1240
rect 105280 -1320 105520 -1300
rect 105280 -1380 105290 -1320
rect 105350 -1380 105370 -1320
rect 105430 -1380 105450 -1320
rect 105510 -1380 105520 -1320
rect 105280 -3000 105520 -1380
rect 105980 -1160 106220 -1150
rect 105980 -1220 105990 -1160
rect 106050 -1220 106070 -1160
rect 106130 -1220 106150 -1160
rect 106210 -1220 106220 -1160
rect 105980 -1240 106220 -1220
rect 105980 -1300 105990 -1240
rect 106050 -1300 106070 -1240
rect 106130 -1300 106150 -1240
rect 106210 -1300 106220 -1240
rect 105980 -1320 106220 -1300
rect 105980 -1380 105990 -1320
rect 106050 -1380 106070 -1320
rect 106130 -1380 106150 -1320
rect 106210 -1380 106220 -1320
rect 105980 -3000 106220 -1380
rect 106680 -1160 106920 -1150
rect 106680 -1220 106690 -1160
rect 106750 -1220 106770 -1160
rect 106830 -1220 106850 -1160
rect 106910 -1220 106920 -1160
rect 106680 -1240 106920 -1220
rect 106680 -1300 106690 -1240
rect 106750 -1300 106770 -1240
rect 106830 -1300 106850 -1240
rect 106910 -1300 106920 -1240
rect 106680 -1320 106920 -1300
rect 106680 -1380 106690 -1320
rect 106750 -1380 106770 -1320
rect 106830 -1380 106850 -1320
rect 106910 -1380 106920 -1320
rect 106680 -3000 106920 -1380
rect 107380 -1160 107620 -1150
rect 107380 -1220 107390 -1160
rect 107450 -1220 107470 -1160
rect 107530 -1220 107550 -1160
rect 107610 -1220 107620 -1160
rect 107380 -1240 107620 -1220
rect 107380 -1300 107390 -1240
rect 107450 -1300 107470 -1240
rect 107530 -1300 107550 -1240
rect 107610 -1300 107620 -1240
rect 107380 -1320 107620 -1300
rect 107380 -1380 107390 -1320
rect 107450 -1380 107470 -1320
rect 107530 -1380 107550 -1320
rect 107610 -1380 107620 -1320
rect 107380 -3000 107620 -1380
rect 107680 -1160 107920 2280
rect 107980 4120 108480 5040
rect 109350 5260 110530 5270
rect 109350 5200 109360 5260
rect 109420 5200 109470 5260
rect 109530 5200 109580 5260
rect 109640 5200 109690 5260
rect 109750 5200 109800 5260
rect 109860 5200 109910 5260
rect 109970 5200 110020 5260
rect 110080 5200 110130 5260
rect 110190 5200 110240 5260
rect 110300 5200 110350 5260
rect 110410 5200 110460 5260
rect 110520 5200 110530 5260
rect 109350 5180 110530 5200
rect 109350 5120 109360 5180
rect 109420 5120 109470 5180
rect 109530 5120 109580 5180
rect 109640 5120 109690 5180
rect 109750 5120 109800 5180
rect 109860 5120 109910 5180
rect 109970 5120 110020 5180
rect 110080 5120 110130 5180
rect 110190 5120 110240 5180
rect 110300 5120 110350 5180
rect 110410 5120 110460 5180
rect 110520 5120 110530 5180
rect 109350 5100 110530 5120
rect 109350 5040 109360 5100
rect 109420 5040 109470 5100
rect 109530 5040 109580 5100
rect 109640 5040 109690 5100
rect 109750 5040 109800 5100
rect 109860 5040 109910 5100
rect 109970 5040 110020 5100
rect 110080 5040 110130 5100
rect 110190 5040 110240 5100
rect 110300 5040 110350 5100
rect 110410 5040 110460 5100
rect 110520 5040 110530 5100
rect 109350 5030 110530 5040
rect 110800 5560 111040 6740
rect 110800 5500 110810 5560
rect 110870 5500 110890 5560
rect 110950 5500 110970 5560
rect 111030 5500 111040 5560
rect 110800 5480 111040 5500
rect 110800 5420 110810 5480
rect 110870 5420 110890 5480
rect 110950 5420 110970 5480
rect 111030 5420 111040 5480
rect 110800 5400 111040 5420
rect 110800 5340 110810 5400
rect 110870 5340 110890 5400
rect 110950 5340 110970 5400
rect 111030 5340 111040 5400
rect 109240 4990 109320 5000
rect 109240 4930 109250 4990
rect 109310 4930 109320 4990
rect 109240 4910 109320 4930
rect 109240 4850 109250 4910
rect 109310 4850 109320 4910
rect 109240 4830 109320 4850
rect 109240 4770 109250 4830
rect 109310 4770 109320 4830
rect 109240 4760 109320 4770
rect 110560 4990 110640 5000
rect 110560 4930 110570 4990
rect 110630 4930 110640 4990
rect 110560 4910 110640 4930
rect 110560 4850 110570 4910
rect 110630 4850 110640 4910
rect 110560 4830 110640 4850
rect 110560 4770 110570 4830
rect 110630 4770 110640 4830
rect 110560 4760 110640 4770
rect 107980 4060 108000 4120
rect 108060 4060 108100 4120
rect 108160 4060 108200 4120
rect 108260 4060 108300 4120
rect 108360 4060 108400 4120
rect 108460 4060 108480 4120
rect 107980 4020 108480 4060
rect 107980 3960 108000 4020
rect 108060 3960 108100 4020
rect 108160 3960 108200 4020
rect 108260 3960 108300 4020
rect 108360 3960 108400 4020
rect 108460 3960 108480 4020
rect 109250 4470 109310 4760
rect 109350 4720 109430 4730
rect 109350 4660 109360 4720
rect 109420 4660 109430 4720
rect 109350 4640 109430 4660
rect 109350 4580 109360 4640
rect 109420 4580 109430 4640
rect 109350 4560 109430 4580
rect 109350 4500 109360 4560
rect 109420 4500 109430 4560
rect 109350 4490 109430 4500
rect 109570 4720 109650 4730
rect 109570 4660 109580 4720
rect 109640 4660 109650 4720
rect 109570 4640 109650 4660
rect 109570 4580 109580 4640
rect 109640 4580 109650 4640
rect 109570 4560 109650 4580
rect 109570 4500 109580 4560
rect 109640 4500 109650 4560
rect 109570 4490 109650 4500
rect 109790 4720 109870 4730
rect 109790 4660 109800 4720
rect 109860 4660 109870 4720
rect 109790 4640 109870 4660
rect 109790 4580 109800 4640
rect 109860 4580 109870 4640
rect 109790 4560 109870 4580
rect 109790 4500 109800 4560
rect 109860 4500 109870 4560
rect 109790 4490 109870 4500
rect 110010 4720 110090 4730
rect 110010 4660 110020 4720
rect 110080 4660 110090 4720
rect 110010 4640 110090 4660
rect 110010 4580 110020 4640
rect 110080 4580 110090 4640
rect 110010 4560 110090 4580
rect 110010 4500 110020 4560
rect 110080 4500 110090 4560
rect 110010 4490 110090 4500
rect 110230 4720 110310 4730
rect 110230 4660 110240 4720
rect 110300 4660 110310 4720
rect 110230 4640 110310 4660
rect 110230 4580 110240 4640
rect 110300 4580 110310 4640
rect 110230 4560 110310 4580
rect 110230 4500 110240 4560
rect 110300 4500 110310 4560
rect 110230 4490 110310 4500
rect 110450 4720 110530 4730
rect 110450 4660 110460 4720
rect 110520 4660 110530 4720
rect 110450 4640 110530 4660
rect 110450 4580 110460 4640
rect 110520 4580 110530 4640
rect 110450 4560 110530 4580
rect 110450 4500 110460 4560
rect 110520 4500 110530 4560
rect 110450 4490 110530 4500
rect 109250 4430 109260 4470
rect 109300 4430 109310 4470
rect 109250 4350 109310 4430
rect 109250 4010 109260 4350
rect 109300 4010 109310 4350
rect 109250 3990 109310 4010
rect 109360 4350 109420 4490
rect 109460 4450 109540 4460
rect 109460 4390 109470 4450
rect 109530 4390 109540 4450
rect 109460 4380 109540 4390
rect 109360 4010 109370 4350
rect 109410 4010 109420 4350
rect 109360 3990 109420 4010
rect 109470 4350 109530 4380
rect 109470 4010 109480 4350
rect 109520 4010 109530 4350
rect 107980 3920 108480 3960
rect 109470 3950 109530 4010
rect 109580 4350 109640 4490
rect 109680 4450 109760 4460
rect 109680 4390 109690 4450
rect 109750 4390 109760 4450
rect 109680 4380 109760 4390
rect 109580 4010 109590 4350
rect 109630 4010 109640 4350
rect 109580 3990 109640 4010
rect 109690 4350 109750 4380
rect 109690 4010 109700 4350
rect 109740 4010 109750 4350
rect 109690 3950 109750 4010
rect 109800 4350 109860 4490
rect 109900 4450 109980 4460
rect 109900 4390 109910 4450
rect 109970 4390 109980 4450
rect 109900 4380 109980 4390
rect 109800 4010 109810 4350
rect 109850 4010 109860 4350
rect 109800 3990 109860 4010
rect 109910 4350 109970 4380
rect 109910 4010 109920 4350
rect 109960 4010 109970 4350
rect 109910 3950 109970 4010
rect 110020 4350 110080 4490
rect 110120 4450 110200 4460
rect 110120 4390 110130 4450
rect 110190 4390 110200 4450
rect 110120 4380 110200 4390
rect 110020 4010 110030 4350
rect 110070 4010 110080 4350
rect 110020 3990 110080 4010
rect 110130 4350 110190 4380
rect 110130 4010 110140 4350
rect 110180 4010 110190 4350
rect 110130 3950 110190 4010
rect 110240 4350 110300 4490
rect 110340 4450 110420 4460
rect 110340 4390 110350 4450
rect 110410 4390 110420 4450
rect 110340 4380 110420 4390
rect 110240 4010 110250 4350
rect 110290 4010 110300 4350
rect 110240 3990 110300 4010
rect 110350 4350 110410 4380
rect 110350 4010 110360 4350
rect 110400 4010 110410 4350
rect 110350 3950 110410 4010
rect 110460 4350 110520 4490
rect 110460 4010 110470 4350
rect 110510 4010 110520 4350
rect 110460 3990 110520 4010
rect 110570 4470 110630 4760
rect 110570 4430 110580 4470
rect 110620 4430 110630 4470
rect 110570 4350 110630 4430
rect 110570 4010 110580 4350
rect 110620 4010 110630 4350
rect 110570 3990 110630 4010
rect 107980 3860 108000 3920
rect 108060 3860 108100 3920
rect 108160 3860 108200 3920
rect 108260 3860 108300 3920
rect 108360 3860 108400 3920
rect 108460 3860 108480 3920
rect 108970 3940 109050 3950
rect 108970 3880 108980 3940
rect 109040 3880 109050 3940
rect 108970 3870 109050 3880
rect 109460 3940 109540 3950
rect 109460 3880 109470 3940
rect 109530 3880 109540 3940
rect 109460 3870 109540 3880
rect 109680 3940 109760 3950
rect 109680 3880 109690 3940
rect 109750 3880 109760 3940
rect 109680 3870 109760 3880
rect 109900 3940 109980 3950
rect 109900 3880 109910 3940
rect 109970 3880 109980 3940
rect 109900 3870 109980 3880
rect 110120 3940 110200 3950
rect 110120 3880 110130 3940
rect 110190 3880 110200 3940
rect 110120 3870 110200 3880
rect 110340 3940 110420 3950
rect 110340 3880 110350 3940
rect 110410 3880 110420 3940
rect 110340 3870 110420 3880
rect 107980 1740 108480 3860
rect 108510 2940 108580 2952
rect 108510 2860 108580 2870
rect 108630 2940 108700 2950
rect 108630 2860 108700 2870
rect 108750 2940 108820 2950
rect 108750 2860 108820 2870
rect 108870 2940 108940 2950
rect 108870 2860 108940 2870
rect 108530 2240 108570 2860
rect 108770 2800 108810 2860
rect 108990 2800 109030 3870
rect 110230 3810 110310 3820
rect 110230 3750 110240 3810
rect 110300 3750 110310 3810
rect 110230 3730 110310 3750
rect 110230 3670 110240 3730
rect 110300 3670 110310 3730
rect 110230 3660 110310 3670
rect 110800 3810 111040 5340
rect 110800 3750 110810 3810
rect 110870 3750 110890 3810
rect 110950 3750 110970 3810
rect 111030 3750 111040 3810
rect 110800 3730 111040 3750
rect 110800 3670 110810 3730
rect 110870 3670 110890 3730
rect 110950 3670 110970 3730
rect 111030 3670 111040 3730
rect 109060 3570 109140 3580
rect 109060 3510 109070 3570
rect 109130 3510 109140 3570
rect 109060 3500 109140 3510
rect 109460 3570 109540 3580
rect 109460 3510 109470 3570
rect 109530 3510 109540 3570
rect 109460 3500 109540 3510
rect 109680 3570 109760 3580
rect 109680 3510 109690 3570
rect 109750 3510 109760 3570
rect 109680 3500 109760 3510
rect 109900 3570 109980 3580
rect 109900 3510 109910 3570
rect 109970 3510 109980 3570
rect 109900 3500 109980 3510
rect 110120 3570 110200 3580
rect 110120 3510 110130 3570
rect 110190 3510 110200 3570
rect 110120 3500 110200 3510
rect 110340 3570 110420 3580
rect 110340 3510 110350 3570
rect 110410 3510 110420 3570
rect 110340 3500 110420 3510
rect 109080 2940 109120 3500
rect 109250 3470 109310 3490
rect 109060 2930 109140 2940
rect 109060 2870 109070 2930
rect 109130 2870 109140 2930
rect 109060 2860 109140 2870
rect 109250 2930 109260 3470
rect 109300 2930 109310 3470
rect 109250 2850 109310 2930
rect 109250 2810 109260 2850
rect 109300 2810 109310 2850
rect 108750 2790 108830 2800
rect 108750 2730 108760 2790
rect 108820 2730 108830 2790
rect 108750 2720 108830 2730
rect 108970 2790 109050 2800
rect 108970 2730 108980 2790
rect 109040 2730 109050 2790
rect 108970 2720 109050 2730
rect 109250 2510 109310 2810
rect 109360 3470 109420 3490
rect 109360 2930 109370 3470
rect 109410 2930 109420 3470
rect 109360 2790 109420 2930
rect 109470 3470 109530 3500
rect 109470 2930 109480 3470
rect 109520 2930 109530 3470
rect 109470 2900 109530 2930
rect 109580 3470 109640 3490
rect 109580 2930 109590 3470
rect 109630 2930 109640 3470
rect 109460 2890 109540 2900
rect 109460 2830 109470 2890
rect 109530 2830 109540 2890
rect 109460 2820 109540 2830
rect 109580 2790 109640 2930
rect 109690 3470 109750 3500
rect 109690 2930 109700 3470
rect 109740 2930 109750 3470
rect 109690 2900 109750 2930
rect 109800 3470 109860 3490
rect 109800 2930 109810 3470
rect 109850 2930 109860 3470
rect 109680 2890 109760 2900
rect 109680 2830 109690 2890
rect 109750 2830 109760 2890
rect 109680 2820 109760 2830
rect 109800 2790 109860 2930
rect 109910 3470 109970 3500
rect 109910 2930 109920 3470
rect 109960 2930 109970 3470
rect 109910 2900 109970 2930
rect 110020 3470 110080 3490
rect 110020 2930 110030 3470
rect 110070 2930 110080 3470
rect 109900 2890 109980 2900
rect 109900 2830 109910 2890
rect 109970 2830 109980 2890
rect 109900 2820 109980 2830
rect 110020 2790 110080 2930
rect 110130 3470 110190 3500
rect 110130 2930 110140 3470
rect 110180 2930 110190 3470
rect 110130 2900 110190 2930
rect 110240 3470 110300 3490
rect 110240 2930 110250 3470
rect 110290 2930 110300 3470
rect 110120 2890 110200 2900
rect 110120 2830 110130 2890
rect 110190 2830 110200 2890
rect 110120 2820 110200 2830
rect 110240 2790 110300 2930
rect 110350 3470 110410 3500
rect 110350 2930 110360 3470
rect 110400 2930 110410 3470
rect 110350 2900 110410 2930
rect 110460 3470 110520 3490
rect 110460 2930 110470 3470
rect 110510 2930 110520 3470
rect 110340 2890 110420 2900
rect 110340 2830 110350 2890
rect 110410 2830 110420 2890
rect 110340 2820 110420 2830
rect 110460 2790 110520 2930
rect 110570 3470 110630 3490
rect 110570 2930 110580 3470
rect 110620 2930 110630 3470
rect 110570 2850 110630 2930
rect 110570 2810 110580 2850
rect 110620 2810 110630 2850
rect 110800 3050 111040 3670
rect 110800 2990 110810 3050
rect 110870 2990 110890 3050
rect 110950 2990 110970 3050
rect 111030 2990 111040 3050
rect 110800 2970 111040 2990
rect 110800 2910 110810 2970
rect 110870 2910 110890 2970
rect 110950 2910 110970 2970
rect 111030 2910 111040 2970
rect 110800 2890 111040 2910
rect 110800 2830 110810 2890
rect 110870 2830 110890 2890
rect 110950 2830 110970 2890
rect 111030 2830 111040 2890
rect 110800 2820 111040 2830
rect 111070 7350 111310 8240
rect 111360 7470 111400 8610
rect 113020 8460 113100 8470
rect 113020 8400 113030 8460
rect 113090 8400 113100 8460
rect 113020 8380 113100 8400
rect 113020 8320 113030 8380
rect 113090 8320 113100 8380
rect 113020 8300 113100 8320
rect 113020 8240 113030 8300
rect 113090 8240 113100 8300
rect 113020 8230 113100 8240
rect 113360 8460 113420 8470
rect 113360 8380 113420 8400
rect 113360 8300 113420 8320
rect 113360 8230 113420 8240
rect 113680 8460 113920 9200
rect 114260 9470 114320 9530
rect 114260 8830 114270 9470
rect 114310 8830 114320 9470
rect 114260 8810 114320 8830
rect 114380 9470 114440 9800
rect 114490 9760 114570 9770
rect 114490 9700 114500 9760
rect 114560 9700 114570 9760
rect 114490 9680 114570 9700
rect 114490 9620 114500 9680
rect 114560 9620 114570 9680
rect 114490 9600 114570 9620
rect 114490 9540 114500 9600
rect 114560 9540 114570 9600
rect 114490 9530 114570 9540
rect 114610 9760 114690 9770
rect 114610 9700 114620 9760
rect 114680 9700 114690 9760
rect 114610 9680 114690 9700
rect 114610 9620 114620 9680
rect 114680 9620 114690 9680
rect 114610 9600 114690 9620
rect 114610 9540 114620 9600
rect 114680 9540 114690 9600
rect 114610 9530 114690 9540
rect 114380 8830 114390 9470
rect 114430 8830 114440 9470
rect 114380 8800 114440 8830
rect 114500 9470 114560 9530
rect 114500 8830 114510 9470
rect 114550 8830 114560 9470
rect 114500 8810 114560 8830
rect 114620 9470 114680 9530
rect 114620 8830 114630 9470
rect 114670 8830 114680 9470
rect 114620 8810 114680 8830
rect 114370 8790 114450 8800
rect 114370 8730 114380 8790
rect 114440 8730 114450 8790
rect 114370 8720 114450 8730
rect 114480 8670 114540 8690
rect 114480 8630 114490 8670
rect 114530 8630 114540 8670
rect 114480 8580 114540 8630
rect 114470 8570 114550 8580
rect 114470 8510 114480 8570
rect 114540 8510 114550 8570
rect 114470 8500 114550 8510
rect 114900 8570 114980 9920
rect 116970 9980 117030 9990
rect 116970 9910 117030 9920
rect 117090 9980 117150 9990
rect 117090 9910 117150 9920
rect 117210 9980 117270 9990
rect 117210 9910 117270 9920
rect 117330 9980 117390 9990
rect 117330 9910 117390 9920
rect 117450 9980 117630 9990
rect 117510 9920 117570 9980
rect 117450 9910 117630 9920
rect 117690 9980 117750 9990
rect 117690 9910 117750 9920
rect 117810 9980 117870 9990
rect 117810 9910 117870 9920
rect 117930 9980 117990 9990
rect 117930 9910 117990 9920
rect 118050 9980 118110 9990
rect 118050 9910 118110 9920
rect 115310 9870 115390 9880
rect 115310 9810 115320 9870
rect 115380 9810 115390 9870
rect 115190 9600 115270 9610
rect 115190 9540 115200 9600
rect 115260 9540 115270 9600
rect 115190 9530 115270 9540
rect 115310 9600 115390 9810
rect 116900 9870 116980 9880
rect 116900 9810 116910 9870
rect 116970 9810 116980 9870
rect 116900 9800 116980 9810
rect 117140 9870 117220 9880
rect 117140 9810 117150 9870
rect 117210 9810 117220 9870
rect 117140 9800 117220 9810
rect 117380 9870 117460 9880
rect 117380 9810 117390 9870
rect 117450 9810 117460 9870
rect 117380 9800 117460 9810
rect 117620 9870 117700 9880
rect 117620 9810 117630 9870
rect 117690 9810 117700 9870
rect 117620 9800 117700 9810
rect 117860 9870 117940 9880
rect 117860 9810 117870 9870
rect 117930 9810 117940 9870
rect 117860 9800 117940 9810
rect 118100 9870 118180 9880
rect 118100 9810 118110 9870
rect 118170 9810 118180 9870
rect 118100 9800 118180 9810
rect 116790 9770 116850 9790
rect 115310 9540 115320 9600
rect 115380 9540 115390 9600
rect 115310 9530 115390 9540
rect 115550 9600 115630 9610
rect 115550 9540 115560 9600
rect 115620 9540 115630 9600
rect 115550 9530 115630 9540
rect 115200 9470 115260 9530
rect 115200 8830 115210 9470
rect 115250 8830 115260 9470
rect 115200 8810 115260 8830
rect 115320 9470 115380 9530
rect 115320 8830 115330 9470
rect 115370 8830 115380 9470
rect 115320 8800 115380 8830
rect 115440 9470 115500 9490
rect 115440 8830 115450 9470
rect 115490 8830 115500 9470
rect 115310 8790 115390 8800
rect 115310 8730 115320 8790
rect 115380 8730 115390 8790
rect 115310 8720 115390 8730
rect 115352 8680 115412 8690
rect 115352 8610 115412 8620
rect 115440 8580 115500 8830
rect 115560 9470 115620 9530
rect 115560 8830 115570 9470
rect 115610 8830 115620 9470
rect 116790 9130 116800 9770
rect 116840 9130 116850 9770
rect 116790 9070 116850 9130
rect 116910 9770 116970 9800
rect 116910 9130 116920 9770
rect 116960 9130 116970 9770
rect 115560 8810 115620 8830
rect 116290 9060 116530 9070
rect 116290 9000 116300 9060
rect 116360 9000 116380 9060
rect 116440 9000 116460 9060
rect 116520 9000 116530 9060
rect 116180 8680 116260 8690
rect 116180 8620 116190 8680
rect 116250 8620 116260 8680
rect 116180 8610 116260 8620
rect 114900 8510 114910 8570
rect 114970 8510 114980 8570
rect 114900 8500 114980 8510
rect 115430 8570 115510 8580
rect 115430 8510 115440 8570
rect 115500 8510 115510 8570
rect 115430 8500 115510 8510
rect 113680 8400 113690 8460
rect 113750 8400 113850 8460
rect 113910 8400 113920 8460
rect 113680 8380 113920 8400
rect 113680 8320 113690 8380
rect 113750 8320 113850 8380
rect 113910 8320 113920 8380
rect 113680 8300 113920 8320
rect 113680 8240 113690 8300
rect 113750 8240 113850 8300
rect 113910 8240 113920 8300
rect 113680 8230 113920 8240
rect 114180 8460 114240 8470
rect 114180 8380 114240 8400
rect 114180 8300 114240 8320
rect 114180 8230 114240 8240
rect 114500 8460 114580 8470
rect 114500 8400 114510 8460
rect 114570 8400 114580 8460
rect 114500 8380 114580 8400
rect 114500 8320 114510 8380
rect 114570 8320 114580 8380
rect 114500 8300 114580 8320
rect 114500 8240 114510 8300
rect 114570 8240 114580 8300
rect 114500 8230 114580 8240
rect 113240 8170 113320 8180
rect 113240 8110 113250 8170
rect 113310 8110 113320 8170
rect 113240 8100 113320 8110
rect 113460 8170 113540 8180
rect 113460 8110 113470 8170
rect 113530 8110 113540 8170
rect 113460 8100 113540 8110
rect 114060 8170 114140 8180
rect 114060 8110 114070 8170
rect 114130 8110 114140 8170
rect 114060 8100 114140 8110
rect 114280 8170 114360 8180
rect 114280 8110 114290 8170
rect 114350 8110 114360 8170
rect 114280 8100 114360 8110
rect 113120 7550 113180 7560
rect 113600 7550 113660 7560
rect 113120 7480 113180 7490
rect 113214 7520 113274 7540
rect 113214 7480 113224 7520
rect 113264 7480 113274 7520
rect 111340 7460 111420 7470
rect 113214 7460 113274 7480
rect 113350 7530 113430 7540
rect 113350 7470 113360 7530
rect 113420 7470 113430 7530
rect 113350 7460 113430 7470
rect 113506 7520 113566 7540
rect 113506 7480 113516 7520
rect 113556 7480 113566 7520
rect 113600 7480 113660 7490
rect 113940 7540 114000 7560
rect 114420 7540 114480 7560
rect 113940 7500 113950 7540
rect 113990 7500 114000 7540
rect 113940 7480 114000 7500
rect 114034 7520 114094 7540
rect 114034 7480 114044 7520
rect 114084 7480 114094 7520
rect 113506 7460 113566 7480
rect 111340 7400 111350 7460
rect 111410 7400 111420 7460
rect 113220 7420 113260 7460
rect 111340 7390 111420 7400
rect 113200 7410 113280 7420
rect 111070 7290 111080 7350
rect 111140 7290 111160 7350
rect 111220 7290 111240 7350
rect 111300 7290 111310 7350
rect 113200 7350 113210 7410
rect 113270 7350 113280 7410
rect 113200 7340 113280 7350
rect 113520 7300 113560 7460
rect 111070 7270 111310 7290
rect 111070 7210 111080 7270
rect 111140 7210 111160 7270
rect 111220 7210 111240 7270
rect 111300 7210 111310 7270
rect 111070 7190 111310 7210
rect 111070 7130 111080 7190
rect 111140 7130 111160 7190
rect 111220 7130 111240 7190
rect 111300 7130 111310 7190
rect 111070 4990 111310 7130
rect 111900 7290 111980 7300
rect 111900 7230 111910 7290
rect 111970 7230 111980 7290
rect 111900 7220 111980 7230
rect 113490 7290 113570 7300
rect 113490 7230 113500 7290
rect 113560 7230 113570 7290
rect 113490 7220 113570 7230
rect 111070 4930 111080 4990
rect 111140 4930 111160 4990
rect 111220 4930 111240 4990
rect 111300 4930 111310 4990
rect 111070 4910 111310 4930
rect 111070 4850 111080 4910
rect 111140 4850 111160 4910
rect 111220 4850 111240 4910
rect 111300 4850 111310 4910
rect 111070 4830 111310 4850
rect 111070 4770 111080 4830
rect 111140 4770 111160 4830
rect 111220 4770 111240 4830
rect 111300 4770 111310 4830
rect 109350 2780 109430 2790
rect 109350 2720 109360 2780
rect 109420 2720 109430 2780
rect 109350 2700 109430 2720
rect 109350 2640 109360 2700
rect 109420 2640 109430 2700
rect 109350 2620 109430 2640
rect 109350 2560 109360 2620
rect 109420 2560 109430 2620
rect 109350 2550 109430 2560
rect 109570 2780 109650 2790
rect 109570 2720 109580 2780
rect 109640 2720 109650 2780
rect 109570 2700 109650 2720
rect 109570 2640 109580 2700
rect 109640 2640 109650 2700
rect 109570 2620 109650 2640
rect 109570 2560 109580 2620
rect 109640 2560 109650 2620
rect 109570 2550 109650 2560
rect 109790 2780 109870 2790
rect 109790 2720 109800 2780
rect 109860 2720 109870 2780
rect 109790 2700 109870 2720
rect 109790 2640 109800 2700
rect 109860 2640 109870 2700
rect 109790 2620 109870 2640
rect 109790 2560 109800 2620
rect 109860 2560 109870 2620
rect 109790 2550 109870 2560
rect 110010 2780 110090 2790
rect 110010 2720 110020 2780
rect 110080 2720 110090 2780
rect 110010 2700 110090 2720
rect 110010 2640 110020 2700
rect 110080 2640 110090 2700
rect 110010 2620 110090 2640
rect 110010 2560 110020 2620
rect 110080 2560 110090 2620
rect 110010 2550 110090 2560
rect 110230 2780 110310 2790
rect 110230 2720 110240 2780
rect 110300 2720 110310 2780
rect 110230 2700 110310 2720
rect 110230 2640 110240 2700
rect 110300 2640 110310 2700
rect 110230 2620 110310 2640
rect 110230 2560 110240 2620
rect 110300 2560 110310 2620
rect 110230 2550 110310 2560
rect 110450 2780 110530 2790
rect 110450 2720 110460 2780
rect 110520 2720 110530 2780
rect 110450 2700 110530 2720
rect 110450 2640 110460 2700
rect 110520 2640 110530 2700
rect 110450 2620 110530 2640
rect 110450 2560 110460 2620
rect 110520 2560 110530 2620
rect 110450 2550 110530 2560
rect 110570 2510 110630 2810
rect 111070 2780 111310 4770
rect 111340 6320 111580 6330
rect 111340 6260 111350 6320
rect 111410 6260 111430 6320
rect 111490 6260 111510 6320
rect 111570 6260 111580 6320
rect 111340 6240 111580 6260
rect 111340 6180 111350 6240
rect 111410 6180 111430 6240
rect 111490 6180 111510 6240
rect 111570 6180 111580 6240
rect 111340 6160 111580 6180
rect 111340 6100 111350 6160
rect 111410 6100 111430 6160
rect 111490 6100 111510 6160
rect 111570 6100 111580 6160
rect 111340 6020 111580 6100
rect 111340 5960 111350 6020
rect 111410 5960 111430 6020
rect 111490 5960 111510 6020
rect 111570 5960 111580 6020
rect 111340 5940 111580 5960
rect 111340 5880 111350 5940
rect 111410 5880 111430 5940
rect 111490 5880 111510 5940
rect 111570 5880 111580 5940
rect 111340 5860 111580 5880
rect 111340 5800 111350 5860
rect 111410 5800 111430 5860
rect 111490 5800 111510 5860
rect 111570 5800 111580 5860
rect 111340 5200 111580 5800
rect 111340 5140 111350 5200
rect 111410 5140 111430 5200
rect 111490 5140 111510 5200
rect 111570 5140 111580 5200
rect 111340 5120 111580 5140
rect 111340 5060 111350 5120
rect 111410 5060 111430 5120
rect 111490 5060 111510 5120
rect 111570 5060 111580 5120
rect 111340 5040 111580 5060
rect 111340 4980 111350 5040
rect 111410 4980 111430 5040
rect 111490 4980 111510 5040
rect 111570 4980 111580 5040
rect 111340 4720 111580 4980
rect 111340 4660 111350 4720
rect 111410 4660 111430 4720
rect 111490 4660 111510 4720
rect 111570 4660 111580 4720
rect 111340 4640 111580 4660
rect 111340 4580 111350 4640
rect 111410 4580 111430 4640
rect 111490 4580 111510 4640
rect 111570 4580 111580 4640
rect 111340 4560 111580 4580
rect 111340 4500 111350 4560
rect 111410 4500 111430 4560
rect 111490 4500 111510 4560
rect 111570 4500 111580 4560
rect 111340 4490 111580 4500
rect 111690 5830 111770 5840
rect 111690 5770 111700 5830
rect 111760 5770 111770 5830
rect 111070 2720 111080 2780
rect 111140 2720 111160 2780
rect 111220 2720 111240 2780
rect 111300 2720 111310 2780
rect 111070 2700 111310 2720
rect 111070 2640 111080 2700
rect 111140 2640 111160 2700
rect 111220 2640 111240 2700
rect 111300 2640 111310 2700
rect 111070 2620 111310 2640
rect 111070 2560 111080 2620
rect 111140 2560 111160 2620
rect 111220 2560 111240 2620
rect 111300 2560 111310 2620
rect 111070 2550 111310 2560
rect 111340 4390 111580 4400
rect 111340 4330 111350 4390
rect 111410 4330 111430 4390
rect 111490 4330 111510 4390
rect 111570 4330 111580 4390
rect 111340 4310 111580 4330
rect 111340 4250 111350 4310
rect 111410 4250 111430 4310
rect 111490 4250 111510 4310
rect 111570 4250 111580 4310
rect 111340 4230 111580 4250
rect 111340 4170 111350 4230
rect 111410 4170 111430 4230
rect 111490 4170 111510 4230
rect 111570 4170 111580 4230
rect 109240 2500 109320 2510
rect 109240 2440 109250 2500
rect 109310 2440 109320 2500
rect 109240 2420 109320 2440
rect 109240 2360 109250 2420
rect 109310 2360 109320 2420
rect 109240 2340 109320 2360
rect 109240 2280 109250 2340
rect 109310 2280 109320 2340
rect 109240 2270 109320 2280
rect 110560 2500 110640 2510
rect 110560 2440 110570 2500
rect 110630 2440 110640 2500
rect 110560 2420 110640 2440
rect 110560 2360 110570 2420
rect 110630 2360 110640 2420
rect 110560 2340 110640 2360
rect 110560 2280 110570 2340
rect 110630 2280 110640 2340
rect 110560 2270 110640 2280
rect 108510 2230 108590 2240
rect 108510 2170 108520 2230
rect 108580 2170 108590 2230
rect 108510 2160 108590 2170
rect 107980 1680 107990 1740
rect 108050 1680 108070 1740
rect 108130 1680 108160 1740
rect 108220 1680 108240 1740
rect 108300 1680 108330 1740
rect 108390 1680 108410 1740
rect 108470 1680 108480 1740
rect 107980 1660 108480 1680
rect 107980 1600 107990 1660
rect 108050 1600 108070 1660
rect 108130 1600 108160 1660
rect 108220 1600 108240 1660
rect 108300 1600 108330 1660
rect 108390 1600 108410 1660
rect 108470 1600 108480 1660
rect 107980 1580 108480 1600
rect 107980 1520 107990 1580
rect 108050 1520 108070 1580
rect 108130 1520 108160 1580
rect 108220 1520 108240 1580
rect 108300 1520 108330 1580
rect 108390 1520 108410 1580
rect 108470 1520 108480 1580
rect 107980 1510 108480 1520
rect 108640 1850 108720 1860
rect 108640 1790 108650 1850
rect 108710 1790 108720 1850
rect 108640 1470 108720 1790
rect 108640 1410 108650 1470
rect 108710 1410 108720 1470
rect 108640 1370 108720 1410
rect 108650 1360 108720 1370
rect 108650 1280 108720 1290
rect 108770 1740 108850 1750
rect 108770 1680 108780 1740
rect 108840 1680 108850 1740
rect 108770 1660 108850 1680
rect 108770 1600 108780 1660
rect 108840 1600 108850 1660
rect 108770 1580 108850 1600
rect 108770 1520 108780 1580
rect 108840 1520 108850 1580
rect 108770 1510 108850 1520
rect 109500 1740 110380 1750
rect 109500 1680 109510 1740
rect 109570 1680 109590 1740
rect 109650 1680 109670 1740
rect 109730 1680 109750 1740
rect 109810 1680 109830 1740
rect 109890 1680 109910 1740
rect 109970 1680 109990 1740
rect 110050 1680 110070 1740
rect 110130 1680 110150 1740
rect 110210 1680 110230 1740
rect 110290 1680 110310 1740
rect 110370 1680 110380 1740
rect 109500 1660 110380 1680
rect 109500 1600 109510 1660
rect 109570 1600 109590 1660
rect 109650 1600 109670 1660
rect 109730 1600 109750 1660
rect 109810 1600 109830 1660
rect 109890 1600 109910 1660
rect 109970 1600 109990 1660
rect 110050 1600 110070 1660
rect 110130 1600 110150 1660
rect 110210 1600 110230 1660
rect 110290 1600 110310 1660
rect 110370 1600 110380 1660
rect 109500 1580 110380 1600
rect 109500 1520 109510 1580
rect 109570 1520 109590 1580
rect 109650 1520 109670 1580
rect 109730 1520 109750 1580
rect 109810 1520 109830 1580
rect 109890 1520 109910 1580
rect 109970 1520 109990 1580
rect 110050 1520 110070 1580
rect 110130 1520 110150 1580
rect 110210 1520 110230 1580
rect 110290 1520 110310 1580
rect 110370 1520 110380 1580
rect 109500 1510 110380 1520
rect 108770 1360 108840 1510
rect 108770 1280 108840 1290
rect 109310 1350 109370 1370
rect 109310 10 109320 1350
rect 109360 10 109370 1350
rect 109310 -70 109370 10
rect 109510 1350 109570 1510
rect 109600 1470 109680 1480
rect 109600 1410 109610 1470
rect 109670 1410 109680 1470
rect 109600 1400 109680 1410
rect 109800 1470 109880 1480
rect 109800 1410 109810 1470
rect 109870 1410 109880 1470
rect 109800 1400 109880 1410
rect 109510 10 109520 1350
rect 109560 10 109570 1350
rect 109510 -20 109570 10
rect 109710 1350 109770 1370
rect 109710 10 109720 1350
rect 109760 10 109770 1350
rect 109310 -110 109320 -70
rect 109360 -110 109370 -70
rect 109500 -30 109580 -20
rect 109500 -90 109510 -30
rect 109570 -90 109580 -30
rect 109500 -100 109580 -90
rect 109310 -1150 109370 -110
rect 109710 -1150 109770 10
rect 109910 1350 109970 1510
rect 110000 1470 110080 1480
rect 110000 1410 110010 1470
rect 110070 1410 110080 1470
rect 110000 1400 110080 1410
rect 110200 1470 110280 1480
rect 110200 1410 110210 1470
rect 110270 1410 110280 1470
rect 110200 1400 110280 1410
rect 109910 10 109920 1350
rect 109960 10 109970 1350
rect 109910 -20 109970 10
rect 110110 1350 110170 1370
rect 110110 10 110120 1350
rect 110160 10 110170 1350
rect 109900 -30 109980 -20
rect 109900 -90 109910 -30
rect 109970 -90 109980 -30
rect 109900 -100 109980 -90
rect 107680 -1220 107690 -1160
rect 107750 -1220 107770 -1160
rect 107830 -1220 107850 -1160
rect 107910 -1220 107920 -1160
rect 107680 -1240 107920 -1220
rect 107680 -1300 107690 -1240
rect 107750 -1300 107770 -1240
rect 107830 -1300 107850 -1240
rect 107910 -1300 107920 -1240
rect 107680 -1320 107920 -1300
rect 107680 -1380 107690 -1320
rect 107750 -1380 107770 -1320
rect 107830 -1380 107850 -1320
rect 107910 -1380 107920 -1320
rect 107680 -1390 107920 -1380
rect 108080 -1160 108320 -1150
rect 108080 -1220 108090 -1160
rect 108150 -1220 108170 -1160
rect 108230 -1220 108250 -1160
rect 108310 -1220 108320 -1160
rect 108080 -1240 108320 -1220
rect 108080 -1300 108090 -1240
rect 108150 -1300 108170 -1240
rect 108230 -1300 108250 -1240
rect 108310 -1300 108320 -1240
rect 108080 -1320 108320 -1300
rect 108080 -1380 108090 -1320
rect 108150 -1380 108170 -1320
rect 108230 -1380 108250 -1320
rect 108310 -1380 108320 -1320
rect 108080 -3000 108320 -1380
rect 108780 -1160 109020 -1150
rect 108780 -1220 108790 -1160
rect 108850 -1220 108870 -1160
rect 108930 -1220 108950 -1160
rect 109010 -1220 109020 -1160
rect 108780 -1240 109020 -1220
rect 108780 -1300 108790 -1240
rect 108850 -1300 108870 -1240
rect 108930 -1300 108950 -1240
rect 109010 -1300 109020 -1240
rect 108780 -1320 109020 -1300
rect 108780 -1380 108790 -1320
rect 108850 -1380 108870 -1320
rect 108930 -1380 108950 -1320
rect 109010 -1380 109020 -1320
rect 108780 -3000 109020 -1380
rect 109300 -1160 109380 -1150
rect 109300 -1220 109310 -1160
rect 109370 -1220 109380 -1160
rect 109300 -1240 109380 -1220
rect 109300 -1300 109310 -1240
rect 109370 -1300 109380 -1240
rect 109300 -1320 109380 -1300
rect 109300 -1380 109310 -1320
rect 109370 -1380 109380 -1320
rect 109300 -1390 109380 -1380
rect 109480 -1160 109770 -1150
rect 109480 -1220 109490 -1160
rect 109550 -1220 109570 -1160
rect 109630 -1220 109650 -1160
rect 109710 -1220 109770 -1160
rect 109480 -1240 109770 -1220
rect 109480 -1300 109490 -1240
rect 109550 -1300 109570 -1240
rect 109630 -1300 109650 -1240
rect 109710 -1300 109770 -1240
rect 109480 -1320 109770 -1300
rect 109480 -1380 109490 -1320
rect 109550 -1380 109570 -1320
rect 109630 -1380 109650 -1320
rect 109710 -1380 109770 -1320
rect 109480 -1390 109770 -1380
rect 110110 -1150 110170 10
rect 110310 1350 110370 1510
rect 110310 10 110320 1350
rect 110360 10 110370 1350
rect 110310 -20 110370 10
rect 110510 1350 110570 1370
rect 110510 10 110520 1350
rect 110560 10 110570 1350
rect 111340 580 111580 4170
rect 111340 520 111350 580
rect 111410 520 111430 580
rect 111490 520 111510 580
rect 111570 520 111580 580
rect 111340 500 111580 520
rect 111340 440 111350 500
rect 111410 440 111430 500
rect 111490 440 111510 500
rect 111570 440 111580 500
rect 111340 420 111580 440
rect 111340 360 111350 420
rect 111410 360 111430 420
rect 111490 360 111510 420
rect 111570 360 111580 420
rect 111340 350 111580 360
rect 111690 200 111770 5770
rect 111900 2240 111940 7220
rect 113940 7190 113980 7480
rect 114034 7460 114094 7480
rect 114170 7530 114250 7540
rect 114170 7470 114180 7530
rect 114240 7470 114250 7530
rect 114170 7460 114250 7470
rect 114326 7520 114386 7540
rect 114326 7480 114336 7520
rect 114376 7480 114386 7520
rect 114420 7500 114430 7540
rect 114470 7500 114480 7540
rect 114420 7480 114480 7500
rect 114326 7460 114386 7480
rect 114040 7300 114080 7460
rect 114340 7420 114380 7460
rect 114320 7410 114400 7420
rect 114320 7350 114330 7410
rect 114390 7350 114400 7410
rect 114320 7340 114400 7350
rect 114030 7290 114110 7300
rect 114030 7230 114040 7290
rect 114100 7230 114110 7290
rect 114030 7220 114110 7230
rect 113700 7180 113780 7190
rect 113700 7120 113710 7180
rect 113770 7120 113780 7180
rect 113700 7110 113780 7120
rect 113920 7180 114000 7190
rect 113920 7120 113930 7180
rect 113990 7120 114000 7180
rect 113920 7110 114000 7120
rect 113720 6970 113760 7110
rect 114440 7080 114480 7480
rect 116200 7470 116240 8610
rect 116290 8460 116530 9000
rect 116780 9060 116860 9070
rect 116780 9000 116790 9060
rect 116850 9000 116860 9060
rect 116780 8990 116860 9000
rect 116910 8960 116970 9130
rect 117030 9770 117090 9790
rect 117030 9130 117040 9770
rect 117080 9130 117090 9770
rect 117030 9070 117090 9130
rect 117150 9770 117210 9800
rect 117150 9130 117160 9770
rect 117200 9130 117210 9770
rect 117020 9060 117100 9070
rect 117020 9000 117030 9060
rect 117090 9000 117100 9060
rect 117020 8990 117100 9000
rect 117150 8960 117210 9130
rect 117270 9770 117330 9790
rect 117270 9130 117280 9770
rect 117320 9130 117330 9770
rect 117270 9070 117330 9130
rect 117390 9770 117450 9800
rect 117390 9130 117400 9770
rect 117440 9130 117450 9770
rect 117260 9060 117340 9070
rect 117260 9000 117270 9060
rect 117330 9000 117340 9060
rect 117260 8990 117340 9000
rect 117390 8960 117450 9130
rect 117510 9770 117570 9790
rect 117510 9130 117520 9770
rect 117560 9130 117570 9770
rect 117510 9070 117570 9130
rect 117630 9770 117690 9800
rect 117630 9130 117640 9770
rect 117680 9130 117690 9770
rect 117500 9060 117580 9070
rect 117500 9000 117510 9060
rect 117570 9000 117580 9060
rect 117500 8990 117580 9000
rect 117630 8960 117690 9130
rect 117750 9770 117810 9790
rect 117750 9130 117760 9770
rect 117800 9130 117810 9770
rect 117750 9070 117810 9130
rect 117870 9770 117930 9800
rect 117870 9130 117880 9770
rect 117920 9130 117930 9770
rect 117740 9060 117820 9070
rect 117740 9000 117750 9060
rect 117810 9000 117820 9060
rect 117740 8990 117820 9000
rect 117870 8960 117930 9130
rect 117990 9770 118050 9790
rect 117990 9130 118000 9770
rect 118040 9130 118050 9770
rect 117990 9070 118050 9130
rect 118110 9770 118170 9800
rect 118110 9130 118120 9770
rect 118160 9130 118170 9770
rect 117980 9060 118060 9070
rect 117980 9000 117990 9060
rect 118050 9000 118060 9060
rect 117980 8990 118060 9000
rect 118110 8960 118170 9130
rect 118230 9770 118290 9790
rect 118230 9130 118240 9770
rect 118280 9130 118290 9770
rect 118230 9070 118290 9130
rect 119280 9340 119520 12220
rect 119280 9280 119290 9340
rect 119350 9280 119370 9340
rect 119430 9280 119450 9340
rect 119510 9280 119520 9340
rect 119280 9260 119520 9280
rect 119280 9200 119290 9260
rect 119350 9200 119370 9260
rect 119430 9200 119450 9260
rect 119510 9200 119520 9260
rect 119280 9180 119520 9200
rect 119280 9120 119290 9180
rect 119350 9120 119370 9180
rect 119430 9120 119450 9180
rect 119510 9120 119520 9180
rect 118220 9060 118300 9070
rect 118220 9000 118230 9060
rect 118290 9000 118300 9060
rect 118220 8990 118300 9000
rect 116290 8400 116300 8460
rect 116360 8400 116380 8460
rect 116440 8400 116460 8460
rect 116520 8400 116530 8460
rect 116900 8950 118420 8960
rect 116900 8890 116910 8950
rect 116970 8890 117150 8950
rect 117210 8890 117390 8950
rect 117450 8890 117630 8950
rect 117690 8890 117870 8950
rect 117930 8890 118110 8950
rect 118170 8890 118350 8950
rect 118410 8890 118420 8950
rect 116900 8870 118420 8890
rect 116900 8810 116910 8870
rect 116970 8810 117150 8870
rect 117210 8810 117390 8870
rect 117450 8810 117630 8870
rect 117690 8810 117870 8870
rect 117930 8810 118110 8870
rect 118170 8810 118350 8870
rect 118410 8810 118420 8870
rect 116900 8790 118420 8810
rect 116900 8730 116910 8790
rect 116970 8730 117150 8790
rect 117210 8730 117390 8790
rect 117450 8730 117630 8790
rect 117690 8730 117870 8790
rect 117930 8730 118110 8790
rect 118170 8730 118350 8790
rect 118410 8730 118420 8790
rect 116900 8710 118420 8730
rect 116900 8650 116910 8710
rect 116970 8650 117150 8710
rect 117210 8650 117390 8710
rect 117450 8650 117630 8710
rect 117690 8650 117870 8710
rect 117930 8650 118110 8710
rect 118170 8650 118350 8710
rect 118410 8650 118420 8710
rect 116900 8630 118420 8650
rect 116900 8570 116910 8630
rect 116970 8570 117150 8630
rect 117210 8570 117390 8630
rect 117450 8570 117630 8630
rect 117690 8570 117870 8630
rect 117930 8570 118110 8630
rect 118170 8570 118350 8630
rect 118410 8570 118420 8630
rect 116900 8550 118420 8570
rect 116900 8490 116910 8550
rect 116970 8490 117150 8550
rect 117210 8490 117390 8550
rect 117450 8490 117630 8550
rect 117690 8490 117870 8550
rect 117930 8490 118110 8550
rect 118170 8490 118350 8550
rect 118410 8490 118420 8550
rect 116900 8470 118420 8490
rect 116900 8410 116910 8470
rect 116970 8410 117150 8470
rect 117210 8410 117390 8470
rect 117450 8410 117630 8470
rect 117690 8410 117870 8470
rect 117930 8410 118110 8470
rect 118170 8410 118350 8470
rect 118410 8410 118420 8470
rect 116900 8400 118420 8410
rect 116290 8380 116530 8400
rect 116290 8320 116300 8380
rect 116360 8320 116380 8380
rect 116440 8320 116460 8380
rect 116520 8320 116530 8380
rect 116290 8300 116530 8320
rect 116290 8240 116300 8300
rect 116360 8240 116380 8300
rect 116440 8240 116460 8300
rect 116520 8240 116530 8300
rect 116180 7460 116260 7470
rect 116180 7400 116190 7460
rect 116250 7400 116260 7460
rect 116180 7390 116260 7400
rect 116290 7350 116530 8240
rect 116910 8370 116970 8400
rect 116910 8330 116920 8370
rect 116960 8330 116970 8370
rect 116910 8250 116970 8330
rect 117020 8350 117100 8360
rect 117020 8290 117030 8350
rect 117090 8290 117100 8350
rect 117020 8280 117100 8290
rect 116910 7610 116920 8250
rect 116960 7610 116970 8250
rect 116910 7590 116970 7610
rect 117030 8250 117090 8280
rect 117030 7610 117040 8250
rect 117080 7610 117090 8250
rect 117030 7580 117090 7610
rect 117150 8250 117210 8400
rect 117260 8350 117340 8360
rect 117260 8290 117270 8350
rect 117330 8290 117340 8350
rect 117260 8280 117340 8290
rect 117150 7610 117160 8250
rect 117200 7610 117210 8250
rect 117150 7590 117210 7610
rect 117270 8250 117330 8280
rect 117270 7610 117280 8250
rect 117320 7610 117330 8250
rect 117270 7580 117330 7610
rect 117390 8250 117450 8400
rect 117500 8350 117580 8360
rect 117500 8290 117510 8350
rect 117570 8290 117580 8350
rect 117500 8280 117580 8290
rect 117390 7610 117400 8250
rect 117440 7610 117450 8250
rect 117390 7590 117450 7610
rect 117510 8250 117570 8280
rect 117510 7610 117520 8250
rect 117560 7610 117570 8250
rect 117510 7580 117570 7610
rect 117630 8250 117690 8400
rect 117740 8350 117820 8360
rect 117740 8290 117750 8350
rect 117810 8290 117820 8350
rect 117740 8280 117820 8290
rect 117630 7610 117640 8250
rect 117680 7610 117690 8250
rect 117630 7590 117690 7610
rect 117750 8250 117810 8280
rect 117750 7610 117760 8250
rect 117800 7610 117810 8250
rect 117750 7580 117810 7610
rect 117870 8250 117930 8400
rect 117980 8350 118060 8360
rect 117980 8290 117990 8350
rect 118050 8290 118060 8350
rect 117980 8280 118060 8290
rect 117870 7610 117880 8250
rect 117920 7610 117930 8250
rect 117870 7590 117930 7610
rect 117990 8250 118050 8280
rect 117990 7610 118000 8250
rect 118040 7610 118050 8250
rect 117990 7580 118050 7610
rect 118110 8250 118170 8400
rect 118350 8370 118410 8400
rect 118220 8350 118300 8360
rect 118220 8290 118230 8350
rect 118290 8290 118300 8350
rect 118220 8280 118300 8290
rect 118350 8330 118360 8370
rect 118400 8330 118410 8370
rect 118110 7610 118120 8250
rect 118160 7610 118170 8250
rect 118110 7590 118170 7610
rect 118230 8250 118290 8280
rect 118230 7610 118240 8250
rect 118280 7610 118290 8250
rect 118230 7580 118290 7610
rect 118350 8250 118410 8330
rect 118350 7610 118360 8250
rect 118400 7610 118410 8250
rect 118350 7590 118410 7610
rect 119010 7670 119090 7680
rect 119010 7610 119020 7670
rect 119080 7610 119090 7670
rect 115630 7290 115710 7300
rect 115630 7230 115640 7290
rect 115700 7230 115710 7290
rect 115630 7220 115710 7230
rect 116290 7290 116300 7350
rect 116360 7290 116380 7350
rect 116440 7290 116460 7350
rect 116520 7290 116530 7350
rect 116290 7270 116530 7290
rect 113870 7070 113950 7080
rect 113870 7010 113880 7070
rect 113940 7010 113950 7070
rect 113870 7000 113950 7010
rect 114420 7070 114500 7080
rect 114420 7010 114430 7070
rect 114490 7010 114500 7070
rect 114420 7000 114500 7010
rect 113890 6970 113930 7000
rect 112170 6960 113350 6970
rect 112170 6900 112180 6960
rect 112240 6900 112290 6960
rect 112350 6900 112400 6960
rect 112460 6900 112510 6960
rect 112570 6900 112620 6960
rect 112680 6900 112730 6960
rect 112790 6900 112840 6960
rect 112900 6900 112950 6960
rect 113010 6900 113060 6960
rect 113120 6900 113170 6960
rect 113230 6900 113280 6960
rect 113340 6900 113350 6960
rect 112170 6880 113350 6900
rect 112170 6820 112180 6880
rect 112240 6820 112290 6880
rect 112350 6820 112400 6880
rect 112460 6820 112510 6880
rect 112570 6820 112620 6880
rect 112680 6820 112730 6880
rect 112790 6820 112840 6880
rect 112900 6820 112950 6880
rect 113010 6820 113060 6880
rect 113120 6820 113170 6880
rect 113230 6820 113280 6880
rect 113340 6820 113350 6880
rect 113660 6960 113780 6970
rect 113660 6900 113710 6960
rect 113770 6900 113780 6960
rect 113660 6890 113780 6900
rect 113870 6950 113950 6970
rect 113870 6910 113890 6950
rect 113930 6910 113950 6950
rect 113870 6890 113950 6910
rect 114250 6960 115430 6970
rect 114250 6900 114260 6960
rect 114320 6900 114370 6960
rect 114430 6900 114480 6960
rect 114540 6900 114590 6960
rect 114650 6900 114700 6960
rect 114760 6900 114810 6960
rect 114870 6900 114920 6960
rect 114980 6900 115030 6960
rect 115090 6900 115140 6960
rect 115200 6900 115250 6960
rect 115310 6900 115360 6960
rect 115420 6900 115430 6960
rect 112170 6800 113350 6820
rect 112170 6740 112180 6800
rect 112240 6740 112290 6800
rect 112350 6740 112400 6800
rect 112460 6740 112510 6800
rect 112570 6740 112620 6800
rect 112680 6740 112730 6800
rect 112790 6740 112840 6800
rect 112900 6740 112950 6800
rect 113010 6740 113060 6800
rect 113120 6740 113170 6800
rect 113230 6740 113280 6800
rect 113340 6740 113350 6800
rect 112170 6730 113350 6740
rect 112170 5940 112250 6730
rect 112170 5880 112180 5940
rect 112240 5880 112250 5940
rect 112170 5870 112250 5880
rect 112390 5940 112470 6730
rect 112390 5880 112400 5940
rect 112460 5880 112470 5940
rect 112390 5870 112470 5880
rect 112610 5940 112690 6730
rect 112610 5880 112620 5940
rect 112680 5880 112690 5940
rect 112610 5870 112690 5880
rect 112830 5940 112910 6730
rect 112830 5880 112840 5940
rect 112900 5880 112910 5940
rect 112830 5870 112910 5880
rect 113050 5940 113130 6730
rect 113050 5880 113060 5940
rect 113120 5880 113130 5940
rect 113050 5870 113130 5880
rect 113270 5940 113350 6730
rect 113550 6830 113610 6850
rect 113550 6390 113560 6830
rect 113600 6390 113610 6830
rect 113550 6330 113610 6390
rect 113660 6830 113720 6890
rect 113660 6390 113670 6830
rect 113710 6390 113720 6830
rect 113660 6370 113720 6390
rect 113770 6830 113830 6850
rect 113770 6390 113780 6830
rect 113820 6390 113830 6830
rect 113770 6330 113830 6390
rect 113880 6830 113940 6890
rect 114250 6880 115430 6900
rect 113880 6390 113890 6830
rect 113930 6390 113940 6830
rect 113880 6370 113940 6390
rect 113990 6830 114050 6850
rect 113990 6390 114000 6830
rect 114040 6390 114050 6830
rect 113990 6330 114050 6390
rect 114250 6820 114260 6880
rect 114320 6820 114370 6880
rect 114430 6820 114480 6880
rect 114540 6820 114590 6880
rect 114650 6820 114700 6880
rect 114760 6820 114810 6880
rect 114870 6820 114920 6880
rect 114980 6820 115030 6880
rect 115090 6820 115140 6880
rect 115200 6820 115250 6880
rect 115310 6820 115360 6880
rect 115420 6820 115430 6880
rect 114250 6800 115430 6820
rect 114250 6740 114260 6800
rect 114320 6740 114370 6800
rect 114430 6740 114480 6800
rect 114540 6740 114590 6800
rect 114650 6740 114700 6800
rect 114760 6740 114810 6800
rect 114870 6740 114920 6800
rect 114980 6740 115030 6800
rect 115090 6740 115140 6800
rect 115200 6740 115250 6800
rect 115310 6740 115360 6800
rect 115420 6740 115430 6800
rect 114250 6730 115430 6740
rect 113540 6320 113620 6330
rect 113540 6260 113550 6320
rect 113610 6260 113620 6320
rect 113540 6240 113620 6260
rect 113540 6180 113550 6240
rect 113610 6180 113620 6240
rect 113540 6160 113620 6180
rect 113540 6100 113550 6160
rect 113610 6100 113620 6160
rect 113540 6090 113620 6100
rect 113760 6320 113840 6330
rect 113760 6260 113770 6320
rect 113830 6260 113840 6320
rect 113760 6240 113840 6260
rect 113760 6180 113770 6240
rect 113830 6180 113840 6240
rect 113760 6160 113840 6180
rect 113760 6100 113770 6160
rect 113830 6100 113840 6160
rect 113760 6090 113840 6100
rect 113980 6320 114060 6330
rect 113980 6260 113990 6320
rect 114050 6260 114060 6320
rect 113980 6240 114060 6260
rect 113980 6180 113990 6240
rect 114050 6180 114060 6240
rect 113980 6160 114060 6180
rect 113980 6100 113990 6160
rect 114050 6100 114060 6160
rect 113980 6090 114060 6100
rect 113270 5880 113280 5940
rect 113340 5880 113350 5940
rect 113270 5870 113350 5880
rect 113570 5940 113650 5950
rect 113570 5880 113580 5940
rect 113640 5880 113650 5940
rect 112232 5830 112298 5840
rect 112232 5770 112238 5830
rect 112292 5770 112298 5830
rect 112232 5760 112298 5770
rect 112342 5830 112408 5840
rect 112342 5770 112348 5830
rect 112402 5770 112408 5830
rect 112342 5760 112408 5770
rect 112452 5830 112518 5840
rect 112452 5770 112458 5830
rect 112512 5770 112518 5830
rect 112452 5760 112518 5770
rect 112562 5830 112628 5840
rect 112562 5770 112568 5830
rect 112622 5770 112628 5830
rect 112562 5760 112628 5770
rect 112672 5830 112738 5840
rect 112672 5770 112678 5830
rect 112732 5770 112738 5830
rect 112672 5760 112738 5770
rect 112782 5830 112848 5840
rect 112782 5770 112788 5830
rect 112842 5770 112848 5830
rect 112782 5760 112848 5770
rect 112892 5830 112958 5840
rect 112892 5770 112898 5830
rect 112952 5770 112958 5830
rect 112892 5760 112958 5770
rect 113002 5830 113068 5840
rect 113002 5770 113008 5830
rect 113062 5770 113068 5830
rect 113002 5760 113068 5770
rect 113112 5830 113178 5840
rect 113112 5770 113118 5830
rect 113172 5770 113178 5830
rect 113112 5760 113178 5770
rect 113222 5830 113288 5840
rect 113222 5770 113228 5830
rect 113282 5770 113288 5830
rect 113222 5760 113288 5770
rect 112060 5700 112130 5720
rect 112060 5460 112080 5700
rect 112120 5460 112130 5700
rect 112060 5440 112130 5460
rect 112070 5430 112130 5440
rect 112180 5700 112240 5730
rect 112180 5460 112190 5700
rect 112230 5460 112240 5700
rect 112070 5380 112130 5400
rect 112070 5340 112080 5380
rect 112120 5340 112130 5380
rect 112070 5210 112130 5340
rect 112180 5320 112240 5460
rect 112290 5700 112350 5730
rect 112290 5460 112300 5700
rect 112340 5460 112350 5700
rect 112290 5430 112350 5460
rect 112400 5700 112460 5730
rect 112400 5460 112410 5700
rect 112450 5460 112460 5700
rect 112280 5420 112360 5430
rect 112280 5360 112290 5420
rect 112350 5360 112360 5420
rect 112280 5350 112360 5360
rect 112170 5310 112250 5320
rect 112170 5250 112180 5310
rect 112240 5250 112250 5310
rect 112170 5240 112250 5250
rect 112060 5200 112140 5210
rect 112060 5140 112070 5200
rect 112130 5140 112140 5200
rect 112060 5120 112140 5140
rect 112060 5060 112070 5120
rect 112130 5060 112140 5120
rect 112060 5040 112140 5060
rect 112060 4980 112070 5040
rect 112130 4980 112140 5040
rect 112060 4970 112140 4980
rect 112290 4050 112350 5350
rect 112400 5320 112460 5460
rect 112510 5700 112570 5730
rect 112510 5460 112520 5700
rect 112560 5460 112570 5700
rect 112510 5430 112570 5460
rect 112620 5700 112680 5730
rect 112620 5460 112630 5700
rect 112670 5460 112680 5700
rect 112500 5420 112580 5430
rect 112500 5360 112510 5420
rect 112570 5360 112580 5420
rect 112500 5350 112580 5360
rect 112390 5310 112470 5320
rect 112390 5250 112400 5310
rect 112460 5250 112470 5310
rect 112390 5240 112470 5250
rect 112170 4030 112250 4040
rect 112080 4010 112140 4020
rect 112170 3970 112180 4030
rect 112240 3970 112250 4030
rect 112510 4050 112570 5350
rect 112620 5320 112680 5460
rect 112730 5700 112790 5730
rect 112730 5460 112740 5700
rect 112780 5460 112790 5700
rect 112730 5430 112790 5460
rect 112840 5700 112900 5730
rect 112840 5460 112850 5700
rect 112890 5460 112900 5700
rect 112720 5420 112800 5430
rect 112720 5360 112730 5420
rect 112790 5360 112800 5420
rect 112720 5350 112800 5360
rect 112610 5310 112690 5320
rect 112610 5250 112620 5310
rect 112680 5250 112690 5310
rect 112610 5240 112690 5250
rect 112290 3980 112350 3990
rect 112390 4030 112470 4040
rect 112170 3960 112250 3970
rect 112390 3970 112400 4030
rect 112460 3970 112470 4030
rect 112730 4050 112790 5350
rect 112840 5320 112900 5460
rect 112950 5700 113010 5730
rect 112950 5460 112960 5700
rect 113000 5460 113010 5700
rect 112950 5430 113010 5460
rect 113060 5700 113120 5730
rect 113060 5460 113070 5700
rect 113110 5460 113120 5700
rect 112940 5420 113020 5430
rect 112940 5360 112950 5420
rect 113010 5360 113020 5420
rect 112940 5350 113020 5360
rect 112830 5310 112910 5320
rect 112830 5250 112840 5310
rect 112900 5250 112910 5310
rect 112830 5240 112910 5250
rect 112510 3980 112570 3990
rect 112610 4030 112690 4040
rect 112390 3960 112470 3970
rect 112610 3970 112620 4030
rect 112680 3970 112690 4030
rect 112950 4050 113010 5350
rect 113060 5320 113120 5460
rect 113170 5700 113230 5730
rect 113170 5460 113180 5700
rect 113220 5460 113230 5700
rect 113170 5430 113230 5460
rect 113280 5700 113340 5730
rect 113280 5460 113290 5700
rect 113330 5460 113340 5700
rect 113160 5420 113240 5430
rect 113160 5360 113170 5420
rect 113230 5360 113240 5420
rect 113160 5350 113240 5360
rect 113050 5310 113130 5320
rect 113050 5250 113060 5310
rect 113120 5250 113130 5310
rect 113050 5240 113130 5250
rect 112730 3980 112790 3990
rect 112830 4030 112910 4040
rect 112610 3960 112690 3970
rect 112830 3970 112840 4030
rect 112900 3970 112910 4030
rect 113170 4050 113230 5350
rect 113280 5320 113340 5460
rect 113390 5700 113530 5720
rect 113390 5460 113400 5700
rect 113440 5460 113530 5700
rect 113390 5440 113530 5460
rect 113390 5380 113450 5440
rect 113390 5340 113400 5380
rect 113440 5340 113450 5380
rect 113270 5310 113350 5320
rect 113270 5250 113280 5310
rect 113340 5250 113350 5310
rect 113270 5240 113350 5250
rect 113390 5210 113450 5340
rect 113570 5310 113650 5880
rect 113570 5250 113580 5310
rect 113640 5250 113650 5310
rect 113570 5240 113650 5250
rect 113950 5940 114030 5950
rect 113950 5880 113960 5940
rect 114020 5880 114030 5940
rect 113950 5310 114030 5880
rect 114250 5940 114330 6730
rect 114250 5880 114260 5940
rect 114320 5880 114330 5940
rect 114250 5870 114330 5880
rect 114470 5940 114550 6730
rect 114470 5880 114480 5940
rect 114540 5880 114550 5940
rect 114470 5870 114550 5880
rect 114690 5940 114770 6730
rect 114690 5880 114700 5940
rect 114760 5880 114770 5940
rect 114690 5870 114770 5880
rect 114910 5940 114990 6730
rect 114910 5880 114920 5940
rect 114980 5880 114990 5940
rect 114910 5870 114990 5880
rect 115130 5940 115210 6730
rect 115130 5880 115140 5940
rect 115200 5880 115210 5940
rect 115130 5870 115210 5880
rect 115350 5940 115430 6730
rect 115350 5880 115360 5940
rect 115420 5880 115430 5940
rect 115350 5870 115430 5880
rect 114312 5830 114378 5840
rect 114312 5770 114318 5830
rect 114372 5770 114378 5830
rect 114312 5760 114378 5770
rect 114422 5830 114488 5840
rect 114422 5770 114428 5830
rect 114482 5770 114488 5830
rect 114422 5760 114488 5770
rect 114532 5830 114598 5840
rect 114532 5770 114538 5830
rect 114592 5770 114598 5830
rect 114532 5760 114598 5770
rect 114642 5830 114708 5840
rect 114642 5770 114648 5830
rect 114702 5770 114708 5830
rect 114642 5760 114708 5770
rect 114752 5830 114818 5840
rect 114752 5770 114758 5830
rect 114812 5770 114818 5830
rect 114752 5760 114818 5770
rect 114862 5830 114928 5840
rect 114862 5770 114868 5830
rect 114922 5770 114928 5830
rect 114862 5760 114928 5770
rect 114972 5830 115038 5840
rect 114972 5770 114978 5830
rect 115032 5770 115038 5830
rect 114972 5760 115038 5770
rect 115082 5830 115148 5840
rect 115082 5770 115088 5830
rect 115142 5770 115148 5830
rect 115082 5760 115148 5770
rect 115192 5830 115258 5840
rect 115192 5770 115198 5830
rect 115252 5770 115258 5830
rect 115192 5760 115258 5770
rect 115302 5830 115368 5840
rect 115302 5770 115308 5830
rect 115362 5770 115368 5830
rect 115302 5760 115368 5770
rect 114070 5700 114210 5720
rect 114070 5460 114160 5700
rect 114200 5460 114210 5700
rect 114070 5440 114210 5460
rect 113950 5250 113960 5310
rect 114020 5250 114030 5310
rect 113950 5240 114030 5250
rect 114150 5380 114210 5440
rect 114150 5340 114160 5380
rect 114200 5340 114210 5380
rect 114150 5210 114210 5340
rect 114260 5700 114320 5730
rect 114260 5460 114270 5700
rect 114310 5460 114320 5700
rect 114260 5320 114320 5460
rect 114370 5700 114430 5730
rect 114370 5460 114380 5700
rect 114420 5460 114430 5700
rect 114370 5430 114430 5460
rect 114480 5700 114540 5730
rect 114480 5460 114490 5700
rect 114530 5460 114540 5700
rect 114360 5420 114440 5430
rect 114360 5360 114370 5420
rect 114430 5360 114440 5420
rect 114360 5350 114440 5360
rect 114250 5310 114330 5320
rect 114250 5250 114260 5310
rect 114320 5250 114330 5310
rect 114250 5240 114330 5250
rect 113380 5200 113460 5210
rect 113380 5140 113390 5200
rect 113450 5140 113460 5200
rect 113380 5120 113460 5140
rect 113380 5060 113390 5120
rect 113450 5060 113460 5120
rect 113380 5040 113460 5060
rect 113380 4980 113390 5040
rect 113450 4980 113460 5040
rect 113380 4970 113460 4980
rect 114140 5200 114220 5210
rect 114140 5140 114150 5200
rect 114210 5140 114220 5200
rect 114140 5120 114220 5140
rect 114140 5060 114150 5120
rect 114210 5060 114220 5120
rect 114140 5040 114220 5060
rect 114140 4980 114150 5040
rect 114210 4980 114220 5040
rect 114140 4970 114220 4980
rect 113760 4390 113840 4400
rect 113760 4330 113770 4390
rect 113830 4330 113840 4390
rect 113760 4310 113840 4330
rect 113760 4250 113770 4310
rect 113830 4250 113840 4310
rect 113760 4230 113840 4250
rect 113760 4170 113770 4230
rect 113830 4170 113840 4230
rect 113760 4160 113840 4170
rect 112950 3980 113010 3990
rect 113050 4030 113130 4040
rect 112830 3960 112910 3970
rect 113050 3970 113060 4030
rect 113120 3970 113130 4030
rect 113170 3980 113230 3990
rect 113270 4030 113350 4040
rect 113050 3960 113130 3970
rect 113270 3970 113280 4030
rect 113340 3970 113350 4030
rect 113270 3960 113350 3970
rect 113380 4030 113440 4040
rect 113380 3960 113440 3970
rect 113680 4030 113740 4040
rect 113680 3960 113740 3970
rect 112080 3940 112140 3950
rect 112070 3830 112130 3850
rect 112070 3590 112080 3830
rect 112120 3590 112130 3830
rect 112070 3570 112130 3590
rect 112180 3830 112240 3960
rect 112280 3940 112360 3950
rect 112280 3880 112290 3940
rect 112350 3880 112360 3940
rect 112280 3870 112360 3880
rect 112180 3590 112190 3830
rect 112230 3590 112240 3830
rect 112180 3560 112240 3590
rect 112290 3830 112350 3870
rect 112290 3590 112300 3830
rect 112340 3590 112350 3830
rect 112170 3550 112250 3560
rect 112070 3510 112130 3530
rect 112070 3470 112080 3510
rect 112120 3470 112130 3510
rect 112170 3490 112180 3550
rect 112240 3490 112250 3550
rect 112170 3480 112250 3490
rect 112070 3450 112130 3470
rect 112080 2510 112120 3450
rect 112290 3420 112350 3590
rect 112400 3830 112460 3960
rect 112500 3940 112580 3950
rect 112500 3880 112510 3940
rect 112570 3880 112580 3940
rect 112500 3870 112580 3880
rect 112400 3590 112410 3830
rect 112450 3590 112460 3830
rect 112400 3560 112460 3590
rect 112510 3830 112570 3870
rect 112510 3590 112520 3830
rect 112560 3590 112570 3830
rect 112390 3550 112470 3560
rect 112390 3490 112400 3550
rect 112460 3490 112470 3550
rect 112390 3480 112470 3490
rect 112510 3420 112570 3590
rect 112620 3830 112680 3960
rect 112720 3940 112800 3950
rect 112720 3880 112730 3940
rect 112790 3880 112800 3940
rect 112720 3870 112800 3880
rect 112620 3590 112630 3830
rect 112670 3590 112680 3830
rect 112620 3560 112680 3590
rect 112730 3830 112790 3870
rect 112730 3590 112740 3830
rect 112780 3590 112790 3830
rect 112610 3550 112690 3560
rect 112610 3490 112620 3550
rect 112680 3490 112690 3550
rect 112610 3480 112690 3490
rect 112730 3420 112790 3590
rect 112840 3830 112900 3960
rect 112940 3940 113020 3950
rect 112940 3880 112950 3940
rect 113010 3880 113020 3940
rect 112940 3870 113020 3880
rect 112840 3590 112850 3830
rect 112890 3590 112900 3830
rect 112840 3560 112900 3590
rect 112950 3830 113010 3870
rect 112950 3590 112960 3830
rect 113000 3590 113010 3830
rect 112830 3550 112910 3560
rect 112830 3490 112840 3550
rect 112900 3490 112910 3550
rect 112830 3480 112910 3490
rect 112950 3420 113010 3590
rect 113060 3830 113120 3960
rect 113160 3940 113240 3950
rect 113160 3880 113170 3940
rect 113230 3880 113240 3940
rect 113160 3870 113240 3880
rect 113060 3590 113070 3830
rect 113110 3590 113120 3830
rect 113060 3560 113120 3590
rect 113170 3830 113230 3870
rect 113170 3590 113180 3830
rect 113220 3590 113230 3830
rect 113050 3550 113130 3560
rect 113050 3490 113060 3550
rect 113120 3490 113130 3550
rect 113050 3480 113130 3490
rect 113170 3420 113230 3590
rect 113280 3830 113340 3960
rect 113280 3590 113290 3830
rect 113330 3590 113340 3830
rect 113280 3560 113340 3590
rect 113390 3830 113610 3850
rect 113390 3590 113400 3830
rect 113440 3590 113560 3830
rect 113600 3590 113610 3830
rect 113390 3570 113610 3590
rect 113660 3830 113720 3850
rect 113660 3590 113670 3830
rect 113710 3590 113720 3830
rect 113270 3550 113350 3560
rect 113270 3490 113280 3550
rect 113340 3490 113350 3550
rect 113480 3530 113520 3570
rect 113660 3560 113720 3590
rect 113770 3830 113830 4160
rect 114370 4050 114430 5350
rect 114480 5320 114540 5460
rect 114590 5700 114650 5730
rect 114590 5460 114600 5700
rect 114640 5460 114650 5700
rect 114590 5430 114650 5460
rect 114700 5700 114760 5730
rect 114700 5460 114710 5700
rect 114750 5460 114760 5700
rect 114580 5420 114660 5430
rect 114580 5360 114590 5420
rect 114650 5360 114660 5420
rect 114580 5350 114660 5360
rect 114470 5310 114550 5320
rect 114470 5250 114480 5310
rect 114540 5250 114550 5310
rect 114470 5240 114550 5250
rect 113860 4030 113920 4040
rect 113860 3960 113920 3970
rect 114160 4030 114220 4040
rect 114160 3960 114220 3970
rect 114250 4030 114330 4040
rect 114250 3970 114260 4030
rect 114320 3970 114330 4030
rect 114590 4050 114650 5350
rect 114700 5320 114760 5460
rect 114810 5700 114870 5730
rect 114810 5460 114820 5700
rect 114860 5460 114870 5700
rect 114810 5430 114870 5460
rect 114920 5700 114980 5730
rect 114920 5460 114930 5700
rect 114970 5460 114980 5700
rect 114800 5420 114880 5430
rect 114800 5360 114810 5420
rect 114870 5360 114880 5420
rect 114800 5350 114880 5360
rect 114690 5310 114770 5320
rect 114690 5250 114700 5310
rect 114760 5250 114770 5310
rect 114690 5240 114770 5250
rect 114370 3980 114430 3990
rect 114470 4030 114550 4040
rect 114250 3960 114330 3970
rect 114470 3970 114480 4030
rect 114540 3970 114550 4030
rect 114810 4050 114870 5350
rect 114920 5320 114980 5460
rect 115030 5700 115090 5730
rect 115030 5460 115040 5700
rect 115080 5460 115090 5700
rect 115030 5430 115090 5460
rect 115140 5700 115200 5730
rect 115140 5460 115150 5700
rect 115190 5460 115200 5700
rect 115020 5420 115100 5430
rect 115020 5360 115030 5420
rect 115090 5360 115100 5420
rect 115020 5350 115100 5360
rect 114910 5310 114990 5320
rect 114910 5250 114920 5310
rect 114980 5250 114990 5310
rect 114910 5240 114990 5250
rect 114590 3980 114650 3990
rect 114690 4030 114770 4040
rect 114470 3960 114550 3970
rect 114690 3970 114700 4030
rect 114760 3970 114770 4030
rect 115030 4050 115090 5350
rect 115140 5320 115200 5460
rect 115250 5700 115310 5730
rect 115250 5460 115260 5700
rect 115300 5460 115310 5700
rect 115250 5430 115310 5460
rect 115360 5700 115420 5730
rect 115360 5460 115370 5700
rect 115410 5460 115420 5700
rect 115240 5420 115320 5430
rect 115240 5360 115250 5420
rect 115310 5360 115320 5420
rect 115240 5350 115320 5360
rect 115130 5310 115210 5320
rect 115130 5250 115140 5310
rect 115200 5250 115210 5310
rect 115130 5240 115210 5250
rect 114810 3980 114870 3990
rect 114910 4030 114990 4040
rect 114690 3960 114770 3970
rect 114910 3970 114920 4030
rect 114980 3970 114990 4030
rect 115250 4050 115310 5350
rect 115360 5320 115420 5460
rect 115470 5700 115530 5720
rect 115470 5460 115480 5700
rect 115520 5460 115530 5700
rect 115470 5440 115530 5460
rect 115470 5380 115530 5400
rect 115470 5340 115480 5380
rect 115520 5340 115530 5380
rect 115350 5310 115430 5320
rect 115350 5250 115360 5310
rect 115420 5250 115430 5310
rect 115350 5240 115430 5250
rect 115470 5210 115530 5340
rect 115460 5200 115540 5210
rect 115460 5140 115470 5200
rect 115530 5140 115540 5200
rect 115460 5120 115540 5140
rect 115460 5060 115470 5120
rect 115530 5060 115540 5120
rect 115460 5040 115540 5060
rect 115460 4980 115470 5040
rect 115530 4980 115540 5040
rect 115460 4970 115540 4980
rect 115030 3980 115090 3990
rect 115130 4030 115210 4040
rect 114910 3960 114990 3970
rect 115130 3970 115140 4030
rect 115200 3970 115210 4030
rect 115250 3980 115310 3990
rect 115350 4030 115430 4040
rect 115130 3960 115210 3970
rect 115350 3970 115360 4030
rect 115420 3970 115430 4030
rect 115350 3960 115430 3970
rect 115460 4010 115520 4020
rect 113770 3590 113780 3830
rect 113820 3590 113830 3830
rect 113770 3570 113830 3590
rect 113880 3830 113940 3850
rect 113880 3590 113890 3830
rect 113930 3590 113940 3830
rect 113880 3560 113940 3590
rect 113990 3830 114210 3850
rect 113990 3590 114000 3830
rect 114040 3590 114160 3830
rect 114200 3590 114210 3830
rect 113990 3570 114210 3590
rect 114260 3830 114320 3960
rect 114360 3940 114440 3950
rect 114360 3880 114370 3940
rect 114430 3880 114440 3940
rect 114360 3870 114440 3880
rect 114260 3590 114270 3830
rect 114310 3590 114320 3830
rect 113650 3550 113730 3560
rect 113270 3480 113350 3490
rect 113470 3510 113530 3530
rect 113470 3470 113480 3510
rect 113520 3470 113530 3510
rect 113470 3450 113530 3470
rect 113650 3490 113660 3550
rect 113720 3490 113730 3550
rect 112280 3410 112360 3420
rect 112280 3350 112290 3410
rect 112350 3350 112360 3410
rect 112280 3340 112360 3350
rect 112500 3410 112580 3420
rect 112500 3350 112510 3410
rect 112570 3350 112580 3410
rect 112500 3340 112580 3350
rect 112720 3410 112800 3420
rect 112720 3350 112730 3410
rect 112790 3350 112800 3410
rect 112720 3340 112800 3350
rect 112880 3410 113400 3420
rect 112880 3350 112950 3410
rect 113010 3350 113170 3410
rect 113230 3350 113400 3410
rect 112060 2500 112140 2510
rect 112060 2440 112070 2500
rect 112130 2440 112140 2500
rect 112060 2420 112140 2440
rect 112060 2360 112070 2420
rect 112130 2360 112140 2420
rect 112060 2340 112140 2360
rect 112060 2280 112070 2340
rect 112130 2280 112140 2340
rect 112060 2270 112140 2280
rect 111880 2230 111960 2240
rect 111880 2170 111890 2230
rect 111950 2170 111960 2230
rect 111880 2160 111960 2170
rect 112880 1730 113400 3350
rect 113480 2510 113520 3450
rect 113460 2500 113540 2510
rect 113460 2440 113470 2500
rect 113530 2440 113540 2500
rect 113460 2420 113540 2440
rect 113460 2360 113470 2420
rect 113530 2360 113540 2420
rect 113460 2340 113540 2360
rect 113460 2280 113470 2340
rect 113530 2280 113540 2340
rect 113460 2270 113540 2280
rect 112880 1670 112890 1730
rect 112950 1670 113110 1730
rect 113170 1670 113330 1730
rect 113390 1670 113400 1730
rect 112880 1660 113400 1670
rect 113540 1730 113620 1740
rect 113540 1670 113550 1730
rect 113610 1670 113620 1730
rect 113540 1660 113620 1670
rect 113650 1700 113730 3490
rect 113870 3550 113950 3560
rect 113870 3490 113880 3550
rect 113940 3490 113950 3550
rect 114080 3530 114120 3570
rect 114260 3560 114320 3590
rect 114370 3830 114430 3870
rect 114370 3590 114380 3830
rect 114420 3590 114430 3830
rect 114250 3550 114330 3560
rect 113650 1660 113670 1700
rect 113710 1660 113730 1700
rect 113760 1730 113840 1740
rect 113760 1670 113770 1730
rect 113830 1670 113840 1730
rect 113760 1660 113840 1670
rect 113870 1700 113950 3490
rect 114070 3510 114130 3530
rect 114070 3470 114080 3510
rect 114120 3470 114130 3510
rect 114250 3490 114260 3550
rect 114320 3490 114330 3550
rect 114250 3480 114330 3490
rect 114070 3450 114130 3470
rect 114080 2510 114120 3450
rect 114370 3420 114430 3590
rect 114480 3830 114540 3960
rect 114580 3940 114660 3950
rect 114580 3880 114590 3940
rect 114650 3880 114660 3940
rect 114580 3870 114660 3880
rect 114480 3590 114490 3830
rect 114530 3590 114540 3830
rect 114480 3560 114540 3590
rect 114590 3830 114650 3870
rect 114590 3590 114600 3830
rect 114640 3590 114650 3830
rect 114470 3550 114550 3560
rect 114470 3490 114480 3550
rect 114540 3490 114550 3550
rect 114470 3480 114550 3490
rect 114590 3420 114650 3590
rect 114700 3830 114760 3960
rect 114800 3940 114880 3950
rect 114800 3880 114810 3940
rect 114870 3880 114880 3940
rect 114800 3870 114880 3880
rect 114700 3590 114710 3830
rect 114750 3590 114760 3830
rect 114700 3560 114760 3590
rect 114810 3830 114870 3870
rect 114810 3590 114820 3830
rect 114860 3590 114870 3830
rect 114690 3550 114770 3560
rect 114690 3490 114700 3550
rect 114760 3490 114770 3550
rect 114690 3480 114770 3490
rect 114810 3420 114870 3590
rect 114920 3830 114980 3960
rect 115020 3940 115100 3950
rect 115020 3880 115030 3940
rect 115090 3880 115100 3940
rect 115020 3870 115100 3880
rect 114920 3590 114930 3830
rect 114970 3590 114980 3830
rect 114920 3560 114980 3590
rect 115030 3830 115090 3870
rect 115030 3590 115040 3830
rect 115080 3590 115090 3830
rect 114910 3550 114990 3560
rect 114910 3490 114920 3550
rect 114980 3490 114990 3550
rect 114910 3480 114990 3490
rect 115030 3420 115090 3590
rect 115140 3830 115200 3960
rect 115240 3940 115320 3950
rect 115240 3880 115250 3940
rect 115310 3880 115320 3940
rect 115240 3870 115320 3880
rect 115140 3590 115150 3830
rect 115190 3590 115200 3830
rect 115140 3560 115200 3590
rect 115250 3830 115310 3870
rect 115250 3590 115260 3830
rect 115300 3590 115310 3830
rect 115130 3550 115210 3560
rect 115130 3490 115140 3550
rect 115200 3490 115210 3550
rect 115130 3480 115210 3490
rect 115250 3420 115310 3590
rect 115360 3830 115420 3960
rect 115460 3940 115520 3950
rect 115360 3590 115370 3830
rect 115410 3590 115420 3830
rect 115360 3560 115420 3590
rect 115470 3830 115530 3850
rect 115470 3590 115480 3830
rect 115520 3590 115530 3830
rect 115470 3570 115530 3590
rect 115350 3550 115430 3560
rect 115350 3490 115360 3550
rect 115420 3490 115430 3550
rect 115350 3480 115430 3490
rect 115470 3510 115530 3530
rect 115470 3470 115480 3510
rect 115520 3470 115530 3510
rect 115470 3450 115530 3470
rect 114200 3410 114720 3420
rect 114200 3350 114370 3410
rect 114430 3350 114590 3410
rect 114650 3350 114720 3410
rect 114060 2500 114140 2510
rect 114060 2440 114070 2500
rect 114130 2440 114140 2500
rect 114060 2420 114140 2440
rect 114060 2360 114070 2420
rect 114130 2360 114140 2420
rect 114060 2340 114140 2360
rect 114060 2280 114070 2340
rect 114130 2280 114140 2340
rect 114060 2270 114140 2280
rect 113870 1660 113890 1700
rect 113930 1660 113950 1700
rect 113980 1730 114060 1740
rect 113980 1670 113990 1730
rect 114050 1670 114060 1730
rect 113980 1660 114060 1670
rect 114200 1730 114720 3350
rect 114800 3410 114880 3420
rect 114800 3350 114810 3410
rect 114870 3350 114880 3410
rect 114800 3340 114880 3350
rect 115020 3410 115100 3420
rect 115020 3350 115030 3410
rect 115090 3350 115100 3410
rect 115020 3340 115100 3350
rect 115240 3410 115320 3420
rect 115240 3350 115250 3410
rect 115310 3350 115320 3410
rect 115240 3340 115320 3350
rect 115480 2510 115520 3450
rect 115460 2500 115540 2510
rect 115460 2440 115470 2500
rect 115530 2440 115540 2500
rect 115460 2420 115540 2440
rect 115460 2360 115470 2420
rect 115530 2360 115540 2420
rect 115460 2340 115540 2360
rect 115460 2280 115470 2340
rect 115530 2280 115540 2340
rect 115460 2270 115540 2280
rect 115650 2240 115690 7220
rect 116290 7210 116300 7270
rect 116360 7210 116380 7270
rect 116440 7210 116460 7270
rect 116520 7210 116530 7270
rect 116290 7190 116530 7210
rect 116290 7130 116300 7190
rect 116360 7130 116380 7190
rect 116440 7130 116460 7190
rect 116520 7130 116530 7190
rect 115720 7070 115800 7080
rect 115720 7010 115730 7070
rect 115790 7010 115800 7070
rect 115720 7000 115800 7010
rect 115630 2230 115710 2240
rect 115630 2170 115640 2230
rect 115700 2170 115710 2230
rect 115630 2160 115710 2170
rect 114200 1670 114210 1730
rect 114270 1670 114430 1730
rect 114490 1670 114650 1730
rect 114710 1670 114720 1730
rect 114200 1660 114720 1670
rect 114860 1730 114940 1740
rect 114860 1670 114870 1730
rect 114930 1670 114940 1730
rect 114860 1660 114940 1670
rect 112370 1580 112510 1600
rect 112370 1140 112460 1580
rect 112500 1140 112510 1580
rect 112370 1120 112510 1140
rect 112450 1080 112510 1120
rect 112560 1580 112620 1600
rect 112560 1140 112570 1580
rect 112610 1140 112620 1580
rect 112560 1080 112620 1140
rect 112670 1580 112730 1600
rect 112670 1140 112680 1580
rect 112720 1140 112730 1580
rect 111690 140 111700 200
rect 111760 140 111770 200
rect 111690 130 111770 140
rect 112440 1070 112520 1080
rect 112440 1010 112450 1070
rect 112510 1010 112520 1070
rect 110300 -30 110380 -20
rect 110300 -90 110310 -30
rect 110370 -90 110380 -30
rect 110300 -100 110380 -90
rect 110510 -70 110570 10
rect 110510 -110 110520 -70
rect 110560 -110 110570 -70
rect 110510 -1150 110570 -110
rect 112440 -240 112520 1010
rect 112550 1070 112630 1080
rect 112550 1010 112560 1070
rect 112620 1010 112630 1070
rect 112550 1000 112630 1010
rect 112670 590 112730 1140
rect 112780 1580 112840 1600
rect 112780 1140 112790 1580
rect 112830 1140 112840 1580
rect 112780 1080 112840 1140
rect 112890 1580 112950 1660
rect 112890 1140 112900 1580
rect 112940 1140 112950 1580
rect 112770 1070 112850 1080
rect 112770 1010 112780 1070
rect 112840 1010 112850 1070
rect 112770 1000 112850 1010
rect 112890 970 112950 1140
rect 113000 1580 113060 1600
rect 113000 1140 113010 1580
rect 113050 1140 113060 1580
rect 113000 1080 113060 1140
rect 113110 1580 113170 1660
rect 113110 1140 113120 1580
rect 113160 1140 113170 1580
rect 112990 1070 113070 1080
rect 112990 1010 113000 1070
rect 113060 1010 113070 1070
rect 112990 1000 113070 1010
rect 113110 970 113170 1140
rect 113220 1580 113280 1600
rect 113220 1140 113230 1580
rect 113270 1140 113280 1580
rect 113220 1080 113280 1140
rect 113330 1580 113390 1660
rect 113330 1140 113340 1580
rect 113380 1140 113390 1580
rect 113210 1070 113290 1080
rect 113210 1010 113220 1070
rect 113280 1010 113290 1070
rect 113210 1000 113290 1010
rect 113330 970 113390 1140
rect 113440 1580 113500 1600
rect 113440 1140 113450 1580
rect 113490 1140 113500 1580
rect 113440 1080 113500 1140
rect 113550 1580 113610 1660
rect 113650 1640 113730 1660
rect 113550 1140 113560 1580
rect 113600 1140 113610 1580
rect 113430 1070 113510 1080
rect 113430 1010 113440 1070
rect 113500 1010 113510 1070
rect 113430 1000 113510 1010
rect 113550 970 113610 1140
rect 113660 1580 113720 1600
rect 113660 1140 113670 1580
rect 113710 1140 113720 1580
rect 113660 1080 113720 1140
rect 113770 1580 113830 1660
rect 113870 1640 113950 1660
rect 113770 1140 113780 1580
rect 113820 1140 113830 1580
rect 113650 1070 113730 1080
rect 113650 1010 113660 1070
rect 113720 1010 113730 1070
rect 113650 1000 113730 1010
rect 113770 970 113830 1140
rect 113880 1580 113940 1600
rect 113880 1140 113890 1580
rect 113930 1140 113940 1580
rect 113880 1080 113940 1140
rect 113990 1580 114050 1660
rect 113990 1140 114000 1580
rect 114040 1140 114050 1580
rect 113870 1070 113950 1080
rect 113870 1010 113880 1070
rect 113940 1010 113950 1070
rect 113870 1000 113950 1010
rect 113990 970 114050 1140
rect 114100 1580 114160 1600
rect 114100 1140 114110 1580
rect 114150 1140 114160 1580
rect 114100 1080 114160 1140
rect 114210 1580 114270 1660
rect 114210 1140 114220 1580
rect 114260 1140 114270 1580
rect 114090 1070 114170 1080
rect 114090 1010 114100 1070
rect 114160 1010 114170 1070
rect 114090 1000 114170 1010
rect 114210 970 114270 1140
rect 114320 1580 114380 1600
rect 114320 1140 114330 1580
rect 114370 1140 114380 1580
rect 114320 1080 114380 1140
rect 114430 1580 114490 1660
rect 114430 1140 114440 1580
rect 114480 1140 114490 1580
rect 114310 1070 114390 1080
rect 114310 1010 114320 1070
rect 114380 1010 114390 1070
rect 114310 1000 114390 1010
rect 114430 970 114490 1140
rect 114540 1580 114600 1600
rect 114540 1140 114550 1580
rect 114590 1140 114600 1580
rect 114540 1080 114600 1140
rect 114650 1580 114710 1660
rect 114650 1140 114660 1580
rect 114700 1140 114710 1580
rect 114530 1070 114610 1080
rect 114530 1010 114540 1070
rect 114600 1010 114610 1070
rect 114530 1000 114610 1010
rect 114650 970 114710 1140
rect 114760 1580 114820 1600
rect 114760 1140 114770 1580
rect 114810 1140 114820 1580
rect 114760 1080 114820 1140
rect 114870 1580 114930 1660
rect 114870 1140 114880 1580
rect 114920 1140 114930 1580
rect 114750 1070 114830 1080
rect 114750 1010 114760 1070
rect 114820 1010 114830 1070
rect 114750 1000 114830 1010
rect 114870 970 114930 1140
rect 114980 1580 115040 1600
rect 114980 1140 114990 1580
rect 115030 1140 115040 1580
rect 114980 1080 115040 1140
rect 114970 1070 115050 1080
rect 114970 1010 114980 1070
rect 115040 1010 115050 1070
rect 112880 960 112960 970
rect 112880 900 112890 960
rect 112950 900 112960 960
rect 112880 880 112960 900
rect 112880 820 112890 880
rect 112950 820 112960 880
rect 112880 800 112960 820
rect 112880 740 112890 800
rect 112950 740 112960 800
rect 112880 730 112960 740
rect 113100 960 113180 970
rect 113100 900 113110 960
rect 113170 900 113180 960
rect 113100 880 113180 900
rect 113100 820 113110 880
rect 113170 820 113180 880
rect 113100 800 113180 820
rect 113100 740 113110 800
rect 113170 740 113180 800
rect 113100 730 113180 740
rect 113320 960 113400 970
rect 113320 900 113330 960
rect 113390 900 113400 960
rect 113320 880 113400 900
rect 113320 820 113330 880
rect 113390 820 113400 880
rect 113320 800 113400 820
rect 113320 740 113330 800
rect 113390 740 113400 800
rect 113320 730 113400 740
rect 113540 960 113620 970
rect 113540 900 113550 960
rect 113610 900 113620 960
rect 113540 880 113620 900
rect 113540 820 113550 880
rect 113610 820 113620 880
rect 113540 800 113620 820
rect 113540 740 113550 800
rect 113610 740 113620 800
rect 113540 730 113620 740
rect 113760 960 113840 970
rect 113760 900 113770 960
rect 113830 900 113840 960
rect 113760 880 113840 900
rect 113760 820 113770 880
rect 113830 820 113840 880
rect 113760 800 113840 820
rect 113760 740 113770 800
rect 113830 740 113840 800
rect 113760 730 113840 740
rect 113980 960 114060 970
rect 113980 900 113990 960
rect 114050 900 114060 960
rect 113980 880 114060 900
rect 113980 820 113990 880
rect 114050 820 114060 880
rect 113980 800 114060 820
rect 113980 740 113990 800
rect 114050 740 114060 800
rect 113980 730 114060 740
rect 114200 960 114280 970
rect 114200 900 114210 960
rect 114270 900 114280 960
rect 114200 880 114280 900
rect 114200 820 114210 880
rect 114270 820 114280 880
rect 114200 800 114280 820
rect 114200 740 114210 800
rect 114270 740 114280 800
rect 114200 730 114280 740
rect 114420 960 114500 970
rect 114420 900 114430 960
rect 114490 900 114500 960
rect 114420 880 114500 900
rect 114420 820 114430 880
rect 114490 820 114500 880
rect 114420 800 114500 820
rect 114420 740 114430 800
rect 114490 740 114500 800
rect 114420 730 114500 740
rect 114640 960 114720 970
rect 114640 900 114650 960
rect 114710 900 114720 960
rect 114640 880 114720 900
rect 114640 820 114650 880
rect 114710 820 114720 880
rect 114640 800 114720 820
rect 114640 740 114650 800
rect 114710 740 114720 800
rect 114640 730 114720 740
rect 114860 960 114940 970
rect 114860 900 114870 960
rect 114930 900 114940 960
rect 114860 880 114940 900
rect 114860 820 114870 880
rect 114930 820 114940 880
rect 114860 800 114940 820
rect 114860 740 114870 800
rect 114930 740 114940 800
rect 114860 730 114940 740
rect 114830 690 114910 700
rect 114830 630 114840 690
rect 114900 630 114910 690
rect 114830 620 114910 630
rect 112660 580 112740 590
rect 112660 520 112670 580
rect 112730 520 112740 580
rect 112660 500 112740 520
rect 112660 440 112670 500
rect 112730 440 112740 500
rect 112660 420 112740 440
rect 112660 360 112670 420
rect 112730 360 112740 420
rect 112660 350 112740 360
rect 112440 -300 112450 -240
rect 112510 -300 112520 -240
rect 112440 -1150 112520 -300
rect 113240 310 113320 320
rect 113240 250 113250 310
rect 113310 250 113320 310
rect 113240 -460 113320 250
rect 113650 310 113730 320
rect 113650 250 113660 310
rect 113720 250 113730 310
rect 113650 240 113730 250
rect 113870 310 113950 320
rect 113870 250 113880 310
rect 113940 250 113950 310
rect 113870 240 113950 250
rect 113540 200 113620 210
rect 113540 140 113550 200
rect 113610 140 113620 200
rect 113540 130 113620 140
rect 113360 70 113500 90
rect 113360 -170 113450 70
rect 113490 -170 113500 70
rect 113360 -190 113500 -170
rect 113440 -250 113500 -190
rect 113550 70 113610 130
rect 113550 -170 113560 70
rect 113600 -170 113610 70
rect 113550 -230 113610 -170
rect 113660 70 113720 240
rect 113760 200 113840 210
rect 113760 140 113770 200
rect 113830 140 113840 200
rect 113760 130 113840 140
rect 113660 -170 113670 70
rect 113710 -170 113720 70
rect 113660 -190 113720 -170
rect 113770 70 113830 130
rect 113770 -170 113780 70
rect 113820 -170 113830 70
rect 113770 -230 113830 -170
rect 113880 70 113940 240
rect 113980 200 114060 210
rect 113980 140 113990 200
rect 114050 140 114060 200
rect 113980 130 114060 140
rect 113880 -170 113890 70
rect 113930 -170 113940 70
rect 113880 -190 113940 -170
rect 113990 70 114050 130
rect 113990 -170 114000 70
rect 114040 -170 114050 70
rect 113990 -230 114050 -170
rect 114100 70 114240 90
rect 114100 -170 114110 70
rect 114150 -170 114240 70
rect 114100 -190 114240 -170
rect 113440 -290 113450 -250
rect 113490 -290 113500 -250
rect 113440 -310 113500 -290
rect 113540 -240 113620 -230
rect 113540 -300 113550 -240
rect 113610 -300 113620 -240
rect 113540 -310 113620 -300
rect 113760 -240 113840 -230
rect 113760 -300 113770 -240
rect 113830 -300 113840 -240
rect 113760 -320 113840 -300
rect 113980 -240 114060 -230
rect 113980 -300 113990 -240
rect 114050 -300 114060 -240
rect 113980 -310 114060 -300
rect 114100 -240 114160 -190
rect 114100 -310 114160 -300
rect 114970 -240 115050 1010
rect 114970 -300 114980 -240
rect 115040 -300 115050 -240
rect 113760 -380 113770 -320
rect 113830 -380 113840 -320
rect 113760 -390 113840 -380
rect 113240 -520 113250 -460
rect 113310 -520 113320 -460
rect 113240 -540 113320 -520
rect 113240 -600 113250 -540
rect 113310 -600 113320 -540
rect 113240 -620 113320 -600
rect 113240 -680 113250 -620
rect 113310 -680 113320 -620
rect 113240 -690 113320 -680
rect 113430 -450 113490 -430
rect 113430 -710 113490 -690
rect 114110 -450 114170 -430
rect 114110 -710 114170 -690
rect 110110 -1160 110420 -1150
rect 110110 -1220 110190 -1160
rect 110250 -1220 110270 -1160
rect 110330 -1220 110350 -1160
rect 110410 -1220 110420 -1160
rect 110110 -1240 110420 -1220
rect 110110 -1300 110190 -1240
rect 110250 -1300 110270 -1240
rect 110330 -1300 110350 -1240
rect 110410 -1300 110420 -1240
rect 110110 -1320 110420 -1300
rect 110110 -1380 110190 -1320
rect 110250 -1380 110270 -1320
rect 110330 -1380 110350 -1320
rect 110410 -1380 110420 -1320
rect 110110 -1390 110420 -1380
rect 110500 -1160 110580 -1150
rect 110500 -1220 110510 -1160
rect 110570 -1220 110580 -1160
rect 110500 -1240 110580 -1220
rect 110500 -1300 110510 -1240
rect 110570 -1300 110580 -1240
rect 110500 -1320 110580 -1300
rect 110500 -1380 110510 -1320
rect 110570 -1380 110580 -1320
rect 110500 -1390 110580 -1380
rect 110880 -1160 111120 -1150
rect 110880 -1220 110890 -1160
rect 110950 -1220 110970 -1160
rect 111030 -1220 111050 -1160
rect 111110 -1220 111120 -1160
rect 110880 -1240 111120 -1220
rect 110880 -1300 110890 -1240
rect 110950 -1300 110970 -1240
rect 111030 -1300 111050 -1240
rect 111110 -1300 111120 -1240
rect 110880 -1320 111120 -1300
rect 110880 -1380 110890 -1320
rect 110950 -1380 110970 -1320
rect 111030 -1380 111050 -1320
rect 111110 -1380 111120 -1320
rect 109480 -3000 109720 -1390
rect 110180 -3000 110420 -1390
rect 110880 -3000 111120 -1380
rect 111580 -1160 111820 -1150
rect 111580 -1220 111590 -1160
rect 111650 -1220 111670 -1160
rect 111730 -1220 111750 -1160
rect 111810 -1220 111820 -1160
rect 111580 -1240 111820 -1220
rect 111580 -1300 111590 -1240
rect 111650 -1300 111670 -1240
rect 111730 -1300 111750 -1240
rect 111810 -1300 111820 -1240
rect 111580 -1320 111820 -1300
rect 111580 -1380 111590 -1320
rect 111650 -1380 111670 -1320
rect 111730 -1380 111750 -1320
rect 111810 -1380 111820 -1320
rect 111580 -3000 111820 -1380
rect 112280 -1160 112520 -1150
rect 112280 -1220 112290 -1160
rect 112350 -1220 112370 -1160
rect 112430 -1220 112450 -1160
rect 112510 -1220 112520 -1160
rect 112280 -1240 112520 -1220
rect 112280 -1300 112290 -1240
rect 112350 -1300 112370 -1240
rect 112430 -1300 112450 -1240
rect 112510 -1300 112520 -1240
rect 112280 -1320 112520 -1300
rect 112280 -1380 112290 -1320
rect 112350 -1380 112370 -1320
rect 112430 -1380 112450 -1320
rect 112510 -1380 112520 -1320
rect 112280 -3000 112520 -1380
rect 112980 -1160 113220 -1150
rect 112980 -1220 112990 -1160
rect 113050 -1220 113070 -1160
rect 113130 -1220 113150 -1160
rect 113210 -1220 113220 -1160
rect 112980 -1240 113220 -1220
rect 112980 -1300 112990 -1240
rect 113050 -1300 113070 -1240
rect 113130 -1300 113150 -1240
rect 113210 -1300 113220 -1240
rect 112980 -1320 113220 -1300
rect 112980 -1380 112990 -1320
rect 113050 -1380 113070 -1320
rect 113130 -1380 113150 -1320
rect 113210 -1380 113220 -1320
rect 112980 -3000 113220 -1380
rect 113680 -1160 113920 -1150
rect 113680 -1220 113690 -1160
rect 113750 -1220 113770 -1160
rect 113830 -1220 113850 -1160
rect 113910 -1220 113920 -1160
rect 113680 -1240 113920 -1220
rect 113680 -1300 113690 -1240
rect 113750 -1300 113770 -1240
rect 113830 -1300 113850 -1240
rect 113910 -1300 113920 -1240
rect 113680 -1320 113920 -1300
rect 113680 -1380 113690 -1320
rect 113750 -1380 113770 -1320
rect 113830 -1380 113850 -1320
rect 113910 -1380 113920 -1320
rect 113680 -3000 113920 -1380
rect 114380 -1160 114620 -1150
rect 114380 -1220 114390 -1160
rect 114450 -1220 114470 -1160
rect 114530 -1220 114550 -1160
rect 114610 -1220 114620 -1160
rect 114380 -1240 114620 -1220
rect 114380 -1300 114390 -1240
rect 114450 -1300 114470 -1240
rect 114530 -1300 114550 -1240
rect 114610 -1300 114620 -1240
rect 114380 -1320 114620 -1300
rect 114380 -1380 114390 -1320
rect 114450 -1380 114470 -1320
rect 114530 -1380 114550 -1320
rect 114610 -1380 114620 -1320
rect 114380 -3000 114620 -1380
rect 114970 -1160 115050 -300
rect 115080 960 115320 970
rect 115080 900 115090 960
rect 115150 900 115170 960
rect 115230 900 115250 960
rect 115310 900 115320 960
rect 115080 880 115320 900
rect 115080 820 115090 880
rect 115150 820 115170 880
rect 115230 820 115250 880
rect 115310 820 115320 880
rect 115080 800 115320 820
rect 115080 740 115090 800
rect 115150 740 115170 800
rect 115230 740 115250 800
rect 115310 740 115320 800
rect 115080 -460 115320 740
rect 115740 700 115780 7000
rect 116020 6320 116260 6330
rect 116020 6260 116030 6320
rect 116090 6260 116110 6320
rect 116170 6260 116190 6320
rect 116250 6260 116260 6320
rect 116020 6240 116260 6260
rect 116020 6180 116030 6240
rect 116090 6180 116110 6240
rect 116170 6180 116190 6240
rect 116250 6180 116260 6240
rect 116020 6160 116260 6180
rect 116020 6100 116030 6160
rect 116090 6100 116110 6160
rect 116170 6100 116190 6160
rect 116250 6100 116260 6160
rect 116020 6020 116260 6100
rect 116020 5960 116030 6020
rect 116090 5960 116110 6020
rect 116170 5960 116190 6020
rect 116250 5960 116260 6020
rect 116020 5940 116260 5960
rect 116020 5880 116030 5940
rect 116090 5880 116110 5940
rect 116170 5880 116190 5940
rect 116250 5880 116260 5940
rect 116020 5860 116260 5880
rect 115830 5830 115910 5840
rect 115830 5770 115840 5830
rect 115900 5770 115910 5830
rect 115720 690 115800 700
rect 115720 630 115730 690
rect 115790 630 115800 690
rect 115720 620 115800 630
rect 115830 200 115910 5770
rect 116020 5800 116030 5860
rect 116090 5800 116110 5860
rect 116170 5800 116190 5860
rect 116250 5800 116260 5860
rect 116020 5200 116260 5800
rect 116020 5140 116030 5200
rect 116090 5140 116110 5200
rect 116170 5140 116190 5200
rect 116250 5140 116260 5200
rect 116020 5120 116260 5140
rect 116020 5060 116030 5120
rect 116090 5060 116110 5120
rect 116170 5060 116190 5120
rect 116250 5060 116260 5120
rect 116020 5040 116260 5060
rect 116020 4980 116030 5040
rect 116090 4980 116110 5040
rect 116170 4980 116190 5040
rect 116250 4980 116260 5040
rect 116020 4720 116260 4980
rect 116020 4660 116030 4720
rect 116090 4660 116110 4720
rect 116170 4660 116190 4720
rect 116250 4660 116260 4720
rect 116020 4640 116260 4660
rect 116020 4580 116030 4640
rect 116090 4580 116110 4640
rect 116170 4580 116190 4640
rect 116250 4580 116260 4640
rect 116020 4560 116260 4580
rect 116020 4500 116030 4560
rect 116090 4500 116110 4560
rect 116170 4500 116190 4560
rect 116250 4500 116260 4560
rect 116020 4490 116260 4500
rect 116290 4990 116530 7130
rect 116290 4930 116300 4990
rect 116360 4930 116380 4990
rect 116440 4930 116460 4990
rect 116520 4930 116530 4990
rect 116290 4910 116530 4930
rect 116290 4850 116300 4910
rect 116360 4850 116380 4910
rect 116440 4850 116460 4910
rect 116520 4850 116530 4910
rect 116290 4830 116530 4850
rect 116290 4770 116300 4830
rect 116360 4770 116380 4830
rect 116440 4770 116460 4830
rect 116520 4770 116530 4830
rect 116020 4390 116260 4400
rect 116020 4330 116030 4390
rect 116090 4330 116110 4390
rect 116170 4330 116190 4390
rect 116250 4330 116260 4390
rect 116020 4310 116260 4330
rect 116020 4250 116030 4310
rect 116090 4250 116110 4310
rect 116170 4250 116190 4310
rect 116250 4250 116260 4310
rect 116020 4230 116260 4250
rect 116020 4170 116030 4230
rect 116090 4170 116110 4230
rect 116170 4170 116190 4230
rect 116250 4170 116260 4230
rect 116020 580 116260 4170
rect 116290 2780 116530 4770
rect 116560 7570 116800 7580
rect 116560 7510 116570 7570
rect 116630 7510 116650 7570
rect 116710 7510 116730 7570
rect 116790 7510 116800 7570
rect 116560 6960 116800 7510
rect 117020 7570 117100 7580
rect 117020 7510 117030 7570
rect 117090 7510 117100 7570
rect 117020 7500 117100 7510
rect 117260 7570 117340 7580
rect 117260 7510 117270 7570
rect 117330 7510 117340 7570
rect 117260 7500 117340 7510
rect 117500 7570 117580 7580
rect 117500 7510 117510 7570
rect 117570 7510 117580 7570
rect 117500 7500 117580 7510
rect 117740 7570 117820 7580
rect 117740 7510 117750 7570
rect 117810 7510 117820 7570
rect 117740 7500 117820 7510
rect 117980 7570 118060 7580
rect 117980 7510 117990 7570
rect 118050 7510 118060 7570
rect 117980 7500 118060 7510
rect 118220 7570 118300 7580
rect 118220 7510 118230 7570
rect 118290 7510 118300 7570
rect 118220 7500 118300 7510
rect 117090 7460 117150 7470
rect 117090 7390 117150 7400
rect 117210 7460 117270 7470
rect 117210 7390 117270 7400
rect 117330 7460 117390 7470
rect 117330 7390 117390 7400
rect 117450 7460 117510 7470
rect 117450 7390 117510 7400
rect 117570 7460 117630 7470
rect 117570 7390 117630 7400
rect 117690 7460 117750 7470
rect 117690 7390 117750 7400
rect 117810 7460 117870 7470
rect 117810 7390 117870 7400
rect 117930 7460 117990 7470
rect 117930 7390 117990 7400
rect 118050 7460 118110 7470
rect 118050 7390 118110 7400
rect 118170 7460 118230 7470
rect 118170 7390 118230 7400
rect 116960 7350 117040 7360
rect 116960 7290 116970 7350
rect 117030 7290 117040 7350
rect 116960 7270 117040 7290
rect 116960 7210 116970 7270
rect 117030 7210 117040 7270
rect 116960 7190 117040 7210
rect 116960 7130 116970 7190
rect 117030 7130 117040 7190
rect 116960 7120 117040 7130
rect 117180 7350 117260 7360
rect 117180 7290 117190 7350
rect 117250 7290 117260 7350
rect 117180 7270 117260 7290
rect 117180 7210 117190 7270
rect 117250 7210 117260 7270
rect 117180 7190 117260 7210
rect 117180 7130 117190 7190
rect 117250 7130 117260 7190
rect 117180 7120 117260 7130
rect 117400 7350 117480 7360
rect 117400 7290 117410 7350
rect 117470 7290 117480 7350
rect 117400 7270 117480 7290
rect 117400 7210 117410 7270
rect 117470 7210 117480 7270
rect 117400 7190 117480 7210
rect 117400 7130 117410 7190
rect 117470 7130 117480 7190
rect 117400 7120 117480 7130
rect 117620 7350 117700 7360
rect 117620 7290 117630 7350
rect 117690 7290 117700 7350
rect 117620 7270 117700 7290
rect 117620 7210 117630 7270
rect 117690 7210 117700 7270
rect 117620 7190 117700 7210
rect 117620 7130 117630 7190
rect 117690 7130 117700 7190
rect 117620 7120 117700 7130
rect 117840 7350 117920 7360
rect 117840 7290 117850 7350
rect 117910 7290 117920 7350
rect 117840 7270 117920 7290
rect 117840 7210 117850 7270
rect 117910 7210 117920 7270
rect 117840 7190 117920 7210
rect 117840 7130 117850 7190
rect 117910 7130 117920 7190
rect 117840 7120 117920 7130
rect 118060 7350 118140 7360
rect 118060 7290 118070 7350
rect 118130 7290 118140 7350
rect 118060 7270 118140 7290
rect 118060 7210 118070 7270
rect 118130 7210 118140 7270
rect 118060 7190 118140 7210
rect 118060 7130 118070 7190
rect 118130 7130 118140 7190
rect 118060 7120 118140 7130
rect 118280 7350 118360 7360
rect 118280 7290 118290 7350
rect 118350 7290 118360 7350
rect 118280 7270 118360 7290
rect 118280 7210 118290 7270
rect 118350 7210 118360 7270
rect 118280 7190 118360 7210
rect 118280 7130 118290 7190
rect 118350 7130 118360 7190
rect 118280 7120 118360 7130
rect 116560 6900 116570 6960
rect 116630 6900 116650 6960
rect 116710 6900 116730 6960
rect 116790 6900 116800 6960
rect 116560 6880 116800 6900
rect 116560 6820 116570 6880
rect 116630 6820 116650 6880
rect 116710 6820 116730 6880
rect 116790 6820 116800 6880
rect 116560 6800 116800 6820
rect 116560 6740 116570 6800
rect 116630 6740 116650 6800
rect 116710 6740 116730 6800
rect 116790 6740 116800 6800
rect 116560 5560 116800 6740
rect 116970 7020 117030 7120
rect 116970 6980 116980 7020
rect 117020 6980 117030 7020
rect 116970 6900 117030 6980
rect 117070 7000 117150 7010
rect 117070 6940 117080 7000
rect 117140 6940 117150 7000
rect 117070 6930 117150 6940
rect 116970 5760 116980 6900
rect 117020 5760 117030 6900
rect 116970 5740 117030 5760
rect 117080 6900 117140 6930
rect 117080 5760 117090 6900
rect 117130 5760 117140 6900
rect 117080 5730 117140 5760
rect 117190 6900 117250 7120
rect 117290 7000 117370 7010
rect 117290 6940 117300 7000
rect 117360 6940 117370 7000
rect 117290 6930 117370 6940
rect 117190 5760 117200 6900
rect 117240 5760 117250 6900
rect 117190 5740 117250 5760
rect 117300 6900 117360 6930
rect 117300 5760 117310 6900
rect 117350 5760 117360 6900
rect 117300 5730 117360 5760
rect 117410 6900 117470 7120
rect 117510 7000 117590 7010
rect 117510 6940 117520 7000
rect 117580 6940 117590 7000
rect 117510 6930 117590 6940
rect 117410 5760 117420 6900
rect 117460 5760 117470 6900
rect 117410 5740 117470 5760
rect 117520 6900 117580 6930
rect 117520 5760 117530 6900
rect 117570 5760 117580 6900
rect 117520 5730 117580 5760
rect 117630 6900 117690 7120
rect 117730 7000 117810 7010
rect 117730 6940 117740 7000
rect 117800 6940 117810 7000
rect 117730 6930 117810 6940
rect 117630 5760 117640 6900
rect 117680 5760 117690 6900
rect 117630 5740 117690 5760
rect 117740 6900 117800 6930
rect 117740 5760 117750 6900
rect 117790 5760 117800 6900
rect 117740 5730 117800 5760
rect 117850 6900 117910 7120
rect 117950 7000 118030 7010
rect 117950 6940 117960 7000
rect 118020 6940 118030 7000
rect 117950 6930 118030 6940
rect 117850 5760 117860 6900
rect 117900 5760 117910 6900
rect 117850 5740 117910 5760
rect 117960 6900 118020 6930
rect 117960 5760 117970 6900
rect 118010 5760 118020 6900
rect 117960 5730 118020 5760
rect 118070 6900 118130 7120
rect 118290 7020 118350 7120
rect 119010 7020 119090 7610
rect 119280 7350 119520 9120
rect 120680 9340 120920 12220
rect 120680 9280 120690 9340
rect 120750 9280 120770 9340
rect 120830 9280 120850 9340
rect 120910 9280 120920 9340
rect 120680 9260 120920 9280
rect 120680 9200 120690 9260
rect 120750 9200 120770 9260
rect 120830 9200 120850 9260
rect 120910 9200 120920 9260
rect 120680 9180 120920 9200
rect 120680 9120 120690 9180
rect 120750 9120 120770 9180
rect 120830 9120 120850 9180
rect 120910 9120 120920 9180
rect 120680 9110 120920 9120
rect 121380 9340 121620 12220
rect 121380 9280 121390 9340
rect 121450 9280 121470 9340
rect 121530 9280 121550 9340
rect 121610 9280 121620 9340
rect 121380 9260 121620 9280
rect 121380 9200 121390 9260
rect 121450 9200 121470 9260
rect 121530 9200 121550 9260
rect 121610 9200 121620 9260
rect 121380 9180 121620 9200
rect 121380 9120 121390 9180
rect 121450 9120 121470 9180
rect 121530 9120 121550 9180
rect 121610 9120 121620 9180
rect 121380 9110 121620 9120
rect 122080 9340 122320 12220
rect 122080 9280 122090 9340
rect 122150 9280 122170 9340
rect 122230 9280 122250 9340
rect 122310 9280 122320 9340
rect 122080 9260 122320 9280
rect 122080 9200 122090 9260
rect 122150 9200 122170 9260
rect 122230 9200 122250 9260
rect 122310 9200 122320 9260
rect 122080 9180 122320 9200
rect 122080 9120 122090 9180
rect 122150 9120 122170 9180
rect 122230 9120 122250 9180
rect 122310 9120 122320 9180
rect 122080 9110 122320 9120
rect 122780 9340 123020 12220
rect 122780 9280 122790 9340
rect 122850 9280 122870 9340
rect 122930 9280 122950 9340
rect 123010 9280 123020 9340
rect 122780 9260 123020 9280
rect 122780 9200 122790 9260
rect 122850 9200 122870 9260
rect 122930 9200 122950 9260
rect 123010 9200 123020 9260
rect 122780 9180 123020 9200
rect 122780 9120 122790 9180
rect 122850 9120 122870 9180
rect 122930 9120 122950 9180
rect 123010 9120 123020 9180
rect 122780 9110 123020 9120
rect 119280 7290 119290 7350
rect 119350 7290 119370 7350
rect 119430 7290 119450 7350
rect 119510 7290 119520 7350
rect 119280 7270 119520 7290
rect 119280 7210 119290 7270
rect 119350 7210 119370 7270
rect 119430 7210 119450 7270
rect 119510 7210 119520 7270
rect 119280 7190 119520 7210
rect 119280 7130 119290 7190
rect 119350 7130 119370 7190
rect 119430 7130 119450 7190
rect 119510 7130 119520 7190
rect 119280 7120 119520 7130
rect 118170 7000 118250 7010
rect 118170 6940 118180 7000
rect 118240 6940 118250 7000
rect 118170 6930 118250 6940
rect 118290 6980 118300 7020
rect 118340 6980 118350 7020
rect 118070 5760 118080 6900
rect 118120 5760 118130 6900
rect 118070 5740 118130 5760
rect 118180 6900 118240 6930
rect 118180 5760 118190 6900
rect 118230 5760 118240 6900
rect 118180 5730 118240 5760
rect 118290 6900 118350 6980
rect 118910 7000 119192 7020
rect 118910 6960 118920 7000
rect 118960 6960 119030 7000
rect 119070 6960 119140 7000
rect 119180 6960 119192 7000
rect 118910 6940 119192 6960
rect 118290 5760 118300 6900
rect 118340 5760 118350 6900
rect 118290 5740 118350 5760
rect 118910 5790 119192 5810
rect 118910 5750 118920 5790
rect 118960 5750 119030 5790
rect 119070 5750 119140 5790
rect 119180 5750 119192 5790
rect 118910 5730 119192 5750
rect 116560 5500 116570 5560
rect 116630 5500 116650 5560
rect 116710 5500 116730 5560
rect 116790 5500 116800 5560
rect 116560 5480 116800 5500
rect 116560 5420 116570 5480
rect 116630 5420 116650 5480
rect 116710 5420 116730 5480
rect 116790 5420 116800 5480
rect 116560 5400 116800 5420
rect 116560 5340 116570 5400
rect 116630 5340 116650 5400
rect 116710 5340 116730 5400
rect 116790 5340 116800 5400
rect 116560 3810 116800 5340
rect 117070 5720 117150 5730
rect 117070 5660 117080 5720
rect 117140 5660 117150 5720
rect 117070 5270 117150 5660
rect 117290 5720 117370 5730
rect 117290 5660 117300 5720
rect 117360 5660 117370 5720
rect 117290 5270 117370 5660
rect 117510 5720 117590 5730
rect 117510 5660 117520 5720
rect 117580 5660 117590 5720
rect 117510 5270 117590 5660
rect 117730 5720 117810 5730
rect 117730 5660 117740 5720
rect 117800 5660 117810 5720
rect 117620 5560 117700 5570
rect 117620 5500 117630 5560
rect 117690 5500 117700 5560
rect 117620 5480 117700 5500
rect 117620 5420 117630 5480
rect 117690 5420 117700 5480
rect 117620 5400 117700 5420
rect 117620 5340 117630 5400
rect 117690 5340 117700 5400
rect 117620 5330 117700 5340
rect 117730 5270 117810 5660
rect 117950 5720 118030 5730
rect 117950 5660 117960 5720
rect 118020 5660 118030 5720
rect 117950 5270 118030 5660
rect 118170 5720 118250 5730
rect 118170 5660 118180 5720
rect 118240 5660 118250 5720
rect 118170 5270 118250 5660
rect 118930 5560 119170 5730
rect 118930 5500 118940 5560
rect 119000 5500 119020 5560
rect 119080 5500 119100 5560
rect 119160 5500 119170 5560
rect 118930 5480 119170 5500
rect 118930 5420 118940 5480
rect 119000 5420 119020 5480
rect 119080 5420 119100 5480
rect 119160 5420 119170 5480
rect 118930 5400 119170 5420
rect 118930 5340 118940 5400
rect 119000 5340 119020 5400
rect 119080 5340 119100 5400
rect 119160 5340 119170 5400
rect 118930 5330 119170 5340
rect 117070 5260 118250 5270
rect 117070 5200 117080 5260
rect 117140 5200 117190 5260
rect 117250 5200 117300 5260
rect 117360 5200 117410 5260
rect 117470 5200 117520 5260
rect 117580 5200 117630 5260
rect 117690 5200 117740 5260
rect 117800 5200 117850 5260
rect 117910 5200 117960 5260
rect 118020 5200 118070 5260
rect 118130 5200 118180 5260
rect 118240 5200 118250 5260
rect 117070 5180 118250 5200
rect 117070 5120 117080 5180
rect 117140 5120 117190 5180
rect 117250 5120 117300 5180
rect 117360 5120 117410 5180
rect 117470 5120 117520 5180
rect 117580 5120 117630 5180
rect 117690 5120 117740 5180
rect 117800 5120 117850 5180
rect 117910 5120 117960 5180
rect 118020 5120 118070 5180
rect 118130 5120 118180 5180
rect 118240 5120 118250 5180
rect 117070 5100 118250 5120
rect 117070 5040 117080 5100
rect 117140 5040 117190 5100
rect 117250 5040 117300 5100
rect 117360 5040 117410 5100
rect 117470 5040 117520 5100
rect 117580 5040 117630 5100
rect 117690 5040 117740 5100
rect 117800 5040 117850 5100
rect 117910 5040 117960 5100
rect 118020 5040 118070 5100
rect 118130 5040 118180 5100
rect 118240 5040 118250 5100
rect 117070 5030 118250 5040
rect 119120 5260 119620 5270
rect 119120 5200 119130 5260
rect 119190 5200 119210 5260
rect 119270 5200 119300 5260
rect 119360 5200 119380 5260
rect 119440 5200 119470 5260
rect 119530 5200 119550 5260
rect 119610 5200 119620 5260
rect 119120 5180 119620 5200
rect 119120 5120 119130 5180
rect 119190 5120 119210 5180
rect 119270 5120 119300 5180
rect 119360 5120 119380 5180
rect 119440 5120 119470 5180
rect 119530 5120 119550 5180
rect 119610 5120 119620 5180
rect 119120 5100 119620 5120
rect 119120 5040 119130 5100
rect 119190 5040 119210 5100
rect 119270 5040 119300 5100
rect 119360 5040 119380 5100
rect 119440 5040 119470 5100
rect 119530 5040 119550 5100
rect 119610 5040 119620 5100
rect 116960 4990 117040 5000
rect 116960 4930 116970 4990
rect 117030 4930 117040 4990
rect 116960 4910 117040 4930
rect 116960 4850 116970 4910
rect 117030 4850 117040 4910
rect 116960 4830 117040 4850
rect 116960 4770 116970 4830
rect 117030 4770 117040 4830
rect 116960 4760 117040 4770
rect 118280 4990 118360 5000
rect 118280 4930 118290 4990
rect 118350 4930 118360 4990
rect 118280 4910 118360 4930
rect 118280 4850 118290 4910
rect 118350 4850 118360 4910
rect 118280 4830 118360 4850
rect 118280 4770 118290 4830
rect 118350 4770 118360 4830
rect 118280 4760 118360 4770
rect 116970 4470 117030 4760
rect 117070 4720 117150 4730
rect 117070 4660 117080 4720
rect 117140 4660 117150 4720
rect 117070 4640 117150 4660
rect 117070 4580 117080 4640
rect 117140 4580 117150 4640
rect 117070 4560 117150 4580
rect 117070 4500 117080 4560
rect 117140 4500 117150 4560
rect 117070 4490 117150 4500
rect 117290 4720 117370 4730
rect 117290 4660 117300 4720
rect 117360 4660 117370 4720
rect 117290 4640 117370 4660
rect 117290 4580 117300 4640
rect 117360 4580 117370 4640
rect 117290 4560 117370 4580
rect 117290 4500 117300 4560
rect 117360 4500 117370 4560
rect 117290 4490 117370 4500
rect 117510 4720 117590 4730
rect 117510 4660 117520 4720
rect 117580 4660 117590 4720
rect 117510 4640 117590 4660
rect 117510 4580 117520 4640
rect 117580 4580 117590 4640
rect 117510 4560 117590 4580
rect 117510 4500 117520 4560
rect 117580 4500 117590 4560
rect 117510 4490 117590 4500
rect 117730 4720 117810 4730
rect 117730 4660 117740 4720
rect 117800 4660 117810 4720
rect 117730 4640 117810 4660
rect 117730 4580 117740 4640
rect 117800 4580 117810 4640
rect 117730 4560 117810 4580
rect 117730 4500 117740 4560
rect 117800 4500 117810 4560
rect 117730 4490 117810 4500
rect 117950 4720 118030 4730
rect 117950 4660 117960 4720
rect 118020 4660 118030 4720
rect 117950 4640 118030 4660
rect 117950 4580 117960 4640
rect 118020 4580 118030 4640
rect 117950 4560 118030 4580
rect 117950 4500 117960 4560
rect 118020 4500 118030 4560
rect 117950 4490 118030 4500
rect 118170 4720 118250 4730
rect 118170 4660 118180 4720
rect 118240 4660 118250 4720
rect 118170 4640 118250 4660
rect 118170 4580 118180 4640
rect 118240 4580 118250 4640
rect 118170 4560 118250 4580
rect 118170 4500 118180 4560
rect 118240 4500 118250 4560
rect 118170 4490 118250 4500
rect 116970 4430 116980 4470
rect 117020 4430 117030 4470
rect 116970 4350 117030 4430
rect 116970 4010 116980 4350
rect 117020 4010 117030 4350
rect 116970 3990 117030 4010
rect 117080 4350 117140 4490
rect 117180 4450 117260 4460
rect 117180 4390 117190 4450
rect 117250 4390 117260 4450
rect 117180 4380 117260 4390
rect 117080 4010 117090 4350
rect 117130 4010 117140 4350
rect 117080 3990 117140 4010
rect 117190 4350 117250 4380
rect 117190 4010 117200 4350
rect 117240 4010 117250 4350
rect 117190 3950 117250 4010
rect 117300 4350 117360 4490
rect 117400 4450 117480 4460
rect 117400 4390 117410 4450
rect 117470 4390 117480 4450
rect 117400 4380 117480 4390
rect 117300 4010 117310 4350
rect 117350 4010 117360 4350
rect 117300 3990 117360 4010
rect 117410 4350 117470 4380
rect 117410 4010 117420 4350
rect 117460 4010 117470 4350
rect 117410 3950 117470 4010
rect 117520 4350 117580 4490
rect 117620 4450 117700 4460
rect 117620 4390 117630 4450
rect 117690 4390 117700 4450
rect 117620 4380 117700 4390
rect 117520 4010 117530 4350
rect 117570 4010 117580 4350
rect 117520 3990 117580 4010
rect 117630 4350 117690 4380
rect 117630 4010 117640 4350
rect 117680 4010 117690 4350
rect 117630 3950 117690 4010
rect 117740 4350 117800 4490
rect 117840 4450 117920 4460
rect 117840 4390 117850 4450
rect 117910 4390 117920 4450
rect 117840 4380 117920 4390
rect 117740 4010 117750 4350
rect 117790 4010 117800 4350
rect 117740 3990 117800 4010
rect 117850 4350 117910 4380
rect 117850 4010 117860 4350
rect 117900 4010 117910 4350
rect 117850 3950 117910 4010
rect 117960 4350 118020 4490
rect 118060 4450 118140 4460
rect 118060 4390 118070 4450
rect 118130 4390 118140 4450
rect 118060 4380 118140 4390
rect 117960 4010 117970 4350
rect 118010 4010 118020 4350
rect 117960 3990 118020 4010
rect 118070 4350 118130 4380
rect 118070 4010 118080 4350
rect 118120 4010 118130 4350
rect 118070 3950 118130 4010
rect 118180 4350 118240 4490
rect 118180 4010 118190 4350
rect 118230 4010 118240 4350
rect 118180 3990 118240 4010
rect 118290 4470 118350 4760
rect 118290 4430 118300 4470
rect 118340 4430 118350 4470
rect 118290 4350 118350 4430
rect 118290 4010 118300 4350
rect 118340 4010 118350 4350
rect 118290 3990 118350 4010
rect 119120 4120 119620 5040
rect 119120 4060 119140 4120
rect 119200 4060 119240 4120
rect 119300 4060 119340 4120
rect 119400 4060 119440 4120
rect 119500 4060 119540 4120
rect 119600 4060 119620 4120
rect 119120 4020 119620 4060
rect 119120 3960 119140 4020
rect 119200 3960 119240 4020
rect 119300 3960 119340 4020
rect 119400 3960 119440 4020
rect 119500 3960 119540 4020
rect 119600 3960 119620 4020
rect 117180 3940 117260 3950
rect 117180 3880 117190 3940
rect 117250 3880 117260 3940
rect 117180 3870 117260 3880
rect 117400 3940 117480 3950
rect 117400 3880 117410 3940
rect 117470 3880 117480 3940
rect 117400 3870 117480 3880
rect 117620 3940 117700 3950
rect 117620 3880 117630 3940
rect 117690 3880 117700 3940
rect 117620 3870 117700 3880
rect 117840 3940 117920 3950
rect 117840 3880 117850 3940
rect 117910 3880 117920 3940
rect 117840 3870 117920 3880
rect 118060 3940 118140 3950
rect 118060 3880 118070 3940
rect 118130 3880 118140 3940
rect 118060 3870 118140 3880
rect 118550 3940 118630 3950
rect 118550 3880 118560 3940
rect 118620 3880 118630 3940
rect 118550 3870 118630 3880
rect 119120 3920 119620 3960
rect 116560 3750 116570 3810
rect 116630 3750 116650 3810
rect 116710 3750 116730 3810
rect 116790 3750 116800 3810
rect 116560 3730 116800 3750
rect 116560 3670 116570 3730
rect 116630 3670 116650 3730
rect 116710 3670 116730 3730
rect 116790 3670 116800 3730
rect 116560 3050 116800 3670
rect 117290 3810 117370 3820
rect 117290 3750 117300 3810
rect 117360 3750 117370 3810
rect 117290 3730 117370 3750
rect 117290 3670 117300 3730
rect 117360 3670 117370 3730
rect 117290 3660 117370 3670
rect 117180 3570 117260 3580
rect 117180 3510 117190 3570
rect 117250 3510 117260 3570
rect 117180 3500 117260 3510
rect 117400 3570 117480 3580
rect 117400 3510 117410 3570
rect 117470 3510 117480 3570
rect 117400 3500 117480 3510
rect 117620 3570 117700 3580
rect 117620 3510 117630 3570
rect 117690 3510 117700 3570
rect 117620 3500 117700 3510
rect 117840 3570 117920 3580
rect 117840 3510 117850 3570
rect 117910 3510 117920 3570
rect 117840 3500 117920 3510
rect 118060 3570 118140 3580
rect 118060 3510 118070 3570
rect 118130 3510 118140 3570
rect 118060 3500 118140 3510
rect 118460 3570 118540 3580
rect 118460 3510 118470 3570
rect 118530 3510 118540 3570
rect 118460 3500 118540 3510
rect 116560 2990 116570 3050
rect 116630 2990 116650 3050
rect 116710 2990 116730 3050
rect 116790 2990 116800 3050
rect 116560 2970 116800 2990
rect 116560 2910 116570 2970
rect 116630 2910 116650 2970
rect 116710 2910 116730 2970
rect 116790 2910 116800 2970
rect 116560 2890 116800 2910
rect 116560 2830 116570 2890
rect 116630 2830 116650 2890
rect 116710 2830 116730 2890
rect 116790 2830 116800 2890
rect 116560 2820 116800 2830
rect 116970 3470 117030 3490
rect 116970 2930 116980 3470
rect 117020 2930 117030 3470
rect 116970 2850 117030 2930
rect 116290 2720 116300 2780
rect 116360 2720 116380 2780
rect 116440 2720 116460 2780
rect 116520 2720 116530 2780
rect 116290 2700 116530 2720
rect 116290 2640 116300 2700
rect 116360 2640 116380 2700
rect 116440 2640 116460 2700
rect 116520 2640 116530 2700
rect 116290 2620 116530 2640
rect 116290 2560 116300 2620
rect 116360 2560 116380 2620
rect 116440 2560 116460 2620
rect 116520 2560 116530 2620
rect 116290 2550 116530 2560
rect 116970 2810 116980 2850
rect 117020 2810 117030 2850
rect 116970 2510 117030 2810
rect 117080 3470 117140 3490
rect 117080 2930 117090 3470
rect 117130 2930 117140 3470
rect 117080 2790 117140 2930
rect 117190 3470 117250 3500
rect 117190 2930 117200 3470
rect 117240 2930 117250 3470
rect 117190 2900 117250 2930
rect 117300 3470 117360 3490
rect 117300 2930 117310 3470
rect 117350 2930 117360 3470
rect 117180 2890 117260 2900
rect 117180 2830 117190 2890
rect 117250 2830 117260 2890
rect 117180 2820 117260 2830
rect 117300 2790 117360 2930
rect 117410 3470 117470 3500
rect 117410 2930 117420 3470
rect 117460 2930 117470 3470
rect 117410 2900 117470 2930
rect 117520 3470 117580 3490
rect 117520 2930 117530 3470
rect 117570 2930 117580 3470
rect 117400 2890 117480 2900
rect 117400 2830 117410 2890
rect 117470 2830 117480 2890
rect 117400 2820 117480 2830
rect 117520 2790 117580 2930
rect 117630 3470 117690 3500
rect 117630 2930 117640 3470
rect 117680 2930 117690 3470
rect 117630 2900 117690 2930
rect 117740 3470 117800 3490
rect 117740 2930 117750 3470
rect 117790 2930 117800 3470
rect 117620 2890 117700 2900
rect 117620 2830 117630 2890
rect 117690 2830 117700 2890
rect 117620 2820 117700 2830
rect 117740 2790 117800 2930
rect 117850 3470 117910 3500
rect 117850 2930 117860 3470
rect 117900 2930 117910 3470
rect 117850 2900 117910 2930
rect 117960 3470 118020 3490
rect 117960 2930 117970 3470
rect 118010 2930 118020 3470
rect 117840 2890 117920 2900
rect 117840 2830 117850 2890
rect 117910 2830 117920 2890
rect 117840 2820 117920 2830
rect 117960 2790 118020 2930
rect 118070 3470 118130 3500
rect 118070 2930 118080 3470
rect 118120 2930 118130 3470
rect 118070 2900 118130 2930
rect 118180 3470 118240 3490
rect 118180 2930 118190 3470
rect 118230 2930 118240 3470
rect 118060 2890 118140 2900
rect 118060 2830 118070 2890
rect 118130 2830 118140 2890
rect 118060 2820 118140 2830
rect 118180 2790 118240 2930
rect 118290 3470 118350 3490
rect 118290 2930 118300 3470
rect 118340 2930 118350 3470
rect 118480 2940 118520 3500
rect 118290 2850 118350 2930
rect 118460 2930 118540 2940
rect 118460 2870 118470 2930
rect 118530 2870 118540 2930
rect 118460 2860 118540 2870
rect 118290 2810 118300 2850
rect 118340 2810 118350 2850
rect 117070 2780 117150 2790
rect 117070 2720 117080 2780
rect 117140 2720 117150 2780
rect 117070 2700 117150 2720
rect 117070 2640 117080 2700
rect 117140 2640 117150 2700
rect 117070 2620 117150 2640
rect 117070 2560 117080 2620
rect 117140 2560 117150 2620
rect 117070 2550 117150 2560
rect 117290 2780 117370 2790
rect 117290 2720 117300 2780
rect 117360 2720 117370 2780
rect 117290 2700 117370 2720
rect 117290 2640 117300 2700
rect 117360 2640 117370 2700
rect 117290 2620 117370 2640
rect 117290 2560 117300 2620
rect 117360 2560 117370 2620
rect 117290 2550 117370 2560
rect 117510 2780 117590 2790
rect 117510 2720 117520 2780
rect 117580 2720 117590 2780
rect 117510 2700 117590 2720
rect 117510 2640 117520 2700
rect 117580 2640 117590 2700
rect 117510 2620 117590 2640
rect 117510 2560 117520 2620
rect 117580 2560 117590 2620
rect 117510 2550 117590 2560
rect 117730 2780 117810 2790
rect 117730 2720 117740 2780
rect 117800 2720 117810 2780
rect 117730 2700 117810 2720
rect 117730 2640 117740 2700
rect 117800 2640 117810 2700
rect 117730 2620 117810 2640
rect 117730 2560 117740 2620
rect 117800 2560 117810 2620
rect 117730 2550 117810 2560
rect 117950 2780 118030 2790
rect 117950 2720 117960 2780
rect 118020 2720 118030 2780
rect 117950 2700 118030 2720
rect 117950 2640 117960 2700
rect 118020 2640 118030 2700
rect 117950 2620 118030 2640
rect 117950 2560 117960 2620
rect 118020 2560 118030 2620
rect 117950 2550 118030 2560
rect 118170 2780 118250 2790
rect 118170 2720 118180 2780
rect 118240 2720 118250 2780
rect 118170 2700 118250 2720
rect 118170 2640 118180 2700
rect 118240 2640 118250 2700
rect 118170 2620 118250 2640
rect 118170 2560 118180 2620
rect 118240 2560 118250 2620
rect 118170 2550 118250 2560
rect 118290 2510 118350 2810
rect 118570 2800 118610 3870
rect 119120 3860 119140 3920
rect 119200 3860 119240 3920
rect 119300 3860 119340 3920
rect 119400 3860 119440 3920
rect 119500 3860 119540 3920
rect 119600 3860 119620 3920
rect 118660 2940 118730 2950
rect 118660 2860 118730 2870
rect 118780 2940 118850 2950
rect 118780 2860 118850 2870
rect 118900 2940 118970 2950
rect 118900 2860 118970 2870
rect 119020 2940 119090 2952
rect 119020 2860 119090 2870
rect 118790 2800 118830 2860
rect 118550 2790 118630 2800
rect 118550 2730 118560 2790
rect 118620 2730 118630 2790
rect 118550 2720 118630 2730
rect 118770 2790 118850 2800
rect 118770 2730 118780 2790
rect 118840 2730 118850 2790
rect 118770 2720 118850 2730
rect 116960 2500 117040 2510
rect 116960 2440 116970 2500
rect 117030 2440 117040 2500
rect 116960 2420 117040 2440
rect 116960 2360 116970 2420
rect 117030 2360 117040 2420
rect 116960 2340 117040 2360
rect 116960 2280 116970 2340
rect 117030 2280 117040 2340
rect 116960 2270 117040 2280
rect 118280 2500 118360 2510
rect 118280 2440 118290 2500
rect 118350 2440 118360 2500
rect 118280 2420 118360 2440
rect 118280 2360 118290 2420
rect 118350 2360 118360 2420
rect 118280 2340 118360 2360
rect 118280 2280 118290 2340
rect 118350 2280 118360 2340
rect 118280 2270 118360 2280
rect 119030 2240 119070 2860
rect 119010 2230 119090 2240
rect 119010 2170 119020 2230
rect 119080 2170 119090 2230
rect 119010 2160 119090 2170
rect 118880 1850 118960 1860
rect 118880 1790 118890 1850
rect 118950 1790 118960 1850
rect 117220 1740 118100 1750
rect 117220 1680 117230 1740
rect 117290 1680 117310 1740
rect 117370 1680 117390 1740
rect 117450 1680 117470 1740
rect 117530 1680 117550 1740
rect 117610 1680 117630 1740
rect 117690 1680 117710 1740
rect 117770 1680 117790 1740
rect 117850 1680 117870 1740
rect 117930 1680 117950 1740
rect 118010 1680 118030 1740
rect 118090 1680 118100 1740
rect 117220 1660 118100 1680
rect 117220 1600 117230 1660
rect 117290 1600 117310 1660
rect 117370 1600 117390 1660
rect 117450 1600 117470 1660
rect 117530 1600 117550 1660
rect 117610 1600 117630 1660
rect 117690 1600 117710 1660
rect 117770 1600 117790 1660
rect 117850 1600 117870 1660
rect 117930 1600 117950 1660
rect 118010 1600 118030 1660
rect 118090 1600 118100 1660
rect 117220 1580 118100 1600
rect 117220 1520 117230 1580
rect 117290 1520 117310 1580
rect 117370 1520 117390 1580
rect 117450 1520 117470 1580
rect 117530 1520 117550 1580
rect 117610 1520 117630 1580
rect 117690 1520 117710 1580
rect 117770 1520 117790 1580
rect 117850 1520 117870 1580
rect 117930 1520 117950 1580
rect 118010 1520 118030 1580
rect 118090 1520 118100 1580
rect 117220 1510 118100 1520
rect 118750 1740 118830 1750
rect 118750 1680 118760 1740
rect 118820 1680 118830 1740
rect 118750 1660 118830 1680
rect 118750 1600 118760 1660
rect 118820 1600 118830 1660
rect 118750 1580 118830 1600
rect 118750 1520 118760 1580
rect 118820 1520 118830 1580
rect 118750 1510 118830 1520
rect 116020 520 116030 580
rect 116090 520 116110 580
rect 116170 520 116190 580
rect 116250 520 116260 580
rect 116020 500 116260 520
rect 116020 440 116030 500
rect 116090 440 116110 500
rect 116170 440 116190 500
rect 116250 440 116260 500
rect 116020 420 116260 440
rect 116020 360 116030 420
rect 116090 360 116110 420
rect 116170 360 116190 420
rect 116250 360 116260 420
rect 116020 350 116260 360
rect 117030 1350 117090 1370
rect 115830 140 115840 200
rect 115900 140 115910 200
rect 115830 130 115910 140
rect 115080 -520 115090 -460
rect 115150 -520 115170 -460
rect 115230 -520 115250 -460
rect 115310 -520 115320 -460
rect 115080 -540 115320 -520
rect 115080 -600 115090 -540
rect 115150 -600 115170 -540
rect 115230 -600 115250 -540
rect 115310 -600 115320 -540
rect 115080 -620 115320 -600
rect 115080 -680 115090 -620
rect 115150 -680 115170 -620
rect 115230 -680 115250 -620
rect 115310 -680 115320 -620
rect 115080 -690 115320 -680
rect 117030 10 117040 1350
rect 117080 10 117090 1350
rect 117030 -70 117090 10
rect 117230 1350 117290 1510
rect 117320 1470 117400 1480
rect 117320 1410 117330 1470
rect 117390 1410 117400 1470
rect 117320 1400 117400 1410
rect 117520 1470 117600 1480
rect 117520 1410 117530 1470
rect 117590 1410 117600 1470
rect 117520 1400 117600 1410
rect 117230 10 117240 1350
rect 117280 10 117290 1350
rect 117230 -20 117290 10
rect 117430 1350 117490 1370
rect 117430 10 117440 1350
rect 117480 10 117490 1350
rect 117030 -110 117040 -70
rect 117080 -110 117090 -70
rect 117220 -30 117300 -20
rect 117220 -90 117230 -30
rect 117290 -90 117300 -30
rect 117220 -100 117300 -90
rect 117030 -1150 117090 -110
rect 117430 -1150 117490 10
rect 117630 1350 117690 1510
rect 117720 1470 117800 1480
rect 117720 1410 117730 1470
rect 117790 1410 117800 1470
rect 117720 1400 117800 1410
rect 117920 1470 118000 1480
rect 117920 1410 117930 1470
rect 117990 1410 118000 1470
rect 117920 1400 118000 1410
rect 117630 10 117640 1350
rect 117680 10 117690 1350
rect 117630 -20 117690 10
rect 117830 1350 117890 1370
rect 117830 10 117840 1350
rect 117880 10 117890 1350
rect 117620 -30 117700 -20
rect 117620 -90 117630 -30
rect 117690 -90 117700 -30
rect 117620 -100 117700 -90
rect 114970 -1220 114980 -1160
rect 115040 -1220 115050 -1160
rect 114970 -1240 115050 -1220
rect 114970 -1300 114980 -1240
rect 115040 -1300 115050 -1240
rect 114970 -1320 115050 -1300
rect 114970 -1380 114980 -1320
rect 115040 -1380 115050 -1320
rect 114970 -1390 115050 -1380
rect 115080 -1160 115320 -1150
rect 115080 -1220 115090 -1160
rect 115150 -1220 115170 -1160
rect 115230 -1220 115250 -1160
rect 115310 -1220 115320 -1160
rect 115080 -1240 115320 -1220
rect 115080 -1300 115090 -1240
rect 115150 -1300 115170 -1240
rect 115230 -1300 115250 -1240
rect 115310 -1300 115320 -1240
rect 115080 -1320 115320 -1300
rect 115080 -1380 115090 -1320
rect 115150 -1380 115170 -1320
rect 115230 -1380 115250 -1320
rect 115310 -1380 115320 -1320
rect 115080 -3000 115320 -1380
rect 115780 -1160 116020 -1150
rect 115780 -1220 115790 -1160
rect 115850 -1220 115870 -1160
rect 115930 -1220 115950 -1160
rect 116010 -1220 116020 -1160
rect 115780 -1240 116020 -1220
rect 115780 -1300 115790 -1240
rect 115850 -1300 115870 -1240
rect 115930 -1300 115950 -1240
rect 116010 -1300 116020 -1240
rect 115780 -1320 116020 -1300
rect 115780 -1380 115790 -1320
rect 115850 -1380 115870 -1320
rect 115930 -1380 115950 -1320
rect 116010 -1380 116020 -1320
rect 115780 -3000 116020 -1380
rect 116480 -1160 116720 -1150
rect 116480 -1220 116490 -1160
rect 116550 -1220 116570 -1160
rect 116630 -1220 116650 -1160
rect 116710 -1220 116720 -1160
rect 116480 -1240 116720 -1220
rect 116480 -1300 116490 -1240
rect 116550 -1300 116570 -1240
rect 116630 -1300 116650 -1240
rect 116710 -1300 116720 -1240
rect 116480 -1320 116720 -1300
rect 116480 -1380 116490 -1320
rect 116550 -1380 116570 -1320
rect 116630 -1380 116650 -1320
rect 116710 -1380 116720 -1320
rect 116480 -3000 116720 -1380
rect 117020 -1160 117100 -1150
rect 117020 -1220 117030 -1160
rect 117090 -1220 117100 -1160
rect 117020 -1240 117100 -1220
rect 117020 -1300 117030 -1240
rect 117090 -1300 117100 -1240
rect 117020 -1320 117100 -1300
rect 117020 -1380 117030 -1320
rect 117090 -1380 117100 -1320
rect 117020 -1390 117100 -1380
rect 117180 -1160 117490 -1150
rect 117180 -1220 117190 -1160
rect 117250 -1220 117270 -1160
rect 117330 -1220 117350 -1160
rect 117410 -1220 117490 -1160
rect 117180 -1240 117490 -1220
rect 117180 -1300 117190 -1240
rect 117250 -1300 117270 -1240
rect 117330 -1300 117350 -1240
rect 117410 -1300 117490 -1240
rect 117180 -1320 117490 -1300
rect 117180 -1380 117190 -1320
rect 117250 -1380 117270 -1320
rect 117330 -1380 117350 -1320
rect 117410 -1380 117490 -1320
rect 117180 -1390 117490 -1380
rect 117830 -1150 117890 10
rect 118030 1350 118090 1510
rect 118030 10 118040 1350
rect 118080 10 118090 1350
rect 118030 -20 118090 10
rect 118230 1350 118290 1370
rect 118230 10 118240 1350
rect 118280 10 118290 1350
rect 118760 1360 118830 1510
rect 118760 1280 118830 1290
rect 118880 1470 118960 1790
rect 119120 1740 119620 3860
rect 119120 1680 119130 1740
rect 119190 1680 119210 1740
rect 119270 1680 119300 1740
rect 119360 1680 119380 1740
rect 119440 1680 119470 1740
rect 119530 1680 119550 1740
rect 119610 1680 119620 1740
rect 119120 1660 119620 1680
rect 119120 1600 119130 1660
rect 119190 1600 119210 1660
rect 119270 1600 119300 1660
rect 119360 1600 119380 1660
rect 119440 1600 119470 1660
rect 119530 1600 119550 1660
rect 119610 1600 119620 1660
rect 119120 1580 119620 1600
rect 119120 1520 119130 1580
rect 119190 1520 119210 1580
rect 119270 1520 119300 1580
rect 119360 1520 119380 1580
rect 119440 1520 119470 1580
rect 119530 1520 119550 1580
rect 119610 1520 119620 1580
rect 119120 1510 119620 1520
rect 119680 4710 119920 4720
rect 119680 4650 119690 4710
rect 119750 4650 119770 4710
rect 119830 4650 119850 4710
rect 119910 4650 119920 4710
rect 119680 4630 119920 4650
rect 119680 4570 119690 4630
rect 119750 4570 119770 4630
rect 119830 4570 119850 4630
rect 119910 4570 119920 4630
rect 119680 4550 119920 4570
rect 119680 4490 119690 4550
rect 119750 4490 119770 4550
rect 119830 4490 119850 4550
rect 119910 4490 119920 4550
rect 119680 2500 119920 4490
rect 119680 2440 119690 2500
rect 119750 2440 119770 2500
rect 119830 2440 119850 2500
rect 119910 2440 119920 2500
rect 119680 2420 119920 2440
rect 119680 2360 119690 2420
rect 119750 2360 119770 2420
rect 119830 2360 119850 2420
rect 119910 2360 119920 2420
rect 119680 2340 119920 2360
rect 119680 2280 119690 2340
rect 119750 2280 119770 2340
rect 119830 2280 119850 2340
rect 119910 2280 119920 2340
rect 118880 1410 118890 1470
rect 118950 1410 118960 1470
rect 118880 1370 118960 1410
rect 118880 1360 118950 1370
rect 118880 1280 118950 1290
rect 118020 -30 118100 -20
rect 118020 -90 118030 -30
rect 118090 -90 118100 -30
rect 118020 -100 118100 -90
rect 118230 -70 118290 10
rect 118230 -110 118240 -70
rect 118280 -110 118290 -70
rect 118230 -1150 118290 -110
rect 117830 -1160 118120 -1150
rect 117830 -1220 117890 -1160
rect 117950 -1220 117970 -1160
rect 118030 -1220 118050 -1160
rect 118110 -1220 118120 -1160
rect 117830 -1240 118120 -1220
rect 117830 -1300 117890 -1240
rect 117950 -1300 117970 -1240
rect 118030 -1300 118050 -1240
rect 118110 -1300 118120 -1240
rect 117830 -1320 118120 -1300
rect 117830 -1380 117890 -1320
rect 117950 -1380 117970 -1320
rect 118030 -1380 118050 -1320
rect 118110 -1380 118120 -1320
rect 117830 -1390 118120 -1380
rect 118220 -1160 118300 -1150
rect 118220 -1220 118230 -1160
rect 118290 -1220 118300 -1160
rect 118220 -1240 118300 -1220
rect 118220 -1300 118230 -1240
rect 118290 -1300 118300 -1240
rect 118220 -1320 118300 -1300
rect 118220 -1380 118230 -1320
rect 118290 -1380 118300 -1320
rect 118220 -1390 118300 -1380
rect 118740 -1160 118980 -1150
rect 118740 -1220 118750 -1160
rect 118810 -1220 118830 -1160
rect 118890 -1220 118910 -1160
rect 118970 -1220 118980 -1160
rect 118740 -1240 118980 -1220
rect 118740 -1300 118750 -1240
rect 118810 -1300 118830 -1240
rect 118890 -1300 118910 -1240
rect 118970 -1300 118980 -1240
rect 118740 -1320 118980 -1300
rect 118740 -1380 118750 -1320
rect 118810 -1380 118830 -1320
rect 118890 -1380 118910 -1320
rect 118970 -1380 118980 -1320
rect 118740 -1390 118980 -1380
rect 119280 -1160 119520 -1150
rect 119280 -1220 119290 -1160
rect 119350 -1220 119370 -1160
rect 119430 -1220 119450 -1160
rect 119510 -1220 119520 -1160
rect 119280 -1240 119520 -1220
rect 119280 -1300 119290 -1240
rect 119350 -1300 119370 -1240
rect 119430 -1300 119450 -1240
rect 119510 -1300 119520 -1240
rect 119280 -1320 119520 -1300
rect 119280 -1380 119290 -1320
rect 119350 -1380 119370 -1320
rect 119430 -1380 119450 -1320
rect 119510 -1380 119520 -1320
rect 117180 -3000 117420 -1390
rect 117880 -3000 118120 -1390
rect 118580 -3000 118820 -1390
rect 119280 -3000 119520 -1380
rect 119680 -1160 119920 2280
rect 119680 -1220 119690 -1160
rect 119750 -1220 119770 -1160
rect 119830 -1220 119850 -1160
rect 119910 -1220 119920 -1160
rect 119680 -1240 119920 -1220
rect 119680 -1300 119690 -1240
rect 119750 -1300 119770 -1240
rect 119830 -1300 119850 -1240
rect 119910 -1300 119920 -1240
rect 119680 -1320 119920 -1300
rect 119680 -1380 119690 -1320
rect 119750 -1380 119770 -1320
rect 119830 -1380 119850 -1320
rect 119910 -1380 119920 -1320
rect 119680 -1390 119920 -1380
rect 119980 -1160 120220 -1150
rect 119980 -1220 119990 -1160
rect 120050 -1220 120070 -1160
rect 120130 -1220 120150 -1160
rect 120210 -1220 120220 -1160
rect 119980 -1240 120220 -1220
rect 119980 -1300 119990 -1240
rect 120050 -1300 120070 -1240
rect 120130 -1300 120150 -1240
rect 120210 -1300 120220 -1240
rect 119980 -1320 120220 -1300
rect 119980 -1380 119990 -1320
rect 120050 -1380 120070 -1320
rect 120130 -1380 120150 -1320
rect 120210 -1380 120220 -1320
rect 119980 -3000 120220 -1380
rect 120680 -1160 120920 -1150
rect 120680 -1220 120690 -1160
rect 120750 -1220 120770 -1160
rect 120830 -1220 120850 -1160
rect 120910 -1220 120920 -1160
rect 120680 -1240 120920 -1220
rect 120680 -1300 120690 -1240
rect 120750 -1300 120770 -1240
rect 120830 -1300 120850 -1240
rect 120910 -1300 120920 -1240
rect 120680 -1320 120920 -1300
rect 120680 -1380 120690 -1320
rect 120750 -1380 120770 -1320
rect 120830 -1380 120850 -1320
rect 120910 -1380 120920 -1320
rect 120680 -3000 120920 -1380
rect 121380 -1160 121620 -1150
rect 121380 -1220 121390 -1160
rect 121450 -1220 121470 -1160
rect 121530 -1220 121550 -1160
rect 121610 -1220 121620 -1160
rect 121380 -1240 121620 -1220
rect 121380 -1300 121390 -1240
rect 121450 -1300 121470 -1240
rect 121530 -1300 121550 -1240
rect 121610 -1300 121620 -1240
rect 121380 -1320 121620 -1300
rect 121380 -1380 121390 -1320
rect 121450 -1380 121470 -1320
rect 121530 -1380 121550 -1320
rect 121610 -1380 121620 -1320
rect 121380 -3000 121620 -1380
rect 122080 -1160 122320 -1150
rect 122080 -1220 122090 -1160
rect 122150 -1220 122170 -1160
rect 122230 -1220 122250 -1160
rect 122310 -1220 122320 -1160
rect 122080 -1240 122320 -1220
rect 122080 -1300 122090 -1240
rect 122150 -1300 122170 -1240
rect 122230 -1300 122250 -1240
rect 122310 -1300 122320 -1240
rect 122080 -1320 122320 -1300
rect 122080 -1380 122090 -1320
rect 122150 -1380 122170 -1320
rect 122230 -1380 122250 -1320
rect 122310 -1380 122320 -1320
rect 122080 -3000 122320 -1380
rect 122780 -1160 123020 -1150
rect 122780 -1220 122790 -1160
rect 122850 -1220 122870 -1160
rect 122930 -1220 122950 -1160
rect 123010 -1220 123020 -1160
rect 122780 -1240 123020 -1220
rect 122780 -1300 122790 -1240
rect 122850 -1300 122870 -1240
rect 122930 -1300 122950 -1240
rect 123010 -1300 123020 -1240
rect 122780 -1320 123020 -1300
rect 122780 -1380 122790 -1320
rect 122850 -1380 122870 -1320
rect 122930 -1380 122950 -1320
rect 123010 -1380 123020 -1320
rect 122780 -3000 123020 -1380
<< via1 >>
rect 104590 9280 104650 9340
rect 104670 9280 104730 9340
rect 104750 9280 104810 9340
rect 104590 9200 104650 9260
rect 104670 9200 104730 9260
rect 104750 9200 104810 9260
rect 104590 9120 104650 9180
rect 104670 9120 104730 9180
rect 104750 9120 104810 9180
rect 105290 9280 105350 9340
rect 105370 9280 105430 9340
rect 105450 9280 105510 9340
rect 105290 9200 105350 9260
rect 105370 9200 105430 9260
rect 105450 9200 105510 9260
rect 105290 9120 105350 9180
rect 105370 9120 105430 9180
rect 105450 9120 105510 9180
rect 105990 9280 106050 9340
rect 106070 9280 106130 9340
rect 106150 9280 106210 9340
rect 105990 9200 106050 9260
rect 106070 9200 106130 9260
rect 106150 9200 106210 9260
rect 105990 9120 106050 9180
rect 106070 9120 106130 9180
rect 106150 9120 106210 9180
rect 106690 9280 106750 9340
rect 106770 9280 106830 9340
rect 106850 9280 106910 9340
rect 106690 9200 106750 9260
rect 106770 9200 106830 9260
rect 106850 9200 106910 9260
rect 106690 9120 106750 9180
rect 106770 9120 106830 9180
rect 106850 9120 106910 9180
rect 109490 9970 109550 9980
rect 109490 9930 109500 9970
rect 109500 9930 109540 9970
rect 109540 9930 109550 9970
rect 109490 9920 109550 9930
rect 109610 9970 109670 9980
rect 109610 9930 109620 9970
rect 109620 9930 109660 9970
rect 109660 9930 109670 9970
rect 109610 9920 109670 9930
rect 109730 9970 109790 9980
rect 109730 9930 109740 9970
rect 109740 9930 109780 9970
rect 109780 9930 109790 9970
rect 109730 9920 109790 9930
rect 109850 9970 109910 9980
rect 109850 9930 109860 9970
rect 109860 9930 109900 9970
rect 109900 9930 109910 9970
rect 109850 9920 109910 9930
rect 109970 9970 110030 9980
rect 109970 9930 109980 9970
rect 109980 9930 110020 9970
rect 110020 9930 110030 9970
rect 109970 9920 110030 9930
rect 110090 9970 110150 9980
rect 110090 9930 110100 9970
rect 110100 9930 110140 9970
rect 110140 9930 110150 9970
rect 110090 9920 110150 9930
rect 110210 9970 110270 9980
rect 110210 9930 110220 9970
rect 110220 9930 110260 9970
rect 110260 9930 110270 9970
rect 110210 9920 110270 9930
rect 110330 9970 110390 9980
rect 110330 9930 110340 9970
rect 110340 9930 110380 9970
rect 110380 9930 110390 9970
rect 110330 9920 110390 9930
rect 110450 9970 110510 9980
rect 110450 9930 110460 9970
rect 110460 9930 110500 9970
rect 110500 9930 110510 9970
rect 110450 9920 110510 9930
rect 110570 9970 110630 9980
rect 110570 9930 110580 9970
rect 110580 9930 110620 9970
rect 110620 9930 110630 9970
rect 110570 9920 110630 9930
rect 114910 9920 114970 9980
rect 109430 9810 109490 9870
rect 109670 9810 109730 9870
rect 109910 9810 109970 9870
rect 110150 9810 110210 9870
rect 110390 9810 110450 9870
rect 110630 9810 110690 9870
rect 112220 9810 112280 9870
rect 108090 9280 108150 9340
rect 108170 9280 108230 9340
rect 108250 9280 108310 9340
rect 108090 9200 108150 9260
rect 108170 9200 108230 9260
rect 108250 9200 108310 9260
rect 108090 9120 108150 9180
rect 108170 9120 108230 9180
rect 108250 9120 108310 9180
rect 109310 9050 109370 9060
rect 109310 9010 109320 9050
rect 109320 9010 109360 9050
rect 109360 9010 109370 9050
rect 109310 9000 109370 9010
rect 109550 9000 109610 9060
rect 109790 9000 109850 9060
rect 110030 9000 110090 9060
rect 110270 9000 110330 9060
rect 110510 9000 110570 9060
rect 111980 9590 112040 9600
rect 111980 9550 111990 9590
rect 111990 9550 112030 9590
rect 112030 9550 112040 9590
rect 111980 9540 112040 9550
rect 113160 9810 113220 9870
rect 114380 9810 114440 9870
rect 112220 9540 112280 9600
rect 112340 9590 112400 9600
rect 112340 9550 112350 9590
rect 112350 9550 112390 9590
rect 112390 9550 112400 9590
rect 112340 9540 112400 9550
rect 110750 9050 110810 9060
rect 110750 9010 110760 9050
rect 110760 9010 110800 9050
rect 110800 9010 110810 9050
rect 110750 9000 110810 9010
rect 111080 9000 111140 9060
rect 111160 9000 111220 9060
rect 111240 9000 111300 9060
rect 109190 8890 109250 8950
rect 109430 8890 109490 8950
rect 109670 8890 109730 8950
rect 109910 8890 109970 8950
rect 110150 8890 110210 8950
rect 110390 8890 110450 8950
rect 110630 8890 110690 8950
rect 109190 8810 109250 8870
rect 109430 8810 109490 8870
rect 109670 8810 109730 8870
rect 109910 8810 109970 8870
rect 110150 8810 110210 8870
rect 110390 8810 110450 8870
rect 110630 8810 110690 8870
rect 109190 8730 109250 8790
rect 109430 8730 109490 8790
rect 109670 8730 109730 8790
rect 109910 8730 109970 8790
rect 110150 8730 110210 8790
rect 110390 8730 110450 8790
rect 110630 8730 110690 8790
rect 109190 8650 109250 8710
rect 109430 8650 109490 8710
rect 109670 8650 109730 8710
rect 109910 8650 109970 8710
rect 110150 8650 110210 8710
rect 110390 8650 110450 8710
rect 110630 8650 110690 8710
rect 109190 8570 109250 8630
rect 109430 8570 109490 8630
rect 109670 8570 109730 8630
rect 109910 8570 109970 8630
rect 110150 8570 110210 8630
rect 110390 8570 110450 8630
rect 110630 8570 110690 8630
rect 109190 8490 109250 8550
rect 109430 8490 109490 8550
rect 109670 8490 109730 8550
rect 109910 8490 109970 8550
rect 110150 8490 110210 8550
rect 110390 8490 110450 8550
rect 110630 8490 110690 8550
rect 109190 8410 109250 8470
rect 109430 8410 109490 8470
rect 109670 8410 109730 8470
rect 109910 8410 109970 8470
rect 110150 8410 110210 8470
rect 110390 8410 110450 8470
rect 110630 8410 110690 8470
rect 112920 9360 112980 9420
rect 112920 9280 112980 9340
rect 112920 9250 112980 9260
rect 112920 9210 112930 9250
rect 112930 9210 112970 9250
rect 112970 9210 112980 9250
rect 112920 9200 112980 9210
rect 113040 9360 113100 9420
rect 113040 9280 113100 9340
rect 113040 9200 113100 9260
rect 113690 9700 113750 9760
rect 113770 9700 113830 9760
rect 113850 9700 113910 9760
rect 113690 9620 113750 9680
rect 113770 9620 113830 9680
rect 113850 9620 113910 9680
rect 113690 9540 113750 9600
rect 113770 9540 113830 9600
rect 113850 9540 113910 9600
rect 113280 9360 113340 9420
rect 113280 9280 113340 9340
rect 113280 9250 113340 9260
rect 113280 9210 113290 9250
rect 113290 9210 113330 9250
rect 113330 9210 113340 9250
rect 113280 9200 113340 9210
rect 114260 9700 114320 9760
rect 114260 9620 114320 9680
rect 114260 9590 114320 9600
rect 114260 9550 114270 9590
rect 114270 9550 114310 9590
rect 114310 9550 114320 9590
rect 114260 9540 114320 9550
rect 113690 9360 113750 9420
rect 113770 9360 113830 9420
rect 113850 9360 113910 9420
rect 113690 9280 113750 9340
rect 113770 9280 113830 9340
rect 113850 9280 113910 9340
rect 113690 9200 113750 9260
rect 113770 9200 113830 9260
rect 113850 9200 113910 9260
rect 112220 8730 112280 8790
rect 113160 8730 113220 8790
rect 111350 8620 111410 8680
rect 112110 8670 112170 8680
rect 112110 8630 112120 8670
rect 112120 8630 112160 8670
rect 112160 8630 112170 8670
rect 112110 8620 112170 8630
rect 113060 8670 113120 8680
rect 113060 8630 113070 8670
rect 113070 8630 113110 8670
rect 113110 8630 113120 8670
rect 113060 8620 113120 8630
rect 111080 8400 111140 8460
rect 111160 8400 111220 8460
rect 111240 8400 111300 8460
rect 109310 8290 109370 8350
rect 108090 7290 108150 7350
rect 108170 7290 108230 7350
rect 108250 7290 108310 7350
rect 108090 7210 108150 7270
rect 108170 7210 108230 7270
rect 108250 7210 108310 7270
rect 108090 7130 108150 7190
rect 108170 7130 108230 7190
rect 108250 7130 108310 7190
rect 108520 7610 108580 7670
rect 109550 8290 109610 8350
rect 109790 8290 109850 8350
rect 110030 8290 110090 8350
rect 110270 8290 110330 8350
rect 110510 8290 110570 8350
rect 111080 8320 111140 8380
rect 111160 8320 111220 8380
rect 111240 8320 111300 8380
rect 111080 8240 111140 8300
rect 111160 8240 111220 8300
rect 111240 8240 111300 8300
rect 109310 7510 109370 7570
rect 109550 7510 109610 7570
rect 109790 7510 109850 7570
rect 110030 7510 110090 7570
rect 110270 7510 110330 7570
rect 110510 7510 110570 7570
rect 110810 7510 110870 7570
rect 110890 7510 110950 7570
rect 110970 7510 111030 7570
rect 109370 7450 109430 7460
rect 109370 7410 109380 7450
rect 109380 7410 109420 7450
rect 109420 7410 109430 7450
rect 109370 7400 109430 7410
rect 109490 7450 109550 7460
rect 109490 7410 109500 7450
rect 109500 7410 109540 7450
rect 109540 7410 109550 7450
rect 109490 7400 109550 7410
rect 109610 7450 109670 7460
rect 109610 7410 109620 7450
rect 109620 7410 109660 7450
rect 109660 7410 109670 7450
rect 109610 7400 109670 7410
rect 109730 7450 109790 7460
rect 109730 7410 109740 7450
rect 109740 7410 109780 7450
rect 109780 7410 109790 7450
rect 109730 7400 109790 7410
rect 109850 7450 109910 7460
rect 109850 7410 109860 7450
rect 109860 7410 109900 7450
rect 109900 7410 109910 7450
rect 109850 7400 109910 7410
rect 109970 7450 110030 7460
rect 109970 7410 109980 7450
rect 109980 7410 110020 7450
rect 110020 7410 110030 7450
rect 109970 7400 110030 7410
rect 110090 7450 110150 7460
rect 110090 7410 110100 7450
rect 110100 7410 110140 7450
rect 110140 7410 110150 7450
rect 110090 7400 110150 7410
rect 110210 7450 110270 7460
rect 110210 7410 110220 7450
rect 110220 7410 110260 7450
rect 110260 7410 110270 7450
rect 110210 7400 110270 7410
rect 110330 7450 110390 7460
rect 110330 7410 110340 7450
rect 110340 7410 110380 7450
rect 110380 7410 110390 7450
rect 110330 7400 110390 7410
rect 110450 7450 110510 7460
rect 110450 7410 110460 7450
rect 110460 7410 110500 7450
rect 110500 7410 110510 7450
rect 110450 7400 110510 7410
rect 109250 7290 109310 7350
rect 109250 7210 109310 7270
rect 109250 7130 109310 7190
rect 109470 7290 109530 7350
rect 109470 7210 109530 7270
rect 109470 7130 109530 7190
rect 109690 7290 109750 7350
rect 109690 7210 109750 7270
rect 109690 7130 109750 7190
rect 109910 7290 109970 7350
rect 109910 7210 109970 7270
rect 109910 7130 109970 7190
rect 110130 7290 110190 7350
rect 110130 7210 110190 7270
rect 110130 7130 110190 7190
rect 110350 7290 110410 7350
rect 110350 7210 110410 7270
rect 110350 7130 110410 7190
rect 110570 7290 110630 7350
rect 110570 7210 110630 7270
rect 110570 7130 110630 7190
rect 109360 6940 109420 7000
rect 109580 6940 109640 7000
rect 109800 6940 109860 7000
rect 110020 6940 110080 7000
rect 110240 6940 110300 7000
rect 110460 6940 110520 7000
rect 110810 6900 110870 6960
rect 110890 6900 110950 6960
rect 110970 6900 111030 6960
rect 110810 6820 110870 6880
rect 110890 6820 110950 6880
rect 110970 6820 111030 6880
rect 110810 6740 110870 6800
rect 110890 6740 110950 6800
rect 110970 6740 111030 6800
rect 108440 5500 108500 5560
rect 108520 5500 108580 5560
rect 108600 5500 108660 5560
rect 108440 5420 108500 5480
rect 108520 5420 108580 5480
rect 108600 5420 108660 5480
rect 108440 5340 108500 5400
rect 108520 5340 108580 5400
rect 108600 5340 108660 5400
rect 109360 5660 109420 5720
rect 109580 5660 109640 5720
rect 109800 5660 109860 5720
rect 110020 5660 110080 5720
rect 109910 5550 109970 5560
rect 109910 5510 109920 5550
rect 109920 5510 109960 5550
rect 109960 5510 109970 5550
rect 109910 5500 109970 5510
rect 109910 5470 109970 5480
rect 109910 5430 109920 5470
rect 109920 5430 109960 5470
rect 109960 5430 109970 5470
rect 109910 5420 109970 5430
rect 109910 5390 109970 5400
rect 109910 5350 109920 5390
rect 109920 5350 109960 5390
rect 109960 5350 109970 5390
rect 109910 5340 109970 5350
rect 110240 5660 110300 5720
rect 110460 5660 110520 5720
rect 107990 5200 108050 5260
rect 108070 5200 108130 5260
rect 108160 5200 108220 5260
rect 108240 5200 108300 5260
rect 108330 5200 108390 5260
rect 108410 5200 108470 5260
rect 107990 5120 108050 5180
rect 108070 5120 108130 5180
rect 108160 5120 108220 5180
rect 108240 5120 108300 5180
rect 108330 5120 108390 5180
rect 108410 5120 108470 5180
rect 107990 5040 108050 5100
rect 108070 5040 108130 5100
rect 108160 5040 108220 5100
rect 108240 5040 108300 5100
rect 108330 5040 108390 5100
rect 108410 5040 108470 5100
rect 107690 4660 107750 4720
rect 107770 4660 107830 4720
rect 107850 4660 107910 4720
rect 107690 4580 107750 4640
rect 107770 4580 107830 4640
rect 107850 4580 107910 4640
rect 107690 4500 107750 4560
rect 107770 4500 107830 4560
rect 107850 4500 107910 4560
rect 107690 2440 107750 2500
rect 107770 2440 107830 2500
rect 107850 2440 107910 2500
rect 107690 2360 107750 2420
rect 107770 2360 107830 2420
rect 107850 2360 107910 2420
rect 107690 2280 107750 2340
rect 107770 2280 107830 2340
rect 107850 2280 107910 2340
rect 104590 -1220 104650 -1160
rect 104670 -1220 104730 -1160
rect 104750 -1220 104810 -1160
rect 104590 -1300 104650 -1240
rect 104670 -1300 104730 -1240
rect 104750 -1300 104810 -1240
rect 104590 -1380 104650 -1320
rect 104670 -1380 104730 -1320
rect 104750 -1380 104810 -1320
rect 105290 -1220 105350 -1160
rect 105370 -1220 105430 -1160
rect 105450 -1220 105510 -1160
rect 105290 -1300 105350 -1240
rect 105370 -1300 105430 -1240
rect 105450 -1300 105510 -1240
rect 105290 -1380 105350 -1320
rect 105370 -1380 105430 -1320
rect 105450 -1380 105510 -1320
rect 105990 -1220 106050 -1160
rect 106070 -1220 106130 -1160
rect 106150 -1220 106210 -1160
rect 105990 -1300 106050 -1240
rect 106070 -1300 106130 -1240
rect 106150 -1300 106210 -1240
rect 105990 -1380 106050 -1320
rect 106070 -1380 106130 -1320
rect 106150 -1380 106210 -1320
rect 106690 -1220 106750 -1160
rect 106770 -1220 106830 -1160
rect 106850 -1220 106910 -1160
rect 106690 -1300 106750 -1240
rect 106770 -1300 106830 -1240
rect 106850 -1300 106910 -1240
rect 106690 -1380 106750 -1320
rect 106770 -1380 106830 -1320
rect 106850 -1380 106910 -1320
rect 107390 -1220 107450 -1160
rect 107470 -1220 107530 -1160
rect 107550 -1220 107610 -1160
rect 107390 -1300 107450 -1240
rect 107470 -1300 107530 -1240
rect 107550 -1300 107610 -1240
rect 107390 -1380 107450 -1320
rect 107470 -1380 107530 -1320
rect 107550 -1380 107610 -1320
rect 109360 5200 109420 5260
rect 109470 5200 109530 5260
rect 109580 5200 109640 5260
rect 109690 5200 109750 5260
rect 109800 5200 109860 5260
rect 109910 5200 109970 5260
rect 110020 5200 110080 5260
rect 110130 5200 110190 5260
rect 110240 5200 110300 5260
rect 110350 5200 110410 5260
rect 110460 5200 110520 5260
rect 109360 5120 109420 5180
rect 109470 5120 109530 5180
rect 109580 5120 109640 5180
rect 109690 5120 109750 5180
rect 109800 5120 109860 5180
rect 109910 5120 109970 5180
rect 110020 5120 110080 5180
rect 110130 5120 110190 5180
rect 110240 5120 110300 5180
rect 110350 5120 110410 5180
rect 110460 5120 110520 5180
rect 109360 5040 109420 5100
rect 109470 5040 109530 5100
rect 109580 5040 109640 5100
rect 109690 5040 109750 5100
rect 109800 5040 109860 5100
rect 109910 5040 109970 5100
rect 110020 5040 110080 5100
rect 110130 5040 110190 5100
rect 110240 5040 110300 5100
rect 110350 5040 110410 5100
rect 110460 5040 110520 5100
rect 110810 5500 110870 5560
rect 110890 5500 110950 5560
rect 110970 5500 111030 5560
rect 110810 5420 110870 5480
rect 110890 5420 110950 5480
rect 110970 5420 111030 5480
rect 110810 5340 110870 5400
rect 110890 5340 110950 5400
rect 110970 5340 111030 5400
rect 109250 4930 109310 4990
rect 109250 4850 109310 4910
rect 109250 4770 109310 4830
rect 110570 4930 110630 4990
rect 110570 4850 110630 4910
rect 110570 4770 110630 4830
rect 108000 4060 108060 4120
rect 108100 4060 108160 4120
rect 108200 4060 108260 4120
rect 108300 4060 108360 4120
rect 108400 4060 108460 4120
rect 108000 3960 108060 4020
rect 108100 3960 108160 4020
rect 108200 3960 108260 4020
rect 108300 3960 108360 4020
rect 108400 3960 108460 4020
rect 109360 4660 109420 4720
rect 109360 4580 109420 4640
rect 109360 4500 109420 4560
rect 109580 4660 109640 4720
rect 109580 4580 109640 4640
rect 109580 4500 109640 4560
rect 109800 4660 109860 4720
rect 109800 4580 109860 4640
rect 109800 4500 109860 4560
rect 110020 4660 110080 4720
rect 110020 4580 110080 4640
rect 110020 4500 110080 4560
rect 110240 4660 110300 4720
rect 110240 4580 110300 4640
rect 110240 4500 110300 4560
rect 110460 4660 110520 4720
rect 110460 4580 110520 4640
rect 110460 4500 110520 4560
rect 109470 4390 109530 4450
rect 109690 4390 109750 4450
rect 109910 4390 109970 4450
rect 110130 4390 110190 4450
rect 110350 4390 110410 4450
rect 108000 3860 108060 3920
rect 108100 3860 108160 3920
rect 108200 3860 108260 3920
rect 108300 3860 108360 3920
rect 108400 3860 108460 3920
rect 108980 3880 109040 3940
rect 109470 3930 109530 3940
rect 109470 3890 109480 3930
rect 109480 3890 109520 3930
rect 109520 3890 109530 3930
rect 109470 3880 109530 3890
rect 109690 3930 109750 3940
rect 109690 3890 109700 3930
rect 109700 3890 109740 3930
rect 109740 3890 109750 3930
rect 109690 3880 109750 3890
rect 109910 3930 109970 3940
rect 109910 3890 109920 3930
rect 109920 3890 109960 3930
rect 109960 3890 109970 3930
rect 109910 3880 109970 3890
rect 110130 3930 110190 3940
rect 110130 3890 110140 3930
rect 110140 3890 110180 3930
rect 110180 3890 110190 3930
rect 110130 3880 110190 3890
rect 110350 3930 110410 3940
rect 110350 3890 110360 3930
rect 110360 3890 110400 3930
rect 110400 3890 110410 3930
rect 110350 3880 110410 3890
rect 108510 2930 108580 2940
rect 108510 2880 108520 2930
rect 108520 2880 108570 2930
rect 108570 2880 108580 2930
rect 108510 2870 108580 2880
rect 108630 2930 108700 2940
rect 108630 2880 108640 2930
rect 108640 2880 108690 2930
rect 108690 2880 108700 2930
rect 108630 2870 108700 2880
rect 108750 2930 108820 2940
rect 108750 2880 108760 2930
rect 108760 2880 108810 2930
rect 108810 2880 108820 2930
rect 108750 2870 108820 2880
rect 108870 2930 108940 2940
rect 108870 2880 108880 2930
rect 108880 2880 108930 2930
rect 108930 2880 108940 2930
rect 108870 2870 108940 2880
rect 110240 3800 110300 3810
rect 110240 3760 110250 3800
rect 110250 3760 110290 3800
rect 110290 3760 110300 3800
rect 110240 3750 110300 3760
rect 110240 3720 110300 3730
rect 110240 3680 110250 3720
rect 110250 3680 110290 3720
rect 110290 3680 110300 3720
rect 110240 3670 110300 3680
rect 110810 3750 110870 3810
rect 110890 3750 110950 3810
rect 110970 3750 111030 3810
rect 110810 3670 110870 3730
rect 110890 3670 110950 3730
rect 110970 3670 111030 3730
rect 109070 3510 109130 3570
rect 109470 3510 109530 3570
rect 109690 3510 109750 3570
rect 109910 3510 109970 3570
rect 110130 3510 110190 3570
rect 110350 3510 110410 3570
rect 109070 2870 109130 2930
rect 108760 2730 108820 2790
rect 108980 2730 109040 2790
rect 109470 2830 109530 2890
rect 109690 2830 109750 2890
rect 109910 2830 109970 2890
rect 110130 2830 110190 2890
rect 110350 2830 110410 2890
rect 110810 2990 110870 3050
rect 110890 2990 110950 3050
rect 110970 2990 111030 3050
rect 110810 2910 110870 2970
rect 110890 2910 110950 2970
rect 110970 2910 111030 2970
rect 110810 2830 110870 2890
rect 110890 2830 110950 2890
rect 110970 2830 111030 2890
rect 113030 8400 113090 8460
rect 113030 8320 113090 8380
rect 113030 8290 113090 8300
rect 113030 8250 113040 8290
rect 113040 8250 113080 8290
rect 113080 8250 113090 8290
rect 113030 8240 113090 8250
rect 113360 8400 113420 8460
rect 113360 8320 113420 8380
rect 113360 8290 113420 8300
rect 113360 8250 113370 8290
rect 113370 8250 113410 8290
rect 113410 8250 113420 8290
rect 113360 8240 113420 8250
rect 114500 9700 114560 9760
rect 114500 9620 114560 9680
rect 114500 9540 114560 9600
rect 114620 9700 114680 9760
rect 114620 9620 114680 9680
rect 114620 9590 114680 9600
rect 114620 9550 114630 9590
rect 114630 9550 114670 9590
rect 114670 9550 114680 9590
rect 114620 9540 114680 9550
rect 114380 8730 114440 8790
rect 114480 8510 114540 8570
rect 116970 9970 117030 9980
rect 116970 9930 116980 9970
rect 116980 9930 117020 9970
rect 117020 9930 117030 9970
rect 116970 9920 117030 9930
rect 117090 9970 117150 9980
rect 117090 9930 117100 9970
rect 117100 9930 117140 9970
rect 117140 9930 117150 9970
rect 117090 9920 117150 9930
rect 117210 9970 117270 9980
rect 117210 9930 117220 9970
rect 117220 9930 117260 9970
rect 117260 9930 117270 9970
rect 117210 9920 117270 9930
rect 117330 9970 117390 9980
rect 117330 9930 117340 9970
rect 117340 9930 117380 9970
rect 117380 9930 117390 9970
rect 117330 9920 117390 9930
rect 117450 9970 117510 9980
rect 117450 9930 117460 9970
rect 117460 9930 117500 9970
rect 117500 9930 117510 9970
rect 117450 9920 117510 9930
rect 117570 9970 117630 9980
rect 117570 9930 117580 9970
rect 117580 9930 117620 9970
rect 117620 9930 117630 9970
rect 117570 9920 117630 9930
rect 117690 9970 117750 9980
rect 117690 9930 117700 9970
rect 117700 9930 117740 9970
rect 117740 9930 117750 9970
rect 117690 9920 117750 9930
rect 117810 9970 117870 9980
rect 117810 9930 117820 9970
rect 117820 9930 117860 9970
rect 117860 9930 117870 9970
rect 117810 9920 117870 9930
rect 117930 9970 117990 9980
rect 117930 9930 117940 9970
rect 117940 9930 117980 9970
rect 117980 9930 117990 9970
rect 117930 9920 117990 9930
rect 118050 9970 118110 9980
rect 118050 9930 118060 9970
rect 118060 9930 118100 9970
rect 118100 9930 118110 9970
rect 118050 9920 118110 9930
rect 115320 9810 115380 9870
rect 115200 9590 115260 9600
rect 115200 9550 115210 9590
rect 115210 9550 115250 9590
rect 115250 9550 115260 9590
rect 115200 9540 115260 9550
rect 116910 9810 116970 9870
rect 117150 9810 117210 9870
rect 117390 9810 117450 9870
rect 117630 9810 117690 9870
rect 117870 9810 117930 9870
rect 118110 9810 118170 9870
rect 115320 9540 115380 9600
rect 115560 9590 115620 9600
rect 115560 9550 115570 9590
rect 115570 9550 115610 9590
rect 115610 9550 115620 9590
rect 115560 9540 115620 9550
rect 115320 8730 115380 8790
rect 115352 8670 115412 8680
rect 115352 8630 115362 8670
rect 115362 8630 115402 8670
rect 115402 8630 115412 8670
rect 115352 8620 115412 8630
rect 116300 9000 116360 9060
rect 116380 9000 116440 9060
rect 116460 9000 116520 9060
rect 116190 8620 116250 8680
rect 114910 8510 114970 8570
rect 115440 8510 115500 8570
rect 113690 8400 113750 8460
rect 113850 8400 113910 8460
rect 113690 8320 113750 8380
rect 113850 8320 113910 8380
rect 113690 8290 113750 8300
rect 113690 8250 113700 8290
rect 113700 8250 113740 8290
rect 113740 8250 113750 8290
rect 113690 8240 113750 8250
rect 113850 8290 113910 8300
rect 113850 8250 113860 8290
rect 113860 8250 113900 8290
rect 113900 8250 113910 8290
rect 113850 8240 113910 8250
rect 114180 8400 114240 8460
rect 114180 8320 114240 8380
rect 114180 8290 114240 8300
rect 114180 8250 114190 8290
rect 114190 8250 114230 8290
rect 114230 8250 114240 8290
rect 114180 8240 114240 8250
rect 114510 8400 114570 8460
rect 114510 8320 114570 8380
rect 114510 8290 114570 8300
rect 114510 8250 114520 8290
rect 114520 8250 114560 8290
rect 114560 8250 114570 8290
rect 114510 8240 114570 8250
rect 113250 8160 113310 8170
rect 113250 8120 113260 8160
rect 113260 8120 113300 8160
rect 113300 8120 113310 8160
rect 113250 8110 113310 8120
rect 113470 8160 113530 8170
rect 113470 8120 113480 8160
rect 113480 8120 113520 8160
rect 113520 8120 113530 8160
rect 113470 8110 113530 8120
rect 114070 8160 114130 8170
rect 114070 8120 114080 8160
rect 114080 8120 114120 8160
rect 114120 8120 114130 8160
rect 114070 8110 114130 8120
rect 114290 8160 114350 8170
rect 114290 8120 114300 8160
rect 114300 8120 114340 8160
rect 114340 8120 114350 8160
rect 114290 8110 114350 8120
rect 113120 7540 113180 7550
rect 113600 7540 113660 7550
rect 113120 7500 113130 7540
rect 113130 7500 113170 7540
rect 113170 7500 113180 7540
rect 113120 7490 113180 7500
rect 113360 7520 113420 7530
rect 113360 7480 113370 7520
rect 113370 7480 113410 7520
rect 113410 7480 113420 7520
rect 113360 7470 113420 7480
rect 113600 7500 113610 7540
rect 113610 7500 113650 7540
rect 113650 7500 113660 7540
rect 113600 7490 113660 7500
rect 111350 7400 111410 7460
rect 111080 7290 111140 7350
rect 111160 7290 111220 7350
rect 111240 7290 111300 7350
rect 113210 7400 113270 7410
rect 113210 7360 113220 7400
rect 113220 7360 113260 7400
rect 113260 7360 113270 7400
rect 113210 7350 113270 7360
rect 111080 7210 111140 7270
rect 111160 7210 111220 7270
rect 111240 7210 111300 7270
rect 111080 7130 111140 7190
rect 111160 7130 111220 7190
rect 111240 7130 111300 7190
rect 111910 7230 111970 7290
rect 113500 7230 113560 7290
rect 111080 4930 111140 4990
rect 111160 4930 111220 4990
rect 111240 4930 111300 4990
rect 111080 4850 111140 4910
rect 111160 4850 111220 4910
rect 111240 4850 111300 4910
rect 111080 4770 111140 4830
rect 111160 4770 111220 4830
rect 111240 4770 111300 4830
rect 109360 2720 109420 2780
rect 109360 2640 109420 2700
rect 109360 2560 109420 2620
rect 109580 2720 109640 2780
rect 109580 2640 109640 2700
rect 109580 2560 109640 2620
rect 109800 2720 109860 2780
rect 109800 2640 109860 2700
rect 109800 2560 109860 2620
rect 110020 2720 110080 2780
rect 110020 2640 110080 2700
rect 110020 2560 110080 2620
rect 110240 2720 110300 2780
rect 110240 2640 110300 2700
rect 110240 2560 110300 2620
rect 110460 2720 110520 2780
rect 110460 2640 110520 2700
rect 110460 2560 110520 2620
rect 111350 6260 111410 6320
rect 111430 6260 111490 6320
rect 111510 6260 111570 6320
rect 111350 6180 111410 6240
rect 111430 6180 111490 6240
rect 111510 6180 111570 6240
rect 111350 6100 111410 6160
rect 111430 6100 111490 6160
rect 111510 6100 111570 6160
rect 111350 5960 111410 6020
rect 111430 5960 111490 6020
rect 111510 5960 111570 6020
rect 111350 5880 111410 5940
rect 111430 5880 111490 5940
rect 111510 5880 111570 5940
rect 111350 5800 111410 5860
rect 111430 5800 111490 5860
rect 111510 5800 111570 5860
rect 111350 5140 111410 5200
rect 111430 5140 111490 5200
rect 111510 5140 111570 5200
rect 111350 5060 111410 5120
rect 111430 5060 111490 5120
rect 111510 5060 111570 5120
rect 111350 4980 111410 5040
rect 111430 4980 111490 5040
rect 111510 4980 111570 5040
rect 111350 4660 111410 4720
rect 111430 4660 111490 4720
rect 111510 4660 111570 4720
rect 111350 4580 111410 4640
rect 111430 4580 111490 4640
rect 111510 4580 111570 4640
rect 111350 4500 111410 4560
rect 111430 4500 111490 4560
rect 111510 4500 111570 4560
rect 111700 5770 111760 5830
rect 111080 2720 111140 2780
rect 111160 2720 111220 2780
rect 111240 2720 111300 2780
rect 111080 2640 111140 2700
rect 111160 2640 111220 2700
rect 111240 2640 111300 2700
rect 111080 2560 111140 2620
rect 111160 2560 111220 2620
rect 111240 2560 111300 2620
rect 111350 4330 111410 4390
rect 111430 4330 111490 4390
rect 111510 4330 111570 4390
rect 111350 4250 111410 4310
rect 111430 4250 111490 4310
rect 111510 4250 111570 4310
rect 111350 4170 111410 4230
rect 111430 4170 111490 4230
rect 111510 4170 111570 4230
rect 109250 2440 109310 2500
rect 109250 2360 109310 2420
rect 109250 2280 109310 2340
rect 110570 2440 110630 2500
rect 110570 2360 110630 2420
rect 110570 2280 110630 2340
rect 108520 2170 108580 2230
rect 107990 1680 108050 1740
rect 108070 1680 108130 1740
rect 108160 1680 108220 1740
rect 108240 1680 108300 1740
rect 108330 1680 108390 1740
rect 108410 1680 108470 1740
rect 107990 1600 108050 1660
rect 108070 1600 108130 1660
rect 108160 1600 108220 1660
rect 108240 1600 108300 1660
rect 108330 1600 108390 1660
rect 108410 1600 108470 1660
rect 107990 1520 108050 1580
rect 108070 1520 108130 1580
rect 108160 1520 108220 1580
rect 108240 1520 108300 1580
rect 108330 1520 108390 1580
rect 108410 1520 108470 1580
rect 108650 1790 108710 1850
rect 108650 1410 108710 1470
rect 108650 1350 108720 1360
rect 108650 1300 108660 1350
rect 108660 1300 108710 1350
rect 108710 1300 108720 1350
rect 108650 1290 108720 1300
rect 108780 1680 108840 1740
rect 108780 1600 108840 1660
rect 108780 1520 108840 1580
rect 109510 1680 109570 1740
rect 109590 1680 109650 1740
rect 109670 1680 109730 1740
rect 109750 1680 109810 1740
rect 109830 1680 109890 1740
rect 109910 1680 109970 1740
rect 109990 1680 110050 1740
rect 110070 1680 110130 1740
rect 110150 1680 110210 1740
rect 110230 1680 110290 1740
rect 110310 1680 110370 1740
rect 109510 1600 109570 1660
rect 109590 1600 109650 1660
rect 109670 1600 109730 1660
rect 109750 1600 109810 1660
rect 109830 1600 109890 1660
rect 109910 1600 109970 1660
rect 109990 1600 110050 1660
rect 110070 1600 110130 1660
rect 110150 1600 110210 1660
rect 110230 1600 110290 1660
rect 110310 1600 110370 1660
rect 109510 1520 109570 1580
rect 109590 1520 109650 1580
rect 109670 1520 109730 1580
rect 109750 1520 109810 1580
rect 109830 1520 109890 1580
rect 109910 1520 109970 1580
rect 109990 1520 110050 1580
rect 110070 1520 110130 1580
rect 110150 1520 110210 1580
rect 110230 1520 110290 1580
rect 110310 1520 110370 1580
rect 108770 1350 108840 1360
rect 108770 1300 108780 1350
rect 108780 1300 108830 1350
rect 108830 1300 108840 1350
rect 108770 1290 108840 1300
rect 109610 1460 109670 1470
rect 109610 1420 109620 1460
rect 109620 1420 109660 1460
rect 109660 1420 109670 1460
rect 109610 1410 109670 1420
rect 109810 1460 109870 1470
rect 109810 1420 109820 1460
rect 109820 1420 109860 1460
rect 109860 1420 109870 1460
rect 109810 1410 109870 1420
rect 109510 -90 109570 -30
rect 110010 1460 110070 1470
rect 110010 1420 110020 1460
rect 110020 1420 110060 1460
rect 110060 1420 110070 1460
rect 110010 1410 110070 1420
rect 110210 1460 110270 1470
rect 110210 1420 110220 1460
rect 110220 1420 110260 1460
rect 110260 1420 110270 1460
rect 110210 1410 110270 1420
rect 109910 -90 109970 -30
rect 107690 -1220 107750 -1160
rect 107770 -1220 107830 -1160
rect 107850 -1220 107910 -1160
rect 107690 -1300 107750 -1240
rect 107770 -1300 107830 -1240
rect 107850 -1300 107910 -1240
rect 107690 -1380 107750 -1320
rect 107770 -1380 107830 -1320
rect 107850 -1380 107910 -1320
rect 108090 -1220 108150 -1160
rect 108170 -1220 108230 -1160
rect 108250 -1220 108310 -1160
rect 108090 -1300 108150 -1240
rect 108170 -1300 108230 -1240
rect 108250 -1300 108310 -1240
rect 108090 -1380 108150 -1320
rect 108170 -1380 108230 -1320
rect 108250 -1380 108310 -1320
rect 108790 -1220 108850 -1160
rect 108870 -1220 108930 -1160
rect 108950 -1220 109010 -1160
rect 108790 -1300 108850 -1240
rect 108870 -1300 108930 -1240
rect 108950 -1300 109010 -1240
rect 108790 -1380 108850 -1320
rect 108870 -1380 108930 -1320
rect 108950 -1380 109010 -1320
rect 109310 -1220 109370 -1160
rect 109310 -1300 109370 -1240
rect 109310 -1380 109370 -1320
rect 109490 -1220 109550 -1160
rect 109570 -1220 109630 -1160
rect 109650 -1220 109710 -1160
rect 109490 -1300 109550 -1240
rect 109570 -1300 109630 -1240
rect 109650 -1300 109710 -1240
rect 109490 -1380 109550 -1320
rect 109570 -1380 109630 -1320
rect 109650 -1380 109710 -1320
rect 111350 520 111410 580
rect 111430 520 111490 580
rect 111510 520 111570 580
rect 111350 440 111410 500
rect 111430 440 111490 500
rect 111510 440 111570 500
rect 111350 360 111410 420
rect 111430 360 111490 420
rect 111510 360 111570 420
rect 114180 7520 114240 7530
rect 114180 7480 114190 7520
rect 114190 7480 114230 7520
rect 114230 7480 114240 7520
rect 114180 7470 114240 7480
rect 114330 7400 114390 7410
rect 114330 7360 114340 7400
rect 114340 7360 114380 7400
rect 114380 7360 114390 7400
rect 114330 7350 114390 7360
rect 114040 7230 114100 7290
rect 113710 7120 113770 7180
rect 113930 7120 113990 7180
rect 116790 9050 116850 9060
rect 116790 9010 116800 9050
rect 116800 9010 116840 9050
rect 116840 9010 116850 9050
rect 116790 9000 116850 9010
rect 117030 9000 117090 9060
rect 117270 9000 117330 9060
rect 117510 9000 117570 9060
rect 117750 9000 117810 9060
rect 117990 9000 118050 9060
rect 119290 9280 119350 9340
rect 119370 9280 119430 9340
rect 119450 9280 119510 9340
rect 119290 9200 119350 9260
rect 119370 9200 119430 9260
rect 119450 9200 119510 9260
rect 119290 9120 119350 9180
rect 119370 9120 119430 9180
rect 119450 9120 119510 9180
rect 118230 9050 118290 9060
rect 118230 9010 118240 9050
rect 118240 9010 118280 9050
rect 118280 9010 118290 9050
rect 118230 9000 118290 9010
rect 116300 8400 116360 8460
rect 116380 8400 116440 8460
rect 116460 8400 116520 8460
rect 116910 8890 116970 8950
rect 117150 8890 117210 8950
rect 117390 8890 117450 8950
rect 117630 8890 117690 8950
rect 117870 8890 117930 8950
rect 118110 8890 118170 8950
rect 118350 8890 118410 8950
rect 116910 8810 116970 8870
rect 117150 8810 117210 8870
rect 117390 8810 117450 8870
rect 117630 8810 117690 8870
rect 117870 8810 117930 8870
rect 118110 8810 118170 8870
rect 118350 8810 118410 8870
rect 116910 8730 116970 8790
rect 117150 8730 117210 8790
rect 117390 8730 117450 8790
rect 117630 8730 117690 8790
rect 117870 8730 117930 8790
rect 118110 8730 118170 8790
rect 118350 8730 118410 8790
rect 116910 8650 116970 8710
rect 117150 8650 117210 8710
rect 117390 8650 117450 8710
rect 117630 8650 117690 8710
rect 117870 8650 117930 8710
rect 118110 8650 118170 8710
rect 118350 8650 118410 8710
rect 116910 8570 116970 8630
rect 117150 8570 117210 8630
rect 117390 8570 117450 8630
rect 117630 8570 117690 8630
rect 117870 8570 117930 8630
rect 118110 8570 118170 8630
rect 118350 8570 118410 8630
rect 116910 8490 116970 8550
rect 117150 8490 117210 8550
rect 117390 8490 117450 8550
rect 117630 8490 117690 8550
rect 117870 8490 117930 8550
rect 118110 8490 118170 8550
rect 118350 8490 118410 8550
rect 116910 8410 116970 8470
rect 117150 8410 117210 8470
rect 117390 8410 117450 8470
rect 117630 8410 117690 8470
rect 117870 8410 117930 8470
rect 118110 8410 118170 8470
rect 118350 8410 118410 8470
rect 116300 8320 116360 8380
rect 116380 8320 116440 8380
rect 116460 8320 116520 8380
rect 116300 8240 116360 8300
rect 116380 8240 116440 8300
rect 116460 8240 116520 8300
rect 116190 7400 116250 7460
rect 117030 8290 117090 8350
rect 117270 8290 117330 8350
rect 117510 8290 117570 8350
rect 117750 8290 117810 8350
rect 117990 8290 118050 8350
rect 118230 8290 118290 8350
rect 119020 7610 119080 7670
rect 115640 7230 115700 7290
rect 116300 7290 116360 7350
rect 116380 7290 116440 7350
rect 116460 7290 116520 7350
rect 113880 7010 113940 7070
rect 114430 7010 114490 7070
rect 112180 6900 112240 6960
rect 112290 6900 112350 6960
rect 112400 6900 112460 6960
rect 112510 6900 112570 6960
rect 112620 6900 112680 6960
rect 112730 6900 112790 6960
rect 112840 6900 112900 6960
rect 112950 6900 113010 6960
rect 113060 6900 113120 6960
rect 113170 6900 113230 6960
rect 113280 6900 113340 6960
rect 112180 6820 112240 6880
rect 112290 6820 112350 6880
rect 112400 6820 112460 6880
rect 112510 6820 112570 6880
rect 112620 6820 112680 6880
rect 112730 6820 112790 6880
rect 112840 6820 112900 6880
rect 112950 6820 113010 6880
rect 113060 6820 113120 6880
rect 113170 6820 113230 6880
rect 113280 6820 113340 6880
rect 113710 6950 113770 6960
rect 113710 6910 113720 6950
rect 113720 6910 113760 6950
rect 113760 6910 113770 6950
rect 113710 6900 113770 6910
rect 114260 6900 114320 6960
rect 114370 6900 114430 6960
rect 114480 6900 114540 6960
rect 114590 6900 114650 6960
rect 114700 6900 114760 6960
rect 114810 6900 114870 6960
rect 114920 6900 114980 6960
rect 115030 6900 115090 6960
rect 115140 6900 115200 6960
rect 115250 6900 115310 6960
rect 115360 6900 115420 6960
rect 112180 6740 112240 6800
rect 112290 6740 112350 6800
rect 112400 6740 112460 6800
rect 112510 6740 112570 6800
rect 112620 6740 112680 6800
rect 112730 6740 112790 6800
rect 112840 6740 112900 6800
rect 112950 6740 113010 6800
rect 113060 6740 113120 6800
rect 113170 6740 113230 6800
rect 113280 6740 113340 6800
rect 112180 5880 112240 5940
rect 112400 5880 112460 5940
rect 112620 5880 112680 5940
rect 112840 5880 112900 5940
rect 113060 5880 113120 5940
rect 114260 6820 114320 6880
rect 114370 6820 114430 6880
rect 114480 6820 114540 6880
rect 114590 6820 114650 6880
rect 114700 6820 114760 6880
rect 114810 6820 114870 6880
rect 114920 6820 114980 6880
rect 115030 6820 115090 6880
rect 115140 6820 115200 6880
rect 115250 6820 115310 6880
rect 115360 6820 115420 6880
rect 114260 6740 114320 6800
rect 114370 6740 114430 6800
rect 114480 6740 114540 6800
rect 114590 6740 114650 6800
rect 114700 6740 114760 6800
rect 114810 6740 114870 6800
rect 114920 6740 114980 6800
rect 115030 6740 115090 6800
rect 115140 6740 115200 6800
rect 115250 6740 115310 6800
rect 115360 6740 115420 6800
rect 113550 6310 113610 6320
rect 113550 6270 113560 6310
rect 113560 6270 113600 6310
rect 113600 6270 113610 6310
rect 113550 6260 113610 6270
rect 113550 6180 113610 6240
rect 113550 6100 113610 6160
rect 113770 6260 113830 6320
rect 113770 6180 113830 6240
rect 113770 6100 113830 6160
rect 113990 6310 114050 6320
rect 113990 6270 114000 6310
rect 114000 6270 114040 6310
rect 114040 6270 114050 6310
rect 113990 6260 114050 6270
rect 113990 6180 114050 6240
rect 113990 6100 114050 6160
rect 113280 5880 113340 5940
rect 113580 5880 113640 5940
rect 112238 5820 112292 5830
rect 112238 5780 112245 5820
rect 112245 5780 112285 5820
rect 112285 5780 112292 5820
rect 112238 5770 112292 5780
rect 112348 5820 112402 5830
rect 112348 5780 112355 5820
rect 112355 5780 112395 5820
rect 112395 5780 112402 5820
rect 112348 5770 112402 5780
rect 112458 5820 112512 5830
rect 112458 5780 112465 5820
rect 112465 5780 112505 5820
rect 112505 5780 112512 5820
rect 112458 5770 112512 5780
rect 112568 5820 112622 5830
rect 112568 5780 112575 5820
rect 112575 5780 112615 5820
rect 112615 5780 112622 5820
rect 112568 5770 112622 5780
rect 112678 5820 112732 5830
rect 112678 5780 112685 5820
rect 112685 5780 112725 5820
rect 112725 5780 112732 5820
rect 112678 5770 112732 5780
rect 112788 5820 112842 5830
rect 112788 5780 112795 5820
rect 112795 5780 112835 5820
rect 112835 5780 112842 5820
rect 112788 5770 112842 5780
rect 112898 5820 112952 5830
rect 112898 5780 112905 5820
rect 112905 5780 112945 5820
rect 112945 5780 112952 5820
rect 112898 5770 112952 5780
rect 113008 5820 113062 5830
rect 113008 5780 113015 5820
rect 113015 5780 113055 5820
rect 113055 5780 113062 5820
rect 113008 5770 113062 5780
rect 113118 5820 113172 5830
rect 113118 5780 113125 5820
rect 113125 5780 113165 5820
rect 113165 5780 113172 5820
rect 113118 5770 113172 5780
rect 113228 5820 113282 5830
rect 113228 5780 113235 5820
rect 113235 5780 113275 5820
rect 113275 5780 113282 5820
rect 113228 5770 113282 5780
rect 112290 5360 112350 5420
rect 112180 5250 112240 5310
rect 112070 5140 112130 5200
rect 112070 5060 112130 5120
rect 112070 4980 112130 5040
rect 112510 5360 112570 5420
rect 112400 5250 112460 5310
rect 112080 4000 112140 4010
rect 112080 3960 112090 4000
rect 112090 3960 112130 4000
rect 112130 3960 112140 4000
rect 112180 3970 112240 4030
rect 112290 3990 112350 4050
rect 112730 5360 112790 5420
rect 112620 5250 112680 5310
rect 112400 3970 112460 4030
rect 112510 3990 112570 4050
rect 112950 5360 113010 5420
rect 112840 5250 112900 5310
rect 112620 3970 112680 4030
rect 112730 3990 112790 4050
rect 113170 5360 113230 5420
rect 113060 5250 113120 5310
rect 112840 3970 112900 4030
rect 112950 3990 113010 4050
rect 113280 5250 113340 5310
rect 113580 5250 113640 5310
rect 113960 5880 114020 5940
rect 114260 5880 114320 5940
rect 114480 5880 114540 5940
rect 114700 5880 114760 5940
rect 114920 5880 114980 5940
rect 115140 5880 115200 5940
rect 115360 5880 115420 5940
rect 114318 5820 114372 5830
rect 114318 5780 114325 5820
rect 114325 5780 114365 5820
rect 114365 5780 114372 5820
rect 114318 5770 114372 5780
rect 114428 5820 114482 5830
rect 114428 5780 114435 5820
rect 114435 5780 114475 5820
rect 114475 5780 114482 5820
rect 114428 5770 114482 5780
rect 114538 5820 114592 5830
rect 114538 5780 114545 5820
rect 114545 5780 114585 5820
rect 114585 5780 114592 5820
rect 114538 5770 114592 5780
rect 114648 5820 114702 5830
rect 114648 5780 114655 5820
rect 114655 5780 114695 5820
rect 114695 5780 114702 5820
rect 114648 5770 114702 5780
rect 114758 5820 114812 5830
rect 114758 5780 114765 5820
rect 114765 5780 114805 5820
rect 114805 5780 114812 5820
rect 114758 5770 114812 5780
rect 114868 5820 114922 5830
rect 114868 5780 114875 5820
rect 114875 5780 114915 5820
rect 114915 5780 114922 5820
rect 114868 5770 114922 5780
rect 114978 5820 115032 5830
rect 114978 5780 114985 5820
rect 114985 5780 115025 5820
rect 115025 5780 115032 5820
rect 114978 5770 115032 5780
rect 115088 5820 115142 5830
rect 115088 5780 115095 5820
rect 115095 5780 115135 5820
rect 115135 5780 115142 5820
rect 115088 5770 115142 5780
rect 115198 5820 115252 5830
rect 115198 5780 115205 5820
rect 115205 5780 115245 5820
rect 115245 5780 115252 5820
rect 115198 5770 115252 5780
rect 115308 5820 115362 5830
rect 115308 5780 115315 5820
rect 115315 5780 115355 5820
rect 115355 5780 115362 5820
rect 115308 5770 115362 5780
rect 113960 5250 114020 5310
rect 114370 5360 114430 5420
rect 114260 5250 114320 5310
rect 113390 5140 113450 5200
rect 113390 5060 113450 5120
rect 113390 4980 113450 5040
rect 114150 5140 114210 5200
rect 114150 5060 114210 5120
rect 114150 4980 114210 5040
rect 113770 4330 113830 4390
rect 113770 4250 113830 4310
rect 113770 4170 113830 4230
rect 113060 3970 113120 4030
rect 113170 3990 113230 4050
rect 113280 3970 113340 4030
rect 113380 4020 113440 4030
rect 113380 3980 113390 4020
rect 113390 3980 113430 4020
rect 113430 3980 113440 4020
rect 113380 3970 113440 3980
rect 113680 4020 113740 4030
rect 113680 3980 113690 4020
rect 113690 3980 113730 4020
rect 113730 3980 113740 4020
rect 113680 3970 113740 3980
rect 112080 3950 112140 3960
rect 112290 3880 112350 3940
rect 112180 3490 112240 3550
rect 112510 3880 112570 3940
rect 112400 3490 112460 3550
rect 112730 3880 112790 3940
rect 112620 3490 112680 3550
rect 112950 3880 113010 3940
rect 112840 3490 112900 3550
rect 113170 3880 113230 3940
rect 113060 3490 113120 3550
rect 113280 3490 113340 3550
rect 114590 5360 114650 5420
rect 114480 5250 114540 5310
rect 113860 4020 113920 4030
rect 113860 3980 113870 4020
rect 113870 3980 113910 4020
rect 113910 3980 113920 4020
rect 113860 3970 113920 3980
rect 114160 4020 114220 4030
rect 114160 3980 114170 4020
rect 114170 3980 114210 4020
rect 114210 3980 114220 4020
rect 114160 3970 114220 3980
rect 114260 3970 114320 4030
rect 114370 3990 114430 4050
rect 114810 5360 114870 5420
rect 114700 5250 114760 5310
rect 114480 3970 114540 4030
rect 114590 3990 114650 4050
rect 115030 5360 115090 5420
rect 114920 5250 114980 5310
rect 114700 3970 114760 4030
rect 114810 3990 114870 4050
rect 115250 5360 115310 5420
rect 115140 5250 115200 5310
rect 114920 3970 114980 4030
rect 115030 3990 115090 4050
rect 115360 5250 115420 5310
rect 115470 5140 115530 5200
rect 115470 5060 115530 5120
rect 115470 4980 115530 5040
rect 115140 3970 115200 4030
rect 115250 3990 115310 4050
rect 115360 3970 115420 4030
rect 115460 4000 115520 4010
rect 115460 3960 115470 4000
rect 115470 3960 115510 4000
rect 115510 3960 115520 4000
rect 114370 3880 114430 3940
rect 113660 3490 113720 3550
rect 112290 3350 112350 3410
rect 112510 3350 112570 3410
rect 112730 3350 112790 3410
rect 112950 3350 113010 3410
rect 113170 3350 113230 3410
rect 112070 2440 112130 2500
rect 112070 2360 112130 2420
rect 112070 2280 112130 2340
rect 111890 2170 111950 2230
rect 113470 2440 113530 2500
rect 113470 2360 113530 2420
rect 113470 2280 113530 2340
rect 112890 1670 112950 1730
rect 113110 1670 113170 1730
rect 113330 1670 113390 1730
rect 113550 1670 113610 1730
rect 113880 3490 113940 3550
rect 113770 1670 113830 1730
rect 114260 3490 114320 3550
rect 114590 3880 114650 3940
rect 114480 3490 114540 3550
rect 114810 3880 114870 3940
rect 114700 3490 114760 3550
rect 115030 3880 115090 3940
rect 114920 3490 114980 3550
rect 115250 3880 115310 3940
rect 115140 3490 115200 3550
rect 115460 3950 115520 3960
rect 115360 3490 115420 3550
rect 114370 3350 114430 3410
rect 114590 3350 114650 3410
rect 114070 2440 114130 2500
rect 114070 2360 114130 2420
rect 114070 2280 114130 2340
rect 113990 1670 114050 1730
rect 114810 3350 114870 3410
rect 115030 3350 115090 3410
rect 115250 3350 115310 3410
rect 115470 2440 115530 2500
rect 115470 2360 115530 2420
rect 115470 2280 115530 2340
rect 116300 7210 116360 7270
rect 116380 7210 116440 7270
rect 116460 7210 116520 7270
rect 116300 7130 116360 7190
rect 116380 7130 116440 7190
rect 116460 7130 116520 7190
rect 115730 7010 115790 7070
rect 115640 2170 115700 2230
rect 114210 1670 114270 1730
rect 114430 1670 114490 1730
rect 114650 1670 114710 1730
rect 114870 1670 114930 1730
rect 111700 140 111760 200
rect 112450 1060 112510 1070
rect 112450 1020 112460 1060
rect 112460 1020 112500 1060
rect 112500 1020 112510 1060
rect 112450 1010 112510 1020
rect 110310 -90 110370 -30
rect 112560 1010 112620 1070
rect 112780 1010 112840 1070
rect 113000 1010 113060 1070
rect 113220 1010 113280 1070
rect 113440 1010 113500 1070
rect 113660 1010 113720 1070
rect 113880 1010 113940 1070
rect 114100 1010 114160 1070
rect 114320 1010 114380 1070
rect 114540 1010 114600 1070
rect 114760 1010 114820 1070
rect 114980 1060 115040 1070
rect 114980 1020 114990 1060
rect 114990 1020 115030 1060
rect 115030 1020 115040 1060
rect 114980 1010 115040 1020
rect 112890 900 112950 960
rect 112890 820 112950 880
rect 112890 740 112950 800
rect 113110 900 113170 960
rect 113110 820 113170 880
rect 113110 740 113170 800
rect 113330 900 113390 960
rect 113330 820 113390 880
rect 113330 740 113390 800
rect 113550 900 113610 960
rect 113550 820 113610 880
rect 113550 740 113610 800
rect 113770 900 113830 960
rect 113770 820 113830 880
rect 113770 740 113830 800
rect 113990 900 114050 960
rect 113990 820 114050 880
rect 113990 740 114050 800
rect 114210 900 114270 960
rect 114210 820 114270 880
rect 114210 740 114270 800
rect 114430 900 114490 960
rect 114430 820 114490 880
rect 114430 740 114490 800
rect 114650 900 114710 960
rect 114650 820 114710 880
rect 114650 740 114710 800
rect 114870 900 114930 960
rect 114870 820 114930 880
rect 114870 740 114930 800
rect 114840 680 114900 690
rect 114840 640 114850 680
rect 114850 640 114890 680
rect 114890 640 114900 680
rect 114840 630 114900 640
rect 112670 520 112730 580
rect 112670 440 112730 500
rect 112670 360 112730 420
rect 112450 -300 112510 -240
rect 113250 250 113310 310
rect 113660 250 113720 310
rect 113880 250 113940 310
rect 113550 140 113610 200
rect 113770 190 113830 200
rect 113770 150 113780 190
rect 113780 150 113820 190
rect 113820 150 113830 190
rect 113770 140 113830 150
rect 113990 140 114050 200
rect 113550 -300 113610 -240
rect 113770 -300 113830 -240
rect 113990 -300 114050 -240
rect 114100 -250 114160 -240
rect 114100 -290 114110 -250
rect 114110 -290 114150 -250
rect 114150 -290 114160 -250
rect 114100 -300 114160 -290
rect 114980 -300 115040 -240
rect 113770 -330 113830 -320
rect 113770 -370 113780 -330
rect 113780 -370 113820 -330
rect 113820 -370 113830 -330
rect 113770 -380 113830 -370
rect 113250 -520 113310 -460
rect 113250 -600 113310 -540
rect 113250 -680 113310 -620
rect 113430 -690 113440 -450
rect 113440 -690 113480 -450
rect 113480 -690 113490 -450
rect 114110 -690 114120 -450
rect 114120 -690 114160 -450
rect 114160 -690 114170 -450
rect 110190 -1220 110250 -1160
rect 110270 -1220 110330 -1160
rect 110350 -1220 110410 -1160
rect 110190 -1300 110250 -1240
rect 110270 -1300 110330 -1240
rect 110350 -1300 110410 -1240
rect 110190 -1380 110250 -1320
rect 110270 -1380 110330 -1320
rect 110350 -1380 110410 -1320
rect 110510 -1220 110570 -1160
rect 110510 -1300 110570 -1240
rect 110510 -1380 110570 -1320
rect 110890 -1220 110950 -1160
rect 110970 -1220 111030 -1160
rect 111050 -1220 111110 -1160
rect 110890 -1300 110950 -1240
rect 110970 -1300 111030 -1240
rect 111050 -1300 111110 -1240
rect 110890 -1380 110950 -1320
rect 110970 -1380 111030 -1320
rect 111050 -1380 111110 -1320
rect 111590 -1220 111650 -1160
rect 111670 -1220 111730 -1160
rect 111750 -1220 111810 -1160
rect 111590 -1300 111650 -1240
rect 111670 -1300 111730 -1240
rect 111750 -1300 111810 -1240
rect 111590 -1380 111650 -1320
rect 111670 -1380 111730 -1320
rect 111750 -1380 111810 -1320
rect 112290 -1220 112350 -1160
rect 112370 -1220 112430 -1160
rect 112450 -1220 112510 -1160
rect 112290 -1300 112350 -1240
rect 112370 -1300 112430 -1240
rect 112450 -1300 112510 -1240
rect 112290 -1380 112350 -1320
rect 112370 -1380 112430 -1320
rect 112450 -1380 112510 -1320
rect 112990 -1220 113050 -1160
rect 113070 -1220 113130 -1160
rect 113150 -1220 113210 -1160
rect 112990 -1300 113050 -1240
rect 113070 -1300 113130 -1240
rect 113150 -1300 113210 -1240
rect 112990 -1380 113050 -1320
rect 113070 -1380 113130 -1320
rect 113150 -1380 113210 -1320
rect 113690 -1220 113750 -1160
rect 113770 -1220 113830 -1160
rect 113850 -1220 113910 -1160
rect 113690 -1300 113750 -1240
rect 113770 -1300 113830 -1240
rect 113850 -1300 113910 -1240
rect 113690 -1380 113750 -1320
rect 113770 -1380 113830 -1320
rect 113850 -1380 113910 -1320
rect 114390 -1220 114450 -1160
rect 114470 -1220 114530 -1160
rect 114550 -1220 114610 -1160
rect 114390 -1300 114450 -1240
rect 114470 -1300 114530 -1240
rect 114550 -1300 114610 -1240
rect 114390 -1380 114450 -1320
rect 114470 -1380 114530 -1320
rect 114550 -1380 114610 -1320
rect 115090 900 115150 960
rect 115170 900 115230 960
rect 115250 900 115310 960
rect 115090 820 115150 880
rect 115170 820 115230 880
rect 115250 820 115310 880
rect 115090 740 115150 800
rect 115170 740 115230 800
rect 115250 740 115310 800
rect 116030 6260 116090 6320
rect 116110 6260 116170 6320
rect 116190 6260 116250 6320
rect 116030 6180 116090 6240
rect 116110 6180 116170 6240
rect 116190 6180 116250 6240
rect 116030 6100 116090 6160
rect 116110 6100 116170 6160
rect 116190 6100 116250 6160
rect 116030 5960 116090 6020
rect 116110 5960 116170 6020
rect 116190 5960 116250 6020
rect 116030 5880 116090 5940
rect 116110 5880 116170 5940
rect 116190 5880 116250 5940
rect 115840 5770 115900 5830
rect 115730 630 115790 690
rect 116030 5800 116090 5860
rect 116110 5800 116170 5860
rect 116190 5800 116250 5860
rect 116030 5140 116090 5200
rect 116110 5140 116170 5200
rect 116190 5140 116250 5200
rect 116030 5060 116090 5120
rect 116110 5060 116170 5120
rect 116190 5060 116250 5120
rect 116030 4980 116090 5040
rect 116110 4980 116170 5040
rect 116190 4980 116250 5040
rect 116030 4660 116090 4720
rect 116110 4660 116170 4720
rect 116190 4660 116250 4720
rect 116030 4580 116090 4640
rect 116110 4580 116170 4640
rect 116190 4580 116250 4640
rect 116030 4500 116090 4560
rect 116110 4500 116170 4560
rect 116190 4500 116250 4560
rect 116300 4930 116360 4990
rect 116380 4930 116440 4990
rect 116460 4930 116520 4990
rect 116300 4850 116360 4910
rect 116380 4850 116440 4910
rect 116460 4850 116520 4910
rect 116300 4770 116360 4830
rect 116380 4770 116440 4830
rect 116460 4770 116520 4830
rect 116030 4330 116090 4390
rect 116110 4330 116170 4390
rect 116190 4330 116250 4390
rect 116030 4250 116090 4310
rect 116110 4250 116170 4310
rect 116190 4250 116250 4310
rect 116030 4170 116090 4230
rect 116110 4170 116170 4230
rect 116190 4170 116250 4230
rect 116570 7510 116630 7570
rect 116650 7510 116710 7570
rect 116730 7510 116790 7570
rect 117030 7510 117090 7570
rect 117270 7510 117330 7570
rect 117510 7510 117570 7570
rect 117750 7510 117810 7570
rect 117990 7510 118050 7570
rect 118230 7510 118290 7570
rect 117090 7450 117150 7460
rect 117090 7410 117100 7450
rect 117100 7410 117140 7450
rect 117140 7410 117150 7450
rect 117090 7400 117150 7410
rect 117210 7450 117270 7460
rect 117210 7410 117220 7450
rect 117220 7410 117260 7450
rect 117260 7410 117270 7450
rect 117210 7400 117270 7410
rect 117330 7450 117390 7460
rect 117330 7410 117340 7450
rect 117340 7410 117380 7450
rect 117380 7410 117390 7450
rect 117330 7400 117390 7410
rect 117450 7450 117510 7460
rect 117450 7410 117460 7450
rect 117460 7410 117500 7450
rect 117500 7410 117510 7450
rect 117450 7400 117510 7410
rect 117570 7450 117630 7460
rect 117570 7410 117580 7450
rect 117580 7410 117620 7450
rect 117620 7410 117630 7450
rect 117570 7400 117630 7410
rect 117690 7450 117750 7460
rect 117690 7410 117700 7450
rect 117700 7410 117740 7450
rect 117740 7410 117750 7450
rect 117690 7400 117750 7410
rect 117810 7450 117870 7460
rect 117810 7410 117820 7450
rect 117820 7410 117860 7450
rect 117860 7410 117870 7450
rect 117810 7400 117870 7410
rect 117930 7450 117990 7460
rect 117930 7410 117940 7450
rect 117940 7410 117980 7450
rect 117980 7410 117990 7450
rect 117930 7400 117990 7410
rect 118050 7450 118110 7460
rect 118050 7410 118060 7450
rect 118060 7410 118100 7450
rect 118100 7410 118110 7450
rect 118050 7400 118110 7410
rect 118170 7450 118230 7460
rect 118170 7410 118180 7450
rect 118180 7410 118220 7450
rect 118220 7410 118230 7450
rect 118170 7400 118230 7410
rect 116970 7290 117030 7350
rect 116970 7210 117030 7270
rect 116970 7130 117030 7190
rect 117190 7290 117250 7350
rect 117190 7210 117250 7270
rect 117190 7130 117250 7190
rect 117410 7290 117470 7350
rect 117410 7210 117470 7270
rect 117410 7130 117470 7190
rect 117630 7290 117690 7350
rect 117630 7210 117690 7270
rect 117630 7130 117690 7190
rect 117850 7290 117910 7350
rect 117850 7210 117910 7270
rect 117850 7130 117910 7190
rect 118070 7290 118130 7350
rect 118070 7210 118130 7270
rect 118070 7130 118130 7190
rect 118290 7290 118350 7350
rect 118290 7210 118350 7270
rect 118290 7130 118350 7190
rect 116570 6900 116630 6960
rect 116650 6900 116710 6960
rect 116730 6900 116790 6960
rect 116570 6820 116630 6880
rect 116650 6820 116710 6880
rect 116730 6820 116790 6880
rect 116570 6740 116630 6800
rect 116650 6740 116710 6800
rect 116730 6740 116790 6800
rect 117080 6940 117140 7000
rect 117300 6940 117360 7000
rect 117520 6940 117580 7000
rect 117740 6940 117800 7000
rect 117960 6940 118020 7000
rect 120690 9280 120750 9340
rect 120770 9280 120830 9340
rect 120850 9280 120910 9340
rect 120690 9200 120750 9260
rect 120770 9200 120830 9260
rect 120850 9200 120910 9260
rect 120690 9120 120750 9180
rect 120770 9120 120830 9180
rect 120850 9120 120910 9180
rect 121390 9280 121450 9340
rect 121470 9280 121530 9340
rect 121550 9280 121610 9340
rect 121390 9200 121450 9260
rect 121470 9200 121530 9260
rect 121550 9200 121610 9260
rect 121390 9120 121450 9180
rect 121470 9120 121530 9180
rect 121550 9120 121610 9180
rect 122090 9280 122150 9340
rect 122170 9280 122230 9340
rect 122250 9280 122310 9340
rect 122090 9200 122150 9260
rect 122170 9200 122230 9260
rect 122250 9200 122310 9260
rect 122090 9120 122150 9180
rect 122170 9120 122230 9180
rect 122250 9120 122310 9180
rect 122790 9280 122850 9340
rect 122870 9280 122930 9340
rect 122950 9280 123010 9340
rect 122790 9200 122850 9260
rect 122870 9200 122930 9260
rect 122950 9200 123010 9260
rect 122790 9120 122850 9180
rect 122870 9120 122930 9180
rect 122950 9120 123010 9180
rect 119290 7290 119350 7350
rect 119370 7290 119430 7350
rect 119450 7290 119510 7350
rect 119290 7210 119350 7270
rect 119370 7210 119430 7270
rect 119450 7210 119510 7270
rect 119290 7130 119350 7190
rect 119370 7130 119430 7190
rect 119450 7130 119510 7190
rect 118180 6940 118240 7000
rect 116570 5500 116630 5560
rect 116650 5500 116710 5560
rect 116730 5500 116790 5560
rect 116570 5420 116630 5480
rect 116650 5420 116710 5480
rect 116730 5420 116790 5480
rect 116570 5340 116630 5400
rect 116650 5340 116710 5400
rect 116730 5340 116790 5400
rect 117080 5660 117140 5720
rect 117300 5660 117360 5720
rect 117520 5660 117580 5720
rect 117740 5660 117800 5720
rect 117630 5550 117690 5560
rect 117630 5510 117640 5550
rect 117640 5510 117680 5550
rect 117680 5510 117690 5550
rect 117630 5500 117690 5510
rect 117630 5470 117690 5480
rect 117630 5430 117640 5470
rect 117640 5430 117680 5470
rect 117680 5430 117690 5470
rect 117630 5420 117690 5430
rect 117630 5390 117690 5400
rect 117630 5350 117640 5390
rect 117640 5350 117680 5390
rect 117680 5350 117690 5390
rect 117630 5340 117690 5350
rect 117960 5660 118020 5720
rect 118180 5660 118240 5720
rect 118940 5500 119000 5560
rect 119020 5500 119080 5560
rect 119100 5500 119160 5560
rect 118940 5420 119000 5480
rect 119020 5420 119080 5480
rect 119100 5420 119160 5480
rect 118940 5340 119000 5400
rect 119020 5340 119080 5400
rect 119100 5340 119160 5400
rect 117080 5200 117140 5260
rect 117190 5200 117250 5260
rect 117300 5200 117360 5260
rect 117410 5200 117470 5260
rect 117520 5200 117580 5260
rect 117630 5200 117690 5260
rect 117740 5200 117800 5260
rect 117850 5200 117910 5260
rect 117960 5200 118020 5260
rect 118070 5200 118130 5260
rect 118180 5200 118240 5260
rect 117080 5120 117140 5180
rect 117190 5120 117250 5180
rect 117300 5120 117360 5180
rect 117410 5120 117470 5180
rect 117520 5120 117580 5180
rect 117630 5120 117690 5180
rect 117740 5120 117800 5180
rect 117850 5120 117910 5180
rect 117960 5120 118020 5180
rect 118070 5120 118130 5180
rect 118180 5120 118240 5180
rect 117080 5040 117140 5100
rect 117190 5040 117250 5100
rect 117300 5040 117360 5100
rect 117410 5040 117470 5100
rect 117520 5040 117580 5100
rect 117630 5040 117690 5100
rect 117740 5040 117800 5100
rect 117850 5040 117910 5100
rect 117960 5040 118020 5100
rect 118070 5040 118130 5100
rect 118180 5040 118240 5100
rect 119130 5200 119190 5260
rect 119210 5200 119270 5260
rect 119300 5200 119360 5260
rect 119380 5200 119440 5260
rect 119470 5200 119530 5260
rect 119550 5200 119610 5260
rect 119130 5120 119190 5180
rect 119210 5120 119270 5180
rect 119300 5120 119360 5180
rect 119380 5120 119440 5180
rect 119470 5120 119530 5180
rect 119550 5120 119610 5180
rect 119130 5040 119190 5100
rect 119210 5040 119270 5100
rect 119300 5040 119360 5100
rect 119380 5040 119440 5100
rect 119470 5040 119530 5100
rect 119550 5040 119610 5100
rect 116970 4930 117030 4990
rect 116970 4850 117030 4910
rect 116970 4770 117030 4830
rect 118290 4930 118350 4990
rect 118290 4850 118350 4910
rect 118290 4770 118350 4830
rect 117080 4660 117140 4720
rect 117080 4580 117140 4640
rect 117080 4500 117140 4560
rect 117300 4660 117360 4720
rect 117300 4580 117360 4640
rect 117300 4500 117360 4560
rect 117520 4660 117580 4720
rect 117520 4580 117580 4640
rect 117520 4500 117580 4560
rect 117740 4660 117800 4720
rect 117740 4580 117800 4640
rect 117740 4500 117800 4560
rect 117960 4660 118020 4720
rect 117960 4580 118020 4640
rect 117960 4500 118020 4560
rect 118180 4660 118240 4720
rect 118180 4580 118240 4640
rect 118180 4500 118240 4560
rect 117190 4390 117250 4450
rect 117410 4390 117470 4450
rect 117630 4390 117690 4450
rect 117850 4390 117910 4450
rect 118070 4390 118130 4450
rect 119140 4060 119200 4120
rect 119240 4060 119300 4120
rect 119340 4060 119400 4120
rect 119440 4060 119500 4120
rect 119540 4060 119600 4120
rect 119140 3960 119200 4020
rect 119240 3960 119300 4020
rect 119340 3960 119400 4020
rect 119440 3960 119500 4020
rect 119540 3960 119600 4020
rect 117190 3930 117250 3940
rect 117190 3890 117200 3930
rect 117200 3890 117240 3930
rect 117240 3890 117250 3930
rect 117190 3880 117250 3890
rect 117410 3930 117470 3940
rect 117410 3890 117420 3930
rect 117420 3890 117460 3930
rect 117460 3890 117470 3930
rect 117410 3880 117470 3890
rect 117630 3930 117690 3940
rect 117630 3890 117640 3930
rect 117640 3890 117680 3930
rect 117680 3890 117690 3930
rect 117630 3880 117690 3890
rect 117850 3930 117910 3940
rect 117850 3890 117860 3930
rect 117860 3890 117900 3930
rect 117900 3890 117910 3930
rect 117850 3880 117910 3890
rect 118070 3930 118130 3940
rect 118070 3890 118080 3930
rect 118080 3890 118120 3930
rect 118120 3890 118130 3930
rect 118070 3880 118130 3890
rect 118560 3880 118620 3940
rect 116570 3750 116630 3810
rect 116650 3750 116710 3810
rect 116730 3750 116790 3810
rect 116570 3670 116630 3730
rect 116650 3670 116710 3730
rect 116730 3670 116790 3730
rect 117300 3800 117360 3810
rect 117300 3760 117310 3800
rect 117310 3760 117350 3800
rect 117350 3760 117360 3800
rect 117300 3750 117360 3760
rect 117300 3720 117360 3730
rect 117300 3680 117310 3720
rect 117310 3680 117350 3720
rect 117350 3680 117360 3720
rect 117300 3670 117360 3680
rect 117190 3510 117250 3570
rect 117410 3510 117470 3570
rect 117630 3510 117690 3570
rect 117850 3510 117910 3570
rect 118070 3510 118130 3570
rect 118470 3510 118530 3570
rect 116570 2990 116630 3050
rect 116650 2990 116710 3050
rect 116730 2990 116790 3050
rect 116570 2910 116630 2970
rect 116650 2910 116710 2970
rect 116730 2910 116790 2970
rect 116570 2830 116630 2890
rect 116650 2830 116710 2890
rect 116730 2830 116790 2890
rect 116300 2720 116360 2780
rect 116380 2720 116440 2780
rect 116460 2720 116520 2780
rect 116300 2640 116360 2700
rect 116380 2640 116440 2700
rect 116460 2640 116520 2700
rect 116300 2560 116360 2620
rect 116380 2560 116440 2620
rect 116460 2560 116520 2620
rect 117190 2830 117250 2890
rect 117410 2830 117470 2890
rect 117630 2830 117690 2890
rect 117850 2830 117910 2890
rect 118070 2830 118130 2890
rect 118470 2870 118530 2930
rect 117080 2720 117140 2780
rect 117080 2640 117140 2700
rect 117080 2560 117140 2620
rect 117300 2720 117360 2780
rect 117300 2640 117360 2700
rect 117300 2560 117360 2620
rect 117520 2720 117580 2780
rect 117520 2640 117580 2700
rect 117520 2560 117580 2620
rect 117740 2720 117800 2780
rect 117740 2640 117800 2700
rect 117740 2560 117800 2620
rect 117960 2720 118020 2780
rect 117960 2640 118020 2700
rect 117960 2560 118020 2620
rect 118180 2720 118240 2780
rect 118180 2640 118240 2700
rect 118180 2560 118240 2620
rect 119140 3860 119200 3920
rect 119240 3860 119300 3920
rect 119340 3860 119400 3920
rect 119440 3860 119500 3920
rect 119540 3860 119600 3920
rect 118660 2930 118730 2940
rect 118660 2880 118670 2930
rect 118670 2880 118720 2930
rect 118720 2880 118730 2930
rect 118660 2870 118730 2880
rect 118780 2930 118850 2940
rect 118780 2880 118790 2930
rect 118790 2880 118840 2930
rect 118840 2880 118850 2930
rect 118780 2870 118850 2880
rect 118900 2930 118970 2940
rect 118900 2880 118910 2930
rect 118910 2880 118960 2930
rect 118960 2880 118970 2930
rect 118900 2870 118970 2880
rect 119020 2930 119090 2940
rect 119020 2880 119030 2930
rect 119030 2880 119080 2930
rect 119080 2880 119090 2930
rect 119020 2870 119090 2880
rect 118560 2730 118620 2790
rect 118780 2730 118840 2790
rect 116970 2440 117030 2500
rect 116970 2360 117030 2420
rect 116970 2280 117030 2340
rect 118290 2440 118350 2500
rect 118290 2360 118350 2420
rect 118290 2280 118350 2340
rect 119020 2170 119080 2230
rect 118890 1790 118950 1850
rect 117230 1680 117290 1740
rect 117310 1680 117370 1740
rect 117390 1680 117450 1740
rect 117470 1680 117530 1740
rect 117550 1680 117610 1740
rect 117630 1680 117690 1740
rect 117710 1680 117770 1740
rect 117790 1680 117850 1740
rect 117870 1680 117930 1740
rect 117950 1680 118010 1740
rect 118030 1680 118090 1740
rect 117230 1600 117290 1660
rect 117310 1600 117370 1660
rect 117390 1600 117450 1660
rect 117470 1600 117530 1660
rect 117550 1600 117610 1660
rect 117630 1600 117690 1660
rect 117710 1600 117770 1660
rect 117790 1600 117850 1660
rect 117870 1600 117930 1660
rect 117950 1600 118010 1660
rect 118030 1600 118090 1660
rect 117230 1520 117290 1580
rect 117310 1520 117370 1580
rect 117390 1520 117450 1580
rect 117470 1520 117530 1580
rect 117550 1520 117610 1580
rect 117630 1520 117690 1580
rect 117710 1520 117770 1580
rect 117790 1520 117850 1580
rect 117870 1520 117930 1580
rect 117950 1520 118010 1580
rect 118030 1520 118090 1580
rect 118760 1680 118820 1740
rect 118760 1600 118820 1660
rect 118760 1520 118820 1580
rect 116030 520 116090 580
rect 116110 520 116170 580
rect 116190 520 116250 580
rect 116030 440 116090 500
rect 116110 440 116170 500
rect 116190 440 116250 500
rect 116030 360 116090 420
rect 116110 360 116170 420
rect 116190 360 116250 420
rect 115840 140 115900 200
rect 115090 -520 115150 -460
rect 115170 -520 115230 -460
rect 115250 -520 115310 -460
rect 115090 -600 115150 -540
rect 115170 -600 115230 -540
rect 115250 -600 115310 -540
rect 115090 -680 115150 -620
rect 115170 -680 115230 -620
rect 115250 -680 115310 -620
rect 117330 1460 117390 1470
rect 117330 1420 117340 1460
rect 117340 1420 117380 1460
rect 117380 1420 117390 1460
rect 117330 1410 117390 1420
rect 117530 1460 117590 1470
rect 117530 1420 117540 1460
rect 117540 1420 117580 1460
rect 117580 1420 117590 1460
rect 117530 1410 117590 1420
rect 117230 -90 117290 -30
rect 117730 1460 117790 1470
rect 117730 1420 117740 1460
rect 117740 1420 117780 1460
rect 117780 1420 117790 1460
rect 117730 1410 117790 1420
rect 117930 1460 117990 1470
rect 117930 1420 117940 1460
rect 117940 1420 117980 1460
rect 117980 1420 117990 1460
rect 117930 1410 117990 1420
rect 117630 -90 117690 -30
rect 114980 -1220 115040 -1160
rect 114980 -1300 115040 -1240
rect 114980 -1380 115040 -1320
rect 115090 -1220 115150 -1160
rect 115170 -1220 115230 -1160
rect 115250 -1220 115310 -1160
rect 115090 -1300 115150 -1240
rect 115170 -1300 115230 -1240
rect 115250 -1300 115310 -1240
rect 115090 -1380 115150 -1320
rect 115170 -1380 115230 -1320
rect 115250 -1380 115310 -1320
rect 115790 -1220 115850 -1160
rect 115870 -1220 115930 -1160
rect 115950 -1220 116010 -1160
rect 115790 -1300 115850 -1240
rect 115870 -1300 115930 -1240
rect 115950 -1300 116010 -1240
rect 115790 -1380 115850 -1320
rect 115870 -1380 115930 -1320
rect 115950 -1380 116010 -1320
rect 116490 -1220 116550 -1160
rect 116570 -1220 116630 -1160
rect 116650 -1220 116710 -1160
rect 116490 -1300 116550 -1240
rect 116570 -1300 116630 -1240
rect 116650 -1300 116710 -1240
rect 116490 -1380 116550 -1320
rect 116570 -1380 116630 -1320
rect 116650 -1380 116710 -1320
rect 117030 -1220 117090 -1160
rect 117030 -1300 117090 -1240
rect 117030 -1380 117090 -1320
rect 117190 -1220 117250 -1160
rect 117270 -1220 117330 -1160
rect 117350 -1220 117410 -1160
rect 117190 -1300 117250 -1240
rect 117270 -1300 117330 -1240
rect 117350 -1300 117410 -1240
rect 117190 -1380 117250 -1320
rect 117270 -1380 117330 -1320
rect 117350 -1380 117410 -1320
rect 118760 1350 118830 1360
rect 118760 1300 118770 1350
rect 118770 1300 118820 1350
rect 118820 1300 118830 1350
rect 118760 1290 118830 1300
rect 119130 1680 119190 1740
rect 119210 1680 119270 1740
rect 119300 1680 119360 1740
rect 119380 1680 119440 1740
rect 119470 1680 119530 1740
rect 119550 1680 119610 1740
rect 119130 1600 119190 1660
rect 119210 1600 119270 1660
rect 119300 1600 119360 1660
rect 119380 1600 119440 1660
rect 119470 1600 119530 1660
rect 119550 1600 119610 1660
rect 119130 1520 119190 1580
rect 119210 1520 119270 1580
rect 119300 1520 119360 1580
rect 119380 1520 119440 1580
rect 119470 1520 119530 1580
rect 119550 1520 119610 1580
rect 119690 4650 119750 4710
rect 119770 4650 119830 4710
rect 119850 4650 119910 4710
rect 119690 4570 119750 4630
rect 119770 4570 119830 4630
rect 119850 4570 119910 4630
rect 119690 4490 119750 4550
rect 119770 4490 119830 4550
rect 119850 4490 119910 4550
rect 119690 2440 119750 2500
rect 119770 2440 119830 2500
rect 119850 2440 119910 2500
rect 119690 2360 119750 2420
rect 119770 2360 119830 2420
rect 119850 2360 119910 2420
rect 119690 2280 119750 2340
rect 119770 2280 119830 2340
rect 119850 2280 119910 2340
rect 118890 1410 118950 1470
rect 118880 1350 118950 1360
rect 118880 1300 118890 1350
rect 118890 1300 118940 1350
rect 118940 1300 118950 1350
rect 118880 1290 118950 1300
rect 118030 -90 118090 -30
rect 117890 -1220 117950 -1160
rect 117970 -1220 118030 -1160
rect 118050 -1220 118110 -1160
rect 117890 -1300 117950 -1240
rect 117970 -1300 118030 -1240
rect 118050 -1300 118110 -1240
rect 117890 -1380 117950 -1320
rect 117970 -1380 118030 -1320
rect 118050 -1380 118110 -1320
rect 118230 -1220 118290 -1160
rect 118230 -1300 118290 -1240
rect 118230 -1380 118290 -1320
rect 118750 -1220 118810 -1160
rect 118830 -1220 118890 -1160
rect 118910 -1220 118970 -1160
rect 118750 -1300 118810 -1240
rect 118830 -1300 118890 -1240
rect 118910 -1300 118970 -1240
rect 118750 -1380 118810 -1320
rect 118830 -1380 118890 -1320
rect 118910 -1380 118970 -1320
rect 119290 -1220 119350 -1160
rect 119370 -1220 119430 -1160
rect 119450 -1220 119510 -1160
rect 119290 -1300 119350 -1240
rect 119370 -1300 119430 -1240
rect 119450 -1300 119510 -1240
rect 119290 -1380 119350 -1320
rect 119370 -1380 119430 -1320
rect 119450 -1380 119510 -1320
rect 119690 -1220 119750 -1160
rect 119770 -1220 119830 -1160
rect 119850 -1220 119910 -1160
rect 119690 -1300 119750 -1240
rect 119770 -1300 119830 -1240
rect 119850 -1300 119910 -1240
rect 119690 -1380 119750 -1320
rect 119770 -1380 119830 -1320
rect 119850 -1380 119910 -1320
rect 119990 -1220 120050 -1160
rect 120070 -1220 120130 -1160
rect 120150 -1220 120210 -1160
rect 119990 -1300 120050 -1240
rect 120070 -1300 120130 -1240
rect 120150 -1300 120210 -1240
rect 119990 -1380 120050 -1320
rect 120070 -1380 120130 -1320
rect 120150 -1380 120210 -1320
rect 120690 -1220 120750 -1160
rect 120770 -1220 120830 -1160
rect 120850 -1220 120910 -1160
rect 120690 -1300 120750 -1240
rect 120770 -1300 120830 -1240
rect 120850 -1300 120910 -1240
rect 120690 -1380 120750 -1320
rect 120770 -1380 120830 -1320
rect 120850 -1380 120910 -1320
rect 121390 -1220 121450 -1160
rect 121470 -1220 121530 -1160
rect 121550 -1220 121610 -1160
rect 121390 -1300 121450 -1240
rect 121470 -1300 121530 -1240
rect 121550 -1300 121610 -1240
rect 121390 -1380 121450 -1320
rect 121470 -1380 121530 -1320
rect 121550 -1380 121610 -1320
rect 122090 -1220 122150 -1160
rect 122170 -1220 122230 -1160
rect 122250 -1220 122310 -1160
rect 122090 -1300 122150 -1240
rect 122170 -1300 122230 -1240
rect 122250 -1300 122310 -1240
rect 122090 -1380 122150 -1320
rect 122170 -1380 122230 -1320
rect 122250 -1380 122310 -1320
rect 122790 -1220 122850 -1160
rect 122870 -1220 122930 -1160
rect 122950 -1220 123010 -1160
rect 122790 -1300 122850 -1240
rect 122870 -1300 122930 -1240
rect 122950 -1300 123010 -1240
rect 122790 -1380 122850 -1320
rect 122870 -1380 122930 -1320
rect 122950 -1380 123010 -1320
<< metal2 >>
rect 109490 9980 118110 9990
rect 109550 9920 109610 9980
rect 109670 9920 109730 9980
rect 109790 9920 109850 9980
rect 109910 9920 109970 9980
rect 110030 9920 110090 9980
rect 110150 9920 110210 9980
rect 110270 9920 110330 9980
rect 110390 9920 110450 9980
rect 110510 9920 110570 9980
rect 110630 9920 114910 9980
rect 114970 9920 116970 9980
rect 117030 9920 117090 9980
rect 117150 9920 117210 9980
rect 117270 9920 117330 9980
rect 117390 9920 117450 9980
rect 117510 9920 117570 9980
rect 117630 9920 117690 9980
rect 117750 9920 117810 9980
rect 117870 9920 117930 9980
rect 117990 9920 118050 9980
rect 109490 9910 118110 9920
rect 109420 9870 110700 9880
rect 109420 9810 109430 9870
rect 109490 9810 109670 9870
rect 109730 9810 109910 9870
rect 109970 9810 110150 9870
rect 110210 9810 110390 9870
rect 110450 9810 110630 9870
rect 110690 9810 110700 9870
rect 109420 9800 110700 9810
rect 112210 9870 112290 9880
rect 112210 9810 112220 9870
rect 112280 9860 112290 9870
rect 113150 9870 113230 9880
rect 113150 9860 113160 9870
rect 112280 9810 113160 9860
rect 113220 9810 113230 9870
rect 112210 9800 112290 9810
rect 113150 9800 113230 9810
rect 114370 9870 114450 9880
rect 114370 9810 114380 9870
rect 114440 9860 114450 9870
rect 115310 9870 115390 9880
rect 115310 9860 115320 9870
rect 114440 9810 115320 9860
rect 115380 9810 115390 9870
rect 114370 9800 114450 9810
rect 115310 9800 115390 9810
rect 116900 9870 118180 9880
rect 116900 9810 116910 9870
rect 116970 9810 117150 9870
rect 117210 9810 117390 9870
rect 117450 9810 117630 9870
rect 117690 9810 117870 9870
rect 117930 9810 118110 9870
rect 118170 9810 118180 9870
rect 116900 9800 118180 9810
rect 113680 9760 114690 9770
rect 113680 9700 113690 9760
rect 113750 9700 113770 9760
rect 113830 9700 113850 9760
rect 113910 9700 114260 9760
rect 114320 9700 114500 9760
rect 114560 9700 114620 9760
rect 114680 9700 114690 9760
rect 113680 9680 114690 9700
rect 113680 9620 113690 9680
rect 113750 9620 113770 9680
rect 113830 9620 113850 9680
rect 113910 9620 114260 9680
rect 114320 9620 114500 9680
rect 114560 9620 114620 9680
rect 114680 9620 114690 9680
rect 111970 9600 112050 9610
rect 111970 9540 111980 9600
rect 112040 9590 112050 9600
rect 112210 9600 112290 9610
rect 112210 9590 112220 9600
rect 112040 9550 112220 9590
rect 112040 9540 112050 9550
rect 111970 9530 112050 9540
rect 112210 9540 112220 9550
rect 112280 9590 112290 9600
rect 112330 9600 112410 9610
rect 112330 9590 112340 9600
rect 112280 9550 112340 9590
rect 112280 9540 112290 9550
rect 112210 9530 112290 9540
rect 112330 9540 112340 9550
rect 112400 9540 112410 9600
rect 112330 9530 112410 9540
rect 113680 9600 114690 9620
rect 113680 9540 113690 9600
rect 113750 9540 113770 9600
rect 113830 9540 113850 9600
rect 113910 9540 114260 9600
rect 114320 9540 114500 9600
rect 114560 9540 114620 9600
rect 114680 9540 114690 9600
rect 113680 9530 114690 9540
rect 115190 9600 115270 9610
rect 115190 9540 115200 9600
rect 115260 9590 115270 9600
rect 115310 9600 115390 9610
rect 115310 9590 115320 9600
rect 115260 9550 115320 9590
rect 115260 9540 115270 9550
rect 115190 9530 115270 9540
rect 115310 9540 115320 9550
rect 115380 9590 115390 9600
rect 115550 9600 115630 9610
rect 115550 9590 115560 9600
rect 115380 9550 115560 9590
rect 115380 9540 115390 9550
rect 115310 9530 115390 9540
rect 115550 9540 115560 9550
rect 115620 9540 115630 9600
rect 115550 9530 115630 9540
rect 112910 9420 113920 9430
rect 112910 9360 112920 9420
rect 112980 9360 113040 9420
rect 113100 9360 113280 9420
rect 113340 9360 113690 9420
rect 113750 9360 113770 9420
rect 113830 9360 113850 9420
rect 113910 9360 113920 9420
rect 104580 9340 108320 9350
rect 104580 9280 104590 9340
rect 104650 9280 104670 9340
rect 104730 9280 104750 9340
rect 104810 9280 105290 9340
rect 105350 9280 105370 9340
rect 105430 9280 105450 9340
rect 105510 9280 105990 9340
rect 106050 9280 106070 9340
rect 106130 9280 106150 9340
rect 106210 9280 106690 9340
rect 106750 9280 106770 9340
rect 106830 9280 106850 9340
rect 106910 9280 108090 9340
rect 108150 9280 108170 9340
rect 108230 9280 108250 9340
rect 108310 9280 108320 9340
rect 104580 9260 108320 9280
rect 104580 9200 104590 9260
rect 104650 9200 104670 9260
rect 104730 9200 104750 9260
rect 104810 9200 105290 9260
rect 105350 9200 105370 9260
rect 105430 9200 105450 9260
rect 105510 9200 105990 9260
rect 106050 9200 106070 9260
rect 106130 9200 106150 9260
rect 106210 9200 106690 9260
rect 106750 9200 106770 9260
rect 106830 9200 106850 9260
rect 106910 9200 108090 9260
rect 108150 9200 108170 9260
rect 108230 9200 108250 9260
rect 108310 9200 108320 9260
rect 104580 9180 108320 9200
rect 112910 9340 113920 9360
rect 112910 9280 112920 9340
rect 112980 9280 113040 9340
rect 113100 9280 113280 9340
rect 113340 9280 113690 9340
rect 113750 9280 113770 9340
rect 113830 9280 113850 9340
rect 113910 9280 113920 9340
rect 112910 9260 113920 9280
rect 112910 9200 112920 9260
rect 112980 9200 113040 9260
rect 113100 9200 113280 9260
rect 113340 9200 113690 9260
rect 113750 9200 113770 9260
rect 113830 9200 113850 9260
rect 113910 9200 113920 9260
rect 112910 9190 113920 9200
rect 119280 9340 123020 9350
rect 119280 9280 119290 9340
rect 119350 9280 119370 9340
rect 119430 9280 119450 9340
rect 119510 9280 120690 9340
rect 120750 9280 120770 9340
rect 120830 9280 120850 9340
rect 120910 9280 121390 9340
rect 121450 9280 121470 9340
rect 121530 9280 121550 9340
rect 121610 9280 122090 9340
rect 122150 9280 122170 9340
rect 122230 9280 122250 9340
rect 122310 9280 122790 9340
rect 122850 9280 122870 9340
rect 122930 9280 122950 9340
rect 123010 9280 123020 9340
rect 119280 9260 123020 9280
rect 119280 9200 119290 9260
rect 119350 9200 119370 9260
rect 119430 9200 119450 9260
rect 119510 9200 120690 9260
rect 120750 9200 120770 9260
rect 120830 9200 120850 9260
rect 120910 9200 121390 9260
rect 121450 9200 121470 9260
rect 121530 9200 121550 9260
rect 121610 9200 122090 9260
rect 122150 9200 122170 9260
rect 122230 9200 122250 9260
rect 122310 9200 122790 9260
rect 122850 9200 122870 9260
rect 122930 9200 122950 9260
rect 123010 9200 123020 9260
rect 104580 9120 104590 9180
rect 104650 9120 104670 9180
rect 104730 9120 104750 9180
rect 104810 9120 105290 9180
rect 105350 9120 105370 9180
rect 105430 9120 105450 9180
rect 105510 9120 105990 9180
rect 106050 9120 106070 9180
rect 106130 9120 106150 9180
rect 106210 9120 106690 9180
rect 106750 9120 106770 9180
rect 106830 9120 106850 9180
rect 106910 9120 108090 9180
rect 108150 9120 108170 9180
rect 108230 9120 108250 9180
rect 108310 9120 108320 9180
rect 104580 9110 108320 9120
rect 119280 9180 123020 9200
rect 119280 9120 119290 9180
rect 119350 9120 119370 9180
rect 119430 9120 119450 9180
rect 119510 9120 120690 9180
rect 120750 9120 120770 9180
rect 120830 9120 120850 9180
rect 120910 9120 121390 9180
rect 121450 9120 121470 9180
rect 121530 9120 121550 9180
rect 121610 9120 122090 9180
rect 122150 9120 122170 9180
rect 122230 9120 122250 9180
rect 122310 9120 122790 9180
rect 122850 9120 122870 9180
rect 122930 9120 122950 9180
rect 123010 9120 123020 9180
rect 119280 9110 123020 9120
rect 109300 9060 111310 9070
rect 109300 9000 109310 9060
rect 109370 9000 109550 9060
rect 109610 9000 109790 9060
rect 109850 9000 110030 9060
rect 110090 9000 110270 9060
rect 110330 9000 110510 9060
rect 110570 9000 110750 9060
rect 110810 9000 111080 9060
rect 111140 9000 111160 9060
rect 111220 9000 111240 9060
rect 111300 9000 111310 9060
rect 109300 8990 111310 9000
rect 116290 9060 118300 9070
rect 116290 9000 116300 9060
rect 116360 9000 116380 9060
rect 116440 9000 116460 9060
rect 116520 9000 116790 9060
rect 116850 9000 117030 9060
rect 117090 9000 117270 9060
rect 117330 9000 117510 9060
rect 117570 9000 117750 9060
rect 117810 9000 117990 9060
rect 118050 9000 118230 9060
rect 118290 9000 118300 9060
rect 116290 8990 118300 9000
rect 109180 8950 110700 8960
rect 109180 8890 109190 8950
rect 109250 8890 109430 8950
rect 109490 8890 109670 8950
rect 109730 8890 109910 8950
rect 109970 8890 110150 8950
rect 110210 8890 110390 8950
rect 110450 8890 110630 8950
rect 110690 8890 110700 8950
rect 109180 8870 110700 8890
rect 109180 8810 109190 8870
rect 109250 8810 109430 8870
rect 109490 8810 109670 8870
rect 109730 8810 109910 8870
rect 109970 8810 110150 8870
rect 110210 8810 110390 8870
rect 110450 8810 110630 8870
rect 110690 8810 110700 8870
rect 109180 8790 110700 8810
rect 116900 8950 118420 8960
rect 116900 8890 116910 8950
rect 116970 8890 117150 8950
rect 117210 8890 117390 8950
rect 117450 8890 117630 8950
rect 117690 8890 117870 8950
rect 117930 8890 118110 8950
rect 118170 8890 118350 8950
rect 118410 8890 118420 8950
rect 116900 8870 118420 8890
rect 116900 8810 116910 8870
rect 116970 8810 117150 8870
rect 117210 8810 117390 8870
rect 117450 8810 117630 8870
rect 117690 8810 117870 8870
rect 117930 8810 118110 8870
rect 118170 8810 118350 8870
rect 118410 8810 118420 8870
rect 109180 8730 109190 8790
rect 109250 8730 109430 8790
rect 109490 8730 109670 8790
rect 109730 8730 109910 8790
rect 109970 8730 110150 8790
rect 110210 8730 110390 8790
rect 110450 8730 110630 8790
rect 110690 8730 110700 8790
rect 109180 8710 110700 8730
rect 112210 8790 112290 8800
rect 112210 8730 112220 8790
rect 112280 8780 112290 8790
rect 113150 8790 113230 8800
rect 113150 8780 113160 8790
rect 112280 8740 113160 8780
rect 112280 8730 112290 8740
rect 112210 8720 112290 8730
rect 113150 8730 113160 8740
rect 113220 8730 113230 8790
rect 113150 8720 113230 8730
rect 114370 8790 114450 8800
rect 114370 8730 114380 8790
rect 114440 8780 114450 8790
rect 115310 8790 115390 8800
rect 115310 8780 115320 8790
rect 114440 8740 115320 8780
rect 114440 8730 114450 8740
rect 114370 8720 114450 8730
rect 115310 8730 115320 8740
rect 115380 8730 115390 8790
rect 115310 8720 115390 8730
rect 116900 8790 118420 8810
rect 116900 8730 116910 8790
rect 116970 8730 117150 8790
rect 117210 8730 117390 8790
rect 117450 8730 117630 8790
rect 117690 8730 117870 8790
rect 117930 8730 118110 8790
rect 118170 8730 118350 8790
rect 118410 8730 118420 8790
rect 109180 8650 109190 8710
rect 109250 8650 109430 8710
rect 109490 8650 109670 8710
rect 109730 8650 109910 8710
rect 109970 8650 110150 8710
rect 110210 8650 110390 8710
rect 110450 8650 110630 8710
rect 110690 8650 110700 8710
rect 116900 8710 118420 8730
rect 109180 8630 110700 8650
rect 109180 8570 109190 8630
rect 109250 8570 109430 8630
rect 109490 8570 109670 8630
rect 109730 8570 109910 8630
rect 109970 8570 110150 8630
rect 110210 8570 110390 8630
rect 110450 8570 110630 8630
rect 110690 8570 110700 8630
rect 111340 8680 111420 8690
rect 111340 8620 111350 8680
rect 111410 8670 111420 8680
rect 112100 8680 112180 8690
rect 112100 8670 112110 8680
rect 111410 8630 112110 8670
rect 111410 8620 111420 8630
rect 111340 8610 111420 8620
rect 112100 8620 112110 8630
rect 112170 8670 112180 8680
rect 113060 8680 113120 8690
rect 112170 8630 113060 8670
rect 112170 8620 112180 8630
rect 112100 8610 112180 8620
rect 115352 8680 115412 8690
rect 113120 8630 115352 8670
rect 113060 8610 113120 8620
rect 116180 8680 116260 8690
rect 116180 8670 116190 8680
rect 115412 8630 116190 8670
rect 115352 8610 115412 8620
rect 116180 8620 116190 8630
rect 116250 8620 116260 8680
rect 116180 8610 116260 8620
rect 116900 8650 116910 8710
rect 116970 8650 117150 8710
rect 117210 8650 117390 8710
rect 117450 8650 117630 8710
rect 117690 8650 117870 8710
rect 117930 8650 118110 8710
rect 118170 8650 118350 8710
rect 118410 8650 118420 8710
rect 116900 8630 118420 8650
rect 109180 8550 110700 8570
rect 109180 8490 109190 8550
rect 109250 8490 109430 8550
rect 109490 8490 109670 8550
rect 109730 8490 109910 8550
rect 109970 8490 110150 8550
rect 110210 8490 110390 8550
rect 110450 8490 110630 8550
rect 110690 8490 110700 8550
rect 114470 8570 115510 8580
rect 114470 8510 114480 8570
rect 114540 8510 114910 8570
rect 114970 8510 115440 8570
rect 115500 8510 115510 8570
rect 114470 8500 115510 8510
rect 116900 8570 116910 8630
rect 116970 8570 117150 8630
rect 117210 8570 117390 8630
rect 117450 8570 117630 8630
rect 117690 8570 117870 8630
rect 117930 8570 118110 8630
rect 118170 8570 118350 8630
rect 118410 8570 118420 8630
rect 116900 8550 118420 8570
rect 109180 8470 110700 8490
rect 116900 8490 116910 8550
rect 116970 8490 117150 8550
rect 117210 8490 117390 8550
rect 117450 8490 117630 8550
rect 117690 8490 117870 8550
rect 117930 8490 118110 8550
rect 118170 8490 118350 8550
rect 118410 8490 118420 8550
rect 116900 8470 118420 8490
rect 109180 8410 109190 8470
rect 109250 8410 109430 8470
rect 109490 8410 109670 8470
rect 109730 8410 109910 8470
rect 109970 8410 110150 8470
rect 110210 8410 110390 8470
rect 110450 8410 110630 8470
rect 110690 8410 110700 8470
rect 109180 8400 110700 8410
rect 111070 8460 116530 8470
rect 111070 8400 111080 8460
rect 111140 8400 111160 8460
rect 111220 8400 111240 8460
rect 111300 8400 113030 8460
rect 113090 8400 113360 8460
rect 113420 8400 113690 8460
rect 113750 8400 113850 8460
rect 113910 8400 114180 8460
rect 114240 8400 114510 8460
rect 114570 8400 116300 8460
rect 116360 8400 116380 8460
rect 116440 8400 116460 8460
rect 116520 8400 116530 8460
rect 116900 8410 116910 8470
rect 116970 8410 117150 8470
rect 117210 8410 117390 8470
rect 117450 8410 117630 8470
rect 117690 8410 117870 8470
rect 117930 8410 118110 8470
rect 118170 8410 118350 8470
rect 118410 8410 118420 8470
rect 116900 8400 118420 8410
rect 111070 8380 116530 8400
rect 109300 8350 110580 8360
rect 109300 8290 109310 8350
rect 109370 8290 109550 8350
rect 109610 8290 109790 8350
rect 109850 8290 110030 8350
rect 110090 8290 110270 8350
rect 110330 8290 110510 8350
rect 110570 8290 110580 8350
rect 109300 8280 110580 8290
rect 111070 8320 111080 8380
rect 111140 8320 111160 8380
rect 111220 8320 111240 8380
rect 111300 8320 113030 8380
rect 113090 8320 113360 8380
rect 113420 8320 113690 8380
rect 113750 8320 113850 8380
rect 113910 8320 114180 8380
rect 114240 8320 114510 8380
rect 114570 8320 116300 8380
rect 116360 8320 116380 8380
rect 116440 8320 116460 8380
rect 116520 8320 116530 8380
rect 111070 8300 116530 8320
rect 111070 8240 111080 8300
rect 111140 8240 111160 8300
rect 111220 8240 111240 8300
rect 111300 8240 113030 8300
rect 113090 8240 113360 8300
rect 113420 8240 113690 8300
rect 113750 8240 113850 8300
rect 113910 8240 114180 8300
rect 114240 8240 114510 8300
rect 114570 8240 116300 8300
rect 116360 8240 116380 8300
rect 116440 8240 116460 8300
rect 116520 8240 116530 8300
rect 117020 8350 118300 8360
rect 117020 8290 117030 8350
rect 117090 8290 117270 8350
rect 117330 8290 117510 8350
rect 117570 8290 117750 8350
rect 117810 8290 117990 8350
rect 118050 8290 118230 8350
rect 118290 8290 118300 8350
rect 117020 8280 118300 8290
rect 111070 8230 116530 8240
rect 113240 8170 113320 8180
rect 113240 8110 113250 8170
rect 113310 8160 113320 8170
rect 113460 8170 113540 8180
rect 113460 8160 113470 8170
rect 113310 8120 113470 8160
rect 113310 8110 113320 8120
rect 113240 8100 113320 8110
rect 113460 8110 113470 8120
rect 113530 8110 113540 8170
rect 113460 8100 113540 8110
rect 114060 8170 114140 8180
rect 114060 8110 114070 8170
rect 114130 8160 114140 8170
rect 114280 8170 114360 8180
rect 114280 8160 114290 8170
rect 114130 8120 114290 8160
rect 114130 8110 114140 8120
rect 114060 8100 114140 8110
rect 114280 8110 114290 8120
rect 114350 8110 114360 8170
rect 114280 8100 114360 8110
rect 108510 7670 108590 7680
rect 108510 7610 108520 7670
rect 108580 7610 108590 7670
rect 108510 7600 108590 7610
rect 119010 7670 119090 7680
rect 119010 7610 119020 7670
rect 119080 7610 119090 7670
rect 119010 7600 119090 7610
rect 109300 7570 111040 7580
rect 109300 7510 109310 7570
rect 109370 7510 109550 7570
rect 109610 7510 109790 7570
rect 109850 7510 110030 7570
rect 110090 7510 110270 7570
rect 110330 7510 110510 7570
rect 110570 7510 110810 7570
rect 110870 7510 110890 7570
rect 110950 7510 110970 7570
rect 111030 7510 111040 7570
rect 116560 7570 118300 7580
rect 109300 7500 111040 7510
rect 113120 7550 113180 7560
rect 113600 7550 113660 7560
rect 113350 7530 113430 7540
rect 113350 7520 113360 7530
rect 113180 7490 113360 7520
rect 113120 7480 113360 7490
rect 113350 7470 113360 7480
rect 113420 7520 113430 7530
rect 113420 7490 113600 7520
rect 114170 7530 114250 7540
rect 114170 7520 114180 7530
rect 113660 7490 114180 7520
rect 113420 7480 114180 7490
rect 113420 7470 113430 7480
rect 109370 7460 109430 7470
rect 109490 7460 109550 7470
rect 109430 7410 109490 7450
rect 109370 7390 109430 7400
rect 109610 7460 109670 7470
rect 109550 7410 109610 7450
rect 109490 7390 109550 7400
rect 109730 7460 109790 7470
rect 109670 7410 109730 7450
rect 109610 7390 109670 7400
rect 109850 7460 109910 7470
rect 109790 7410 109850 7450
rect 109730 7390 109790 7400
rect 109970 7460 110030 7470
rect 109910 7410 109970 7450
rect 109850 7390 109910 7400
rect 110090 7460 110150 7470
rect 110030 7410 110090 7450
rect 109970 7390 110030 7400
rect 110210 7460 110270 7470
rect 110150 7410 110210 7450
rect 110090 7390 110150 7400
rect 110330 7460 110390 7470
rect 110270 7410 110330 7450
rect 110210 7390 110270 7400
rect 110450 7460 110510 7470
rect 110390 7410 110450 7450
rect 110330 7390 110390 7400
rect 111340 7460 111420 7470
rect 113350 7460 113430 7470
rect 114170 7470 114180 7480
rect 114240 7520 114250 7530
rect 114240 7480 114260 7520
rect 116560 7510 116570 7570
rect 116630 7510 116650 7570
rect 116710 7510 116730 7570
rect 116790 7510 117030 7570
rect 117090 7510 117270 7570
rect 117330 7510 117510 7570
rect 117570 7510 117750 7570
rect 117810 7510 117990 7570
rect 118050 7510 118230 7570
rect 118290 7510 118300 7570
rect 116560 7500 118300 7510
rect 114240 7470 114250 7480
rect 114170 7460 114250 7470
rect 116180 7460 116260 7470
rect 111340 7450 111350 7460
rect 110510 7410 111350 7450
rect 110450 7390 110510 7400
rect 111340 7400 111350 7410
rect 111410 7400 111420 7460
rect 113200 7410 113280 7420
rect 113200 7400 113210 7410
rect 111340 7390 111420 7400
rect 112730 7360 113210 7400
rect 108080 7350 111310 7360
rect 108080 7290 108090 7350
rect 108150 7290 108170 7350
rect 108230 7290 108250 7350
rect 108310 7290 109250 7350
rect 109310 7290 109470 7350
rect 109530 7290 109690 7350
rect 109750 7290 109910 7350
rect 109970 7290 110130 7350
rect 110190 7290 110350 7350
rect 110410 7290 110570 7350
rect 110630 7290 111080 7350
rect 111140 7290 111160 7350
rect 111220 7290 111240 7350
rect 111300 7290 111310 7350
rect 113200 7350 113210 7360
rect 113270 7400 113280 7410
rect 114320 7410 114400 7420
rect 114320 7400 114330 7410
rect 113270 7360 114330 7400
rect 113270 7350 113280 7360
rect 113200 7340 113280 7350
rect 114320 7350 114330 7360
rect 114390 7350 114400 7410
rect 116180 7400 116190 7460
rect 116250 7450 116260 7460
rect 117090 7460 117150 7470
rect 116250 7410 117090 7450
rect 116250 7400 116260 7410
rect 116180 7390 116260 7400
rect 117210 7460 117270 7470
rect 117150 7410 117210 7450
rect 117090 7390 117150 7400
rect 117330 7460 117390 7470
rect 117270 7410 117330 7450
rect 117210 7390 117270 7400
rect 117450 7460 117510 7470
rect 117390 7410 117450 7450
rect 117330 7390 117390 7400
rect 117570 7460 117630 7470
rect 117510 7410 117570 7450
rect 117450 7390 117510 7400
rect 117690 7460 117750 7470
rect 117630 7410 117690 7450
rect 117570 7390 117630 7400
rect 117810 7460 117870 7470
rect 117750 7410 117810 7450
rect 117690 7390 117750 7400
rect 117930 7460 117990 7470
rect 117870 7410 117930 7450
rect 117810 7390 117870 7400
rect 118050 7460 118110 7470
rect 117990 7410 118050 7450
rect 117930 7390 117990 7400
rect 118170 7460 118230 7470
rect 118110 7410 118170 7450
rect 118050 7390 118110 7400
rect 118170 7390 118230 7400
rect 114320 7340 114400 7350
rect 116290 7350 119520 7360
rect 108080 7270 111310 7290
rect 108080 7210 108090 7270
rect 108150 7210 108170 7270
rect 108230 7210 108250 7270
rect 108310 7210 109250 7270
rect 109310 7210 109470 7270
rect 109530 7210 109690 7270
rect 109750 7210 109910 7270
rect 109970 7210 110130 7270
rect 110190 7210 110350 7270
rect 110410 7210 110570 7270
rect 110630 7210 111080 7270
rect 111140 7210 111160 7270
rect 111220 7210 111240 7270
rect 111300 7210 111310 7270
rect 111900 7290 111980 7300
rect 111900 7230 111910 7290
rect 111970 7280 111980 7290
rect 113490 7290 113570 7300
rect 113490 7280 113500 7290
rect 111970 7240 113500 7280
rect 111970 7230 111980 7240
rect 111900 7220 111980 7230
rect 113490 7230 113500 7240
rect 113560 7280 113570 7290
rect 114030 7290 114110 7300
rect 114030 7280 114040 7290
rect 113560 7240 114040 7280
rect 113560 7230 113570 7240
rect 113490 7220 113570 7230
rect 114030 7230 114040 7240
rect 114100 7280 114110 7290
rect 115630 7290 115710 7300
rect 115630 7280 115640 7290
rect 114100 7240 115640 7280
rect 114100 7230 114110 7240
rect 114030 7220 114110 7230
rect 115630 7230 115640 7240
rect 115700 7230 115710 7290
rect 115630 7220 115710 7230
rect 116290 7290 116300 7350
rect 116360 7290 116380 7350
rect 116440 7290 116460 7350
rect 116520 7290 116970 7350
rect 117030 7290 117190 7350
rect 117250 7290 117410 7350
rect 117470 7290 117630 7350
rect 117690 7290 117850 7350
rect 117910 7290 118070 7350
rect 118130 7290 118290 7350
rect 118350 7290 119290 7350
rect 119350 7290 119370 7350
rect 119430 7290 119450 7350
rect 119510 7290 119520 7350
rect 116290 7270 119520 7290
rect 108080 7190 111310 7210
rect 116290 7210 116300 7270
rect 116360 7210 116380 7270
rect 116440 7210 116460 7270
rect 116520 7210 116970 7270
rect 117030 7210 117190 7270
rect 117250 7210 117410 7270
rect 117470 7210 117630 7270
rect 117690 7210 117850 7270
rect 117910 7210 118070 7270
rect 118130 7210 118290 7270
rect 118350 7210 119290 7270
rect 119350 7210 119370 7270
rect 119430 7210 119450 7270
rect 119510 7210 119520 7270
rect 116290 7190 119520 7210
rect 108080 7130 108090 7190
rect 108150 7130 108170 7190
rect 108230 7130 108250 7190
rect 108310 7130 109250 7190
rect 109310 7130 109470 7190
rect 109530 7130 109690 7190
rect 109750 7130 109910 7190
rect 109970 7130 110130 7190
rect 110190 7130 110350 7190
rect 110410 7130 110570 7190
rect 110630 7130 111080 7190
rect 111140 7130 111160 7190
rect 111220 7130 111240 7190
rect 111300 7130 111310 7190
rect 108080 7120 111310 7130
rect 113700 7180 113780 7190
rect 113700 7120 113710 7180
rect 113770 7170 113780 7180
rect 113920 7180 114000 7190
rect 113920 7170 113930 7180
rect 113770 7130 113930 7170
rect 113770 7120 113780 7130
rect 113700 7110 113780 7120
rect 113920 7120 113930 7130
rect 113990 7120 114000 7180
rect 116290 7130 116300 7190
rect 116360 7130 116380 7190
rect 116440 7130 116460 7190
rect 116520 7130 116970 7190
rect 117030 7130 117190 7190
rect 117250 7130 117410 7190
rect 117470 7130 117630 7190
rect 117690 7130 117850 7190
rect 117910 7130 118070 7190
rect 118130 7130 118290 7190
rect 118350 7130 119290 7190
rect 119350 7130 119370 7190
rect 119430 7130 119450 7190
rect 119510 7130 119520 7190
rect 116290 7120 119520 7130
rect 113920 7110 114000 7120
rect 113870 7070 113950 7080
rect 113870 7010 113880 7070
rect 113940 7060 113950 7070
rect 114420 7070 114500 7080
rect 114420 7060 114430 7070
rect 113940 7020 114430 7060
rect 113940 7010 113950 7020
rect 109350 7000 109430 7010
rect 109350 6940 109360 7000
rect 109420 6990 109430 7000
rect 109570 7000 109650 7010
rect 109570 6990 109580 7000
rect 109420 6950 109580 6990
rect 109420 6940 109430 6950
rect 109350 6930 109430 6940
rect 109570 6940 109580 6950
rect 109640 6990 109650 7000
rect 109790 7000 109870 7010
rect 109790 6990 109800 7000
rect 109640 6950 109800 6990
rect 109640 6940 109650 6950
rect 109570 6930 109650 6940
rect 109790 6940 109800 6950
rect 109860 6990 109870 7000
rect 110010 7000 110090 7010
rect 110010 6990 110020 7000
rect 109860 6950 110020 6990
rect 109860 6940 109870 6950
rect 109790 6930 109870 6940
rect 110010 6940 110020 6950
rect 110080 6990 110090 7000
rect 110230 7000 110310 7010
rect 110230 6990 110240 7000
rect 110080 6950 110240 6990
rect 110080 6940 110090 6950
rect 110010 6930 110090 6940
rect 110230 6940 110240 6950
rect 110300 6990 110310 7000
rect 110450 7000 110530 7010
rect 113870 7000 113950 7010
rect 114420 7010 114430 7020
rect 114490 7060 114500 7070
rect 115720 7070 115800 7080
rect 115720 7060 115730 7070
rect 114490 7020 115730 7060
rect 114490 7010 114500 7020
rect 114420 7000 114500 7010
rect 115720 7010 115730 7020
rect 115790 7010 115800 7070
rect 115720 7000 115800 7010
rect 117070 7000 117150 7010
rect 110450 6990 110460 7000
rect 110300 6950 110460 6990
rect 110300 6940 110310 6950
rect 110230 6930 110310 6940
rect 110450 6940 110460 6950
rect 110520 6940 110530 7000
rect 110450 6930 110530 6940
rect 110800 6960 113350 6970
rect 110800 6900 110810 6960
rect 110870 6900 110890 6960
rect 110950 6900 110970 6960
rect 111030 6900 112180 6960
rect 112240 6900 112290 6960
rect 112350 6900 112400 6960
rect 112460 6900 112510 6960
rect 112570 6900 112620 6960
rect 112680 6900 112730 6960
rect 112790 6900 112840 6960
rect 112900 6900 112950 6960
rect 113010 6900 113060 6960
rect 113120 6900 113170 6960
rect 113230 6900 113280 6960
rect 113340 6900 113350 6960
rect 110800 6880 113350 6900
rect 113700 6960 113780 6970
rect 113700 6900 113710 6960
rect 113770 6900 113780 6960
rect 113700 6890 113780 6900
rect 114250 6960 116800 6970
rect 114250 6900 114260 6960
rect 114320 6900 114370 6960
rect 114430 6900 114480 6960
rect 114540 6900 114590 6960
rect 114650 6900 114700 6960
rect 114760 6900 114810 6960
rect 114870 6900 114920 6960
rect 114980 6900 115030 6960
rect 115090 6900 115140 6960
rect 115200 6900 115250 6960
rect 115310 6900 115360 6960
rect 115420 6900 116570 6960
rect 116630 6900 116650 6960
rect 116710 6900 116730 6960
rect 116790 6900 116800 6960
rect 117070 6940 117080 7000
rect 117140 6990 117150 7000
rect 117290 7000 117370 7010
rect 117290 6990 117300 7000
rect 117140 6950 117300 6990
rect 117140 6940 117150 6950
rect 117070 6930 117150 6940
rect 117290 6940 117300 6950
rect 117360 6990 117370 7000
rect 117510 7000 117590 7010
rect 117510 6990 117520 7000
rect 117360 6950 117520 6990
rect 117360 6940 117370 6950
rect 117290 6930 117370 6940
rect 117510 6940 117520 6950
rect 117580 6990 117590 7000
rect 117730 7000 117810 7010
rect 117730 6990 117740 7000
rect 117580 6950 117740 6990
rect 117580 6940 117590 6950
rect 117510 6930 117590 6940
rect 117730 6940 117740 6950
rect 117800 6990 117810 7000
rect 117950 7000 118030 7010
rect 117950 6990 117960 7000
rect 117800 6950 117960 6990
rect 117800 6940 117810 6950
rect 117730 6930 117810 6940
rect 117950 6940 117960 6950
rect 118020 6990 118030 7000
rect 118170 7000 118250 7010
rect 118170 6990 118180 7000
rect 118020 6950 118180 6990
rect 118020 6940 118030 6950
rect 117950 6930 118030 6940
rect 118170 6940 118180 6950
rect 118240 6940 118250 7000
rect 118170 6930 118250 6940
rect 110800 6820 110810 6880
rect 110870 6820 110890 6880
rect 110950 6820 110970 6880
rect 111030 6820 112180 6880
rect 112240 6820 112290 6880
rect 112350 6820 112400 6880
rect 112460 6820 112510 6880
rect 112570 6820 112620 6880
rect 112680 6820 112730 6880
rect 112790 6820 112840 6880
rect 112900 6820 112950 6880
rect 113010 6820 113060 6880
rect 113120 6820 113170 6880
rect 113230 6820 113280 6880
rect 113340 6820 113350 6880
rect 110800 6800 113350 6820
rect 110800 6740 110810 6800
rect 110870 6740 110890 6800
rect 110950 6740 110970 6800
rect 111030 6740 112180 6800
rect 112240 6740 112290 6800
rect 112350 6740 112400 6800
rect 112460 6740 112510 6800
rect 112570 6740 112620 6800
rect 112680 6740 112730 6800
rect 112790 6740 112840 6800
rect 112900 6740 112950 6800
rect 113010 6740 113060 6800
rect 113120 6740 113170 6800
rect 113230 6740 113280 6800
rect 113340 6740 113350 6800
rect 110800 6730 113350 6740
rect 114250 6880 116800 6900
rect 114250 6820 114260 6880
rect 114320 6820 114370 6880
rect 114430 6820 114480 6880
rect 114540 6820 114590 6880
rect 114650 6820 114700 6880
rect 114760 6820 114810 6880
rect 114870 6820 114920 6880
rect 114980 6820 115030 6880
rect 115090 6820 115140 6880
rect 115200 6820 115250 6880
rect 115310 6820 115360 6880
rect 115420 6820 116570 6880
rect 116630 6820 116650 6880
rect 116710 6820 116730 6880
rect 116790 6820 116800 6880
rect 114250 6800 116800 6820
rect 114250 6740 114260 6800
rect 114320 6740 114370 6800
rect 114430 6740 114480 6800
rect 114540 6740 114590 6800
rect 114650 6740 114700 6800
rect 114760 6740 114810 6800
rect 114870 6740 114920 6800
rect 114980 6740 115030 6800
rect 115090 6740 115140 6800
rect 115200 6740 115250 6800
rect 115310 6740 115360 6800
rect 115420 6740 116570 6800
rect 116630 6740 116650 6800
rect 116710 6740 116730 6800
rect 116790 6740 116800 6800
rect 114250 6730 116800 6740
rect 111340 6320 116260 6330
rect 111340 6260 111350 6320
rect 111410 6260 111430 6320
rect 111490 6260 111510 6320
rect 111570 6260 113550 6320
rect 113610 6260 113770 6320
rect 113830 6260 113990 6320
rect 114050 6260 116030 6320
rect 116090 6260 116110 6320
rect 116170 6260 116190 6320
rect 116250 6260 116260 6320
rect 111340 6240 116260 6260
rect 111340 6180 111350 6240
rect 111410 6180 111430 6240
rect 111490 6180 111510 6240
rect 111570 6180 113550 6240
rect 113610 6180 113770 6240
rect 113830 6180 113990 6240
rect 114050 6180 116030 6240
rect 116090 6180 116110 6240
rect 116170 6180 116190 6240
rect 116250 6180 116260 6240
rect 111340 6160 116260 6180
rect 111340 6100 111350 6160
rect 111410 6100 111430 6160
rect 111490 6100 111510 6160
rect 111570 6100 113550 6160
rect 113610 6100 113770 6160
rect 113830 6100 113990 6160
rect 114050 6100 116030 6160
rect 116090 6100 116110 6160
rect 116170 6100 116190 6160
rect 116250 6100 116260 6160
rect 111340 6090 116260 6100
rect 111340 6020 111580 6030
rect 111340 5960 111350 6020
rect 111410 5960 111430 6020
rect 111490 5960 111510 6020
rect 111570 5960 111580 6020
rect 111340 5940 111580 5960
rect 116020 6020 116260 6030
rect 116020 5960 116030 6020
rect 116090 5960 116110 6020
rect 116170 5960 116190 6020
rect 116250 5960 116260 6020
rect 111340 5880 111350 5940
rect 111410 5880 111430 5940
rect 111490 5880 111510 5940
rect 111570 5880 111580 5940
rect 111340 5860 111580 5880
rect 112170 5940 113650 5950
rect 112170 5880 112180 5940
rect 112240 5880 112400 5940
rect 112460 5880 112620 5940
rect 112680 5880 112840 5940
rect 112900 5880 113060 5940
rect 113120 5880 113280 5940
rect 113340 5880 113580 5940
rect 113640 5880 113650 5940
rect 112170 5870 113650 5880
rect 113950 5940 115430 5950
rect 113950 5880 113960 5940
rect 114020 5880 114260 5940
rect 114320 5880 114480 5940
rect 114540 5880 114700 5940
rect 114760 5880 114920 5940
rect 114980 5880 115140 5940
rect 115200 5880 115360 5940
rect 115420 5880 115430 5940
rect 113950 5870 115430 5880
rect 116020 5940 116260 5960
rect 116020 5880 116030 5940
rect 116090 5880 116110 5940
rect 116170 5880 116190 5940
rect 116250 5880 116260 5940
rect 111340 5800 111350 5860
rect 111410 5800 111430 5860
rect 111490 5800 111510 5860
rect 111570 5800 111580 5860
rect 116020 5860 116260 5880
rect 111340 5790 111580 5800
rect 111690 5830 115910 5840
rect 111690 5770 111700 5830
rect 111760 5770 112238 5830
rect 112292 5770 112348 5830
rect 112402 5770 112458 5830
rect 112512 5770 112568 5830
rect 112622 5770 112678 5830
rect 112732 5770 112788 5830
rect 112842 5770 112898 5830
rect 112952 5770 113008 5830
rect 113062 5770 113118 5830
rect 113172 5770 113228 5830
rect 113282 5770 114318 5830
rect 114372 5770 114428 5830
rect 114482 5770 114538 5830
rect 114592 5770 114648 5830
rect 114702 5770 114758 5830
rect 114812 5770 114868 5830
rect 114922 5770 114978 5830
rect 115032 5770 115088 5830
rect 115142 5770 115198 5830
rect 115252 5770 115308 5830
rect 115362 5770 115840 5830
rect 115900 5770 115910 5830
rect 116020 5800 116030 5860
rect 116090 5800 116110 5860
rect 116170 5800 116190 5860
rect 116250 5800 116260 5860
rect 116020 5790 116260 5800
rect 111690 5760 115910 5770
rect 109350 5720 109430 5730
rect 109350 5660 109360 5720
rect 109420 5710 109430 5720
rect 109570 5720 109650 5730
rect 109570 5710 109580 5720
rect 109420 5670 109580 5710
rect 109420 5660 109430 5670
rect 109350 5650 109430 5660
rect 109570 5660 109580 5670
rect 109640 5710 109650 5720
rect 109790 5720 109870 5730
rect 109790 5710 109800 5720
rect 109640 5670 109800 5710
rect 109640 5660 109650 5670
rect 109570 5650 109650 5660
rect 109790 5660 109800 5670
rect 109860 5710 109870 5720
rect 110010 5720 110090 5730
rect 110010 5710 110020 5720
rect 109860 5670 110020 5710
rect 109860 5660 109870 5670
rect 109790 5650 109870 5660
rect 110010 5660 110020 5670
rect 110080 5710 110090 5720
rect 110230 5720 110310 5730
rect 110230 5710 110240 5720
rect 110080 5670 110240 5710
rect 110080 5660 110090 5670
rect 110010 5650 110090 5660
rect 110230 5660 110240 5670
rect 110300 5710 110310 5720
rect 110450 5720 110530 5730
rect 110450 5710 110460 5720
rect 110300 5670 110460 5710
rect 110300 5660 110310 5670
rect 110230 5650 110310 5660
rect 110450 5660 110460 5670
rect 110520 5660 110530 5720
rect 110450 5650 110530 5660
rect 117070 5720 117150 5730
rect 117070 5660 117080 5720
rect 117140 5710 117150 5720
rect 117290 5720 117370 5730
rect 117290 5710 117300 5720
rect 117140 5670 117300 5710
rect 117140 5660 117150 5670
rect 117070 5650 117150 5660
rect 117290 5660 117300 5670
rect 117360 5710 117370 5720
rect 117510 5720 117590 5730
rect 117510 5710 117520 5720
rect 117360 5670 117520 5710
rect 117360 5660 117370 5670
rect 117290 5650 117370 5660
rect 117510 5660 117520 5670
rect 117580 5710 117590 5720
rect 117730 5720 117810 5730
rect 117730 5710 117740 5720
rect 117580 5670 117740 5710
rect 117580 5660 117590 5670
rect 117510 5650 117590 5660
rect 117730 5660 117740 5670
rect 117800 5710 117810 5720
rect 117950 5720 118030 5730
rect 117950 5710 117960 5720
rect 117800 5670 117960 5710
rect 117800 5660 117810 5670
rect 117730 5650 117810 5660
rect 117950 5660 117960 5670
rect 118020 5710 118030 5720
rect 118170 5720 118250 5730
rect 118170 5710 118180 5720
rect 118020 5670 118180 5710
rect 118020 5660 118030 5670
rect 117950 5650 118030 5660
rect 118170 5660 118180 5670
rect 118240 5660 118250 5720
rect 118170 5650 118250 5660
rect 108430 5560 111040 5570
rect 108430 5500 108440 5560
rect 108500 5500 108520 5560
rect 108580 5500 108600 5560
rect 108660 5500 109910 5560
rect 109970 5500 110810 5560
rect 110870 5500 110890 5560
rect 110950 5500 110970 5560
rect 111030 5500 111040 5560
rect 108430 5480 111040 5500
rect 108430 5420 108440 5480
rect 108500 5420 108520 5480
rect 108580 5420 108600 5480
rect 108660 5420 109910 5480
rect 109970 5420 110810 5480
rect 110870 5420 110890 5480
rect 110950 5420 110970 5480
rect 111030 5420 111040 5480
rect 116560 5560 119170 5570
rect 116560 5500 116570 5560
rect 116630 5500 116650 5560
rect 116710 5500 116730 5560
rect 116790 5500 117630 5560
rect 117690 5500 118940 5560
rect 119000 5500 119020 5560
rect 119080 5500 119100 5560
rect 119160 5500 119170 5560
rect 116560 5480 119170 5500
rect 108430 5400 111040 5420
rect 108430 5340 108440 5400
rect 108500 5340 108520 5400
rect 108580 5340 108600 5400
rect 108660 5340 109910 5400
rect 109970 5340 110810 5400
rect 110870 5340 110890 5400
rect 110950 5340 110970 5400
rect 111030 5340 111040 5400
rect 112280 5420 112360 5430
rect 112280 5360 112290 5420
rect 112350 5410 112360 5420
rect 112500 5420 112580 5430
rect 112500 5410 112510 5420
rect 112350 5370 112510 5410
rect 112350 5360 112360 5370
rect 112280 5350 112360 5360
rect 112500 5360 112510 5370
rect 112570 5410 112580 5420
rect 112720 5420 112800 5430
rect 112720 5410 112730 5420
rect 112570 5370 112730 5410
rect 112570 5360 112580 5370
rect 112500 5350 112580 5360
rect 112720 5360 112730 5370
rect 112790 5410 112800 5420
rect 112940 5420 113020 5430
rect 112940 5410 112950 5420
rect 112790 5370 112950 5410
rect 112790 5360 112800 5370
rect 112720 5350 112800 5360
rect 112940 5360 112950 5370
rect 113010 5410 113020 5420
rect 113160 5420 113240 5430
rect 113160 5410 113170 5420
rect 113010 5370 113170 5410
rect 113010 5360 113020 5370
rect 112940 5350 113020 5360
rect 113160 5360 113170 5370
rect 113230 5360 113240 5420
rect 113160 5350 113240 5360
rect 114360 5420 114440 5430
rect 114360 5360 114370 5420
rect 114430 5410 114440 5420
rect 114580 5420 114660 5430
rect 114580 5410 114590 5420
rect 114430 5370 114590 5410
rect 114430 5360 114440 5370
rect 114360 5350 114440 5360
rect 114580 5360 114590 5370
rect 114650 5410 114660 5420
rect 114800 5420 114880 5430
rect 114800 5410 114810 5420
rect 114650 5370 114810 5410
rect 114650 5360 114660 5370
rect 114580 5350 114660 5360
rect 114800 5360 114810 5370
rect 114870 5410 114880 5420
rect 115020 5420 115100 5430
rect 115020 5410 115030 5420
rect 114870 5370 115030 5410
rect 114870 5360 114880 5370
rect 114800 5350 114880 5360
rect 115020 5360 115030 5370
rect 115090 5410 115100 5420
rect 115240 5420 115320 5430
rect 115240 5410 115250 5420
rect 115090 5370 115250 5410
rect 115090 5360 115100 5370
rect 115020 5350 115100 5360
rect 115240 5360 115250 5370
rect 115310 5360 115320 5420
rect 115240 5350 115320 5360
rect 116560 5420 116570 5480
rect 116630 5420 116650 5480
rect 116710 5420 116730 5480
rect 116790 5420 117630 5480
rect 117690 5420 118940 5480
rect 119000 5420 119020 5480
rect 119080 5420 119100 5480
rect 119160 5420 119170 5480
rect 116560 5400 119170 5420
rect 108430 5330 111040 5340
rect 116560 5340 116570 5400
rect 116630 5340 116650 5400
rect 116710 5340 116730 5400
rect 116790 5340 117630 5400
rect 117690 5340 118940 5400
rect 119000 5340 119020 5400
rect 119080 5340 119100 5400
rect 119160 5340 119170 5400
rect 116560 5330 119170 5340
rect 112170 5310 113650 5320
rect 107980 5260 110530 5270
rect 107980 5200 107990 5260
rect 108050 5200 108070 5260
rect 108130 5200 108160 5260
rect 108220 5200 108240 5260
rect 108300 5200 108330 5260
rect 108390 5200 108410 5260
rect 108470 5200 109360 5260
rect 109420 5200 109470 5260
rect 109530 5200 109580 5260
rect 109640 5200 109690 5260
rect 109750 5200 109800 5260
rect 109860 5200 109910 5260
rect 109970 5200 110020 5260
rect 110080 5200 110130 5260
rect 110190 5200 110240 5260
rect 110300 5200 110350 5260
rect 110410 5200 110460 5260
rect 110520 5200 110530 5260
rect 112170 5250 112180 5310
rect 112240 5250 112400 5310
rect 112460 5250 112620 5310
rect 112680 5250 112840 5310
rect 112900 5250 113060 5310
rect 113120 5250 113280 5310
rect 113340 5250 113580 5310
rect 113640 5250 113650 5310
rect 112170 5240 113650 5250
rect 113950 5310 115430 5320
rect 113950 5250 113960 5310
rect 114020 5250 114260 5310
rect 114320 5250 114480 5310
rect 114540 5250 114700 5310
rect 114760 5250 114920 5310
rect 114980 5250 115140 5310
rect 115200 5250 115360 5310
rect 115420 5250 115430 5310
rect 113950 5240 115430 5250
rect 117070 5260 119620 5270
rect 107980 5180 110530 5200
rect 107980 5120 107990 5180
rect 108050 5120 108070 5180
rect 108130 5120 108160 5180
rect 108220 5120 108240 5180
rect 108300 5120 108330 5180
rect 108390 5120 108410 5180
rect 108470 5120 109360 5180
rect 109420 5120 109470 5180
rect 109530 5120 109580 5180
rect 109640 5120 109690 5180
rect 109750 5120 109800 5180
rect 109860 5120 109910 5180
rect 109970 5120 110020 5180
rect 110080 5120 110130 5180
rect 110190 5120 110240 5180
rect 110300 5120 110350 5180
rect 110410 5120 110460 5180
rect 110520 5120 110530 5180
rect 107980 5100 110530 5120
rect 107980 5040 107990 5100
rect 108050 5040 108070 5100
rect 108130 5040 108160 5100
rect 108220 5040 108240 5100
rect 108300 5040 108330 5100
rect 108390 5040 108410 5100
rect 108470 5040 109360 5100
rect 109420 5040 109470 5100
rect 109530 5040 109580 5100
rect 109640 5040 109690 5100
rect 109750 5040 109800 5100
rect 109860 5040 109910 5100
rect 109970 5040 110020 5100
rect 110080 5040 110130 5100
rect 110190 5040 110240 5100
rect 110300 5040 110350 5100
rect 110410 5040 110460 5100
rect 110520 5040 110530 5100
rect 107980 5030 110530 5040
rect 111340 5200 116260 5210
rect 111340 5140 111350 5200
rect 111410 5140 111430 5200
rect 111490 5140 111510 5200
rect 111570 5140 112070 5200
rect 112130 5140 113390 5200
rect 113450 5140 114150 5200
rect 114210 5140 115470 5200
rect 115530 5140 116030 5200
rect 116090 5140 116110 5200
rect 116170 5140 116190 5200
rect 116250 5140 116260 5200
rect 111340 5120 116260 5140
rect 111340 5060 111350 5120
rect 111410 5060 111430 5120
rect 111490 5060 111510 5120
rect 111570 5060 112070 5120
rect 112130 5060 113390 5120
rect 113450 5060 114150 5120
rect 114210 5060 115470 5120
rect 115530 5060 116030 5120
rect 116090 5060 116110 5120
rect 116170 5060 116190 5120
rect 116250 5060 116260 5120
rect 111340 5040 116260 5060
rect 109240 4990 111310 5000
rect 109240 4930 109250 4990
rect 109310 4930 110570 4990
rect 110630 4930 111080 4990
rect 111140 4930 111160 4990
rect 111220 4930 111240 4990
rect 111300 4930 111310 4990
rect 111340 4980 111350 5040
rect 111410 4980 111430 5040
rect 111490 4980 111510 5040
rect 111570 4980 112070 5040
rect 112130 4980 113390 5040
rect 113450 4980 114150 5040
rect 114210 4980 115470 5040
rect 115530 4980 116030 5040
rect 116090 4980 116110 5040
rect 116170 4980 116190 5040
rect 116250 4980 116260 5040
rect 117070 5200 117080 5260
rect 117140 5200 117190 5260
rect 117250 5200 117300 5260
rect 117360 5200 117410 5260
rect 117470 5200 117520 5260
rect 117580 5200 117630 5260
rect 117690 5200 117740 5260
rect 117800 5200 117850 5260
rect 117910 5200 117960 5260
rect 118020 5200 118070 5260
rect 118130 5200 118180 5260
rect 118240 5200 119130 5260
rect 119190 5200 119210 5260
rect 119270 5200 119300 5260
rect 119360 5200 119380 5260
rect 119440 5200 119470 5260
rect 119530 5200 119550 5260
rect 119610 5200 119620 5260
rect 117070 5180 119620 5200
rect 117070 5120 117080 5180
rect 117140 5120 117190 5180
rect 117250 5120 117300 5180
rect 117360 5120 117410 5180
rect 117470 5120 117520 5180
rect 117580 5120 117630 5180
rect 117690 5120 117740 5180
rect 117800 5120 117850 5180
rect 117910 5120 117960 5180
rect 118020 5120 118070 5180
rect 118130 5120 118180 5180
rect 118240 5120 119130 5180
rect 119190 5120 119210 5180
rect 119270 5120 119300 5180
rect 119360 5120 119380 5180
rect 119440 5120 119470 5180
rect 119530 5120 119550 5180
rect 119610 5120 119620 5180
rect 117070 5100 119620 5120
rect 117070 5040 117080 5100
rect 117140 5040 117190 5100
rect 117250 5040 117300 5100
rect 117360 5040 117410 5100
rect 117470 5040 117520 5100
rect 117580 5040 117630 5100
rect 117690 5040 117740 5100
rect 117800 5040 117850 5100
rect 117910 5040 117960 5100
rect 118020 5040 118070 5100
rect 118130 5040 118180 5100
rect 118240 5040 119130 5100
rect 119190 5040 119210 5100
rect 119270 5040 119300 5100
rect 119360 5040 119380 5100
rect 119440 5040 119470 5100
rect 119530 5040 119550 5100
rect 119610 5040 119620 5100
rect 117070 5030 119620 5040
rect 111340 4970 116260 4980
rect 116290 4990 118360 5000
rect 109240 4910 111310 4930
rect 109240 4850 109250 4910
rect 109310 4850 110570 4910
rect 110630 4850 111080 4910
rect 111140 4850 111160 4910
rect 111220 4850 111240 4910
rect 111300 4850 111310 4910
rect 109240 4830 111310 4850
rect 109240 4770 109250 4830
rect 109310 4770 110570 4830
rect 110630 4770 111080 4830
rect 111140 4770 111160 4830
rect 111220 4770 111240 4830
rect 111300 4770 111310 4830
rect 109240 4760 111310 4770
rect 116290 4930 116300 4990
rect 116360 4930 116380 4990
rect 116440 4930 116460 4990
rect 116520 4930 116970 4990
rect 117030 4930 118290 4990
rect 118350 4930 118360 4990
rect 116290 4910 118360 4930
rect 116290 4850 116300 4910
rect 116360 4850 116380 4910
rect 116440 4850 116460 4910
rect 116520 4850 116970 4910
rect 117030 4850 118290 4910
rect 118350 4850 118360 4910
rect 116290 4830 118360 4850
rect 116290 4770 116300 4830
rect 116360 4770 116380 4830
rect 116440 4770 116460 4830
rect 116520 4770 116970 4830
rect 117030 4770 118290 4830
rect 118350 4770 118360 4830
rect 116290 4760 118360 4770
rect 107680 4720 111580 4730
rect 107680 4660 107690 4720
rect 107750 4660 107770 4720
rect 107830 4660 107850 4720
rect 107910 4660 109360 4720
rect 109420 4660 109580 4720
rect 109640 4660 109800 4720
rect 109860 4660 110020 4720
rect 110080 4660 110240 4720
rect 110300 4660 110460 4720
rect 110520 4660 111350 4720
rect 111410 4660 111430 4720
rect 111490 4660 111510 4720
rect 111570 4660 111580 4720
rect 107680 4640 111580 4660
rect 107680 4580 107690 4640
rect 107750 4580 107770 4640
rect 107830 4580 107850 4640
rect 107910 4580 109360 4640
rect 109420 4580 109580 4640
rect 109640 4580 109800 4640
rect 109860 4580 110020 4640
rect 110080 4580 110240 4640
rect 110300 4580 110460 4640
rect 110520 4580 111350 4640
rect 111410 4580 111430 4640
rect 111490 4580 111510 4640
rect 111570 4580 111580 4640
rect 107680 4560 111580 4580
rect 107680 4500 107690 4560
rect 107750 4500 107770 4560
rect 107830 4500 107850 4560
rect 107910 4500 109360 4560
rect 109420 4500 109580 4560
rect 109640 4500 109800 4560
rect 109860 4500 110020 4560
rect 110080 4500 110240 4560
rect 110300 4500 110460 4560
rect 110520 4500 111350 4560
rect 111410 4500 111430 4560
rect 111490 4500 111510 4560
rect 111570 4500 111580 4560
rect 107680 4490 111580 4500
rect 116020 4720 119630 4730
rect 116020 4660 116030 4720
rect 116090 4660 116110 4720
rect 116170 4660 116190 4720
rect 116250 4660 117080 4720
rect 117140 4660 117300 4720
rect 117360 4660 117520 4720
rect 117580 4660 117740 4720
rect 117800 4660 117960 4720
rect 118020 4660 118180 4720
rect 118240 4710 119920 4720
rect 118240 4660 119690 4710
rect 116020 4650 119690 4660
rect 119750 4650 119770 4710
rect 119830 4650 119850 4710
rect 119910 4650 119920 4710
rect 116020 4640 119920 4650
rect 116020 4580 116030 4640
rect 116090 4580 116110 4640
rect 116170 4580 116190 4640
rect 116250 4580 117080 4640
rect 117140 4580 117300 4640
rect 117360 4580 117520 4640
rect 117580 4580 117740 4640
rect 117800 4580 117960 4640
rect 118020 4580 118180 4640
rect 118240 4630 119920 4640
rect 118240 4580 119690 4630
rect 116020 4570 119690 4580
rect 119750 4570 119770 4630
rect 119830 4570 119850 4630
rect 119910 4570 119920 4630
rect 116020 4560 119920 4570
rect 116020 4500 116030 4560
rect 116090 4500 116110 4560
rect 116170 4500 116190 4560
rect 116250 4500 117080 4560
rect 117140 4500 117300 4560
rect 117360 4500 117520 4560
rect 117580 4500 117740 4560
rect 117800 4500 117960 4560
rect 118020 4500 118180 4560
rect 118240 4550 119920 4560
rect 118240 4500 119690 4550
rect 116020 4490 119690 4500
rect 119750 4490 119770 4550
rect 119830 4490 119850 4550
rect 119910 4490 119920 4550
rect 119630 4480 119920 4490
rect 109460 4450 109540 4460
rect 109460 4390 109470 4450
rect 109530 4440 109540 4450
rect 109680 4450 109760 4460
rect 109680 4440 109690 4450
rect 109530 4400 109690 4440
rect 109530 4390 109540 4400
rect 109460 4380 109540 4390
rect 109680 4390 109690 4400
rect 109750 4440 109760 4450
rect 109900 4450 109980 4460
rect 109900 4440 109910 4450
rect 109750 4400 109910 4440
rect 109750 4390 109760 4400
rect 109680 4380 109760 4390
rect 109900 4390 109910 4400
rect 109970 4440 109980 4450
rect 110120 4450 110200 4460
rect 110120 4440 110130 4450
rect 109970 4400 110130 4440
rect 109970 4390 109980 4400
rect 109900 4380 109980 4390
rect 110120 4390 110130 4400
rect 110190 4440 110200 4450
rect 110340 4450 110420 4460
rect 110340 4440 110350 4450
rect 110190 4400 110350 4440
rect 110190 4390 110200 4400
rect 110120 4380 110200 4390
rect 110340 4390 110350 4400
rect 110410 4390 110420 4450
rect 117180 4450 117260 4460
rect 110340 4380 110420 4390
rect 111340 4390 116260 4400
rect 111340 4330 111350 4390
rect 111410 4330 111430 4390
rect 111490 4330 111510 4390
rect 111570 4330 113770 4390
rect 113830 4330 116030 4390
rect 116090 4330 116110 4390
rect 116170 4330 116190 4390
rect 116250 4330 116260 4390
rect 117180 4390 117190 4450
rect 117250 4440 117260 4450
rect 117400 4450 117480 4460
rect 117400 4440 117410 4450
rect 117250 4400 117410 4440
rect 117250 4390 117260 4400
rect 117180 4380 117260 4390
rect 117400 4390 117410 4400
rect 117470 4440 117480 4450
rect 117620 4450 117700 4460
rect 117620 4440 117630 4450
rect 117470 4400 117630 4440
rect 117470 4390 117480 4400
rect 117400 4380 117480 4390
rect 117620 4390 117630 4400
rect 117690 4440 117700 4450
rect 117840 4450 117920 4460
rect 117840 4440 117850 4450
rect 117690 4400 117850 4440
rect 117690 4390 117700 4400
rect 117620 4380 117700 4390
rect 117840 4390 117850 4400
rect 117910 4440 117920 4450
rect 118060 4450 118140 4460
rect 118060 4440 118070 4450
rect 117910 4400 118070 4440
rect 117910 4390 117920 4400
rect 117840 4380 117920 4390
rect 118060 4390 118070 4400
rect 118130 4390 118140 4450
rect 118060 4380 118140 4390
rect 111340 4310 116260 4330
rect 111340 4250 111350 4310
rect 111410 4250 111430 4310
rect 111490 4250 111510 4310
rect 111570 4250 113770 4310
rect 113830 4250 116030 4310
rect 116090 4250 116110 4310
rect 116170 4250 116190 4310
rect 116250 4250 116260 4310
rect 111340 4230 116260 4250
rect 111340 4170 111350 4230
rect 111410 4170 111430 4230
rect 111490 4170 111510 4230
rect 111570 4170 113770 4230
rect 113830 4170 116030 4230
rect 116090 4170 116110 4230
rect 116170 4170 116190 4230
rect 116250 4170 116260 4230
rect 111340 4160 116260 4170
rect 107980 4120 108480 4140
rect 107980 4060 108000 4120
rect 108060 4060 108100 4120
rect 108160 4060 108200 4120
rect 108260 4060 108300 4120
rect 108360 4060 108400 4120
rect 108460 4060 108480 4120
rect 119120 4120 119620 4140
rect 119120 4060 119140 4120
rect 119200 4060 119240 4120
rect 119300 4060 119340 4120
rect 119400 4060 119440 4120
rect 119500 4060 119540 4120
rect 119600 4060 119620 4120
rect 107980 4020 108480 4060
rect 112290 4050 112350 4060
rect 112170 4030 112250 4040
rect 107980 3960 108000 4020
rect 108060 3960 108100 4020
rect 108160 3960 108200 4020
rect 108260 3960 108300 4020
rect 108360 3960 108400 4020
rect 108460 3960 108480 4020
rect 112080 4010 112140 4020
rect 112060 3960 112080 4000
rect 107980 3920 108480 3960
rect 112170 3970 112180 4030
rect 112240 4020 112250 4030
rect 112240 3990 112290 4020
rect 112510 4050 112570 4060
rect 112390 4030 112470 4040
rect 112390 4020 112400 4030
rect 112350 3990 112400 4020
rect 112240 3980 112400 3990
rect 112240 3970 112250 3980
rect 112170 3960 112250 3970
rect 112390 3970 112400 3980
rect 112460 4020 112470 4030
rect 112460 3990 112510 4020
rect 112730 4050 112790 4060
rect 112610 4030 112690 4040
rect 112610 4020 112620 4030
rect 112570 3990 112620 4020
rect 112460 3980 112620 3990
rect 112460 3970 112470 3980
rect 112390 3960 112470 3970
rect 112610 3970 112620 3980
rect 112680 4020 112690 4030
rect 112680 3990 112730 4020
rect 112950 4050 113010 4060
rect 112830 4030 112910 4040
rect 112830 4020 112840 4030
rect 112790 3990 112840 4020
rect 112680 3980 112840 3990
rect 112680 3970 112690 3980
rect 112610 3960 112690 3970
rect 112830 3970 112840 3980
rect 112900 4020 112910 4030
rect 112900 3990 112950 4020
rect 113170 4050 113230 4060
rect 113050 4030 113130 4040
rect 113050 4020 113060 4030
rect 113010 3990 113060 4020
rect 112900 3980 113060 3990
rect 112900 3970 112910 3980
rect 112830 3960 112910 3970
rect 113050 3970 113060 3980
rect 113120 4020 113130 4030
rect 113120 3990 113170 4020
rect 114370 4050 114430 4060
rect 113270 4030 113350 4040
rect 113270 4020 113280 4030
rect 113230 3990 113280 4020
rect 113120 3980 113280 3990
rect 113120 3970 113130 3980
rect 113050 3960 113130 3970
rect 113270 3970 113280 3980
rect 113340 3970 113350 4030
rect 113270 3960 113350 3970
rect 113380 4030 113440 4040
rect 113680 4030 113740 4040
rect 113440 3980 113680 4020
rect 113380 3960 113440 3970
rect 113680 3960 113740 3970
rect 113860 4030 113920 4040
rect 114160 4030 114220 4040
rect 113920 3980 114160 4020
rect 113860 3960 113920 3970
rect 114160 3960 114220 3970
rect 114250 4030 114330 4040
rect 114250 3970 114260 4030
rect 114320 4020 114330 4030
rect 114320 3990 114370 4020
rect 114590 4050 114650 4060
rect 114470 4030 114550 4040
rect 114470 4020 114480 4030
rect 114430 3990 114480 4020
rect 114320 3980 114480 3990
rect 114320 3970 114330 3980
rect 114250 3960 114330 3970
rect 114470 3970 114480 3980
rect 114540 4020 114550 4030
rect 114540 3990 114590 4020
rect 114810 4050 114870 4060
rect 114690 4030 114770 4040
rect 114690 4020 114700 4030
rect 114650 3990 114700 4020
rect 114540 3980 114700 3990
rect 114540 3970 114550 3980
rect 114470 3960 114550 3970
rect 114690 3970 114700 3980
rect 114760 4020 114770 4030
rect 114760 3990 114810 4020
rect 115030 4050 115090 4060
rect 114910 4030 114990 4040
rect 114910 4020 114920 4030
rect 114870 3990 114920 4020
rect 114760 3980 114920 3990
rect 114760 3970 114770 3980
rect 114690 3960 114770 3970
rect 114910 3970 114920 3980
rect 114980 4020 114990 4030
rect 114980 3990 115030 4020
rect 115250 4050 115310 4060
rect 115130 4030 115210 4040
rect 115130 4020 115140 4030
rect 115090 3990 115140 4020
rect 114980 3980 115140 3990
rect 114980 3970 114990 3980
rect 114910 3960 114990 3970
rect 115130 3970 115140 3980
rect 115200 4020 115210 4030
rect 115200 3990 115250 4020
rect 115350 4030 115430 4040
rect 115350 4020 115360 4030
rect 115310 3990 115360 4020
rect 115200 3980 115360 3990
rect 115200 3970 115210 3980
rect 115130 3960 115210 3970
rect 115350 3970 115360 3980
rect 115420 3970 115430 4030
rect 119120 4020 119620 4060
rect 115350 3960 115430 3970
rect 115460 4010 115520 4020
rect 115520 3960 115540 4000
rect 119120 3960 119140 4020
rect 119200 3960 119240 4020
rect 119300 3960 119340 4020
rect 119400 3960 119440 4020
rect 119500 3960 119540 4020
rect 119600 3960 119620 4020
rect 107980 3860 108000 3920
rect 108060 3860 108100 3920
rect 108160 3860 108200 3920
rect 108260 3860 108300 3920
rect 108360 3860 108400 3920
rect 108460 3860 108480 3920
rect 108970 3940 109050 3950
rect 108970 3880 108980 3940
rect 109040 3930 109050 3940
rect 109460 3940 109540 3950
rect 109460 3930 109470 3940
rect 109040 3890 109470 3930
rect 109040 3880 109050 3890
rect 108970 3870 109050 3880
rect 109460 3880 109470 3890
rect 109530 3930 109540 3940
rect 109680 3940 109760 3950
rect 109680 3930 109690 3940
rect 109530 3890 109690 3930
rect 109530 3880 109540 3890
rect 109460 3870 109540 3880
rect 109680 3880 109690 3890
rect 109750 3930 109760 3940
rect 109900 3940 109980 3950
rect 109900 3930 109910 3940
rect 109750 3890 109910 3930
rect 109750 3880 109760 3890
rect 109680 3870 109760 3880
rect 109900 3880 109910 3890
rect 109970 3930 109980 3940
rect 110120 3940 110200 3950
rect 110120 3930 110130 3940
rect 109970 3890 110130 3930
rect 109970 3880 109980 3890
rect 109900 3870 109980 3880
rect 110120 3880 110130 3890
rect 110190 3930 110200 3940
rect 110340 3940 110420 3950
rect 112080 3940 112140 3950
rect 112280 3940 112360 3950
rect 110340 3930 110350 3940
rect 110190 3890 110350 3930
rect 110190 3880 110200 3890
rect 110120 3870 110200 3880
rect 110340 3880 110350 3890
rect 110410 3880 110420 3940
rect 110340 3870 110420 3880
rect 112280 3880 112290 3940
rect 112350 3930 112360 3940
rect 112500 3940 112580 3950
rect 112500 3930 112510 3940
rect 112350 3890 112510 3930
rect 112350 3880 112360 3890
rect 112280 3870 112360 3880
rect 112500 3880 112510 3890
rect 112570 3930 112580 3940
rect 112720 3940 112800 3950
rect 112720 3930 112730 3940
rect 112570 3890 112730 3930
rect 112570 3880 112580 3890
rect 112500 3870 112580 3880
rect 112720 3880 112730 3890
rect 112790 3930 112800 3940
rect 112940 3940 113020 3950
rect 112940 3930 112950 3940
rect 112790 3890 112950 3930
rect 112790 3880 112800 3890
rect 112720 3870 112800 3880
rect 112940 3880 112950 3890
rect 113010 3930 113020 3940
rect 113160 3940 113240 3950
rect 113160 3930 113170 3940
rect 113010 3890 113170 3930
rect 113010 3880 113020 3890
rect 112940 3870 113020 3880
rect 113160 3880 113170 3890
rect 113230 3930 113240 3940
rect 114360 3940 114440 3950
rect 114360 3930 114370 3940
rect 113230 3890 114370 3930
rect 113230 3880 113240 3890
rect 113160 3870 113240 3880
rect 114360 3880 114370 3890
rect 114430 3930 114440 3940
rect 114580 3940 114660 3950
rect 114580 3930 114590 3940
rect 114430 3890 114590 3930
rect 114430 3880 114440 3890
rect 114360 3870 114440 3880
rect 114580 3880 114590 3890
rect 114650 3930 114660 3940
rect 114800 3940 114880 3950
rect 114800 3930 114810 3940
rect 114650 3890 114810 3930
rect 114650 3880 114660 3890
rect 114580 3870 114660 3880
rect 114800 3880 114810 3890
rect 114870 3930 114880 3940
rect 115020 3940 115100 3950
rect 115020 3930 115030 3940
rect 114870 3890 115030 3930
rect 114870 3880 114880 3890
rect 114800 3870 114880 3880
rect 115020 3880 115030 3890
rect 115090 3930 115100 3940
rect 115240 3940 115320 3950
rect 115460 3940 115520 3950
rect 117180 3940 117260 3950
rect 115240 3930 115250 3940
rect 115090 3890 115250 3930
rect 115090 3880 115100 3890
rect 115020 3870 115100 3880
rect 115240 3880 115250 3890
rect 115310 3880 115320 3940
rect 115240 3870 115320 3880
rect 117180 3880 117190 3940
rect 117250 3930 117260 3940
rect 117400 3940 117480 3950
rect 117400 3930 117410 3940
rect 117250 3890 117410 3930
rect 117250 3880 117260 3890
rect 117180 3870 117260 3880
rect 117400 3880 117410 3890
rect 117470 3930 117480 3940
rect 117620 3940 117700 3950
rect 117620 3930 117630 3940
rect 117470 3890 117630 3930
rect 117470 3880 117480 3890
rect 117400 3870 117480 3880
rect 117620 3880 117630 3890
rect 117690 3930 117700 3940
rect 117840 3940 117920 3950
rect 117840 3930 117850 3940
rect 117690 3890 117850 3930
rect 117690 3880 117700 3890
rect 117620 3870 117700 3880
rect 117840 3880 117850 3890
rect 117910 3930 117920 3940
rect 118060 3940 118140 3950
rect 118060 3930 118070 3940
rect 117910 3890 118070 3930
rect 117910 3880 117920 3890
rect 117840 3870 117920 3880
rect 118060 3880 118070 3890
rect 118130 3930 118140 3940
rect 118550 3940 118630 3950
rect 118550 3930 118560 3940
rect 118130 3890 118560 3930
rect 118130 3880 118140 3890
rect 118060 3870 118140 3880
rect 118550 3880 118560 3890
rect 118620 3880 118630 3940
rect 118550 3870 118630 3880
rect 119120 3920 119620 3960
rect 107980 3840 108480 3860
rect 119120 3860 119140 3920
rect 119200 3860 119240 3920
rect 119300 3860 119340 3920
rect 119400 3860 119440 3920
rect 119500 3860 119540 3920
rect 119600 3860 119620 3920
rect 119120 3840 119620 3860
rect 110230 3810 111040 3820
rect 110230 3750 110240 3810
rect 110300 3750 110810 3810
rect 110870 3750 110890 3810
rect 110950 3750 110970 3810
rect 111030 3750 111040 3810
rect 110230 3730 111040 3750
rect 110230 3670 110240 3730
rect 110300 3670 110810 3730
rect 110870 3670 110890 3730
rect 110950 3670 110970 3730
rect 111030 3670 111040 3730
rect 110230 3660 111040 3670
rect 116560 3810 117370 3820
rect 116560 3750 116570 3810
rect 116630 3750 116650 3810
rect 116710 3750 116730 3810
rect 116790 3750 117300 3810
rect 117360 3750 117370 3810
rect 116560 3730 117370 3750
rect 116560 3670 116570 3730
rect 116630 3670 116650 3730
rect 116710 3670 116730 3730
rect 116790 3670 117300 3730
rect 117360 3670 117370 3730
rect 116560 3660 117370 3670
rect 109060 3570 109140 3580
rect 109060 3510 109070 3570
rect 109130 3560 109140 3570
rect 109460 3570 109540 3580
rect 109460 3560 109470 3570
rect 109130 3520 109470 3560
rect 109130 3510 109140 3520
rect 109060 3500 109140 3510
rect 109460 3510 109470 3520
rect 109530 3560 109540 3570
rect 109680 3570 109760 3580
rect 109680 3560 109690 3570
rect 109530 3520 109690 3560
rect 109530 3510 109540 3520
rect 109460 3500 109540 3510
rect 109680 3510 109690 3520
rect 109750 3560 109760 3570
rect 109900 3570 109980 3580
rect 109900 3560 109910 3570
rect 109750 3520 109910 3560
rect 109750 3510 109760 3520
rect 109680 3500 109760 3510
rect 109900 3510 109910 3520
rect 109970 3560 109980 3570
rect 110120 3570 110200 3580
rect 110120 3560 110130 3570
rect 109970 3520 110130 3560
rect 109970 3510 109980 3520
rect 109900 3500 109980 3510
rect 110120 3510 110130 3520
rect 110190 3560 110200 3570
rect 110340 3570 110420 3580
rect 110340 3560 110350 3570
rect 110190 3520 110350 3560
rect 110190 3510 110200 3520
rect 110120 3500 110200 3510
rect 110340 3510 110350 3520
rect 110410 3510 110420 3570
rect 117180 3570 117260 3580
rect 110340 3500 110420 3510
rect 112170 3550 112250 3560
rect 112170 3490 112180 3550
rect 112240 3540 112250 3550
rect 112390 3550 112470 3560
rect 112390 3540 112400 3550
rect 112240 3500 112400 3540
rect 112240 3490 112250 3500
rect 112170 3480 112250 3490
rect 112390 3490 112400 3500
rect 112460 3540 112470 3550
rect 112610 3550 112690 3560
rect 112610 3540 112620 3550
rect 112460 3500 112620 3540
rect 112460 3490 112470 3500
rect 112390 3480 112470 3490
rect 112610 3490 112620 3500
rect 112680 3540 112690 3550
rect 112830 3550 112910 3560
rect 112830 3540 112840 3550
rect 112680 3500 112840 3540
rect 112680 3490 112690 3500
rect 112610 3480 112690 3490
rect 112830 3490 112840 3500
rect 112900 3540 112910 3550
rect 113050 3550 113130 3560
rect 113050 3540 113060 3550
rect 112900 3500 113060 3540
rect 112900 3490 112910 3500
rect 112830 3480 112910 3490
rect 113050 3490 113060 3500
rect 113120 3540 113130 3550
rect 113270 3550 113350 3560
rect 113270 3540 113280 3550
rect 113120 3500 113280 3540
rect 113120 3490 113130 3500
rect 113050 3480 113130 3490
rect 113270 3490 113280 3500
rect 113340 3490 113350 3550
rect 113270 3480 113350 3490
rect 113650 3550 113730 3560
rect 113650 3490 113660 3550
rect 113720 3540 113730 3550
rect 113870 3550 113950 3560
rect 113870 3540 113880 3550
rect 113720 3500 113880 3540
rect 113720 3490 113730 3500
rect 113650 3480 113730 3490
rect 113870 3490 113880 3500
rect 113940 3490 113950 3550
rect 113870 3480 113950 3490
rect 114250 3550 114330 3560
rect 114250 3490 114260 3550
rect 114320 3540 114330 3550
rect 114470 3550 114550 3560
rect 114470 3540 114480 3550
rect 114320 3500 114480 3540
rect 114320 3490 114330 3500
rect 114250 3480 114330 3490
rect 114470 3490 114480 3500
rect 114540 3540 114550 3550
rect 114690 3550 114770 3560
rect 114690 3540 114700 3550
rect 114540 3500 114700 3540
rect 114540 3490 114550 3500
rect 114470 3480 114550 3490
rect 114690 3490 114700 3500
rect 114760 3540 114770 3550
rect 114910 3550 114990 3560
rect 114910 3540 114920 3550
rect 114760 3500 114920 3540
rect 114760 3490 114770 3500
rect 114690 3480 114770 3490
rect 114910 3490 114920 3500
rect 114980 3540 114990 3550
rect 115130 3550 115210 3560
rect 115130 3540 115140 3550
rect 114980 3500 115140 3540
rect 114980 3490 114990 3500
rect 114910 3480 114990 3490
rect 115130 3490 115140 3500
rect 115200 3540 115210 3550
rect 115350 3550 115430 3560
rect 115350 3540 115360 3550
rect 115200 3500 115360 3540
rect 115200 3490 115210 3500
rect 115130 3480 115210 3490
rect 115350 3490 115360 3500
rect 115420 3490 115430 3550
rect 117180 3510 117190 3570
rect 117250 3560 117260 3570
rect 117400 3570 117480 3580
rect 117400 3560 117410 3570
rect 117250 3520 117410 3560
rect 117250 3510 117260 3520
rect 117180 3500 117260 3510
rect 117400 3510 117410 3520
rect 117470 3560 117480 3570
rect 117620 3570 117700 3580
rect 117620 3560 117630 3570
rect 117470 3520 117630 3560
rect 117470 3510 117480 3520
rect 117400 3500 117480 3510
rect 117620 3510 117630 3520
rect 117690 3560 117700 3570
rect 117840 3570 117920 3580
rect 117840 3560 117850 3570
rect 117690 3520 117850 3560
rect 117690 3510 117700 3520
rect 117620 3500 117700 3510
rect 117840 3510 117850 3520
rect 117910 3560 117920 3570
rect 118060 3570 118140 3580
rect 118060 3560 118070 3570
rect 117910 3520 118070 3560
rect 117910 3510 117920 3520
rect 117840 3500 117920 3510
rect 118060 3510 118070 3520
rect 118130 3560 118140 3570
rect 118460 3570 118540 3580
rect 118460 3560 118470 3570
rect 118130 3520 118470 3560
rect 118130 3510 118140 3520
rect 118060 3500 118140 3510
rect 118460 3510 118470 3520
rect 118530 3510 118540 3570
rect 118460 3500 118540 3510
rect 115350 3480 115430 3490
rect 112280 3410 115320 3420
rect 112280 3350 112290 3410
rect 112350 3350 112510 3410
rect 112570 3350 112730 3410
rect 112790 3350 112950 3410
rect 113010 3350 113170 3410
rect 113230 3350 114370 3410
rect 114430 3350 114590 3410
rect 114650 3350 114810 3410
rect 114870 3350 115030 3410
rect 115090 3350 115250 3410
rect 115310 3350 115320 3410
rect 112280 3340 115320 3350
rect 110800 3050 111040 3060
rect 110800 2990 110810 3050
rect 110870 2990 110890 3050
rect 110950 2990 110970 3050
rect 111030 2990 111040 3050
rect 110800 2970 111040 2990
rect 108510 2950 108580 2952
rect 108510 2940 108700 2950
rect 108580 2870 108630 2940
rect 108510 2860 108700 2870
rect 108750 2940 108820 2950
rect 108750 2860 108820 2870
rect 108870 2940 108940 2950
rect 109060 2930 109140 2940
rect 109060 2920 109070 2930
rect 108940 2880 109070 2920
rect 108870 2860 108940 2870
rect 109060 2870 109070 2880
rect 109130 2870 109140 2930
rect 110800 2910 110810 2970
rect 110870 2910 110890 2970
rect 110950 2910 110970 2970
rect 111030 2910 111040 2970
rect 109060 2860 109140 2870
rect 109460 2890 109540 2900
rect 109460 2830 109470 2890
rect 109530 2880 109540 2890
rect 109680 2890 109760 2900
rect 109680 2880 109690 2890
rect 109530 2840 109690 2880
rect 109530 2830 109540 2840
rect 109460 2820 109540 2830
rect 109680 2830 109690 2840
rect 109750 2880 109760 2890
rect 109900 2890 109980 2900
rect 109900 2880 109910 2890
rect 109750 2840 109910 2880
rect 109750 2830 109760 2840
rect 109680 2820 109760 2830
rect 109900 2830 109910 2840
rect 109970 2880 109980 2890
rect 110120 2890 110200 2900
rect 110120 2880 110130 2890
rect 109970 2840 110130 2880
rect 109970 2830 109980 2840
rect 109900 2820 109980 2830
rect 110120 2830 110130 2840
rect 110190 2880 110200 2890
rect 110340 2890 110420 2900
rect 110340 2880 110350 2890
rect 110190 2840 110350 2880
rect 110190 2830 110200 2840
rect 110120 2820 110200 2830
rect 110340 2830 110350 2840
rect 110410 2830 110420 2890
rect 110340 2820 110420 2830
rect 110800 2890 111040 2910
rect 110800 2830 110810 2890
rect 110870 2830 110890 2890
rect 110950 2830 110970 2890
rect 111030 2830 111040 2890
rect 110800 2820 111040 2830
rect 116560 3050 116800 3060
rect 116560 2990 116570 3050
rect 116630 2990 116650 3050
rect 116710 2990 116730 3050
rect 116790 2990 116800 3050
rect 116560 2970 116800 2990
rect 116560 2910 116570 2970
rect 116630 2910 116650 2970
rect 116710 2910 116730 2970
rect 116790 2910 116800 2970
rect 119020 2950 119090 2952
rect 118660 2940 118730 2950
rect 116560 2890 116800 2910
rect 118460 2930 118540 2940
rect 116560 2830 116570 2890
rect 116630 2830 116650 2890
rect 116710 2830 116730 2890
rect 116790 2830 116800 2890
rect 116560 2820 116800 2830
rect 117180 2890 117260 2900
rect 117180 2830 117190 2890
rect 117250 2880 117260 2890
rect 117400 2890 117480 2900
rect 117400 2880 117410 2890
rect 117250 2840 117410 2880
rect 117250 2830 117260 2840
rect 117180 2820 117260 2830
rect 117400 2830 117410 2840
rect 117470 2880 117480 2890
rect 117620 2890 117700 2900
rect 117620 2880 117630 2890
rect 117470 2840 117630 2880
rect 117470 2830 117480 2840
rect 117400 2820 117480 2830
rect 117620 2830 117630 2840
rect 117690 2880 117700 2890
rect 117840 2890 117920 2900
rect 117840 2880 117850 2890
rect 117690 2840 117850 2880
rect 117690 2830 117700 2840
rect 117620 2820 117700 2830
rect 117840 2830 117850 2840
rect 117910 2880 117920 2890
rect 118060 2890 118140 2900
rect 118060 2880 118070 2890
rect 117910 2840 118070 2880
rect 117910 2830 117920 2840
rect 117840 2820 117920 2830
rect 118060 2830 118070 2840
rect 118130 2830 118140 2890
rect 118460 2870 118470 2930
rect 118530 2920 118540 2930
rect 118530 2880 118660 2920
rect 118530 2870 118540 2880
rect 118460 2860 118540 2870
rect 118660 2860 118730 2870
rect 118780 2940 118850 2950
rect 118780 2860 118850 2870
rect 118900 2940 119090 2950
rect 118970 2870 119020 2940
rect 118900 2860 119090 2870
rect 118060 2820 118140 2830
rect 108750 2790 108830 2800
rect 108750 2730 108760 2790
rect 108820 2770 108830 2790
rect 108970 2790 109050 2800
rect 118550 2790 118630 2800
rect 108970 2770 108980 2790
rect 108820 2740 108980 2770
rect 108820 2730 108830 2740
rect 108750 2720 108830 2730
rect 108970 2730 108980 2740
rect 109040 2730 109050 2790
rect 108970 2720 109050 2730
rect 109350 2780 111310 2790
rect 109350 2720 109360 2780
rect 109420 2720 109580 2780
rect 109640 2720 109800 2780
rect 109860 2720 110020 2780
rect 110080 2720 110240 2780
rect 110300 2720 110460 2780
rect 110520 2720 111080 2780
rect 111140 2720 111160 2780
rect 111220 2720 111240 2780
rect 111300 2720 111310 2780
rect 109350 2700 111310 2720
rect 109350 2640 109360 2700
rect 109420 2640 109580 2700
rect 109640 2640 109800 2700
rect 109860 2640 110020 2700
rect 110080 2640 110240 2700
rect 110300 2640 110460 2700
rect 110520 2640 111080 2700
rect 111140 2640 111160 2700
rect 111220 2640 111240 2700
rect 111300 2640 111310 2700
rect 109350 2620 111310 2640
rect 109350 2560 109360 2620
rect 109420 2560 109580 2620
rect 109640 2560 109800 2620
rect 109860 2560 110020 2620
rect 110080 2560 110240 2620
rect 110300 2560 110460 2620
rect 110520 2560 111080 2620
rect 111140 2560 111160 2620
rect 111220 2560 111240 2620
rect 111300 2560 111310 2620
rect 109350 2550 111310 2560
rect 116290 2780 118250 2790
rect 116290 2720 116300 2780
rect 116360 2720 116380 2780
rect 116440 2720 116460 2780
rect 116520 2720 117080 2780
rect 117140 2720 117300 2780
rect 117360 2720 117520 2780
rect 117580 2720 117740 2780
rect 117800 2720 117960 2780
rect 118020 2720 118180 2780
rect 118240 2720 118250 2780
rect 118550 2730 118560 2790
rect 118620 2780 118630 2790
rect 118770 2790 118850 2800
rect 118770 2780 118780 2790
rect 118620 2740 118780 2780
rect 118620 2730 118630 2740
rect 118550 2720 118630 2730
rect 118770 2730 118780 2740
rect 118840 2730 118850 2790
rect 118770 2720 118850 2730
rect 116290 2700 118250 2720
rect 116290 2640 116300 2700
rect 116360 2640 116380 2700
rect 116440 2640 116460 2700
rect 116520 2640 117080 2700
rect 117140 2640 117300 2700
rect 117360 2640 117520 2700
rect 117580 2640 117740 2700
rect 117800 2640 117960 2700
rect 118020 2640 118180 2700
rect 118240 2640 118250 2700
rect 116290 2620 118250 2640
rect 116290 2560 116300 2620
rect 116360 2560 116380 2620
rect 116440 2560 116460 2620
rect 116520 2560 117080 2620
rect 117140 2560 117300 2620
rect 117360 2560 117520 2620
rect 117580 2560 117740 2620
rect 117800 2560 117960 2620
rect 118020 2560 118180 2620
rect 118240 2560 118250 2620
rect 116290 2550 118250 2560
rect 107680 2500 119920 2510
rect 107680 2440 107690 2500
rect 107750 2440 107770 2500
rect 107830 2440 107850 2500
rect 107910 2440 109250 2500
rect 109310 2440 110570 2500
rect 110630 2440 112070 2500
rect 112130 2440 113470 2500
rect 113530 2440 114070 2500
rect 114130 2440 115470 2500
rect 115530 2440 116970 2500
rect 117030 2440 118290 2500
rect 118350 2440 119690 2500
rect 119750 2440 119770 2500
rect 119830 2440 119850 2500
rect 119910 2440 119920 2500
rect 107680 2420 119920 2440
rect 107680 2360 107690 2420
rect 107750 2360 107770 2420
rect 107830 2360 107850 2420
rect 107910 2360 109250 2420
rect 109310 2360 110570 2420
rect 110630 2360 112070 2420
rect 112130 2360 113470 2420
rect 113530 2360 114070 2420
rect 114130 2360 115470 2420
rect 115530 2360 116970 2420
rect 117030 2360 118290 2420
rect 118350 2360 119690 2420
rect 119750 2360 119770 2420
rect 119830 2360 119850 2420
rect 119910 2360 119920 2420
rect 107680 2340 119920 2360
rect 107680 2280 107690 2340
rect 107750 2280 107770 2340
rect 107830 2280 107850 2340
rect 107910 2280 109250 2340
rect 109310 2280 110570 2340
rect 110630 2280 112070 2340
rect 112130 2280 113470 2340
rect 113530 2280 114070 2340
rect 114130 2280 115470 2340
rect 115530 2280 116970 2340
rect 117030 2280 118290 2340
rect 118350 2280 119690 2340
rect 119750 2280 119770 2340
rect 119830 2280 119850 2340
rect 119910 2280 119920 2340
rect 107680 2270 119920 2280
rect 108510 2230 108590 2240
rect 108510 2170 108520 2230
rect 108580 2220 108590 2230
rect 111880 2230 111960 2240
rect 111880 2220 111890 2230
rect 108580 2180 111890 2220
rect 108580 2170 108590 2180
rect 108510 2160 108590 2170
rect 111880 2170 111890 2180
rect 111950 2170 111960 2230
rect 111880 2160 111960 2170
rect 115630 2230 115710 2240
rect 115630 2170 115640 2230
rect 115700 2220 115710 2230
rect 119010 2230 119090 2240
rect 119010 2220 119020 2230
rect 115700 2180 119020 2220
rect 115700 2170 115710 2180
rect 115630 2160 115710 2170
rect 119010 2170 119020 2180
rect 119080 2170 119090 2230
rect 119010 2160 119090 2170
rect 108640 1850 118960 1860
rect 108640 1790 108650 1850
rect 108710 1790 118890 1850
rect 118950 1790 118960 1850
rect 108640 1780 118960 1790
rect 107980 1740 110380 1750
rect 117220 1740 119620 1750
rect 107980 1680 107990 1740
rect 108050 1680 108070 1740
rect 108130 1680 108160 1740
rect 108220 1680 108240 1740
rect 108300 1680 108330 1740
rect 108390 1680 108410 1740
rect 108470 1680 108780 1740
rect 108840 1680 109510 1740
rect 109570 1680 109590 1740
rect 109650 1680 109670 1740
rect 109730 1680 109750 1740
rect 109810 1680 109830 1740
rect 109890 1680 109910 1740
rect 109970 1680 109990 1740
rect 110050 1680 110070 1740
rect 110130 1680 110150 1740
rect 110210 1680 110230 1740
rect 110290 1680 110310 1740
rect 110370 1680 110380 1740
rect 107980 1660 110380 1680
rect 112880 1730 114940 1740
rect 112880 1670 112890 1730
rect 112950 1670 113110 1730
rect 113170 1670 113330 1730
rect 113390 1670 113550 1730
rect 113610 1670 113770 1730
rect 113830 1670 113990 1730
rect 114050 1670 114210 1730
rect 114270 1670 114430 1730
rect 114490 1670 114650 1730
rect 114710 1670 114870 1730
rect 114930 1670 114940 1730
rect 112880 1660 114940 1670
rect 117220 1680 117230 1740
rect 117290 1680 117310 1740
rect 117370 1680 117390 1740
rect 117450 1680 117470 1740
rect 117530 1680 117550 1740
rect 117610 1680 117630 1740
rect 117690 1680 117710 1740
rect 117770 1680 117790 1740
rect 117850 1680 117870 1740
rect 117930 1680 117950 1740
rect 118010 1680 118030 1740
rect 118090 1680 118760 1740
rect 118820 1680 119130 1740
rect 119190 1680 119210 1740
rect 119270 1680 119300 1740
rect 119360 1680 119380 1740
rect 119440 1680 119470 1740
rect 119530 1680 119550 1740
rect 119610 1680 119620 1740
rect 117220 1660 119620 1680
rect 107980 1600 107990 1660
rect 108050 1600 108070 1660
rect 108130 1600 108160 1660
rect 108220 1600 108240 1660
rect 108300 1600 108330 1660
rect 108390 1600 108410 1660
rect 108470 1600 108780 1660
rect 108840 1600 109510 1660
rect 109570 1600 109590 1660
rect 109650 1600 109670 1660
rect 109730 1600 109750 1660
rect 109810 1600 109830 1660
rect 109890 1600 109910 1660
rect 109970 1600 109990 1660
rect 110050 1600 110070 1660
rect 110130 1600 110150 1660
rect 110210 1600 110230 1660
rect 110290 1600 110310 1660
rect 110370 1600 110380 1660
rect 107980 1580 110380 1600
rect 107980 1520 107990 1580
rect 108050 1520 108070 1580
rect 108130 1520 108160 1580
rect 108220 1520 108240 1580
rect 108300 1520 108330 1580
rect 108390 1520 108410 1580
rect 108470 1520 108780 1580
rect 108840 1520 109510 1580
rect 109570 1520 109590 1580
rect 109650 1520 109670 1580
rect 109730 1520 109750 1580
rect 109810 1520 109830 1580
rect 109890 1520 109910 1580
rect 109970 1520 109990 1580
rect 110050 1520 110070 1580
rect 110130 1520 110150 1580
rect 110210 1520 110230 1580
rect 110290 1520 110310 1580
rect 110370 1520 110380 1580
rect 107980 1510 110380 1520
rect 117220 1600 117230 1660
rect 117290 1600 117310 1660
rect 117370 1600 117390 1660
rect 117450 1600 117470 1660
rect 117530 1600 117550 1660
rect 117610 1600 117630 1660
rect 117690 1600 117710 1660
rect 117770 1600 117790 1660
rect 117850 1600 117870 1660
rect 117930 1600 117950 1660
rect 118010 1600 118030 1660
rect 118090 1600 118760 1660
rect 118820 1600 119130 1660
rect 119190 1600 119210 1660
rect 119270 1600 119300 1660
rect 119360 1600 119380 1660
rect 119440 1600 119470 1660
rect 119530 1600 119550 1660
rect 119610 1600 119620 1660
rect 117220 1580 119620 1600
rect 117220 1520 117230 1580
rect 117290 1520 117310 1580
rect 117370 1520 117390 1580
rect 117450 1520 117470 1580
rect 117530 1520 117550 1580
rect 117610 1520 117630 1580
rect 117690 1520 117710 1580
rect 117770 1520 117790 1580
rect 117850 1520 117870 1580
rect 117930 1520 117950 1580
rect 118010 1520 118030 1580
rect 118090 1520 118760 1580
rect 118820 1520 119130 1580
rect 119190 1520 119210 1580
rect 119270 1520 119300 1580
rect 119360 1520 119380 1580
rect 119440 1520 119470 1580
rect 119530 1520 119550 1580
rect 119610 1520 119620 1580
rect 117220 1510 119620 1520
rect 108640 1470 110280 1480
rect 108640 1410 108650 1470
rect 108710 1410 109610 1470
rect 109670 1410 109810 1470
rect 109870 1410 110010 1470
rect 110070 1410 110210 1470
rect 110270 1410 110280 1470
rect 108640 1400 110280 1410
rect 117320 1470 118960 1480
rect 117320 1410 117330 1470
rect 117390 1410 117530 1470
rect 117590 1410 117730 1470
rect 117790 1410 117930 1470
rect 117990 1410 118890 1470
rect 118950 1410 118960 1470
rect 117320 1400 118960 1410
rect 108650 1360 108720 1370
rect 108650 1280 108720 1290
rect 108770 1360 108840 1370
rect 108770 1280 108840 1290
rect 118760 1360 118830 1370
rect 118760 1280 118830 1290
rect 118880 1360 118950 1370
rect 118880 1280 118950 1290
rect 112440 1070 112520 1080
rect 112440 1010 112450 1070
rect 112510 1060 112520 1070
rect 112550 1070 112630 1080
rect 112550 1060 112560 1070
rect 112510 1020 112560 1060
rect 112510 1010 112520 1020
rect 112440 1000 112520 1010
rect 112550 1010 112560 1020
rect 112620 1060 112630 1070
rect 112770 1070 112850 1080
rect 112770 1060 112780 1070
rect 112620 1020 112780 1060
rect 112620 1010 112630 1020
rect 112550 1000 112630 1010
rect 112770 1010 112780 1020
rect 112840 1060 112850 1070
rect 112990 1070 113070 1080
rect 112990 1060 113000 1070
rect 112840 1020 113000 1060
rect 112840 1010 112850 1020
rect 112770 1000 112850 1010
rect 112990 1010 113000 1020
rect 113060 1060 113070 1070
rect 113210 1070 113290 1080
rect 113210 1060 113220 1070
rect 113060 1020 113220 1060
rect 113060 1010 113070 1020
rect 112990 1000 113070 1010
rect 113210 1010 113220 1020
rect 113280 1060 113290 1070
rect 113430 1070 113510 1080
rect 113430 1060 113440 1070
rect 113280 1020 113440 1060
rect 113280 1010 113290 1020
rect 113210 1000 113290 1010
rect 113430 1010 113440 1020
rect 113500 1060 113510 1070
rect 113650 1070 113730 1080
rect 113650 1060 113660 1070
rect 113500 1020 113660 1060
rect 113500 1010 113510 1020
rect 113430 1000 113510 1010
rect 113650 1010 113660 1020
rect 113720 1060 113730 1070
rect 113870 1070 113950 1080
rect 113870 1060 113880 1070
rect 113720 1020 113880 1060
rect 113720 1010 113730 1020
rect 113650 1000 113730 1010
rect 113870 1010 113880 1020
rect 113940 1060 113950 1070
rect 114090 1070 114170 1080
rect 114090 1060 114100 1070
rect 113940 1020 114100 1060
rect 113940 1010 113950 1020
rect 113870 1000 113950 1010
rect 114090 1010 114100 1020
rect 114160 1060 114170 1070
rect 114310 1070 114390 1080
rect 114310 1060 114320 1070
rect 114160 1020 114320 1060
rect 114160 1010 114170 1020
rect 114090 1000 114170 1010
rect 114310 1010 114320 1020
rect 114380 1060 114390 1070
rect 114530 1070 114610 1080
rect 114530 1060 114540 1070
rect 114380 1020 114540 1060
rect 114380 1010 114390 1020
rect 114310 1000 114390 1010
rect 114530 1010 114540 1020
rect 114600 1060 114610 1070
rect 114750 1070 114830 1080
rect 114750 1060 114760 1070
rect 114600 1020 114760 1060
rect 114600 1010 114610 1020
rect 114530 1000 114610 1010
rect 114750 1010 114760 1020
rect 114820 1060 114830 1070
rect 114970 1070 115050 1080
rect 114970 1060 114980 1070
rect 114820 1020 114980 1060
rect 114820 1010 114830 1020
rect 114750 1000 114830 1010
rect 114970 1010 114980 1020
rect 115040 1010 115050 1070
rect 114970 1000 115050 1010
rect 112880 960 115320 970
rect 112880 900 112890 960
rect 112950 900 113110 960
rect 113170 900 113330 960
rect 113390 900 113550 960
rect 113610 900 113770 960
rect 113830 900 113990 960
rect 114050 900 114210 960
rect 114270 900 114430 960
rect 114490 900 114650 960
rect 114710 900 114870 960
rect 114930 900 115090 960
rect 115150 900 115170 960
rect 115230 900 115250 960
rect 115310 900 115320 960
rect 112880 880 115320 900
rect 112880 820 112890 880
rect 112950 820 113110 880
rect 113170 820 113330 880
rect 113390 820 113550 880
rect 113610 820 113770 880
rect 113830 820 113990 880
rect 114050 820 114210 880
rect 114270 820 114430 880
rect 114490 820 114650 880
rect 114710 820 114870 880
rect 114930 820 115090 880
rect 115150 820 115170 880
rect 115230 820 115250 880
rect 115310 820 115320 880
rect 112880 800 115320 820
rect 112880 740 112890 800
rect 112950 740 113110 800
rect 113170 740 113330 800
rect 113390 740 113550 800
rect 113610 740 113770 800
rect 113830 740 113990 800
rect 114050 740 114210 800
rect 114270 740 114430 800
rect 114490 740 114650 800
rect 114710 740 114870 800
rect 114930 740 115090 800
rect 115150 740 115170 800
rect 115230 740 115250 800
rect 115310 740 115320 800
rect 112880 730 115320 740
rect 114830 690 114910 700
rect 114830 630 114840 690
rect 114900 680 114910 690
rect 115720 690 115800 700
rect 115720 680 115730 690
rect 114900 640 115730 680
rect 114900 630 114910 640
rect 114830 620 114910 630
rect 115720 630 115730 640
rect 115790 630 115800 690
rect 115720 620 115800 630
rect 111340 580 116260 590
rect 111340 520 111350 580
rect 111410 520 111430 580
rect 111490 520 111510 580
rect 111570 520 112670 580
rect 112730 520 116030 580
rect 116090 520 116110 580
rect 116170 520 116190 580
rect 116250 520 116260 580
rect 111340 500 116260 520
rect 111340 440 111350 500
rect 111410 440 111430 500
rect 111490 440 111510 500
rect 111570 440 112670 500
rect 112730 440 116030 500
rect 116090 440 116110 500
rect 116170 440 116190 500
rect 116250 440 116260 500
rect 111340 420 116260 440
rect 111340 360 111350 420
rect 111410 360 111430 420
rect 111490 360 111510 420
rect 111570 360 112670 420
rect 112730 360 116030 420
rect 116090 360 116110 420
rect 116170 360 116190 420
rect 116250 360 116260 420
rect 111340 350 116260 360
rect 113240 310 113950 320
rect 113240 250 113250 310
rect 113310 250 113660 310
rect 113720 250 113880 310
rect 113940 250 113950 310
rect 113240 240 113950 250
rect 111690 200 115910 210
rect 111690 140 111700 200
rect 111760 140 113550 200
rect 113610 140 113770 200
rect 113830 140 113990 200
rect 114050 140 115840 200
rect 115900 140 115910 200
rect 111690 130 115910 140
rect 109500 -30 110380 -20
rect 109500 -90 109510 -30
rect 109570 -90 109910 -30
rect 109970 -90 110310 -30
rect 110370 -90 110380 -30
rect 109500 -100 110380 -90
rect 117220 -30 118100 -20
rect 117220 -90 117230 -30
rect 117290 -90 117630 -30
rect 117690 -90 118030 -30
rect 118090 -90 118100 -30
rect 117220 -100 118100 -90
rect 112440 -240 113500 -230
rect 112440 -300 112450 -240
rect 112510 -300 113500 -240
rect 112440 -310 113500 -300
rect 113540 -240 114060 -230
rect 113540 -300 113550 -240
rect 113610 -300 113770 -240
rect 113830 -300 113990 -240
rect 114050 -300 114060 -240
rect 113540 -310 114060 -300
rect 114100 -240 115050 -230
rect 114160 -300 114980 -240
rect 115040 -300 115050 -240
rect 114100 -310 115050 -300
rect 113760 -320 113840 -310
rect 113760 -380 113770 -320
rect 113830 -380 113840 -320
rect 113760 -390 113840 -380
rect 113240 -460 113430 -450
rect 113240 -520 113250 -460
rect 113310 -520 113430 -460
rect 113240 -540 113430 -520
rect 113240 -600 113250 -540
rect 113310 -600 113430 -540
rect 113240 -620 113430 -600
rect 113240 -680 113250 -620
rect 113310 -680 113430 -620
rect 113240 -690 113430 -680
rect 113490 -690 113500 -450
rect 114100 -690 114110 -450
rect 114170 -460 115320 -450
rect 114170 -520 115090 -460
rect 115150 -520 115170 -460
rect 115230 -520 115250 -460
rect 115310 -520 115320 -460
rect 114170 -540 115320 -520
rect 114170 -600 115090 -540
rect 115150 -600 115170 -540
rect 115230 -600 115250 -540
rect 115310 -600 115320 -540
rect 114170 -620 115320 -600
rect 114170 -680 115090 -620
rect 115150 -680 115170 -620
rect 115230 -680 115250 -620
rect 115310 -680 115320 -620
rect 114170 -690 115320 -680
rect 104580 -1160 123020 -1150
rect 104580 -1220 104590 -1160
rect 104650 -1220 104670 -1160
rect 104730 -1220 104750 -1160
rect 104810 -1220 105290 -1160
rect 105350 -1220 105370 -1160
rect 105430 -1220 105450 -1160
rect 105510 -1220 105990 -1160
rect 106050 -1220 106070 -1160
rect 106130 -1220 106150 -1160
rect 106210 -1220 106690 -1160
rect 106750 -1220 106770 -1160
rect 106830 -1220 106850 -1160
rect 106910 -1220 107390 -1160
rect 107450 -1220 107470 -1160
rect 107530 -1220 107550 -1160
rect 107610 -1220 107690 -1160
rect 107750 -1220 107770 -1160
rect 107830 -1220 107850 -1160
rect 107910 -1220 108090 -1160
rect 108150 -1220 108170 -1160
rect 108230 -1220 108250 -1160
rect 108310 -1220 108790 -1160
rect 108850 -1220 108870 -1160
rect 108930 -1220 108950 -1160
rect 109010 -1220 109310 -1160
rect 109370 -1220 109490 -1160
rect 109550 -1220 109570 -1160
rect 109630 -1220 109650 -1160
rect 109710 -1220 110190 -1160
rect 110250 -1220 110270 -1160
rect 110330 -1220 110350 -1160
rect 110410 -1220 110510 -1160
rect 110570 -1220 110890 -1160
rect 110950 -1220 110970 -1160
rect 111030 -1220 111050 -1160
rect 111110 -1220 111590 -1160
rect 111650 -1220 111670 -1160
rect 111730 -1220 111750 -1160
rect 111810 -1220 112290 -1160
rect 112350 -1220 112370 -1160
rect 112430 -1220 112450 -1160
rect 112510 -1220 112990 -1160
rect 113050 -1220 113070 -1160
rect 113130 -1220 113150 -1160
rect 113210 -1220 113690 -1160
rect 113750 -1220 113770 -1160
rect 113830 -1220 113850 -1160
rect 113910 -1220 114390 -1160
rect 114450 -1220 114470 -1160
rect 114530 -1220 114550 -1160
rect 114610 -1220 114980 -1160
rect 115040 -1220 115090 -1160
rect 115150 -1220 115170 -1160
rect 115230 -1220 115250 -1160
rect 115310 -1220 115790 -1160
rect 115850 -1220 115870 -1160
rect 115930 -1220 115950 -1160
rect 116010 -1220 116490 -1160
rect 116550 -1220 116570 -1160
rect 116630 -1220 116650 -1160
rect 116710 -1220 117030 -1160
rect 117090 -1220 117190 -1160
rect 117250 -1220 117270 -1160
rect 117330 -1220 117350 -1160
rect 117410 -1220 117890 -1160
rect 117950 -1220 117970 -1160
rect 118030 -1220 118050 -1160
rect 118110 -1220 118230 -1160
rect 118290 -1220 118750 -1160
rect 118810 -1220 118830 -1160
rect 118890 -1220 118910 -1160
rect 118970 -1220 119290 -1160
rect 119350 -1220 119370 -1160
rect 119430 -1220 119450 -1160
rect 119510 -1220 119690 -1160
rect 119750 -1220 119770 -1160
rect 119830 -1220 119850 -1160
rect 119910 -1220 119990 -1160
rect 120050 -1220 120070 -1160
rect 120130 -1220 120150 -1160
rect 120210 -1220 120690 -1160
rect 120750 -1220 120770 -1160
rect 120830 -1220 120850 -1160
rect 120910 -1220 121390 -1160
rect 121450 -1220 121470 -1160
rect 121530 -1220 121550 -1160
rect 121610 -1220 122090 -1160
rect 122150 -1220 122170 -1160
rect 122230 -1220 122250 -1160
rect 122310 -1220 122790 -1160
rect 122850 -1220 122870 -1160
rect 122930 -1220 122950 -1160
rect 123010 -1220 123020 -1160
rect 104580 -1240 123020 -1220
rect 104580 -1300 104590 -1240
rect 104650 -1300 104670 -1240
rect 104730 -1300 104750 -1240
rect 104810 -1300 105290 -1240
rect 105350 -1300 105370 -1240
rect 105430 -1300 105450 -1240
rect 105510 -1300 105990 -1240
rect 106050 -1300 106070 -1240
rect 106130 -1300 106150 -1240
rect 106210 -1300 106690 -1240
rect 106750 -1300 106770 -1240
rect 106830 -1300 106850 -1240
rect 106910 -1300 107390 -1240
rect 107450 -1300 107470 -1240
rect 107530 -1300 107550 -1240
rect 107610 -1300 107690 -1240
rect 107750 -1300 107770 -1240
rect 107830 -1300 107850 -1240
rect 107910 -1300 108090 -1240
rect 108150 -1300 108170 -1240
rect 108230 -1300 108250 -1240
rect 108310 -1300 108790 -1240
rect 108850 -1300 108870 -1240
rect 108930 -1300 108950 -1240
rect 109010 -1300 109310 -1240
rect 109370 -1300 109490 -1240
rect 109550 -1300 109570 -1240
rect 109630 -1300 109650 -1240
rect 109710 -1300 110190 -1240
rect 110250 -1300 110270 -1240
rect 110330 -1300 110350 -1240
rect 110410 -1300 110510 -1240
rect 110570 -1300 110890 -1240
rect 110950 -1300 110970 -1240
rect 111030 -1300 111050 -1240
rect 111110 -1300 111590 -1240
rect 111650 -1300 111670 -1240
rect 111730 -1300 111750 -1240
rect 111810 -1300 112290 -1240
rect 112350 -1300 112370 -1240
rect 112430 -1300 112450 -1240
rect 112510 -1300 112990 -1240
rect 113050 -1300 113070 -1240
rect 113130 -1300 113150 -1240
rect 113210 -1300 113690 -1240
rect 113750 -1300 113770 -1240
rect 113830 -1300 113850 -1240
rect 113910 -1300 114390 -1240
rect 114450 -1300 114470 -1240
rect 114530 -1300 114550 -1240
rect 114610 -1300 114980 -1240
rect 115040 -1300 115090 -1240
rect 115150 -1300 115170 -1240
rect 115230 -1300 115250 -1240
rect 115310 -1300 115790 -1240
rect 115850 -1300 115870 -1240
rect 115930 -1300 115950 -1240
rect 116010 -1300 116490 -1240
rect 116550 -1300 116570 -1240
rect 116630 -1300 116650 -1240
rect 116710 -1300 117030 -1240
rect 117090 -1300 117190 -1240
rect 117250 -1300 117270 -1240
rect 117330 -1300 117350 -1240
rect 117410 -1300 117890 -1240
rect 117950 -1300 117970 -1240
rect 118030 -1300 118050 -1240
rect 118110 -1300 118230 -1240
rect 118290 -1300 118750 -1240
rect 118810 -1300 118830 -1240
rect 118890 -1300 118910 -1240
rect 118970 -1300 119290 -1240
rect 119350 -1300 119370 -1240
rect 119430 -1300 119450 -1240
rect 119510 -1300 119690 -1240
rect 119750 -1300 119770 -1240
rect 119830 -1300 119850 -1240
rect 119910 -1300 119990 -1240
rect 120050 -1300 120070 -1240
rect 120130 -1300 120150 -1240
rect 120210 -1300 120690 -1240
rect 120750 -1300 120770 -1240
rect 120830 -1300 120850 -1240
rect 120910 -1300 121390 -1240
rect 121450 -1300 121470 -1240
rect 121530 -1300 121550 -1240
rect 121610 -1300 122090 -1240
rect 122150 -1300 122170 -1240
rect 122230 -1300 122250 -1240
rect 122310 -1300 122790 -1240
rect 122850 -1300 122870 -1240
rect 122930 -1300 122950 -1240
rect 123010 -1300 123020 -1240
rect 104580 -1320 123020 -1300
rect 104580 -1380 104590 -1320
rect 104650 -1380 104670 -1320
rect 104730 -1380 104750 -1320
rect 104810 -1380 105290 -1320
rect 105350 -1380 105370 -1320
rect 105430 -1380 105450 -1320
rect 105510 -1380 105990 -1320
rect 106050 -1380 106070 -1320
rect 106130 -1380 106150 -1320
rect 106210 -1380 106690 -1320
rect 106750 -1380 106770 -1320
rect 106830 -1380 106850 -1320
rect 106910 -1380 107390 -1320
rect 107450 -1380 107470 -1320
rect 107530 -1380 107550 -1320
rect 107610 -1380 107690 -1320
rect 107750 -1380 107770 -1320
rect 107830 -1380 107850 -1320
rect 107910 -1380 108090 -1320
rect 108150 -1380 108170 -1320
rect 108230 -1380 108250 -1320
rect 108310 -1380 108790 -1320
rect 108850 -1380 108870 -1320
rect 108930 -1380 108950 -1320
rect 109010 -1380 109310 -1320
rect 109370 -1380 109490 -1320
rect 109550 -1380 109570 -1320
rect 109630 -1380 109650 -1320
rect 109710 -1380 110190 -1320
rect 110250 -1380 110270 -1320
rect 110330 -1380 110350 -1320
rect 110410 -1380 110510 -1320
rect 110570 -1380 110890 -1320
rect 110950 -1380 110970 -1320
rect 111030 -1380 111050 -1320
rect 111110 -1380 111590 -1320
rect 111650 -1380 111670 -1320
rect 111730 -1380 111750 -1320
rect 111810 -1380 112290 -1320
rect 112350 -1380 112370 -1320
rect 112430 -1380 112450 -1320
rect 112510 -1380 112990 -1320
rect 113050 -1380 113070 -1320
rect 113130 -1380 113150 -1320
rect 113210 -1380 113690 -1320
rect 113750 -1380 113770 -1320
rect 113830 -1380 113850 -1320
rect 113910 -1380 114390 -1320
rect 114450 -1380 114470 -1320
rect 114530 -1380 114550 -1320
rect 114610 -1380 114980 -1320
rect 115040 -1380 115090 -1320
rect 115150 -1380 115170 -1320
rect 115230 -1380 115250 -1320
rect 115310 -1380 115790 -1320
rect 115850 -1380 115870 -1320
rect 115930 -1380 115950 -1320
rect 116010 -1380 116490 -1320
rect 116550 -1380 116570 -1320
rect 116630 -1380 116650 -1320
rect 116710 -1380 117030 -1320
rect 117090 -1380 117190 -1320
rect 117250 -1380 117270 -1320
rect 117330 -1380 117350 -1320
rect 117410 -1380 117890 -1320
rect 117950 -1380 117970 -1320
rect 118030 -1380 118050 -1320
rect 118110 -1380 118230 -1320
rect 118290 -1380 118750 -1320
rect 118810 -1380 118830 -1320
rect 118890 -1380 118910 -1320
rect 118970 -1380 119290 -1320
rect 119350 -1380 119370 -1320
rect 119430 -1380 119450 -1320
rect 119510 -1380 119690 -1320
rect 119750 -1380 119770 -1320
rect 119830 -1380 119850 -1320
rect 119910 -1380 119990 -1320
rect 120050 -1380 120070 -1320
rect 120130 -1380 120150 -1320
rect 120210 -1380 120690 -1320
rect 120750 -1380 120770 -1320
rect 120830 -1380 120850 -1320
rect 120910 -1380 121390 -1320
rect 121450 -1380 121470 -1320
rect 121530 -1380 121550 -1320
rect 121610 -1380 122090 -1320
rect 122150 -1380 122170 -1320
rect 122230 -1380 122250 -1320
rect 122310 -1380 122790 -1320
rect 122850 -1380 122870 -1320
rect 122930 -1380 122950 -1320
rect 123010 -1380 123020 -1320
rect 104580 -1390 123020 -1380
<< via2 >>
rect 108520 7610 108580 7670
rect 119020 7610 119080 7670
rect 108000 4060 108060 4120
rect 108100 4060 108160 4120
rect 108200 4060 108260 4120
rect 108300 4060 108360 4120
rect 108400 4060 108460 4120
rect 119140 4060 119200 4120
rect 119240 4060 119300 4120
rect 119340 4060 119400 4120
rect 119440 4060 119500 4120
rect 119540 4060 119600 4120
rect 108000 3960 108060 4020
rect 108100 3960 108160 4020
rect 108200 3960 108260 4020
rect 108300 3960 108360 4020
rect 108400 3960 108460 4020
rect 119140 3960 119200 4020
rect 119240 3960 119300 4020
rect 119340 3960 119400 4020
rect 119440 3960 119500 4020
rect 119540 3960 119600 4020
rect 108000 3860 108060 3920
rect 108100 3860 108160 3920
rect 108200 3860 108260 3920
rect 108300 3860 108360 3920
rect 108400 3860 108460 3920
rect 119140 3860 119200 3920
rect 119240 3860 119300 3920
rect 119340 3860 119400 3920
rect 119440 3860 119500 3920
rect 119540 3860 119600 3920
<< metal3 >>
rect 105700 11210 105800 11300
rect 121800 11210 121900 11290
rect 104120 11040 104580 11210
rect 104820 11040 105280 11210
rect 105520 11040 105980 11210
rect 106220 11040 106680 11210
rect 106920 11040 107380 11210
rect 107620 11040 108080 11210
rect 108320 11040 108780 11210
rect 109020 11040 109480 11210
rect 109720 11040 110180 11210
rect 110420 11040 110880 11210
rect 111120 11040 111580 11210
rect 111820 11040 112280 11210
rect 112520 11040 112980 11210
rect 113220 11040 113680 11210
rect 104120 10940 113680 11040
rect 104120 10750 104580 10940
rect 104820 10750 105280 10940
rect 105520 10750 105980 10940
rect 106220 10750 106680 10940
rect 106920 10750 107380 10940
rect 107620 10750 108080 10940
rect 108320 10750 108780 10940
rect 109020 10750 109480 10940
rect 109720 10750 110180 10940
rect 110420 10750 110880 10940
rect 111120 10750 111580 10940
rect 111820 10750 112280 10940
rect 112520 10750 112980 10940
rect 113220 10750 113680 10940
rect 113920 11040 114380 11210
rect 114620 11040 115080 11210
rect 115320 11040 115780 11210
rect 116020 11040 116480 11210
rect 116720 11040 117180 11210
rect 117420 11040 117880 11210
rect 118120 11040 118580 11210
rect 118820 11040 119280 11210
rect 119520 11040 119980 11210
rect 120220 11040 120680 11210
rect 120920 11040 121380 11210
rect 121620 11040 122080 11210
rect 122320 11040 122780 11210
rect 123020 11040 123480 11210
rect 113920 10940 123480 11040
rect 113920 10750 114380 10940
rect 114620 10750 115080 10940
rect 115320 10750 115780 10940
rect 116020 10750 116480 10940
rect 116720 10750 117180 10940
rect 117420 10750 117880 10940
rect 118120 10750 118580 10940
rect 118820 10750 119280 10940
rect 119520 10750 119980 10940
rect 120220 10750 120680 10940
rect 120920 10750 121380 10940
rect 121620 10750 122080 10940
rect 122320 10750 122780 10940
rect 123020 10750 123480 10940
rect 105700 10510 105800 10750
rect 107800 10510 107900 10750
rect 108500 10510 108600 10750
rect 109200 10510 109300 10750
rect 109900 10510 110000 10750
rect 110600 10510 110700 10750
rect 111300 10510 111400 10750
rect 112000 10510 112100 10750
rect 112700 10510 112800 10750
rect 113400 10510 113500 10750
rect 114100 10510 114200 10750
rect 114800 10510 114900 10750
rect 115500 10510 115600 10750
rect 116200 10510 116300 10750
rect 116900 10510 117000 10750
rect 117600 10510 117700 10750
rect 118300 10510 118400 10750
rect 119000 10510 119100 10750
rect 119700 10510 119800 10750
rect 121800 10510 121900 10750
rect 104120 10340 104580 10510
rect 104820 10340 105280 10510
rect 105520 10340 105980 10510
rect 106220 10340 106680 10510
rect 106920 10340 107380 10510
rect 104120 10240 107380 10340
rect 104120 10050 104580 10240
rect 104820 10050 105280 10240
rect 105520 10050 105980 10240
rect 106220 10050 106680 10240
rect 106920 10050 107380 10240
rect 107620 10050 108080 10510
rect 108320 10050 108780 10510
rect 109020 10050 109480 10510
rect 109720 10050 110180 10510
rect 110420 10050 110880 10510
rect 111120 10050 111580 10510
rect 111820 10050 112280 10510
rect 112520 10050 112980 10510
rect 113220 10050 113680 10510
rect 113920 10050 114380 10510
rect 114620 10050 115080 10510
rect 115320 10050 115780 10510
rect 116020 10050 116480 10510
rect 116720 10050 117180 10510
rect 117420 10050 117880 10510
rect 118120 10050 118580 10510
rect 118820 10050 119280 10510
rect 119520 10050 119980 10510
rect 120220 10340 120680 10510
rect 120920 10340 121380 10510
rect 121620 10340 122080 10510
rect 122320 10340 122780 10510
rect 123020 10340 123480 10510
rect 120220 10240 123480 10340
rect 120220 10050 120680 10240
rect 120920 10050 121380 10240
rect 121620 10050 122080 10240
rect 122320 10050 122780 10240
rect 123020 10050 123480 10240
rect 105700 9810 105800 10050
rect 107800 9810 107900 10050
rect 108500 9810 108600 10050
rect 119000 9810 119100 10050
rect 119700 9810 119800 10050
rect 121800 9810 121900 10050
rect 104120 9640 104580 9810
rect 104820 9640 105280 9810
rect 105520 9640 105980 9810
rect 106220 9640 106680 9810
rect 106920 9640 107380 9810
rect 104120 9540 107380 9640
rect 104120 9350 104580 9540
rect 104820 9350 105280 9540
rect 105520 9350 105980 9540
rect 106220 9350 106680 9540
rect 106920 9350 107380 9540
rect 107620 9350 108080 9810
rect 108320 9350 108780 9810
rect 118820 9350 119280 9810
rect 119520 9350 119980 9810
rect 120220 9640 120680 9810
rect 120920 9640 121380 9810
rect 121620 9640 122080 9810
rect 122320 9640 122780 9810
rect 123020 9640 123480 9810
rect 120220 9540 123480 9640
rect 120220 9350 120680 9540
rect 120920 9350 121380 9540
rect 121620 9350 122080 9540
rect 122320 9350 122780 9540
rect 123020 9350 123480 9540
rect 105700 9110 105800 9350
rect 104120 8940 104580 9110
rect 104820 8940 105280 9110
rect 105520 8940 105980 9110
rect 106220 8940 106680 9110
rect 106920 8940 107380 9110
rect 104120 8840 107380 8940
rect 104120 8650 104580 8840
rect 104820 8650 105280 8840
rect 105520 8650 105980 8840
rect 106220 8650 106680 8840
rect 106920 8650 107380 8840
rect 105700 8410 105800 8650
rect 104120 8240 104580 8410
rect 104820 8240 105280 8410
rect 105520 8240 105980 8410
rect 106220 8240 106680 8410
rect 106920 8240 107380 8410
rect 104120 8140 107380 8240
rect 104120 7950 104580 8140
rect 104820 7950 105280 8140
rect 105520 7950 105980 8140
rect 106220 7950 106680 8140
rect 106920 7950 107380 8140
rect 105700 7710 105800 7950
rect 104120 7540 104580 7710
rect 104820 7540 105280 7710
rect 105520 7540 105980 7710
rect 106220 7540 106680 7710
rect 106920 7540 107380 7710
rect 108510 7670 108590 9350
rect 108510 7610 108520 7670
rect 108580 7610 108590 7670
rect 108510 7600 108590 7610
rect 119010 7670 119090 9350
rect 121800 9110 121900 9350
rect 120220 8940 120680 9110
rect 120920 8940 121380 9110
rect 121620 8940 122080 9110
rect 122320 8940 122780 9110
rect 123020 8940 123480 9110
rect 120220 8840 123480 8940
rect 120220 8650 120680 8840
rect 120920 8650 121380 8840
rect 121620 8650 122080 8840
rect 122320 8650 122780 8840
rect 123020 8650 123480 8840
rect 121800 8410 121900 8650
rect 120220 8240 120680 8410
rect 120920 8240 121380 8410
rect 121620 8240 122080 8410
rect 122320 8240 122780 8410
rect 123020 8240 123480 8410
rect 120220 8140 123480 8240
rect 120220 7950 120680 8140
rect 120920 7950 121380 8140
rect 121620 7950 122080 8140
rect 122320 7950 122780 8140
rect 123020 7950 123480 8140
rect 121800 7710 121900 7950
rect 119010 7610 119020 7670
rect 119080 7610 119090 7670
rect 119010 7600 119090 7610
rect 104120 7440 107380 7540
rect 104120 7250 104580 7440
rect 104820 7250 105280 7440
rect 105520 7250 105980 7440
rect 106220 7250 106680 7440
rect 106920 7250 107380 7440
rect 120220 7540 120680 7710
rect 120920 7540 121380 7710
rect 121620 7540 122080 7710
rect 122320 7540 122780 7710
rect 123020 7540 123480 7710
rect 120220 7440 123480 7540
rect 120220 7250 120680 7440
rect 120920 7250 121380 7440
rect 121620 7250 122080 7440
rect 122320 7250 122780 7440
rect 123020 7250 123480 7440
rect 105700 7010 105800 7250
rect 121800 7010 121900 7250
rect 104120 6840 104580 7010
rect 104820 6840 105280 7010
rect 105520 6840 105980 7010
rect 106220 6840 106680 7010
rect 106920 6840 107380 7010
rect 104120 6740 107380 6840
rect 104120 6550 104580 6740
rect 104820 6550 105280 6740
rect 105520 6550 105980 6740
rect 106220 6550 106680 6740
rect 106920 6550 107380 6740
rect 120220 6840 120680 7010
rect 120920 6840 121380 7010
rect 121620 6840 122080 7010
rect 122320 6840 122780 7010
rect 123020 6840 123480 7010
rect 120220 6740 123480 6840
rect 120220 6550 120680 6740
rect 120920 6550 121380 6740
rect 121620 6550 122080 6740
rect 122320 6550 122780 6740
rect 123020 6550 123480 6740
rect 105700 6310 105800 6550
rect 121800 6310 121900 6550
rect 104120 6140 104580 6310
rect 104820 6140 105280 6310
rect 105520 6140 105980 6310
rect 106220 6140 106680 6310
rect 106920 6140 107380 6310
rect 104120 6040 107380 6140
rect 104120 5850 104580 6040
rect 104820 5850 105280 6040
rect 105520 5850 105980 6040
rect 106220 5850 106680 6040
rect 106920 5850 107380 6040
rect 120220 6140 120680 6310
rect 120920 6140 121380 6310
rect 121620 6140 122080 6310
rect 122320 6140 122780 6310
rect 123020 6140 123480 6310
rect 120220 6040 123480 6140
rect 120220 5850 120680 6040
rect 120920 5850 121380 6040
rect 121620 5850 122080 6040
rect 122320 5850 122780 6040
rect 123020 5850 123480 6040
rect 105700 5610 105800 5850
rect 121800 5610 121900 5850
rect 104120 5440 104580 5610
rect 104820 5440 105280 5610
rect 105520 5440 105980 5610
rect 106220 5440 106680 5610
rect 106920 5440 107380 5610
rect 104120 5340 107380 5440
rect 104120 5150 104580 5340
rect 104820 5150 105280 5340
rect 105520 5150 105980 5340
rect 106220 5150 106680 5340
rect 106920 5150 107380 5340
rect 120220 5440 120680 5610
rect 120920 5440 121380 5610
rect 121620 5440 122080 5610
rect 122320 5440 122780 5610
rect 123020 5440 123480 5610
rect 120220 5340 123480 5440
rect 120220 5150 120680 5340
rect 120920 5150 121380 5340
rect 121620 5150 122080 5340
rect 122320 5150 122780 5340
rect 123020 5150 123480 5340
rect 105700 4910 105800 5150
rect 121800 4910 121900 5150
rect 104120 4740 104580 4910
rect 104820 4740 105280 4910
rect 105520 4740 105980 4910
rect 106220 4740 106680 4910
rect 106920 4740 107380 4910
rect 104120 4640 107380 4740
rect 104120 4450 104580 4640
rect 104820 4450 105280 4640
rect 105520 4450 105980 4640
rect 106220 4450 106680 4640
rect 106920 4450 107380 4640
rect 120220 4740 120680 4910
rect 120920 4740 121380 4910
rect 121620 4740 122080 4910
rect 122320 4740 122780 4910
rect 123020 4740 123480 4910
rect 120220 4640 123480 4740
rect 120220 4450 120680 4640
rect 120920 4450 121380 4640
rect 121620 4450 122080 4640
rect 122320 4450 122780 4640
rect 123020 4450 123480 4640
rect 105700 4210 105800 4450
rect 121800 4210 121900 4450
rect 104120 4040 104580 4210
rect 104820 4040 105280 4210
rect 105520 4040 105980 4210
rect 106220 4040 106680 4210
rect 106920 4040 107380 4210
rect 104120 3940 107380 4040
rect 104120 3750 104580 3940
rect 104820 3750 105280 3940
rect 105520 3750 105980 3940
rect 106220 3750 106680 3940
rect 106920 3750 107380 3940
rect 107980 4130 108480 4140
rect 107980 4050 107990 4130
rect 108070 4050 108090 4130
rect 108170 4050 108190 4130
rect 108270 4050 108290 4130
rect 108370 4050 108390 4130
rect 108470 4050 108480 4130
rect 107980 4030 108480 4050
rect 107980 3950 107990 4030
rect 108070 3950 108090 4030
rect 108170 3950 108190 4030
rect 108270 3950 108290 4030
rect 108370 3950 108390 4030
rect 108470 3950 108480 4030
rect 107980 3930 108480 3950
rect 107980 3850 107990 3930
rect 108070 3850 108090 3930
rect 108170 3850 108190 3930
rect 108270 3850 108290 3930
rect 108370 3850 108390 3930
rect 108470 3850 108480 3930
rect 107980 3840 108480 3850
rect 119120 4130 119620 4140
rect 119120 4050 119130 4130
rect 119210 4050 119230 4130
rect 119310 4050 119330 4130
rect 119410 4050 119430 4130
rect 119510 4050 119530 4130
rect 119610 4050 119620 4130
rect 119120 4030 119620 4050
rect 119120 3950 119130 4030
rect 119210 3950 119230 4030
rect 119310 3950 119330 4030
rect 119410 3950 119430 4030
rect 119510 3950 119530 4030
rect 119610 3950 119620 4030
rect 119120 3930 119620 3950
rect 119120 3850 119130 3930
rect 119210 3850 119230 3930
rect 119310 3850 119330 3930
rect 119410 3850 119430 3930
rect 119510 3850 119530 3930
rect 119610 3850 119620 3930
rect 119120 3840 119620 3850
rect 120220 4040 120680 4210
rect 120920 4040 121380 4210
rect 121620 4040 122080 4210
rect 122320 4040 122780 4210
rect 123020 4040 123480 4210
rect 120220 3940 123480 4040
rect 120220 3750 120680 3940
rect 120920 3750 121380 3940
rect 121620 3750 122080 3940
rect 122320 3750 122780 3940
rect 123020 3750 123480 3940
rect 105700 3510 105800 3750
rect 121800 3510 121900 3750
rect 104120 3340 104580 3510
rect 104820 3340 105280 3510
rect 105520 3340 105980 3510
rect 106220 3340 106680 3510
rect 106920 3340 107380 3510
rect 104120 3240 107380 3340
rect 104120 3050 104580 3240
rect 104820 3050 105280 3240
rect 105520 3050 105980 3240
rect 106220 3050 106680 3240
rect 106920 3050 107380 3240
rect 120220 3340 120680 3510
rect 120920 3340 121380 3510
rect 121620 3340 122080 3510
rect 122320 3340 122780 3510
rect 123020 3340 123480 3510
rect 120220 3240 123480 3340
rect 120220 3050 120680 3240
rect 120920 3050 121380 3240
rect 121620 3050 122080 3240
rect 122320 3050 122780 3240
rect 123020 3050 123480 3240
rect 105700 2810 105800 3050
rect 121800 2810 121900 3050
rect 104120 2640 104580 2810
rect 104820 2640 105280 2810
rect 105520 2640 105980 2810
rect 106220 2640 106680 2810
rect 106920 2640 107380 2810
rect 104120 2540 107380 2640
rect 104120 2350 104580 2540
rect 104820 2350 105280 2540
rect 105520 2350 105980 2540
rect 106220 2350 106680 2540
rect 106920 2350 107380 2540
rect 120220 2640 120680 2810
rect 120920 2640 121380 2810
rect 121620 2640 122080 2810
rect 122320 2640 122780 2810
rect 123020 2640 123480 2810
rect 120220 2540 123480 2640
rect 120220 2350 120680 2540
rect 120920 2350 121380 2540
rect 121620 2350 122080 2540
rect 122320 2350 122780 2540
rect 123020 2350 123480 2540
rect 105700 2110 105800 2350
rect 121800 2110 121900 2350
rect 104120 1940 104580 2110
rect 104820 1940 105280 2110
rect 105520 1940 105980 2110
rect 106220 1940 106680 2110
rect 106920 1940 107380 2110
rect 104120 1840 107380 1940
rect 104120 1650 104580 1840
rect 104820 1650 105280 1840
rect 105520 1650 105980 1840
rect 106220 1650 106680 1840
rect 106920 1650 107380 1840
rect 120220 1940 120680 2110
rect 120920 1940 121380 2110
rect 121620 1940 122080 2110
rect 122320 1940 122780 2110
rect 123020 1940 123480 2110
rect 120220 1840 123480 1940
rect 120220 1650 120680 1840
rect 120920 1650 121380 1840
rect 121620 1650 122080 1840
rect 122320 1650 122780 1840
rect 123020 1650 123480 1840
rect 105700 1410 105800 1650
rect 121800 1410 121900 1650
rect 104120 1240 104580 1410
rect 104820 1240 105280 1410
rect 105520 1240 105980 1410
rect 106220 1240 106680 1410
rect 106920 1240 107380 1410
rect 104120 1140 107380 1240
rect 104120 950 104580 1140
rect 104820 950 105280 1140
rect 105520 950 105980 1140
rect 106220 950 106680 1140
rect 106920 950 107380 1140
rect 120220 1240 120680 1410
rect 120920 1240 121380 1410
rect 121620 1240 122080 1410
rect 122320 1240 122780 1410
rect 123020 1240 123480 1410
rect 120220 1140 123480 1240
rect 120220 950 120680 1140
rect 120920 950 121380 1140
rect 121620 950 122080 1140
rect 122320 950 122780 1140
rect 123020 950 123480 1140
rect 105700 710 105800 950
rect 121800 710 121900 950
rect 104120 540 104580 710
rect 104820 540 105280 710
rect 105520 540 105980 710
rect 106220 540 106680 710
rect 106920 540 107380 710
rect 104120 440 107380 540
rect 104120 250 104580 440
rect 104820 250 105280 440
rect 105520 250 105980 440
rect 106220 250 106680 440
rect 106920 250 107380 440
rect 120220 540 120680 710
rect 120920 540 121380 710
rect 121620 540 122080 710
rect 122320 540 122780 710
rect 123020 540 123480 710
rect 120220 440 123480 540
rect 120220 250 120680 440
rect 120920 250 121380 440
rect 121620 250 122080 440
rect 122320 250 122780 440
rect 123020 250 123480 440
rect 105700 10 105800 250
rect 121800 10 121900 250
rect 104120 -160 104580 10
rect 104820 -160 105280 10
rect 105520 -160 105980 10
rect 106220 -160 106680 10
rect 106920 -160 107380 10
rect 104120 -260 107380 -160
rect 104120 -450 104580 -260
rect 104820 -450 105280 -260
rect 105520 -450 105980 -260
rect 106220 -450 106680 -260
rect 106920 -450 107380 -260
rect 120220 -160 120680 10
rect 120920 -160 121380 10
rect 121620 -160 122080 10
rect 122320 -160 122780 10
rect 123020 -160 123480 10
rect 120220 -260 123480 -160
rect 120220 -450 120680 -260
rect 120920 -450 121380 -260
rect 121620 -450 122080 -260
rect 122320 -450 122780 -260
rect 123020 -450 123480 -260
rect 105700 -690 105800 -450
rect 121800 -690 121900 -450
rect 104120 -860 104580 -690
rect 104820 -860 105280 -690
rect 105520 -860 105980 -690
rect 106220 -860 106680 -690
rect 106920 -860 107380 -690
rect 104120 -960 107380 -860
rect 104120 -1150 104580 -960
rect 104820 -1150 105280 -960
rect 105520 -1150 105980 -960
rect 106220 -1150 106680 -960
rect 106920 -1150 107380 -960
rect 120220 -860 120680 -690
rect 120920 -860 121380 -690
rect 121620 -860 122080 -690
rect 122320 -860 122780 -690
rect 123020 -860 123480 -690
rect 120220 -960 123480 -860
rect 120220 -1150 120680 -960
rect 120920 -1150 121380 -960
rect 121620 -1150 122080 -960
rect 122320 -1150 122780 -960
rect 123020 -1150 123480 -960
rect 105700 -1390 105800 -1150
rect 121800 -1390 121900 -1150
rect 104120 -1560 104580 -1390
rect 104820 -1560 105280 -1390
rect 105520 -1560 105980 -1390
rect 106220 -1560 106680 -1390
rect 106920 -1560 107380 -1390
rect 107620 -1560 108080 -1390
rect 108320 -1560 108780 -1390
rect 109020 -1560 109480 -1390
rect 109720 -1560 110180 -1390
rect 110420 -1560 110880 -1390
rect 111120 -1560 111580 -1390
rect 111820 -1560 112280 -1390
rect 112520 -1560 112980 -1390
rect 113220 -1560 113680 -1390
rect 104120 -1660 113680 -1560
rect 104120 -1850 104580 -1660
rect 104820 -1850 105280 -1660
rect 105520 -1850 105980 -1660
rect 106220 -1850 106680 -1660
rect 106920 -1850 107380 -1660
rect 107620 -1850 108080 -1660
rect 108320 -1850 108780 -1660
rect 109020 -1850 109480 -1660
rect 109720 -1850 110180 -1660
rect 110420 -1850 110880 -1660
rect 111120 -1850 111580 -1660
rect 111820 -1850 112280 -1660
rect 112520 -1850 112980 -1660
rect 113220 -1850 113680 -1660
rect 113920 -1560 114380 -1390
rect 114620 -1560 115080 -1390
rect 115320 -1560 115780 -1390
rect 116020 -1560 116480 -1390
rect 116720 -1560 117180 -1390
rect 117420 -1560 117880 -1390
rect 118120 -1560 118580 -1390
rect 118820 -1560 119280 -1390
rect 119520 -1560 119980 -1390
rect 120220 -1560 120680 -1390
rect 120920 -1560 121380 -1390
rect 121620 -1560 122080 -1390
rect 122320 -1560 122780 -1390
rect 123020 -1560 123480 -1390
rect 113920 -1660 123480 -1560
rect 113920 -1850 114380 -1660
rect 114620 -1850 115080 -1660
rect 115320 -1850 115780 -1660
rect 116020 -1850 116480 -1660
rect 116720 -1850 117180 -1660
rect 117420 -1850 117880 -1660
rect 118120 -1850 118580 -1660
rect 118820 -1850 119280 -1660
rect 119520 -1850 119980 -1660
rect 120220 -1850 120680 -1660
rect 120920 -1850 121380 -1660
rect 121620 -1850 122080 -1660
rect 122320 -1850 122780 -1660
rect 123020 -1850 123480 -1660
rect 105700 -2090 105800 -1850
rect 106400 -2090 106500 -1850
rect 107100 -2090 107200 -1850
rect 107800 -2090 107900 -1850
rect 108500 -2090 108600 -1850
rect 109200 -2090 109300 -1850
rect 109900 -2090 110000 -1850
rect 110600 -2090 110700 -1850
rect 111300 -2090 111400 -1850
rect 112000 -2090 112100 -1850
rect 112700 -2090 112800 -1850
rect 113400 -2090 113500 -1850
rect 114100 -2090 114200 -1850
rect 114800 -2090 114900 -1850
rect 115500 -2090 115600 -1850
rect 116200 -2090 116300 -1850
rect 116900 -2090 117000 -1850
rect 117600 -2090 117700 -1850
rect 118300 -2090 118400 -1850
rect 119000 -2090 119100 -1850
rect 119700 -2090 119800 -1850
rect 120400 -2090 120500 -1850
rect 121100 -2090 121200 -1850
rect 121800 -2090 121900 -1850
rect 104120 -2260 104580 -2090
rect 104820 -2260 105280 -2090
rect 105520 -2260 105980 -2090
rect 104120 -2360 105980 -2260
rect 104120 -2550 104580 -2360
rect 104820 -2550 105280 -2360
rect 105520 -2550 105980 -2360
rect 106220 -2550 106680 -2090
rect 106920 -2550 107380 -2090
rect 107620 -2550 108080 -2090
rect 108320 -2550 108780 -2090
rect 109020 -2550 109480 -2090
rect 109720 -2550 110180 -2090
rect 110420 -2550 110880 -2090
rect 111120 -2550 111580 -2090
rect 111820 -2550 112280 -2090
rect 112520 -2550 112980 -2090
rect 113220 -2550 113680 -2090
rect 113920 -2550 114380 -2090
rect 114620 -2550 115080 -2090
rect 115320 -2550 115780 -2090
rect 116020 -2550 116480 -2090
rect 116720 -2550 117180 -2090
rect 117420 -2550 117880 -2090
rect 118120 -2550 118580 -2090
rect 118820 -2550 119280 -2090
rect 119520 -2550 119980 -2090
rect 120220 -2550 120680 -2090
rect 120920 -2550 121380 -2090
rect 121620 -2260 122080 -2090
rect 122320 -2260 122780 -2090
rect 123020 -2260 123480 -2090
rect 121620 -2360 123480 -2260
rect 121620 -2550 122080 -2360
rect 122320 -2550 122780 -2360
rect 123020 -2550 123480 -2360
<< via3 >>
rect 107990 4120 108070 4130
rect 107990 4060 108000 4120
rect 108000 4060 108060 4120
rect 108060 4060 108070 4120
rect 107990 4050 108070 4060
rect 108090 4120 108170 4130
rect 108090 4060 108100 4120
rect 108100 4060 108160 4120
rect 108160 4060 108170 4120
rect 108090 4050 108170 4060
rect 108190 4120 108270 4130
rect 108190 4060 108200 4120
rect 108200 4060 108260 4120
rect 108260 4060 108270 4120
rect 108190 4050 108270 4060
rect 108290 4120 108370 4130
rect 108290 4060 108300 4120
rect 108300 4060 108360 4120
rect 108360 4060 108370 4120
rect 108290 4050 108370 4060
rect 108390 4120 108470 4130
rect 108390 4060 108400 4120
rect 108400 4060 108460 4120
rect 108460 4060 108470 4120
rect 108390 4050 108470 4060
rect 107990 4020 108070 4030
rect 107990 3960 108000 4020
rect 108000 3960 108060 4020
rect 108060 3960 108070 4020
rect 107990 3950 108070 3960
rect 108090 4020 108170 4030
rect 108090 3960 108100 4020
rect 108100 3960 108160 4020
rect 108160 3960 108170 4020
rect 108090 3950 108170 3960
rect 108190 4020 108270 4030
rect 108190 3960 108200 4020
rect 108200 3960 108260 4020
rect 108260 3960 108270 4020
rect 108190 3950 108270 3960
rect 108290 4020 108370 4030
rect 108290 3960 108300 4020
rect 108300 3960 108360 4020
rect 108360 3960 108370 4020
rect 108290 3950 108370 3960
rect 108390 4020 108470 4030
rect 108390 3960 108400 4020
rect 108400 3960 108460 4020
rect 108460 3960 108470 4020
rect 108390 3950 108470 3960
rect 107990 3920 108070 3930
rect 107990 3860 108000 3920
rect 108000 3860 108060 3920
rect 108060 3860 108070 3920
rect 107990 3850 108070 3860
rect 108090 3920 108170 3930
rect 108090 3860 108100 3920
rect 108100 3860 108160 3920
rect 108160 3860 108170 3920
rect 108090 3850 108170 3860
rect 108190 3920 108270 3930
rect 108190 3860 108200 3920
rect 108200 3860 108260 3920
rect 108260 3860 108270 3920
rect 108190 3850 108270 3860
rect 108290 3920 108370 3930
rect 108290 3860 108300 3920
rect 108300 3860 108360 3920
rect 108360 3860 108370 3920
rect 108290 3850 108370 3860
rect 108390 3920 108470 3930
rect 108390 3860 108400 3920
rect 108400 3860 108460 3920
rect 108460 3860 108470 3920
rect 108390 3850 108470 3860
rect 119130 4120 119210 4130
rect 119130 4060 119140 4120
rect 119140 4060 119200 4120
rect 119200 4060 119210 4120
rect 119130 4050 119210 4060
rect 119230 4120 119310 4130
rect 119230 4060 119240 4120
rect 119240 4060 119300 4120
rect 119300 4060 119310 4120
rect 119230 4050 119310 4060
rect 119330 4120 119410 4130
rect 119330 4060 119340 4120
rect 119340 4060 119400 4120
rect 119400 4060 119410 4120
rect 119330 4050 119410 4060
rect 119430 4120 119510 4130
rect 119430 4060 119440 4120
rect 119440 4060 119500 4120
rect 119500 4060 119510 4120
rect 119430 4050 119510 4060
rect 119530 4120 119610 4130
rect 119530 4060 119540 4120
rect 119540 4060 119600 4120
rect 119600 4060 119610 4120
rect 119530 4050 119610 4060
rect 119130 4020 119210 4030
rect 119130 3960 119140 4020
rect 119140 3960 119200 4020
rect 119200 3960 119210 4020
rect 119130 3950 119210 3960
rect 119230 4020 119310 4030
rect 119230 3960 119240 4020
rect 119240 3960 119300 4020
rect 119300 3960 119310 4020
rect 119230 3950 119310 3960
rect 119330 4020 119410 4030
rect 119330 3960 119340 4020
rect 119340 3960 119400 4020
rect 119400 3960 119410 4020
rect 119330 3950 119410 3960
rect 119430 4020 119510 4030
rect 119430 3960 119440 4020
rect 119440 3960 119500 4020
rect 119500 3960 119510 4020
rect 119430 3950 119510 3960
rect 119530 4020 119610 4030
rect 119530 3960 119540 4020
rect 119540 3960 119600 4020
rect 119600 3960 119610 4020
rect 119530 3950 119610 3960
rect 119130 3920 119210 3930
rect 119130 3860 119140 3920
rect 119140 3860 119200 3920
rect 119200 3860 119210 3920
rect 119130 3850 119210 3860
rect 119230 3920 119310 3930
rect 119230 3860 119240 3920
rect 119240 3860 119300 3920
rect 119300 3860 119310 3920
rect 119230 3850 119310 3860
rect 119330 3920 119410 3930
rect 119330 3860 119340 3920
rect 119340 3860 119400 3920
rect 119400 3860 119410 3920
rect 119330 3850 119410 3860
rect 119430 3920 119510 3930
rect 119430 3860 119440 3920
rect 119440 3860 119500 3920
rect 119500 3860 119510 3920
rect 119430 3850 119510 3860
rect 119530 3920 119610 3930
rect 119530 3860 119540 3920
rect 119540 3860 119600 3920
rect 119600 3860 119610 3920
rect 119530 3850 119610 3860
<< mimcap >>
rect 104150 11030 104550 11180
rect 104150 10950 104310 11030
rect 104390 10950 104550 11030
rect 104150 10780 104550 10950
rect 104850 11030 105250 11180
rect 104850 10950 105010 11030
rect 105090 10950 105250 11030
rect 104850 10780 105250 10950
rect 105550 11030 105950 11180
rect 105550 10950 105710 11030
rect 105790 10950 105950 11030
rect 105550 10780 105950 10950
rect 106250 11030 106650 11180
rect 106250 10950 106410 11030
rect 106490 10950 106650 11030
rect 106250 10780 106650 10950
rect 106950 11030 107350 11180
rect 106950 10950 107110 11030
rect 107190 10950 107350 11030
rect 106950 10780 107350 10950
rect 107650 11030 108050 11180
rect 107650 10950 107810 11030
rect 107890 10950 108050 11030
rect 107650 10780 108050 10950
rect 108350 11030 108750 11180
rect 108350 10950 108510 11030
rect 108590 10950 108750 11030
rect 108350 10780 108750 10950
rect 109050 11030 109450 11180
rect 109050 10950 109210 11030
rect 109290 10950 109450 11030
rect 109050 10780 109450 10950
rect 109750 11030 110150 11180
rect 109750 10950 109910 11030
rect 109990 10950 110150 11030
rect 109750 10780 110150 10950
rect 110450 11030 110850 11180
rect 110450 10950 110610 11030
rect 110690 10950 110850 11030
rect 110450 10780 110850 10950
rect 111150 11030 111550 11180
rect 111150 10950 111310 11030
rect 111390 10950 111550 11030
rect 111150 10780 111550 10950
rect 111850 11030 112250 11180
rect 111850 10950 112010 11030
rect 112090 10950 112250 11030
rect 111850 10780 112250 10950
rect 112550 11030 112950 11180
rect 112550 10950 112710 11030
rect 112790 10950 112950 11030
rect 112550 10780 112950 10950
rect 113250 11030 113650 11180
rect 113250 10950 113410 11030
rect 113490 10950 113650 11030
rect 113250 10780 113650 10950
rect 113950 11030 114350 11180
rect 113950 10950 114110 11030
rect 114190 10950 114350 11030
rect 113950 10780 114350 10950
rect 114650 11030 115050 11180
rect 114650 10950 114810 11030
rect 114890 10950 115050 11030
rect 114650 10780 115050 10950
rect 115350 11030 115750 11180
rect 115350 10950 115510 11030
rect 115590 10950 115750 11030
rect 115350 10780 115750 10950
rect 116050 11030 116450 11180
rect 116050 10950 116210 11030
rect 116290 10950 116450 11030
rect 116050 10780 116450 10950
rect 116750 11030 117150 11180
rect 116750 10950 116910 11030
rect 116990 10950 117150 11030
rect 116750 10780 117150 10950
rect 117450 11030 117850 11180
rect 117450 10950 117610 11030
rect 117690 10950 117850 11030
rect 117450 10780 117850 10950
rect 118150 11030 118550 11180
rect 118150 10950 118310 11030
rect 118390 10950 118550 11030
rect 118150 10780 118550 10950
rect 118850 11030 119250 11180
rect 118850 10950 119010 11030
rect 119090 10950 119250 11030
rect 118850 10780 119250 10950
rect 119550 11030 119950 11180
rect 119550 10950 119710 11030
rect 119790 10950 119950 11030
rect 119550 10780 119950 10950
rect 120250 11030 120650 11180
rect 120250 10950 120410 11030
rect 120490 10950 120650 11030
rect 120250 10780 120650 10950
rect 120950 11030 121350 11180
rect 120950 10950 121110 11030
rect 121190 10950 121350 11030
rect 120950 10780 121350 10950
rect 121650 11030 122050 11180
rect 121650 10950 121810 11030
rect 121890 10950 122050 11030
rect 121650 10780 122050 10950
rect 122350 11030 122750 11180
rect 122350 10950 122510 11030
rect 122590 10950 122750 11030
rect 122350 10780 122750 10950
rect 123050 11030 123450 11180
rect 123050 10950 123210 11030
rect 123290 10950 123450 11030
rect 123050 10780 123450 10950
rect 104150 10330 104550 10480
rect 104150 10250 104310 10330
rect 104390 10250 104550 10330
rect 104150 10080 104550 10250
rect 104850 10330 105250 10480
rect 104850 10250 105010 10330
rect 105090 10250 105250 10330
rect 104850 10080 105250 10250
rect 105550 10330 105950 10480
rect 105550 10250 105710 10330
rect 105790 10250 105950 10330
rect 105550 10080 105950 10250
rect 106250 10330 106650 10480
rect 106250 10250 106410 10330
rect 106490 10250 106650 10330
rect 106250 10080 106650 10250
rect 106950 10330 107350 10480
rect 106950 10250 107110 10330
rect 107190 10250 107350 10330
rect 106950 10080 107350 10250
rect 107650 10330 108050 10480
rect 107650 10250 107810 10330
rect 107890 10250 108050 10330
rect 107650 10080 108050 10250
rect 108350 10330 108750 10480
rect 108350 10250 108510 10330
rect 108590 10250 108750 10330
rect 108350 10080 108750 10250
rect 109050 10330 109450 10480
rect 109050 10250 109210 10330
rect 109290 10250 109450 10330
rect 109050 10080 109450 10250
rect 109750 10330 110150 10480
rect 109750 10250 109910 10330
rect 109990 10250 110150 10330
rect 109750 10080 110150 10250
rect 110450 10310 110850 10480
rect 110450 10230 110610 10310
rect 110690 10230 110850 10310
rect 110450 10080 110850 10230
rect 111150 10310 111550 10480
rect 111150 10230 111310 10310
rect 111390 10230 111550 10310
rect 111150 10080 111550 10230
rect 111850 10330 112250 10480
rect 111850 10250 112010 10330
rect 112090 10250 112250 10330
rect 111850 10080 112250 10250
rect 112550 10310 112950 10480
rect 112550 10230 112710 10310
rect 112790 10230 112950 10310
rect 112550 10080 112950 10230
rect 113250 10310 113650 10480
rect 113250 10230 113410 10310
rect 113490 10230 113650 10310
rect 113250 10080 113650 10230
rect 113950 10310 114350 10480
rect 113950 10230 114110 10310
rect 114190 10230 114350 10310
rect 113950 10080 114350 10230
rect 114650 10310 115050 10480
rect 114650 10240 114810 10310
rect 114890 10240 115050 10310
rect 114650 10080 115050 10240
rect 115350 10330 115750 10480
rect 115350 10250 115510 10330
rect 115590 10250 115750 10330
rect 115350 10080 115750 10250
rect 116050 10310 116450 10480
rect 116050 10230 116210 10310
rect 116290 10230 116450 10310
rect 116050 10080 116450 10230
rect 116750 10310 117150 10480
rect 116750 10240 116910 10310
rect 116990 10240 117150 10310
rect 116750 10080 117150 10240
rect 117450 10330 117850 10480
rect 117450 10250 117610 10330
rect 117690 10250 117850 10330
rect 117450 10080 117850 10250
rect 118150 10330 118550 10480
rect 118150 10250 118310 10330
rect 118390 10250 118550 10330
rect 118150 10080 118550 10250
rect 118850 10330 119250 10480
rect 118850 10250 119010 10330
rect 119090 10250 119250 10330
rect 118850 10080 119250 10250
rect 119550 10330 119950 10480
rect 119550 10250 119710 10330
rect 119790 10250 119950 10330
rect 119550 10080 119950 10250
rect 120250 10330 120650 10480
rect 120250 10250 120410 10330
rect 120490 10250 120650 10330
rect 120250 10080 120650 10250
rect 120950 10330 121350 10480
rect 120950 10250 121110 10330
rect 121190 10250 121350 10330
rect 120950 10080 121350 10250
rect 121650 10330 122050 10480
rect 121650 10250 121810 10330
rect 121890 10250 122050 10330
rect 121650 10080 122050 10250
rect 122350 10330 122750 10480
rect 122350 10250 122510 10330
rect 122590 10250 122750 10330
rect 122350 10080 122750 10250
rect 123050 10330 123450 10480
rect 123050 10250 123210 10330
rect 123290 10250 123450 10330
rect 123050 10080 123450 10250
rect 104150 9630 104550 9780
rect 104150 9550 104310 9630
rect 104390 9550 104550 9630
rect 104150 9380 104550 9550
rect 104850 9630 105250 9780
rect 104850 9550 105010 9630
rect 105090 9550 105250 9630
rect 104850 9380 105250 9550
rect 105550 9630 105950 9780
rect 105550 9550 105710 9630
rect 105790 9550 105950 9630
rect 105550 9380 105950 9550
rect 106250 9630 106650 9780
rect 106250 9550 106410 9630
rect 106490 9550 106650 9630
rect 106250 9380 106650 9550
rect 106950 9630 107350 9780
rect 106950 9550 107110 9630
rect 107190 9550 107350 9630
rect 106950 9380 107350 9550
rect 107650 9630 108050 9780
rect 107650 9550 107810 9630
rect 107890 9550 108050 9630
rect 107650 9380 108050 9550
rect 108350 9630 108750 9780
rect 108350 9550 108510 9630
rect 108590 9550 108750 9630
rect 108350 9380 108750 9550
rect 118850 9630 119250 9780
rect 118850 9550 119010 9630
rect 119090 9550 119250 9630
rect 118850 9380 119250 9550
rect 119550 9630 119950 9780
rect 119550 9550 119710 9630
rect 119790 9550 119950 9630
rect 119550 9380 119950 9550
rect 120250 9630 120650 9780
rect 120250 9550 120410 9630
rect 120490 9550 120650 9630
rect 120250 9380 120650 9550
rect 120950 9630 121350 9780
rect 120950 9550 121110 9630
rect 121190 9550 121350 9630
rect 120950 9380 121350 9550
rect 121650 9630 122050 9780
rect 121650 9550 121810 9630
rect 121890 9550 122050 9630
rect 121650 9380 122050 9550
rect 122350 9630 122750 9780
rect 122350 9550 122510 9630
rect 122590 9550 122750 9630
rect 122350 9380 122750 9550
rect 123050 9630 123450 9780
rect 123050 9550 123210 9630
rect 123290 9550 123450 9630
rect 123050 9380 123450 9550
rect 104150 8930 104550 9080
rect 104150 8850 104310 8930
rect 104390 8850 104550 8930
rect 104150 8680 104550 8850
rect 104850 8930 105250 9080
rect 104850 8850 105010 8930
rect 105090 8850 105250 8930
rect 104850 8680 105250 8850
rect 105550 8930 105950 9080
rect 105550 8850 105710 8930
rect 105790 8850 105950 8930
rect 105550 8680 105950 8850
rect 106250 8930 106650 9080
rect 106250 8850 106410 8930
rect 106490 8850 106650 8930
rect 106250 8680 106650 8850
rect 106950 8930 107350 9080
rect 106950 8850 107110 8930
rect 107190 8850 107350 8930
rect 106950 8680 107350 8850
rect 120250 8930 120650 9080
rect 120250 8850 120410 8930
rect 120490 8850 120650 8930
rect 120250 8680 120650 8850
rect 120950 8930 121350 9080
rect 120950 8850 121110 8930
rect 121190 8850 121350 8930
rect 120950 8680 121350 8850
rect 121650 8930 122050 9080
rect 121650 8850 121810 8930
rect 121890 8850 122050 8930
rect 121650 8680 122050 8850
rect 122350 8930 122750 9080
rect 122350 8850 122510 8930
rect 122590 8850 122750 8930
rect 122350 8680 122750 8850
rect 123050 8930 123450 9080
rect 123050 8850 123210 8930
rect 123290 8850 123450 8930
rect 123050 8680 123450 8850
rect 104150 8230 104550 8380
rect 104150 8150 104310 8230
rect 104390 8150 104550 8230
rect 104150 7980 104550 8150
rect 104850 8230 105250 8380
rect 104850 8150 105010 8230
rect 105090 8150 105250 8230
rect 104850 7980 105250 8150
rect 105550 8230 105950 8380
rect 105550 8150 105710 8230
rect 105790 8150 105950 8230
rect 105550 7980 105950 8150
rect 106250 8230 106650 8380
rect 106250 8150 106410 8230
rect 106490 8150 106650 8230
rect 106250 7980 106650 8150
rect 106950 8230 107350 8380
rect 106950 8150 107110 8230
rect 107190 8150 107350 8230
rect 106950 7980 107350 8150
rect 120250 8230 120650 8380
rect 120250 8150 120410 8230
rect 120490 8150 120650 8230
rect 120250 7980 120650 8150
rect 120950 8230 121350 8380
rect 120950 8150 121110 8230
rect 121190 8150 121350 8230
rect 120950 7980 121350 8150
rect 121650 8230 122050 8380
rect 121650 8150 121810 8230
rect 121890 8150 122050 8230
rect 121650 7980 122050 8150
rect 122350 8230 122750 8380
rect 122350 8150 122510 8230
rect 122590 8150 122750 8230
rect 122350 7980 122750 8150
rect 123050 8230 123450 8380
rect 123050 8150 123210 8230
rect 123290 8150 123450 8230
rect 123050 7980 123450 8150
rect 104150 7530 104550 7680
rect 104150 7450 104310 7530
rect 104390 7450 104550 7530
rect 104150 7280 104550 7450
rect 104850 7530 105250 7680
rect 104850 7450 105010 7530
rect 105090 7450 105250 7530
rect 104850 7280 105250 7450
rect 105550 7530 105950 7680
rect 105550 7450 105710 7530
rect 105790 7450 105950 7530
rect 105550 7280 105950 7450
rect 106250 7530 106650 7680
rect 106250 7450 106410 7530
rect 106490 7450 106650 7530
rect 106250 7280 106650 7450
rect 106950 7530 107350 7680
rect 106950 7450 107110 7530
rect 107190 7450 107350 7530
rect 106950 7280 107350 7450
rect 120250 7530 120650 7680
rect 120250 7450 120410 7530
rect 120490 7450 120650 7530
rect 120250 7280 120650 7450
rect 120950 7530 121350 7680
rect 120950 7450 121110 7530
rect 121190 7450 121350 7530
rect 120950 7280 121350 7450
rect 121650 7530 122050 7680
rect 121650 7450 121810 7530
rect 121890 7450 122050 7530
rect 121650 7280 122050 7450
rect 122350 7530 122750 7680
rect 122350 7450 122510 7530
rect 122590 7450 122750 7530
rect 122350 7280 122750 7450
rect 123050 7530 123450 7680
rect 123050 7450 123210 7530
rect 123290 7450 123450 7530
rect 123050 7280 123450 7450
rect 104150 6830 104550 6980
rect 104150 6750 104310 6830
rect 104390 6750 104550 6830
rect 104150 6580 104550 6750
rect 104850 6830 105250 6980
rect 104850 6750 105010 6830
rect 105090 6750 105250 6830
rect 104850 6580 105250 6750
rect 105550 6830 105950 6980
rect 105550 6750 105710 6830
rect 105790 6750 105950 6830
rect 105550 6580 105950 6750
rect 106250 6830 106650 6980
rect 106250 6750 106410 6830
rect 106490 6750 106650 6830
rect 106250 6580 106650 6750
rect 106950 6830 107350 6980
rect 106950 6750 107110 6830
rect 107190 6750 107350 6830
rect 106950 6580 107350 6750
rect 120250 6830 120650 6980
rect 120250 6750 120410 6830
rect 120490 6750 120650 6830
rect 120250 6580 120650 6750
rect 120950 6830 121350 6980
rect 120950 6750 121110 6830
rect 121190 6750 121350 6830
rect 120950 6580 121350 6750
rect 121650 6830 122050 6980
rect 121650 6750 121810 6830
rect 121890 6750 122050 6830
rect 121650 6580 122050 6750
rect 122350 6830 122750 6980
rect 122350 6750 122510 6830
rect 122590 6750 122750 6830
rect 122350 6580 122750 6750
rect 123050 6830 123450 6980
rect 123050 6750 123210 6830
rect 123290 6750 123450 6830
rect 123050 6580 123450 6750
rect 104150 6130 104550 6280
rect 104150 6050 104310 6130
rect 104390 6050 104550 6130
rect 104150 5880 104550 6050
rect 104850 6130 105250 6280
rect 104850 6050 105010 6130
rect 105090 6050 105250 6130
rect 104850 5880 105250 6050
rect 105550 6130 105950 6280
rect 105550 6050 105710 6130
rect 105790 6050 105950 6130
rect 105550 5880 105950 6050
rect 106250 6130 106650 6280
rect 106250 6050 106410 6130
rect 106490 6050 106650 6130
rect 106250 5880 106650 6050
rect 106950 6130 107350 6280
rect 106950 6050 107110 6130
rect 107190 6050 107350 6130
rect 106950 5880 107350 6050
rect 120250 6130 120650 6280
rect 120250 6050 120410 6130
rect 120490 6050 120650 6130
rect 120250 5880 120650 6050
rect 120950 6130 121350 6280
rect 120950 6050 121110 6130
rect 121190 6050 121350 6130
rect 120950 5880 121350 6050
rect 121650 6130 122050 6280
rect 121650 6050 121810 6130
rect 121890 6050 122050 6130
rect 121650 5880 122050 6050
rect 122350 6130 122750 6280
rect 122350 6050 122510 6130
rect 122590 6050 122750 6130
rect 122350 5880 122750 6050
rect 123050 6130 123450 6280
rect 123050 6050 123210 6130
rect 123290 6050 123450 6130
rect 123050 5880 123450 6050
rect 104150 5430 104550 5580
rect 104150 5350 104310 5430
rect 104390 5350 104550 5430
rect 104150 5180 104550 5350
rect 104850 5430 105250 5580
rect 104850 5350 105010 5430
rect 105090 5350 105250 5430
rect 104850 5180 105250 5350
rect 105550 5430 105950 5580
rect 105550 5350 105710 5430
rect 105790 5350 105950 5430
rect 105550 5180 105950 5350
rect 106250 5430 106650 5580
rect 106250 5350 106410 5430
rect 106490 5350 106650 5430
rect 106250 5180 106650 5350
rect 106950 5430 107350 5580
rect 106950 5350 107110 5430
rect 107190 5350 107350 5430
rect 106950 5180 107350 5350
rect 120250 5430 120650 5580
rect 120250 5350 120410 5430
rect 120490 5350 120650 5430
rect 120250 5180 120650 5350
rect 120950 5430 121350 5580
rect 120950 5350 121110 5430
rect 121190 5350 121350 5430
rect 120950 5180 121350 5350
rect 121650 5430 122050 5580
rect 121650 5350 121810 5430
rect 121890 5350 122050 5430
rect 121650 5180 122050 5350
rect 122350 5430 122750 5580
rect 122350 5350 122510 5430
rect 122590 5350 122750 5430
rect 122350 5180 122750 5350
rect 123050 5430 123450 5580
rect 123050 5350 123210 5430
rect 123290 5350 123450 5430
rect 123050 5180 123450 5350
rect 104150 4730 104550 4880
rect 104150 4650 104310 4730
rect 104390 4650 104550 4730
rect 104150 4480 104550 4650
rect 104850 4730 105250 4880
rect 104850 4650 105010 4730
rect 105090 4650 105250 4730
rect 104850 4480 105250 4650
rect 105550 4730 105950 4880
rect 105550 4650 105710 4730
rect 105790 4650 105950 4730
rect 105550 4480 105950 4650
rect 106250 4730 106650 4880
rect 106250 4650 106410 4730
rect 106490 4650 106650 4730
rect 106250 4480 106650 4650
rect 106950 4730 107350 4880
rect 106950 4650 107110 4730
rect 107190 4650 107350 4730
rect 106950 4480 107350 4650
rect 120250 4730 120650 4880
rect 120250 4650 120410 4730
rect 120490 4650 120650 4730
rect 120250 4480 120650 4650
rect 120950 4730 121350 4880
rect 120950 4650 121110 4730
rect 121190 4650 121350 4730
rect 120950 4480 121350 4650
rect 121650 4730 122050 4880
rect 121650 4650 121810 4730
rect 121890 4650 122050 4730
rect 121650 4480 122050 4650
rect 122350 4730 122750 4880
rect 122350 4650 122510 4730
rect 122590 4650 122750 4730
rect 122350 4480 122750 4650
rect 123050 4730 123450 4880
rect 123050 4650 123210 4730
rect 123290 4650 123450 4730
rect 123050 4480 123450 4650
rect 104150 4030 104550 4180
rect 104150 3950 104310 4030
rect 104390 3950 104550 4030
rect 104150 3780 104550 3950
rect 104850 4030 105250 4180
rect 104850 3950 105010 4030
rect 105090 3950 105250 4030
rect 104850 3780 105250 3950
rect 105550 4030 105950 4180
rect 105550 3950 105710 4030
rect 105790 3950 105950 4030
rect 105550 3780 105950 3950
rect 106250 4030 106650 4180
rect 106250 3950 106410 4030
rect 106490 3950 106650 4030
rect 106250 3780 106650 3950
rect 106950 4030 107350 4180
rect 106950 3950 107110 4030
rect 107190 3950 107350 4030
rect 106950 3780 107350 3950
rect 120250 4030 120650 4180
rect 120250 3950 120410 4030
rect 120490 3950 120650 4030
rect 120250 3780 120650 3950
rect 120950 4030 121350 4180
rect 120950 3950 121110 4030
rect 121190 3950 121350 4030
rect 120950 3780 121350 3950
rect 121650 4030 122050 4180
rect 121650 3950 121810 4030
rect 121890 3950 122050 4030
rect 121650 3780 122050 3950
rect 122350 4030 122750 4180
rect 122350 3950 122510 4030
rect 122590 3950 122750 4030
rect 122350 3780 122750 3950
rect 123050 4030 123450 4180
rect 123050 3950 123210 4030
rect 123290 3950 123450 4030
rect 123050 3780 123450 3950
rect 104150 3330 104550 3480
rect 104150 3250 104310 3330
rect 104390 3250 104550 3330
rect 104150 3080 104550 3250
rect 104850 3330 105250 3480
rect 104850 3250 105010 3330
rect 105090 3250 105250 3330
rect 104850 3080 105250 3250
rect 105550 3330 105950 3480
rect 105550 3250 105710 3330
rect 105790 3250 105950 3330
rect 105550 3080 105950 3250
rect 106250 3330 106650 3480
rect 106250 3250 106410 3330
rect 106490 3250 106650 3330
rect 106250 3080 106650 3250
rect 106950 3330 107350 3480
rect 106950 3250 107110 3330
rect 107190 3250 107350 3330
rect 106950 3080 107350 3250
rect 120250 3330 120650 3480
rect 120250 3250 120410 3330
rect 120490 3250 120650 3330
rect 120250 3080 120650 3250
rect 120950 3330 121350 3480
rect 120950 3250 121110 3330
rect 121190 3250 121350 3330
rect 120950 3080 121350 3250
rect 121650 3330 122050 3480
rect 121650 3250 121810 3330
rect 121890 3250 122050 3330
rect 121650 3080 122050 3250
rect 122350 3330 122750 3480
rect 122350 3250 122510 3330
rect 122590 3250 122750 3330
rect 122350 3080 122750 3250
rect 123050 3330 123450 3480
rect 123050 3250 123210 3330
rect 123290 3250 123450 3330
rect 123050 3080 123450 3250
rect 104150 2630 104550 2780
rect 104150 2550 104310 2630
rect 104390 2550 104550 2630
rect 104150 2380 104550 2550
rect 104850 2630 105250 2780
rect 104850 2550 105010 2630
rect 105090 2550 105250 2630
rect 104850 2380 105250 2550
rect 105550 2630 105950 2780
rect 105550 2550 105710 2630
rect 105790 2550 105950 2630
rect 105550 2380 105950 2550
rect 106250 2630 106650 2780
rect 106250 2550 106410 2630
rect 106490 2550 106650 2630
rect 106250 2380 106650 2550
rect 106950 2630 107350 2780
rect 106950 2550 107110 2630
rect 107190 2550 107350 2630
rect 106950 2380 107350 2550
rect 120250 2630 120650 2780
rect 120250 2550 120410 2630
rect 120490 2550 120650 2630
rect 120250 2380 120650 2550
rect 120950 2630 121350 2780
rect 120950 2550 121110 2630
rect 121190 2550 121350 2630
rect 120950 2380 121350 2550
rect 121650 2630 122050 2780
rect 121650 2550 121810 2630
rect 121890 2550 122050 2630
rect 121650 2380 122050 2550
rect 122350 2630 122750 2780
rect 122350 2550 122510 2630
rect 122590 2550 122750 2630
rect 122350 2380 122750 2550
rect 123050 2630 123450 2780
rect 123050 2550 123210 2630
rect 123290 2550 123450 2630
rect 123050 2380 123450 2550
rect 104150 1930 104550 2080
rect 104150 1850 104310 1930
rect 104390 1850 104550 1930
rect 104150 1680 104550 1850
rect 104850 1930 105250 2080
rect 104850 1850 105010 1930
rect 105090 1850 105250 1930
rect 104850 1680 105250 1850
rect 105550 1930 105950 2080
rect 105550 1850 105710 1930
rect 105790 1850 105950 1930
rect 105550 1680 105950 1850
rect 106250 1930 106650 2080
rect 106250 1850 106410 1930
rect 106490 1850 106650 1930
rect 106250 1680 106650 1850
rect 106950 1930 107350 2080
rect 106950 1850 107110 1930
rect 107190 1850 107350 1930
rect 106950 1680 107350 1850
rect 120250 1930 120650 2080
rect 120250 1850 120410 1930
rect 120490 1850 120650 1930
rect 120250 1680 120650 1850
rect 120950 1930 121350 2080
rect 120950 1850 121110 1930
rect 121190 1850 121350 1930
rect 120950 1680 121350 1850
rect 121650 1930 122050 2080
rect 121650 1850 121810 1930
rect 121890 1850 122050 1930
rect 121650 1680 122050 1850
rect 122350 1930 122750 2080
rect 122350 1850 122510 1930
rect 122590 1850 122750 1930
rect 122350 1680 122750 1850
rect 123050 1930 123450 2080
rect 123050 1850 123210 1930
rect 123290 1850 123450 1930
rect 123050 1680 123450 1850
rect 104150 1230 104550 1380
rect 104150 1150 104310 1230
rect 104390 1150 104550 1230
rect 104150 980 104550 1150
rect 104850 1230 105250 1380
rect 104850 1150 105010 1230
rect 105090 1150 105250 1230
rect 104850 980 105250 1150
rect 105550 1230 105950 1380
rect 105550 1150 105710 1230
rect 105790 1150 105950 1230
rect 105550 980 105950 1150
rect 106250 1230 106650 1380
rect 106250 1150 106410 1230
rect 106490 1150 106650 1230
rect 106250 980 106650 1150
rect 106950 1230 107350 1380
rect 106950 1150 107110 1230
rect 107190 1150 107350 1230
rect 106950 980 107350 1150
rect 120250 1230 120650 1380
rect 120250 1150 120410 1230
rect 120490 1150 120650 1230
rect 120250 980 120650 1150
rect 120950 1230 121350 1380
rect 120950 1150 121110 1230
rect 121190 1150 121350 1230
rect 120950 980 121350 1150
rect 121650 1230 122050 1380
rect 121650 1150 121810 1230
rect 121890 1150 122050 1230
rect 121650 980 122050 1150
rect 122350 1230 122750 1380
rect 122350 1150 122510 1230
rect 122590 1150 122750 1230
rect 122350 980 122750 1150
rect 123050 1230 123450 1380
rect 123050 1150 123210 1230
rect 123290 1150 123450 1230
rect 123050 980 123450 1150
rect 104150 530 104550 680
rect 104150 450 104310 530
rect 104390 450 104550 530
rect 104150 280 104550 450
rect 104850 530 105250 680
rect 104850 450 105010 530
rect 105090 450 105250 530
rect 104850 280 105250 450
rect 105550 530 105950 680
rect 105550 450 105710 530
rect 105790 450 105950 530
rect 105550 280 105950 450
rect 106250 530 106650 680
rect 106250 450 106410 530
rect 106490 450 106650 530
rect 106250 280 106650 450
rect 106950 530 107350 680
rect 106950 450 107110 530
rect 107190 450 107350 530
rect 106950 280 107350 450
rect 120250 530 120650 680
rect 120250 450 120410 530
rect 120490 450 120650 530
rect 120250 280 120650 450
rect 120950 530 121350 680
rect 120950 450 121110 530
rect 121190 450 121350 530
rect 120950 280 121350 450
rect 121650 530 122050 680
rect 121650 450 121810 530
rect 121890 450 122050 530
rect 121650 280 122050 450
rect 122350 530 122750 680
rect 122350 450 122510 530
rect 122590 450 122750 530
rect 122350 280 122750 450
rect 123050 530 123450 680
rect 123050 450 123210 530
rect 123290 450 123450 530
rect 123050 280 123450 450
rect 104150 -170 104550 -20
rect 104150 -250 104310 -170
rect 104390 -250 104550 -170
rect 104150 -420 104550 -250
rect 104850 -170 105250 -20
rect 104850 -250 105010 -170
rect 105090 -250 105250 -170
rect 104850 -420 105250 -250
rect 105550 -170 105950 -20
rect 105550 -250 105710 -170
rect 105790 -250 105950 -170
rect 105550 -420 105950 -250
rect 106250 -170 106650 -20
rect 106250 -250 106410 -170
rect 106490 -250 106650 -170
rect 106250 -420 106650 -250
rect 106950 -170 107350 -20
rect 106950 -250 107110 -170
rect 107190 -250 107350 -170
rect 106950 -420 107350 -250
rect 120250 -170 120650 -20
rect 120250 -250 120410 -170
rect 120490 -250 120650 -170
rect 120250 -420 120650 -250
rect 120950 -170 121350 -20
rect 120950 -250 121110 -170
rect 121190 -250 121350 -170
rect 120950 -420 121350 -250
rect 121650 -170 122050 -20
rect 121650 -250 121810 -170
rect 121890 -250 122050 -170
rect 121650 -420 122050 -250
rect 122350 -170 122750 -20
rect 122350 -250 122510 -170
rect 122590 -250 122750 -170
rect 122350 -420 122750 -250
rect 123050 -170 123450 -20
rect 123050 -250 123210 -170
rect 123290 -250 123450 -170
rect 123050 -420 123450 -250
rect 104150 -870 104550 -720
rect 104150 -950 104310 -870
rect 104390 -950 104550 -870
rect 104150 -1120 104550 -950
rect 104850 -870 105250 -720
rect 104850 -950 105010 -870
rect 105090 -950 105250 -870
rect 104850 -1120 105250 -950
rect 105550 -870 105950 -720
rect 105550 -950 105710 -870
rect 105790 -950 105950 -870
rect 105550 -1120 105950 -950
rect 106250 -870 106650 -720
rect 106250 -950 106410 -870
rect 106490 -950 106650 -870
rect 106250 -1120 106650 -950
rect 106950 -870 107350 -720
rect 106950 -950 107110 -870
rect 107190 -950 107350 -870
rect 106950 -1120 107350 -950
rect 120250 -870 120650 -720
rect 120250 -950 120410 -870
rect 120490 -950 120650 -870
rect 120250 -1120 120650 -950
rect 120950 -870 121350 -720
rect 120950 -950 121110 -870
rect 121190 -950 121350 -870
rect 120950 -1120 121350 -950
rect 121650 -870 122050 -720
rect 121650 -950 121810 -870
rect 121890 -950 122050 -870
rect 121650 -1120 122050 -950
rect 122350 -870 122750 -720
rect 122350 -950 122510 -870
rect 122590 -950 122750 -870
rect 122350 -1120 122750 -950
rect 123050 -870 123450 -720
rect 123050 -950 123210 -870
rect 123290 -950 123450 -870
rect 123050 -1120 123450 -950
rect 104150 -1570 104550 -1420
rect 104150 -1650 104310 -1570
rect 104390 -1650 104550 -1570
rect 104150 -1820 104550 -1650
rect 104850 -1570 105250 -1420
rect 104850 -1650 105010 -1570
rect 105090 -1650 105250 -1570
rect 104850 -1820 105250 -1650
rect 105550 -1570 105950 -1420
rect 105550 -1650 105710 -1570
rect 105790 -1650 105950 -1570
rect 105550 -1820 105950 -1650
rect 106250 -1570 106650 -1420
rect 106250 -1650 106410 -1570
rect 106490 -1650 106650 -1570
rect 106250 -1820 106650 -1650
rect 106950 -1570 107350 -1420
rect 106950 -1650 107110 -1570
rect 107190 -1650 107350 -1570
rect 106950 -1820 107350 -1650
rect 107650 -1570 108050 -1420
rect 107650 -1650 107810 -1570
rect 107890 -1650 108050 -1570
rect 107650 -1820 108050 -1650
rect 108350 -1570 108750 -1420
rect 108350 -1650 108510 -1570
rect 108590 -1650 108750 -1570
rect 108350 -1820 108750 -1650
rect 109050 -1570 109450 -1420
rect 109050 -1650 109210 -1570
rect 109290 -1650 109450 -1570
rect 109050 -1820 109450 -1650
rect 109750 -1570 110150 -1420
rect 109750 -1650 109910 -1570
rect 109990 -1650 110150 -1570
rect 109750 -1820 110150 -1650
rect 110450 -1570 110850 -1420
rect 110450 -1650 110610 -1570
rect 110690 -1650 110850 -1570
rect 110450 -1820 110850 -1650
rect 111150 -1570 111550 -1420
rect 111150 -1650 111310 -1570
rect 111390 -1650 111550 -1570
rect 111150 -1820 111550 -1650
rect 111850 -1570 112250 -1420
rect 111850 -1650 112010 -1570
rect 112090 -1650 112250 -1570
rect 111850 -1820 112250 -1650
rect 112550 -1570 112950 -1420
rect 112550 -1650 112710 -1570
rect 112790 -1650 112950 -1570
rect 112550 -1820 112950 -1650
rect 113250 -1570 113650 -1420
rect 113250 -1650 113410 -1570
rect 113490 -1650 113650 -1570
rect 113250 -1820 113650 -1650
rect 113950 -1570 114350 -1420
rect 113950 -1650 114110 -1570
rect 114190 -1650 114350 -1570
rect 113950 -1820 114350 -1650
rect 114650 -1570 115050 -1420
rect 114650 -1650 114810 -1570
rect 114890 -1650 115050 -1570
rect 114650 -1820 115050 -1650
rect 115350 -1570 115750 -1420
rect 115350 -1650 115510 -1570
rect 115590 -1650 115750 -1570
rect 115350 -1820 115750 -1650
rect 116050 -1570 116450 -1420
rect 116050 -1650 116210 -1570
rect 116290 -1650 116450 -1570
rect 116050 -1820 116450 -1650
rect 116750 -1570 117150 -1420
rect 116750 -1650 116910 -1570
rect 116990 -1650 117150 -1570
rect 116750 -1820 117150 -1650
rect 117450 -1570 117850 -1420
rect 117450 -1650 117610 -1570
rect 117690 -1650 117850 -1570
rect 117450 -1820 117850 -1650
rect 118150 -1570 118550 -1420
rect 118150 -1650 118310 -1570
rect 118390 -1650 118550 -1570
rect 118150 -1820 118550 -1650
rect 118850 -1570 119250 -1420
rect 118850 -1650 119010 -1570
rect 119090 -1650 119250 -1570
rect 118850 -1820 119250 -1650
rect 119550 -1570 119950 -1420
rect 119550 -1650 119710 -1570
rect 119790 -1650 119950 -1570
rect 119550 -1820 119950 -1650
rect 120250 -1570 120650 -1420
rect 120250 -1650 120410 -1570
rect 120490 -1650 120650 -1570
rect 120250 -1820 120650 -1650
rect 120950 -1570 121350 -1420
rect 120950 -1650 121110 -1570
rect 121190 -1650 121350 -1570
rect 120950 -1820 121350 -1650
rect 121650 -1570 122050 -1420
rect 121650 -1650 121810 -1570
rect 121890 -1650 122050 -1570
rect 121650 -1820 122050 -1650
rect 122350 -1570 122750 -1420
rect 122350 -1650 122510 -1570
rect 122590 -1650 122750 -1570
rect 122350 -1820 122750 -1650
rect 123050 -1570 123450 -1420
rect 123050 -1650 123210 -1570
rect 123290 -1650 123450 -1570
rect 123050 -1820 123450 -1650
rect 104150 -2270 104550 -2120
rect 104150 -2350 104310 -2270
rect 104390 -2350 104550 -2270
rect 104150 -2520 104550 -2350
rect 104850 -2270 105250 -2120
rect 104850 -2350 105010 -2270
rect 105090 -2350 105250 -2270
rect 104850 -2520 105250 -2350
rect 105550 -2270 105950 -2120
rect 105550 -2350 105710 -2270
rect 105790 -2350 105950 -2270
rect 105550 -2520 105950 -2350
rect 106250 -2270 106650 -2120
rect 106250 -2350 106410 -2270
rect 106490 -2350 106650 -2270
rect 106250 -2520 106650 -2350
rect 106950 -2270 107350 -2120
rect 106950 -2350 107110 -2270
rect 107190 -2350 107350 -2270
rect 106950 -2520 107350 -2350
rect 107650 -2270 108050 -2120
rect 107650 -2350 107810 -2270
rect 107890 -2350 108050 -2270
rect 107650 -2520 108050 -2350
rect 108350 -2270 108750 -2120
rect 108350 -2350 108510 -2270
rect 108590 -2350 108750 -2270
rect 108350 -2520 108750 -2350
rect 109050 -2270 109450 -2120
rect 109050 -2350 109210 -2270
rect 109290 -2350 109450 -2270
rect 109050 -2520 109450 -2350
rect 109750 -2270 110150 -2120
rect 109750 -2350 109910 -2270
rect 109990 -2350 110150 -2270
rect 109750 -2520 110150 -2350
rect 110450 -2270 110850 -2120
rect 110450 -2350 110610 -2270
rect 110690 -2350 110850 -2270
rect 110450 -2520 110850 -2350
rect 111150 -2270 111550 -2120
rect 111150 -2350 111310 -2270
rect 111390 -2350 111550 -2270
rect 111150 -2520 111550 -2350
rect 111850 -2270 112250 -2120
rect 111850 -2350 112010 -2270
rect 112090 -2350 112250 -2270
rect 111850 -2520 112250 -2350
rect 112550 -2270 112950 -2120
rect 112550 -2350 112710 -2270
rect 112790 -2350 112950 -2270
rect 112550 -2520 112950 -2350
rect 113250 -2270 113650 -2120
rect 113250 -2350 113410 -2270
rect 113490 -2350 113650 -2270
rect 113250 -2520 113650 -2350
rect 113950 -2270 114350 -2120
rect 113950 -2350 114110 -2270
rect 114190 -2350 114350 -2270
rect 113950 -2520 114350 -2350
rect 114650 -2270 115050 -2120
rect 114650 -2350 114810 -2270
rect 114890 -2350 115050 -2270
rect 114650 -2520 115050 -2350
rect 115350 -2270 115750 -2120
rect 115350 -2350 115510 -2270
rect 115590 -2350 115750 -2270
rect 115350 -2520 115750 -2350
rect 116050 -2270 116450 -2120
rect 116050 -2350 116210 -2270
rect 116290 -2350 116450 -2270
rect 116050 -2520 116450 -2350
rect 116750 -2270 117150 -2120
rect 116750 -2350 116910 -2270
rect 116990 -2350 117150 -2270
rect 116750 -2520 117150 -2350
rect 117450 -2270 117850 -2120
rect 117450 -2350 117610 -2270
rect 117690 -2350 117850 -2270
rect 117450 -2520 117850 -2350
rect 118150 -2270 118550 -2120
rect 118150 -2350 118310 -2270
rect 118390 -2350 118550 -2270
rect 118150 -2520 118550 -2350
rect 118850 -2270 119250 -2120
rect 118850 -2350 119010 -2270
rect 119090 -2350 119250 -2270
rect 118850 -2520 119250 -2350
rect 119550 -2270 119950 -2120
rect 119550 -2350 119710 -2270
rect 119790 -2350 119950 -2270
rect 119550 -2520 119950 -2350
rect 120250 -2270 120650 -2120
rect 120250 -2350 120410 -2270
rect 120490 -2350 120650 -2270
rect 120250 -2520 120650 -2350
rect 120950 -2270 121350 -2120
rect 120950 -2350 121110 -2270
rect 121190 -2350 121350 -2270
rect 120950 -2520 121350 -2350
rect 121650 -2270 122050 -2120
rect 121650 -2350 121810 -2270
rect 121890 -2350 122050 -2270
rect 121650 -2520 122050 -2350
rect 122350 -2270 122750 -2120
rect 122350 -2350 122510 -2270
rect 122590 -2350 122750 -2270
rect 122350 -2520 122750 -2350
rect 123050 -2270 123450 -2120
rect 123050 -2350 123210 -2270
rect 123290 -2350 123450 -2270
rect 123050 -2520 123450 -2350
<< mimcapcontact >>
rect 104310 10950 104390 11030
rect 105010 10950 105090 11030
rect 105710 10950 105790 11030
rect 106410 10950 106490 11030
rect 107110 10950 107190 11030
rect 107810 10950 107890 11030
rect 108510 10950 108590 11030
rect 109210 10950 109290 11030
rect 109910 10950 109990 11030
rect 110610 10950 110690 11030
rect 111310 10950 111390 11030
rect 112010 10950 112090 11030
rect 112710 10950 112790 11030
rect 113410 10950 113490 11030
rect 114110 10950 114190 11030
rect 114810 10950 114890 11030
rect 115510 10950 115590 11030
rect 116210 10950 116290 11030
rect 116910 10950 116990 11030
rect 117610 10950 117690 11030
rect 118310 10950 118390 11030
rect 119010 10950 119090 11030
rect 119710 10950 119790 11030
rect 120410 10950 120490 11030
rect 121110 10950 121190 11030
rect 121810 10950 121890 11030
rect 122510 10950 122590 11030
rect 123210 10950 123290 11030
rect 104310 10250 104390 10330
rect 105010 10250 105090 10330
rect 105710 10250 105790 10330
rect 106410 10250 106490 10330
rect 107110 10250 107190 10330
rect 107810 10250 107890 10330
rect 108510 10250 108590 10330
rect 109210 10250 109290 10330
rect 109910 10250 109990 10330
rect 110610 10230 110690 10310
rect 111310 10230 111390 10310
rect 112010 10250 112090 10330
rect 112710 10230 112790 10310
rect 113410 10230 113490 10310
rect 114110 10230 114190 10310
rect 114810 10240 114890 10310
rect 115510 10250 115590 10330
rect 116210 10230 116290 10310
rect 116910 10240 116990 10310
rect 117610 10250 117690 10330
rect 118310 10250 118390 10330
rect 119010 10250 119090 10330
rect 119710 10250 119790 10330
rect 120410 10250 120490 10330
rect 121110 10250 121190 10330
rect 121810 10250 121890 10330
rect 122510 10250 122590 10330
rect 123210 10250 123290 10330
rect 104310 9550 104390 9630
rect 105010 9550 105090 9630
rect 105710 9550 105790 9630
rect 106410 9550 106490 9630
rect 107110 9550 107190 9630
rect 107810 9550 107890 9630
rect 108510 9550 108590 9630
rect 119010 9550 119090 9630
rect 119710 9550 119790 9630
rect 120410 9550 120490 9630
rect 121110 9550 121190 9630
rect 121810 9550 121890 9630
rect 122510 9550 122590 9630
rect 123210 9550 123290 9630
rect 104310 8850 104390 8930
rect 105010 8850 105090 8930
rect 105710 8850 105790 8930
rect 106410 8850 106490 8930
rect 107110 8850 107190 8930
rect 120410 8850 120490 8930
rect 121110 8850 121190 8930
rect 121810 8850 121890 8930
rect 122510 8850 122590 8930
rect 123210 8850 123290 8930
rect 104310 8150 104390 8230
rect 105010 8150 105090 8230
rect 105710 8150 105790 8230
rect 106410 8150 106490 8230
rect 107110 8150 107190 8230
rect 120410 8150 120490 8230
rect 121110 8150 121190 8230
rect 121810 8150 121890 8230
rect 122510 8150 122590 8230
rect 123210 8150 123290 8230
rect 104310 7450 104390 7530
rect 105010 7450 105090 7530
rect 105710 7450 105790 7530
rect 106410 7450 106490 7530
rect 107110 7450 107190 7530
rect 120410 7450 120490 7530
rect 121110 7450 121190 7530
rect 121810 7450 121890 7530
rect 122510 7450 122590 7530
rect 123210 7450 123290 7530
rect 104310 6750 104390 6830
rect 105010 6750 105090 6830
rect 105710 6750 105790 6830
rect 106410 6750 106490 6830
rect 107110 6750 107190 6830
rect 120410 6750 120490 6830
rect 121110 6750 121190 6830
rect 121810 6750 121890 6830
rect 122510 6750 122590 6830
rect 123210 6750 123290 6830
rect 104310 6050 104390 6130
rect 105010 6050 105090 6130
rect 105710 6050 105790 6130
rect 106410 6050 106490 6130
rect 107110 6050 107190 6130
rect 120410 6050 120490 6130
rect 121110 6050 121190 6130
rect 121810 6050 121890 6130
rect 122510 6050 122590 6130
rect 123210 6050 123290 6130
rect 104310 5350 104390 5430
rect 105010 5350 105090 5430
rect 105710 5350 105790 5430
rect 106410 5350 106490 5430
rect 107110 5350 107190 5430
rect 120410 5350 120490 5430
rect 121110 5350 121190 5430
rect 121810 5350 121890 5430
rect 122510 5350 122590 5430
rect 123210 5350 123290 5430
rect 104310 4650 104390 4730
rect 105010 4650 105090 4730
rect 105710 4650 105790 4730
rect 106410 4650 106490 4730
rect 107110 4650 107190 4730
rect 120410 4650 120490 4730
rect 121110 4650 121190 4730
rect 121810 4650 121890 4730
rect 122510 4650 122590 4730
rect 123210 4650 123290 4730
rect 104310 3950 104390 4030
rect 105010 3950 105090 4030
rect 105710 3950 105790 4030
rect 106410 3950 106490 4030
rect 107110 3950 107190 4030
rect 120410 3950 120490 4030
rect 121110 3950 121190 4030
rect 121810 3950 121890 4030
rect 122510 3950 122590 4030
rect 123210 3950 123290 4030
rect 104310 3250 104390 3330
rect 105010 3250 105090 3330
rect 105710 3250 105790 3330
rect 106410 3250 106490 3330
rect 107110 3250 107190 3330
rect 120410 3250 120490 3330
rect 121110 3250 121190 3330
rect 121810 3250 121890 3330
rect 122510 3250 122590 3330
rect 123210 3250 123290 3330
rect 104310 2550 104390 2630
rect 105010 2550 105090 2630
rect 105710 2550 105790 2630
rect 106410 2550 106490 2630
rect 107110 2550 107190 2630
rect 120410 2550 120490 2630
rect 121110 2550 121190 2630
rect 121810 2550 121890 2630
rect 122510 2550 122590 2630
rect 123210 2550 123290 2630
rect 104310 1850 104390 1930
rect 105010 1850 105090 1930
rect 105710 1850 105790 1930
rect 106410 1850 106490 1930
rect 107110 1850 107190 1930
rect 120410 1850 120490 1930
rect 121110 1850 121190 1930
rect 121810 1850 121890 1930
rect 122510 1850 122590 1930
rect 123210 1850 123290 1930
rect 104310 1150 104390 1230
rect 105010 1150 105090 1230
rect 105710 1150 105790 1230
rect 106410 1150 106490 1230
rect 107110 1150 107190 1230
rect 120410 1150 120490 1230
rect 121110 1150 121190 1230
rect 121810 1150 121890 1230
rect 122510 1150 122590 1230
rect 123210 1150 123290 1230
rect 104310 450 104390 530
rect 105010 450 105090 530
rect 105710 450 105790 530
rect 106410 450 106490 530
rect 107110 450 107190 530
rect 120410 450 120490 530
rect 121110 450 121190 530
rect 121810 450 121890 530
rect 122510 450 122590 530
rect 123210 450 123290 530
rect 104310 -250 104390 -170
rect 105010 -250 105090 -170
rect 105710 -250 105790 -170
rect 106410 -250 106490 -170
rect 107110 -250 107190 -170
rect 120410 -250 120490 -170
rect 121110 -250 121190 -170
rect 121810 -250 121890 -170
rect 122510 -250 122590 -170
rect 123210 -250 123290 -170
rect 104310 -950 104390 -870
rect 105010 -950 105090 -870
rect 105710 -950 105790 -870
rect 106410 -950 106490 -870
rect 107110 -950 107190 -870
rect 120410 -950 120490 -870
rect 121110 -950 121190 -870
rect 121810 -950 121890 -870
rect 122510 -950 122590 -870
rect 123210 -950 123290 -870
rect 104310 -1650 104390 -1570
rect 105010 -1650 105090 -1570
rect 105710 -1650 105790 -1570
rect 106410 -1650 106490 -1570
rect 107110 -1650 107190 -1570
rect 107810 -1650 107890 -1570
rect 108510 -1650 108590 -1570
rect 109210 -1650 109290 -1570
rect 109910 -1650 109990 -1570
rect 110610 -1650 110690 -1570
rect 111310 -1650 111390 -1570
rect 112010 -1650 112090 -1570
rect 112710 -1650 112790 -1570
rect 113410 -1650 113490 -1570
rect 114110 -1650 114190 -1570
rect 114810 -1650 114890 -1570
rect 115510 -1650 115590 -1570
rect 116210 -1650 116290 -1570
rect 116910 -1650 116990 -1570
rect 117610 -1650 117690 -1570
rect 118310 -1650 118390 -1570
rect 119010 -1650 119090 -1570
rect 119710 -1650 119790 -1570
rect 120410 -1650 120490 -1570
rect 121110 -1650 121190 -1570
rect 121810 -1650 121890 -1570
rect 122510 -1650 122590 -1570
rect 123210 -1650 123290 -1570
rect 104310 -2350 104390 -2270
rect 105010 -2350 105090 -2270
rect 105710 -2350 105790 -2270
rect 106410 -2350 106490 -2270
rect 107110 -2350 107190 -2270
rect 107810 -2350 107890 -2270
rect 108510 -2350 108590 -2270
rect 109210 -2350 109290 -2270
rect 109910 -2350 109990 -2270
rect 110610 -2350 110690 -2270
rect 111310 -2350 111390 -2270
rect 112010 -2350 112090 -2270
rect 112710 -2350 112790 -2270
rect 113410 -2350 113490 -2270
rect 114110 -2350 114190 -2270
rect 114810 -2350 114890 -2270
rect 115510 -2350 115590 -2270
rect 116210 -2350 116290 -2270
rect 116910 -2350 116990 -2270
rect 117610 -2350 117690 -2270
rect 118310 -2350 118390 -2270
rect 119010 -2350 119090 -2270
rect 119710 -2350 119790 -2270
rect 120410 -2350 120490 -2270
rect 121110 -2350 121190 -2270
rect 121810 -2350 121890 -2270
rect 122510 -2350 122590 -2270
rect 123210 -2350 123290 -2270
<< metal4 >>
rect 105700 11040 105800 11300
rect 121800 11040 121900 11290
rect 104300 11030 113500 11040
rect 104300 10950 104310 11030
rect 104390 10950 105010 11030
rect 105090 10950 105710 11030
rect 105790 10950 106410 11030
rect 106490 10950 107110 11030
rect 107190 10950 107810 11030
rect 107890 10950 108510 11030
rect 108590 10950 109210 11030
rect 109290 10950 109910 11030
rect 109990 10950 110610 11030
rect 110690 10950 111310 11030
rect 111390 10950 112010 11030
rect 112090 10950 112710 11030
rect 112790 10950 113410 11030
rect 113490 10950 113500 11030
rect 104300 10940 113500 10950
rect 105700 10340 105800 10940
rect 104300 10330 107200 10340
rect 104300 10250 104310 10330
rect 104390 10250 105010 10330
rect 105090 10250 105710 10330
rect 105790 10250 106410 10330
rect 106490 10250 107110 10330
rect 107190 10250 107200 10330
rect 104300 10240 107200 10250
rect 107800 10330 107900 10940
rect 107800 10250 107810 10330
rect 107890 10250 107900 10330
rect 105700 9640 105800 10240
rect 104300 9630 107200 9640
rect 104300 9550 104310 9630
rect 104390 9550 105010 9630
rect 105090 9550 105710 9630
rect 105790 9550 106410 9630
rect 106490 9550 107110 9630
rect 107190 9550 107200 9630
rect 104300 9540 107200 9550
rect 107800 9630 107900 10250
rect 107800 9550 107810 9630
rect 107890 9550 107900 9630
rect 107800 9540 107900 9550
rect 108500 10330 108600 10940
rect 108500 10250 108510 10330
rect 108590 10250 108600 10330
rect 108500 9630 108600 10250
rect 109200 10330 109300 10940
rect 109200 10250 109210 10330
rect 109290 10250 109300 10330
rect 109200 10220 109300 10250
rect 109900 10330 110000 10940
rect 109900 10250 109910 10330
rect 109990 10250 110000 10330
rect 109900 10220 110000 10250
rect 110600 10310 110700 10940
rect 110600 10230 110610 10310
rect 110690 10230 110700 10310
rect 110600 10220 110700 10230
rect 111300 10310 111400 10940
rect 111300 10230 111310 10310
rect 111390 10230 111400 10310
rect 111300 10220 111400 10230
rect 112000 10330 112100 10940
rect 112000 10250 112010 10330
rect 112090 10250 112100 10330
rect 112000 10220 112100 10250
rect 112700 10310 112800 10940
rect 112700 10230 112710 10310
rect 112790 10230 112800 10310
rect 112700 10220 112800 10230
rect 113400 10310 113500 10940
rect 113400 10230 113410 10310
rect 113490 10230 113500 10310
rect 113400 10220 113500 10230
rect 114100 11030 123300 11040
rect 114100 10950 114110 11030
rect 114190 10950 114810 11030
rect 114890 10950 115510 11030
rect 115590 10950 116210 11030
rect 116290 10950 116910 11030
rect 116990 10950 117610 11030
rect 117690 10950 118310 11030
rect 118390 10950 119010 11030
rect 119090 10950 119710 11030
rect 119790 10950 120410 11030
rect 120490 10950 121110 11030
rect 121190 10950 121810 11030
rect 121890 10950 122510 11030
rect 122590 10950 123210 11030
rect 123290 10950 123300 11030
rect 114100 10940 123300 10950
rect 114100 10310 114200 10940
rect 114100 10230 114110 10310
rect 114190 10230 114200 10310
rect 114800 10310 114900 10940
rect 114800 10240 114810 10310
rect 114890 10240 114900 10310
rect 115500 10330 115600 10940
rect 115500 10250 115510 10330
rect 115590 10250 115600 10330
rect 115500 10240 115600 10250
rect 116200 10310 116300 10940
rect 114100 10220 114200 10230
rect 116200 10230 116210 10310
rect 116290 10230 116300 10310
rect 116900 10310 117000 10940
rect 116900 10240 116910 10310
rect 116990 10240 117000 10310
rect 117600 10330 117700 10940
rect 117600 10250 117610 10330
rect 117690 10250 117700 10330
rect 117600 10240 117700 10250
rect 118300 10330 118400 10940
rect 118300 10250 118310 10330
rect 118390 10250 118400 10330
rect 118300 10240 118400 10250
rect 119000 10330 119100 10940
rect 119000 10250 119010 10330
rect 119090 10250 119100 10330
rect 116200 10220 116300 10230
rect 108500 9550 108510 9630
rect 108590 9550 108600 9630
rect 108500 9540 108600 9550
rect 119000 9630 119100 10250
rect 119000 9550 119010 9630
rect 119090 9550 119100 9630
rect 119000 9540 119100 9550
rect 119700 10330 119800 10940
rect 121800 10340 121900 10940
rect 119700 10250 119710 10330
rect 119790 10250 119800 10330
rect 119700 9630 119800 10250
rect 120400 10330 123300 10340
rect 120400 10250 120410 10330
rect 120490 10250 121110 10330
rect 121190 10250 121810 10330
rect 121890 10250 122510 10330
rect 122590 10250 123210 10330
rect 123290 10250 123300 10330
rect 120400 10240 123300 10250
rect 121800 9640 121900 10240
rect 119700 9550 119710 9630
rect 119790 9550 119800 9630
rect 119700 9540 119800 9550
rect 120400 9630 123300 9640
rect 120400 9550 120410 9630
rect 120490 9550 121110 9630
rect 121190 9550 121810 9630
rect 121890 9550 122510 9630
rect 122590 9550 123210 9630
rect 123290 9550 123300 9630
rect 120400 9540 123300 9550
rect 105700 8940 105800 9540
rect 121800 8940 121900 9540
rect 104300 8930 107200 8940
rect 104300 8850 104310 8930
rect 104390 8850 105010 8930
rect 105090 8850 105710 8930
rect 105790 8850 106410 8930
rect 106490 8850 107110 8930
rect 107190 8850 107200 8930
rect 104300 8840 107200 8850
rect 120400 8930 123300 8940
rect 120400 8850 120410 8930
rect 120490 8850 121110 8930
rect 121190 8850 121810 8930
rect 121890 8850 122510 8930
rect 122590 8850 123210 8930
rect 123290 8850 123300 8930
rect 120400 8840 123300 8850
rect 105700 8240 105800 8840
rect 121800 8240 121900 8840
rect 104300 8230 107200 8240
rect 104300 8150 104310 8230
rect 104390 8150 105010 8230
rect 105090 8150 105710 8230
rect 105790 8150 106410 8230
rect 106490 8150 107110 8230
rect 107190 8150 107200 8230
rect 104300 8140 107200 8150
rect 120400 8230 123300 8240
rect 120400 8150 120410 8230
rect 120490 8150 121110 8230
rect 121190 8150 121810 8230
rect 121890 8150 122510 8230
rect 122590 8150 123210 8230
rect 123290 8150 123300 8230
rect 120400 8140 123300 8150
rect 105700 7540 105800 8140
rect 121800 7540 121900 8140
rect 104300 7530 107200 7540
rect 104300 7450 104310 7530
rect 104390 7450 105010 7530
rect 105090 7450 105710 7530
rect 105790 7450 106410 7530
rect 106490 7450 107110 7530
rect 107190 7450 107200 7530
rect 104300 7440 107200 7450
rect 120400 7530 123300 7540
rect 120400 7450 120410 7530
rect 120490 7450 121110 7530
rect 121190 7450 121810 7530
rect 121890 7450 122510 7530
rect 122590 7450 123210 7530
rect 123290 7450 123300 7530
rect 120400 7440 123300 7450
rect 105700 6840 105800 7440
rect 121800 6840 121900 7440
rect 104300 6830 107200 6840
rect 104300 6750 104310 6830
rect 104390 6750 105010 6830
rect 105090 6750 105710 6830
rect 105790 6750 106410 6830
rect 106490 6750 107110 6830
rect 107190 6750 107200 6830
rect 104300 6740 107200 6750
rect 120400 6830 123300 6840
rect 120400 6750 120410 6830
rect 120490 6750 121110 6830
rect 121190 6750 121810 6830
rect 121890 6750 122510 6830
rect 122590 6750 123210 6830
rect 123290 6750 123300 6830
rect 120400 6740 123300 6750
rect 105700 6140 105800 6740
rect 121800 6140 121900 6740
rect 104300 6130 107200 6140
rect 104300 6050 104310 6130
rect 104390 6050 105010 6130
rect 105090 6050 105710 6130
rect 105790 6050 106410 6130
rect 106490 6050 107110 6130
rect 107190 6050 107200 6130
rect 104300 6040 107200 6050
rect 120400 6130 123300 6140
rect 120400 6050 120410 6130
rect 120490 6050 121110 6130
rect 121190 6050 121810 6130
rect 121890 6050 122510 6130
rect 122590 6050 123210 6130
rect 123290 6050 123300 6130
rect 120400 6040 123300 6050
rect 105700 5440 105800 6040
rect 121800 5440 121900 6040
rect 104300 5430 107200 5440
rect 104300 5350 104310 5430
rect 104390 5350 105010 5430
rect 105090 5350 105710 5430
rect 105790 5350 106410 5430
rect 106490 5350 107110 5430
rect 107190 5350 107200 5430
rect 104300 5340 107200 5350
rect 120400 5430 123300 5440
rect 120400 5350 120410 5430
rect 120490 5350 121110 5430
rect 121190 5350 121810 5430
rect 121890 5350 122510 5430
rect 122590 5350 123210 5430
rect 123290 5350 123300 5430
rect 120400 5340 123300 5350
rect 105700 4740 105800 5340
rect 121800 4740 121900 5340
rect 104300 4730 107200 4740
rect 104300 4650 104310 4730
rect 104390 4650 105010 4730
rect 105090 4650 105710 4730
rect 105790 4650 106410 4730
rect 106490 4650 107110 4730
rect 107190 4650 107200 4730
rect 104300 4640 107200 4650
rect 120400 4730 123300 4740
rect 120400 4650 120410 4730
rect 120490 4650 121110 4730
rect 121190 4650 121810 4730
rect 121890 4650 122510 4730
rect 122590 4650 123210 4730
rect 123290 4650 123300 4730
rect 120400 4640 123300 4650
rect 105700 4040 105800 4640
rect 107100 4130 108480 4140
rect 107100 4050 107990 4130
rect 108070 4050 108090 4130
rect 108170 4050 108190 4130
rect 108270 4050 108290 4130
rect 108370 4050 108390 4130
rect 108470 4050 108480 4130
rect 107100 4040 108480 4050
rect 104300 4030 108480 4040
rect 104300 3950 104310 4030
rect 104390 3950 105010 4030
rect 105090 3950 105710 4030
rect 105790 3950 106410 4030
rect 106490 3950 107110 4030
rect 107190 3950 107990 4030
rect 108070 3950 108090 4030
rect 108170 3950 108190 4030
rect 108270 3950 108290 4030
rect 108370 3950 108390 4030
rect 108470 3950 108480 4030
rect 104300 3940 108480 3950
rect 105700 3340 105800 3940
rect 107100 3930 108480 3940
rect 107100 3850 107990 3930
rect 108070 3850 108090 3930
rect 108170 3850 108190 3930
rect 108270 3850 108290 3930
rect 108370 3850 108390 3930
rect 108470 3850 108480 3930
rect 107100 3840 108480 3850
rect 119120 4130 120510 4140
rect 119120 4050 119130 4130
rect 119210 4050 119230 4130
rect 119310 4050 119330 4130
rect 119410 4050 119430 4130
rect 119510 4050 119530 4130
rect 119610 4050 120510 4130
rect 119120 4040 120510 4050
rect 121800 4040 121900 4640
rect 119120 4030 123300 4040
rect 119120 3950 119130 4030
rect 119210 3950 119230 4030
rect 119310 3950 119330 4030
rect 119410 3950 119430 4030
rect 119510 3950 119530 4030
rect 119610 3950 120410 4030
rect 120490 3950 121110 4030
rect 121190 3950 121810 4030
rect 121890 3950 122510 4030
rect 122590 3950 123210 4030
rect 123290 3950 123300 4030
rect 119120 3940 123300 3950
rect 119120 3930 120510 3940
rect 119120 3850 119130 3930
rect 119210 3850 119230 3930
rect 119310 3850 119330 3930
rect 119410 3850 119430 3930
rect 119510 3850 119530 3930
rect 119610 3850 120510 3930
rect 119120 3840 120510 3850
rect 121800 3340 121900 3940
rect 104300 3330 107200 3340
rect 104300 3250 104310 3330
rect 104390 3250 105010 3330
rect 105090 3250 105710 3330
rect 105790 3250 106410 3330
rect 106490 3250 107110 3330
rect 107190 3250 107200 3330
rect 104300 3240 107200 3250
rect 120400 3330 123300 3340
rect 120400 3250 120410 3330
rect 120490 3250 121110 3330
rect 121190 3250 121810 3330
rect 121890 3250 122510 3330
rect 122590 3250 123210 3330
rect 123290 3250 123300 3330
rect 120400 3240 123300 3250
rect 105700 2640 105800 3240
rect 121800 2640 121900 3240
rect 104300 2630 107200 2640
rect 104300 2550 104310 2630
rect 104390 2550 105010 2630
rect 105090 2550 105710 2630
rect 105790 2550 106410 2630
rect 106490 2550 107110 2630
rect 107190 2550 107200 2630
rect 104300 2540 107200 2550
rect 120400 2630 123300 2640
rect 120400 2550 120410 2630
rect 120490 2550 121110 2630
rect 121190 2550 121810 2630
rect 121890 2550 122510 2630
rect 122590 2550 123210 2630
rect 123290 2550 123300 2630
rect 120400 2540 123300 2550
rect 105700 1940 105800 2540
rect 121800 1940 121900 2540
rect 104300 1930 107200 1940
rect 104300 1850 104310 1930
rect 104390 1850 105010 1930
rect 105090 1850 105710 1930
rect 105790 1850 106410 1930
rect 106490 1850 107110 1930
rect 107190 1850 107200 1930
rect 104300 1840 107200 1850
rect 120400 1930 123300 1940
rect 120400 1850 120410 1930
rect 120490 1850 121110 1930
rect 121190 1850 121810 1930
rect 121890 1850 122510 1930
rect 122590 1850 123210 1930
rect 123290 1850 123300 1930
rect 120400 1840 123300 1850
rect 105700 1240 105800 1840
rect 121800 1240 121900 1840
rect 104300 1230 107200 1240
rect 104300 1150 104310 1230
rect 104390 1150 105010 1230
rect 105090 1150 105710 1230
rect 105790 1150 106410 1230
rect 106490 1150 107110 1230
rect 107190 1150 107200 1230
rect 104300 1140 107200 1150
rect 120400 1230 123300 1240
rect 120400 1150 120410 1230
rect 120490 1150 121110 1230
rect 121190 1150 121810 1230
rect 121890 1150 122510 1230
rect 122590 1150 123210 1230
rect 123290 1150 123300 1230
rect 120400 1140 123300 1150
rect 105700 540 105800 1140
rect 121800 540 121900 1140
rect 104300 530 107200 540
rect 104300 450 104310 530
rect 104390 450 105010 530
rect 105090 450 105710 530
rect 105790 450 106410 530
rect 106490 450 107110 530
rect 107190 450 107200 530
rect 104300 440 107200 450
rect 120400 530 123300 540
rect 120400 450 120410 530
rect 120490 450 121110 530
rect 121190 450 121810 530
rect 121890 450 122510 530
rect 122590 450 123210 530
rect 123290 450 123300 530
rect 120400 440 123300 450
rect 105700 -160 105800 440
rect 121800 -160 121900 440
rect 104300 -170 107200 -160
rect 104300 -250 104310 -170
rect 104390 -250 105010 -170
rect 105090 -250 105710 -170
rect 105790 -250 106410 -170
rect 106490 -250 107110 -170
rect 107190 -250 107200 -170
rect 104300 -260 107200 -250
rect 120400 -170 123300 -160
rect 120400 -250 120410 -170
rect 120490 -250 121110 -170
rect 121190 -250 121810 -170
rect 121890 -250 122510 -170
rect 122590 -250 123210 -170
rect 123290 -250 123300 -170
rect 120400 -260 123300 -250
rect 105700 -860 105800 -260
rect 121800 -860 121900 -260
rect 104300 -870 107200 -860
rect 104300 -950 104310 -870
rect 104390 -950 105010 -870
rect 105090 -950 105710 -870
rect 105790 -950 106410 -870
rect 106490 -950 107110 -870
rect 107190 -950 107200 -870
rect 104300 -960 107200 -950
rect 120400 -870 123300 -860
rect 120400 -950 120410 -870
rect 120490 -950 121110 -870
rect 121190 -950 121810 -870
rect 121890 -950 122510 -870
rect 122590 -950 123210 -870
rect 123290 -950 123300 -870
rect 120400 -960 123300 -950
rect 105700 -1560 105800 -960
rect 121800 -1560 121900 -960
rect 104300 -1570 113500 -1560
rect 104300 -1650 104310 -1570
rect 104390 -1650 105010 -1570
rect 105090 -1650 105710 -1570
rect 105790 -1650 106410 -1570
rect 106490 -1650 107110 -1570
rect 107190 -1650 107810 -1570
rect 107890 -1650 108510 -1570
rect 108590 -1650 109210 -1570
rect 109290 -1650 109910 -1570
rect 109990 -1650 110610 -1570
rect 110690 -1650 111310 -1570
rect 111390 -1650 112010 -1570
rect 112090 -1650 112710 -1570
rect 112790 -1650 113410 -1570
rect 113490 -1650 113500 -1570
rect 104300 -1660 113500 -1650
rect 105700 -2260 105800 -1660
rect 104300 -2270 105800 -2260
rect 104300 -2350 104310 -2270
rect 104390 -2350 105010 -2270
rect 105090 -2350 105710 -2270
rect 105790 -2350 105800 -2270
rect 104300 -2360 105800 -2350
rect 106400 -2270 106500 -1660
rect 106400 -2350 106410 -2270
rect 106490 -2350 106500 -2270
rect 106400 -2360 106500 -2350
rect 107100 -2270 107200 -1660
rect 107100 -2350 107110 -2270
rect 107190 -2350 107200 -2270
rect 107100 -2360 107200 -2350
rect 107800 -2270 107900 -1660
rect 107800 -2350 107810 -2270
rect 107890 -2350 107900 -2270
rect 107800 -2360 107900 -2350
rect 108500 -2270 108600 -1660
rect 108500 -2350 108510 -2270
rect 108590 -2350 108600 -2270
rect 108500 -2360 108600 -2350
rect 109200 -2270 109300 -1660
rect 109200 -2350 109210 -2270
rect 109290 -2350 109300 -2270
rect 109200 -2360 109300 -2350
rect 109900 -2270 110000 -1660
rect 109900 -2350 109910 -2270
rect 109990 -2350 110000 -2270
rect 109900 -2360 110000 -2350
rect 110600 -2270 110700 -1660
rect 110600 -2350 110610 -2270
rect 110690 -2350 110700 -2270
rect 110600 -2360 110700 -2350
rect 111300 -2270 111400 -1660
rect 111300 -2350 111310 -2270
rect 111390 -2350 111400 -2270
rect 111300 -2360 111400 -2350
rect 112000 -2270 112100 -1660
rect 112000 -2350 112010 -2270
rect 112090 -2350 112100 -2270
rect 112000 -2360 112100 -2350
rect 112700 -2270 112800 -1660
rect 112700 -2350 112710 -2270
rect 112790 -2350 112800 -2270
rect 112700 -2360 112800 -2350
rect 113400 -2270 113500 -1660
rect 113400 -2350 113410 -2270
rect 113490 -2350 113500 -2270
rect 113400 -2360 113500 -2350
rect 114100 -1570 123300 -1560
rect 114100 -1650 114110 -1570
rect 114190 -1650 114810 -1570
rect 114890 -1650 115510 -1570
rect 115590 -1650 116210 -1570
rect 116290 -1650 116910 -1570
rect 116990 -1650 117610 -1570
rect 117690 -1650 118310 -1570
rect 118390 -1650 119010 -1570
rect 119090 -1650 119710 -1570
rect 119790 -1650 120410 -1570
rect 120490 -1650 121110 -1570
rect 121190 -1650 121810 -1570
rect 121890 -1650 122510 -1570
rect 122590 -1650 123210 -1570
rect 123290 -1650 123300 -1570
rect 114100 -1660 123300 -1650
rect 114100 -2270 114200 -1660
rect 114100 -2350 114110 -2270
rect 114190 -2350 114200 -2270
rect 114100 -2360 114200 -2350
rect 114800 -2270 114900 -1660
rect 114800 -2350 114810 -2270
rect 114890 -2350 114900 -2270
rect 114800 -2360 114900 -2350
rect 115500 -2270 115600 -1660
rect 115500 -2350 115510 -2270
rect 115590 -2350 115600 -2270
rect 115500 -2360 115600 -2350
rect 116200 -2270 116300 -1660
rect 116200 -2350 116210 -2270
rect 116290 -2350 116300 -2270
rect 116200 -2360 116300 -2350
rect 116900 -2270 117000 -1660
rect 116900 -2350 116910 -2270
rect 116990 -2350 117000 -2270
rect 116900 -2360 117000 -2350
rect 117600 -2270 117700 -1660
rect 117600 -2350 117610 -2270
rect 117690 -2350 117700 -2270
rect 117600 -2360 117700 -2350
rect 118300 -2270 118400 -1660
rect 118300 -2350 118310 -2270
rect 118390 -2350 118400 -2270
rect 118300 -2360 118400 -2350
rect 119000 -2270 119100 -1660
rect 119000 -2350 119010 -2270
rect 119090 -2350 119100 -2270
rect 119000 -2360 119100 -2350
rect 119700 -2270 119800 -1660
rect 119700 -2350 119710 -2270
rect 119790 -2350 119800 -2270
rect 119700 -2360 119800 -2350
rect 120400 -2270 120500 -1660
rect 120400 -2350 120410 -2270
rect 120490 -2350 120500 -2270
rect 120400 -2360 120500 -2350
rect 121100 -2270 121200 -1660
rect 121100 -2350 121110 -2270
rect 121190 -2350 121200 -2270
rect 121100 -2360 121200 -2350
rect 121800 -2260 121900 -1660
rect 121800 -2270 123300 -2260
rect 121800 -2350 121810 -2270
rect 121890 -2350 122510 -2270
rect 122590 -2350 123210 -2270
rect 123290 -2350 123300 -2270
rect 121800 -2360 123300 -2350
<< labels >>
flabel metal2 110600 8420 110600 8420 5 FreeSans 480 0 0 -160 VD4
flabel metal2 117000 8420 117000 8420 5 FreeSans 480 0 0 -160 VD3
flabel metal2 112710 9860 112710 9860 1 FreeSans 480 0 0 160 Vb2_2
flabel metal2 114930 9860 114930 9860 1 FreeSans 480 0 0 160 Vb2_Vb3
flabel metal2 114800 8500 114800 8500 5 FreeSans 400 0 0 -160 Vb3
port 4 s
flabel metal1 111380 7390 111380 7390 5 FreeSans 400 0 0 -160 Vb2
port 5 s
flabel metal2 114360 8140 114360 8140 3 FreeSans 480 0 160 0 V_err_p
flabel metal1 113240 8140 113240 8140 7 FreeSans 480 0 -160 0 V_err_mir_p
flabel metal2 114250 7500 114250 7500 3 FreeSans 480 0 160 0 V_err_gate
port 13 e
flabel metal2 112730 7380 112730 7380 7 FreeSans 480 0 -160 0 V_err_amp_ref
port 12 w
flabel metal3 119080 7790 119080 7790 3 FreeSans 480 0 160 0 cap_res_X
flabel metal3 108510 7790 108510 7790 7 FreeSans 480 0 -160 0 cap_res_Y
flabel metal2 109100 3580 109100 3580 1 FreeSans 480 0 0 160 V_CMFB_S4
port 8 n
flabel metal1 112740 4070 112740 4070 7 FreeSans 480 0 -160 0 VD2
flabel metal1 114860 4070 114860 4070 3 FreeSans 480 0 160 0 VD1
flabel metal2 112060 3980 112060 3980 7 FreeSans 480 0 -160 0 VIN+
flabel metal2 115540 3980 115540 3980 3 FreeSans 480 0 160 0 VIN-
flabel metal2 114910 6950 114910 6950 7 FreeSans 480 0 -160 0 X
flabel metal1 112690 6930 112690 6930 3 FreeSans 480 0 160 0 Y
flabel metal2 115050 7060 115050 7060 1 FreeSans 480 0 0 160 err_amp_out
flabel metal2 114000 7150 114000 7150 3 FreeSans 480 0 160 0 err_amp_mir
flabel metal2 115160 7280 115160 7280 1 FreeSans 480 0 0 320 V_tot
flabel metal1 118590 3950 118590 3950 1 FreeSans 480 0 0 160 V_CMFB_S1
port 2 n
flabel metal1 118500 3580 118500 3580 1 FreeSans 480 0 0 160 V_CMFB_S2
port 7 n
flabel metal2 109010 3950 109010 3950 1 FreeSans 480 0 0 160 V_CMFB_S3
port 3 n
flabel metal1 113890 2120 113890 2120 7 FreeSans 480 0 -160 0 V_tail_gate
port 11 w
flabel metal2 112920 590 112920 590 1 FreeSans 480 0 0 160 V_p_mir
flabel metal1 114440 1950 114440 1950 3 FreeSans 480 0 160 0 V_source
flabel metal1 119410 1510 119410 1510 5 FreeSans 480 0 0 -160 VOUT-
port 9 s
flabel metal2 115440 1800 115440 1800 5 FreeSans 400 0 0 -160 V_b_2nd_stage
flabel metal2 108190 1510 108190 1510 5 FreeSans 480 0 0 -160 VOUT+
port 10 s
flabel metal2 113800 300 113800 300 1 FreeSans 480 0 0 160 Vb1_2
flabel metal2 113800 5790 113800 5790 5 FreeSans 480 0 0 -160 Vb1
<< end >>
