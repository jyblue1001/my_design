** sch_path: /foss/designs/my_design/projects/pnp/xschem_ngspice/tb_pnp.sch
**.subckt tb_pnp
Ve EMITTER GND 0.7
XQ1 EMITTER GND GND sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ2 EMITTER GND GND sky130_fd_pr__pnp_05v5_W0p68L0p68
**** begin user architecture code



.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.subckt sky130_fd_pr__pnp_05v5_W0p68L0p68.model emitter base collector
.include /foss/pdks/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pnp_05v5_W0p68L0p68.model.spice
.ends

.control
dc ve 0.3 0.8 0.001
plot i(ve)
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
