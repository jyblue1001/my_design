f.end
