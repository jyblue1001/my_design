magic
tech sky130A
timestamp 1739761143
<< nwell >>
rect 800 -4355 2310 -3735
<< nmos >>
rect 900 -3645 915 -3545
rect 955 -3645 970 -3545
rect 1160 -3645 1175 -3545
rect 1215 -3645 1230 -3545
rect 1350 -3645 1365 -3545
rect 1405 -3645 1420 -3545
rect 1610 -3645 1625 -3545
rect 1665 -3645 1680 -3545
rect 1830 -3645 1845 -3545
rect 1885 -3645 1900 -3545
rect 2050 -3645 2065 -3545
rect 2215 -3645 2230 -3545
rect 900 -4545 915 -4445
rect 955 -4545 970 -4445
rect 1160 -4545 1175 -4445
rect 1215 -4545 1230 -4445
rect 1350 -4545 1365 -4445
rect 1405 -4545 1420 -4445
rect 1610 -4545 1625 -4445
rect 1665 -4545 1680 -4445
rect 1865 -4545 1880 -4445
rect 2030 -4545 2045 -4445
rect 2195 -4545 2210 -4445
<< pmos >>
rect 900 -3955 915 -3755
rect 955 -3955 970 -3755
rect 1160 -3955 1175 -3755
rect 1215 -3955 1230 -3755
rect 1350 -3955 1365 -3755
rect 1405 -3955 1420 -3755
rect 1610 -3955 1625 -3755
rect 1665 -3955 1680 -3755
rect 1830 -3955 1845 -3755
rect 1885 -3955 1900 -3755
rect 2050 -3955 2065 -3755
rect 2215 -3955 2230 -3755
rect 900 -4335 915 -4135
rect 955 -4335 970 -4135
rect 1160 -4335 1175 -4135
rect 1215 -4335 1230 -4135
rect 1350 -4335 1365 -4135
rect 1405 -4335 1420 -4135
rect 1610 -4335 1625 -4135
rect 1665 -4335 1680 -4135
rect 1865 -4335 1880 -4135
rect 2030 -4335 2045 -4135
rect 2195 -4335 2210 -4135
<< ndiff >>
rect 860 -3560 900 -3545
rect 860 -3580 870 -3560
rect 890 -3580 900 -3560
rect 860 -3610 900 -3580
rect 860 -3630 870 -3610
rect 890 -3630 900 -3610
rect 860 -3645 900 -3630
rect 915 -3560 955 -3545
rect 915 -3580 925 -3560
rect 945 -3580 955 -3560
rect 915 -3610 955 -3580
rect 915 -3630 925 -3610
rect 945 -3630 955 -3610
rect 915 -3645 955 -3630
rect 970 -3560 1010 -3545
rect 970 -3580 980 -3560
rect 1000 -3580 1010 -3560
rect 970 -3610 1010 -3580
rect 970 -3630 980 -3610
rect 1000 -3630 1010 -3610
rect 970 -3645 1010 -3630
rect 1120 -3560 1160 -3545
rect 1120 -3580 1130 -3560
rect 1150 -3580 1160 -3560
rect 1120 -3610 1160 -3580
rect 1120 -3630 1130 -3610
rect 1150 -3630 1160 -3610
rect 1120 -3645 1160 -3630
rect 1175 -3560 1215 -3545
rect 1175 -3580 1185 -3560
rect 1205 -3580 1215 -3560
rect 1175 -3610 1215 -3580
rect 1175 -3630 1185 -3610
rect 1205 -3630 1215 -3610
rect 1175 -3645 1215 -3630
rect 1230 -3560 1270 -3545
rect 1310 -3560 1350 -3545
rect 1230 -3580 1240 -3560
rect 1260 -3580 1270 -3560
rect 1310 -3580 1320 -3560
rect 1340 -3580 1350 -3560
rect 1230 -3610 1270 -3580
rect 1310 -3610 1350 -3580
rect 1230 -3630 1240 -3610
rect 1260 -3630 1270 -3610
rect 1310 -3630 1320 -3610
rect 1340 -3630 1350 -3610
rect 1230 -3645 1270 -3630
rect 1310 -3645 1350 -3630
rect 1365 -3560 1405 -3545
rect 1365 -3580 1375 -3560
rect 1395 -3580 1405 -3560
rect 1365 -3610 1405 -3580
rect 1365 -3630 1375 -3610
rect 1395 -3630 1405 -3610
rect 1365 -3645 1405 -3630
rect 1420 -3560 1460 -3545
rect 1420 -3580 1430 -3560
rect 1450 -3580 1460 -3560
rect 1420 -3610 1460 -3580
rect 1420 -3630 1430 -3610
rect 1450 -3630 1460 -3610
rect 1420 -3645 1460 -3630
rect 1570 -3560 1610 -3545
rect 1570 -3580 1580 -3560
rect 1600 -3580 1610 -3560
rect 1570 -3610 1610 -3580
rect 1570 -3630 1580 -3610
rect 1600 -3630 1610 -3610
rect 1570 -3645 1610 -3630
rect 1625 -3560 1665 -3545
rect 1625 -3580 1635 -3560
rect 1655 -3580 1665 -3560
rect 1625 -3610 1665 -3580
rect 1625 -3630 1635 -3610
rect 1655 -3630 1665 -3610
rect 1625 -3645 1665 -3630
rect 1680 -3560 1720 -3545
rect 1680 -3580 1690 -3560
rect 1710 -3580 1720 -3560
rect 1680 -3610 1720 -3580
rect 1680 -3630 1690 -3610
rect 1710 -3630 1720 -3610
rect 1680 -3645 1720 -3630
rect 1790 -3560 1830 -3545
rect 1790 -3580 1800 -3560
rect 1820 -3580 1830 -3560
rect 1790 -3610 1830 -3580
rect 1790 -3630 1800 -3610
rect 1820 -3630 1830 -3610
rect 1790 -3645 1830 -3630
rect 1845 -3560 1885 -3545
rect 1845 -3580 1855 -3560
rect 1875 -3580 1885 -3560
rect 1845 -3610 1885 -3580
rect 1845 -3630 1855 -3610
rect 1875 -3630 1885 -3610
rect 1845 -3645 1885 -3630
rect 1900 -3560 1940 -3545
rect 1900 -3580 1910 -3560
rect 1930 -3580 1940 -3560
rect 1900 -3610 1940 -3580
rect 1900 -3630 1910 -3610
rect 1930 -3630 1940 -3610
rect 1900 -3645 1940 -3630
rect 2010 -3560 2050 -3545
rect 2010 -3580 2020 -3560
rect 2040 -3580 2050 -3560
rect 2010 -3610 2050 -3580
rect 2010 -3630 2020 -3610
rect 2040 -3630 2050 -3610
rect 2010 -3645 2050 -3630
rect 2065 -3560 2105 -3545
rect 2065 -3580 2075 -3560
rect 2095 -3580 2105 -3560
rect 2065 -3610 2105 -3580
rect 2065 -3630 2075 -3610
rect 2095 -3630 2105 -3610
rect 2065 -3645 2105 -3630
rect 2175 -3560 2215 -3545
rect 2175 -3580 2185 -3560
rect 2205 -3580 2215 -3560
rect 2175 -3610 2215 -3580
rect 2175 -3630 2185 -3610
rect 2205 -3630 2215 -3610
rect 2175 -3645 2215 -3630
rect 2230 -3560 2270 -3545
rect 2230 -3580 2240 -3560
rect 2260 -3580 2270 -3560
rect 2230 -3610 2270 -3580
rect 2230 -3630 2240 -3610
rect 2260 -3630 2270 -3610
rect 2230 -3645 2270 -3630
rect 860 -4460 900 -4445
rect 860 -4480 870 -4460
rect 890 -4480 900 -4460
rect 860 -4510 900 -4480
rect 860 -4530 870 -4510
rect 890 -4530 900 -4510
rect 860 -4545 900 -4530
rect 915 -4460 955 -4445
rect 915 -4480 925 -4460
rect 945 -4480 955 -4460
rect 915 -4510 955 -4480
rect 915 -4530 925 -4510
rect 945 -4530 955 -4510
rect 915 -4545 955 -4530
rect 970 -4460 1010 -4445
rect 970 -4480 980 -4460
rect 1000 -4480 1010 -4460
rect 970 -4510 1010 -4480
rect 970 -4530 980 -4510
rect 1000 -4530 1010 -4510
rect 970 -4545 1010 -4530
rect 1120 -4460 1160 -4445
rect 1120 -4480 1130 -4460
rect 1150 -4480 1160 -4460
rect 1120 -4510 1160 -4480
rect 1120 -4530 1130 -4510
rect 1150 -4530 1160 -4510
rect 1120 -4545 1160 -4530
rect 1175 -4460 1215 -4445
rect 1175 -4480 1185 -4460
rect 1205 -4480 1215 -4460
rect 1175 -4510 1215 -4480
rect 1175 -4530 1185 -4510
rect 1205 -4530 1215 -4510
rect 1175 -4545 1215 -4530
rect 1230 -4460 1270 -4445
rect 1310 -4460 1350 -4445
rect 1230 -4480 1240 -4460
rect 1260 -4480 1270 -4460
rect 1310 -4480 1320 -4460
rect 1340 -4480 1350 -4460
rect 1230 -4510 1270 -4480
rect 1310 -4510 1350 -4480
rect 1230 -4530 1240 -4510
rect 1260 -4530 1270 -4510
rect 1310 -4530 1320 -4510
rect 1340 -4530 1350 -4510
rect 1230 -4545 1270 -4530
rect 1310 -4545 1350 -4530
rect 1365 -4460 1405 -4445
rect 1365 -4480 1375 -4460
rect 1395 -4480 1405 -4460
rect 1365 -4510 1405 -4480
rect 1365 -4530 1375 -4510
rect 1395 -4530 1405 -4510
rect 1365 -4545 1405 -4530
rect 1420 -4460 1460 -4445
rect 1420 -4480 1430 -4460
rect 1450 -4480 1460 -4460
rect 1420 -4510 1460 -4480
rect 1420 -4530 1430 -4510
rect 1450 -4530 1460 -4510
rect 1420 -4545 1460 -4530
rect 1570 -4460 1610 -4445
rect 1570 -4480 1580 -4460
rect 1600 -4480 1610 -4460
rect 1570 -4510 1610 -4480
rect 1570 -4530 1580 -4510
rect 1600 -4530 1610 -4510
rect 1570 -4545 1610 -4530
rect 1625 -4460 1665 -4445
rect 1625 -4480 1635 -4460
rect 1655 -4480 1665 -4460
rect 1625 -4510 1665 -4480
rect 1625 -4530 1635 -4510
rect 1655 -4530 1665 -4510
rect 1625 -4545 1665 -4530
rect 1680 -4460 1720 -4445
rect 1680 -4480 1690 -4460
rect 1710 -4480 1720 -4460
rect 1680 -4510 1720 -4480
rect 1680 -4530 1690 -4510
rect 1710 -4530 1720 -4510
rect 1680 -4545 1720 -4530
rect 1825 -4460 1865 -4445
rect 1825 -4480 1835 -4460
rect 1855 -4480 1865 -4460
rect 1825 -4510 1865 -4480
rect 1825 -4530 1835 -4510
rect 1855 -4530 1865 -4510
rect 1825 -4545 1865 -4530
rect 1880 -4460 1920 -4445
rect 1880 -4480 1890 -4460
rect 1910 -4480 1920 -4460
rect 1880 -4510 1920 -4480
rect 1880 -4530 1890 -4510
rect 1910 -4530 1920 -4510
rect 1880 -4545 1920 -4530
rect 1990 -4460 2030 -4445
rect 1990 -4480 2000 -4460
rect 2020 -4480 2030 -4460
rect 1990 -4510 2030 -4480
rect 1990 -4530 2000 -4510
rect 2020 -4530 2030 -4510
rect 1990 -4545 2030 -4530
rect 2045 -4460 2085 -4445
rect 2045 -4480 2055 -4460
rect 2075 -4480 2085 -4460
rect 2045 -4510 2085 -4480
rect 2045 -4530 2055 -4510
rect 2075 -4530 2085 -4510
rect 2045 -4545 2085 -4530
rect 2155 -4460 2195 -4445
rect 2155 -4480 2165 -4460
rect 2185 -4480 2195 -4460
rect 2155 -4510 2195 -4480
rect 2155 -4530 2165 -4510
rect 2185 -4530 2195 -4510
rect 2155 -4545 2195 -4530
rect 2210 -4460 2250 -4445
rect 2210 -4480 2220 -4460
rect 2240 -4480 2250 -4460
rect 2210 -4510 2250 -4480
rect 2210 -4530 2220 -4510
rect 2240 -4530 2250 -4510
rect 2210 -4545 2250 -4530
<< pdiff >>
rect 860 -3770 900 -3755
rect 860 -3790 870 -3770
rect 890 -3790 900 -3770
rect 860 -3820 900 -3790
rect 860 -3840 870 -3820
rect 890 -3840 900 -3820
rect 860 -3870 900 -3840
rect 860 -3890 870 -3870
rect 890 -3890 900 -3870
rect 860 -3920 900 -3890
rect 860 -3940 870 -3920
rect 890 -3940 900 -3920
rect 860 -3955 900 -3940
rect 915 -3770 955 -3755
rect 915 -3790 925 -3770
rect 945 -3790 955 -3770
rect 915 -3820 955 -3790
rect 915 -3840 925 -3820
rect 945 -3840 955 -3820
rect 915 -3870 955 -3840
rect 915 -3890 925 -3870
rect 945 -3890 955 -3870
rect 915 -3920 955 -3890
rect 915 -3940 925 -3920
rect 945 -3940 955 -3920
rect 915 -3955 955 -3940
rect 970 -3770 1010 -3755
rect 970 -3790 980 -3770
rect 1000 -3790 1010 -3770
rect 970 -3820 1010 -3790
rect 970 -3840 980 -3820
rect 1000 -3840 1010 -3820
rect 970 -3870 1010 -3840
rect 970 -3890 980 -3870
rect 1000 -3890 1010 -3870
rect 970 -3920 1010 -3890
rect 970 -3940 980 -3920
rect 1000 -3940 1010 -3920
rect 970 -3955 1010 -3940
rect 1120 -3770 1160 -3755
rect 1120 -3790 1130 -3770
rect 1150 -3790 1160 -3770
rect 1120 -3820 1160 -3790
rect 1120 -3840 1130 -3820
rect 1150 -3840 1160 -3820
rect 1120 -3870 1160 -3840
rect 1120 -3890 1130 -3870
rect 1150 -3890 1160 -3870
rect 1120 -3920 1160 -3890
rect 1120 -3940 1130 -3920
rect 1150 -3940 1160 -3920
rect 1120 -3955 1160 -3940
rect 1175 -3770 1215 -3755
rect 1175 -3790 1185 -3770
rect 1205 -3790 1215 -3770
rect 1175 -3820 1215 -3790
rect 1175 -3840 1185 -3820
rect 1205 -3840 1215 -3820
rect 1175 -3870 1215 -3840
rect 1175 -3890 1185 -3870
rect 1205 -3890 1215 -3870
rect 1175 -3920 1215 -3890
rect 1175 -3940 1185 -3920
rect 1205 -3940 1215 -3920
rect 1175 -3955 1215 -3940
rect 1230 -3770 1270 -3755
rect 1310 -3770 1350 -3755
rect 1230 -3790 1240 -3770
rect 1260 -3790 1270 -3770
rect 1310 -3790 1320 -3770
rect 1340 -3790 1350 -3770
rect 1230 -3820 1270 -3790
rect 1310 -3820 1350 -3790
rect 1230 -3840 1240 -3820
rect 1260 -3840 1270 -3820
rect 1310 -3840 1320 -3820
rect 1340 -3840 1350 -3820
rect 1230 -3870 1270 -3840
rect 1310 -3870 1350 -3840
rect 1230 -3890 1240 -3870
rect 1260 -3890 1270 -3870
rect 1310 -3890 1320 -3870
rect 1340 -3890 1350 -3870
rect 1230 -3920 1270 -3890
rect 1310 -3920 1350 -3890
rect 1230 -3940 1240 -3920
rect 1260 -3940 1270 -3920
rect 1310 -3940 1320 -3920
rect 1340 -3940 1350 -3920
rect 1230 -3955 1270 -3940
rect 1310 -3955 1350 -3940
rect 1365 -3770 1405 -3755
rect 1365 -3790 1375 -3770
rect 1395 -3790 1405 -3770
rect 1365 -3820 1405 -3790
rect 1365 -3840 1375 -3820
rect 1395 -3840 1405 -3820
rect 1365 -3870 1405 -3840
rect 1365 -3890 1375 -3870
rect 1395 -3890 1405 -3870
rect 1365 -3920 1405 -3890
rect 1365 -3940 1375 -3920
rect 1395 -3940 1405 -3920
rect 1365 -3955 1405 -3940
rect 1420 -3770 1460 -3755
rect 1420 -3790 1430 -3770
rect 1450 -3790 1460 -3770
rect 1420 -3820 1460 -3790
rect 1420 -3840 1430 -3820
rect 1450 -3840 1460 -3820
rect 1420 -3870 1460 -3840
rect 1420 -3890 1430 -3870
rect 1450 -3890 1460 -3870
rect 1420 -3920 1460 -3890
rect 1420 -3940 1430 -3920
rect 1450 -3940 1460 -3920
rect 1420 -3955 1460 -3940
rect 1570 -3770 1610 -3755
rect 1570 -3790 1580 -3770
rect 1600 -3790 1610 -3770
rect 1570 -3820 1610 -3790
rect 1570 -3840 1580 -3820
rect 1600 -3840 1610 -3820
rect 1570 -3870 1610 -3840
rect 1570 -3890 1580 -3870
rect 1600 -3890 1610 -3870
rect 1570 -3920 1610 -3890
rect 1570 -3940 1580 -3920
rect 1600 -3940 1610 -3920
rect 1570 -3955 1610 -3940
rect 1625 -3770 1665 -3755
rect 1625 -3790 1635 -3770
rect 1655 -3790 1665 -3770
rect 1625 -3820 1665 -3790
rect 1625 -3840 1635 -3820
rect 1655 -3840 1665 -3820
rect 1625 -3870 1665 -3840
rect 1625 -3890 1635 -3870
rect 1655 -3890 1665 -3870
rect 1625 -3920 1665 -3890
rect 1625 -3940 1635 -3920
rect 1655 -3940 1665 -3920
rect 1625 -3955 1665 -3940
rect 1680 -3770 1720 -3755
rect 1680 -3790 1690 -3770
rect 1710 -3790 1720 -3770
rect 1680 -3820 1720 -3790
rect 1680 -3840 1690 -3820
rect 1710 -3840 1720 -3820
rect 1680 -3870 1720 -3840
rect 1680 -3890 1690 -3870
rect 1710 -3890 1720 -3870
rect 1680 -3920 1720 -3890
rect 1680 -3940 1690 -3920
rect 1710 -3940 1720 -3920
rect 1680 -3955 1720 -3940
rect 1790 -3770 1830 -3755
rect 1790 -3790 1800 -3770
rect 1820 -3790 1830 -3770
rect 1790 -3820 1830 -3790
rect 1790 -3840 1800 -3820
rect 1820 -3840 1830 -3820
rect 1790 -3870 1830 -3840
rect 1790 -3890 1800 -3870
rect 1820 -3890 1830 -3870
rect 1790 -3920 1830 -3890
rect 1790 -3940 1800 -3920
rect 1820 -3940 1830 -3920
rect 1790 -3955 1830 -3940
rect 1845 -3770 1885 -3755
rect 1845 -3790 1855 -3770
rect 1875 -3790 1885 -3770
rect 1845 -3820 1885 -3790
rect 1845 -3840 1855 -3820
rect 1875 -3840 1885 -3820
rect 1845 -3870 1885 -3840
rect 1845 -3890 1855 -3870
rect 1875 -3890 1885 -3870
rect 1845 -3920 1885 -3890
rect 1845 -3940 1855 -3920
rect 1875 -3940 1885 -3920
rect 1845 -3955 1885 -3940
rect 1900 -3770 1940 -3755
rect 1900 -3790 1910 -3770
rect 1930 -3790 1940 -3770
rect 1900 -3820 1940 -3790
rect 1900 -3840 1910 -3820
rect 1930 -3840 1940 -3820
rect 1900 -3870 1940 -3840
rect 1900 -3890 1910 -3870
rect 1930 -3890 1940 -3870
rect 1900 -3920 1940 -3890
rect 1900 -3940 1910 -3920
rect 1930 -3940 1940 -3920
rect 1900 -3955 1940 -3940
rect 2010 -3770 2050 -3755
rect 2010 -3790 2020 -3770
rect 2040 -3790 2050 -3770
rect 2010 -3820 2050 -3790
rect 2010 -3840 2020 -3820
rect 2040 -3840 2050 -3820
rect 2010 -3870 2050 -3840
rect 2010 -3890 2020 -3870
rect 2040 -3890 2050 -3870
rect 2010 -3920 2050 -3890
rect 2010 -3940 2020 -3920
rect 2040 -3940 2050 -3920
rect 2010 -3955 2050 -3940
rect 2065 -3770 2105 -3755
rect 2065 -3790 2075 -3770
rect 2095 -3790 2105 -3770
rect 2065 -3820 2105 -3790
rect 2065 -3840 2075 -3820
rect 2095 -3840 2105 -3820
rect 2065 -3870 2105 -3840
rect 2065 -3890 2075 -3870
rect 2095 -3890 2105 -3870
rect 2065 -3920 2105 -3890
rect 2065 -3940 2075 -3920
rect 2095 -3940 2105 -3920
rect 2065 -3955 2105 -3940
rect 2175 -3770 2215 -3755
rect 2175 -3790 2185 -3770
rect 2205 -3790 2215 -3770
rect 2175 -3820 2215 -3790
rect 2175 -3840 2185 -3820
rect 2205 -3840 2215 -3820
rect 2175 -3870 2215 -3840
rect 2175 -3890 2185 -3870
rect 2205 -3890 2215 -3870
rect 2175 -3920 2215 -3890
rect 2175 -3940 2185 -3920
rect 2205 -3940 2215 -3920
rect 2175 -3955 2215 -3940
rect 2230 -3770 2270 -3755
rect 2230 -3790 2240 -3770
rect 2260 -3790 2270 -3770
rect 2230 -3820 2270 -3790
rect 2230 -3840 2240 -3820
rect 2260 -3840 2270 -3820
rect 2230 -3870 2270 -3840
rect 2230 -3890 2240 -3870
rect 2260 -3890 2270 -3870
rect 2230 -3920 2270 -3890
rect 2230 -3940 2240 -3920
rect 2260 -3940 2270 -3920
rect 2230 -3955 2270 -3940
rect 860 -4150 900 -4135
rect 860 -4170 870 -4150
rect 890 -4170 900 -4150
rect 860 -4200 900 -4170
rect 860 -4220 870 -4200
rect 890 -4220 900 -4200
rect 860 -4250 900 -4220
rect 860 -4270 870 -4250
rect 890 -4270 900 -4250
rect 860 -4300 900 -4270
rect 860 -4320 870 -4300
rect 890 -4320 900 -4300
rect 860 -4335 900 -4320
rect 915 -4150 955 -4135
rect 915 -4170 925 -4150
rect 945 -4170 955 -4150
rect 915 -4200 955 -4170
rect 915 -4220 925 -4200
rect 945 -4220 955 -4200
rect 915 -4250 955 -4220
rect 915 -4270 925 -4250
rect 945 -4270 955 -4250
rect 915 -4300 955 -4270
rect 915 -4320 925 -4300
rect 945 -4320 955 -4300
rect 915 -4335 955 -4320
rect 970 -4150 1010 -4135
rect 970 -4170 980 -4150
rect 1000 -4170 1010 -4150
rect 970 -4200 1010 -4170
rect 970 -4220 980 -4200
rect 1000 -4220 1010 -4200
rect 970 -4250 1010 -4220
rect 970 -4270 980 -4250
rect 1000 -4270 1010 -4250
rect 970 -4300 1010 -4270
rect 970 -4320 980 -4300
rect 1000 -4320 1010 -4300
rect 970 -4335 1010 -4320
rect 1120 -4150 1160 -4135
rect 1120 -4170 1130 -4150
rect 1150 -4170 1160 -4150
rect 1120 -4200 1160 -4170
rect 1120 -4220 1130 -4200
rect 1150 -4220 1160 -4200
rect 1120 -4250 1160 -4220
rect 1120 -4270 1130 -4250
rect 1150 -4270 1160 -4250
rect 1120 -4300 1160 -4270
rect 1120 -4320 1130 -4300
rect 1150 -4320 1160 -4300
rect 1120 -4335 1160 -4320
rect 1175 -4150 1215 -4135
rect 1175 -4170 1185 -4150
rect 1205 -4170 1215 -4150
rect 1175 -4200 1215 -4170
rect 1175 -4220 1185 -4200
rect 1205 -4220 1215 -4200
rect 1175 -4250 1215 -4220
rect 1175 -4270 1185 -4250
rect 1205 -4270 1215 -4250
rect 1175 -4300 1215 -4270
rect 1175 -4320 1185 -4300
rect 1205 -4320 1215 -4300
rect 1175 -4335 1215 -4320
rect 1230 -4150 1270 -4135
rect 1310 -4150 1350 -4135
rect 1230 -4170 1240 -4150
rect 1260 -4170 1270 -4150
rect 1310 -4170 1320 -4150
rect 1340 -4170 1350 -4150
rect 1230 -4200 1270 -4170
rect 1310 -4200 1350 -4170
rect 1230 -4220 1240 -4200
rect 1260 -4220 1270 -4200
rect 1310 -4220 1320 -4200
rect 1340 -4220 1350 -4200
rect 1230 -4250 1270 -4220
rect 1310 -4250 1350 -4220
rect 1230 -4270 1240 -4250
rect 1260 -4270 1270 -4250
rect 1310 -4270 1320 -4250
rect 1340 -4270 1350 -4250
rect 1230 -4300 1270 -4270
rect 1310 -4300 1350 -4270
rect 1230 -4320 1240 -4300
rect 1260 -4320 1270 -4300
rect 1310 -4320 1320 -4300
rect 1340 -4320 1350 -4300
rect 1230 -4335 1270 -4320
rect 1310 -4335 1350 -4320
rect 1365 -4150 1405 -4135
rect 1365 -4170 1375 -4150
rect 1395 -4170 1405 -4150
rect 1365 -4200 1405 -4170
rect 1365 -4220 1375 -4200
rect 1395 -4220 1405 -4200
rect 1365 -4250 1405 -4220
rect 1365 -4270 1375 -4250
rect 1395 -4270 1405 -4250
rect 1365 -4300 1405 -4270
rect 1365 -4320 1375 -4300
rect 1395 -4320 1405 -4300
rect 1365 -4335 1405 -4320
rect 1420 -4150 1460 -4135
rect 1420 -4170 1430 -4150
rect 1450 -4170 1460 -4150
rect 1420 -4200 1460 -4170
rect 1420 -4220 1430 -4200
rect 1450 -4220 1460 -4200
rect 1420 -4250 1460 -4220
rect 1420 -4270 1430 -4250
rect 1450 -4270 1460 -4250
rect 1420 -4300 1460 -4270
rect 1420 -4320 1430 -4300
rect 1450 -4320 1460 -4300
rect 1420 -4335 1460 -4320
rect 1570 -4150 1610 -4135
rect 1570 -4170 1580 -4150
rect 1600 -4170 1610 -4150
rect 1570 -4200 1610 -4170
rect 1570 -4220 1580 -4200
rect 1600 -4220 1610 -4200
rect 1570 -4250 1610 -4220
rect 1570 -4270 1580 -4250
rect 1600 -4270 1610 -4250
rect 1570 -4300 1610 -4270
rect 1570 -4320 1580 -4300
rect 1600 -4320 1610 -4300
rect 1570 -4335 1610 -4320
rect 1625 -4150 1665 -4135
rect 1625 -4170 1635 -4150
rect 1655 -4170 1665 -4150
rect 1625 -4200 1665 -4170
rect 1625 -4220 1635 -4200
rect 1655 -4220 1665 -4200
rect 1625 -4250 1665 -4220
rect 1625 -4270 1635 -4250
rect 1655 -4270 1665 -4250
rect 1625 -4300 1665 -4270
rect 1625 -4320 1635 -4300
rect 1655 -4320 1665 -4300
rect 1625 -4335 1665 -4320
rect 1680 -4150 1720 -4135
rect 1680 -4170 1690 -4150
rect 1710 -4170 1720 -4150
rect 1680 -4200 1720 -4170
rect 1680 -4220 1690 -4200
rect 1710 -4220 1720 -4200
rect 1680 -4250 1720 -4220
rect 1680 -4270 1690 -4250
rect 1710 -4270 1720 -4250
rect 1680 -4300 1720 -4270
rect 1680 -4320 1690 -4300
rect 1710 -4320 1720 -4300
rect 1680 -4335 1720 -4320
rect 1825 -4150 1865 -4135
rect 1825 -4170 1835 -4150
rect 1855 -4170 1865 -4150
rect 1825 -4200 1865 -4170
rect 1825 -4220 1835 -4200
rect 1855 -4220 1865 -4200
rect 1825 -4250 1865 -4220
rect 1825 -4270 1835 -4250
rect 1855 -4270 1865 -4250
rect 1825 -4300 1865 -4270
rect 1825 -4320 1835 -4300
rect 1855 -4320 1865 -4300
rect 1825 -4335 1865 -4320
rect 1880 -4150 1920 -4135
rect 1880 -4170 1890 -4150
rect 1910 -4170 1920 -4150
rect 1880 -4200 1920 -4170
rect 1880 -4220 1890 -4200
rect 1910 -4220 1920 -4200
rect 1880 -4250 1920 -4220
rect 1880 -4270 1890 -4250
rect 1910 -4270 1920 -4250
rect 1880 -4300 1920 -4270
rect 1880 -4320 1890 -4300
rect 1910 -4320 1920 -4300
rect 1880 -4335 1920 -4320
rect 1990 -4150 2030 -4135
rect 1990 -4170 2000 -4150
rect 2020 -4170 2030 -4150
rect 1990 -4200 2030 -4170
rect 1990 -4220 2000 -4200
rect 2020 -4220 2030 -4200
rect 1990 -4250 2030 -4220
rect 1990 -4270 2000 -4250
rect 2020 -4270 2030 -4250
rect 1990 -4300 2030 -4270
rect 1990 -4320 2000 -4300
rect 2020 -4320 2030 -4300
rect 1990 -4335 2030 -4320
rect 2045 -4150 2085 -4135
rect 2045 -4170 2055 -4150
rect 2075 -4170 2085 -4150
rect 2045 -4200 2085 -4170
rect 2045 -4220 2055 -4200
rect 2075 -4220 2085 -4200
rect 2045 -4250 2085 -4220
rect 2045 -4270 2055 -4250
rect 2075 -4270 2085 -4250
rect 2045 -4300 2085 -4270
rect 2045 -4320 2055 -4300
rect 2075 -4320 2085 -4300
rect 2045 -4335 2085 -4320
rect 2155 -4150 2195 -4135
rect 2155 -4170 2165 -4150
rect 2185 -4170 2195 -4150
rect 2155 -4200 2195 -4170
rect 2155 -4220 2165 -4200
rect 2185 -4220 2195 -4200
rect 2155 -4250 2195 -4220
rect 2155 -4270 2165 -4250
rect 2185 -4270 2195 -4250
rect 2155 -4300 2195 -4270
rect 2155 -4320 2165 -4300
rect 2185 -4320 2195 -4300
rect 2155 -4335 2195 -4320
rect 2210 -4150 2250 -4135
rect 2210 -4170 2220 -4150
rect 2240 -4170 2250 -4150
rect 2210 -4200 2250 -4170
rect 2210 -4220 2220 -4200
rect 2240 -4220 2250 -4200
rect 2210 -4250 2250 -4220
rect 2210 -4270 2220 -4250
rect 2240 -4270 2250 -4250
rect 2210 -4300 2250 -4270
rect 2210 -4320 2220 -4300
rect 2240 -4320 2250 -4300
rect 2210 -4335 2250 -4320
<< ndiffc >>
rect 870 -3580 890 -3560
rect 870 -3630 890 -3610
rect 925 -3580 945 -3560
rect 925 -3630 945 -3610
rect 980 -3580 1000 -3560
rect 980 -3630 1000 -3610
rect 1130 -3580 1150 -3560
rect 1130 -3630 1150 -3610
rect 1185 -3580 1205 -3560
rect 1185 -3630 1205 -3610
rect 1240 -3580 1260 -3560
rect 1320 -3580 1340 -3560
rect 1240 -3630 1260 -3610
rect 1320 -3630 1340 -3610
rect 1375 -3580 1395 -3560
rect 1375 -3630 1395 -3610
rect 1430 -3580 1450 -3560
rect 1430 -3630 1450 -3610
rect 1580 -3580 1600 -3560
rect 1580 -3630 1600 -3610
rect 1635 -3580 1655 -3560
rect 1635 -3630 1655 -3610
rect 1690 -3580 1710 -3560
rect 1690 -3630 1710 -3610
rect 1800 -3580 1820 -3560
rect 1800 -3630 1820 -3610
rect 1855 -3580 1875 -3560
rect 1855 -3630 1875 -3610
rect 1910 -3580 1930 -3560
rect 1910 -3630 1930 -3610
rect 2020 -3580 2040 -3560
rect 2020 -3630 2040 -3610
rect 2075 -3580 2095 -3560
rect 2075 -3630 2095 -3610
rect 2185 -3580 2205 -3560
rect 2185 -3630 2205 -3610
rect 2240 -3580 2260 -3560
rect 2240 -3630 2260 -3610
rect 870 -4480 890 -4460
rect 870 -4530 890 -4510
rect 925 -4480 945 -4460
rect 925 -4530 945 -4510
rect 980 -4480 1000 -4460
rect 980 -4530 1000 -4510
rect 1130 -4480 1150 -4460
rect 1130 -4530 1150 -4510
rect 1185 -4480 1205 -4460
rect 1185 -4530 1205 -4510
rect 1240 -4480 1260 -4460
rect 1320 -4480 1340 -4460
rect 1240 -4530 1260 -4510
rect 1320 -4530 1340 -4510
rect 1375 -4480 1395 -4460
rect 1375 -4530 1395 -4510
rect 1430 -4480 1450 -4460
rect 1430 -4530 1450 -4510
rect 1580 -4480 1600 -4460
rect 1580 -4530 1600 -4510
rect 1635 -4480 1655 -4460
rect 1635 -4530 1655 -4510
rect 1690 -4480 1710 -4460
rect 1690 -4530 1710 -4510
rect 1835 -4480 1855 -4460
rect 1835 -4530 1855 -4510
rect 1890 -4480 1910 -4460
rect 1890 -4530 1910 -4510
rect 2000 -4480 2020 -4460
rect 2000 -4530 2020 -4510
rect 2055 -4480 2075 -4460
rect 2055 -4530 2075 -4510
rect 2165 -4480 2185 -4460
rect 2165 -4530 2185 -4510
rect 2220 -4480 2240 -4460
rect 2220 -4530 2240 -4510
<< pdiffc >>
rect 870 -3790 890 -3770
rect 870 -3840 890 -3820
rect 870 -3890 890 -3870
rect 870 -3940 890 -3920
rect 925 -3790 945 -3770
rect 925 -3840 945 -3820
rect 925 -3890 945 -3870
rect 925 -3940 945 -3920
rect 980 -3790 1000 -3770
rect 980 -3840 1000 -3820
rect 980 -3890 1000 -3870
rect 980 -3940 1000 -3920
rect 1130 -3790 1150 -3770
rect 1130 -3840 1150 -3820
rect 1130 -3890 1150 -3870
rect 1130 -3940 1150 -3920
rect 1185 -3790 1205 -3770
rect 1185 -3840 1205 -3820
rect 1185 -3890 1205 -3870
rect 1185 -3940 1205 -3920
rect 1240 -3790 1260 -3770
rect 1320 -3790 1340 -3770
rect 1240 -3840 1260 -3820
rect 1320 -3840 1340 -3820
rect 1240 -3890 1260 -3870
rect 1320 -3890 1340 -3870
rect 1240 -3940 1260 -3920
rect 1320 -3940 1340 -3920
rect 1375 -3790 1395 -3770
rect 1375 -3840 1395 -3820
rect 1375 -3890 1395 -3870
rect 1375 -3940 1395 -3920
rect 1430 -3790 1450 -3770
rect 1430 -3840 1450 -3820
rect 1430 -3890 1450 -3870
rect 1430 -3940 1450 -3920
rect 1580 -3790 1600 -3770
rect 1580 -3840 1600 -3820
rect 1580 -3890 1600 -3870
rect 1580 -3940 1600 -3920
rect 1635 -3790 1655 -3770
rect 1635 -3840 1655 -3820
rect 1635 -3890 1655 -3870
rect 1635 -3940 1655 -3920
rect 1690 -3790 1710 -3770
rect 1690 -3840 1710 -3820
rect 1690 -3890 1710 -3870
rect 1690 -3940 1710 -3920
rect 1800 -3790 1820 -3770
rect 1800 -3840 1820 -3820
rect 1800 -3890 1820 -3870
rect 1800 -3940 1820 -3920
rect 1855 -3790 1875 -3770
rect 1855 -3840 1875 -3820
rect 1855 -3890 1875 -3870
rect 1855 -3940 1875 -3920
rect 1910 -3790 1930 -3770
rect 1910 -3840 1930 -3820
rect 1910 -3890 1930 -3870
rect 1910 -3940 1930 -3920
rect 2020 -3790 2040 -3770
rect 2020 -3840 2040 -3820
rect 2020 -3890 2040 -3870
rect 2020 -3940 2040 -3920
rect 2075 -3790 2095 -3770
rect 2075 -3840 2095 -3820
rect 2075 -3890 2095 -3870
rect 2075 -3940 2095 -3920
rect 2185 -3790 2205 -3770
rect 2185 -3840 2205 -3820
rect 2185 -3890 2205 -3870
rect 2185 -3940 2205 -3920
rect 2240 -3790 2260 -3770
rect 2240 -3840 2260 -3820
rect 2240 -3890 2260 -3870
rect 2240 -3940 2260 -3920
rect 870 -4170 890 -4150
rect 870 -4220 890 -4200
rect 870 -4270 890 -4250
rect 870 -4320 890 -4300
rect 925 -4170 945 -4150
rect 925 -4220 945 -4200
rect 925 -4270 945 -4250
rect 925 -4320 945 -4300
rect 980 -4170 1000 -4150
rect 980 -4220 1000 -4200
rect 980 -4270 1000 -4250
rect 980 -4320 1000 -4300
rect 1130 -4170 1150 -4150
rect 1130 -4220 1150 -4200
rect 1130 -4270 1150 -4250
rect 1130 -4320 1150 -4300
rect 1185 -4170 1205 -4150
rect 1185 -4220 1205 -4200
rect 1185 -4270 1205 -4250
rect 1185 -4320 1205 -4300
rect 1240 -4170 1260 -4150
rect 1320 -4170 1340 -4150
rect 1240 -4220 1260 -4200
rect 1320 -4220 1340 -4200
rect 1240 -4270 1260 -4250
rect 1320 -4270 1340 -4250
rect 1240 -4320 1260 -4300
rect 1320 -4320 1340 -4300
rect 1375 -4170 1395 -4150
rect 1375 -4220 1395 -4200
rect 1375 -4270 1395 -4250
rect 1375 -4320 1395 -4300
rect 1430 -4170 1450 -4150
rect 1430 -4220 1450 -4200
rect 1430 -4270 1450 -4250
rect 1430 -4320 1450 -4300
rect 1580 -4170 1600 -4150
rect 1580 -4220 1600 -4200
rect 1580 -4270 1600 -4250
rect 1580 -4320 1600 -4300
rect 1635 -4170 1655 -4150
rect 1635 -4220 1655 -4200
rect 1635 -4270 1655 -4250
rect 1635 -4320 1655 -4300
rect 1690 -4170 1710 -4150
rect 1690 -4220 1710 -4200
rect 1690 -4270 1710 -4250
rect 1690 -4320 1710 -4300
rect 1835 -4170 1855 -4150
rect 1835 -4220 1855 -4200
rect 1835 -4270 1855 -4250
rect 1835 -4320 1855 -4300
rect 1890 -4170 1910 -4150
rect 1890 -4220 1910 -4200
rect 1890 -4270 1910 -4250
rect 1890 -4320 1910 -4300
rect 2000 -4170 2020 -4150
rect 2000 -4220 2020 -4200
rect 2000 -4270 2020 -4250
rect 2000 -4320 2020 -4300
rect 2055 -4170 2075 -4150
rect 2055 -4220 2075 -4200
rect 2055 -4270 2075 -4250
rect 2055 -4320 2075 -4300
rect 2165 -4170 2185 -4150
rect 2165 -4220 2185 -4200
rect 2165 -4270 2185 -4250
rect 2165 -4320 2185 -4300
rect 2220 -4170 2240 -4150
rect 2220 -4220 2240 -4200
rect 2220 -4270 2240 -4250
rect 2220 -4320 2240 -4300
<< psubdiff >>
rect 820 -3560 860 -3545
rect 820 -3580 830 -3560
rect 850 -3580 860 -3560
rect 820 -3610 860 -3580
rect 820 -3630 830 -3610
rect 850 -3630 860 -3610
rect 820 -3645 860 -3630
rect 1270 -3560 1310 -3545
rect 1270 -3580 1280 -3560
rect 1300 -3580 1310 -3560
rect 1270 -3610 1310 -3580
rect 1270 -3630 1280 -3610
rect 1300 -3630 1310 -3610
rect 1270 -3645 1310 -3630
rect 1720 -3560 1760 -3545
rect 1720 -3580 1730 -3560
rect 1750 -3580 1760 -3560
rect 1720 -3610 1760 -3580
rect 1720 -3630 1730 -3610
rect 1750 -3630 1760 -3610
rect 1720 -3645 1760 -3630
rect 1970 -3560 2010 -3545
rect 1970 -3580 1980 -3560
rect 2000 -3580 2010 -3560
rect 1970 -3610 2010 -3580
rect 1970 -3630 1980 -3610
rect 2000 -3630 2010 -3610
rect 1970 -3645 2010 -3630
rect 2135 -3560 2175 -3545
rect 2135 -3580 2145 -3560
rect 2165 -3580 2175 -3560
rect 2135 -3610 2175 -3580
rect 2135 -3630 2145 -3610
rect 2165 -3630 2175 -3610
rect 2135 -3645 2175 -3630
rect 820 -4460 860 -4445
rect 820 -4480 830 -4460
rect 850 -4480 860 -4460
rect 820 -4510 860 -4480
rect 820 -4530 830 -4510
rect 850 -4530 860 -4510
rect 820 -4545 860 -4530
rect 1270 -4460 1310 -4445
rect 1270 -4480 1280 -4460
rect 1300 -4480 1310 -4460
rect 1270 -4510 1310 -4480
rect 1270 -4530 1280 -4510
rect 1300 -4530 1310 -4510
rect 1270 -4545 1310 -4530
rect 1720 -4460 1760 -4445
rect 1720 -4480 1730 -4460
rect 1750 -4480 1760 -4460
rect 1720 -4510 1760 -4480
rect 1720 -4530 1730 -4510
rect 1750 -4530 1760 -4510
rect 1720 -4545 1760 -4530
rect 1920 -4460 1960 -4445
rect 1920 -4480 1930 -4460
rect 1950 -4480 1960 -4460
rect 1920 -4510 1960 -4480
rect 1920 -4530 1930 -4510
rect 1950 -4530 1960 -4510
rect 1920 -4545 1960 -4530
rect 2085 -4460 2125 -4445
rect 2085 -4480 2095 -4460
rect 2115 -4480 2125 -4460
rect 2085 -4510 2125 -4480
rect 2085 -4530 2095 -4510
rect 2115 -4530 2125 -4510
rect 2085 -4545 2125 -4530
rect 2250 -4460 2290 -4445
rect 2250 -4480 2260 -4460
rect 2280 -4480 2290 -4460
rect 2250 -4510 2290 -4480
rect 2250 -4530 2260 -4510
rect 2280 -4530 2290 -4510
rect 2250 -4545 2290 -4530
<< nsubdiff >>
rect 820 -3770 860 -3755
rect 820 -3790 830 -3770
rect 850 -3790 860 -3770
rect 820 -3820 860 -3790
rect 820 -3840 830 -3820
rect 850 -3840 860 -3820
rect 820 -3870 860 -3840
rect 820 -3890 830 -3870
rect 850 -3890 860 -3870
rect 820 -3920 860 -3890
rect 820 -3940 830 -3920
rect 850 -3940 860 -3920
rect 820 -3955 860 -3940
rect 1270 -3770 1310 -3755
rect 1270 -3790 1280 -3770
rect 1300 -3790 1310 -3770
rect 1270 -3820 1310 -3790
rect 1270 -3840 1280 -3820
rect 1300 -3840 1310 -3820
rect 1270 -3870 1310 -3840
rect 1270 -3890 1280 -3870
rect 1300 -3890 1310 -3870
rect 1270 -3920 1310 -3890
rect 1270 -3940 1280 -3920
rect 1300 -3940 1310 -3920
rect 1270 -3955 1310 -3940
rect 1720 -3770 1760 -3755
rect 1720 -3790 1730 -3770
rect 1750 -3790 1760 -3770
rect 1720 -3820 1760 -3790
rect 1720 -3840 1730 -3820
rect 1750 -3840 1760 -3820
rect 1720 -3870 1760 -3840
rect 1720 -3890 1730 -3870
rect 1750 -3890 1760 -3870
rect 1720 -3920 1760 -3890
rect 1720 -3940 1730 -3920
rect 1750 -3940 1760 -3920
rect 1720 -3955 1760 -3940
rect 1970 -3770 2010 -3755
rect 1970 -3790 1980 -3770
rect 2000 -3790 2010 -3770
rect 1970 -3820 2010 -3790
rect 1970 -3840 1980 -3820
rect 2000 -3840 2010 -3820
rect 1970 -3870 2010 -3840
rect 1970 -3890 1980 -3870
rect 2000 -3890 2010 -3870
rect 1970 -3920 2010 -3890
rect 1970 -3940 1980 -3920
rect 2000 -3940 2010 -3920
rect 1970 -3955 2010 -3940
rect 2135 -3770 2175 -3755
rect 2135 -3790 2145 -3770
rect 2165 -3790 2175 -3770
rect 2135 -3820 2175 -3790
rect 2135 -3840 2145 -3820
rect 2165 -3840 2175 -3820
rect 2135 -3870 2175 -3840
rect 2135 -3890 2145 -3870
rect 2165 -3890 2175 -3870
rect 2135 -3920 2175 -3890
rect 2135 -3940 2145 -3920
rect 2165 -3940 2175 -3920
rect 2135 -3955 2175 -3940
rect 820 -4150 860 -4135
rect 820 -4170 830 -4150
rect 850 -4170 860 -4150
rect 820 -4200 860 -4170
rect 820 -4220 830 -4200
rect 850 -4220 860 -4200
rect 820 -4250 860 -4220
rect 820 -4270 830 -4250
rect 850 -4270 860 -4250
rect 820 -4300 860 -4270
rect 820 -4320 830 -4300
rect 850 -4320 860 -4300
rect 820 -4335 860 -4320
rect 1270 -4150 1310 -4135
rect 1270 -4170 1280 -4150
rect 1300 -4170 1310 -4150
rect 1270 -4200 1310 -4170
rect 1270 -4220 1280 -4200
rect 1300 -4220 1310 -4200
rect 1270 -4250 1310 -4220
rect 1270 -4270 1280 -4250
rect 1300 -4270 1310 -4250
rect 1270 -4300 1310 -4270
rect 1270 -4320 1280 -4300
rect 1300 -4320 1310 -4300
rect 1270 -4335 1310 -4320
rect 1720 -4150 1760 -4135
rect 1720 -4170 1730 -4150
rect 1750 -4170 1760 -4150
rect 1720 -4200 1760 -4170
rect 1720 -4220 1730 -4200
rect 1750 -4220 1760 -4200
rect 1720 -4250 1760 -4220
rect 1720 -4270 1730 -4250
rect 1750 -4270 1760 -4250
rect 1720 -4300 1760 -4270
rect 1720 -4320 1730 -4300
rect 1750 -4320 1760 -4300
rect 1720 -4335 1760 -4320
rect 1920 -4150 1960 -4135
rect 1920 -4170 1930 -4150
rect 1950 -4170 1960 -4150
rect 1920 -4200 1960 -4170
rect 1920 -4220 1930 -4200
rect 1950 -4220 1960 -4200
rect 1920 -4250 1960 -4220
rect 1920 -4270 1930 -4250
rect 1950 -4270 1960 -4250
rect 1920 -4300 1960 -4270
rect 1920 -4320 1930 -4300
rect 1950 -4320 1960 -4300
rect 1920 -4335 1960 -4320
rect 2085 -4150 2125 -4135
rect 2085 -4170 2095 -4150
rect 2115 -4170 2125 -4150
rect 2085 -4200 2125 -4170
rect 2085 -4220 2095 -4200
rect 2115 -4220 2125 -4200
rect 2085 -4250 2125 -4220
rect 2085 -4270 2095 -4250
rect 2115 -4270 2125 -4250
rect 2085 -4300 2125 -4270
rect 2085 -4320 2095 -4300
rect 2115 -4320 2125 -4300
rect 2085 -4335 2125 -4320
rect 2250 -4150 2290 -4135
rect 2250 -4170 2260 -4150
rect 2280 -4170 2290 -4150
rect 2250 -4200 2290 -4170
rect 2250 -4220 2260 -4200
rect 2280 -4220 2290 -4200
rect 2250 -4250 2290 -4220
rect 2250 -4270 2260 -4250
rect 2280 -4270 2290 -4250
rect 2250 -4300 2290 -4270
rect 2250 -4320 2260 -4300
rect 2280 -4320 2290 -4300
rect 2250 -4335 2290 -4320
<< psubdiffcont >>
rect 830 -3580 850 -3560
rect 830 -3630 850 -3610
rect 1280 -3580 1300 -3560
rect 1280 -3630 1300 -3610
rect 1730 -3580 1750 -3560
rect 1730 -3630 1750 -3610
rect 1980 -3580 2000 -3560
rect 1980 -3630 2000 -3610
rect 2145 -3580 2165 -3560
rect 2145 -3630 2165 -3610
rect 830 -4480 850 -4460
rect 830 -4530 850 -4510
rect 1280 -4480 1300 -4460
rect 1280 -4530 1300 -4510
rect 1730 -4480 1750 -4460
rect 1730 -4530 1750 -4510
rect 1930 -4480 1950 -4460
rect 1930 -4530 1950 -4510
rect 2095 -4480 2115 -4460
rect 2095 -4530 2115 -4510
rect 2260 -4480 2280 -4460
rect 2260 -4530 2280 -4510
<< nsubdiffcont >>
rect 830 -3790 850 -3770
rect 830 -3840 850 -3820
rect 830 -3890 850 -3870
rect 830 -3940 850 -3920
rect 1280 -3790 1300 -3770
rect 1280 -3840 1300 -3820
rect 1280 -3890 1300 -3870
rect 1280 -3940 1300 -3920
rect 1730 -3790 1750 -3770
rect 1730 -3840 1750 -3820
rect 1730 -3890 1750 -3870
rect 1730 -3940 1750 -3920
rect 1980 -3790 2000 -3770
rect 1980 -3840 2000 -3820
rect 1980 -3890 2000 -3870
rect 1980 -3940 2000 -3920
rect 2145 -3790 2165 -3770
rect 2145 -3840 2165 -3820
rect 2145 -3890 2165 -3870
rect 2145 -3940 2165 -3920
rect 830 -4170 850 -4150
rect 830 -4220 850 -4200
rect 830 -4270 850 -4250
rect 830 -4320 850 -4300
rect 1280 -4170 1300 -4150
rect 1280 -4220 1300 -4200
rect 1280 -4270 1300 -4250
rect 1280 -4320 1300 -4300
rect 1730 -4170 1750 -4150
rect 1730 -4220 1750 -4200
rect 1730 -4270 1750 -4250
rect 1730 -4320 1750 -4300
rect 1930 -4170 1950 -4150
rect 1930 -4220 1950 -4200
rect 1930 -4270 1950 -4250
rect 1930 -4320 1950 -4300
rect 2095 -4170 2115 -4150
rect 2095 -4220 2115 -4200
rect 2095 -4270 2115 -4250
rect 2095 -4320 2115 -4300
rect 2260 -4170 2280 -4150
rect 2260 -4220 2280 -4200
rect 2260 -4270 2280 -4250
rect 2260 -4320 2280 -4300
<< poly >>
rect 1160 -3505 1365 -3490
rect 900 -3545 915 -3530
rect 955 -3545 970 -3530
rect 1160 -3545 1175 -3505
rect 1215 -3545 1230 -3530
rect 1350 -3545 1365 -3505
rect 1885 -3500 1925 -3490
rect 1885 -3520 1895 -3500
rect 1915 -3520 1925 -3500
rect 1885 -3530 1925 -3520
rect 1405 -3545 1420 -3530
rect 1610 -3545 1625 -3530
rect 1665 -3545 1680 -3530
rect 1830 -3545 1845 -3530
rect 1885 -3545 1900 -3530
rect 2050 -3545 2065 -3530
rect 2215 -3545 2230 -3530
rect 900 -3680 915 -3645
rect 840 -3695 915 -3680
rect 900 -3755 915 -3695
rect 955 -3660 970 -3645
rect 955 -3670 1005 -3660
rect 1160 -3665 1175 -3645
rect 955 -3690 975 -3670
rect 995 -3690 1005 -3670
rect 955 -3700 1005 -3690
rect 1050 -3680 1175 -3665
rect 955 -3755 970 -3700
rect 1050 -3910 1065 -3680
rect 1160 -3755 1175 -3680
rect 1215 -3700 1230 -3645
rect 1215 -3710 1265 -3700
rect 1215 -3730 1235 -3710
rect 1255 -3730 1265 -3710
rect 1215 -3740 1265 -3730
rect 1215 -3755 1230 -3740
rect 1350 -3755 1365 -3645
rect 1405 -3660 1420 -3645
rect 1405 -3670 1455 -3660
rect 1610 -3665 1625 -3645
rect 1405 -3690 1425 -3670
rect 1445 -3690 1455 -3670
rect 1405 -3700 1455 -3690
rect 1500 -3680 1625 -3665
rect 1405 -3755 1420 -3700
rect 1025 -3920 1065 -3910
rect 1025 -3940 1035 -3920
rect 1055 -3940 1065 -3920
rect 1025 -3950 1065 -3940
rect 1500 -3910 1515 -3680
rect 1610 -3755 1625 -3680
rect 1665 -3665 1680 -3645
rect 1665 -3675 1750 -3665
rect 1665 -3680 1720 -3675
rect 1665 -3755 1680 -3680
rect 1710 -3695 1720 -3680
rect 1740 -3695 1750 -3675
rect 1710 -3705 1750 -3695
rect 1830 -3755 1845 -3645
rect 1885 -3755 1900 -3645
rect 1925 -3695 1965 -3685
rect 2050 -3695 2065 -3645
rect 1925 -3715 1935 -3695
rect 1955 -3710 2065 -3695
rect 1955 -3715 1965 -3710
rect 1925 -3725 1965 -3715
rect 2050 -3755 2065 -3710
rect 2090 -3695 2130 -3685
rect 2215 -3695 2230 -3645
rect 2090 -3715 2100 -3695
rect 2120 -3710 2230 -3695
rect 2120 -3715 2130 -3710
rect 2090 -3725 2130 -3715
rect 2215 -3755 2230 -3710
rect 2255 -3695 2295 -3685
rect 2255 -3715 2265 -3695
rect 2285 -3715 2295 -3695
rect 2255 -3725 2295 -3715
rect 1475 -3920 1515 -3910
rect 1475 -3940 1485 -3920
rect 1505 -3940 1515 -3920
rect 1475 -3950 1515 -3940
rect 900 -3970 915 -3955
rect 955 -3970 970 -3955
rect 1160 -3970 1175 -3955
rect 1215 -3970 1230 -3955
rect 1350 -3970 1365 -3955
rect 1405 -3970 1420 -3955
rect 1610 -3970 1625 -3955
rect 1665 -3970 1680 -3955
rect 1830 -3970 1845 -3955
rect 1885 -3970 1900 -3955
rect 2050 -3970 2065 -3955
rect 2215 -3970 2230 -3955
rect 1800 -3980 1845 -3970
rect 1800 -4000 1810 -3980
rect 1830 -4000 1845 -3980
rect 1800 -4010 1845 -4000
rect 900 -4135 915 -4120
rect 955 -4135 970 -4120
rect 1160 -4135 1175 -4120
rect 1215 -4135 1230 -4120
rect 1350 -4135 1365 -4120
rect 1405 -4135 1420 -4120
rect 1610 -4135 1625 -4120
rect 1665 -4135 1680 -4120
rect 1865 -4135 1880 -4120
rect 2030 -4135 2045 -4120
rect 2195 -4135 2210 -4120
rect 1025 -4150 1065 -4140
rect 1025 -4170 1035 -4150
rect 1055 -4170 1065 -4150
rect 1025 -4180 1065 -4170
rect 900 -4395 915 -4335
rect 840 -4410 915 -4395
rect 900 -4445 915 -4410
rect 955 -4390 970 -4335
rect 955 -4400 1005 -4390
rect 955 -4420 975 -4400
rect 995 -4420 1005 -4400
rect 955 -4430 1005 -4420
rect 1050 -4410 1065 -4180
rect 1475 -4150 1515 -4140
rect 1475 -4170 1485 -4150
rect 1505 -4170 1515 -4150
rect 1475 -4180 1515 -4170
rect 1160 -4410 1175 -4335
rect 1050 -4425 1175 -4410
rect 955 -4445 970 -4430
rect 1160 -4445 1175 -4425
rect 1215 -4350 1230 -4335
rect 1215 -4360 1265 -4350
rect 1215 -4380 1235 -4360
rect 1255 -4380 1265 -4360
rect 1215 -4390 1265 -4380
rect 1215 -4445 1230 -4390
rect 1350 -4445 1365 -4335
rect 1405 -4390 1420 -4335
rect 1405 -4400 1455 -4390
rect 1405 -4420 1425 -4400
rect 1445 -4420 1455 -4400
rect 1405 -4430 1455 -4420
rect 1500 -4410 1515 -4180
rect 1610 -4410 1625 -4335
rect 1500 -4425 1625 -4410
rect 1405 -4445 1420 -4430
rect 1610 -4445 1625 -4425
rect 1665 -4365 1680 -4335
rect 1665 -4375 1840 -4365
rect 1665 -4380 1730 -4375
rect 1665 -4445 1680 -4380
rect 1720 -4395 1730 -4380
rect 1750 -4380 1810 -4375
rect 1750 -4395 1760 -4380
rect 1720 -4405 1760 -4395
rect 1800 -4395 1810 -4380
rect 1830 -4395 1840 -4375
rect 1800 -4405 1840 -4395
rect 1865 -4380 1880 -4335
rect 1965 -4375 2005 -4365
rect 1965 -4380 1975 -4375
rect 1865 -4395 1975 -4380
rect 1995 -4395 2005 -4375
rect 1865 -4445 1880 -4395
rect 1965 -4405 2005 -4395
rect 2030 -4380 2045 -4335
rect 2130 -4375 2170 -4365
rect 2130 -4380 2140 -4375
rect 2030 -4395 2140 -4380
rect 2160 -4395 2170 -4375
rect 2030 -4445 2045 -4395
rect 2130 -4405 2170 -4395
rect 2195 -4380 2210 -4335
rect 2260 -4375 2300 -4365
rect 2260 -4380 2270 -4375
rect 2195 -4395 2270 -4380
rect 2290 -4395 2300 -4375
rect 2195 -4445 2210 -4395
rect 2260 -4405 2300 -4395
rect 900 -4560 915 -4545
rect 955 -4560 970 -4545
rect 1160 -4585 1175 -4545
rect 1215 -4560 1230 -4545
rect 1350 -4585 1365 -4545
rect 1405 -4560 1420 -4545
rect 1610 -4560 1625 -4545
rect 1665 -4560 1680 -4545
rect 1865 -4560 1880 -4545
rect 2030 -4560 2045 -4545
rect 2195 -4560 2210 -4545
rect 1160 -4600 1365 -4585
<< polycont >>
rect 1895 -3520 1915 -3500
rect 975 -3690 995 -3670
rect 1235 -3730 1255 -3710
rect 1425 -3690 1445 -3670
rect 1035 -3940 1055 -3920
rect 1720 -3695 1740 -3675
rect 1935 -3715 1955 -3695
rect 2100 -3715 2120 -3695
rect 2265 -3715 2285 -3695
rect 1485 -3940 1505 -3920
rect 1810 -4000 1830 -3980
rect 1035 -4170 1055 -4150
rect 975 -4420 995 -4400
rect 1485 -4170 1505 -4150
rect 1235 -4380 1255 -4360
rect 1425 -4420 1445 -4400
rect 1730 -4395 1750 -4375
rect 1810 -4395 1830 -4375
rect 1975 -4395 1995 -4375
rect 2140 -4395 2160 -4375
rect 2270 -4395 2290 -4375
<< locali >>
rect 650 -3445 700 -3435
rect 650 -3450 730 -3445
rect 650 -3470 665 -3450
rect 685 -3465 730 -3450
rect 750 -3465 780 -3445
rect 800 -3465 830 -3445
rect 850 -3465 880 -3445
rect 900 -3465 930 -3445
rect 950 -3465 980 -3445
rect 1000 -3465 1030 -3445
rect 1050 -3465 1080 -3445
rect 1100 -3465 1130 -3445
rect 1150 -3465 1180 -3445
rect 1200 -3465 1230 -3445
rect 1250 -3465 1280 -3445
rect 1300 -3465 1330 -3445
rect 1350 -3465 1380 -3445
rect 1400 -3465 1430 -3445
rect 1450 -3465 1480 -3445
rect 1500 -3465 1530 -3445
rect 1550 -3465 1580 -3445
rect 1600 -3465 1630 -3445
rect 1650 -3465 1680 -3445
rect 1700 -3465 1730 -3445
rect 1750 -3465 1780 -3445
rect 1800 -3465 1830 -3445
rect 1850 -3465 1880 -3445
rect 1900 -3465 1930 -3445
rect 1950 -3465 1980 -3445
rect 2000 -3465 2030 -3445
rect 2050 -3465 2080 -3445
rect 2100 -3465 2130 -3445
rect 2150 -3465 2180 -3445
rect 2200 -3465 2230 -3445
rect 2250 -3465 2280 -3445
rect 2300 -3465 2310 -3445
rect 685 -3470 700 -3465
rect 650 -3485 700 -3470
rect 870 -3550 890 -3465
rect 980 -3550 1000 -3465
rect 1065 -3500 1105 -3490
rect 1065 -3520 1075 -3500
rect 1095 -3520 1105 -3500
rect 1065 -3530 1105 -3520
rect 825 -3560 895 -3550
rect 825 -3580 830 -3560
rect 850 -3580 870 -3560
rect 890 -3580 895 -3560
rect 825 -3610 895 -3580
rect 825 -3630 830 -3610
rect 850 -3630 870 -3610
rect 890 -3630 895 -3610
rect 825 -3640 895 -3630
rect 920 -3560 950 -3550
rect 920 -3580 925 -3560
rect 945 -3580 950 -3560
rect 920 -3610 950 -3580
rect 920 -3630 925 -3610
rect 945 -3630 950 -3610
rect 920 -3640 950 -3630
rect 975 -3560 1005 -3550
rect 975 -3580 980 -3560
rect 1000 -3580 1005 -3560
rect 975 -3610 1005 -3580
rect 975 -3630 980 -3610
rect 1000 -3630 1005 -3610
rect 975 -3640 1005 -3630
rect 920 -3720 940 -3640
rect 965 -3670 1005 -3660
rect 965 -3690 975 -3670
rect 995 -3680 1005 -3670
rect 1085 -3680 1105 -3530
rect 1130 -3550 1150 -3465
rect 1240 -3550 1260 -3465
rect 1320 -3550 1340 -3465
rect 1430 -3550 1450 -3465
rect 1580 -3550 1600 -3465
rect 1690 -3550 1710 -3465
rect 1800 -3550 1820 -3465
rect 1885 -3500 1925 -3490
rect 1885 -3520 1895 -3500
rect 1915 -3520 1925 -3500
rect 1885 -3530 1925 -3520
rect 2020 -3550 2040 -3465
rect 2185 -3550 2205 -3465
rect 1125 -3560 1155 -3550
rect 1125 -3580 1130 -3560
rect 1150 -3580 1155 -3560
rect 1125 -3610 1155 -3580
rect 1125 -3630 1130 -3610
rect 1150 -3630 1155 -3610
rect 1125 -3640 1155 -3630
rect 1180 -3560 1210 -3550
rect 1180 -3580 1185 -3560
rect 1205 -3580 1210 -3560
rect 1180 -3610 1210 -3580
rect 1180 -3630 1185 -3610
rect 1205 -3630 1210 -3610
rect 1180 -3640 1210 -3630
rect 1235 -3560 1345 -3550
rect 1235 -3580 1240 -3560
rect 1260 -3580 1280 -3560
rect 1300 -3580 1320 -3560
rect 1340 -3580 1345 -3560
rect 1235 -3610 1345 -3580
rect 1235 -3630 1240 -3610
rect 1260 -3630 1280 -3610
rect 1300 -3630 1320 -3610
rect 1340 -3630 1345 -3610
rect 1235 -3640 1345 -3630
rect 1370 -3560 1400 -3550
rect 1370 -3580 1375 -3560
rect 1395 -3580 1400 -3560
rect 1370 -3610 1400 -3580
rect 1370 -3630 1375 -3610
rect 1395 -3630 1400 -3610
rect 1370 -3640 1400 -3630
rect 1425 -3560 1455 -3550
rect 1425 -3580 1430 -3560
rect 1450 -3580 1455 -3560
rect 1425 -3610 1455 -3580
rect 1425 -3630 1430 -3610
rect 1450 -3630 1455 -3610
rect 1425 -3640 1455 -3630
rect 1575 -3560 1605 -3550
rect 1575 -3580 1580 -3560
rect 1600 -3580 1605 -3560
rect 1575 -3610 1605 -3580
rect 1575 -3630 1580 -3610
rect 1600 -3630 1605 -3610
rect 1575 -3640 1605 -3630
rect 1630 -3560 1660 -3550
rect 1630 -3580 1635 -3560
rect 1655 -3580 1660 -3560
rect 1630 -3610 1660 -3580
rect 1630 -3630 1635 -3610
rect 1655 -3630 1660 -3610
rect 1630 -3640 1660 -3630
rect 1685 -3560 1755 -3550
rect 1685 -3580 1690 -3560
rect 1710 -3580 1730 -3560
rect 1750 -3580 1755 -3560
rect 1685 -3610 1755 -3580
rect 1685 -3630 1690 -3610
rect 1710 -3630 1730 -3610
rect 1750 -3630 1755 -3610
rect 1685 -3640 1755 -3630
rect 1795 -3560 1825 -3550
rect 1795 -3580 1800 -3560
rect 1820 -3580 1825 -3560
rect 1795 -3610 1825 -3580
rect 1795 -3630 1800 -3610
rect 1820 -3630 1825 -3610
rect 1795 -3640 1825 -3630
rect 1850 -3560 1880 -3550
rect 1850 -3580 1855 -3560
rect 1875 -3580 1880 -3560
rect 1850 -3610 1880 -3580
rect 1850 -3630 1855 -3610
rect 1875 -3630 1880 -3610
rect 1850 -3640 1880 -3630
rect 1905 -3560 1935 -3550
rect 1905 -3580 1910 -3560
rect 1930 -3580 1935 -3560
rect 1905 -3610 1935 -3580
rect 1905 -3630 1910 -3610
rect 1930 -3630 1935 -3610
rect 1905 -3640 1935 -3630
rect 1975 -3560 2045 -3550
rect 1975 -3580 1980 -3560
rect 2000 -3580 2020 -3560
rect 2040 -3580 2045 -3560
rect 1975 -3610 2045 -3580
rect 1975 -3630 1980 -3610
rect 2000 -3630 2020 -3610
rect 2040 -3630 2045 -3610
rect 1975 -3640 2045 -3630
rect 2070 -3560 2100 -3550
rect 2070 -3580 2075 -3560
rect 2095 -3580 2100 -3560
rect 2070 -3610 2100 -3580
rect 2070 -3630 2075 -3610
rect 2095 -3630 2100 -3610
rect 2070 -3640 2100 -3630
rect 2140 -3560 2210 -3550
rect 2140 -3580 2145 -3560
rect 2165 -3580 2185 -3560
rect 2205 -3580 2210 -3560
rect 2140 -3610 2210 -3580
rect 2140 -3630 2145 -3610
rect 2165 -3630 2185 -3610
rect 2205 -3630 2210 -3610
rect 2140 -3640 2210 -3630
rect 2235 -3560 2265 -3550
rect 2235 -3580 2240 -3560
rect 2260 -3580 2265 -3560
rect 2235 -3610 2265 -3580
rect 2235 -3630 2240 -3610
rect 2260 -3630 2265 -3610
rect 2235 -3640 2265 -3630
rect 995 -3690 1105 -3680
rect 965 -3700 1105 -3690
rect 920 -3740 1000 -3720
rect 980 -3760 1000 -3740
rect 825 -3770 895 -3760
rect 825 -3790 830 -3770
rect 850 -3790 870 -3770
rect 890 -3790 895 -3770
rect 825 -3820 895 -3790
rect 825 -3840 830 -3820
rect 850 -3840 870 -3820
rect 890 -3840 895 -3820
rect 825 -3870 895 -3840
rect 825 -3890 830 -3870
rect 850 -3890 870 -3870
rect 890 -3890 895 -3870
rect 825 -3920 895 -3890
rect 825 -3940 830 -3920
rect 850 -3940 870 -3920
rect 890 -3940 895 -3920
rect 825 -3950 895 -3940
rect 920 -3770 950 -3760
rect 920 -3790 925 -3770
rect 945 -3790 950 -3770
rect 920 -3820 950 -3790
rect 920 -3840 925 -3820
rect 945 -3840 950 -3820
rect 920 -3870 950 -3840
rect 920 -3890 925 -3870
rect 945 -3890 950 -3870
rect 920 -3920 950 -3890
rect 920 -3940 925 -3920
rect 945 -3940 950 -3920
rect 920 -3950 950 -3940
rect 975 -3770 1005 -3760
rect 975 -3790 980 -3770
rect 1000 -3790 1005 -3770
rect 975 -3820 1005 -3790
rect 975 -3840 980 -3820
rect 1000 -3840 1005 -3820
rect 975 -3870 1005 -3840
rect 975 -3890 980 -3870
rect 1000 -3890 1005 -3870
rect 975 -3920 1005 -3890
rect 975 -3940 980 -3920
rect 1000 -3925 1005 -3920
rect 1025 -3920 1065 -3910
rect 1025 -3925 1035 -3920
rect 1000 -3940 1035 -3925
rect 1055 -3940 1065 -3920
rect 975 -3950 1065 -3940
rect 1085 -3930 1105 -3700
rect 1185 -3720 1205 -3640
rect 1130 -3740 1205 -3720
rect 1225 -3710 1265 -3700
rect 1225 -3730 1235 -3710
rect 1255 -3720 1265 -3710
rect 1370 -3720 1390 -3640
rect 1415 -3670 1455 -3660
rect 1415 -3690 1425 -3670
rect 1445 -3680 1455 -3670
rect 1445 -3690 1555 -3680
rect 1415 -3700 1555 -3690
rect 1255 -3730 1450 -3720
rect 1225 -3740 1450 -3730
rect 1130 -3760 1150 -3740
rect 1430 -3760 1450 -3740
rect 1125 -3770 1155 -3760
rect 1125 -3790 1130 -3770
rect 1150 -3790 1155 -3770
rect 1125 -3820 1155 -3790
rect 1125 -3840 1130 -3820
rect 1150 -3840 1155 -3820
rect 1125 -3870 1155 -3840
rect 1125 -3890 1130 -3870
rect 1150 -3890 1155 -3870
rect 1125 -3920 1155 -3890
rect 1125 -3930 1130 -3920
rect 1085 -3940 1130 -3930
rect 1150 -3940 1155 -3920
rect 1085 -3950 1155 -3940
rect 1180 -3770 1210 -3760
rect 1180 -3790 1185 -3770
rect 1205 -3790 1210 -3770
rect 1180 -3820 1210 -3790
rect 1180 -3840 1185 -3820
rect 1205 -3840 1210 -3820
rect 1180 -3870 1210 -3840
rect 1180 -3890 1185 -3870
rect 1205 -3890 1210 -3870
rect 1180 -3920 1210 -3890
rect 1180 -3940 1185 -3920
rect 1205 -3940 1210 -3920
rect 1180 -3950 1210 -3940
rect 1235 -3770 1345 -3760
rect 1235 -3790 1240 -3770
rect 1260 -3790 1280 -3770
rect 1300 -3790 1320 -3770
rect 1340 -3790 1345 -3770
rect 1235 -3820 1345 -3790
rect 1235 -3840 1240 -3820
rect 1260 -3840 1280 -3820
rect 1300 -3840 1320 -3820
rect 1340 -3840 1345 -3820
rect 1235 -3870 1345 -3840
rect 1235 -3890 1240 -3870
rect 1260 -3890 1280 -3870
rect 1300 -3890 1320 -3870
rect 1340 -3890 1345 -3870
rect 1235 -3920 1345 -3890
rect 1235 -3940 1240 -3920
rect 1260 -3940 1280 -3920
rect 1300 -3940 1320 -3920
rect 1340 -3940 1345 -3920
rect 1235 -3950 1345 -3940
rect 1370 -3770 1400 -3760
rect 1370 -3790 1375 -3770
rect 1395 -3790 1400 -3770
rect 1370 -3820 1400 -3790
rect 1370 -3840 1375 -3820
rect 1395 -3840 1400 -3820
rect 1370 -3870 1400 -3840
rect 1370 -3890 1375 -3870
rect 1395 -3890 1400 -3870
rect 1370 -3920 1400 -3890
rect 1370 -3940 1375 -3920
rect 1395 -3940 1400 -3920
rect 1370 -3950 1400 -3940
rect 1425 -3770 1455 -3760
rect 1425 -3790 1430 -3770
rect 1450 -3790 1455 -3770
rect 1425 -3820 1455 -3790
rect 1425 -3840 1430 -3820
rect 1450 -3840 1455 -3820
rect 1425 -3870 1455 -3840
rect 1425 -3890 1430 -3870
rect 1450 -3890 1455 -3870
rect 1425 -3920 1455 -3890
rect 1425 -3940 1430 -3920
rect 1450 -3925 1455 -3920
rect 1475 -3920 1515 -3910
rect 1475 -3925 1485 -3920
rect 1450 -3940 1485 -3925
rect 1505 -3940 1515 -3920
rect 1425 -3950 1515 -3940
rect 1535 -3930 1555 -3700
rect 1635 -3720 1655 -3640
rect 1710 -3675 1750 -3665
rect 1710 -3695 1720 -3675
rect 1740 -3695 1750 -3675
rect 1710 -3705 1750 -3695
rect 1910 -3685 1930 -3640
rect 2080 -3685 2100 -3640
rect 2245 -3685 2265 -3640
rect 1910 -3695 1965 -3685
rect 1910 -3715 1935 -3695
rect 1955 -3715 1965 -3695
rect 1910 -3720 1965 -3715
rect 1580 -3740 1655 -3720
rect 1800 -3725 1965 -3720
rect 2080 -3695 2130 -3685
rect 2080 -3715 2100 -3695
rect 2120 -3715 2130 -3695
rect 2080 -3725 2130 -3715
rect 2245 -3695 2295 -3685
rect 2245 -3715 2265 -3695
rect 2285 -3715 2295 -3695
rect 2245 -3725 2295 -3715
rect 1800 -3740 1930 -3725
rect 1580 -3760 1600 -3740
rect 1800 -3760 1820 -3740
rect 1910 -3760 1930 -3740
rect 2080 -3760 2100 -3725
rect 2245 -3760 2265 -3725
rect 1575 -3770 1605 -3760
rect 1575 -3790 1580 -3770
rect 1600 -3790 1605 -3770
rect 1575 -3820 1605 -3790
rect 1575 -3840 1580 -3820
rect 1600 -3840 1605 -3820
rect 1575 -3870 1605 -3840
rect 1575 -3890 1580 -3870
rect 1600 -3890 1605 -3870
rect 1575 -3920 1605 -3890
rect 1575 -3930 1580 -3920
rect 1535 -3940 1580 -3930
rect 1600 -3940 1605 -3920
rect 1535 -3950 1605 -3940
rect 1630 -3770 1660 -3760
rect 1630 -3790 1635 -3770
rect 1655 -3790 1660 -3770
rect 1630 -3820 1660 -3790
rect 1630 -3840 1635 -3820
rect 1655 -3840 1660 -3820
rect 1630 -3870 1660 -3840
rect 1630 -3890 1635 -3870
rect 1655 -3890 1660 -3870
rect 1630 -3920 1660 -3890
rect 1630 -3940 1635 -3920
rect 1655 -3940 1660 -3920
rect 1630 -3950 1660 -3940
rect 1685 -3770 1755 -3760
rect 1685 -3790 1690 -3770
rect 1710 -3790 1730 -3770
rect 1750 -3790 1755 -3770
rect 1685 -3820 1755 -3790
rect 1685 -3840 1690 -3820
rect 1710 -3840 1730 -3820
rect 1750 -3840 1755 -3820
rect 1685 -3870 1755 -3840
rect 1685 -3890 1690 -3870
rect 1710 -3890 1730 -3870
rect 1750 -3890 1755 -3870
rect 1685 -3920 1755 -3890
rect 1685 -3940 1690 -3920
rect 1710 -3940 1730 -3920
rect 1750 -3940 1755 -3920
rect 1685 -3950 1755 -3940
rect 1795 -3770 1825 -3760
rect 1795 -3790 1800 -3770
rect 1820 -3790 1825 -3770
rect 1795 -3820 1825 -3790
rect 1795 -3840 1800 -3820
rect 1820 -3840 1825 -3820
rect 1795 -3870 1825 -3840
rect 1795 -3890 1800 -3870
rect 1820 -3890 1825 -3870
rect 1795 -3920 1825 -3890
rect 1795 -3940 1800 -3920
rect 1820 -3940 1825 -3920
rect 1795 -3950 1825 -3940
rect 1850 -3770 1880 -3760
rect 1850 -3790 1855 -3770
rect 1875 -3790 1880 -3770
rect 1850 -3820 1880 -3790
rect 1850 -3840 1855 -3820
rect 1875 -3840 1880 -3820
rect 1850 -3870 1880 -3840
rect 1850 -3890 1855 -3870
rect 1875 -3890 1880 -3870
rect 1850 -3920 1880 -3890
rect 1850 -3940 1855 -3920
rect 1875 -3940 1880 -3920
rect 1850 -3950 1880 -3940
rect 1905 -3770 1935 -3760
rect 1905 -3790 1910 -3770
rect 1930 -3790 1935 -3770
rect 1905 -3820 1935 -3790
rect 1905 -3840 1910 -3820
rect 1930 -3840 1935 -3820
rect 1905 -3870 1935 -3840
rect 1905 -3890 1910 -3870
rect 1930 -3890 1935 -3870
rect 1905 -3920 1935 -3890
rect 1905 -3940 1910 -3920
rect 1930 -3940 1935 -3920
rect 1905 -3950 1935 -3940
rect 1975 -3770 2045 -3760
rect 1975 -3790 1980 -3770
rect 2000 -3790 2020 -3770
rect 2040 -3790 2045 -3770
rect 1975 -3820 2045 -3790
rect 1975 -3840 1980 -3820
rect 2000 -3840 2020 -3820
rect 2040 -3840 2045 -3820
rect 1975 -3870 2045 -3840
rect 1975 -3890 1980 -3870
rect 2000 -3890 2020 -3870
rect 2040 -3890 2045 -3870
rect 1975 -3920 2045 -3890
rect 1975 -3940 1980 -3920
rect 2000 -3940 2020 -3920
rect 2040 -3940 2045 -3920
rect 1975 -3950 2045 -3940
rect 2070 -3770 2100 -3760
rect 2070 -3790 2075 -3770
rect 2095 -3790 2100 -3770
rect 2070 -3820 2100 -3790
rect 2070 -3840 2075 -3820
rect 2095 -3840 2100 -3820
rect 2070 -3870 2100 -3840
rect 2070 -3890 2075 -3870
rect 2095 -3890 2100 -3870
rect 2070 -3920 2100 -3890
rect 2070 -3940 2075 -3920
rect 2095 -3940 2100 -3920
rect 2070 -3950 2100 -3940
rect 2140 -3770 2210 -3760
rect 2140 -3790 2145 -3770
rect 2165 -3790 2185 -3770
rect 2205 -3790 2210 -3770
rect 2140 -3820 2210 -3790
rect 2140 -3840 2145 -3820
rect 2165 -3840 2185 -3820
rect 2205 -3840 2210 -3820
rect 2140 -3870 2210 -3840
rect 2140 -3890 2145 -3870
rect 2165 -3890 2185 -3870
rect 2205 -3890 2210 -3870
rect 2140 -3920 2210 -3890
rect 2140 -3940 2145 -3920
rect 2165 -3940 2185 -3920
rect 2205 -3940 2210 -3920
rect 2140 -3950 2210 -3940
rect 2235 -3770 2265 -3760
rect 2235 -3790 2240 -3770
rect 2260 -3790 2265 -3770
rect 2235 -3820 2265 -3790
rect 2235 -3840 2240 -3820
rect 2260 -3840 2265 -3820
rect 2235 -3870 2265 -3840
rect 2235 -3890 2240 -3870
rect 2260 -3890 2265 -3870
rect 2235 -3920 2265 -3890
rect 2235 -3940 2240 -3920
rect 2260 -3940 2265 -3920
rect 2235 -3950 2265 -3940
rect 870 -4035 890 -3950
rect 1240 -4035 1260 -3950
rect 1320 -4035 1340 -3950
rect 1690 -4035 1710 -3950
rect 1800 -3980 1840 -3970
rect 1800 -4000 1810 -3980
rect 1830 -4000 1840 -3980
rect 1800 -4010 1840 -4000
rect 1860 -4035 1880 -3950
rect 2020 -4035 2040 -3950
rect 2185 -4035 2205 -3950
rect 800 -4055 830 -4035
rect 850 -4055 880 -4035
rect 900 -4055 930 -4035
rect 950 -4055 980 -4035
rect 1000 -4055 1030 -4035
rect 1050 -4055 1080 -4035
rect 1100 -4055 1130 -4035
rect 1150 -4055 1180 -4035
rect 1200 -4055 1230 -4035
rect 1250 -4055 1280 -4035
rect 1300 -4055 1330 -4035
rect 1350 -4055 1380 -4035
rect 1400 -4055 1430 -4035
rect 1450 -4055 1480 -4035
rect 1500 -4055 1530 -4035
rect 1550 -4055 1580 -4035
rect 1600 -4055 1630 -4035
rect 1650 -4055 1680 -4035
rect 1700 -4055 1730 -4035
rect 1750 -4055 1780 -4035
rect 1800 -4055 1830 -4035
rect 1850 -4055 1880 -4035
rect 1900 -4055 1930 -4035
rect 1950 -4055 1980 -4035
rect 2000 -4055 2030 -4035
rect 2050 -4055 2080 -4035
rect 2100 -4055 2130 -4035
rect 2150 -4055 2180 -4035
rect 2200 -4055 2230 -4035
rect 2250 -4055 2280 -4035
rect 2300 -4055 2310 -4035
rect 870 -4140 890 -4055
rect 1085 -4090 1125 -4080
rect 1085 -4110 1095 -4090
rect 1115 -4110 1125 -4090
rect 1085 -4120 1125 -4110
rect 1085 -4140 1105 -4120
rect 1240 -4140 1260 -4055
rect 1320 -4140 1340 -4055
rect 1690 -4140 1710 -4055
rect 1890 -4140 1910 -4055
rect 2055 -4140 2075 -4055
rect 2220 -4140 2240 -4055
rect 825 -4150 895 -4140
rect 825 -4170 830 -4150
rect 850 -4170 870 -4150
rect 890 -4170 895 -4150
rect 825 -4200 895 -4170
rect 825 -4220 830 -4200
rect 850 -4220 870 -4200
rect 890 -4220 895 -4200
rect 825 -4250 895 -4220
rect 825 -4270 830 -4250
rect 850 -4270 870 -4250
rect 890 -4270 895 -4250
rect 825 -4300 895 -4270
rect 825 -4320 830 -4300
rect 850 -4320 870 -4300
rect 890 -4320 895 -4300
rect 825 -4330 895 -4320
rect 920 -4150 950 -4140
rect 920 -4170 925 -4150
rect 945 -4170 950 -4150
rect 920 -4200 950 -4170
rect 920 -4220 925 -4200
rect 945 -4220 950 -4200
rect 920 -4250 950 -4220
rect 920 -4270 925 -4250
rect 945 -4270 950 -4250
rect 920 -4300 950 -4270
rect 920 -4320 925 -4300
rect 945 -4320 950 -4300
rect 920 -4330 950 -4320
rect 975 -4150 1065 -4140
rect 975 -4170 980 -4150
rect 1000 -4165 1035 -4150
rect 1000 -4170 1005 -4165
rect 975 -4200 1005 -4170
rect 1025 -4170 1035 -4165
rect 1055 -4170 1065 -4150
rect 1025 -4180 1065 -4170
rect 1085 -4150 1155 -4140
rect 1085 -4160 1130 -4150
rect 975 -4220 980 -4200
rect 1000 -4220 1005 -4200
rect 975 -4250 1005 -4220
rect 975 -4270 980 -4250
rect 1000 -4270 1005 -4250
rect 975 -4300 1005 -4270
rect 975 -4320 980 -4300
rect 1000 -4320 1005 -4300
rect 975 -4330 1005 -4320
rect 980 -4350 1000 -4330
rect 920 -4370 1000 -4350
rect 920 -4450 940 -4370
rect 1085 -4390 1105 -4160
rect 1125 -4170 1130 -4160
rect 1150 -4170 1155 -4150
rect 1125 -4200 1155 -4170
rect 1125 -4220 1130 -4200
rect 1150 -4220 1155 -4200
rect 1125 -4250 1155 -4220
rect 1125 -4270 1130 -4250
rect 1150 -4270 1155 -4250
rect 1125 -4300 1155 -4270
rect 1125 -4320 1130 -4300
rect 1150 -4320 1155 -4300
rect 1125 -4330 1155 -4320
rect 1180 -4150 1210 -4140
rect 1180 -4170 1185 -4150
rect 1205 -4170 1210 -4150
rect 1180 -4200 1210 -4170
rect 1180 -4220 1185 -4200
rect 1205 -4220 1210 -4200
rect 1180 -4250 1210 -4220
rect 1180 -4270 1185 -4250
rect 1205 -4270 1210 -4250
rect 1180 -4300 1210 -4270
rect 1180 -4320 1185 -4300
rect 1205 -4320 1210 -4300
rect 1180 -4330 1210 -4320
rect 1235 -4150 1345 -4140
rect 1235 -4170 1240 -4150
rect 1260 -4170 1280 -4150
rect 1300 -4170 1320 -4150
rect 1340 -4170 1345 -4150
rect 1235 -4200 1345 -4170
rect 1235 -4220 1240 -4200
rect 1260 -4220 1280 -4200
rect 1300 -4220 1320 -4200
rect 1340 -4220 1345 -4200
rect 1235 -4250 1345 -4220
rect 1235 -4270 1240 -4250
rect 1260 -4270 1280 -4250
rect 1300 -4270 1320 -4250
rect 1340 -4270 1345 -4250
rect 1235 -4300 1345 -4270
rect 1235 -4320 1240 -4300
rect 1260 -4320 1280 -4300
rect 1300 -4320 1320 -4300
rect 1340 -4320 1345 -4300
rect 1235 -4330 1345 -4320
rect 1370 -4150 1400 -4140
rect 1370 -4170 1375 -4150
rect 1395 -4170 1400 -4150
rect 1370 -4200 1400 -4170
rect 1370 -4220 1375 -4200
rect 1395 -4220 1400 -4200
rect 1370 -4250 1400 -4220
rect 1370 -4270 1375 -4250
rect 1395 -4270 1400 -4250
rect 1370 -4300 1400 -4270
rect 1370 -4320 1375 -4300
rect 1395 -4320 1400 -4300
rect 1370 -4330 1400 -4320
rect 1425 -4150 1515 -4140
rect 1425 -4170 1430 -4150
rect 1450 -4165 1485 -4150
rect 1450 -4170 1455 -4165
rect 1425 -4200 1455 -4170
rect 1475 -4170 1485 -4165
rect 1505 -4170 1515 -4150
rect 1475 -4180 1515 -4170
rect 1535 -4150 1605 -4140
rect 1535 -4160 1580 -4150
rect 1425 -4220 1430 -4200
rect 1450 -4220 1455 -4200
rect 1425 -4250 1455 -4220
rect 1425 -4270 1430 -4250
rect 1450 -4270 1455 -4250
rect 1425 -4300 1455 -4270
rect 1425 -4320 1430 -4300
rect 1450 -4320 1455 -4300
rect 1425 -4330 1455 -4320
rect 1130 -4350 1150 -4330
rect 1430 -4350 1450 -4330
rect 1130 -4370 1205 -4350
rect 965 -4400 1105 -4390
rect 965 -4420 975 -4400
rect 995 -4410 1105 -4400
rect 995 -4420 1005 -4410
rect 965 -4430 1005 -4420
rect 1185 -4450 1205 -4370
rect 1225 -4360 1450 -4350
rect 1225 -4380 1235 -4360
rect 1255 -4370 1450 -4360
rect 1255 -4380 1265 -4370
rect 1225 -4390 1265 -4380
rect 1370 -4450 1390 -4370
rect 1535 -4390 1555 -4160
rect 1575 -4170 1580 -4160
rect 1600 -4170 1605 -4150
rect 1575 -4200 1605 -4170
rect 1575 -4220 1580 -4200
rect 1600 -4220 1605 -4200
rect 1575 -4250 1605 -4220
rect 1575 -4270 1580 -4250
rect 1600 -4270 1605 -4250
rect 1575 -4300 1605 -4270
rect 1575 -4320 1580 -4300
rect 1600 -4320 1605 -4300
rect 1575 -4330 1605 -4320
rect 1630 -4150 1660 -4140
rect 1630 -4170 1635 -4150
rect 1655 -4170 1660 -4150
rect 1630 -4200 1660 -4170
rect 1630 -4220 1635 -4200
rect 1655 -4220 1660 -4200
rect 1630 -4250 1660 -4220
rect 1630 -4270 1635 -4250
rect 1655 -4270 1660 -4250
rect 1630 -4300 1660 -4270
rect 1630 -4320 1635 -4300
rect 1655 -4320 1660 -4300
rect 1630 -4330 1660 -4320
rect 1685 -4150 1755 -4140
rect 1685 -4170 1690 -4150
rect 1710 -4170 1730 -4150
rect 1750 -4170 1755 -4150
rect 1685 -4200 1755 -4170
rect 1685 -4220 1690 -4200
rect 1710 -4220 1730 -4200
rect 1750 -4220 1755 -4200
rect 1685 -4250 1755 -4220
rect 1685 -4270 1690 -4250
rect 1710 -4270 1730 -4250
rect 1750 -4270 1755 -4250
rect 1685 -4300 1755 -4270
rect 1685 -4320 1690 -4300
rect 1710 -4320 1730 -4300
rect 1750 -4320 1755 -4300
rect 1685 -4330 1755 -4320
rect 1830 -4150 1860 -4140
rect 1830 -4170 1835 -4150
rect 1855 -4170 1860 -4150
rect 1830 -4200 1860 -4170
rect 1830 -4220 1835 -4200
rect 1855 -4220 1860 -4200
rect 1830 -4250 1860 -4220
rect 1830 -4270 1835 -4250
rect 1855 -4270 1860 -4250
rect 1830 -4300 1860 -4270
rect 1830 -4320 1835 -4300
rect 1855 -4320 1860 -4300
rect 1830 -4330 1860 -4320
rect 1885 -4150 1955 -4140
rect 1885 -4170 1890 -4150
rect 1910 -4170 1930 -4150
rect 1950 -4170 1955 -4150
rect 1885 -4200 1955 -4170
rect 1885 -4220 1890 -4200
rect 1910 -4220 1930 -4200
rect 1950 -4220 1955 -4200
rect 1885 -4250 1955 -4220
rect 1885 -4270 1890 -4250
rect 1910 -4270 1930 -4250
rect 1950 -4270 1955 -4250
rect 1885 -4300 1955 -4270
rect 1885 -4320 1890 -4300
rect 1910 -4320 1930 -4300
rect 1950 -4320 1955 -4300
rect 1885 -4330 1955 -4320
rect 1995 -4150 2025 -4140
rect 1995 -4170 2000 -4150
rect 2020 -4170 2025 -4150
rect 1995 -4200 2025 -4170
rect 1995 -4220 2000 -4200
rect 2020 -4220 2025 -4200
rect 1995 -4250 2025 -4220
rect 1995 -4270 2000 -4250
rect 2020 -4270 2025 -4250
rect 1995 -4300 2025 -4270
rect 1995 -4320 2000 -4300
rect 2020 -4320 2025 -4300
rect 1995 -4330 2025 -4320
rect 2050 -4150 2120 -4140
rect 2050 -4170 2055 -4150
rect 2075 -4170 2095 -4150
rect 2115 -4170 2120 -4150
rect 2050 -4200 2120 -4170
rect 2050 -4220 2055 -4200
rect 2075 -4220 2095 -4200
rect 2115 -4220 2120 -4200
rect 2050 -4250 2120 -4220
rect 2050 -4270 2055 -4250
rect 2075 -4270 2095 -4250
rect 2115 -4270 2120 -4250
rect 2050 -4300 2120 -4270
rect 2050 -4320 2055 -4300
rect 2075 -4320 2095 -4300
rect 2115 -4320 2120 -4300
rect 2050 -4330 2120 -4320
rect 2160 -4150 2190 -4140
rect 2160 -4170 2165 -4150
rect 2185 -4170 2190 -4150
rect 2160 -4200 2190 -4170
rect 2160 -4220 2165 -4200
rect 2185 -4220 2190 -4200
rect 2160 -4250 2190 -4220
rect 2160 -4270 2165 -4250
rect 2185 -4270 2190 -4250
rect 2160 -4300 2190 -4270
rect 2160 -4320 2165 -4300
rect 2185 -4320 2190 -4300
rect 2160 -4330 2190 -4320
rect 2215 -4150 2285 -4140
rect 2215 -4170 2220 -4150
rect 2240 -4170 2260 -4150
rect 2280 -4170 2285 -4150
rect 2215 -4200 2285 -4170
rect 2215 -4220 2220 -4200
rect 2240 -4220 2260 -4200
rect 2280 -4220 2285 -4200
rect 2215 -4250 2285 -4220
rect 2215 -4270 2220 -4250
rect 2240 -4270 2260 -4250
rect 2280 -4270 2285 -4250
rect 2215 -4300 2285 -4270
rect 2215 -4320 2220 -4300
rect 2240 -4320 2260 -4300
rect 2280 -4320 2285 -4300
rect 2215 -4330 2285 -4320
rect 1580 -4350 1600 -4330
rect 1580 -4370 1655 -4350
rect 1830 -4365 1850 -4330
rect 1995 -4365 2015 -4330
rect 2160 -4365 2180 -4330
rect 1415 -4400 1555 -4390
rect 1415 -4420 1425 -4400
rect 1445 -4410 1555 -4400
rect 1445 -4420 1455 -4410
rect 1415 -4430 1455 -4420
rect 1635 -4450 1655 -4370
rect 1720 -4375 1760 -4365
rect 1720 -4395 1730 -4375
rect 1750 -4395 1760 -4375
rect 1720 -4405 1760 -4395
rect 1800 -4375 1850 -4365
rect 1800 -4395 1810 -4375
rect 1830 -4395 1850 -4375
rect 1800 -4405 1850 -4395
rect 1965 -4375 2015 -4365
rect 1965 -4395 1975 -4375
rect 1995 -4395 2015 -4375
rect 1965 -4405 2015 -4395
rect 2130 -4375 2180 -4365
rect 2130 -4395 2140 -4375
rect 2160 -4395 2180 -4375
rect 2130 -4405 2180 -4395
rect 2260 -4375 2300 -4365
rect 2260 -4395 2270 -4375
rect 2290 -4395 2300 -4375
rect 2260 -4405 2300 -4395
rect 1830 -4450 1850 -4405
rect 1995 -4450 2015 -4405
rect 2160 -4450 2180 -4405
rect 825 -4460 895 -4450
rect 825 -4480 830 -4460
rect 850 -4480 870 -4460
rect 890 -4480 895 -4460
rect 825 -4510 895 -4480
rect 825 -4530 830 -4510
rect 850 -4530 870 -4510
rect 890 -4530 895 -4510
rect 825 -4540 895 -4530
rect 920 -4460 950 -4450
rect 920 -4480 925 -4460
rect 945 -4480 950 -4460
rect 920 -4510 950 -4480
rect 920 -4530 925 -4510
rect 945 -4530 950 -4510
rect 920 -4540 950 -4530
rect 975 -4460 1005 -4450
rect 975 -4480 980 -4460
rect 1000 -4480 1005 -4460
rect 975 -4510 1005 -4480
rect 975 -4530 980 -4510
rect 1000 -4530 1005 -4510
rect 975 -4540 1005 -4530
rect 1125 -4460 1155 -4450
rect 1125 -4480 1130 -4460
rect 1150 -4480 1155 -4460
rect 1125 -4510 1155 -4480
rect 1125 -4530 1130 -4510
rect 1150 -4530 1155 -4510
rect 1125 -4540 1155 -4530
rect 1180 -4460 1210 -4450
rect 1180 -4480 1185 -4460
rect 1205 -4480 1210 -4460
rect 1180 -4510 1210 -4480
rect 1180 -4530 1185 -4510
rect 1205 -4530 1210 -4510
rect 1180 -4540 1210 -4530
rect 1235 -4460 1345 -4450
rect 1235 -4480 1240 -4460
rect 1260 -4480 1280 -4460
rect 1300 -4480 1320 -4460
rect 1340 -4480 1345 -4460
rect 1235 -4510 1345 -4480
rect 1235 -4530 1240 -4510
rect 1260 -4530 1280 -4510
rect 1300 -4530 1320 -4510
rect 1340 -4530 1345 -4510
rect 1235 -4540 1345 -4530
rect 1370 -4460 1400 -4450
rect 1370 -4480 1375 -4460
rect 1395 -4480 1400 -4460
rect 1370 -4510 1400 -4480
rect 1370 -4530 1375 -4510
rect 1395 -4530 1400 -4510
rect 1370 -4540 1400 -4530
rect 1425 -4460 1455 -4450
rect 1425 -4480 1430 -4460
rect 1450 -4480 1455 -4460
rect 1425 -4510 1455 -4480
rect 1425 -4530 1430 -4510
rect 1450 -4530 1455 -4510
rect 1425 -4540 1455 -4530
rect 1575 -4460 1605 -4450
rect 1575 -4480 1580 -4460
rect 1600 -4480 1605 -4460
rect 1575 -4510 1605 -4480
rect 1575 -4530 1580 -4510
rect 1600 -4530 1605 -4510
rect 1575 -4540 1605 -4530
rect 1630 -4460 1660 -4450
rect 1630 -4480 1635 -4460
rect 1655 -4480 1660 -4460
rect 1630 -4510 1660 -4480
rect 1630 -4530 1635 -4510
rect 1655 -4530 1660 -4510
rect 1630 -4540 1660 -4530
rect 1685 -4460 1755 -4450
rect 1685 -4480 1690 -4460
rect 1710 -4480 1730 -4460
rect 1750 -4480 1755 -4460
rect 1685 -4510 1755 -4480
rect 1685 -4530 1690 -4510
rect 1710 -4530 1730 -4510
rect 1750 -4530 1755 -4510
rect 1685 -4540 1755 -4530
rect 1830 -4460 1860 -4450
rect 1830 -4480 1835 -4460
rect 1855 -4480 1860 -4460
rect 1830 -4510 1860 -4480
rect 1830 -4530 1835 -4510
rect 1855 -4530 1860 -4510
rect 1830 -4540 1860 -4530
rect 1885 -4460 1955 -4450
rect 1885 -4480 1890 -4460
rect 1910 -4480 1930 -4460
rect 1950 -4480 1955 -4460
rect 1885 -4510 1955 -4480
rect 1885 -4530 1890 -4510
rect 1910 -4530 1930 -4510
rect 1950 -4530 1955 -4510
rect 1885 -4540 1955 -4530
rect 1995 -4460 2025 -4450
rect 1995 -4480 2000 -4460
rect 2020 -4480 2025 -4460
rect 1995 -4510 2025 -4480
rect 1995 -4530 2000 -4510
rect 2020 -4530 2025 -4510
rect 1995 -4540 2025 -4530
rect 2050 -4460 2120 -4450
rect 2050 -4480 2055 -4460
rect 2075 -4480 2095 -4460
rect 2115 -4480 2120 -4460
rect 2050 -4510 2120 -4480
rect 2050 -4530 2055 -4510
rect 2075 -4530 2095 -4510
rect 2115 -4530 2120 -4510
rect 2050 -4540 2120 -4530
rect 2160 -4460 2190 -4450
rect 2160 -4480 2165 -4460
rect 2185 -4480 2190 -4460
rect 2160 -4510 2190 -4480
rect 2160 -4530 2165 -4510
rect 2185 -4530 2190 -4510
rect 2160 -4540 2190 -4530
rect 2215 -4460 2285 -4450
rect 2215 -4480 2220 -4460
rect 2240 -4480 2260 -4460
rect 2280 -4480 2285 -4460
rect 2215 -4510 2285 -4480
rect 2215 -4530 2220 -4510
rect 2240 -4530 2260 -4510
rect 2280 -4530 2285 -4510
rect 2215 -4540 2285 -4530
rect 650 -4620 700 -4605
rect 650 -4640 665 -4620
rect 685 -4625 700 -4620
rect 870 -4625 890 -4540
rect 980 -4625 1000 -4540
rect 1130 -4625 1150 -4540
rect 1245 -4625 1265 -4540
rect 1320 -4625 1340 -4540
rect 1430 -4625 1450 -4540
rect 1580 -4625 1600 -4540
rect 1690 -4625 1710 -4540
rect 1890 -4625 1910 -4540
rect 2055 -4625 2075 -4540
rect 2220 -4625 2240 -4540
rect 685 -4640 730 -4625
rect 650 -4645 730 -4640
rect 750 -4645 780 -4625
rect 800 -4645 830 -4625
rect 850 -4645 880 -4625
rect 900 -4645 930 -4625
rect 950 -4645 980 -4625
rect 1000 -4645 1030 -4625
rect 1050 -4645 1080 -4625
rect 1100 -4645 1130 -4625
rect 1150 -4645 1180 -4625
rect 1200 -4645 1230 -4625
rect 1250 -4645 1280 -4625
rect 1300 -4645 1330 -4625
rect 1350 -4645 1380 -4625
rect 1400 -4645 1430 -4625
rect 1450 -4645 1480 -4625
rect 1500 -4645 1530 -4625
rect 1550 -4645 1580 -4625
rect 1600 -4645 1630 -4625
rect 1650 -4645 1680 -4625
rect 1700 -4645 1730 -4625
rect 1750 -4645 1780 -4625
rect 1800 -4645 1830 -4625
rect 1850 -4645 1880 -4625
rect 1900 -4645 1930 -4625
rect 1950 -4645 1980 -4625
rect 2000 -4645 2030 -4625
rect 2050 -4645 2080 -4625
rect 2100 -4645 2130 -4625
rect 2150 -4645 2180 -4625
rect 2200 -4645 2230 -4625
rect 2250 -4645 2280 -4625
rect 2300 -4645 2310 -4625
rect 650 -4655 700 -4645
<< viali >>
rect 665 -3470 685 -3450
rect 730 -3465 750 -3445
rect 780 -3465 800 -3445
rect 830 -3465 850 -3445
rect 880 -3465 900 -3445
rect 930 -3465 950 -3445
rect 980 -3465 1000 -3445
rect 1030 -3465 1050 -3445
rect 1080 -3465 1100 -3445
rect 1130 -3465 1150 -3445
rect 1180 -3465 1200 -3445
rect 1230 -3465 1250 -3445
rect 1280 -3465 1300 -3445
rect 1330 -3465 1350 -3445
rect 1380 -3465 1400 -3445
rect 1430 -3465 1450 -3445
rect 1480 -3465 1500 -3445
rect 1530 -3465 1550 -3445
rect 1580 -3465 1600 -3445
rect 1630 -3465 1650 -3445
rect 1680 -3465 1700 -3445
rect 1730 -3465 1750 -3445
rect 1780 -3465 1800 -3445
rect 1830 -3465 1850 -3445
rect 1880 -3465 1900 -3445
rect 1930 -3465 1950 -3445
rect 1980 -3465 2000 -3445
rect 2030 -3465 2050 -3445
rect 2080 -3465 2100 -3445
rect 2130 -3465 2150 -3445
rect 2180 -3465 2200 -3445
rect 2230 -3465 2250 -3445
rect 2280 -3465 2300 -3445
rect 1075 -3520 1095 -3500
rect 1895 -3520 1915 -3500
rect 1720 -3695 1740 -3675
rect 2265 -3715 2285 -3695
rect 1810 -4000 1830 -3980
rect 830 -4055 850 -4035
rect 880 -4055 900 -4035
rect 930 -4055 950 -4035
rect 980 -4055 1000 -4035
rect 1030 -4055 1050 -4035
rect 1080 -4055 1100 -4035
rect 1130 -4055 1150 -4035
rect 1180 -4055 1200 -4035
rect 1230 -4055 1250 -4035
rect 1280 -4055 1300 -4035
rect 1330 -4055 1350 -4035
rect 1380 -4055 1400 -4035
rect 1430 -4055 1450 -4035
rect 1480 -4055 1500 -4035
rect 1530 -4055 1550 -4035
rect 1580 -4055 1600 -4035
rect 1630 -4055 1650 -4035
rect 1680 -4055 1700 -4035
rect 1730 -4055 1750 -4035
rect 1780 -4055 1800 -4035
rect 1830 -4055 1850 -4035
rect 1880 -4055 1900 -4035
rect 1930 -4055 1950 -4035
rect 1980 -4055 2000 -4035
rect 2030 -4055 2050 -4035
rect 2080 -4055 2100 -4035
rect 2130 -4055 2150 -4035
rect 2180 -4055 2200 -4035
rect 2230 -4055 2250 -4035
rect 2280 -4055 2300 -4035
rect 1095 -4110 1115 -4090
rect 1730 -4395 1750 -4375
rect 2270 -4395 2290 -4375
rect 665 -4640 685 -4620
rect 730 -4645 750 -4625
rect 780 -4645 800 -4625
rect 830 -4645 850 -4625
rect 880 -4645 900 -4625
rect 930 -4645 950 -4625
rect 980 -4645 1000 -4625
rect 1030 -4645 1050 -4625
rect 1080 -4645 1100 -4625
rect 1130 -4645 1150 -4625
rect 1180 -4645 1200 -4625
rect 1230 -4645 1250 -4625
rect 1280 -4645 1300 -4625
rect 1330 -4645 1350 -4625
rect 1380 -4645 1400 -4625
rect 1430 -4645 1450 -4625
rect 1480 -4645 1500 -4625
rect 1530 -4645 1550 -4625
rect 1580 -4645 1600 -4625
rect 1630 -4645 1650 -4625
rect 1680 -4645 1700 -4625
rect 1730 -4645 1750 -4625
rect 1780 -4645 1800 -4625
rect 1830 -4645 1850 -4625
rect 1880 -4645 1900 -4625
rect 1930 -4645 1950 -4625
rect 1980 -4645 2000 -4625
rect 2030 -4645 2050 -4625
rect 2080 -4645 2100 -4625
rect 2130 -4645 2150 -4625
rect 2180 -4645 2200 -4625
rect 2230 -4645 2250 -4625
rect 2280 -4645 2300 -4625
<< metal1 >>
rect 650 -3445 2310 -3435
rect 650 -3475 660 -3445
rect 690 -3465 730 -3445
rect 750 -3465 780 -3445
rect 800 -3465 830 -3445
rect 850 -3465 880 -3445
rect 900 -3465 930 -3445
rect 950 -3465 980 -3445
rect 1000 -3465 1030 -3445
rect 1050 -3465 1080 -3445
rect 1100 -3465 1130 -3445
rect 1150 -3465 1180 -3445
rect 1200 -3465 1230 -3445
rect 1250 -3465 1280 -3445
rect 1300 -3465 1330 -3445
rect 1350 -3465 1380 -3445
rect 1400 -3465 1430 -3445
rect 1450 -3465 1480 -3445
rect 1500 -3465 1530 -3445
rect 1550 -3465 1580 -3445
rect 1600 -3465 1630 -3445
rect 1650 -3465 1680 -3445
rect 1700 -3465 1730 -3445
rect 1750 -3465 1780 -3445
rect 1800 -3465 1830 -3445
rect 1850 -3465 1880 -3445
rect 1900 -3465 1930 -3445
rect 1950 -3465 1980 -3445
rect 2000 -3465 2030 -3445
rect 2050 -3465 2080 -3445
rect 2100 -3465 2130 -3445
rect 2150 -3465 2180 -3445
rect 2200 -3465 2230 -3445
rect 2250 -3465 2280 -3445
rect 2300 -3465 2310 -3445
rect 690 -3475 2310 -3465
rect 650 -3485 700 -3475
rect 1065 -3500 1105 -3490
rect 1065 -3520 1075 -3500
rect 1095 -3510 1105 -3500
rect 1885 -3500 1925 -3490
rect 1885 -3510 1895 -3500
rect 1095 -3520 1895 -3510
rect 1915 -3510 1925 -3500
rect 1915 -3520 2310 -3510
rect 1065 -3530 2310 -3520
rect 1710 -3670 1750 -3665
rect 1710 -3700 1715 -3670
rect 1745 -3700 1750 -3670
rect 1710 -3705 1750 -3700
rect 2255 -3690 2295 -3685
rect 2255 -3720 2260 -3690
rect 2290 -3720 2295 -3690
rect 2255 -3725 2295 -3720
rect 1800 -3975 1840 -3970
rect 1800 -4005 1805 -3975
rect 1835 -4005 1840 -3975
rect 1800 -4010 1840 -4005
rect 800 -4035 2310 -4025
rect 800 -4055 830 -4035
rect 850 -4055 880 -4035
rect 900 -4055 930 -4035
rect 950 -4055 980 -4035
rect 1000 -4055 1030 -4035
rect 1050 -4055 1080 -4035
rect 1100 -4055 1130 -4035
rect 1150 -4055 1180 -4035
rect 1200 -4055 1230 -4035
rect 1250 -4055 1280 -4035
rect 1300 -4055 1330 -4035
rect 1350 -4055 1380 -4035
rect 1400 -4055 1430 -4035
rect 1450 -4055 1480 -4035
rect 1500 -4055 1530 -4035
rect 1550 -4055 1580 -4035
rect 1600 -4055 1630 -4035
rect 1650 -4055 1680 -4035
rect 1700 -4055 1730 -4035
rect 1750 -4055 1780 -4035
rect 1800 -4055 1830 -4035
rect 1850 -4055 1880 -4035
rect 1900 -4055 1930 -4035
rect 1950 -4055 1980 -4035
rect 2000 -4055 2030 -4035
rect 2050 -4055 2080 -4035
rect 2100 -4055 2130 -4035
rect 2150 -4055 2180 -4035
rect 2200 -4055 2230 -4035
rect 2250 -4055 2280 -4035
rect 2300 -4055 2310 -4035
rect 800 -4065 2310 -4055
rect 1085 -4090 1125 -4080
rect 1085 -4110 1095 -4090
rect 1115 -4095 1125 -4090
rect 1115 -4100 2310 -4095
rect 1115 -4110 1775 -4100
rect 1085 -4115 1775 -4110
rect 1085 -4120 1125 -4115
rect 1770 -4130 1775 -4115
rect 1805 -4115 2310 -4100
rect 1805 -4130 1810 -4115
rect 1770 -4135 1810 -4130
rect 1720 -4370 1760 -4365
rect 1720 -4400 1725 -4370
rect 1755 -4400 1760 -4370
rect 1720 -4405 1760 -4400
rect 2260 -4370 2300 -4365
rect 2260 -4400 2265 -4370
rect 2295 -4400 2300 -4370
rect 2260 -4405 2300 -4400
rect 650 -4615 700 -4605
rect 650 -4645 660 -4615
rect 690 -4625 2310 -4615
rect 690 -4645 730 -4625
rect 750 -4645 780 -4625
rect 800 -4645 830 -4625
rect 850 -4645 880 -4625
rect 900 -4645 930 -4625
rect 950 -4645 980 -4625
rect 1000 -4645 1030 -4625
rect 1050 -4645 1080 -4625
rect 1100 -4645 1130 -4625
rect 1150 -4645 1180 -4625
rect 1200 -4645 1230 -4625
rect 1250 -4645 1280 -4625
rect 1300 -4645 1330 -4625
rect 1350 -4645 1380 -4625
rect 1400 -4645 1430 -4625
rect 1450 -4645 1480 -4625
rect 1500 -4645 1530 -4625
rect 1550 -4645 1580 -4625
rect 1600 -4645 1630 -4625
rect 1650 -4645 1680 -4625
rect 1700 -4645 1730 -4625
rect 1750 -4645 1780 -4625
rect 1800 -4645 1830 -4625
rect 1850 -4645 1880 -4625
rect 1900 -4645 1930 -4625
rect 1950 -4645 1980 -4625
rect 2000 -4645 2030 -4625
rect 2050 -4645 2080 -4625
rect 2100 -4645 2130 -4625
rect 2150 -4645 2180 -4625
rect 2200 -4645 2230 -4625
rect 2250 -4645 2280 -4625
rect 2300 -4645 2310 -4625
rect 650 -4655 2310 -4645
<< via1 >>
rect 660 -3450 690 -3445
rect 660 -3470 665 -3450
rect 665 -3470 685 -3450
rect 685 -3470 690 -3450
rect 660 -3475 690 -3470
rect 1715 -3675 1745 -3670
rect 1715 -3695 1720 -3675
rect 1720 -3695 1740 -3675
rect 1740 -3695 1745 -3675
rect 1715 -3700 1745 -3695
rect 2260 -3695 2290 -3690
rect 2260 -3715 2265 -3695
rect 2265 -3715 2285 -3695
rect 2285 -3715 2290 -3695
rect 2260 -3720 2290 -3715
rect 1805 -3980 1835 -3975
rect 1805 -4000 1810 -3980
rect 1810 -4000 1830 -3980
rect 1830 -4000 1835 -3980
rect 1805 -4005 1835 -4000
rect 1775 -4130 1805 -4100
rect 1725 -4375 1755 -4370
rect 1725 -4395 1730 -4375
rect 1730 -4395 1750 -4375
rect 1750 -4395 1755 -4375
rect 1725 -4400 1755 -4395
rect 2265 -4375 2295 -4370
rect 2265 -4395 2270 -4375
rect 2270 -4395 2290 -4375
rect 2290 -4395 2295 -4375
rect 2265 -4400 2295 -4395
rect 660 -4620 690 -4615
rect 660 -4640 665 -4620
rect 665 -4640 685 -4620
rect 685 -4640 690 -4620
rect 660 -4645 690 -4640
<< metal2 >>
rect 650 -3445 700 -3435
rect 650 -3475 660 -3445
rect 690 -3475 700 -3445
rect 650 -3485 700 -3475
rect 1710 -3670 1750 -3665
rect 1710 -3700 1715 -3670
rect 1745 -3700 1750 -3670
rect 1710 -3705 1750 -3700
rect 1730 -4365 1750 -3705
rect 2255 -3690 2300 -3685
rect 2255 -3720 2260 -3690
rect 2290 -3720 2300 -3690
rect 2255 -3725 2300 -3720
rect 1790 -3975 1840 -3970
rect 1790 -4005 1805 -3975
rect 1835 -4005 1840 -3975
rect 1790 -4010 1840 -4005
rect 1790 -4095 1810 -4010
rect 1770 -4100 1810 -4095
rect 1770 -4130 1775 -4100
rect 1805 -4130 1810 -4100
rect 1770 -4135 1810 -4130
rect 2280 -4365 2300 -3725
rect 1720 -4370 1760 -4365
rect 1720 -4400 1725 -4370
rect 1755 -4400 1760 -4370
rect 1720 -4405 1760 -4400
rect 2260 -4370 2300 -4365
rect 2260 -4400 2265 -4370
rect 2295 -4400 2300 -4370
rect 2260 -4405 2300 -4400
rect 650 -4615 700 -4605
rect 650 -4645 660 -4615
rect 690 -4645 700 -4615
rect 650 -4655 700 -4645
<< via2 >>
rect 660 -3475 690 -3445
rect 660 -4645 690 -4615
<< metal3 >>
rect 650 -3440 700 -3435
rect 650 -3480 655 -3440
rect 695 -3480 700 -3440
rect 650 -3485 700 -3480
rect 650 -4610 700 -4605
rect 650 -4650 655 -4610
rect 695 -4650 700 -4610
rect 650 -4655 700 -4650
<< via3 >>
rect 655 -3445 695 -3440
rect 655 -3475 660 -3445
rect 660 -3475 690 -3445
rect 690 -3475 695 -3445
rect 655 -3480 695 -3475
rect 655 -4615 695 -4610
rect 655 -4645 660 -4615
rect 660 -4645 690 -4615
rect 690 -4645 695 -4615
rect 655 -4650 695 -4645
<< metal4 >>
rect 650 -3440 700 -3435
rect 650 -3480 655 -3440
rect 695 -3480 700 -3440
rect 650 -4610 700 -3480
rect 650 -4650 655 -4610
rect 695 -4650 700 -4610
rect 650 -4655 700 -4650
<< labels >>
flabel locali 1085 -4120 1085 -4120 7 FreeSans 160 0 -80 0 QB
port 6 w
flabel locali 1085 -3585 1085 -3585 7 FreeSans 160 0 -80 0 QA
port 5 w
flabel metal1 800 -4045 800 -4045 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel metal4 650 -4520 650 -4520 7 FreeSans 160 0 -80 0 GNDA
port 4 w
flabel locali 1800 -4405 1800 -4405 5 FreeSans 160 0 0 -80 Reset
flabel locali 1655 -4370 1655 -4370 3 FreeSans 160 0 80 0 F_b
flabel locali 1450 -4370 1450 -4370 3 FreeSans 160 0 80 0 F
flabel poly 1050 -4240 1050 -4240 7 FreeSans 160 0 -80 0 QB_b
flabel poly 840 -4405 840 -4405 7 FreeSans 160 0 -80 0 F_VCO
port 2 w
flabel poly 840 -3690 840 -3690 7 FreeSans 160 0 -80 0 F_REF
port 1 w
flabel poly 1050 -3720 1050 -3720 7 FreeSans 160 0 -80 0 QA_b
flabel locali 1655 -3720 1655 -3720 3 FreeSans 160 0 80 0 E_b
flabel locali 1450 -3720 1450 -3720 3 FreeSans 160 0 80 0 E
flabel locali 1965 -3685 1965 -3685 3 FreeSans 160 0 80 0 before_Reset
<< end >>
