magic
tech sky130A
timestamp 1738662969
<< error_p >>
rect 4145 1837 4165 1840
rect 4145 1748 4148 1837
rect 4162 1748 4165 1837
rect 4145 1745 4165 1748
rect 4345 1837 4365 1840
rect 4345 1748 4348 1837
rect 4362 1748 4365 1837
rect 4345 1745 4365 1748
rect 4545 1837 4565 1840
rect 4545 1748 4548 1837
rect 4562 1748 4565 1837
rect 4545 1745 4565 1748
rect 4745 1837 4765 1840
rect 4745 1748 4748 1837
rect 4762 1748 4765 1837
rect 4745 1745 4765 1748
rect 4925 1837 4945 1840
rect 4925 1748 4928 1837
rect 4942 1748 4945 1837
rect 4925 1745 4945 1748
rect 4435 1675 4475 1678
<< nwell >>
rect 4010 2185 5060 2685
<< nmos >>
rect 4080 1975 4095 2025
rect 4145 1975 4160 2025
rect 4210 1975 4225 2025
rect 4275 1975 4290 2025
rect 4440 1975 4455 2025
rect 4505 1975 4520 2025
rect 4570 1975 4585 2025
rect 4635 1975 4650 2025
rect 4780 1975 4795 2025
rect 4845 1975 4860 2025
rect 4910 1975 4925 2025
rect 4975 1975 4990 2025
rect 4080 1730 4130 1855
rect 4180 1730 4230 1855
rect 4280 1730 4330 1855
rect 4380 1730 4430 1855
rect 4480 1730 4530 1855
rect 4580 1730 4630 1855
rect 4680 1730 4730 1855
rect 4780 1730 4830 1855
<< pmos >>
rect 4095 2380 4145 2630
rect 4195 2380 4245 2630
rect 4295 2380 4345 2630
rect 4395 2380 4445 2630
rect 4495 2380 4545 2630
rect 4595 2380 4645 2630
rect 4695 2380 4745 2630
rect 4795 2380 4845 2630
rect 4080 2210 4095 2310
rect 4145 2210 4160 2310
rect 4210 2210 4225 2310
rect 4275 2210 4290 2310
rect 4440 2210 4455 2310
rect 4505 2210 4520 2310
rect 4570 2210 4585 2310
rect 4635 2210 4650 2310
rect 4780 2210 4795 2310
rect 4845 2210 4860 2310
rect 4910 2210 4925 2310
rect 4975 2210 4990 2310
<< ndiff >>
rect 4030 2010 4080 2025
rect 4030 1990 4045 2010
rect 4065 1990 4080 2010
rect 4030 1975 4080 1990
rect 4095 2010 4145 2025
rect 4095 1990 4110 2010
rect 4130 1990 4145 2010
rect 4095 1975 4145 1990
rect 4160 2010 4210 2025
rect 4160 1990 4175 2010
rect 4195 1990 4210 2010
rect 4160 1975 4210 1990
rect 4225 2010 4275 2025
rect 4225 1990 4240 2010
rect 4260 1990 4275 2010
rect 4225 1975 4275 1990
rect 4290 2010 4340 2025
rect 4290 1990 4305 2010
rect 4325 1990 4340 2010
rect 4290 1975 4340 1990
rect 4390 2010 4440 2025
rect 4390 1990 4405 2010
rect 4425 1990 4440 2010
rect 4390 1975 4440 1990
rect 4455 2010 4505 2025
rect 4455 1990 4470 2010
rect 4490 1990 4505 2010
rect 4455 1975 4505 1990
rect 4520 2010 4570 2025
rect 4520 1990 4535 2010
rect 4555 1990 4570 2010
rect 4520 1975 4570 1990
rect 4585 2010 4635 2025
rect 4585 1990 4600 2010
rect 4620 1990 4635 2010
rect 4585 1975 4635 1990
rect 4650 2010 4700 2025
rect 4650 1990 4665 2010
rect 4685 1990 4700 2010
rect 4650 1975 4700 1990
rect 4730 2010 4780 2025
rect 4730 1990 4745 2010
rect 4765 1990 4780 2010
rect 4730 1975 4780 1990
rect 4795 2010 4845 2025
rect 4795 1990 4810 2010
rect 4830 1990 4845 2010
rect 4795 1975 4845 1990
rect 4860 2010 4910 2025
rect 4860 1990 4875 2010
rect 4895 1990 4910 2010
rect 4860 1975 4910 1990
rect 4925 2010 4975 2025
rect 4925 1990 4940 2010
rect 4960 1990 4975 2010
rect 4925 1975 4975 1990
rect 4990 2010 5040 2025
rect 4990 1990 5005 2010
rect 5025 1990 5040 2010
rect 4990 1975 5040 1990
rect 4030 1840 4080 1855
rect 4030 1745 4045 1840
rect 4065 1745 4080 1840
rect 4030 1730 4080 1745
rect 4130 1840 4180 1855
rect 4130 1745 4145 1840
rect 4165 1745 4180 1840
rect 4130 1730 4180 1745
rect 4230 1840 4280 1855
rect 4230 1745 4245 1840
rect 4265 1745 4280 1840
rect 4230 1730 4280 1745
rect 4330 1840 4380 1855
rect 4330 1745 4345 1840
rect 4365 1745 4380 1840
rect 4330 1730 4380 1745
rect 4430 1840 4480 1855
rect 4430 1745 4445 1840
rect 4465 1745 4480 1840
rect 4430 1730 4480 1745
rect 4530 1840 4580 1855
rect 4530 1745 4545 1840
rect 4565 1745 4580 1840
rect 4530 1730 4580 1745
rect 4630 1840 4680 1855
rect 4630 1745 4645 1840
rect 4665 1745 4680 1840
rect 4630 1730 4680 1745
rect 4730 1840 4780 1855
rect 4730 1745 4745 1840
rect 4765 1745 4780 1840
rect 4730 1730 4780 1745
rect 4830 1840 4880 1855
rect 4830 1745 4845 1840
rect 4865 1745 4880 1840
rect 4830 1730 4880 1745
<< pdiff >>
rect 4045 2615 4095 2630
rect 4045 2395 4060 2615
rect 4080 2395 4095 2615
rect 4045 2380 4095 2395
rect 4145 2615 4195 2630
rect 4145 2395 4160 2615
rect 4180 2395 4195 2615
rect 4145 2380 4195 2395
rect 4245 2615 4295 2630
rect 4245 2395 4260 2615
rect 4280 2395 4295 2615
rect 4245 2380 4295 2395
rect 4345 2615 4395 2630
rect 4345 2395 4360 2615
rect 4380 2395 4395 2615
rect 4345 2380 4395 2395
rect 4445 2615 4495 2630
rect 4445 2395 4460 2615
rect 4480 2395 4495 2615
rect 4445 2380 4495 2395
rect 4545 2615 4595 2630
rect 4545 2395 4560 2615
rect 4580 2395 4595 2615
rect 4545 2380 4595 2395
rect 4645 2615 4695 2630
rect 4645 2395 4660 2615
rect 4680 2395 4695 2615
rect 4645 2380 4695 2395
rect 4745 2615 4795 2630
rect 4745 2395 4760 2615
rect 4780 2395 4795 2615
rect 4745 2380 4795 2395
rect 4845 2615 4895 2630
rect 4845 2395 4860 2615
rect 4880 2395 4895 2615
rect 4845 2380 4895 2395
rect 4030 2295 4080 2310
rect 4030 2225 4045 2295
rect 4065 2225 4080 2295
rect 4030 2210 4080 2225
rect 4095 2295 4145 2310
rect 4095 2225 4110 2295
rect 4130 2225 4145 2295
rect 4095 2210 4145 2225
rect 4160 2295 4210 2310
rect 4160 2225 4175 2295
rect 4195 2225 4210 2295
rect 4160 2210 4210 2225
rect 4225 2295 4275 2310
rect 4225 2225 4240 2295
rect 4260 2225 4275 2295
rect 4225 2210 4275 2225
rect 4290 2295 4340 2310
rect 4290 2225 4305 2295
rect 4325 2225 4340 2295
rect 4290 2210 4340 2225
rect 4390 2295 4440 2310
rect 4390 2225 4405 2295
rect 4425 2225 4440 2295
rect 4390 2210 4440 2225
rect 4455 2295 4505 2310
rect 4455 2225 4470 2295
rect 4490 2225 4505 2295
rect 4455 2210 4505 2225
rect 4520 2295 4570 2310
rect 4520 2225 4535 2295
rect 4555 2225 4570 2295
rect 4520 2210 4570 2225
rect 4585 2295 4635 2310
rect 4585 2225 4600 2295
rect 4620 2225 4635 2295
rect 4585 2210 4635 2225
rect 4650 2295 4700 2310
rect 4650 2225 4665 2295
rect 4685 2225 4700 2295
rect 4650 2210 4700 2225
rect 4730 2295 4780 2310
rect 4730 2225 4745 2295
rect 4765 2225 4780 2295
rect 4730 2210 4780 2225
rect 4795 2295 4845 2310
rect 4795 2225 4810 2295
rect 4830 2225 4845 2295
rect 4795 2210 4845 2225
rect 4860 2295 4910 2310
rect 4860 2225 4875 2295
rect 4895 2225 4910 2295
rect 4860 2210 4910 2225
rect 4925 2295 4975 2310
rect 4925 2225 4940 2295
rect 4960 2225 4975 2295
rect 4925 2210 4975 2225
rect 4990 2295 5040 2310
rect 4990 2225 5005 2295
rect 5025 2225 5040 2295
rect 4990 2210 5040 2225
<< ndiffc >>
rect 4045 1990 4065 2010
rect 4110 1990 4130 2010
rect 4175 1990 4195 2010
rect 4240 1990 4260 2010
rect 4305 1990 4325 2010
rect 4405 1990 4425 2010
rect 4470 1990 4490 2010
rect 4535 1990 4555 2010
rect 4600 1990 4620 2010
rect 4665 1990 4685 2010
rect 4745 1990 4765 2010
rect 4810 1990 4830 2010
rect 4875 1990 4895 2010
rect 4940 1990 4960 2010
rect 5005 1990 5025 2010
rect 4045 1745 4065 1840
rect 4145 1745 4165 1840
rect 4245 1745 4265 1840
rect 4345 1745 4365 1840
rect 4445 1745 4465 1840
rect 4545 1745 4565 1840
rect 4645 1745 4665 1840
rect 4745 1745 4765 1840
rect 4845 1745 4865 1840
<< pdiffc >>
rect 4060 2395 4080 2615
rect 4160 2395 4180 2615
rect 4260 2395 4280 2615
rect 4360 2395 4380 2615
rect 4460 2395 4480 2615
rect 4560 2395 4580 2615
rect 4660 2395 4680 2615
rect 4760 2395 4780 2615
rect 4860 2395 4880 2615
rect 4045 2225 4065 2295
rect 4110 2225 4130 2295
rect 4175 2225 4195 2295
rect 4240 2225 4260 2295
rect 4305 2225 4325 2295
rect 4405 2225 4425 2295
rect 4470 2225 4490 2295
rect 4535 2225 4555 2295
rect 4600 2225 4620 2295
rect 4665 2225 4685 2295
rect 4745 2225 4765 2295
rect 4810 2225 4830 2295
rect 4875 2225 4895 2295
rect 4940 2225 4960 2295
rect 5005 2225 5025 2295
<< psubdiff >>
rect 4910 1840 4960 1855
rect 4910 1745 4925 1840
rect 4945 1745 4960 1840
rect 4910 1730 4960 1745
<< nsubdiff >>
rect 4940 2615 4990 2630
rect 4940 2395 4955 2615
rect 4975 2395 4990 2615
rect 4940 2380 4990 2395
<< psubdiffcont >>
rect 4925 1745 4945 1840
<< nsubdiffcont >>
rect 4955 2395 4975 2615
<< poly >>
rect 4075 2675 4115 2685
rect 4075 2655 4085 2675
rect 4105 2655 4115 2675
rect 4450 2675 4490 2685
rect 4450 2655 4460 2675
rect 4480 2655 4490 2675
rect 4830 2675 4870 2685
rect 4830 2655 4840 2675
rect 4860 2655 4870 2675
rect 4075 2645 4870 2655
rect 4095 2640 4845 2645
rect 4095 2630 4145 2640
rect 4195 2630 4245 2640
rect 4295 2630 4345 2640
rect 4395 2630 4445 2640
rect 4495 2630 4545 2640
rect 4595 2630 4645 2640
rect 4695 2630 4745 2640
rect 4795 2630 4845 2640
rect 4095 2365 4145 2380
rect 4195 2365 4245 2380
rect 4295 2365 4345 2380
rect 4395 2365 4445 2380
rect 4495 2365 4545 2380
rect 4595 2365 4645 2380
rect 4695 2365 4745 2380
rect 4795 2365 4845 2380
rect 4080 2310 4095 2325
rect 4145 2310 4160 2325
rect 4210 2310 4225 2325
rect 4275 2310 4290 2325
rect 4440 2310 4455 2325
rect 4505 2310 4520 2325
rect 4570 2310 4585 2325
rect 4635 2310 4650 2325
rect 4780 2310 4795 2325
rect 4845 2310 4860 2325
rect 4910 2310 4925 2325
rect 4975 2310 4990 2325
rect 5060 2215 5100 2225
rect 4080 2200 4095 2210
rect 4145 2200 4160 2210
rect 4080 2185 4160 2200
rect 4210 2200 4225 2210
rect 4275 2200 4290 2210
rect 4210 2195 4290 2200
rect 4440 2200 4455 2210
rect 4505 2200 4520 2210
rect 4570 2200 4585 2210
rect 4635 2200 4650 2210
rect 4210 2185 4315 2195
rect 4440 2185 4650 2200
rect 4780 2200 4795 2210
rect 4845 2200 4860 2210
rect 4910 2200 4925 2210
rect 4975 2200 4990 2210
rect 5060 2200 5070 2215
rect 4780 2195 5070 2200
rect 5090 2195 5100 2215
rect 4780 2185 5100 2195
rect 4080 2120 4095 2185
rect 4275 2165 4285 2185
rect 4305 2165 4315 2185
rect 4275 2155 4315 2165
rect 4460 2180 4500 2185
rect 4460 2160 4470 2180
rect 4490 2160 4500 2180
rect 4460 2150 4500 2160
rect 4590 2180 4630 2185
rect 4590 2160 4600 2180
rect 4620 2160 4630 2180
rect 4590 2150 4630 2160
rect 4780 2165 4790 2185
rect 4810 2165 4820 2185
rect 4780 2155 4820 2165
rect 3990 2105 4455 2120
rect 4100 2070 4140 2080
rect 4100 2050 4110 2070
rect 4130 2050 4140 2070
rect 4230 2070 4270 2080
rect 4230 2050 4240 2070
rect 4260 2050 4270 2070
rect 4440 2050 4455 2105
rect 4545 2075 4585 2085
rect 4545 2055 4555 2075
rect 4575 2055 4585 2075
rect 4545 2050 4585 2055
rect 4080 2035 4290 2050
rect 4080 2025 4095 2035
rect 4145 2025 4160 2035
rect 4210 2025 4225 2035
rect 4275 2025 4290 2035
rect 4440 2035 4520 2050
rect 4545 2045 4650 2050
rect 4440 2025 4455 2035
rect 4505 2025 4520 2035
rect 4570 2035 4650 2045
rect 4570 2025 4585 2035
rect 4635 2025 4650 2035
rect 4780 2035 4990 2050
rect 4780 2025 4795 2035
rect 4845 2025 4860 2035
rect 4910 2025 4925 2035
rect 4975 2025 4990 2035
rect 4080 1960 4095 1975
rect 4145 1960 4160 1975
rect 4210 1960 4225 1975
rect 4275 1960 4290 1975
rect 4440 1960 4455 1975
rect 4505 1960 4520 1975
rect 4570 1960 4585 1975
rect 4635 1960 4650 1975
rect 4780 1960 4795 1975
rect 4845 1960 4860 1975
rect 4910 1960 4925 1975
rect 4975 1935 4990 1975
rect 4165 1925 4990 1935
rect 4165 1905 4175 1925
rect 4195 1920 4990 1925
rect 4195 1905 4205 1920
rect 4165 1895 4205 1905
rect 4975 1915 4990 1920
rect 4975 1905 5015 1915
rect 4975 1885 4985 1905
rect 5005 1885 5015 1905
rect 4975 1875 5015 1885
rect 4080 1855 4130 1870
rect 4180 1855 4230 1870
rect 4280 1855 4330 1870
rect 4380 1855 4430 1870
rect 4480 1855 4530 1870
rect 4580 1855 4630 1870
rect 4680 1855 4730 1870
rect 4780 1855 4830 1870
rect 4080 1720 4130 1730
rect 4180 1720 4230 1730
rect 4280 1720 4330 1730
rect 4380 1720 4430 1730
rect 4480 1720 4530 1730
rect 4580 1720 4630 1730
rect 4680 1720 4730 1730
rect 4780 1720 4830 1730
rect 4080 1710 4830 1720
rect 4080 1705 4095 1710
rect 4085 1690 4095 1705
rect 4115 1705 4795 1710
rect 4115 1690 4125 1705
rect 4085 1680 4125 1690
rect 4435 1685 4445 1705
rect 4465 1685 4475 1705
rect 4435 1675 4475 1685
rect 4785 1690 4795 1705
rect 4815 1705 4830 1710
rect 4815 1690 4825 1705
rect 4785 1680 4825 1690
<< polycont >>
rect 4085 2655 4105 2675
rect 4460 2655 4480 2675
rect 4840 2655 4860 2675
rect 5070 2195 5090 2215
rect 4285 2165 4305 2185
rect 4470 2160 4490 2180
rect 4600 2160 4620 2180
rect 4790 2165 4810 2185
rect 4110 2050 4130 2070
rect 4240 2050 4260 2070
rect 4555 2055 4575 2075
rect 4175 1905 4195 1925
rect 4985 1885 5005 1905
rect 4095 1690 4115 1710
rect 4445 1685 4465 1705
rect 4795 1690 4815 1710
<< xpolycontact >>
rect 4180 1595 4400 1630
rect 4470 1595 4690 1630
rect 5325 1595 5545 1630
rect 5643 1595 5863 1630
<< xpolyres >>
rect 4400 1595 4470 1630
rect 5545 1595 5643 1630
<< locali >>
rect 4075 2675 4115 2685
rect 4075 2670 4085 2675
rect 3940 2655 4085 2670
rect 4105 2670 4115 2675
rect 4450 2675 4490 2685
rect 4450 2670 4460 2675
rect 4105 2655 4460 2670
rect 4480 2670 4490 2675
rect 4830 2675 4870 2685
rect 4830 2670 4840 2675
rect 4480 2655 4840 2670
rect 4860 2670 4870 2675
rect 4860 2655 4880 2670
rect 3940 2650 4880 2655
rect 3940 1815 3960 2650
rect 4060 2645 4115 2650
rect 4450 2645 4490 2650
rect 4830 2645 4880 2650
rect 4060 2625 4080 2645
rect 4460 2625 4480 2645
rect 4860 2625 4880 2645
rect 4045 2615 4090 2625
rect 4045 2395 4060 2615
rect 4080 2395 4090 2615
rect 4045 2385 4090 2395
rect 4150 2615 4190 2625
rect 4150 2395 4160 2615
rect 4180 2395 4190 2615
rect 4150 2385 4190 2395
rect 4250 2615 4290 2625
rect 4250 2395 4260 2615
rect 4280 2395 4290 2615
rect 4250 2385 4290 2395
rect 4350 2615 4390 2625
rect 4350 2395 4360 2615
rect 4380 2395 4390 2615
rect 4350 2385 4390 2395
rect 4450 2615 4490 2625
rect 4450 2395 4460 2615
rect 4480 2395 4490 2615
rect 4450 2385 4490 2395
rect 4550 2615 4590 2625
rect 4550 2395 4560 2615
rect 4580 2395 4590 2615
rect 4550 2385 4590 2395
rect 4650 2615 4690 2625
rect 4650 2395 4660 2615
rect 4680 2395 4690 2615
rect 4650 2385 4690 2395
rect 4750 2615 4790 2625
rect 4750 2395 4760 2615
rect 4780 2395 4790 2615
rect 4750 2385 4790 2395
rect 4850 2615 4890 2625
rect 4850 2395 4860 2615
rect 4880 2395 4890 2615
rect 4850 2385 4890 2395
rect 4945 2615 4985 2625
rect 4945 2395 4955 2615
rect 4975 2395 4985 2615
rect 4945 2385 4985 2395
rect 4260 2365 4280 2385
rect 4660 2365 4680 2385
rect 4260 2345 4680 2365
rect 4045 2325 4325 2345
rect 4045 2305 4065 2325
rect 4175 2305 4195 2325
rect 4305 2305 4325 2325
rect 4745 2325 5025 2345
rect 4745 2305 4765 2325
rect 4875 2305 4895 2325
rect 5005 2305 5025 2325
rect 4035 2295 4075 2305
rect 4035 2225 4045 2295
rect 4065 2225 4075 2295
rect 4035 2215 4075 2225
rect 4100 2295 4140 2305
rect 4100 2225 4110 2295
rect 4130 2225 4140 2295
rect 4100 2215 4140 2225
rect 4165 2295 4205 2305
rect 4165 2225 4175 2295
rect 4195 2225 4205 2295
rect 4165 2215 4205 2225
rect 4230 2295 4270 2305
rect 4230 2225 4240 2295
rect 4260 2225 4270 2295
rect 4230 2215 4270 2225
rect 4295 2295 4340 2305
rect 4295 2225 4305 2295
rect 4325 2225 4340 2295
rect 4295 2215 4340 2225
rect 4395 2295 4435 2305
rect 4395 2225 4405 2295
rect 4425 2225 4435 2295
rect 4395 2215 4435 2225
rect 4460 2295 4500 2305
rect 4460 2225 4470 2295
rect 4490 2225 4500 2295
rect 4460 2215 4500 2225
rect 4525 2295 4565 2305
rect 4525 2225 4535 2295
rect 4555 2225 4565 2295
rect 4525 2215 4565 2225
rect 4590 2295 4635 2305
rect 4590 2225 4600 2295
rect 4620 2225 4635 2295
rect 4590 2215 4635 2225
rect 4655 2295 4695 2305
rect 4655 2225 4665 2295
rect 4685 2225 4695 2295
rect 4655 2215 4695 2225
rect 4735 2295 4775 2305
rect 4735 2225 4745 2295
rect 4765 2225 4775 2295
rect 4735 2215 4775 2225
rect 4800 2295 4840 2305
rect 4800 2225 4810 2295
rect 4830 2225 4840 2295
rect 4800 2215 4840 2225
rect 4865 2295 4905 2305
rect 4865 2225 4875 2295
rect 4895 2225 4905 2295
rect 4865 2215 4905 2225
rect 4930 2295 4970 2305
rect 4930 2225 4940 2295
rect 4960 2225 4970 2295
rect 4930 2215 4970 2225
rect 4995 2295 5035 2305
rect 4995 2225 5005 2295
rect 5025 2225 5035 2295
rect 4995 2215 5035 2225
rect 5060 2215 5100 2225
rect 4110 2080 4130 2215
rect 4230 2195 4250 2215
rect 4175 2175 4250 2195
rect 4275 2185 4315 2195
rect 4100 2070 4140 2080
rect 4045 2050 4110 2070
rect 4130 2050 4140 2070
rect 4045 2020 4065 2050
rect 4100 2040 4140 2050
rect 4175 2020 4195 2175
rect 4275 2165 4285 2185
rect 4305 2165 4315 2185
rect 4275 2155 4315 2165
rect 4405 2180 4425 2215
rect 4460 2180 4500 2190
rect 4405 2160 4470 2180
rect 4490 2160 4500 2180
rect 4460 2150 4500 2160
rect 4230 2070 4270 2080
rect 4230 2050 4240 2070
rect 4260 2050 4325 2070
rect 4230 2040 4270 2050
rect 4305 2020 4325 2050
rect 4470 2020 4490 2150
rect 4535 2130 4555 2215
rect 4590 2180 4630 2190
rect 4665 2180 4685 2215
rect 4590 2160 4600 2180
rect 4620 2160 4685 2180
rect 4780 2185 4820 2195
rect 4780 2165 4790 2185
rect 4810 2165 4820 2185
rect 4590 2150 4630 2160
rect 4780 2155 4820 2165
rect 5005 2165 5025 2215
rect 5060 2195 5070 2215
rect 5090 2205 5100 2215
rect 5090 2195 5180 2205
rect 5060 2185 5180 2195
rect 4780 2130 4800 2155
rect 5005 2145 5140 2165
rect 4535 2110 4800 2130
rect 4545 2075 4585 2085
rect 4545 2055 4555 2075
rect 4575 2055 4585 2075
rect 4545 2045 4585 2055
rect 4610 2020 4630 2110
rect 4035 2010 4075 2020
rect 4035 1990 4045 2010
rect 4065 1990 4075 2010
rect 4035 1980 4075 1990
rect 4100 2010 4140 2020
rect 4100 1990 4110 2010
rect 4130 1990 4140 2010
rect 4100 1980 4140 1990
rect 4165 2010 4205 2020
rect 4165 1990 4175 2010
rect 4195 1990 4205 2010
rect 4165 1980 4205 1990
rect 4230 2010 4270 2020
rect 4230 1990 4240 2010
rect 4260 1990 4270 2010
rect 4230 1980 4270 1990
rect 4295 2010 4335 2020
rect 4295 1990 4305 2010
rect 4325 1990 4335 2010
rect 4295 1980 4335 1990
rect 4395 2010 4435 2020
rect 4395 1990 4405 2010
rect 4425 1990 4435 2010
rect 4395 1980 4435 1990
rect 4460 2010 4500 2020
rect 4460 1990 4470 2010
rect 4490 1990 4500 2010
rect 4460 1980 4500 1990
rect 4525 2010 4565 2020
rect 4525 1990 4535 2010
rect 4555 1990 4565 2010
rect 4525 1980 4565 1990
rect 4590 2010 4630 2020
rect 4590 1990 4600 2010
rect 4620 1990 4630 2010
rect 4590 1980 4630 1990
rect 4655 2010 4695 2020
rect 4655 1990 4665 2010
rect 4685 1990 4695 2010
rect 4655 1980 4695 1990
rect 4735 2010 4775 2020
rect 4735 1990 4745 2010
rect 4765 1990 4775 2010
rect 4735 1980 4775 1990
rect 4800 2010 4840 2020
rect 4800 1990 4810 2010
rect 4830 1990 4840 2010
rect 4800 1980 4840 1990
rect 4865 2010 4905 2020
rect 4865 1990 4875 2010
rect 4895 1990 4905 2010
rect 4865 1980 4905 1990
rect 4930 2010 4970 2020
rect 4930 1990 4940 2010
rect 4960 1990 4970 2010
rect 4930 1980 4970 1990
rect 4995 2010 5035 2020
rect 4995 1990 5005 2010
rect 5025 1990 5035 2010
rect 4995 1980 5035 1990
rect 4175 1935 4195 1980
rect 4405 1960 4425 1980
rect 4535 1960 4555 1980
rect 4665 1960 4685 1980
rect 4405 1940 4685 1960
rect 4745 1960 4765 1980
rect 4875 1960 4895 1980
rect 5005 1960 5025 1980
rect 4745 1955 5025 1960
rect 4165 1925 4205 1935
rect 4165 1905 4175 1925
rect 4195 1905 4205 1925
rect 4165 1895 4205 1905
rect 4535 1890 4555 1940
rect 4745 1935 5060 1955
rect 4975 1905 5020 1915
rect 4245 1870 4665 1890
rect 4975 1885 4985 1905
rect 5005 1885 5020 1905
rect 4975 1875 5020 1885
rect 4245 1850 4265 1870
rect 4645 1850 4665 1870
rect 4035 1840 4075 1850
rect 3940 1795 3980 1815
rect 4035 1745 4045 1840
rect 4065 1745 4075 1840
rect 4035 1735 4075 1745
rect 4135 1840 4175 1850
rect 4135 1745 4145 1840
rect 4165 1745 4175 1840
rect 4135 1735 4175 1745
rect 4235 1840 4275 1850
rect 4235 1745 4245 1840
rect 4265 1745 4275 1840
rect 4235 1735 4275 1745
rect 4335 1840 4375 1850
rect 4335 1745 4345 1840
rect 4365 1745 4375 1840
rect 4335 1735 4375 1745
rect 4435 1840 4475 1850
rect 4435 1745 4445 1840
rect 4465 1745 4475 1840
rect 4435 1735 4475 1745
rect 4535 1840 4575 1850
rect 4535 1745 4545 1840
rect 4565 1745 4575 1840
rect 4535 1735 4575 1745
rect 4635 1840 4675 1850
rect 4635 1745 4645 1840
rect 4665 1745 4675 1840
rect 4635 1735 4675 1745
rect 4735 1840 4775 1850
rect 4735 1745 4745 1840
rect 4765 1745 4775 1840
rect 4735 1735 4775 1745
rect 4835 1840 4875 1850
rect 4835 1745 4845 1840
rect 4865 1745 4875 1840
rect 4835 1735 4875 1745
rect 4915 1840 4955 1850
rect 4915 1745 4925 1840
rect 4945 1745 4955 1840
rect 4915 1735 4955 1745
rect 4045 1715 4065 1735
rect 4085 1715 4125 1720
rect 4445 1715 4465 1735
rect 4785 1715 4825 1720
rect 4845 1715 4865 1735
rect 4045 1710 4865 1715
rect 4045 1695 4095 1710
rect 4085 1690 4095 1695
rect 4115 1705 4795 1710
rect 4115 1695 4445 1705
rect 4115 1690 4125 1695
rect 4085 1680 4125 1690
rect 4435 1685 4445 1695
rect 4465 1695 4795 1705
rect 4465 1685 4475 1695
rect 4435 1675 4475 1685
rect 4785 1690 4795 1695
rect 4815 1695 4865 1710
rect 4815 1690 4825 1695
rect 4785 1680 4825 1690
rect 3985 1595 4180 1615
rect 5000 1615 5020 1875
rect 4690 1595 5020 1615
rect 3985 1575 4005 1595
rect 5040 1575 5060 1935
rect 3965 1565 4015 1575
rect 3965 1535 3975 1565
rect 4005 1535 4015 1565
rect 3965 1525 4015 1535
rect 4930 1565 5060 1575
rect 4930 1530 4940 1565
rect 4975 1555 5060 1565
rect 4975 1530 4985 1555
rect 4930 1520 4985 1530
rect 5040 1490 5060 1555
rect 5120 1575 5140 2145
rect 5160 1615 5180 2185
rect 5160 1595 5325 1615
rect 5863 1595 6180 1615
rect 6160 1575 6180 1595
rect 5120 1565 5235 1575
rect 5120 1555 5190 1565
rect 5120 1490 5140 1555
rect 5180 1530 5190 1555
rect 5225 1530 5235 1565
rect 5180 1520 5235 1530
rect 6150 1565 6200 1575
rect 6150 1535 6160 1565
rect 6190 1535 6200 1565
rect 6150 1525 6200 1535
rect 5040 1471 5140 1490
rect 5040 1470 5105 1471
<< viali >>
rect 4160 2395 4180 2615
rect 4360 2395 4380 2615
rect 4560 2395 4580 2615
rect 4760 2395 4780 2615
rect 4955 2395 4975 2615
rect 4470 2225 4490 2295
rect 4600 2225 4620 2295
rect 4810 2225 4830 2295
rect 4940 2225 4960 2295
rect 4285 2165 4305 2185
rect 4555 2055 4575 2075
rect 4145 1745 4165 1840
rect 4345 1745 4365 1840
rect 4545 1745 4565 1840
rect 4745 1745 4765 1840
rect 4925 1745 4945 1840
rect 3975 1535 4005 1565
rect 4940 1530 4975 1565
rect 5190 1530 5225 1565
rect 6160 1535 6190 1565
<< metal1 >>
rect 3990 2615 5060 2685
rect 3990 2395 4160 2615
rect 4180 2395 4360 2615
rect 4380 2395 4560 2615
rect 4580 2395 4760 2615
rect 4780 2395 4955 2615
rect 4975 2395 5060 2615
rect 3990 2295 5060 2395
rect 3990 2225 4470 2295
rect 4490 2225 4600 2295
rect 4620 2225 4810 2295
rect 4830 2225 4940 2295
rect 4960 2225 5060 2295
rect 3990 2185 5060 2225
rect 4275 2165 4285 2185
rect 4305 2165 4315 2185
rect 4275 2155 4315 2165
rect 4295 2140 4315 2155
rect 3990 2120 4565 2140
rect 4545 2085 4565 2120
rect 4545 2075 4585 2085
rect 4545 2055 4555 2075
rect 4575 2055 4585 2075
rect 4545 2045 4585 2055
rect 4165 1980 4205 2020
rect 3965 1565 4015 1575
rect 3965 1535 3975 1565
rect 4005 1535 4015 1565
rect 3965 1525 4015 1535
rect 4930 1565 4985 1575
rect 4930 1530 4940 1565
rect 4975 1530 4985 1565
rect 4930 1520 4985 1530
rect 5180 1565 5235 1575
rect 5180 1530 5190 1565
rect 5225 1530 5235 1565
rect 5180 1520 5235 1530
rect 6150 1565 6200 1575
rect 6150 1535 6160 1565
rect 6190 1535 6200 1565
rect 6150 1525 6200 1535
<< via1 >>
rect 3975 1535 4005 1565
rect 4940 1530 4975 1565
rect 5190 1530 5225 1565
rect 6160 1535 6190 1565
<< metal2 >>
rect 3965 1565 4015 1575
rect 3965 1535 3975 1565
rect 4005 1535 4015 1565
rect 3965 1525 4015 1535
rect 4930 1565 4985 1575
rect 4930 1530 4940 1565
rect 4975 1530 4985 1565
rect 4930 1520 4985 1530
rect 5180 1565 5235 1575
rect 5180 1530 5190 1565
rect 5225 1530 5235 1565
rect 5180 1520 5235 1530
rect 6150 1565 6200 1575
rect 6150 1535 6160 1565
rect 6190 1535 6200 1565
rect 6150 1525 6200 1535
<< via2 >>
rect 3975 1535 4005 1565
rect 4940 1530 4975 1565
rect 5190 1530 5225 1565
rect 6160 1535 6190 1565
<< metal3 >>
rect 3965 1565 4015 1575
rect 3965 1535 3975 1565
rect 4005 1535 4015 1565
rect 3965 1525 4015 1535
rect 3970 1400 4015 1525
rect 4930 1565 4985 1575
rect 4930 1530 4940 1565
rect 4975 1530 4985 1565
rect 4930 1520 4985 1530
rect 5180 1565 5235 1575
rect 5180 1530 5190 1565
rect 5225 1530 5235 1565
rect 5180 1520 5235 1530
rect 6150 1565 6200 1575
rect 6150 1535 6160 1565
rect 6190 1535 6200 1565
rect 6150 1525 6200 1535
rect 6150 1400 6195 1525
rect 3970 370 5000 1400
rect 5165 370 6195 1400
<< via3 >>
rect 4940 1530 4975 1565
rect 5190 1530 5225 1565
<< mimcap >>
rect 3985 1375 4985 1385
rect 3985 1340 4940 1375
rect 4975 1340 4985 1375
rect 3985 385 4985 1340
rect 5180 1375 6180 1385
rect 5180 1340 5190 1375
rect 5225 1340 6180 1375
rect 5180 385 6180 1340
<< mimcapcontact >>
rect 4940 1340 4975 1375
rect 5190 1340 5225 1375
<< metal4 >>
rect 4930 1565 4985 1575
rect 4930 1530 4940 1565
rect 4975 1530 4985 1565
rect 4930 1375 4985 1530
rect 4930 1340 4940 1375
rect 4975 1340 4985 1375
rect 4930 1335 4985 1340
rect 5180 1565 5235 1575
rect 5180 1530 5190 1565
rect 5225 1530 5235 1565
rect 5180 1375 5235 1530
rect 5180 1340 5190 1375
rect 5225 1340 5235 1375
rect 5180 1335 5235 1340
<< labels >>
flabel locali 4490 2130 4490 2130 3 FreeSans 160 0 80 0 n_left
flabel locali 4630 2130 4630 2130 3 FreeSans 160 0 80 0 n_right
flabel locali 3940 2545 3940 2545 7 FreeSans 160 0 -80 0 p_bias
flabel locali 4680 2345 4680 2345 4 FreeSans 400 0 0 0 v_common_p
flabel locali 4250 2175 4250 2175 3 FreeSans 160 0 80 0 p_right
<< end >>
