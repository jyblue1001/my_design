magic
tech sky130A
timestamp 1756075196
<< metal1 >>
rect 2070 19310 2190 19325
rect 2070 19280 2115 19310
rect 2145 19280 2190 19310
rect 2070 19245 2190 19280
rect 2070 19215 2115 19245
rect 2145 19215 2190 19245
rect 2070 19175 2190 19215
rect 2070 19145 2115 19175
rect 2145 19145 2190 19175
rect 2070 19105 2190 19145
rect 2070 19075 2115 19105
rect 2145 19075 2190 19105
rect 2070 19035 2190 19075
rect 2070 19005 2115 19035
rect 2145 19005 2190 19035
rect 2070 18970 2190 19005
rect 2070 18940 2115 18970
rect 2145 18940 2190 18970
rect 2070 18910 2190 18940
rect 2070 18880 2115 18910
rect 2145 18880 2190 18910
rect 2070 18845 2190 18880
rect 2070 18815 2115 18845
rect 2145 18815 2190 18845
rect 2070 18775 2190 18815
rect 2070 18745 2115 18775
rect 2145 18745 2190 18775
rect 2070 18705 2190 18745
rect 2070 18675 2115 18705
rect 2145 18675 2190 18705
rect 2070 18635 2190 18675
rect 2070 18605 2115 18635
rect 2145 18605 2190 18635
rect 2070 18570 2190 18605
rect 2070 18540 2115 18570
rect 2145 18540 2190 18570
rect 2070 18510 2190 18540
rect 2070 18480 2115 18510
rect 2145 18480 2190 18510
rect 2070 18445 2190 18480
rect 2070 18415 2115 18445
rect 2145 18415 2190 18445
rect 2070 18375 2190 18415
rect 2070 18345 2115 18375
rect 2145 18345 2190 18375
rect 2070 18305 2190 18345
rect 2070 18275 2115 18305
rect 2145 18275 2190 18305
rect 2070 18235 2190 18275
rect 2070 18205 2115 18235
rect 2145 18205 2190 18235
rect 2070 18170 2190 18205
rect 2070 18140 2115 18170
rect 2145 18140 2190 18170
rect 2070 18110 2190 18140
rect 2070 18080 2115 18110
rect 2145 18080 2190 18110
rect 2070 18045 2190 18080
rect 2070 18015 2115 18045
rect 2145 18015 2190 18045
rect 2070 17975 2190 18015
rect 2070 17945 2115 17975
rect 2145 17945 2190 17975
rect 2070 17905 2190 17945
rect 2070 17875 2115 17905
rect 2145 17875 2190 17905
rect 2070 17835 2190 17875
rect 2070 17805 2115 17835
rect 2145 17805 2190 17835
rect 2070 17770 2190 17805
rect 2070 17740 2115 17770
rect 2145 17740 2190 17770
rect 2070 15690 2190 17740
rect 6690 19310 6750 19325
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2070 15660 2075 15690
rect 2105 15660 2115 15690
rect 2145 15660 2155 15690
rect 2185 15660 2190 15690
rect 2070 15650 2190 15660
rect 2070 15620 2075 15650
rect 2105 15620 2115 15650
rect 2145 15620 2155 15650
rect 2185 15620 2190 15650
rect 2070 15610 2190 15620
rect 2070 15580 2075 15610
rect 2105 15580 2115 15610
rect 2145 15580 2155 15610
rect 2185 15580 2190 15610
rect 2070 12710 2190 15580
rect 2070 12680 2075 12710
rect 2105 12680 2115 12710
rect 2145 12680 2155 12710
rect 2185 12680 2190 12710
rect 2070 12670 2190 12680
rect 2070 12640 2075 12670
rect 2105 12640 2115 12670
rect 2145 12640 2155 12670
rect 2185 12640 2190 12670
rect 2070 12550 2190 12640
rect 2070 12520 2075 12550
rect 2105 12520 2115 12550
rect 2145 12520 2155 12550
rect 2185 12520 2190 12550
rect 2070 12510 2190 12520
rect 2070 12480 2075 12510
rect 2105 12480 2115 12510
rect 2145 12480 2155 12510
rect 2185 12480 2190 12510
rect 2070 12470 2190 12480
rect 2070 12440 2075 12470
rect 2105 12440 2115 12470
rect 2145 12440 2155 12470
rect 2185 12440 2190 12470
rect 2070 12435 2190 12440
rect 2205 15925 2325 15930
rect 2205 15895 2210 15925
rect 2240 15895 2250 15925
rect 2280 15895 2290 15925
rect 2320 15895 2325 15925
rect 1280 9635 1400 9650
rect 1280 9605 1325 9635
rect 1355 9605 1400 9635
rect 1280 9570 1400 9605
rect 1280 9540 1325 9570
rect 1355 9540 1400 9570
rect 1280 9500 1400 9540
rect 1280 9470 1325 9500
rect 1355 9470 1400 9500
rect 1280 9430 1400 9470
rect 1280 9400 1325 9430
rect 1355 9400 1400 9430
rect 1280 9360 1400 9400
rect 1280 9330 1325 9360
rect 1355 9330 1400 9360
rect 1280 9295 1400 9330
rect 1280 9265 1325 9295
rect 1355 9265 1400 9295
rect 1280 9235 1400 9265
rect 1280 9205 1325 9235
rect 1355 9205 1400 9235
rect 1280 9170 1400 9205
rect 1280 9140 1325 9170
rect 1355 9140 1400 9170
rect 1280 9100 1400 9140
rect 1280 9070 1325 9100
rect 1355 9070 1400 9100
rect 1280 9030 1400 9070
rect 1280 9000 1325 9030
rect 1355 9000 1400 9030
rect 1280 8960 1400 9000
rect 1280 8930 1325 8960
rect 1355 8930 1400 8960
rect 1280 8895 1400 8930
rect 1280 8865 1325 8895
rect 1355 8865 1400 8895
rect 1280 8835 1400 8865
rect 1280 8805 1325 8835
rect 1355 8805 1400 8835
rect 1280 8770 1400 8805
rect 1280 8740 1325 8770
rect 1355 8740 1400 8770
rect 1280 8700 1400 8740
rect 1280 8670 1325 8700
rect 1355 8670 1400 8700
rect 1280 8630 1400 8670
rect 1280 8600 1325 8630
rect 1355 8600 1400 8630
rect 1280 8560 1400 8600
rect 1280 8530 1325 8560
rect 1355 8530 1400 8560
rect 1280 8495 1400 8530
rect 1280 8465 1325 8495
rect 1355 8465 1400 8495
rect 1280 8435 1400 8465
rect 1280 8405 1325 8435
rect 1355 8405 1400 8435
rect 1280 8370 1400 8405
rect 1280 8340 1325 8370
rect 1355 8340 1400 8370
rect 1280 8300 1400 8340
rect 1280 8270 1325 8300
rect 1355 8270 1400 8300
rect 1280 8230 1400 8270
rect 1280 8200 1325 8230
rect 1355 8200 1400 8230
rect 1280 8160 1400 8200
rect 1280 8130 1325 8160
rect 1355 8130 1400 8160
rect 1280 7740 1400 8130
rect 2205 9635 2325 15895
rect 6660 15595 6780 17725
rect 6660 15565 6665 15595
rect 6695 15565 6705 15595
rect 6735 15565 6745 15595
rect 6775 15565 6780 15595
rect 6660 15555 6780 15565
rect 6660 15525 6665 15555
rect 6695 15525 6705 15555
rect 6735 15525 6745 15555
rect 6775 15525 6780 15555
rect 6660 15515 6780 15525
rect 6660 15485 6665 15515
rect 6695 15485 6705 15515
rect 6735 15485 6745 15515
rect 6775 15485 6780 15515
rect 2205 9605 2250 9635
rect 2280 9605 2325 9635
rect 2205 9570 2325 9605
rect 2205 9540 2250 9570
rect 2280 9540 2325 9570
rect 2205 9500 2325 9540
rect 2205 9470 2250 9500
rect 2280 9470 2325 9500
rect 2205 9430 2325 9470
rect 2205 9400 2250 9430
rect 2280 9400 2325 9430
rect 2205 9360 2325 9400
rect 2205 9330 2250 9360
rect 2280 9330 2325 9360
rect 2205 9295 2325 9330
rect 2205 9265 2250 9295
rect 2280 9265 2325 9295
rect 2205 9235 2325 9265
rect 2205 9205 2250 9235
rect 2280 9205 2325 9235
rect 2205 9170 2325 9205
rect 2205 9140 2250 9170
rect 2280 9140 2325 9170
rect 2205 9100 2325 9140
rect 2205 9070 2250 9100
rect 2280 9070 2325 9100
rect 2205 9030 2325 9070
rect 2205 9000 2250 9030
rect 2280 9000 2325 9030
rect 2205 8960 2325 9000
rect 2205 8930 2250 8960
rect 2280 8930 2325 8960
rect 2205 8895 2325 8930
rect 2205 8865 2250 8895
rect 2280 8865 2325 8895
rect 2205 8835 2325 8865
rect 2205 8805 2250 8835
rect 2280 8805 2325 8835
rect 2205 8770 2325 8805
rect 2205 8740 2250 8770
rect 2280 8740 2325 8770
rect 2205 8700 2325 8740
rect 2205 8670 2250 8700
rect 2280 8670 2325 8700
rect 2205 8630 2325 8670
rect 2205 8600 2250 8630
rect 2280 8600 2325 8630
rect 2205 8560 2325 8600
rect 2205 8530 2250 8560
rect 2280 8530 2325 8560
rect 2205 8495 2325 8530
rect 2205 8465 2250 8495
rect 2280 8465 2325 8495
rect 2205 8435 2325 8465
rect 2205 8405 2250 8435
rect 2280 8405 2325 8435
rect 2205 8370 2325 8405
rect 2205 8340 2250 8370
rect 2280 8340 2325 8370
rect 2205 8300 2325 8340
rect 2205 8270 2250 8300
rect 2280 8270 2325 8300
rect 2205 8230 2325 8270
rect 2205 8200 2250 8230
rect 2280 8200 2325 8230
rect 2205 8160 2325 8200
rect 2205 8130 2250 8160
rect 2280 8130 2325 8160
rect 2205 8105 2325 8130
rect 1980 8070 2100 8075
rect 1980 8040 1985 8070
rect 2015 8040 2025 8070
rect 2055 8040 2065 8070
rect 2095 8040 2100 8070
rect 1630 8015 1750 8020
rect 1630 7985 1635 8015
rect 1665 7985 1675 8015
rect 1705 7985 1715 8015
rect 1745 7985 1750 8015
rect 1630 7740 1750 7985
rect 1980 7740 2100 8040
rect 2475 8070 2515 13175
rect 2475 8040 2480 8070
rect 2510 8040 2515 8070
rect 2475 8035 2515 8040
rect 2725 7855 2745 9735
rect 2855 7965 2875 9735
rect 3175 9650 3215 10325
rect 3165 9635 3225 9650
rect 3165 9605 3180 9635
rect 3210 9605 3225 9635
rect 3165 9570 3225 9605
rect 3165 9540 3180 9570
rect 3210 9540 3225 9570
rect 3165 9500 3225 9540
rect 3165 9470 3180 9500
rect 3210 9470 3225 9500
rect 3165 9430 3225 9470
rect 3165 9400 3180 9430
rect 3210 9400 3225 9430
rect 3165 9360 3225 9400
rect 3165 9330 3180 9360
rect 3210 9330 3225 9360
rect 3165 9295 3225 9330
rect 3165 9265 3180 9295
rect 3210 9265 3225 9295
rect 3165 9235 3225 9265
rect 3165 9205 3180 9235
rect 3210 9205 3225 9235
rect 3165 9170 3225 9205
rect 3165 9140 3180 9170
rect 3210 9140 3225 9170
rect 3165 9100 3225 9140
rect 3165 9070 3180 9100
rect 3210 9070 3225 9100
rect 3165 9030 3225 9070
rect 3165 9000 3180 9030
rect 3210 9000 3225 9030
rect 3165 8960 3225 9000
rect 3165 8930 3180 8960
rect 3210 8930 3225 8960
rect 3165 8895 3225 8930
rect 3165 8865 3180 8895
rect 3210 8865 3225 8895
rect 3165 8835 3225 8865
rect 3165 8805 3180 8835
rect 3210 8805 3225 8835
rect 3165 8770 3225 8805
rect 3165 8740 3180 8770
rect 3210 8740 3225 8770
rect 3165 8700 3225 8740
rect 3165 8670 3180 8700
rect 3210 8670 3225 8700
rect 3165 8630 3225 8670
rect 3165 8600 3180 8630
rect 3210 8600 3225 8630
rect 3165 8560 3225 8600
rect 3165 8530 3180 8560
rect 3210 8530 3225 8560
rect 3165 8495 3225 8530
rect 3165 8465 3180 8495
rect 3210 8465 3225 8495
rect 3165 8435 3225 8465
rect 3165 8405 3180 8435
rect 3210 8405 3225 8435
rect 3165 8370 3225 8405
rect 3165 8340 3180 8370
rect 3210 8340 3225 8370
rect 3165 8300 3225 8340
rect 3165 8270 3180 8300
rect 3210 8270 3225 8300
rect 3165 8230 3225 8270
rect 3165 8200 3180 8230
rect 3210 8200 3225 8230
rect 3165 8160 3225 8200
rect 3165 8130 3180 8160
rect 3210 8130 3225 8160
rect 3165 8105 3225 8130
rect 2845 7960 2885 7965
rect 2845 7930 2850 7960
rect 2880 7930 2885 7960
rect 2845 7925 2885 7930
rect 3290 7870 3330 10660
rect 3630 8015 3670 10100
rect 3630 7985 3635 8015
rect 3665 7985 3670 8015
rect 3630 7980 3670 7985
rect 3850 8015 3890 10100
rect 3850 7985 3855 8015
rect 3885 7985 3890 8015
rect 3850 7980 3890 7985
rect 3385 7960 3420 7965
rect 3415 7930 3420 7960
rect 3385 7925 3420 7930
rect 2715 7850 2755 7855
rect 2715 7820 2720 7850
rect 2750 7820 2755 7850
rect 2715 7815 2755 7820
rect 3075 7850 3115 7855
rect 3075 7820 3080 7850
rect 3110 7820 3115 7850
rect 3075 7815 3115 7820
rect 3290 7840 3295 7870
rect 3325 7840 3330 7870
rect 3290 7830 3330 7840
rect 930 7735 1050 7740
rect 930 7705 935 7735
rect 965 7705 975 7735
rect 1005 7705 1015 7735
rect 1045 7705 1050 7735
rect 930 7695 1050 7705
rect 930 7665 935 7695
rect 965 7665 975 7695
rect 1005 7665 1015 7695
rect 1045 7665 1050 7695
rect 930 7655 1050 7665
rect 930 7625 935 7655
rect 965 7625 975 7655
rect 1005 7625 1015 7655
rect 1045 7625 1050 7655
rect 930 2690 1050 7625
rect 3085 6625 3105 7815
rect 3290 7800 3295 7830
rect 3325 7800 3330 7830
rect 3290 7790 3330 7800
rect 3290 7760 3295 7790
rect 3325 7760 3330 7790
rect 3290 7755 3330 7760
rect 3075 6620 3115 6625
rect 3075 6590 3080 6620
rect 3110 6590 3115 6620
rect 3075 6585 3115 6590
rect 3390 5340 3410 7925
rect 3435 7870 3475 7875
rect 3435 7840 3440 7870
rect 3470 7840 3475 7870
rect 3435 7830 3475 7840
rect 3435 7800 3440 7830
rect 3470 7800 3475 7830
rect 3435 7790 3475 7800
rect 3435 7760 3440 7790
rect 3470 7760 3475 7790
rect 3380 5335 3420 5340
rect 3380 5305 3385 5335
rect 3415 5305 3420 5335
rect 3380 5300 3420 5305
rect 3435 4655 3475 7760
rect 4310 7735 4340 9735
rect 4310 7695 4340 7705
rect 4310 7655 4340 7665
rect 4310 7620 4340 7625
rect 4420 7735 4450 9735
rect 4420 7695 4450 7705
rect 4420 7655 4450 7665
rect 4420 7620 4450 7625
rect 4530 7735 4560 9735
rect 4530 7695 4560 7705
rect 4530 7655 4560 7665
rect 4530 7620 4560 7625
rect 4640 7735 4670 9735
rect 5090 8015 5130 10100
rect 5090 7985 5095 8015
rect 5125 7985 5130 8015
rect 5090 7980 5130 7985
rect 5310 8015 5350 10100
rect 5310 7985 5315 8015
rect 5345 7985 5350 8015
rect 5310 7980 5350 7985
rect 6155 7965 6175 9740
rect 5470 7960 5510 7965
rect 5470 7930 5475 7960
rect 5505 7930 5510 7960
rect 5470 7925 5510 7930
rect 6145 7960 6185 7965
rect 6145 7930 6150 7960
rect 6180 7930 6185 7960
rect 6145 7925 6185 7930
rect 4640 7695 4670 7705
rect 4640 7655 4670 7665
rect 4640 7620 4670 7625
rect 5480 5400 5500 7925
rect 5545 7870 5585 7875
rect 5545 7840 5550 7870
rect 5580 7840 5585 7870
rect 5545 7830 5585 7840
rect 5545 7800 5550 7830
rect 5580 7800 5585 7830
rect 5545 7790 5585 7800
rect 5545 7760 5550 7790
rect 5580 7760 5585 7790
rect 5475 5395 5505 5400
rect 5475 5360 5505 5365
rect 3435 4625 3440 4655
rect 3470 4625 3475 4655
rect 3435 4620 3475 4625
rect 4470 4655 4510 4660
rect 4470 4625 4475 4655
rect 4505 4625 4510 4655
rect 4470 4435 4510 4625
rect 5545 4655 5585 7760
rect 5870 6965 5910 6970
rect 5870 6935 5875 6965
rect 5905 6935 5910 6965
rect 5620 6565 5660 6570
rect 5620 6535 5625 6565
rect 5655 6535 5660 6565
rect 5620 5970 5660 6535
rect 5870 6565 5910 6935
rect 6220 6965 6260 13120
rect 6465 8070 6505 13175
rect 6660 12925 6780 15485
rect 6660 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6745 12925
rect 6775 12895 6780 12925
rect 6660 12885 6780 12895
rect 6660 12855 6665 12885
rect 6695 12855 6705 12885
rect 6735 12855 6745 12885
rect 6775 12855 6780 12885
rect 6660 12845 6780 12855
rect 6660 12815 6665 12845
rect 6695 12815 6705 12845
rect 6735 12815 6745 12845
rect 6775 12815 6780 12845
rect 6660 12810 6780 12815
rect 6660 12150 6780 12155
rect 6660 12120 6665 12150
rect 6695 12120 6705 12150
rect 6735 12120 6745 12150
rect 6775 12120 6780 12150
rect 6660 12110 6780 12120
rect 6660 12080 6665 12110
rect 6695 12080 6705 12110
rect 6735 12080 6745 12110
rect 6775 12080 6780 12110
rect 6660 12070 6780 12080
rect 6660 12040 6665 12070
rect 6695 12040 6705 12070
rect 6735 12040 6745 12070
rect 6775 12040 6780 12070
rect 6660 11165 6780 12040
rect 6660 11135 6665 11165
rect 6695 11135 6705 11165
rect 6735 11135 6745 11165
rect 6775 11135 6780 11165
rect 6660 11125 6780 11135
rect 6660 11095 6665 11125
rect 6695 11095 6705 11125
rect 6735 11095 6745 11125
rect 6775 11095 6780 11125
rect 6660 11085 6780 11095
rect 6660 11055 6665 11085
rect 6695 11055 6705 11085
rect 6735 11055 6745 11085
rect 6775 11055 6780 11085
rect 6660 10440 6780 11055
rect 6660 10410 6665 10440
rect 6695 10410 6705 10440
rect 6735 10410 6745 10440
rect 6775 10410 6780 10440
rect 6660 10400 6780 10410
rect 6660 10370 6665 10400
rect 6695 10370 6705 10400
rect 6735 10370 6745 10400
rect 6775 10370 6780 10400
rect 6660 10360 6780 10370
rect 6660 10330 6665 10360
rect 6695 10330 6705 10360
rect 6735 10330 6745 10360
rect 6775 10330 6780 10360
rect 6660 10080 6780 10330
rect 6660 10050 6665 10080
rect 6695 10050 6705 10080
rect 6735 10050 6745 10080
rect 6775 10050 6780 10080
rect 6660 10040 6780 10050
rect 6660 10010 6665 10040
rect 6695 10010 6705 10040
rect 6735 10010 6745 10040
rect 6775 10010 6780 10040
rect 6660 10000 6780 10010
rect 6660 9970 6665 10000
rect 6695 9970 6705 10000
rect 6735 9970 6745 10000
rect 6775 9970 6780 10000
rect 6660 9570 6780 9970
rect 6660 9540 6705 9570
rect 6735 9540 6780 9570
rect 6660 9500 6780 9540
rect 6660 9470 6705 9500
rect 6735 9470 6780 9500
rect 6660 9430 6780 9470
rect 6660 9400 6705 9430
rect 6735 9400 6780 9430
rect 6660 9360 6780 9400
rect 6660 9330 6705 9360
rect 6735 9330 6780 9360
rect 6660 9295 6780 9330
rect 6660 9265 6705 9295
rect 6735 9265 6780 9295
rect 6660 9235 6780 9265
rect 6660 9205 6705 9235
rect 6735 9205 6780 9235
rect 6660 9170 6780 9205
rect 6660 9140 6705 9170
rect 6735 9140 6780 9170
rect 6660 9100 6780 9140
rect 6660 9070 6705 9100
rect 6735 9070 6780 9100
rect 6660 9030 6780 9070
rect 6660 9000 6705 9030
rect 6735 9000 6780 9030
rect 6660 8960 6780 9000
rect 6660 8930 6705 8960
rect 6735 8930 6780 8960
rect 6660 8895 6780 8930
rect 6660 8865 6705 8895
rect 6735 8865 6780 8895
rect 6660 8835 6780 8865
rect 6660 8805 6705 8835
rect 6735 8805 6780 8835
rect 6660 8770 6780 8805
rect 6660 8740 6705 8770
rect 6735 8740 6780 8770
rect 6660 8700 6780 8740
rect 6660 8670 6705 8700
rect 6735 8670 6780 8700
rect 6660 8630 6780 8670
rect 6660 8600 6705 8630
rect 6735 8600 6780 8630
rect 6660 8560 6780 8600
rect 6660 8530 6705 8560
rect 6735 8530 6780 8560
rect 6660 8495 6780 8530
rect 6660 8465 6705 8495
rect 6735 8465 6780 8495
rect 6660 8435 6780 8465
rect 6660 8405 6705 8435
rect 6735 8405 6780 8435
rect 6660 8370 6780 8405
rect 6660 8340 6705 8370
rect 6735 8340 6780 8370
rect 6660 8300 6780 8340
rect 6660 8270 6705 8300
rect 6735 8270 6780 8300
rect 6660 8230 6780 8270
rect 6660 8200 6705 8230
rect 6735 8200 6780 8230
rect 6660 8160 6780 8200
rect 6660 8130 6705 8160
rect 6735 8130 6780 8160
rect 6660 8105 6780 8130
rect 7580 9635 7700 9650
rect 7580 9605 7625 9635
rect 7655 9605 7700 9635
rect 7580 9570 7700 9605
rect 7580 9540 7625 9570
rect 7655 9540 7700 9570
rect 7580 9500 7700 9540
rect 7580 9470 7625 9500
rect 7655 9470 7700 9500
rect 7580 9430 7700 9470
rect 7580 9400 7625 9430
rect 7655 9400 7700 9430
rect 7580 9360 7700 9400
rect 7580 9330 7625 9360
rect 7655 9330 7700 9360
rect 7580 9295 7700 9330
rect 7580 9265 7625 9295
rect 7655 9265 7700 9295
rect 7580 9235 7700 9265
rect 7580 9205 7625 9235
rect 7655 9205 7700 9235
rect 7580 9170 7700 9205
rect 7580 9140 7625 9170
rect 7655 9140 7700 9170
rect 7580 9100 7700 9140
rect 7580 9070 7625 9100
rect 7655 9070 7700 9100
rect 7580 9030 7700 9070
rect 7580 9000 7625 9030
rect 7655 9000 7700 9030
rect 7580 8960 7700 9000
rect 7580 8930 7625 8960
rect 7655 8930 7700 8960
rect 7580 8895 7700 8930
rect 7580 8865 7625 8895
rect 7655 8865 7700 8895
rect 7580 8835 7700 8865
rect 7580 8805 7625 8835
rect 7655 8805 7700 8835
rect 7580 8770 7700 8805
rect 7580 8740 7625 8770
rect 7655 8740 7700 8770
rect 7580 8700 7700 8740
rect 7580 8670 7625 8700
rect 7655 8670 7700 8700
rect 7580 8630 7700 8670
rect 7580 8600 7625 8630
rect 7655 8600 7700 8630
rect 7580 8560 7700 8600
rect 7580 8530 7625 8560
rect 7655 8530 7700 8560
rect 7580 8495 7700 8530
rect 7580 8465 7625 8495
rect 7655 8465 7700 8495
rect 7580 8435 7700 8465
rect 7580 8405 7625 8435
rect 7655 8405 7700 8435
rect 7580 8370 7700 8405
rect 7580 8340 7625 8370
rect 7655 8340 7700 8370
rect 7580 8300 7700 8340
rect 7580 8270 7625 8300
rect 7655 8270 7700 8300
rect 7580 8230 7700 8270
rect 7580 8200 7625 8230
rect 7655 8200 7700 8230
rect 7580 8160 7700 8200
rect 7580 8130 7625 8160
rect 7655 8130 7700 8160
rect 6465 8040 6470 8070
rect 6500 8040 6505 8070
rect 6465 8035 6505 8040
rect 6880 8070 7000 8075
rect 6880 8040 6885 8070
rect 6915 8040 6925 8070
rect 6955 8040 6965 8070
rect 6995 8040 7000 8070
rect 6880 7740 7000 8040
rect 7230 8015 7350 8020
rect 7230 7985 7235 8015
rect 7265 7985 7275 8015
rect 7305 7985 7315 8015
rect 7345 7985 7350 8015
rect 7230 7740 7350 7985
rect 7580 7740 7700 8130
rect 6220 6935 6225 6965
rect 6255 6935 6260 6965
rect 6220 6930 6260 6935
rect 7930 7735 8050 7740
rect 7930 7705 7935 7735
rect 7965 7705 7975 7735
rect 8005 7705 8015 7735
rect 8045 7705 8050 7735
rect 7930 7695 8050 7705
rect 7930 7665 7935 7695
rect 7965 7665 7975 7695
rect 8005 7665 8015 7695
rect 8045 7665 8050 7695
rect 7930 7655 8050 7665
rect 7930 7625 7935 7655
rect 7965 7625 7975 7655
rect 8005 7625 8015 7655
rect 8045 7625 8050 7655
rect 5870 6535 5875 6565
rect 5905 6535 5910 6565
rect 5870 6530 5910 6535
rect 5620 5940 5625 5970
rect 5655 5940 5660 5970
rect 5620 5935 5660 5940
rect 5545 4625 5550 4655
rect 5580 4625 5585 4655
rect 5545 4620 5585 4625
rect 4470 4405 4475 4435
rect 4505 4405 4510 4435
rect 4470 4400 4510 4405
rect 930 2660 935 2690
rect 965 2660 975 2690
rect 1005 2660 1015 2690
rect 1045 2660 1050 2690
rect 930 2650 1050 2660
rect 930 2620 935 2650
rect 965 2620 975 2650
rect 1005 2620 1015 2650
rect 1045 2620 1050 2650
rect 930 2610 1050 2620
rect 930 2580 935 2610
rect 965 2580 975 2610
rect 1005 2580 1015 2610
rect 1045 2580 1050 2610
rect 930 2575 1050 2580
rect 4415 2690 4455 2695
rect 4415 2660 4420 2690
rect 4450 2660 4455 2690
rect 4415 2650 4455 2660
rect 4415 2620 4420 2650
rect 4450 2620 4455 2650
rect 4415 2610 4455 2620
rect 4415 2580 4420 2610
rect 4450 2580 4455 2610
rect 4415 2575 4455 2580
rect 4525 2690 4565 2695
rect 4525 2660 4530 2690
rect 4560 2660 4565 2690
rect 4525 2650 4565 2660
rect 4525 2620 4530 2650
rect 4560 2620 4565 2650
rect 4525 2610 4565 2620
rect 4525 2580 4530 2610
rect 4560 2580 4565 2610
rect 4525 2575 4565 2580
rect 7930 2690 8050 7625
rect 7930 2660 7935 2690
rect 7965 2660 7975 2690
rect 8005 2660 8015 2690
rect 8045 2660 8050 2690
rect 7930 2650 8050 2660
rect 7930 2620 7935 2650
rect 7965 2620 7975 2650
rect 8005 2620 8015 2650
rect 8045 2620 8050 2650
rect 7930 2610 8050 2620
rect 7930 2580 7935 2610
rect 7965 2580 7975 2610
rect 8005 2580 8015 2610
rect 8045 2580 8050 2610
rect 7930 2575 8050 2580
rect -120 225 0 320
rect -120 195 -75 225
rect -45 195 0 225
rect -120 160 0 195
rect -120 130 -75 160
rect -45 130 0 160
rect -120 90 0 130
rect -120 60 -75 90
rect -45 60 0 90
rect -120 20 0 60
rect -120 -10 -75 20
rect -45 -10 0 20
rect -120 -50 0 -10
rect -120 -80 -75 -50
rect -45 -80 0 -50
rect -120 -115 0 -80
rect -120 -145 -75 -115
rect -45 -145 0 -115
rect -120 -175 0 -145
rect -120 -205 -75 -175
rect -45 -205 0 -175
rect -120 -240 0 -205
rect -120 -270 -75 -240
rect -45 -270 0 -240
rect -120 -310 0 -270
rect -120 -340 -75 -310
rect -45 -340 0 -310
rect -120 -380 0 -340
rect -120 -410 -75 -380
rect -45 -410 0 -380
rect -120 -450 0 -410
rect -120 -480 -75 -450
rect -45 -480 0 -450
rect -120 -515 0 -480
rect -120 -545 -75 -515
rect -45 -545 0 -515
rect -120 -575 0 -545
rect -120 -605 -75 -575
rect -45 -605 0 -575
rect -120 -640 0 -605
rect -120 -670 -75 -640
rect -45 -670 0 -640
rect -120 -710 0 -670
rect -120 -740 -75 -710
rect -45 -740 0 -710
rect -120 -780 0 -740
rect -120 -810 -75 -780
rect -45 -810 0 -780
rect -120 -850 0 -810
rect -120 -880 -75 -850
rect -45 -880 0 -850
rect -120 -915 0 -880
rect -120 -945 -75 -915
rect -45 -945 0 -915
rect -120 -975 0 -945
rect -120 -1005 -75 -975
rect -45 -1005 0 -975
rect -120 -1040 0 -1005
rect -120 -1070 -75 -1040
rect -45 -1070 0 -1040
rect -120 -1110 0 -1070
rect -120 -1140 -75 -1110
rect -45 -1140 0 -1110
rect -120 -1180 0 -1140
rect -120 -1210 -75 -1180
rect -45 -1210 0 -1180
rect -120 -1250 0 -1210
rect -120 -1280 -75 -1250
rect -45 -1280 0 -1250
rect -120 -1315 0 -1280
rect -120 -1345 -75 -1315
rect -45 -1345 0 -1315
rect -120 -1360 0 -1345
rect 230 225 350 320
rect 230 195 275 225
rect 305 195 350 225
rect 230 160 350 195
rect 230 130 275 160
rect 305 130 350 160
rect 230 90 350 130
rect 230 60 275 90
rect 305 60 350 90
rect 230 20 350 60
rect 230 -10 275 20
rect 305 -10 350 20
rect 230 -50 350 -10
rect 230 -80 275 -50
rect 305 -80 350 -50
rect 230 -115 350 -80
rect 230 -145 275 -115
rect 305 -145 350 -115
rect 230 -175 350 -145
rect 230 -205 275 -175
rect 305 -205 350 -175
rect 230 -240 350 -205
rect 230 -270 275 -240
rect 305 -270 350 -240
rect 230 -310 350 -270
rect 230 -340 275 -310
rect 305 -340 350 -310
rect 230 -380 350 -340
rect 230 -410 275 -380
rect 305 -410 350 -380
rect 230 -450 350 -410
rect 230 -480 275 -450
rect 305 -480 350 -450
rect 230 -515 350 -480
rect 230 -545 275 -515
rect 305 -545 350 -515
rect 230 -575 350 -545
rect 230 -605 275 -575
rect 305 -605 350 -575
rect 230 -640 350 -605
rect 230 -670 275 -640
rect 305 -670 350 -640
rect 230 -710 350 -670
rect 230 -740 275 -710
rect 305 -740 350 -710
rect 230 -780 350 -740
rect 230 -810 275 -780
rect 305 -810 350 -780
rect 230 -850 350 -810
rect 230 -880 275 -850
rect 305 -880 350 -850
rect 230 -915 350 -880
rect 230 -945 275 -915
rect 305 -945 350 -915
rect 230 -975 350 -945
rect 230 -1005 275 -975
rect 305 -1005 350 -975
rect 230 -1040 350 -1005
rect 230 -1070 275 -1040
rect 305 -1070 350 -1040
rect 230 -1110 350 -1070
rect 230 -1140 275 -1110
rect 305 -1140 350 -1110
rect 230 -1180 350 -1140
rect 230 -1210 275 -1180
rect 305 -1210 350 -1180
rect 230 -1250 350 -1210
rect 230 -1280 275 -1250
rect 305 -1280 350 -1250
rect 230 -1315 350 -1280
rect 230 -1345 275 -1315
rect 305 -1345 350 -1315
rect 230 -1360 350 -1345
rect 580 225 700 320
rect 580 195 625 225
rect 655 195 700 225
rect 580 160 700 195
rect 580 130 625 160
rect 655 130 700 160
rect 580 90 700 130
rect 580 60 625 90
rect 655 60 700 90
rect 580 20 700 60
rect 580 -10 625 20
rect 655 -10 700 20
rect 580 -50 700 -10
rect 580 -80 625 -50
rect 655 -80 700 -50
rect 580 -115 700 -80
rect 580 -145 625 -115
rect 655 -145 700 -115
rect 580 -175 700 -145
rect 580 -205 625 -175
rect 655 -205 700 -175
rect 580 -240 700 -205
rect 580 -270 625 -240
rect 655 -270 700 -240
rect 580 -310 700 -270
rect 580 -340 625 -310
rect 655 -340 700 -310
rect 580 -380 700 -340
rect 580 -410 625 -380
rect 655 -410 700 -380
rect 580 -450 700 -410
rect 580 -480 625 -450
rect 655 -480 700 -450
rect 580 -515 700 -480
rect 580 -545 625 -515
rect 655 -545 700 -515
rect 580 -575 700 -545
rect 580 -605 625 -575
rect 655 -605 700 -575
rect 580 -640 700 -605
rect 580 -670 625 -640
rect 655 -670 700 -640
rect 580 -710 700 -670
rect 580 -740 625 -710
rect 655 -740 700 -710
rect 580 -780 700 -740
rect 580 -810 625 -780
rect 655 -810 700 -780
rect 580 -850 700 -810
rect 580 -880 625 -850
rect 655 -880 700 -850
rect 580 -915 700 -880
rect 580 -945 625 -915
rect 655 -945 700 -915
rect 580 -975 700 -945
rect 580 -1005 625 -975
rect 655 -1005 700 -975
rect 580 -1040 700 -1005
rect 580 -1070 625 -1040
rect 655 -1070 700 -1040
rect 580 -1110 700 -1070
rect 580 -1140 625 -1110
rect 655 -1140 700 -1110
rect 580 -1180 700 -1140
rect 580 -1210 625 -1180
rect 655 -1210 700 -1180
rect 580 -1250 700 -1210
rect 580 -1280 625 -1250
rect 655 -1280 700 -1250
rect 580 -1315 700 -1280
rect 580 -1345 625 -1315
rect 655 -1345 700 -1315
rect 580 -1360 700 -1345
rect 930 225 1050 320
rect 930 195 975 225
rect 1005 195 1050 225
rect 930 160 1050 195
rect 930 130 975 160
rect 1005 130 1050 160
rect 930 90 1050 130
rect 930 60 975 90
rect 1005 60 1050 90
rect 930 20 1050 60
rect 930 -10 975 20
rect 1005 -10 1050 20
rect 930 -50 1050 -10
rect 930 -80 975 -50
rect 1005 -80 1050 -50
rect 930 -115 1050 -80
rect 930 -145 975 -115
rect 1005 -145 1050 -115
rect 930 -175 1050 -145
rect 930 -205 975 -175
rect 1005 -205 1050 -175
rect 930 -240 1050 -205
rect 930 -270 975 -240
rect 1005 -270 1050 -240
rect 930 -310 1050 -270
rect 930 -340 975 -310
rect 1005 -340 1050 -310
rect 930 -380 1050 -340
rect 930 -410 975 -380
rect 1005 -410 1050 -380
rect 930 -450 1050 -410
rect 930 -480 975 -450
rect 1005 -480 1050 -450
rect 930 -515 1050 -480
rect 930 -545 975 -515
rect 1005 -545 1050 -515
rect 930 -575 1050 -545
rect 930 -605 975 -575
rect 1005 -605 1050 -575
rect 930 -640 1050 -605
rect 930 -670 975 -640
rect 1005 -670 1050 -640
rect 930 -710 1050 -670
rect 930 -740 975 -710
rect 1005 -740 1050 -710
rect 930 -780 1050 -740
rect 930 -810 975 -780
rect 1005 -810 1050 -780
rect 930 -850 1050 -810
rect 930 -880 975 -850
rect 1005 -880 1050 -850
rect 930 -915 1050 -880
rect 930 -945 975 -915
rect 1005 -945 1050 -915
rect 930 -975 1050 -945
rect 930 -1005 975 -975
rect 1005 -1005 1050 -975
rect 930 -1040 1050 -1005
rect 930 -1070 975 -1040
rect 1005 -1070 1050 -1040
rect 930 -1110 1050 -1070
rect 930 -1140 975 -1110
rect 1005 -1140 1050 -1110
rect 930 -1180 1050 -1140
rect 930 -1210 975 -1180
rect 1005 -1210 1050 -1180
rect 930 -1250 1050 -1210
rect 930 -1280 975 -1250
rect 1005 -1280 1050 -1250
rect 930 -1315 1050 -1280
rect 930 -1345 975 -1315
rect 1005 -1345 1050 -1315
rect 930 -1360 1050 -1345
rect 1280 225 1400 320
rect 1280 195 1325 225
rect 1355 195 1400 225
rect 1280 160 1400 195
rect 1280 130 1325 160
rect 1355 130 1400 160
rect 1280 90 1400 130
rect 1280 60 1325 90
rect 1355 60 1400 90
rect 1280 20 1400 60
rect 1280 -10 1325 20
rect 1355 -10 1400 20
rect 1280 -50 1400 -10
rect 1280 -80 1325 -50
rect 1355 -80 1400 -50
rect 1280 -115 1400 -80
rect 1280 -145 1325 -115
rect 1355 -145 1400 -115
rect 1280 -175 1400 -145
rect 1280 -205 1325 -175
rect 1355 -205 1400 -175
rect 1280 -240 1400 -205
rect 1280 -270 1325 -240
rect 1355 -270 1400 -240
rect 1280 -310 1400 -270
rect 1280 -340 1325 -310
rect 1355 -340 1400 -310
rect 1280 -380 1400 -340
rect 1280 -410 1325 -380
rect 1355 -410 1400 -380
rect 1280 -450 1400 -410
rect 1280 -480 1325 -450
rect 1355 -480 1400 -450
rect 1280 -515 1400 -480
rect 1280 -545 1325 -515
rect 1355 -545 1400 -515
rect 1280 -575 1400 -545
rect 1280 -605 1325 -575
rect 1355 -605 1400 -575
rect 1280 -640 1400 -605
rect 1280 -670 1325 -640
rect 1355 -670 1400 -640
rect 1280 -710 1400 -670
rect 1280 -740 1325 -710
rect 1355 -740 1400 -710
rect 1280 -780 1400 -740
rect 1280 -810 1325 -780
rect 1355 -810 1400 -780
rect 1280 -850 1400 -810
rect 1280 -880 1325 -850
rect 1355 -880 1400 -850
rect 1280 -915 1400 -880
rect 1280 -945 1325 -915
rect 1355 -945 1400 -915
rect 1280 -975 1400 -945
rect 1280 -1005 1325 -975
rect 1355 -1005 1400 -975
rect 1280 -1040 1400 -1005
rect 1280 -1070 1325 -1040
rect 1355 -1070 1400 -1040
rect 1280 -1110 1400 -1070
rect 1280 -1140 1325 -1110
rect 1355 -1140 1400 -1110
rect 1280 -1180 1400 -1140
rect 1280 -1210 1325 -1180
rect 1355 -1210 1400 -1180
rect 1280 -1250 1400 -1210
rect 1280 -1280 1325 -1250
rect 1355 -1280 1400 -1250
rect 1280 -1315 1400 -1280
rect 1280 -1345 1325 -1315
rect 1355 -1345 1400 -1315
rect 1280 -1360 1400 -1345
rect 1630 225 1750 320
rect 1630 195 1675 225
rect 1705 195 1750 225
rect 1630 160 1750 195
rect 1630 130 1675 160
rect 1705 130 1750 160
rect 1630 90 1750 130
rect 1630 60 1675 90
rect 1705 60 1750 90
rect 1630 20 1750 60
rect 1630 -10 1675 20
rect 1705 -10 1750 20
rect 1630 -50 1750 -10
rect 1630 -80 1675 -50
rect 1705 -80 1750 -50
rect 1630 -115 1750 -80
rect 1630 -145 1675 -115
rect 1705 -145 1750 -115
rect 1630 -175 1750 -145
rect 1630 -205 1675 -175
rect 1705 -205 1750 -175
rect 1630 -240 1750 -205
rect 1630 -270 1675 -240
rect 1705 -270 1750 -240
rect 1630 -310 1750 -270
rect 1630 -340 1675 -310
rect 1705 -340 1750 -310
rect 1630 -380 1750 -340
rect 1630 -410 1675 -380
rect 1705 -410 1750 -380
rect 1630 -450 1750 -410
rect 1630 -480 1675 -450
rect 1705 -480 1750 -450
rect 1630 -515 1750 -480
rect 1630 -545 1675 -515
rect 1705 -545 1750 -515
rect 1630 -575 1750 -545
rect 1630 -605 1675 -575
rect 1705 -605 1750 -575
rect 1630 -640 1750 -605
rect 1630 -670 1675 -640
rect 1705 -670 1750 -640
rect 1630 -710 1750 -670
rect 1630 -740 1675 -710
rect 1705 -740 1750 -710
rect 1630 -780 1750 -740
rect 1630 -810 1675 -780
rect 1705 -810 1750 -780
rect 1630 -850 1750 -810
rect 1630 -880 1675 -850
rect 1705 -880 1750 -850
rect 1630 -915 1750 -880
rect 1630 -945 1675 -915
rect 1705 -945 1750 -915
rect 1630 -975 1750 -945
rect 1630 -1005 1675 -975
rect 1705 -1005 1750 -975
rect 1630 -1040 1750 -1005
rect 1630 -1070 1675 -1040
rect 1705 -1070 1750 -1040
rect 1630 -1110 1750 -1070
rect 1630 -1140 1675 -1110
rect 1705 -1140 1750 -1110
rect 1630 -1180 1750 -1140
rect 1630 -1210 1675 -1180
rect 1705 -1210 1750 -1180
rect 1630 -1250 1750 -1210
rect 1630 -1280 1675 -1250
rect 1705 -1280 1750 -1250
rect 1630 -1315 1750 -1280
rect 1630 -1345 1675 -1315
rect 1705 -1345 1750 -1315
rect 1630 -1360 1750 -1345
rect 1980 225 2100 320
rect 1980 195 2025 225
rect 2055 195 2100 225
rect 1980 160 2100 195
rect 1980 130 2025 160
rect 2055 130 2100 160
rect 1980 90 2100 130
rect 1980 60 2025 90
rect 2055 60 2100 90
rect 1980 20 2100 60
rect 1980 -10 2025 20
rect 2055 -10 2100 20
rect 1980 -50 2100 -10
rect 1980 -80 2025 -50
rect 2055 -80 2100 -50
rect 1980 -115 2100 -80
rect 1980 -145 2025 -115
rect 2055 -145 2100 -115
rect 1980 -175 2100 -145
rect 1980 -205 2025 -175
rect 2055 -205 2100 -175
rect 1980 -240 2100 -205
rect 1980 -270 2025 -240
rect 2055 -270 2100 -240
rect 1980 -310 2100 -270
rect 1980 -340 2025 -310
rect 2055 -340 2100 -310
rect 1980 -380 2100 -340
rect 1980 -410 2025 -380
rect 2055 -410 2100 -380
rect 1980 -450 2100 -410
rect 1980 -480 2025 -450
rect 2055 -480 2100 -450
rect 1980 -515 2100 -480
rect 1980 -545 2025 -515
rect 2055 -545 2100 -515
rect 1980 -575 2100 -545
rect 1980 -605 2025 -575
rect 2055 -605 2100 -575
rect 1980 -640 2100 -605
rect 1980 -670 2025 -640
rect 2055 -670 2100 -640
rect 1980 -710 2100 -670
rect 1980 -740 2025 -710
rect 2055 -740 2100 -710
rect 1980 -780 2100 -740
rect 1980 -810 2025 -780
rect 2055 -810 2100 -780
rect 1980 -850 2100 -810
rect 1980 -880 2025 -850
rect 2055 -880 2100 -850
rect 1980 -915 2100 -880
rect 1980 -945 2025 -915
rect 2055 -945 2100 -915
rect 1980 -975 2100 -945
rect 1980 -1005 2025 -975
rect 2055 -1005 2100 -975
rect 1980 -1040 2100 -1005
rect 1980 -1070 2025 -1040
rect 2055 -1070 2100 -1040
rect 1980 -1110 2100 -1070
rect 1980 -1140 2025 -1110
rect 2055 -1140 2100 -1110
rect 1980 -1180 2100 -1140
rect 1980 -1210 2025 -1180
rect 2055 -1210 2100 -1180
rect 1980 -1250 2100 -1210
rect 1980 -1280 2025 -1250
rect 2055 -1280 2100 -1250
rect 1980 -1315 2100 -1280
rect 1980 -1345 2025 -1315
rect 2055 -1345 2100 -1315
rect 1980 -1360 2100 -1345
rect 2330 225 2450 320
rect 2330 195 2375 225
rect 2405 195 2450 225
rect 2330 160 2450 195
rect 2330 130 2375 160
rect 2405 130 2450 160
rect 2330 90 2450 130
rect 2330 60 2375 90
rect 2405 60 2450 90
rect 2330 20 2450 60
rect 2330 -10 2375 20
rect 2405 -10 2450 20
rect 2330 -50 2450 -10
rect 2330 -80 2375 -50
rect 2405 -80 2450 -50
rect 2330 -115 2450 -80
rect 2330 -145 2375 -115
rect 2405 -145 2450 -115
rect 2330 -175 2450 -145
rect 2330 -205 2375 -175
rect 2405 -205 2450 -175
rect 2330 -240 2450 -205
rect 2330 -270 2375 -240
rect 2405 -270 2450 -240
rect 2330 -310 2450 -270
rect 2330 -340 2375 -310
rect 2405 -340 2450 -310
rect 2330 -380 2450 -340
rect 2330 -410 2375 -380
rect 2405 -410 2450 -380
rect 2330 -450 2450 -410
rect 2330 -480 2375 -450
rect 2405 -480 2450 -450
rect 2330 -515 2450 -480
rect 2330 -545 2375 -515
rect 2405 -545 2450 -515
rect 2330 -575 2450 -545
rect 2330 -605 2375 -575
rect 2405 -605 2450 -575
rect 2330 -640 2450 -605
rect 2330 -670 2375 -640
rect 2405 -670 2450 -640
rect 2330 -710 2450 -670
rect 2330 -740 2375 -710
rect 2405 -740 2450 -710
rect 2330 -780 2450 -740
rect 2330 -810 2375 -780
rect 2405 -810 2450 -780
rect 2330 -850 2450 -810
rect 2330 -880 2375 -850
rect 2405 -880 2450 -850
rect 2330 -915 2450 -880
rect 2330 -945 2375 -915
rect 2405 -945 2450 -915
rect 2330 -975 2450 -945
rect 2330 -1005 2375 -975
rect 2405 -1005 2450 -975
rect 2330 -1040 2450 -1005
rect 2330 -1070 2375 -1040
rect 2405 -1070 2450 -1040
rect 2330 -1110 2450 -1070
rect 2330 -1140 2375 -1110
rect 2405 -1140 2450 -1110
rect 2330 -1180 2450 -1140
rect 2330 -1210 2375 -1180
rect 2405 -1210 2450 -1180
rect 2330 -1250 2450 -1210
rect 2330 -1280 2375 -1250
rect 2405 -1280 2450 -1250
rect 2330 -1315 2450 -1280
rect 2330 -1345 2375 -1315
rect 2405 -1345 2450 -1315
rect 2330 -1360 2450 -1345
rect 2680 225 2800 320
rect 2680 195 2725 225
rect 2755 195 2800 225
rect 2680 160 2800 195
rect 2680 130 2725 160
rect 2755 130 2800 160
rect 2680 90 2800 130
rect 2680 60 2725 90
rect 2755 60 2800 90
rect 2680 20 2800 60
rect 2680 -10 2725 20
rect 2755 -10 2800 20
rect 2680 -50 2800 -10
rect 2680 -80 2725 -50
rect 2755 -80 2800 -50
rect 2680 -115 2800 -80
rect 2680 -145 2725 -115
rect 2755 -145 2800 -115
rect 2680 -175 2800 -145
rect 2680 -205 2725 -175
rect 2755 -205 2800 -175
rect 2680 -240 2800 -205
rect 2680 -270 2725 -240
rect 2755 -270 2800 -240
rect 2680 -310 2800 -270
rect 2680 -340 2725 -310
rect 2755 -340 2800 -310
rect 2680 -380 2800 -340
rect 2680 -410 2725 -380
rect 2755 -410 2800 -380
rect 2680 -450 2800 -410
rect 2680 -480 2725 -450
rect 2755 -480 2800 -450
rect 2680 -515 2800 -480
rect 2680 -545 2725 -515
rect 2755 -545 2800 -515
rect 2680 -575 2800 -545
rect 2680 -605 2725 -575
rect 2755 -605 2800 -575
rect 2680 -640 2800 -605
rect 2680 -670 2725 -640
rect 2755 -670 2800 -640
rect 2680 -710 2800 -670
rect 2680 -740 2725 -710
rect 2755 -740 2800 -710
rect 2680 -780 2800 -740
rect 2680 -810 2725 -780
rect 2755 -810 2800 -780
rect 2680 -850 2800 -810
rect 2680 -880 2725 -850
rect 2755 -880 2800 -850
rect 2680 -915 2800 -880
rect 2680 -945 2725 -915
rect 2755 -945 2800 -915
rect 2680 -975 2800 -945
rect 2680 -1005 2725 -975
rect 2755 -1005 2800 -975
rect 2680 -1040 2800 -1005
rect 2680 -1070 2725 -1040
rect 2755 -1070 2800 -1040
rect 2680 -1110 2800 -1070
rect 2680 -1140 2725 -1110
rect 2755 -1140 2800 -1110
rect 2680 -1180 2800 -1140
rect 2680 -1210 2725 -1180
rect 2755 -1210 2800 -1180
rect 2680 -1250 2800 -1210
rect 2680 -1280 2725 -1250
rect 2755 -1280 2800 -1250
rect 2680 -1315 2800 -1280
rect 2680 -1345 2725 -1315
rect 2755 -1345 2800 -1315
rect 2680 -1360 2800 -1345
rect 3030 225 3150 320
rect 3030 195 3075 225
rect 3105 195 3150 225
rect 3030 160 3150 195
rect 3030 130 3075 160
rect 3105 130 3150 160
rect 3030 90 3150 130
rect 3030 60 3075 90
rect 3105 60 3150 90
rect 3030 20 3150 60
rect 3030 -10 3075 20
rect 3105 -10 3150 20
rect 3030 -50 3150 -10
rect 3030 -80 3075 -50
rect 3105 -80 3150 -50
rect 3030 -115 3150 -80
rect 3030 -145 3075 -115
rect 3105 -145 3150 -115
rect 3030 -175 3150 -145
rect 3030 -205 3075 -175
rect 3105 -205 3150 -175
rect 3030 -240 3150 -205
rect 3030 -270 3075 -240
rect 3105 -270 3150 -240
rect 3030 -310 3150 -270
rect 3030 -340 3075 -310
rect 3105 -340 3150 -310
rect 3030 -380 3150 -340
rect 3030 -410 3075 -380
rect 3105 -410 3150 -380
rect 3030 -450 3150 -410
rect 3030 -480 3075 -450
rect 3105 -480 3150 -450
rect 3030 -515 3150 -480
rect 3030 -545 3075 -515
rect 3105 -545 3150 -515
rect 3030 -575 3150 -545
rect 3030 -605 3075 -575
rect 3105 -605 3150 -575
rect 3030 -640 3150 -605
rect 3030 -670 3075 -640
rect 3105 -670 3150 -640
rect 3030 -710 3150 -670
rect 3030 -740 3075 -710
rect 3105 -740 3150 -710
rect 3030 -780 3150 -740
rect 3030 -810 3075 -780
rect 3105 -810 3150 -780
rect 3030 -850 3150 -810
rect 3030 -880 3075 -850
rect 3105 -880 3150 -850
rect 3030 -915 3150 -880
rect 3030 -945 3075 -915
rect 3105 -945 3150 -915
rect 3030 -975 3150 -945
rect 3030 -1005 3075 -975
rect 3105 -1005 3150 -975
rect 3030 -1040 3150 -1005
rect 3030 -1070 3075 -1040
rect 3105 -1070 3150 -1040
rect 3030 -1110 3150 -1070
rect 3030 -1140 3075 -1110
rect 3105 -1140 3150 -1110
rect 3030 -1180 3150 -1140
rect 3030 -1210 3075 -1180
rect 3105 -1210 3150 -1180
rect 3030 -1250 3150 -1210
rect 3030 -1280 3075 -1250
rect 3105 -1280 3150 -1250
rect 3030 -1315 3150 -1280
rect 3030 -1345 3075 -1315
rect 3105 -1345 3150 -1315
rect 3030 -1360 3150 -1345
rect 3380 225 3500 295
rect 3380 195 3425 225
rect 3455 195 3500 225
rect 3380 160 3500 195
rect 3380 130 3425 160
rect 3455 130 3500 160
rect 3380 90 3500 130
rect 3380 60 3425 90
rect 3455 60 3500 90
rect 3380 20 3500 60
rect 3380 -10 3425 20
rect 3455 -10 3500 20
rect 3380 -50 3500 -10
rect 3380 -80 3425 -50
rect 3455 -80 3500 -50
rect 3380 -115 3500 -80
rect 3380 -145 3425 -115
rect 3455 -145 3500 -115
rect 3380 -175 3500 -145
rect 3380 -205 3425 -175
rect 3455 -205 3500 -175
rect 3380 -240 3500 -205
rect 3380 -270 3425 -240
rect 3455 -270 3500 -240
rect 3380 -310 3500 -270
rect 3380 -340 3425 -310
rect 3455 -340 3500 -310
rect 3380 -380 3500 -340
rect 3380 -410 3425 -380
rect 3455 -410 3500 -380
rect 3380 -450 3500 -410
rect 3380 -480 3425 -450
rect 3455 -480 3500 -450
rect 3380 -515 3500 -480
rect 3380 -545 3425 -515
rect 3455 -545 3500 -515
rect 3380 -575 3500 -545
rect 3380 -605 3425 -575
rect 3455 -605 3500 -575
rect 3380 -640 3500 -605
rect 3380 -670 3425 -640
rect 3455 -670 3500 -640
rect 3380 -710 3500 -670
rect 3380 -740 3425 -710
rect 3455 -740 3500 -710
rect 3380 -780 3500 -740
rect 3380 -810 3425 -780
rect 3455 -810 3500 -780
rect 3380 -850 3500 -810
rect 3380 -880 3425 -850
rect 3455 -880 3500 -850
rect 3380 -915 3500 -880
rect 3380 -945 3425 -915
rect 3455 -945 3500 -915
rect 3380 -975 3500 -945
rect 3380 -1005 3425 -975
rect 3455 -1005 3500 -975
rect 3380 -1040 3500 -1005
rect 3380 -1070 3425 -1040
rect 3455 -1070 3500 -1040
rect 3380 -1110 3500 -1070
rect 3380 -1140 3425 -1110
rect 3455 -1140 3500 -1110
rect 3380 -1180 3500 -1140
rect 3380 -1210 3425 -1180
rect 3455 -1210 3500 -1180
rect 3380 -1250 3500 -1210
rect 3380 -1280 3425 -1250
rect 3455 -1280 3500 -1250
rect 3380 -1315 3500 -1280
rect 3380 -1345 3425 -1315
rect 3455 -1345 3500 -1315
rect 3380 -1360 3500 -1345
rect 3730 225 3850 295
rect 3730 195 3775 225
rect 3805 195 3850 225
rect 3730 160 3850 195
rect 3730 130 3775 160
rect 3805 130 3850 160
rect 3730 90 3850 130
rect 3730 60 3775 90
rect 3805 60 3850 90
rect 3730 20 3850 60
rect 3730 -10 3775 20
rect 3805 -10 3850 20
rect 3730 -50 3850 -10
rect 3730 -80 3775 -50
rect 3805 -80 3850 -50
rect 3730 -115 3850 -80
rect 3730 -145 3775 -115
rect 3805 -145 3850 -115
rect 3730 -175 3850 -145
rect 3730 -205 3775 -175
rect 3805 -205 3850 -175
rect 3730 -240 3850 -205
rect 3730 -270 3775 -240
rect 3805 -270 3850 -240
rect 3730 -310 3850 -270
rect 3730 -340 3775 -310
rect 3805 -340 3850 -310
rect 3730 -380 3850 -340
rect 3730 -410 3775 -380
rect 3805 -410 3850 -380
rect 3730 -450 3850 -410
rect 3730 -480 3775 -450
rect 3805 -480 3850 -450
rect 3730 -515 3850 -480
rect 3730 -545 3775 -515
rect 3805 -545 3850 -515
rect 3730 -575 3850 -545
rect 3730 -605 3775 -575
rect 3805 -605 3850 -575
rect 3730 -640 3850 -605
rect 3730 -670 3775 -640
rect 3805 -670 3850 -640
rect 3730 -710 3850 -670
rect 3730 -740 3775 -710
rect 3805 -740 3850 -710
rect 3730 -780 3850 -740
rect 3730 -810 3775 -780
rect 3805 -810 3850 -780
rect 3730 -850 3850 -810
rect 3730 -880 3775 -850
rect 3805 -880 3850 -850
rect 3730 -915 3850 -880
rect 3730 -945 3775 -915
rect 3805 -945 3850 -915
rect 3730 -975 3850 -945
rect 3730 -1005 3775 -975
rect 3805 -1005 3850 -975
rect 3730 -1040 3850 -1005
rect 3730 -1070 3775 -1040
rect 3805 -1070 3850 -1040
rect 3730 -1110 3850 -1070
rect 3730 -1140 3775 -1110
rect 3805 -1140 3850 -1110
rect 3730 -1180 3850 -1140
rect 3730 -1210 3775 -1180
rect 3805 -1210 3850 -1180
rect 3730 -1250 3850 -1210
rect 3730 -1280 3775 -1250
rect 3805 -1280 3850 -1250
rect 3730 -1315 3850 -1280
rect 3730 -1345 3775 -1315
rect 3805 -1345 3850 -1315
rect 3730 -1360 3850 -1345
rect 4080 225 4200 295
rect 4080 195 4125 225
rect 4155 195 4200 225
rect 4080 160 4200 195
rect 4080 130 4125 160
rect 4155 130 4200 160
rect 4080 90 4200 130
rect 4080 60 4125 90
rect 4155 60 4200 90
rect 4080 20 4200 60
rect 4080 -10 4125 20
rect 4155 -10 4200 20
rect 4080 -50 4200 -10
rect 4080 -80 4125 -50
rect 4155 -80 4200 -50
rect 4080 -115 4200 -80
rect 4080 -145 4125 -115
rect 4155 -145 4200 -115
rect 4080 -175 4200 -145
rect 4080 -205 4125 -175
rect 4155 -205 4200 -175
rect 4080 -240 4200 -205
rect 4080 -270 4125 -240
rect 4155 -270 4200 -240
rect 4080 -310 4200 -270
rect 4080 -340 4125 -310
rect 4155 -340 4200 -310
rect 4080 -380 4200 -340
rect 4080 -410 4125 -380
rect 4155 -410 4200 -380
rect 4080 -450 4200 -410
rect 4080 -480 4125 -450
rect 4155 -480 4200 -450
rect 4080 -515 4200 -480
rect 4080 -545 4125 -515
rect 4155 -545 4200 -515
rect 4080 -575 4200 -545
rect 4080 -605 4125 -575
rect 4155 -605 4200 -575
rect 4080 -640 4200 -605
rect 4080 -670 4125 -640
rect 4155 -670 4200 -640
rect 4080 -710 4200 -670
rect 4080 -740 4125 -710
rect 4155 -740 4200 -710
rect 4080 -780 4200 -740
rect 4080 -810 4125 -780
rect 4155 -810 4200 -780
rect 4080 -850 4200 -810
rect 4080 -880 4125 -850
rect 4155 -880 4200 -850
rect 4080 -915 4200 -880
rect 4080 -945 4125 -915
rect 4155 -945 4200 -915
rect 4080 -975 4200 -945
rect 4080 -1005 4125 -975
rect 4155 -1005 4200 -975
rect 4080 -1040 4200 -1005
rect 4080 -1070 4125 -1040
rect 4155 -1070 4200 -1040
rect 4080 -1110 4200 -1070
rect 4080 -1140 4125 -1110
rect 4155 -1140 4200 -1110
rect 4080 -1180 4200 -1140
rect 4080 -1210 4125 -1180
rect 4155 -1210 4200 -1180
rect 4080 -1250 4200 -1210
rect 4080 -1280 4125 -1250
rect 4155 -1280 4200 -1250
rect 4080 -1315 4200 -1280
rect 4080 -1345 4125 -1315
rect 4155 -1345 4200 -1315
rect 4080 -1360 4200 -1345
rect 4430 225 4550 295
rect 4430 195 4475 225
rect 4505 195 4550 225
rect 4430 160 4550 195
rect 4430 130 4475 160
rect 4505 130 4550 160
rect 4430 90 4550 130
rect 4430 60 4475 90
rect 4505 60 4550 90
rect 4430 20 4550 60
rect 4430 -10 4475 20
rect 4505 -10 4550 20
rect 4430 -50 4550 -10
rect 4430 -80 4475 -50
rect 4505 -80 4550 -50
rect 4430 -115 4550 -80
rect 4430 -145 4475 -115
rect 4505 -145 4550 -115
rect 4430 -175 4550 -145
rect 4430 -205 4475 -175
rect 4505 -205 4550 -175
rect 4430 -240 4550 -205
rect 4430 -270 4475 -240
rect 4505 -270 4550 -240
rect 4430 -310 4550 -270
rect 4430 -340 4475 -310
rect 4505 -340 4550 -310
rect 4430 -380 4550 -340
rect 4430 -410 4475 -380
rect 4505 -410 4550 -380
rect 4430 -450 4550 -410
rect 4430 -480 4475 -450
rect 4505 -480 4550 -450
rect 4430 -515 4550 -480
rect 4430 -545 4475 -515
rect 4505 -545 4550 -515
rect 4430 -575 4550 -545
rect 4430 -605 4475 -575
rect 4505 -605 4550 -575
rect 4430 -640 4550 -605
rect 4430 -670 4475 -640
rect 4505 -670 4550 -640
rect 4430 -710 4550 -670
rect 4430 -740 4475 -710
rect 4505 -740 4550 -710
rect 4430 -780 4550 -740
rect 4430 -810 4475 -780
rect 4505 -810 4550 -780
rect 4430 -850 4550 -810
rect 4430 -880 4475 -850
rect 4505 -880 4550 -850
rect 4430 -915 4550 -880
rect 4430 -945 4475 -915
rect 4505 -945 4550 -915
rect 4430 -975 4550 -945
rect 4430 -1005 4475 -975
rect 4505 -1005 4550 -975
rect 4430 -1040 4550 -1005
rect 4430 -1070 4475 -1040
rect 4505 -1070 4550 -1040
rect 4430 -1110 4550 -1070
rect 4430 -1140 4475 -1110
rect 4505 -1140 4550 -1110
rect 4430 -1180 4550 -1140
rect 4430 -1210 4475 -1180
rect 4505 -1210 4550 -1180
rect 4430 -1250 4550 -1210
rect 4430 -1280 4475 -1250
rect 4505 -1280 4550 -1250
rect 4430 -1315 4550 -1280
rect 4430 -1345 4475 -1315
rect 4505 -1345 4550 -1315
rect 4430 -1360 4550 -1345
rect 4780 225 4900 295
rect 4780 195 4825 225
rect 4855 195 4900 225
rect 4780 160 4900 195
rect 4780 130 4825 160
rect 4855 130 4900 160
rect 4780 90 4900 130
rect 4780 60 4825 90
rect 4855 60 4900 90
rect 4780 20 4900 60
rect 4780 -10 4825 20
rect 4855 -10 4900 20
rect 4780 -50 4900 -10
rect 4780 -80 4825 -50
rect 4855 -80 4900 -50
rect 4780 -115 4900 -80
rect 4780 -145 4825 -115
rect 4855 -145 4900 -115
rect 4780 -175 4900 -145
rect 4780 -205 4825 -175
rect 4855 -205 4900 -175
rect 4780 -240 4900 -205
rect 4780 -270 4825 -240
rect 4855 -270 4900 -240
rect 4780 -310 4900 -270
rect 4780 -340 4825 -310
rect 4855 -340 4900 -310
rect 4780 -380 4900 -340
rect 4780 -410 4825 -380
rect 4855 -410 4900 -380
rect 4780 -450 4900 -410
rect 4780 -480 4825 -450
rect 4855 -480 4900 -450
rect 4780 -515 4900 -480
rect 4780 -545 4825 -515
rect 4855 -545 4900 -515
rect 4780 -575 4900 -545
rect 4780 -605 4825 -575
rect 4855 -605 4900 -575
rect 4780 -640 4900 -605
rect 4780 -670 4825 -640
rect 4855 -670 4900 -640
rect 4780 -710 4900 -670
rect 4780 -740 4825 -710
rect 4855 -740 4900 -710
rect 4780 -780 4900 -740
rect 4780 -810 4825 -780
rect 4855 -810 4900 -780
rect 4780 -850 4900 -810
rect 4780 -880 4825 -850
rect 4855 -880 4900 -850
rect 4780 -915 4900 -880
rect 4780 -945 4825 -915
rect 4855 -945 4900 -915
rect 4780 -975 4900 -945
rect 4780 -1005 4825 -975
rect 4855 -1005 4900 -975
rect 4780 -1040 4900 -1005
rect 4780 -1070 4825 -1040
rect 4855 -1070 4900 -1040
rect 4780 -1110 4900 -1070
rect 4780 -1140 4825 -1110
rect 4855 -1140 4900 -1110
rect 4780 -1180 4900 -1140
rect 4780 -1210 4825 -1180
rect 4855 -1210 4900 -1180
rect 4780 -1250 4900 -1210
rect 4780 -1280 4825 -1250
rect 4855 -1280 4900 -1250
rect 4780 -1315 4900 -1280
rect 4780 -1345 4825 -1315
rect 4855 -1345 4900 -1315
rect 4780 -1360 4900 -1345
rect 5130 225 5250 295
rect 5130 195 5175 225
rect 5205 195 5250 225
rect 5130 160 5250 195
rect 5130 130 5175 160
rect 5205 130 5250 160
rect 5130 90 5250 130
rect 5130 60 5175 90
rect 5205 60 5250 90
rect 5130 20 5250 60
rect 5130 -10 5175 20
rect 5205 -10 5250 20
rect 5130 -50 5250 -10
rect 5130 -80 5175 -50
rect 5205 -80 5250 -50
rect 5130 -115 5250 -80
rect 5130 -145 5175 -115
rect 5205 -145 5250 -115
rect 5130 -175 5250 -145
rect 5130 -205 5175 -175
rect 5205 -205 5250 -175
rect 5130 -240 5250 -205
rect 5130 -270 5175 -240
rect 5205 -270 5250 -240
rect 5130 -310 5250 -270
rect 5130 -340 5175 -310
rect 5205 -340 5250 -310
rect 5130 -380 5250 -340
rect 5130 -410 5175 -380
rect 5205 -410 5250 -380
rect 5130 -450 5250 -410
rect 5130 -480 5175 -450
rect 5205 -480 5250 -450
rect 5130 -515 5250 -480
rect 5130 -545 5175 -515
rect 5205 -545 5250 -515
rect 5130 -575 5250 -545
rect 5130 -605 5175 -575
rect 5205 -605 5250 -575
rect 5130 -640 5250 -605
rect 5130 -670 5175 -640
rect 5205 -670 5250 -640
rect 5130 -710 5250 -670
rect 5130 -740 5175 -710
rect 5205 -740 5250 -710
rect 5130 -780 5250 -740
rect 5130 -810 5175 -780
rect 5205 -810 5250 -780
rect 5130 -850 5250 -810
rect 5130 -880 5175 -850
rect 5205 -880 5250 -850
rect 5130 -915 5250 -880
rect 5130 -945 5175 -915
rect 5205 -945 5250 -915
rect 5130 -975 5250 -945
rect 5130 -1005 5175 -975
rect 5205 -1005 5250 -975
rect 5130 -1040 5250 -1005
rect 5130 -1070 5175 -1040
rect 5205 -1070 5250 -1040
rect 5130 -1110 5250 -1070
rect 5130 -1140 5175 -1110
rect 5205 -1140 5250 -1110
rect 5130 -1180 5250 -1140
rect 5130 -1210 5175 -1180
rect 5205 -1210 5250 -1180
rect 5130 -1250 5250 -1210
rect 5130 -1280 5175 -1250
rect 5205 -1280 5250 -1250
rect 5130 -1315 5250 -1280
rect 5130 -1345 5175 -1315
rect 5205 -1345 5250 -1315
rect 5130 -1360 5250 -1345
rect 5480 225 5600 295
rect 5480 195 5525 225
rect 5555 195 5600 225
rect 5480 160 5600 195
rect 5480 130 5525 160
rect 5555 130 5600 160
rect 5480 90 5600 130
rect 5480 60 5525 90
rect 5555 60 5600 90
rect 5480 20 5600 60
rect 5480 -10 5525 20
rect 5555 -10 5600 20
rect 5480 -50 5600 -10
rect 5480 -80 5525 -50
rect 5555 -80 5600 -50
rect 5480 -115 5600 -80
rect 5480 -145 5525 -115
rect 5555 -145 5600 -115
rect 5480 -175 5600 -145
rect 5480 -205 5525 -175
rect 5555 -205 5600 -175
rect 5480 -240 5600 -205
rect 5480 -270 5525 -240
rect 5555 -270 5600 -240
rect 5480 -310 5600 -270
rect 5480 -340 5525 -310
rect 5555 -340 5600 -310
rect 5480 -380 5600 -340
rect 5480 -410 5525 -380
rect 5555 -410 5600 -380
rect 5480 -450 5600 -410
rect 5480 -480 5525 -450
rect 5555 -480 5600 -450
rect 5480 -515 5600 -480
rect 5480 -545 5525 -515
rect 5555 -545 5600 -515
rect 5480 -575 5600 -545
rect 5480 -605 5525 -575
rect 5555 -605 5600 -575
rect 5480 -640 5600 -605
rect 5480 -670 5525 -640
rect 5555 -670 5600 -640
rect 5480 -710 5600 -670
rect 5480 -740 5525 -710
rect 5555 -740 5600 -710
rect 5480 -780 5600 -740
rect 5480 -810 5525 -780
rect 5555 -810 5600 -780
rect 5480 -850 5600 -810
rect 5480 -880 5525 -850
rect 5555 -880 5600 -850
rect 5480 -915 5600 -880
rect 5480 -945 5525 -915
rect 5555 -945 5600 -915
rect 5480 -975 5600 -945
rect 5480 -1005 5525 -975
rect 5555 -1005 5600 -975
rect 5480 -1040 5600 -1005
rect 5480 -1070 5525 -1040
rect 5555 -1070 5600 -1040
rect 5480 -1110 5600 -1070
rect 5480 -1140 5525 -1110
rect 5555 -1140 5600 -1110
rect 5480 -1180 5600 -1140
rect 5480 -1210 5525 -1180
rect 5555 -1210 5600 -1180
rect 5480 -1250 5600 -1210
rect 5480 -1280 5525 -1250
rect 5555 -1280 5600 -1250
rect 5480 -1315 5600 -1280
rect 5480 -1345 5525 -1315
rect 5555 -1345 5600 -1315
rect 5480 -1360 5600 -1345
rect 5830 225 5950 320
rect 5830 195 5875 225
rect 5905 195 5950 225
rect 5830 160 5950 195
rect 5830 130 5875 160
rect 5905 130 5950 160
rect 5830 90 5950 130
rect 5830 60 5875 90
rect 5905 60 5950 90
rect 5830 20 5950 60
rect 5830 -10 5875 20
rect 5905 -10 5950 20
rect 5830 -50 5950 -10
rect 5830 -80 5875 -50
rect 5905 -80 5950 -50
rect 5830 -115 5950 -80
rect 5830 -145 5875 -115
rect 5905 -145 5950 -115
rect 5830 -175 5950 -145
rect 5830 -205 5875 -175
rect 5905 -205 5950 -175
rect 5830 -240 5950 -205
rect 5830 -270 5875 -240
rect 5905 -270 5950 -240
rect 5830 -310 5950 -270
rect 5830 -340 5875 -310
rect 5905 -340 5950 -310
rect 5830 -380 5950 -340
rect 5830 -410 5875 -380
rect 5905 -410 5950 -380
rect 5830 -450 5950 -410
rect 5830 -480 5875 -450
rect 5905 -480 5950 -450
rect 5830 -515 5950 -480
rect 5830 -545 5875 -515
rect 5905 -545 5950 -515
rect 5830 -575 5950 -545
rect 5830 -605 5875 -575
rect 5905 -605 5950 -575
rect 5830 -640 5950 -605
rect 5830 -670 5875 -640
rect 5905 -670 5950 -640
rect 5830 -710 5950 -670
rect 5830 -740 5875 -710
rect 5905 -740 5950 -710
rect 5830 -780 5950 -740
rect 5830 -810 5875 -780
rect 5905 -810 5950 -780
rect 5830 -850 5950 -810
rect 5830 -880 5875 -850
rect 5905 -880 5950 -850
rect 5830 -915 5950 -880
rect 5830 -945 5875 -915
rect 5905 -945 5950 -915
rect 5830 -975 5950 -945
rect 5830 -1005 5875 -975
rect 5905 -1005 5950 -975
rect 5830 -1040 5950 -1005
rect 5830 -1070 5875 -1040
rect 5905 -1070 5950 -1040
rect 5830 -1110 5950 -1070
rect 5830 -1140 5875 -1110
rect 5905 -1140 5950 -1110
rect 5830 -1180 5950 -1140
rect 5830 -1210 5875 -1180
rect 5905 -1210 5950 -1180
rect 5830 -1250 5950 -1210
rect 5830 -1280 5875 -1250
rect 5905 -1280 5950 -1250
rect 5830 -1315 5950 -1280
rect 5830 -1345 5875 -1315
rect 5905 -1345 5950 -1315
rect 5830 -1360 5950 -1345
rect 6180 225 6300 320
rect 6180 195 6225 225
rect 6255 195 6300 225
rect 6180 160 6300 195
rect 6180 130 6225 160
rect 6255 130 6300 160
rect 6180 90 6300 130
rect 6180 60 6225 90
rect 6255 60 6300 90
rect 6180 20 6300 60
rect 6180 -10 6225 20
rect 6255 -10 6300 20
rect 6180 -50 6300 -10
rect 6180 -80 6225 -50
rect 6255 -80 6300 -50
rect 6180 -115 6300 -80
rect 6180 -145 6225 -115
rect 6255 -145 6300 -115
rect 6180 -175 6300 -145
rect 6180 -205 6225 -175
rect 6255 -205 6300 -175
rect 6180 -240 6300 -205
rect 6180 -270 6225 -240
rect 6255 -270 6300 -240
rect 6180 -310 6300 -270
rect 6180 -340 6225 -310
rect 6255 -340 6300 -310
rect 6180 -380 6300 -340
rect 6180 -410 6225 -380
rect 6255 -410 6300 -380
rect 6180 -450 6300 -410
rect 6180 -480 6225 -450
rect 6255 -480 6300 -450
rect 6180 -515 6300 -480
rect 6180 -545 6225 -515
rect 6255 -545 6300 -515
rect 6180 -575 6300 -545
rect 6180 -605 6225 -575
rect 6255 -605 6300 -575
rect 6180 -640 6300 -605
rect 6180 -670 6225 -640
rect 6255 -670 6300 -640
rect 6180 -710 6300 -670
rect 6180 -740 6225 -710
rect 6255 -740 6300 -710
rect 6180 -780 6300 -740
rect 6180 -810 6225 -780
rect 6255 -810 6300 -780
rect 6180 -850 6300 -810
rect 6180 -880 6225 -850
rect 6255 -880 6300 -850
rect 6180 -915 6300 -880
rect 6180 -945 6225 -915
rect 6255 -945 6300 -915
rect 6180 -975 6300 -945
rect 6180 -1005 6225 -975
rect 6255 -1005 6300 -975
rect 6180 -1040 6300 -1005
rect 6180 -1070 6225 -1040
rect 6255 -1070 6300 -1040
rect 6180 -1110 6300 -1070
rect 6180 -1140 6225 -1110
rect 6255 -1140 6300 -1110
rect 6180 -1180 6300 -1140
rect 6180 -1210 6225 -1180
rect 6255 -1210 6300 -1180
rect 6180 -1250 6300 -1210
rect 6180 -1280 6225 -1250
rect 6255 -1280 6300 -1250
rect 6180 -1315 6300 -1280
rect 6180 -1345 6225 -1315
rect 6255 -1345 6300 -1315
rect 6180 -1360 6300 -1345
rect 6530 225 6650 320
rect 6530 195 6575 225
rect 6605 195 6650 225
rect 6530 160 6650 195
rect 6530 130 6575 160
rect 6605 130 6650 160
rect 6530 90 6650 130
rect 6530 60 6575 90
rect 6605 60 6650 90
rect 6530 20 6650 60
rect 6530 -10 6575 20
rect 6605 -10 6650 20
rect 6530 -50 6650 -10
rect 6530 -80 6575 -50
rect 6605 -80 6650 -50
rect 6530 -115 6650 -80
rect 6530 -145 6575 -115
rect 6605 -145 6650 -115
rect 6530 -175 6650 -145
rect 6530 -205 6575 -175
rect 6605 -205 6650 -175
rect 6530 -240 6650 -205
rect 6530 -270 6575 -240
rect 6605 -270 6650 -240
rect 6530 -310 6650 -270
rect 6530 -340 6575 -310
rect 6605 -340 6650 -310
rect 6530 -380 6650 -340
rect 6530 -410 6575 -380
rect 6605 -410 6650 -380
rect 6530 -450 6650 -410
rect 6530 -480 6575 -450
rect 6605 -480 6650 -450
rect 6530 -515 6650 -480
rect 6530 -545 6575 -515
rect 6605 -545 6650 -515
rect 6530 -575 6650 -545
rect 6530 -605 6575 -575
rect 6605 -605 6650 -575
rect 6530 -640 6650 -605
rect 6530 -670 6575 -640
rect 6605 -670 6650 -640
rect 6530 -710 6650 -670
rect 6530 -740 6575 -710
rect 6605 -740 6650 -710
rect 6530 -780 6650 -740
rect 6530 -810 6575 -780
rect 6605 -810 6650 -780
rect 6530 -850 6650 -810
rect 6530 -880 6575 -850
rect 6605 -880 6650 -850
rect 6530 -915 6650 -880
rect 6530 -945 6575 -915
rect 6605 -945 6650 -915
rect 6530 -975 6650 -945
rect 6530 -1005 6575 -975
rect 6605 -1005 6650 -975
rect 6530 -1040 6650 -1005
rect 6530 -1070 6575 -1040
rect 6605 -1070 6650 -1040
rect 6530 -1110 6650 -1070
rect 6530 -1140 6575 -1110
rect 6605 -1140 6650 -1110
rect 6530 -1180 6650 -1140
rect 6530 -1210 6575 -1180
rect 6605 -1210 6650 -1180
rect 6530 -1250 6650 -1210
rect 6530 -1280 6575 -1250
rect 6605 -1280 6650 -1250
rect 6530 -1315 6650 -1280
rect 6530 -1345 6575 -1315
rect 6605 -1345 6650 -1315
rect 6530 -1360 6650 -1345
rect 6880 225 7000 320
rect 6880 195 6925 225
rect 6955 195 7000 225
rect 6880 160 7000 195
rect 6880 130 6925 160
rect 6955 130 7000 160
rect 6880 90 7000 130
rect 6880 60 6925 90
rect 6955 60 7000 90
rect 6880 20 7000 60
rect 6880 -10 6925 20
rect 6955 -10 7000 20
rect 6880 -50 7000 -10
rect 6880 -80 6925 -50
rect 6955 -80 7000 -50
rect 6880 -115 7000 -80
rect 6880 -145 6925 -115
rect 6955 -145 7000 -115
rect 6880 -175 7000 -145
rect 6880 -205 6925 -175
rect 6955 -205 7000 -175
rect 6880 -240 7000 -205
rect 6880 -270 6925 -240
rect 6955 -270 7000 -240
rect 6880 -310 7000 -270
rect 6880 -340 6925 -310
rect 6955 -340 7000 -310
rect 6880 -380 7000 -340
rect 6880 -410 6925 -380
rect 6955 -410 7000 -380
rect 6880 -450 7000 -410
rect 6880 -480 6925 -450
rect 6955 -480 7000 -450
rect 6880 -515 7000 -480
rect 6880 -545 6925 -515
rect 6955 -545 7000 -515
rect 6880 -575 7000 -545
rect 6880 -605 6925 -575
rect 6955 -605 7000 -575
rect 6880 -640 7000 -605
rect 6880 -670 6925 -640
rect 6955 -670 7000 -640
rect 6880 -710 7000 -670
rect 6880 -740 6925 -710
rect 6955 -740 7000 -710
rect 6880 -780 7000 -740
rect 6880 -810 6925 -780
rect 6955 -810 7000 -780
rect 6880 -850 7000 -810
rect 6880 -880 6925 -850
rect 6955 -880 7000 -850
rect 6880 -915 7000 -880
rect 6880 -945 6925 -915
rect 6955 -945 7000 -915
rect 6880 -975 7000 -945
rect 6880 -1005 6925 -975
rect 6955 -1005 7000 -975
rect 6880 -1040 7000 -1005
rect 6880 -1070 6925 -1040
rect 6955 -1070 7000 -1040
rect 6880 -1110 7000 -1070
rect 6880 -1140 6925 -1110
rect 6955 -1140 7000 -1110
rect 6880 -1180 7000 -1140
rect 6880 -1210 6925 -1180
rect 6955 -1210 7000 -1180
rect 6880 -1250 7000 -1210
rect 6880 -1280 6925 -1250
rect 6955 -1280 7000 -1250
rect 6880 -1315 7000 -1280
rect 6880 -1345 6925 -1315
rect 6955 -1345 7000 -1315
rect 6880 -1360 7000 -1345
rect 7230 225 7350 320
rect 7230 195 7275 225
rect 7305 195 7350 225
rect 7230 160 7350 195
rect 7230 130 7275 160
rect 7305 130 7350 160
rect 7230 90 7350 130
rect 7230 60 7275 90
rect 7305 60 7350 90
rect 7230 20 7350 60
rect 7230 -10 7275 20
rect 7305 -10 7350 20
rect 7230 -50 7350 -10
rect 7230 -80 7275 -50
rect 7305 -80 7350 -50
rect 7230 -115 7350 -80
rect 7230 -145 7275 -115
rect 7305 -145 7350 -115
rect 7230 -175 7350 -145
rect 7230 -205 7275 -175
rect 7305 -205 7350 -175
rect 7230 -240 7350 -205
rect 7230 -270 7275 -240
rect 7305 -270 7350 -240
rect 7230 -310 7350 -270
rect 7230 -340 7275 -310
rect 7305 -340 7350 -310
rect 7230 -380 7350 -340
rect 7230 -410 7275 -380
rect 7305 -410 7350 -380
rect 7230 -450 7350 -410
rect 7230 -480 7275 -450
rect 7305 -480 7350 -450
rect 7230 -515 7350 -480
rect 7230 -545 7275 -515
rect 7305 -545 7350 -515
rect 7230 -575 7350 -545
rect 7230 -605 7275 -575
rect 7305 -605 7350 -575
rect 7230 -640 7350 -605
rect 7230 -670 7275 -640
rect 7305 -670 7350 -640
rect 7230 -710 7350 -670
rect 7230 -740 7275 -710
rect 7305 -740 7350 -710
rect 7230 -780 7350 -740
rect 7230 -810 7275 -780
rect 7305 -810 7350 -780
rect 7230 -850 7350 -810
rect 7230 -880 7275 -850
rect 7305 -880 7350 -850
rect 7230 -915 7350 -880
rect 7230 -945 7275 -915
rect 7305 -945 7350 -915
rect 7230 -975 7350 -945
rect 7230 -1005 7275 -975
rect 7305 -1005 7350 -975
rect 7230 -1040 7350 -1005
rect 7230 -1070 7275 -1040
rect 7305 -1070 7350 -1040
rect 7230 -1110 7350 -1070
rect 7230 -1140 7275 -1110
rect 7305 -1140 7350 -1110
rect 7230 -1180 7350 -1140
rect 7230 -1210 7275 -1180
rect 7305 -1210 7350 -1180
rect 7230 -1250 7350 -1210
rect 7230 -1280 7275 -1250
rect 7305 -1280 7350 -1250
rect 7230 -1315 7350 -1280
rect 7230 -1345 7275 -1315
rect 7305 -1345 7350 -1315
rect 7230 -1360 7350 -1345
rect 7580 225 7700 320
rect 7580 195 7625 225
rect 7655 195 7700 225
rect 7580 160 7700 195
rect 7580 130 7625 160
rect 7655 130 7700 160
rect 7580 90 7700 130
rect 7580 60 7625 90
rect 7655 60 7700 90
rect 7580 20 7700 60
rect 7580 -10 7625 20
rect 7655 -10 7700 20
rect 7580 -50 7700 -10
rect 7580 -80 7625 -50
rect 7655 -80 7700 -50
rect 7580 -115 7700 -80
rect 7580 -145 7625 -115
rect 7655 -145 7700 -115
rect 7580 -175 7700 -145
rect 7580 -205 7625 -175
rect 7655 -205 7700 -175
rect 7580 -240 7700 -205
rect 7580 -270 7625 -240
rect 7655 -270 7700 -240
rect 7580 -310 7700 -270
rect 7580 -340 7625 -310
rect 7655 -340 7700 -310
rect 7580 -380 7700 -340
rect 7580 -410 7625 -380
rect 7655 -410 7700 -380
rect 7580 -450 7700 -410
rect 7580 -480 7625 -450
rect 7655 -480 7700 -450
rect 7580 -515 7700 -480
rect 7580 -545 7625 -515
rect 7655 -545 7700 -515
rect 7580 -575 7700 -545
rect 7580 -605 7625 -575
rect 7655 -605 7700 -575
rect 7580 -640 7700 -605
rect 7580 -670 7625 -640
rect 7655 -670 7700 -640
rect 7580 -710 7700 -670
rect 7580 -740 7625 -710
rect 7655 -740 7700 -710
rect 7580 -780 7700 -740
rect 7580 -810 7625 -780
rect 7655 -810 7700 -780
rect 7580 -850 7700 -810
rect 7580 -880 7625 -850
rect 7655 -880 7700 -850
rect 7580 -915 7700 -880
rect 7580 -945 7625 -915
rect 7655 -945 7700 -915
rect 7580 -975 7700 -945
rect 7580 -1005 7625 -975
rect 7655 -1005 7700 -975
rect 7580 -1040 7700 -1005
rect 7580 -1070 7625 -1040
rect 7655 -1070 7700 -1040
rect 7580 -1110 7700 -1070
rect 7580 -1140 7625 -1110
rect 7655 -1140 7700 -1110
rect 7580 -1180 7700 -1140
rect 7580 -1210 7625 -1180
rect 7655 -1210 7700 -1180
rect 7580 -1250 7700 -1210
rect 7580 -1280 7625 -1250
rect 7655 -1280 7700 -1250
rect 7580 -1315 7700 -1280
rect 7580 -1345 7625 -1315
rect 7655 -1345 7700 -1315
rect 7580 -1360 7700 -1345
rect 7930 225 8050 320
rect 7930 195 7975 225
rect 8005 195 8050 225
rect 7930 160 8050 195
rect 7930 130 7975 160
rect 8005 130 8050 160
rect 7930 90 8050 130
rect 7930 60 7975 90
rect 8005 60 8050 90
rect 7930 20 8050 60
rect 7930 -10 7975 20
rect 8005 -10 8050 20
rect 7930 -50 8050 -10
rect 7930 -80 7975 -50
rect 8005 -80 8050 -50
rect 7930 -115 8050 -80
rect 7930 -145 7975 -115
rect 8005 -145 8050 -115
rect 7930 -175 8050 -145
rect 7930 -205 7975 -175
rect 8005 -205 8050 -175
rect 7930 -240 8050 -205
rect 7930 -270 7975 -240
rect 8005 -270 8050 -240
rect 7930 -310 8050 -270
rect 7930 -340 7975 -310
rect 8005 -340 8050 -310
rect 7930 -380 8050 -340
rect 7930 -410 7975 -380
rect 8005 -410 8050 -380
rect 7930 -450 8050 -410
rect 7930 -480 7975 -450
rect 8005 -480 8050 -450
rect 7930 -515 8050 -480
rect 7930 -545 7975 -515
rect 8005 -545 8050 -515
rect 7930 -575 8050 -545
rect 7930 -605 7975 -575
rect 8005 -605 8050 -575
rect 7930 -640 8050 -605
rect 7930 -670 7975 -640
rect 8005 -670 8050 -640
rect 7930 -710 8050 -670
rect 7930 -740 7975 -710
rect 8005 -740 8050 -710
rect 7930 -780 8050 -740
rect 7930 -810 7975 -780
rect 8005 -810 8050 -780
rect 7930 -850 8050 -810
rect 7930 -880 7975 -850
rect 8005 -880 8050 -850
rect 7930 -915 8050 -880
rect 7930 -945 7975 -915
rect 8005 -945 8050 -915
rect 7930 -975 8050 -945
rect 7930 -1005 7975 -975
rect 8005 -1005 8050 -975
rect 7930 -1040 8050 -1005
rect 7930 -1070 7975 -1040
rect 8005 -1070 8050 -1040
rect 7930 -1110 8050 -1070
rect 7930 -1140 7975 -1110
rect 8005 -1140 8050 -1110
rect 7930 -1180 8050 -1140
rect 7930 -1210 7975 -1180
rect 8005 -1210 8050 -1180
rect 7930 -1250 8050 -1210
rect 7930 -1280 7975 -1250
rect 8005 -1280 8050 -1250
rect 7930 -1315 8050 -1280
rect 7930 -1345 7975 -1315
rect 8005 -1345 8050 -1315
rect 7930 -1360 8050 -1345
rect 8280 225 8400 320
rect 8280 195 8325 225
rect 8355 195 8400 225
rect 8280 160 8400 195
rect 8280 130 8325 160
rect 8355 130 8400 160
rect 8280 90 8400 130
rect 8280 60 8325 90
rect 8355 60 8400 90
rect 8280 20 8400 60
rect 8280 -10 8325 20
rect 8355 -10 8400 20
rect 8280 -50 8400 -10
rect 8280 -80 8325 -50
rect 8355 -80 8400 -50
rect 8280 -115 8400 -80
rect 8280 -145 8325 -115
rect 8355 -145 8400 -115
rect 8280 -175 8400 -145
rect 8280 -205 8325 -175
rect 8355 -205 8400 -175
rect 8280 -240 8400 -205
rect 8280 -270 8325 -240
rect 8355 -270 8400 -240
rect 8280 -310 8400 -270
rect 8280 -340 8325 -310
rect 8355 -340 8400 -310
rect 8280 -380 8400 -340
rect 8280 -410 8325 -380
rect 8355 -410 8400 -380
rect 8280 -450 8400 -410
rect 8280 -480 8325 -450
rect 8355 -480 8400 -450
rect 8280 -515 8400 -480
rect 8280 -545 8325 -515
rect 8355 -545 8400 -515
rect 8280 -575 8400 -545
rect 8280 -605 8325 -575
rect 8355 -605 8400 -575
rect 8280 -640 8400 -605
rect 8280 -670 8325 -640
rect 8355 -670 8400 -640
rect 8280 -710 8400 -670
rect 8280 -740 8325 -710
rect 8355 -740 8400 -710
rect 8280 -780 8400 -740
rect 8280 -810 8325 -780
rect 8355 -810 8400 -780
rect 8280 -850 8400 -810
rect 8280 -880 8325 -850
rect 8355 -880 8400 -850
rect 8280 -915 8400 -880
rect 8280 -945 8325 -915
rect 8355 -945 8400 -915
rect 8280 -975 8400 -945
rect 8280 -1005 8325 -975
rect 8355 -1005 8400 -975
rect 8280 -1040 8400 -1005
rect 8280 -1070 8325 -1040
rect 8355 -1070 8400 -1040
rect 8280 -1110 8400 -1070
rect 8280 -1140 8325 -1110
rect 8355 -1140 8400 -1110
rect 8280 -1180 8400 -1140
rect 8280 -1210 8325 -1180
rect 8355 -1210 8400 -1180
rect 8280 -1250 8400 -1210
rect 8280 -1280 8325 -1250
rect 8355 -1280 8400 -1250
rect 8280 -1315 8400 -1280
rect 8280 -1345 8325 -1315
rect 8355 -1345 8400 -1315
rect 8280 -1360 8400 -1345
rect 8630 225 8750 320
rect 8630 195 8675 225
rect 8705 195 8750 225
rect 8630 160 8750 195
rect 8630 130 8675 160
rect 8705 130 8750 160
rect 8630 90 8750 130
rect 8630 60 8675 90
rect 8705 60 8750 90
rect 8630 20 8750 60
rect 8630 -10 8675 20
rect 8705 -10 8750 20
rect 8630 -50 8750 -10
rect 8630 -80 8675 -50
rect 8705 -80 8750 -50
rect 8630 -115 8750 -80
rect 8630 -145 8675 -115
rect 8705 -145 8750 -115
rect 8630 -175 8750 -145
rect 8630 -205 8675 -175
rect 8705 -205 8750 -175
rect 8630 -240 8750 -205
rect 8630 -270 8675 -240
rect 8705 -270 8750 -240
rect 8630 -310 8750 -270
rect 8630 -340 8675 -310
rect 8705 -340 8750 -310
rect 8630 -380 8750 -340
rect 8630 -410 8675 -380
rect 8705 -410 8750 -380
rect 8630 -450 8750 -410
rect 8630 -480 8675 -450
rect 8705 -480 8750 -450
rect 8630 -515 8750 -480
rect 8630 -545 8675 -515
rect 8705 -545 8750 -515
rect 8630 -575 8750 -545
rect 8630 -605 8675 -575
rect 8705 -605 8750 -575
rect 8630 -640 8750 -605
rect 8630 -670 8675 -640
rect 8705 -670 8750 -640
rect 8630 -710 8750 -670
rect 8630 -740 8675 -710
rect 8705 -740 8750 -710
rect 8630 -780 8750 -740
rect 8630 -810 8675 -780
rect 8705 -810 8750 -780
rect 8630 -850 8750 -810
rect 8630 -880 8675 -850
rect 8705 -880 8750 -850
rect 8630 -915 8750 -880
rect 8630 -945 8675 -915
rect 8705 -945 8750 -915
rect 8630 -975 8750 -945
rect 8630 -1005 8675 -975
rect 8705 -1005 8750 -975
rect 8630 -1040 8750 -1005
rect 8630 -1070 8675 -1040
rect 8705 -1070 8750 -1040
rect 8630 -1110 8750 -1070
rect 8630 -1140 8675 -1110
rect 8705 -1140 8750 -1110
rect 8630 -1180 8750 -1140
rect 8630 -1210 8675 -1180
rect 8705 -1210 8750 -1180
rect 8630 -1250 8750 -1210
rect 8630 -1280 8675 -1250
rect 8705 -1280 8750 -1250
rect 8630 -1315 8750 -1280
rect 8630 -1345 8675 -1315
rect 8705 -1345 8750 -1315
rect 8630 -1360 8750 -1345
rect 8980 225 9100 320
rect 8980 195 9025 225
rect 9055 195 9100 225
rect 8980 160 9100 195
rect 8980 130 9025 160
rect 9055 130 9100 160
rect 8980 90 9100 130
rect 8980 60 9025 90
rect 9055 60 9100 90
rect 8980 20 9100 60
rect 8980 -10 9025 20
rect 9055 -10 9100 20
rect 8980 -50 9100 -10
rect 8980 -80 9025 -50
rect 9055 -80 9100 -50
rect 8980 -115 9100 -80
rect 8980 -145 9025 -115
rect 9055 -145 9100 -115
rect 8980 -175 9100 -145
rect 8980 -205 9025 -175
rect 9055 -205 9100 -175
rect 8980 -240 9100 -205
rect 8980 -270 9025 -240
rect 9055 -270 9100 -240
rect 8980 -310 9100 -270
rect 8980 -340 9025 -310
rect 9055 -340 9100 -310
rect 8980 -380 9100 -340
rect 8980 -410 9025 -380
rect 9055 -410 9100 -380
rect 8980 -450 9100 -410
rect 8980 -480 9025 -450
rect 9055 -480 9100 -450
rect 8980 -515 9100 -480
rect 8980 -545 9025 -515
rect 9055 -545 9100 -515
rect 8980 -575 9100 -545
rect 8980 -605 9025 -575
rect 9055 -605 9100 -575
rect 8980 -640 9100 -605
rect 8980 -670 9025 -640
rect 9055 -670 9100 -640
rect 8980 -710 9100 -670
rect 8980 -740 9025 -710
rect 9055 -740 9100 -710
rect 8980 -780 9100 -740
rect 8980 -810 9025 -780
rect 9055 -810 9100 -780
rect 8980 -850 9100 -810
rect 8980 -880 9025 -850
rect 9055 -880 9100 -850
rect 8980 -915 9100 -880
rect 8980 -945 9025 -915
rect 9055 -945 9100 -915
rect 8980 -975 9100 -945
rect 8980 -1005 9025 -975
rect 9055 -1005 9100 -975
rect 8980 -1040 9100 -1005
rect 8980 -1070 9025 -1040
rect 9055 -1070 9100 -1040
rect 8980 -1110 9100 -1070
rect 8980 -1140 9025 -1110
rect 9055 -1140 9100 -1110
rect 8980 -1180 9100 -1140
rect 8980 -1210 9025 -1180
rect 9055 -1210 9100 -1180
rect 8980 -1250 9100 -1210
rect 8980 -1280 9025 -1250
rect 9055 -1280 9100 -1250
rect 8980 -1315 9100 -1280
rect 8980 -1345 9025 -1315
rect 9055 -1345 9100 -1315
rect 8980 -1360 9100 -1345
<< via1 >>
rect 2115 19280 2145 19310
rect 2115 19215 2145 19245
rect 2115 19145 2145 19175
rect 2115 19075 2145 19105
rect 2115 19005 2145 19035
rect 2115 18940 2145 18970
rect 2115 18880 2145 18910
rect 2115 18815 2145 18845
rect 2115 18745 2145 18775
rect 2115 18675 2145 18705
rect 2115 18605 2145 18635
rect 2115 18540 2145 18570
rect 2115 18480 2145 18510
rect 2115 18415 2145 18445
rect 2115 18345 2145 18375
rect 2115 18275 2145 18305
rect 2115 18205 2145 18235
rect 2115 18140 2145 18170
rect 2115 18080 2145 18110
rect 2115 18015 2145 18045
rect 2115 17945 2145 17975
rect 2115 17875 2145 17905
rect 2115 17805 2145 17835
rect 2115 17740 2145 17770
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 2075 15660 2105 15690
rect 2115 15660 2145 15690
rect 2155 15660 2185 15690
rect 2075 15620 2105 15650
rect 2115 15620 2145 15650
rect 2155 15620 2185 15650
rect 2075 15580 2105 15610
rect 2115 15580 2145 15610
rect 2155 15580 2185 15610
rect 2075 12680 2105 12710
rect 2115 12680 2145 12710
rect 2155 12680 2185 12710
rect 2075 12640 2105 12670
rect 2115 12640 2145 12670
rect 2155 12640 2185 12670
rect 2075 12520 2105 12550
rect 2115 12520 2145 12550
rect 2155 12520 2185 12550
rect 2075 12480 2105 12510
rect 2115 12480 2145 12510
rect 2155 12480 2185 12510
rect 2075 12440 2105 12470
rect 2115 12440 2145 12470
rect 2155 12440 2185 12470
rect 2210 15895 2240 15925
rect 2250 15895 2280 15925
rect 2290 15895 2320 15925
rect 1325 9605 1355 9635
rect 1325 9540 1355 9570
rect 1325 9470 1355 9500
rect 1325 9400 1355 9430
rect 1325 9330 1355 9360
rect 1325 9265 1355 9295
rect 1325 9205 1355 9235
rect 1325 9140 1355 9170
rect 1325 9070 1355 9100
rect 1325 9000 1355 9030
rect 1325 8930 1355 8960
rect 1325 8865 1355 8895
rect 1325 8805 1355 8835
rect 1325 8740 1355 8770
rect 1325 8670 1355 8700
rect 1325 8600 1355 8630
rect 1325 8530 1355 8560
rect 1325 8465 1355 8495
rect 1325 8405 1355 8435
rect 1325 8340 1355 8370
rect 1325 8270 1355 8300
rect 1325 8200 1355 8230
rect 1325 8130 1355 8160
rect 6665 15565 6695 15595
rect 6705 15565 6735 15595
rect 6745 15565 6775 15595
rect 6665 15525 6695 15555
rect 6705 15525 6735 15555
rect 6745 15525 6775 15555
rect 6665 15485 6695 15515
rect 6705 15485 6735 15515
rect 6745 15485 6775 15515
rect 2250 9605 2280 9635
rect 2250 9540 2280 9570
rect 2250 9470 2280 9500
rect 2250 9400 2280 9430
rect 2250 9330 2280 9360
rect 2250 9265 2280 9295
rect 2250 9205 2280 9235
rect 2250 9140 2280 9170
rect 2250 9070 2280 9100
rect 2250 9000 2280 9030
rect 2250 8930 2280 8960
rect 2250 8865 2280 8895
rect 2250 8805 2280 8835
rect 2250 8740 2280 8770
rect 2250 8670 2280 8700
rect 2250 8600 2280 8630
rect 2250 8530 2280 8560
rect 2250 8465 2280 8495
rect 2250 8405 2280 8435
rect 2250 8340 2280 8370
rect 2250 8270 2280 8300
rect 2250 8200 2280 8230
rect 2250 8130 2280 8160
rect 1985 8040 2015 8070
rect 2025 8040 2055 8070
rect 2065 8040 2095 8070
rect 1635 7985 1665 8015
rect 1675 7985 1705 8015
rect 1715 7985 1745 8015
rect 2480 8040 2510 8070
rect 3180 9605 3210 9635
rect 3180 9540 3210 9570
rect 3180 9470 3210 9500
rect 3180 9400 3210 9430
rect 3180 9330 3210 9360
rect 3180 9265 3210 9295
rect 3180 9205 3210 9235
rect 3180 9140 3210 9170
rect 3180 9070 3210 9100
rect 3180 9000 3210 9030
rect 3180 8930 3210 8960
rect 3180 8865 3210 8895
rect 3180 8805 3210 8835
rect 3180 8740 3210 8770
rect 3180 8670 3210 8700
rect 3180 8600 3210 8630
rect 3180 8530 3210 8560
rect 3180 8465 3210 8495
rect 3180 8405 3210 8435
rect 3180 8340 3210 8370
rect 3180 8270 3210 8300
rect 3180 8200 3210 8230
rect 3180 8130 3210 8160
rect 2850 7930 2880 7960
rect 3635 7985 3665 8015
rect 3855 7985 3885 8015
rect 3385 7930 3415 7960
rect 2720 7820 2750 7850
rect 3080 7820 3110 7850
rect 3295 7840 3325 7870
rect 935 7705 965 7735
rect 975 7705 1005 7735
rect 1015 7705 1045 7735
rect 935 7665 965 7695
rect 975 7665 1005 7695
rect 1015 7665 1045 7695
rect 935 7625 965 7655
rect 975 7625 1005 7655
rect 1015 7625 1045 7655
rect 3295 7800 3325 7830
rect 3295 7760 3325 7790
rect 3080 6590 3110 6620
rect 3440 7840 3470 7870
rect 3440 7800 3470 7830
rect 3440 7760 3470 7790
rect 3385 5305 3415 5335
rect 4310 7705 4340 7735
rect 4310 7665 4340 7695
rect 4310 7625 4340 7655
rect 4420 7705 4450 7735
rect 4420 7665 4450 7695
rect 4420 7625 4450 7655
rect 4530 7705 4560 7735
rect 4530 7665 4560 7695
rect 4530 7625 4560 7655
rect 5095 7985 5125 8015
rect 5315 7985 5345 8015
rect 5475 7930 5505 7960
rect 6150 7930 6180 7960
rect 4640 7705 4670 7735
rect 4640 7665 4670 7695
rect 4640 7625 4670 7655
rect 5550 7840 5580 7870
rect 5550 7800 5580 7830
rect 5550 7760 5580 7790
rect 5475 5365 5505 5395
rect 3440 4625 3470 4655
rect 4475 4625 4505 4655
rect 5875 6935 5905 6965
rect 5625 6535 5655 6565
rect 6665 12895 6695 12925
rect 6705 12895 6735 12925
rect 6745 12895 6775 12925
rect 6665 12855 6695 12885
rect 6705 12855 6735 12885
rect 6745 12855 6775 12885
rect 6665 12815 6695 12845
rect 6705 12815 6735 12845
rect 6745 12815 6775 12845
rect 6665 12120 6695 12150
rect 6705 12120 6735 12150
rect 6745 12120 6775 12150
rect 6665 12080 6695 12110
rect 6705 12080 6735 12110
rect 6745 12080 6775 12110
rect 6665 12040 6695 12070
rect 6705 12040 6735 12070
rect 6745 12040 6775 12070
rect 6665 11135 6695 11165
rect 6705 11135 6735 11165
rect 6745 11135 6775 11165
rect 6665 11095 6695 11125
rect 6705 11095 6735 11125
rect 6745 11095 6775 11125
rect 6665 11055 6695 11085
rect 6705 11055 6735 11085
rect 6745 11055 6775 11085
rect 6665 10410 6695 10440
rect 6705 10410 6735 10440
rect 6745 10410 6775 10440
rect 6665 10370 6695 10400
rect 6705 10370 6735 10400
rect 6745 10370 6775 10400
rect 6665 10330 6695 10360
rect 6705 10330 6735 10360
rect 6745 10330 6775 10360
rect 6665 10050 6695 10080
rect 6705 10050 6735 10080
rect 6745 10050 6775 10080
rect 6665 10010 6695 10040
rect 6705 10010 6735 10040
rect 6745 10010 6775 10040
rect 6665 9970 6695 10000
rect 6705 9970 6735 10000
rect 6745 9970 6775 10000
rect 6705 9540 6735 9570
rect 6705 9470 6735 9500
rect 6705 9400 6735 9430
rect 6705 9330 6735 9360
rect 6705 9265 6735 9295
rect 6705 9205 6735 9235
rect 6705 9140 6735 9170
rect 6705 9070 6735 9100
rect 6705 9000 6735 9030
rect 6705 8930 6735 8960
rect 6705 8865 6735 8895
rect 6705 8805 6735 8835
rect 6705 8740 6735 8770
rect 6705 8670 6735 8700
rect 6705 8600 6735 8630
rect 6705 8530 6735 8560
rect 6705 8465 6735 8495
rect 6705 8405 6735 8435
rect 6705 8340 6735 8370
rect 6705 8270 6735 8300
rect 6705 8200 6735 8230
rect 6705 8130 6735 8160
rect 7625 9605 7655 9635
rect 7625 9540 7655 9570
rect 7625 9470 7655 9500
rect 7625 9400 7655 9430
rect 7625 9330 7655 9360
rect 7625 9265 7655 9295
rect 7625 9205 7655 9235
rect 7625 9140 7655 9170
rect 7625 9070 7655 9100
rect 7625 9000 7655 9030
rect 7625 8930 7655 8960
rect 7625 8865 7655 8895
rect 7625 8805 7655 8835
rect 7625 8740 7655 8770
rect 7625 8670 7655 8700
rect 7625 8600 7655 8630
rect 7625 8530 7655 8560
rect 7625 8465 7655 8495
rect 7625 8405 7655 8435
rect 7625 8340 7655 8370
rect 7625 8270 7655 8300
rect 7625 8200 7655 8230
rect 7625 8130 7655 8160
rect 6470 8040 6500 8070
rect 6885 8040 6915 8070
rect 6925 8040 6955 8070
rect 6965 8040 6995 8070
rect 7235 7985 7265 8015
rect 7275 7985 7305 8015
rect 7315 7985 7345 8015
rect 6225 6935 6255 6965
rect 7935 7705 7965 7735
rect 7975 7705 8005 7735
rect 8015 7705 8045 7735
rect 7935 7665 7965 7695
rect 7975 7665 8005 7695
rect 8015 7665 8045 7695
rect 7935 7625 7965 7655
rect 7975 7625 8005 7655
rect 8015 7625 8045 7655
rect 5875 6535 5905 6565
rect 5625 5940 5655 5970
rect 5550 4625 5580 4655
rect 4475 4405 4505 4435
rect 935 2660 965 2690
rect 975 2660 1005 2690
rect 1015 2660 1045 2690
rect 935 2620 965 2650
rect 975 2620 1005 2650
rect 1015 2620 1045 2650
rect 935 2580 965 2610
rect 975 2580 1005 2610
rect 1015 2580 1045 2610
rect 4420 2660 4450 2690
rect 4420 2620 4450 2650
rect 4420 2580 4450 2610
rect 4530 2660 4560 2690
rect 4530 2620 4560 2650
rect 4530 2580 4560 2610
rect 7935 2660 7965 2690
rect 7975 2660 8005 2690
rect 8015 2660 8045 2690
rect 7935 2620 7965 2650
rect 7975 2620 8005 2650
rect 8015 2620 8045 2650
rect 7935 2580 7965 2610
rect 7975 2580 8005 2610
rect 8015 2580 8045 2610
rect -75 195 -45 225
rect -75 130 -45 160
rect -75 60 -45 90
rect -75 -10 -45 20
rect -75 -80 -45 -50
rect -75 -145 -45 -115
rect -75 -205 -45 -175
rect -75 -270 -45 -240
rect -75 -340 -45 -310
rect -75 -410 -45 -380
rect -75 -480 -45 -450
rect -75 -545 -45 -515
rect -75 -605 -45 -575
rect -75 -670 -45 -640
rect -75 -740 -45 -710
rect -75 -810 -45 -780
rect -75 -880 -45 -850
rect -75 -945 -45 -915
rect -75 -1005 -45 -975
rect -75 -1070 -45 -1040
rect -75 -1140 -45 -1110
rect -75 -1210 -45 -1180
rect -75 -1280 -45 -1250
rect -75 -1345 -45 -1315
rect 275 195 305 225
rect 275 130 305 160
rect 275 60 305 90
rect 275 -10 305 20
rect 275 -80 305 -50
rect 275 -145 305 -115
rect 275 -205 305 -175
rect 275 -270 305 -240
rect 275 -340 305 -310
rect 275 -410 305 -380
rect 275 -480 305 -450
rect 275 -545 305 -515
rect 275 -605 305 -575
rect 275 -670 305 -640
rect 275 -740 305 -710
rect 275 -810 305 -780
rect 275 -880 305 -850
rect 275 -945 305 -915
rect 275 -1005 305 -975
rect 275 -1070 305 -1040
rect 275 -1140 305 -1110
rect 275 -1210 305 -1180
rect 275 -1280 305 -1250
rect 275 -1345 305 -1315
rect 625 195 655 225
rect 625 130 655 160
rect 625 60 655 90
rect 625 -10 655 20
rect 625 -80 655 -50
rect 625 -145 655 -115
rect 625 -205 655 -175
rect 625 -270 655 -240
rect 625 -340 655 -310
rect 625 -410 655 -380
rect 625 -480 655 -450
rect 625 -545 655 -515
rect 625 -605 655 -575
rect 625 -670 655 -640
rect 625 -740 655 -710
rect 625 -810 655 -780
rect 625 -880 655 -850
rect 625 -945 655 -915
rect 625 -1005 655 -975
rect 625 -1070 655 -1040
rect 625 -1140 655 -1110
rect 625 -1210 655 -1180
rect 625 -1280 655 -1250
rect 625 -1345 655 -1315
rect 975 195 1005 225
rect 975 130 1005 160
rect 975 60 1005 90
rect 975 -10 1005 20
rect 975 -80 1005 -50
rect 975 -145 1005 -115
rect 975 -205 1005 -175
rect 975 -270 1005 -240
rect 975 -340 1005 -310
rect 975 -410 1005 -380
rect 975 -480 1005 -450
rect 975 -545 1005 -515
rect 975 -605 1005 -575
rect 975 -670 1005 -640
rect 975 -740 1005 -710
rect 975 -810 1005 -780
rect 975 -880 1005 -850
rect 975 -945 1005 -915
rect 975 -1005 1005 -975
rect 975 -1070 1005 -1040
rect 975 -1140 1005 -1110
rect 975 -1210 1005 -1180
rect 975 -1280 1005 -1250
rect 975 -1345 1005 -1315
rect 1325 195 1355 225
rect 1325 130 1355 160
rect 1325 60 1355 90
rect 1325 -10 1355 20
rect 1325 -80 1355 -50
rect 1325 -145 1355 -115
rect 1325 -205 1355 -175
rect 1325 -270 1355 -240
rect 1325 -340 1355 -310
rect 1325 -410 1355 -380
rect 1325 -480 1355 -450
rect 1325 -545 1355 -515
rect 1325 -605 1355 -575
rect 1325 -670 1355 -640
rect 1325 -740 1355 -710
rect 1325 -810 1355 -780
rect 1325 -880 1355 -850
rect 1325 -945 1355 -915
rect 1325 -1005 1355 -975
rect 1325 -1070 1355 -1040
rect 1325 -1140 1355 -1110
rect 1325 -1210 1355 -1180
rect 1325 -1280 1355 -1250
rect 1325 -1345 1355 -1315
rect 1675 195 1705 225
rect 1675 130 1705 160
rect 1675 60 1705 90
rect 1675 -10 1705 20
rect 1675 -80 1705 -50
rect 1675 -145 1705 -115
rect 1675 -205 1705 -175
rect 1675 -270 1705 -240
rect 1675 -340 1705 -310
rect 1675 -410 1705 -380
rect 1675 -480 1705 -450
rect 1675 -545 1705 -515
rect 1675 -605 1705 -575
rect 1675 -670 1705 -640
rect 1675 -740 1705 -710
rect 1675 -810 1705 -780
rect 1675 -880 1705 -850
rect 1675 -945 1705 -915
rect 1675 -1005 1705 -975
rect 1675 -1070 1705 -1040
rect 1675 -1140 1705 -1110
rect 1675 -1210 1705 -1180
rect 1675 -1280 1705 -1250
rect 1675 -1345 1705 -1315
rect 2025 195 2055 225
rect 2025 130 2055 160
rect 2025 60 2055 90
rect 2025 -10 2055 20
rect 2025 -80 2055 -50
rect 2025 -145 2055 -115
rect 2025 -205 2055 -175
rect 2025 -270 2055 -240
rect 2025 -340 2055 -310
rect 2025 -410 2055 -380
rect 2025 -480 2055 -450
rect 2025 -545 2055 -515
rect 2025 -605 2055 -575
rect 2025 -670 2055 -640
rect 2025 -740 2055 -710
rect 2025 -810 2055 -780
rect 2025 -880 2055 -850
rect 2025 -945 2055 -915
rect 2025 -1005 2055 -975
rect 2025 -1070 2055 -1040
rect 2025 -1140 2055 -1110
rect 2025 -1210 2055 -1180
rect 2025 -1280 2055 -1250
rect 2025 -1345 2055 -1315
rect 2375 195 2405 225
rect 2375 130 2405 160
rect 2375 60 2405 90
rect 2375 -10 2405 20
rect 2375 -80 2405 -50
rect 2375 -145 2405 -115
rect 2375 -205 2405 -175
rect 2375 -270 2405 -240
rect 2375 -340 2405 -310
rect 2375 -410 2405 -380
rect 2375 -480 2405 -450
rect 2375 -545 2405 -515
rect 2375 -605 2405 -575
rect 2375 -670 2405 -640
rect 2375 -740 2405 -710
rect 2375 -810 2405 -780
rect 2375 -880 2405 -850
rect 2375 -945 2405 -915
rect 2375 -1005 2405 -975
rect 2375 -1070 2405 -1040
rect 2375 -1140 2405 -1110
rect 2375 -1210 2405 -1180
rect 2375 -1280 2405 -1250
rect 2375 -1345 2405 -1315
rect 2725 195 2755 225
rect 2725 130 2755 160
rect 2725 60 2755 90
rect 2725 -10 2755 20
rect 2725 -80 2755 -50
rect 2725 -145 2755 -115
rect 2725 -205 2755 -175
rect 2725 -270 2755 -240
rect 2725 -340 2755 -310
rect 2725 -410 2755 -380
rect 2725 -480 2755 -450
rect 2725 -545 2755 -515
rect 2725 -605 2755 -575
rect 2725 -670 2755 -640
rect 2725 -740 2755 -710
rect 2725 -810 2755 -780
rect 2725 -880 2755 -850
rect 2725 -945 2755 -915
rect 2725 -1005 2755 -975
rect 2725 -1070 2755 -1040
rect 2725 -1140 2755 -1110
rect 2725 -1210 2755 -1180
rect 2725 -1280 2755 -1250
rect 2725 -1345 2755 -1315
rect 3075 195 3105 225
rect 3075 130 3105 160
rect 3075 60 3105 90
rect 3075 -10 3105 20
rect 3075 -80 3105 -50
rect 3075 -145 3105 -115
rect 3075 -205 3105 -175
rect 3075 -270 3105 -240
rect 3075 -340 3105 -310
rect 3075 -410 3105 -380
rect 3075 -480 3105 -450
rect 3075 -545 3105 -515
rect 3075 -605 3105 -575
rect 3075 -670 3105 -640
rect 3075 -740 3105 -710
rect 3075 -810 3105 -780
rect 3075 -880 3105 -850
rect 3075 -945 3105 -915
rect 3075 -1005 3105 -975
rect 3075 -1070 3105 -1040
rect 3075 -1140 3105 -1110
rect 3075 -1210 3105 -1180
rect 3075 -1280 3105 -1250
rect 3075 -1345 3105 -1315
rect 3425 195 3455 225
rect 3425 130 3455 160
rect 3425 60 3455 90
rect 3425 -10 3455 20
rect 3425 -80 3455 -50
rect 3425 -145 3455 -115
rect 3425 -205 3455 -175
rect 3425 -270 3455 -240
rect 3425 -340 3455 -310
rect 3425 -410 3455 -380
rect 3425 -480 3455 -450
rect 3425 -545 3455 -515
rect 3425 -605 3455 -575
rect 3425 -670 3455 -640
rect 3425 -740 3455 -710
rect 3425 -810 3455 -780
rect 3425 -880 3455 -850
rect 3425 -945 3455 -915
rect 3425 -1005 3455 -975
rect 3425 -1070 3455 -1040
rect 3425 -1140 3455 -1110
rect 3425 -1210 3455 -1180
rect 3425 -1280 3455 -1250
rect 3425 -1345 3455 -1315
rect 3775 195 3805 225
rect 3775 130 3805 160
rect 3775 60 3805 90
rect 3775 -10 3805 20
rect 3775 -80 3805 -50
rect 3775 -145 3805 -115
rect 3775 -205 3805 -175
rect 3775 -270 3805 -240
rect 3775 -340 3805 -310
rect 3775 -410 3805 -380
rect 3775 -480 3805 -450
rect 3775 -545 3805 -515
rect 3775 -605 3805 -575
rect 3775 -670 3805 -640
rect 3775 -740 3805 -710
rect 3775 -810 3805 -780
rect 3775 -880 3805 -850
rect 3775 -945 3805 -915
rect 3775 -1005 3805 -975
rect 3775 -1070 3805 -1040
rect 3775 -1140 3805 -1110
rect 3775 -1210 3805 -1180
rect 3775 -1280 3805 -1250
rect 3775 -1345 3805 -1315
rect 4125 195 4155 225
rect 4125 130 4155 160
rect 4125 60 4155 90
rect 4125 -10 4155 20
rect 4125 -80 4155 -50
rect 4125 -145 4155 -115
rect 4125 -205 4155 -175
rect 4125 -270 4155 -240
rect 4125 -340 4155 -310
rect 4125 -410 4155 -380
rect 4125 -480 4155 -450
rect 4125 -545 4155 -515
rect 4125 -605 4155 -575
rect 4125 -670 4155 -640
rect 4125 -740 4155 -710
rect 4125 -810 4155 -780
rect 4125 -880 4155 -850
rect 4125 -945 4155 -915
rect 4125 -1005 4155 -975
rect 4125 -1070 4155 -1040
rect 4125 -1140 4155 -1110
rect 4125 -1210 4155 -1180
rect 4125 -1280 4155 -1250
rect 4125 -1345 4155 -1315
rect 4475 195 4505 225
rect 4475 130 4505 160
rect 4475 60 4505 90
rect 4475 -10 4505 20
rect 4475 -80 4505 -50
rect 4475 -145 4505 -115
rect 4475 -205 4505 -175
rect 4475 -270 4505 -240
rect 4475 -340 4505 -310
rect 4475 -410 4505 -380
rect 4475 -480 4505 -450
rect 4475 -545 4505 -515
rect 4475 -605 4505 -575
rect 4475 -670 4505 -640
rect 4475 -740 4505 -710
rect 4475 -810 4505 -780
rect 4475 -880 4505 -850
rect 4475 -945 4505 -915
rect 4475 -1005 4505 -975
rect 4475 -1070 4505 -1040
rect 4475 -1140 4505 -1110
rect 4475 -1210 4505 -1180
rect 4475 -1280 4505 -1250
rect 4475 -1345 4505 -1315
rect 4825 195 4855 225
rect 4825 130 4855 160
rect 4825 60 4855 90
rect 4825 -10 4855 20
rect 4825 -80 4855 -50
rect 4825 -145 4855 -115
rect 4825 -205 4855 -175
rect 4825 -270 4855 -240
rect 4825 -340 4855 -310
rect 4825 -410 4855 -380
rect 4825 -480 4855 -450
rect 4825 -545 4855 -515
rect 4825 -605 4855 -575
rect 4825 -670 4855 -640
rect 4825 -740 4855 -710
rect 4825 -810 4855 -780
rect 4825 -880 4855 -850
rect 4825 -945 4855 -915
rect 4825 -1005 4855 -975
rect 4825 -1070 4855 -1040
rect 4825 -1140 4855 -1110
rect 4825 -1210 4855 -1180
rect 4825 -1280 4855 -1250
rect 4825 -1345 4855 -1315
rect 5175 195 5205 225
rect 5175 130 5205 160
rect 5175 60 5205 90
rect 5175 -10 5205 20
rect 5175 -80 5205 -50
rect 5175 -145 5205 -115
rect 5175 -205 5205 -175
rect 5175 -270 5205 -240
rect 5175 -340 5205 -310
rect 5175 -410 5205 -380
rect 5175 -480 5205 -450
rect 5175 -545 5205 -515
rect 5175 -605 5205 -575
rect 5175 -670 5205 -640
rect 5175 -740 5205 -710
rect 5175 -810 5205 -780
rect 5175 -880 5205 -850
rect 5175 -945 5205 -915
rect 5175 -1005 5205 -975
rect 5175 -1070 5205 -1040
rect 5175 -1140 5205 -1110
rect 5175 -1210 5205 -1180
rect 5175 -1280 5205 -1250
rect 5175 -1345 5205 -1315
rect 5525 195 5555 225
rect 5525 130 5555 160
rect 5525 60 5555 90
rect 5525 -10 5555 20
rect 5525 -80 5555 -50
rect 5525 -145 5555 -115
rect 5525 -205 5555 -175
rect 5525 -270 5555 -240
rect 5525 -340 5555 -310
rect 5525 -410 5555 -380
rect 5525 -480 5555 -450
rect 5525 -545 5555 -515
rect 5525 -605 5555 -575
rect 5525 -670 5555 -640
rect 5525 -740 5555 -710
rect 5525 -810 5555 -780
rect 5525 -880 5555 -850
rect 5525 -945 5555 -915
rect 5525 -1005 5555 -975
rect 5525 -1070 5555 -1040
rect 5525 -1140 5555 -1110
rect 5525 -1210 5555 -1180
rect 5525 -1280 5555 -1250
rect 5525 -1345 5555 -1315
rect 5875 195 5905 225
rect 5875 130 5905 160
rect 5875 60 5905 90
rect 5875 -10 5905 20
rect 5875 -80 5905 -50
rect 5875 -145 5905 -115
rect 5875 -205 5905 -175
rect 5875 -270 5905 -240
rect 5875 -340 5905 -310
rect 5875 -410 5905 -380
rect 5875 -480 5905 -450
rect 5875 -545 5905 -515
rect 5875 -605 5905 -575
rect 5875 -670 5905 -640
rect 5875 -740 5905 -710
rect 5875 -810 5905 -780
rect 5875 -880 5905 -850
rect 5875 -945 5905 -915
rect 5875 -1005 5905 -975
rect 5875 -1070 5905 -1040
rect 5875 -1140 5905 -1110
rect 5875 -1210 5905 -1180
rect 5875 -1280 5905 -1250
rect 5875 -1345 5905 -1315
rect 6225 195 6255 225
rect 6225 130 6255 160
rect 6225 60 6255 90
rect 6225 -10 6255 20
rect 6225 -80 6255 -50
rect 6225 -145 6255 -115
rect 6225 -205 6255 -175
rect 6225 -270 6255 -240
rect 6225 -340 6255 -310
rect 6225 -410 6255 -380
rect 6225 -480 6255 -450
rect 6225 -545 6255 -515
rect 6225 -605 6255 -575
rect 6225 -670 6255 -640
rect 6225 -740 6255 -710
rect 6225 -810 6255 -780
rect 6225 -880 6255 -850
rect 6225 -945 6255 -915
rect 6225 -1005 6255 -975
rect 6225 -1070 6255 -1040
rect 6225 -1140 6255 -1110
rect 6225 -1210 6255 -1180
rect 6225 -1280 6255 -1250
rect 6225 -1345 6255 -1315
rect 6575 195 6605 225
rect 6575 130 6605 160
rect 6575 60 6605 90
rect 6575 -10 6605 20
rect 6575 -80 6605 -50
rect 6575 -145 6605 -115
rect 6575 -205 6605 -175
rect 6575 -270 6605 -240
rect 6575 -340 6605 -310
rect 6575 -410 6605 -380
rect 6575 -480 6605 -450
rect 6575 -545 6605 -515
rect 6575 -605 6605 -575
rect 6575 -670 6605 -640
rect 6575 -740 6605 -710
rect 6575 -810 6605 -780
rect 6575 -880 6605 -850
rect 6575 -945 6605 -915
rect 6575 -1005 6605 -975
rect 6575 -1070 6605 -1040
rect 6575 -1140 6605 -1110
rect 6575 -1210 6605 -1180
rect 6575 -1280 6605 -1250
rect 6575 -1345 6605 -1315
rect 6925 195 6955 225
rect 6925 130 6955 160
rect 6925 60 6955 90
rect 6925 -10 6955 20
rect 6925 -80 6955 -50
rect 6925 -145 6955 -115
rect 6925 -205 6955 -175
rect 6925 -270 6955 -240
rect 6925 -340 6955 -310
rect 6925 -410 6955 -380
rect 6925 -480 6955 -450
rect 6925 -545 6955 -515
rect 6925 -605 6955 -575
rect 6925 -670 6955 -640
rect 6925 -740 6955 -710
rect 6925 -810 6955 -780
rect 6925 -880 6955 -850
rect 6925 -945 6955 -915
rect 6925 -1005 6955 -975
rect 6925 -1070 6955 -1040
rect 6925 -1140 6955 -1110
rect 6925 -1210 6955 -1180
rect 6925 -1280 6955 -1250
rect 6925 -1345 6955 -1315
rect 7275 195 7305 225
rect 7275 130 7305 160
rect 7275 60 7305 90
rect 7275 -10 7305 20
rect 7275 -80 7305 -50
rect 7275 -145 7305 -115
rect 7275 -205 7305 -175
rect 7275 -270 7305 -240
rect 7275 -340 7305 -310
rect 7275 -410 7305 -380
rect 7275 -480 7305 -450
rect 7275 -545 7305 -515
rect 7275 -605 7305 -575
rect 7275 -670 7305 -640
rect 7275 -740 7305 -710
rect 7275 -810 7305 -780
rect 7275 -880 7305 -850
rect 7275 -945 7305 -915
rect 7275 -1005 7305 -975
rect 7275 -1070 7305 -1040
rect 7275 -1140 7305 -1110
rect 7275 -1210 7305 -1180
rect 7275 -1280 7305 -1250
rect 7275 -1345 7305 -1315
rect 7625 195 7655 225
rect 7625 130 7655 160
rect 7625 60 7655 90
rect 7625 -10 7655 20
rect 7625 -80 7655 -50
rect 7625 -145 7655 -115
rect 7625 -205 7655 -175
rect 7625 -270 7655 -240
rect 7625 -340 7655 -310
rect 7625 -410 7655 -380
rect 7625 -480 7655 -450
rect 7625 -545 7655 -515
rect 7625 -605 7655 -575
rect 7625 -670 7655 -640
rect 7625 -740 7655 -710
rect 7625 -810 7655 -780
rect 7625 -880 7655 -850
rect 7625 -945 7655 -915
rect 7625 -1005 7655 -975
rect 7625 -1070 7655 -1040
rect 7625 -1140 7655 -1110
rect 7625 -1210 7655 -1180
rect 7625 -1280 7655 -1250
rect 7625 -1345 7655 -1315
rect 7975 195 8005 225
rect 7975 130 8005 160
rect 7975 60 8005 90
rect 7975 -10 8005 20
rect 7975 -80 8005 -50
rect 7975 -145 8005 -115
rect 7975 -205 8005 -175
rect 7975 -270 8005 -240
rect 7975 -340 8005 -310
rect 7975 -410 8005 -380
rect 7975 -480 8005 -450
rect 7975 -545 8005 -515
rect 7975 -605 8005 -575
rect 7975 -670 8005 -640
rect 7975 -740 8005 -710
rect 7975 -810 8005 -780
rect 7975 -880 8005 -850
rect 7975 -945 8005 -915
rect 7975 -1005 8005 -975
rect 7975 -1070 8005 -1040
rect 7975 -1140 8005 -1110
rect 7975 -1210 8005 -1180
rect 7975 -1280 8005 -1250
rect 7975 -1345 8005 -1315
rect 8325 195 8355 225
rect 8325 130 8355 160
rect 8325 60 8355 90
rect 8325 -10 8355 20
rect 8325 -80 8355 -50
rect 8325 -145 8355 -115
rect 8325 -205 8355 -175
rect 8325 -270 8355 -240
rect 8325 -340 8355 -310
rect 8325 -410 8355 -380
rect 8325 -480 8355 -450
rect 8325 -545 8355 -515
rect 8325 -605 8355 -575
rect 8325 -670 8355 -640
rect 8325 -740 8355 -710
rect 8325 -810 8355 -780
rect 8325 -880 8355 -850
rect 8325 -945 8355 -915
rect 8325 -1005 8355 -975
rect 8325 -1070 8355 -1040
rect 8325 -1140 8355 -1110
rect 8325 -1210 8355 -1180
rect 8325 -1280 8355 -1250
rect 8325 -1345 8355 -1315
rect 8675 195 8705 225
rect 8675 130 8705 160
rect 8675 60 8705 90
rect 8675 -10 8705 20
rect 8675 -80 8705 -50
rect 8675 -145 8705 -115
rect 8675 -205 8705 -175
rect 8675 -270 8705 -240
rect 8675 -340 8705 -310
rect 8675 -410 8705 -380
rect 8675 -480 8705 -450
rect 8675 -545 8705 -515
rect 8675 -605 8705 -575
rect 8675 -670 8705 -640
rect 8675 -740 8705 -710
rect 8675 -810 8705 -780
rect 8675 -880 8705 -850
rect 8675 -945 8705 -915
rect 8675 -1005 8705 -975
rect 8675 -1070 8705 -1040
rect 8675 -1140 8705 -1110
rect 8675 -1210 8705 -1180
rect 8675 -1280 8705 -1250
rect 8675 -1345 8705 -1315
rect 9025 195 9055 225
rect 9025 130 9055 160
rect 9025 60 9055 90
rect 9025 -10 9055 20
rect 9025 -80 9055 -50
rect 9025 -145 9055 -115
rect 9025 -205 9055 -175
rect 9025 -270 9055 -240
rect 9025 -340 9055 -310
rect 9025 -410 9055 -380
rect 9025 -480 9055 -450
rect 9025 -545 9055 -515
rect 9025 -605 9055 -575
rect 9025 -670 9055 -640
rect 9025 -740 9055 -710
rect 9025 -810 9055 -780
rect 9025 -880 9055 -850
rect 9025 -945 9055 -915
rect 9025 -1005 9055 -975
rect 9025 -1070 9055 -1040
rect 9025 -1140 9055 -1110
rect 9025 -1210 9055 -1180
rect 9025 -1280 9055 -1250
rect 9025 -1345 9055 -1315
<< metal2 >>
rect 2100 19310 2160 19325
rect 2100 19280 2115 19310
rect 2145 19280 2160 19310
rect 2100 19245 2160 19280
rect 2100 19215 2115 19245
rect 2145 19215 2160 19245
rect 2100 19175 2160 19215
rect 2100 19145 2115 19175
rect 2145 19145 2160 19175
rect 2100 19105 2160 19145
rect 2100 19075 2115 19105
rect 2145 19075 2160 19105
rect 2100 19035 2160 19075
rect 2100 19005 2115 19035
rect 2145 19005 2160 19035
rect 2100 18970 2160 19005
rect 2100 18940 2115 18970
rect 2145 18940 2160 18970
rect 2100 18910 2160 18940
rect 2100 18880 2115 18910
rect 2145 18880 2160 18910
rect 2100 18845 2160 18880
rect 2100 18815 2115 18845
rect 2145 18815 2160 18845
rect 2100 18775 2160 18815
rect 2100 18745 2115 18775
rect 2145 18745 2160 18775
rect 2100 18705 2160 18745
rect 2100 18675 2115 18705
rect 2145 18675 2160 18705
rect 2100 18635 2160 18675
rect 2100 18605 2115 18635
rect 2145 18605 2160 18635
rect 2100 18570 2160 18605
rect 2100 18540 2115 18570
rect 2145 18540 2160 18570
rect 2100 18510 2160 18540
rect 2100 18480 2115 18510
rect 2145 18480 2160 18510
rect 2100 18445 2160 18480
rect 2100 18415 2115 18445
rect 2145 18415 2160 18445
rect 2100 18375 2160 18415
rect 2100 18345 2115 18375
rect 2145 18345 2160 18375
rect 2100 18305 2160 18345
rect 2100 18275 2115 18305
rect 2145 18275 2160 18305
rect 2100 18235 2160 18275
rect 2100 18205 2115 18235
rect 2145 18205 2160 18235
rect 2100 18170 2160 18205
rect 2100 18140 2115 18170
rect 2145 18140 2160 18170
rect 2100 18110 2160 18140
rect 2100 18080 2115 18110
rect 2145 18080 2160 18110
rect 2100 18045 2160 18080
rect 2100 18015 2115 18045
rect 2145 18015 2160 18045
rect 2100 17975 2160 18015
rect 2100 17945 2115 17975
rect 2145 17945 2160 17975
rect 2100 17905 2160 17945
rect 2100 17875 2115 17905
rect 2145 17875 2160 17905
rect 2100 17835 2160 17875
rect 2100 17805 2115 17835
rect 2145 17805 2160 17835
rect 2100 17770 2160 17805
rect 2100 17740 2115 17770
rect 2145 17740 2160 17770
rect 2100 17725 2160 17740
rect 6690 19310 6750 19325
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2205 15925 2325 15930
rect 2205 15895 2210 15925
rect 2240 15895 2250 15925
rect 2280 15895 2290 15925
rect 2320 15920 2325 15925
rect 2320 15900 2385 15920
rect 2320 15895 2325 15900
rect 2205 15890 2325 15895
rect 2070 15690 2970 15695
rect 2070 15660 2075 15690
rect 2105 15660 2115 15690
rect 2145 15660 2155 15690
rect 2185 15660 2970 15690
rect 2070 15650 2970 15660
rect 2070 15620 2075 15650
rect 2105 15620 2115 15650
rect 2145 15620 2155 15650
rect 2185 15620 2970 15650
rect 2070 15610 2970 15620
rect 2070 15580 2075 15610
rect 2105 15580 2115 15610
rect 2145 15580 2155 15610
rect 2185 15580 2970 15610
rect 2070 15575 2970 15580
rect 6650 15595 6780 15600
rect 6650 15565 6665 15595
rect 6695 15565 6705 15595
rect 6735 15565 6745 15595
rect 6775 15565 6780 15595
rect 6650 15555 6780 15565
rect 6650 15525 6665 15555
rect 6695 15525 6705 15555
rect 6735 15525 6745 15555
rect 6775 15525 6780 15555
rect 6650 15515 6780 15525
rect 6650 15485 6665 15515
rect 6695 15485 6705 15515
rect 6735 15485 6745 15515
rect 6775 15485 6780 15515
rect 6650 15480 6780 15485
rect 5690 12925 6780 12930
rect 5690 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6745 12925
rect 6775 12895 6780 12925
rect 5690 12885 6780 12895
rect 5690 12855 6665 12885
rect 6695 12855 6705 12885
rect 6735 12855 6745 12885
rect 6775 12855 6780 12885
rect 5690 12845 6780 12855
rect 5690 12815 6665 12845
rect 6695 12815 6705 12845
rect 6735 12815 6745 12845
rect 6775 12815 6780 12845
rect 5690 12810 6780 12815
rect 2070 12710 3355 12715
rect 2070 12680 2075 12710
rect 2105 12680 2115 12710
rect 2145 12680 2155 12710
rect 2185 12680 3355 12710
rect 2070 12670 3355 12680
rect 2070 12640 2075 12670
rect 2105 12640 2115 12670
rect 2145 12640 2155 12670
rect 2185 12640 3355 12670
rect 2070 12635 3355 12640
rect 2070 12550 3800 12555
rect 2070 12520 2075 12550
rect 2105 12520 2115 12550
rect 2145 12520 2155 12550
rect 2185 12520 3800 12550
rect 2070 12510 3800 12520
rect 2070 12480 2075 12510
rect 2105 12480 2115 12510
rect 2145 12480 2155 12510
rect 2185 12480 3800 12510
rect 2070 12470 3800 12480
rect 2070 12440 2075 12470
rect 2105 12440 2115 12470
rect 2145 12440 2155 12470
rect 2185 12440 3800 12470
rect 2070 12435 3800 12440
rect 5670 12150 6780 12155
rect 5670 12120 6665 12150
rect 6695 12120 6705 12150
rect 6735 12120 6745 12150
rect 6775 12120 6780 12150
rect 5670 12110 6780 12120
rect 5670 12080 6665 12110
rect 6695 12080 6705 12110
rect 6735 12080 6745 12110
rect 6775 12080 6780 12110
rect 5670 12070 6780 12080
rect 5670 12040 6665 12070
rect 6695 12040 6705 12070
rect 6735 12040 6745 12070
rect 6775 12040 6780 12070
rect 5670 12035 6780 12040
rect 5870 11165 6780 11170
rect 5870 11135 6665 11165
rect 6695 11135 6705 11165
rect 6735 11135 6745 11165
rect 6775 11135 6780 11165
rect 5870 11125 6780 11135
rect 5870 11095 6665 11125
rect 6695 11095 6705 11125
rect 6735 11095 6745 11125
rect 6775 11095 6780 11125
rect 5870 11085 6780 11095
rect 5870 11055 6665 11085
rect 6695 11055 6705 11085
rect 6735 11055 6745 11085
rect 6775 11055 6780 11085
rect 5870 11050 6780 11055
rect 5855 10440 6780 10445
rect 5855 10410 6665 10440
rect 6695 10410 6705 10440
rect 6735 10410 6745 10440
rect 6775 10410 6780 10440
rect 5855 10400 6780 10410
rect 5855 10370 6665 10400
rect 6695 10370 6705 10400
rect 6735 10370 6745 10400
rect 6775 10370 6780 10400
rect 5855 10360 6780 10370
rect 5855 10330 6665 10360
rect 6695 10330 6705 10360
rect 6735 10330 6745 10360
rect 6775 10330 6780 10360
rect 5855 10325 6780 10330
rect 5925 10080 6780 10085
rect 5925 10050 6665 10080
rect 6695 10050 6705 10080
rect 6735 10050 6745 10080
rect 6775 10050 6780 10080
rect 5925 10040 6780 10050
rect 5925 10010 6665 10040
rect 6695 10010 6705 10040
rect 6735 10010 6745 10040
rect 6775 10010 6780 10040
rect 5925 10000 6780 10010
rect 5925 9970 6665 10000
rect 6695 9970 6705 10000
rect 6735 9970 6745 10000
rect 6775 9970 6780 10000
rect 5925 9965 6780 9970
rect 1310 9635 1370 9650
rect 1310 9605 1325 9635
rect 1355 9605 1370 9635
rect 1310 9570 1370 9605
rect 1310 9540 1325 9570
rect 1355 9540 1370 9570
rect 1310 9500 1370 9540
rect 1310 9470 1325 9500
rect 1355 9470 1370 9500
rect 1310 9430 1370 9470
rect 1310 9400 1325 9430
rect 1355 9400 1370 9430
rect 1310 9360 1370 9400
rect 1310 9330 1325 9360
rect 1355 9330 1370 9360
rect 1310 9295 1370 9330
rect 1310 9265 1325 9295
rect 1355 9265 1370 9295
rect 1310 9235 1370 9265
rect 1310 9205 1325 9235
rect 1355 9205 1370 9235
rect 1310 9170 1370 9205
rect 1310 9140 1325 9170
rect 1355 9140 1370 9170
rect 1310 9100 1370 9140
rect 1310 9070 1325 9100
rect 1355 9070 1370 9100
rect 1310 9030 1370 9070
rect 1310 9000 1325 9030
rect 1355 9000 1370 9030
rect 1310 8960 1370 9000
rect 1310 8930 1325 8960
rect 1355 8930 1370 8960
rect 1310 8895 1370 8930
rect 1310 8865 1325 8895
rect 1355 8865 1370 8895
rect 1310 8835 1370 8865
rect 1310 8805 1325 8835
rect 1355 8805 1370 8835
rect 1310 8770 1370 8805
rect 1310 8740 1325 8770
rect 1355 8740 1370 8770
rect 1310 8700 1370 8740
rect 1310 8670 1325 8700
rect 1355 8670 1370 8700
rect 1310 8630 1370 8670
rect 1310 8600 1325 8630
rect 1355 8600 1370 8630
rect 1310 8560 1370 8600
rect 1310 8530 1325 8560
rect 1355 8530 1370 8560
rect 1310 8495 1370 8530
rect 1310 8465 1325 8495
rect 1355 8465 1370 8495
rect 1310 8435 1370 8465
rect 1310 8405 1325 8435
rect 1355 8405 1370 8435
rect 1310 8370 1370 8405
rect 1310 8340 1325 8370
rect 1355 8340 1370 8370
rect 1310 8300 1370 8340
rect 1310 8270 1325 8300
rect 1355 8270 1370 8300
rect 1310 8230 1370 8270
rect 1310 8200 1325 8230
rect 1355 8200 1370 8230
rect 1310 8160 1370 8200
rect 1310 8130 1325 8160
rect 1355 8130 1370 8160
rect 1310 8105 1370 8130
rect 2235 9635 2295 9650
rect 2235 9605 2250 9635
rect 2280 9605 2295 9635
rect 2235 9570 2295 9605
rect 2235 9540 2250 9570
rect 2280 9540 2295 9570
rect 2235 9500 2295 9540
rect 2235 9470 2250 9500
rect 2280 9470 2295 9500
rect 2235 9430 2295 9470
rect 2235 9400 2250 9430
rect 2280 9400 2295 9430
rect 2235 9360 2295 9400
rect 2235 9330 2250 9360
rect 2280 9330 2295 9360
rect 2235 9295 2295 9330
rect 2235 9265 2250 9295
rect 2280 9265 2295 9295
rect 2235 9235 2295 9265
rect 2235 9205 2250 9235
rect 2280 9205 2295 9235
rect 2235 9170 2295 9205
rect 2235 9140 2250 9170
rect 2280 9140 2295 9170
rect 2235 9100 2295 9140
rect 2235 9070 2250 9100
rect 2280 9070 2295 9100
rect 2235 9030 2295 9070
rect 2235 9000 2250 9030
rect 2280 9000 2295 9030
rect 2235 8960 2295 9000
rect 2235 8930 2250 8960
rect 2280 8930 2295 8960
rect 2235 8895 2295 8930
rect 2235 8865 2250 8895
rect 2280 8865 2295 8895
rect 2235 8835 2295 8865
rect 2235 8805 2250 8835
rect 2280 8805 2295 8835
rect 2235 8770 2295 8805
rect 2235 8740 2250 8770
rect 2280 8740 2295 8770
rect 2235 8700 2295 8740
rect 2235 8670 2250 8700
rect 2280 8670 2295 8700
rect 2235 8630 2295 8670
rect 2235 8600 2250 8630
rect 2280 8600 2295 8630
rect 2235 8560 2295 8600
rect 2235 8530 2250 8560
rect 2280 8530 2295 8560
rect 2235 8495 2295 8530
rect 2235 8465 2250 8495
rect 2280 8465 2295 8495
rect 2235 8435 2295 8465
rect 2235 8405 2250 8435
rect 2280 8405 2295 8435
rect 2235 8370 2295 8405
rect 2235 8340 2250 8370
rect 2280 8340 2295 8370
rect 2235 8300 2295 8340
rect 2235 8270 2250 8300
rect 2280 8270 2295 8300
rect 2235 8230 2295 8270
rect 2235 8200 2250 8230
rect 2280 8200 2295 8230
rect 2235 8160 2295 8200
rect 2235 8130 2250 8160
rect 2280 8130 2295 8160
rect 2235 8105 2295 8130
rect 3165 9635 3225 9650
rect 3165 9605 3180 9635
rect 3210 9605 3225 9635
rect 3165 9570 3225 9605
rect 3165 9540 3180 9570
rect 3210 9540 3225 9570
rect 3165 9500 3225 9540
rect 3165 9470 3180 9500
rect 3210 9470 3225 9500
rect 3165 9430 3225 9470
rect 3165 9400 3180 9430
rect 3210 9400 3225 9430
rect 3165 9360 3225 9400
rect 3165 9330 3180 9360
rect 3210 9330 3225 9360
rect 3165 9295 3225 9330
rect 3165 9265 3180 9295
rect 3210 9265 3225 9295
rect 3165 9235 3225 9265
rect 3165 9205 3180 9235
rect 3210 9205 3225 9235
rect 3165 9170 3225 9205
rect 3165 9140 3180 9170
rect 3210 9140 3225 9170
rect 3165 9100 3225 9140
rect 3165 9070 3180 9100
rect 3210 9070 3225 9100
rect 3165 9030 3225 9070
rect 3165 9000 3180 9030
rect 3210 9000 3225 9030
rect 3165 8960 3225 9000
rect 3165 8930 3180 8960
rect 3210 8930 3225 8960
rect 3165 8895 3225 8930
rect 3165 8865 3180 8895
rect 3210 8865 3225 8895
rect 3165 8835 3225 8865
rect 3165 8805 3180 8835
rect 3210 8805 3225 8835
rect 3165 8770 3225 8805
rect 3165 8740 3180 8770
rect 3210 8740 3225 8770
rect 3165 8700 3225 8740
rect 3165 8670 3180 8700
rect 3210 8670 3225 8700
rect 3165 8630 3225 8670
rect 3165 8600 3180 8630
rect 3210 8600 3225 8630
rect 3165 8560 3225 8600
rect 3165 8530 3180 8560
rect 3210 8530 3225 8560
rect 3165 8495 3225 8530
rect 3165 8465 3180 8495
rect 3210 8465 3225 8495
rect 3165 8435 3225 8465
rect 3165 8405 3180 8435
rect 3210 8405 3225 8435
rect 3165 8370 3225 8405
rect 3165 8340 3180 8370
rect 3210 8340 3225 8370
rect 3165 8300 3225 8340
rect 3165 8270 3180 8300
rect 3210 8270 3225 8300
rect 3165 8230 3225 8270
rect 3165 8200 3180 8230
rect 3210 8200 3225 8230
rect 3165 8160 3225 8200
rect 3165 8130 3180 8160
rect 3210 8130 3225 8160
rect 3165 8105 3225 8130
rect 6690 9635 6750 9650
rect 6690 9605 6705 9635
rect 6735 9605 6750 9635
rect 6690 9570 6750 9605
rect 6690 9540 6705 9570
rect 6735 9540 6750 9570
rect 6690 9500 6750 9540
rect 6690 9470 6705 9500
rect 6735 9470 6750 9500
rect 6690 9430 6750 9470
rect 6690 9400 6705 9430
rect 6735 9400 6750 9430
rect 6690 9360 6750 9400
rect 6690 9330 6705 9360
rect 6735 9330 6750 9360
rect 6690 9295 6750 9330
rect 6690 9265 6705 9295
rect 6735 9265 6750 9295
rect 6690 9235 6750 9265
rect 6690 9205 6705 9235
rect 6735 9205 6750 9235
rect 6690 9170 6750 9205
rect 6690 9140 6705 9170
rect 6735 9140 6750 9170
rect 6690 9100 6750 9140
rect 6690 9070 6705 9100
rect 6735 9070 6750 9100
rect 6690 9030 6750 9070
rect 6690 9000 6705 9030
rect 6735 9000 6750 9030
rect 6690 8960 6750 9000
rect 6690 8930 6705 8960
rect 6735 8930 6750 8960
rect 6690 8895 6750 8930
rect 6690 8865 6705 8895
rect 6735 8865 6750 8895
rect 6690 8835 6750 8865
rect 6690 8805 6705 8835
rect 6735 8805 6750 8835
rect 6690 8770 6750 8805
rect 6690 8740 6705 8770
rect 6735 8740 6750 8770
rect 6690 8700 6750 8740
rect 6690 8670 6705 8700
rect 6735 8670 6750 8700
rect 6690 8630 6750 8670
rect 6690 8600 6705 8630
rect 6735 8600 6750 8630
rect 6690 8560 6750 8600
rect 6690 8530 6705 8560
rect 6735 8530 6750 8560
rect 6690 8495 6750 8530
rect 6690 8465 6705 8495
rect 6735 8465 6750 8495
rect 6690 8435 6750 8465
rect 6690 8405 6705 8435
rect 6735 8405 6750 8435
rect 6690 8370 6750 8405
rect 6690 8340 6705 8370
rect 6735 8340 6750 8370
rect 6690 8300 6750 8340
rect 6690 8270 6705 8300
rect 6735 8270 6750 8300
rect 6690 8230 6750 8270
rect 6690 8200 6705 8230
rect 6735 8200 6750 8230
rect 6690 8160 6750 8200
rect 6690 8130 6705 8160
rect 6735 8130 6750 8160
rect 6690 8105 6750 8130
rect 7610 9635 7670 9650
rect 7610 9605 7625 9635
rect 7655 9605 7670 9635
rect 7610 9570 7670 9605
rect 7610 9540 7625 9570
rect 7655 9540 7670 9570
rect 7610 9500 7670 9540
rect 7610 9470 7625 9500
rect 7655 9470 7670 9500
rect 7610 9430 7670 9470
rect 7610 9400 7625 9430
rect 7655 9400 7670 9430
rect 7610 9360 7670 9400
rect 7610 9330 7625 9360
rect 7655 9330 7670 9360
rect 7610 9295 7670 9330
rect 7610 9265 7625 9295
rect 7655 9265 7670 9295
rect 7610 9235 7670 9265
rect 7610 9205 7625 9235
rect 7655 9205 7670 9235
rect 7610 9170 7670 9205
rect 7610 9140 7625 9170
rect 7655 9140 7670 9170
rect 7610 9100 7670 9140
rect 7610 9070 7625 9100
rect 7655 9070 7670 9100
rect 7610 9030 7670 9070
rect 7610 9000 7625 9030
rect 7655 9000 7670 9030
rect 7610 8960 7670 9000
rect 7610 8930 7625 8960
rect 7655 8930 7670 8960
rect 7610 8895 7670 8930
rect 7610 8865 7625 8895
rect 7655 8865 7670 8895
rect 7610 8835 7670 8865
rect 7610 8805 7625 8835
rect 7655 8805 7670 8835
rect 7610 8770 7670 8805
rect 7610 8740 7625 8770
rect 7655 8740 7670 8770
rect 7610 8700 7670 8740
rect 7610 8670 7625 8700
rect 7655 8670 7670 8700
rect 7610 8630 7670 8670
rect 7610 8600 7625 8630
rect 7655 8600 7670 8630
rect 7610 8560 7670 8600
rect 7610 8530 7625 8560
rect 7655 8530 7670 8560
rect 7610 8495 7670 8530
rect 7610 8465 7625 8495
rect 7655 8465 7670 8495
rect 7610 8435 7670 8465
rect 7610 8405 7625 8435
rect 7655 8405 7670 8435
rect 7610 8370 7670 8405
rect 7610 8340 7625 8370
rect 7655 8340 7670 8370
rect 7610 8300 7670 8340
rect 7610 8270 7625 8300
rect 7655 8270 7670 8300
rect 7610 8230 7670 8270
rect 7610 8200 7625 8230
rect 7655 8200 7670 8230
rect 7610 8160 7670 8200
rect 7610 8130 7625 8160
rect 7655 8130 7670 8160
rect 7610 8105 7670 8130
rect 1980 8070 2515 8075
rect 1980 8040 1985 8070
rect 2015 8040 2025 8070
rect 2055 8040 2065 8070
rect 2095 8040 2480 8070
rect 2510 8040 2515 8070
rect 1980 8035 2515 8040
rect 6465 8070 7000 8075
rect 6465 8040 6470 8070
rect 6500 8040 6885 8070
rect 6915 8040 6925 8070
rect 6955 8040 6965 8070
rect 6995 8040 7000 8070
rect 6465 8035 7000 8040
rect 1630 8015 3890 8020
rect 1630 7985 1635 8015
rect 1665 7985 1675 8015
rect 1705 7985 1715 8015
rect 1745 7985 3635 8015
rect 3665 7985 3855 8015
rect 3885 7985 3890 8015
rect 1630 7980 3890 7985
rect 5090 8015 7350 8020
rect 5090 7985 5095 8015
rect 5125 7985 5315 8015
rect 5345 7985 7235 8015
rect 7265 7985 7275 8015
rect 7305 7985 7315 8015
rect 7345 7985 7350 8015
rect 5090 7980 7350 7985
rect 2845 7960 2885 7965
rect 2845 7930 2850 7960
rect 2880 7955 2885 7960
rect 3385 7960 3420 7965
rect 2880 7935 3385 7955
rect 2880 7930 2885 7935
rect 2845 7925 2885 7930
rect 3415 7930 3420 7960
rect 3385 7925 3420 7930
rect 5470 7960 5510 7965
rect 5470 7930 5475 7960
rect 5505 7955 5510 7960
rect 6145 7960 6185 7965
rect 6145 7955 6150 7960
rect 5505 7935 6150 7955
rect 5505 7930 5510 7935
rect 5470 7925 5510 7930
rect 6145 7930 6150 7935
rect 6180 7930 6185 7960
rect 6145 7925 6185 7930
rect 3290 7870 5585 7875
rect 2715 7850 2755 7855
rect 2715 7820 2720 7850
rect 2750 7845 2755 7850
rect 3075 7850 3115 7855
rect 3075 7845 3080 7850
rect 2750 7825 3080 7845
rect 2750 7820 2755 7825
rect 2715 7815 2755 7820
rect 3075 7820 3080 7825
rect 3110 7820 3115 7850
rect 3075 7815 3115 7820
rect 3290 7840 3295 7870
rect 3325 7840 3440 7870
rect 3470 7840 5550 7870
rect 5580 7840 5585 7870
rect 3290 7830 5585 7840
rect 3290 7800 3295 7830
rect 3325 7800 3440 7830
rect 3470 7800 5550 7830
rect 5580 7800 5585 7830
rect 3290 7790 5585 7800
rect 3290 7760 3295 7790
rect 3325 7760 3440 7790
rect 3470 7760 5550 7790
rect 5580 7760 5585 7790
rect 3290 7755 5585 7760
rect 930 7735 8050 7740
rect 930 7705 935 7735
rect 965 7705 975 7735
rect 1005 7705 1015 7735
rect 1045 7705 4310 7735
rect 4340 7705 4420 7735
rect 4450 7705 4530 7735
rect 4560 7705 4640 7735
rect 4670 7705 7935 7735
rect 7965 7705 7975 7735
rect 8005 7705 8015 7735
rect 8045 7705 8050 7735
rect 930 7695 8050 7705
rect 930 7665 935 7695
rect 965 7665 975 7695
rect 1005 7665 1015 7695
rect 1045 7665 4310 7695
rect 4340 7665 4420 7695
rect 4450 7665 4530 7695
rect 4560 7665 4640 7695
rect 4670 7665 7935 7695
rect 7965 7665 7975 7695
rect 8005 7665 8015 7695
rect 8045 7665 8050 7695
rect 930 7655 8050 7665
rect 930 7625 935 7655
rect 965 7625 975 7655
rect 1005 7625 1015 7655
rect 1045 7625 4310 7655
rect 4340 7625 4420 7655
rect 4450 7625 4530 7655
rect 4560 7625 4640 7655
rect 4670 7625 7935 7655
rect 7965 7625 7975 7655
rect 8005 7625 8015 7655
rect 8045 7625 8050 7655
rect 930 7620 8050 7625
rect 5870 6965 6260 6970
rect 5870 6935 5875 6965
rect 5905 6935 6225 6965
rect 6255 6935 6260 6965
rect 5870 6930 6260 6935
rect 3075 6620 3115 6625
rect 3075 6590 3080 6620
rect 3110 6590 3115 6620
rect 3075 6585 3115 6590
rect 5620 6565 5910 6570
rect 5620 6535 5625 6565
rect 5655 6535 5875 6565
rect 5905 6535 5910 6565
rect 5620 6530 5910 6535
rect 5620 5970 5660 5975
rect 5620 5940 5625 5970
rect 5655 5940 5660 5970
rect 5620 5935 5660 5940
rect 5475 5395 5505 5400
rect 4720 5370 5475 5390
rect 5475 5360 5505 5365
rect 3380 5335 3420 5340
rect 3380 5305 3385 5335
rect 3415 5330 3420 5335
rect 3415 5310 3955 5330
rect 3415 5305 3420 5310
rect 3380 5300 3420 5305
rect 3435 4655 5585 4660
rect 3435 4625 3440 4655
rect 3470 4625 4475 4655
rect 4505 4625 5550 4655
rect 5580 4625 5585 4655
rect 3435 4620 5585 4625
rect 4470 4435 4510 4440
rect 4470 4405 4475 4435
rect 4505 4405 4510 4435
rect 4470 4400 4510 4405
rect 2045 3840 2085 3850
rect 2120 3840 2160 3850
rect 2045 3820 2160 3840
rect 2045 3810 2085 3820
rect 2120 3810 2160 3820
rect 2000 3785 2040 3795
rect 2075 3785 2115 3795
rect 2000 3765 2115 3785
rect 2000 3755 2040 3765
rect 2075 3755 2115 3765
rect 3605 3125 3625 3145
rect 5355 3125 5375 3145
rect 930 2690 8050 2695
rect 930 2660 935 2690
rect 965 2660 975 2690
rect 1005 2660 1015 2690
rect 1045 2660 4420 2690
rect 4450 2660 4530 2690
rect 4560 2660 7935 2690
rect 7965 2660 7975 2690
rect 8005 2660 8015 2690
rect 8045 2660 8050 2690
rect 930 2650 8050 2660
rect 930 2620 935 2650
rect 965 2620 975 2650
rect 1005 2620 1015 2650
rect 1045 2620 4420 2650
rect 4450 2620 4530 2650
rect 4560 2620 7935 2650
rect 7965 2620 7975 2650
rect 8005 2620 8015 2650
rect 8045 2620 8050 2650
rect 930 2610 8050 2620
rect 930 2580 935 2610
rect 965 2580 975 2610
rect 1005 2580 1015 2610
rect 1045 2580 4420 2610
rect 4450 2580 4530 2610
rect 4560 2580 7935 2610
rect 7965 2580 7975 2610
rect 8005 2580 8015 2610
rect 8045 2580 8050 2610
rect 930 2575 8050 2580
rect 2175 2385 2195 2405
rect 6785 2385 6805 2405
rect -90 225 -30 240
rect -90 195 -75 225
rect -45 195 -30 225
rect -90 160 -30 195
rect -90 130 -75 160
rect -45 130 -30 160
rect -90 90 -30 130
rect -90 60 -75 90
rect -45 60 -30 90
rect -90 20 -30 60
rect -90 -10 -75 20
rect -45 -10 -30 20
rect -90 -50 -30 -10
rect -90 -80 -75 -50
rect -45 -80 -30 -50
rect -90 -115 -30 -80
rect -90 -145 -75 -115
rect -45 -145 -30 -115
rect -90 -175 -30 -145
rect -90 -205 -75 -175
rect -45 -205 -30 -175
rect -90 -240 -30 -205
rect -90 -270 -75 -240
rect -45 -270 -30 -240
rect -90 -310 -30 -270
rect -90 -340 -75 -310
rect -45 -340 -30 -310
rect -90 -380 -30 -340
rect -90 -410 -75 -380
rect -45 -410 -30 -380
rect -90 -450 -30 -410
rect -90 -480 -75 -450
rect -45 -480 -30 -450
rect -90 -515 -30 -480
rect -90 -545 -75 -515
rect -45 -545 -30 -515
rect -90 -575 -30 -545
rect -90 -605 -75 -575
rect -45 -605 -30 -575
rect -90 -640 -30 -605
rect -90 -670 -75 -640
rect -45 -670 -30 -640
rect -90 -710 -30 -670
rect -90 -740 -75 -710
rect -45 -740 -30 -710
rect -90 -780 -30 -740
rect -90 -810 -75 -780
rect -45 -810 -30 -780
rect -90 -850 -30 -810
rect -90 -880 -75 -850
rect -45 -880 -30 -850
rect -90 -915 -30 -880
rect -90 -945 -75 -915
rect -45 -945 -30 -915
rect -90 -975 -30 -945
rect -90 -1005 -75 -975
rect -45 -1005 -30 -975
rect -90 -1040 -30 -1005
rect -90 -1070 -75 -1040
rect -45 -1070 -30 -1040
rect -90 -1110 -30 -1070
rect -90 -1140 -75 -1110
rect -45 -1140 -30 -1110
rect -90 -1180 -30 -1140
rect -90 -1210 -75 -1180
rect -45 -1210 -30 -1180
rect -90 -1250 -30 -1210
rect -90 -1280 -75 -1250
rect -45 -1280 -30 -1250
rect -90 -1315 -30 -1280
rect -90 -1345 -75 -1315
rect -45 -1345 -30 -1315
rect -90 -1360 -30 -1345
rect 260 225 320 240
rect 260 195 275 225
rect 305 195 320 225
rect 260 160 320 195
rect 260 130 275 160
rect 305 130 320 160
rect 260 90 320 130
rect 260 60 275 90
rect 305 60 320 90
rect 260 20 320 60
rect 260 -10 275 20
rect 305 -10 320 20
rect 260 -50 320 -10
rect 260 -80 275 -50
rect 305 -80 320 -50
rect 260 -115 320 -80
rect 260 -145 275 -115
rect 305 -145 320 -115
rect 260 -175 320 -145
rect 260 -205 275 -175
rect 305 -205 320 -175
rect 260 -240 320 -205
rect 260 -270 275 -240
rect 305 -270 320 -240
rect 260 -310 320 -270
rect 260 -340 275 -310
rect 305 -340 320 -310
rect 260 -380 320 -340
rect 260 -410 275 -380
rect 305 -410 320 -380
rect 260 -450 320 -410
rect 260 -480 275 -450
rect 305 -480 320 -450
rect 260 -515 320 -480
rect 260 -545 275 -515
rect 305 -545 320 -515
rect 260 -575 320 -545
rect 260 -605 275 -575
rect 305 -605 320 -575
rect 260 -640 320 -605
rect 260 -670 275 -640
rect 305 -670 320 -640
rect 260 -710 320 -670
rect 260 -740 275 -710
rect 305 -740 320 -710
rect 260 -780 320 -740
rect 260 -810 275 -780
rect 305 -810 320 -780
rect 260 -850 320 -810
rect 260 -880 275 -850
rect 305 -880 320 -850
rect 260 -915 320 -880
rect 260 -945 275 -915
rect 305 -945 320 -915
rect 260 -975 320 -945
rect 260 -1005 275 -975
rect 305 -1005 320 -975
rect 260 -1040 320 -1005
rect 260 -1070 275 -1040
rect 305 -1070 320 -1040
rect 260 -1110 320 -1070
rect 260 -1140 275 -1110
rect 305 -1140 320 -1110
rect 260 -1180 320 -1140
rect 260 -1210 275 -1180
rect 305 -1210 320 -1180
rect 260 -1250 320 -1210
rect 260 -1280 275 -1250
rect 305 -1280 320 -1250
rect 260 -1315 320 -1280
rect 260 -1345 275 -1315
rect 305 -1345 320 -1315
rect 260 -1360 320 -1345
rect 610 225 670 240
rect 610 195 625 225
rect 655 195 670 225
rect 610 160 670 195
rect 610 130 625 160
rect 655 130 670 160
rect 610 90 670 130
rect 610 60 625 90
rect 655 60 670 90
rect 610 20 670 60
rect 610 -10 625 20
rect 655 -10 670 20
rect 610 -50 670 -10
rect 610 -80 625 -50
rect 655 -80 670 -50
rect 610 -115 670 -80
rect 610 -145 625 -115
rect 655 -145 670 -115
rect 610 -175 670 -145
rect 610 -205 625 -175
rect 655 -205 670 -175
rect 610 -240 670 -205
rect 610 -270 625 -240
rect 655 -270 670 -240
rect 610 -310 670 -270
rect 610 -340 625 -310
rect 655 -340 670 -310
rect 610 -380 670 -340
rect 610 -410 625 -380
rect 655 -410 670 -380
rect 610 -450 670 -410
rect 610 -480 625 -450
rect 655 -480 670 -450
rect 610 -515 670 -480
rect 610 -545 625 -515
rect 655 -545 670 -515
rect 610 -575 670 -545
rect 610 -605 625 -575
rect 655 -605 670 -575
rect 610 -640 670 -605
rect 610 -670 625 -640
rect 655 -670 670 -640
rect 610 -710 670 -670
rect 610 -740 625 -710
rect 655 -740 670 -710
rect 610 -780 670 -740
rect 610 -810 625 -780
rect 655 -810 670 -780
rect 610 -850 670 -810
rect 610 -880 625 -850
rect 655 -880 670 -850
rect 610 -915 670 -880
rect 610 -945 625 -915
rect 655 -945 670 -915
rect 610 -975 670 -945
rect 610 -1005 625 -975
rect 655 -1005 670 -975
rect 610 -1040 670 -1005
rect 610 -1070 625 -1040
rect 655 -1070 670 -1040
rect 610 -1110 670 -1070
rect 610 -1140 625 -1110
rect 655 -1140 670 -1110
rect 610 -1180 670 -1140
rect 610 -1210 625 -1180
rect 655 -1210 670 -1180
rect 610 -1250 670 -1210
rect 610 -1280 625 -1250
rect 655 -1280 670 -1250
rect 610 -1315 670 -1280
rect 610 -1345 625 -1315
rect 655 -1345 670 -1315
rect 610 -1360 670 -1345
rect 960 225 1020 240
rect 960 195 975 225
rect 1005 195 1020 225
rect 960 160 1020 195
rect 960 130 975 160
rect 1005 130 1020 160
rect 960 90 1020 130
rect 960 60 975 90
rect 1005 60 1020 90
rect 960 20 1020 60
rect 960 -10 975 20
rect 1005 -10 1020 20
rect 960 -50 1020 -10
rect 960 -80 975 -50
rect 1005 -80 1020 -50
rect 960 -115 1020 -80
rect 960 -145 975 -115
rect 1005 -145 1020 -115
rect 960 -175 1020 -145
rect 960 -205 975 -175
rect 1005 -205 1020 -175
rect 960 -240 1020 -205
rect 960 -270 975 -240
rect 1005 -270 1020 -240
rect 960 -310 1020 -270
rect 960 -340 975 -310
rect 1005 -340 1020 -310
rect 960 -380 1020 -340
rect 960 -410 975 -380
rect 1005 -410 1020 -380
rect 960 -450 1020 -410
rect 960 -480 975 -450
rect 1005 -480 1020 -450
rect 960 -515 1020 -480
rect 960 -545 975 -515
rect 1005 -545 1020 -515
rect 960 -575 1020 -545
rect 960 -605 975 -575
rect 1005 -605 1020 -575
rect 960 -640 1020 -605
rect 960 -670 975 -640
rect 1005 -670 1020 -640
rect 960 -710 1020 -670
rect 960 -740 975 -710
rect 1005 -740 1020 -710
rect 960 -780 1020 -740
rect 960 -810 975 -780
rect 1005 -810 1020 -780
rect 960 -850 1020 -810
rect 960 -880 975 -850
rect 1005 -880 1020 -850
rect 960 -915 1020 -880
rect 960 -945 975 -915
rect 1005 -945 1020 -915
rect 960 -975 1020 -945
rect 960 -1005 975 -975
rect 1005 -1005 1020 -975
rect 960 -1040 1020 -1005
rect 960 -1070 975 -1040
rect 1005 -1070 1020 -1040
rect 960 -1110 1020 -1070
rect 960 -1140 975 -1110
rect 1005 -1140 1020 -1110
rect 960 -1180 1020 -1140
rect 960 -1210 975 -1180
rect 1005 -1210 1020 -1180
rect 960 -1250 1020 -1210
rect 960 -1280 975 -1250
rect 1005 -1280 1020 -1250
rect 960 -1315 1020 -1280
rect 960 -1345 975 -1315
rect 1005 -1345 1020 -1315
rect 960 -1360 1020 -1345
rect 1310 225 1370 240
rect 1310 195 1325 225
rect 1355 195 1370 225
rect 1310 160 1370 195
rect 1310 130 1325 160
rect 1355 130 1370 160
rect 1310 90 1370 130
rect 1310 60 1325 90
rect 1355 60 1370 90
rect 1310 20 1370 60
rect 1310 -10 1325 20
rect 1355 -10 1370 20
rect 1310 -50 1370 -10
rect 1310 -80 1325 -50
rect 1355 -80 1370 -50
rect 1310 -115 1370 -80
rect 1310 -145 1325 -115
rect 1355 -145 1370 -115
rect 1310 -175 1370 -145
rect 1310 -205 1325 -175
rect 1355 -205 1370 -175
rect 1310 -240 1370 -205
rect 1310 -270 1325 -240
rect 1355 -270 1370 -240
rect 1310 -310 1370 -270
rect 1310 -340 1325 -310
rect 1355 -340 1370 -310
rect 1310 -380 1370 -340
rect 1310 -410 1325 -380
rect 1355 -410 1370 -380
rect 1310 -450 1370 -410
rect 1310 -480 1325 -450
rect 1355 -480 1370 -450
rect 1310 -515 1370 -480
rect 1310 -545 1325 -515
rect 1355 -545 1370 -515
rect 1310 -575 1370 -545
rect 1310 -605 1325 -575
rect 1355 -605 1370 -575
rect 1310 -640 1370 -605
rect 1310 -670 1325 -640
rect 1355 -670 1370 -640
rect 1310 -710 1370 -670
rect 1310 -740 1325 -710
rect 1355 -740 1370 -710
rect 1310 -780 1370 -740
rect 1310 -810 1325 -780
rect 1355 -810 1370 -780
rect 1310 -850 1370 -810
rect 1310 -880 1325 -850
rect 1355 -880 1370 -850
rect 1310 -915 1370 -880
rect 1310 -945 1325 -915
rect 1355 -945 1370 -915
rect 1310 -975 1370 -945
rect 1310 -1005 1325 -975
rect 1355 -1005 1370 -975
rect 1310 -1040 1370 -1005
rect 1310 -1070 1325 -1040
rect 1355 -1070 1370 -1040
rect 1310 -1110 1370 -1070
rect 1310 -1140 1325 -1110
rect 1355 -1140 1370 -1110
rect 1310 -1180 1370 -1140
rect 1310 -1210 1325 -1180
rect 1355 -1210 1370 -1180
rect 1310 -1250 1370 -1210
rect 1310 -1280 1325 -1250
rect 1355 -1280 1370 -1250
rect 1310 -1315 1370 -1280
rect 1310 -1345 1325 -1315
rect 1355 -1345 1370 -1315
rect 1310 -1360 1370 -1345
rect 1660 225 1720 240
rect 1660 195 1675 225
rect 1705 195 1720 225
rect 1660 160 1720 195
rect 1660 130 1675 160
rect 1705 130 1720 160
rect 1660 90 1720 130
rect 1660 60 1675 90
rect 1705 60 1720 90
rect 1660 20 1720 60
rect 1660 -10 1675 20
rect 1705 -10 1720 20
rect 1660 -50 1720 -10
rect 1660 -80 1675 -50
rect 1705 -80 1720 -50
rect 1660 -115 1720 -80
rect 1660 -145 1675 -115
rect 1705 -145 1720 -115
rect 1660 -175 1720 -145
rect 1660 -205 1675 -175
rect 1705 -205 1720 -175
rect 1660 -240 1720 -205
rect 1660 -270 1675 -240
rect 1705 -270 1720 -240
rect 1660 -310 1720 -270
rect 1660 -340 1675 -310
rect 1705 -340 1720 -310
rect 1660 -380 1720 -340
rect 1660 -410 1675 -380
rect 1705 -410 1720 -380
rect 1660 -450 1720 -410
rect 1660 -480 1675 -450
rect 1705 -480 1720 -450
rect 1660 -515 1720 -480
rect 1660 -545 1675 -515
rect 1705 -545 1720 -515
rect 1660 -575 1720 -545
rect 1660 -605 1675 -575
rect 1705 -605 1720 -575
rect 1660 -640 1720 -605
rect 1660 -670 1675 -640
rect 1705 -670 1720 -640
rect 1660 -710 1720 -670
rect 1660 -740 1675 -710
rect 1705 -740 1720 -710
rect 1660 -780 1720 -740
rect 1660 -810 1675 -780
rect 1705 -810 1720 -780
rect 1660 -850 1720 -810
rect 1660 -880 1675 -850
rect 1705 -880 1720 -850
rect 1660 -915 1720 -880
rect 1660 -945 1675 -915
rect 1705 -945 1720 -915
rect 1660 -975 1720 -945
rect 1660 -1005 1675 -975
rect 1705 -1005 1720 -975
rect 1660 -1040 1720 -1005
rect 1660 -1070 1675 -1040
rect 1705 -1070 1720 -1040
rect 1660 -1110 1720 -1070
rect 1660 -1140 1675 -1110
rect 1705 -1140 1720 -1110
rect 1660 -1180 1720 -1140
rect 1660 -1210 1675 -1180
rect 1705 -1210 1720 -1180
rect 1660 -1250 1720 -1210
rect 1660 -1280 1675 -1250
rect 1705 -1280 1720 -1250
rect 1660 -1315 1720 -1280
rect 1660 -1345 1675 -1315
rect 1705 -1345 1720 -1315
rect 1660 -1360 1720 -1345
rect 2010 225 2070 240
rect 2010 195 2025 225
rect 2055 195 2070 225
rect 2010 160 2070 195
rect 2010 130 2025 160
rect 2055 130 2070 160
rect 2010 90 2070 130
rect 2010 60 2025 90
rect 2055 60 2070 90
rect 2010 20 2070 60
rect 2010 -10 2025 20
rect 2055 -10 2070 20
rect 2010 -50 2070 -10
rect 2010 -80 2025 -50
rect 2055 -80 2070 -50
rect 2010 -115 2070 -80
rect 2010 -145 2025 -115
rect 2055 -145 2070 -115
rect 2010 -175 2070 -145
rect 2010 -205 2025 -175
rect 2055 -205 2070 -175
rect 2010 -240 2070 -205
rect 2010 -270 2025 -240
rect 2055 -270 2070 -240
rect 2010 -310 2070 -270
rect 2010 -340 2025 -310
rect 2055 -340 2070 -310
rect 2010 -380 2070 -340
rect 2010 -410 2025 -380
rect 2055 -410 2070 -380
rect 2010 -450 2070 -410
rect 2010 -480 2025 -450
rect 2055 -480 2070 -450
rect 2010 -515 2070 -480
rect 2010 -545 2025 -515
rect 2055 -545 2070 -515
rect 2010 -575 2070 -545
rect 2010 -605 2025 -575
rect 2055 -605 2070 -575
rect 2010 -640 2070 -605
rect 2010 -670 2025 -640
rect 2055 -670 2070 -640
rect 2010 -710 2070 -670
rect 2010 -740 2025 -710
rect 2055 -740 2070 -710
rect 2010 -780 2070 -740
rect 2010 -810 2025 -780
rect 2055 -810 2070 -780
rect 2010 -850 2070 -810
rect 2010 -880 2025 -850
rect 2055 -880 2070 -850
rect 2010 -915 2070 -880
rect 2010 -945 2025 -915
rect 2055 -945 2070 -915
rect 2010 -975 2070 -945
rect 2010 -1005 2025 -975
rect 2055 -1005 2070 -975
rect 2010 -1040 2070 -1005
rect 2010 -1070 2025 -1040
rect 2055 -1070 2070 -1040
rect 2010 -1110 2070 -1070
rect 2010 -1140 2025 -1110
rect 2055 -1140 2070 -1110
rect 2010 -1180 2070 -1140
rect 2010 -1210 2025 -1180
rect 2055 -1210 2070 -1180
rect 2010 -1250 2070 -1210
rect 2010 -1280 2025 -1250
rect 2055 -1280 2070 -1250
rect 2010 -1315 2070 -1280
rect 2010 -1345 2025 -1315
rect 2055 -1345 2070 -1315
rect 2010 -1360 2070 -1345
rect 2360 225 2420 240
rect 2360 195 2375 225
rect 2405 195 2420 225
rect 2360 160 2420 195
rect 2360 130 2375 160
rect 2405 130 2420 160
rect 2360 90 2420 130
rect 2360 60 2375 90
rect 2405 60 2420 90
rect 2360 20 2420 60
rect 2360 -10 2375 20
rect 2405 -10 2420 20
rect 2360 -50 2420 -10
rect 2360 -80 2375 -50
rect 2405 -80 2420 -50
rect 2360 -115 2420 -80
rect 2360 -145 2375 -115
rect 2405 -145 2420 -115
rect 2360 -175 2420 -145
rect 2360 -205 2375 -175
rect 2405 -205 2420 -175
rect 2360 -240 2420 -205
rect 2360 -270 2375 -240
rect 2405 -270 2420 -240
rect 2360 -310 2420 -270
rect 2360 -340 2375 -310
rect 2405 -340 2420 -310
rect 2360 -380 2420 -340
rect 2360 -410 2375 -380
rect 2405 -410 2420 -380
rect 2360 -450 2420 -410
rect 2360 -480 2375 -450
rect 2405 -480 2420 -450
rect 2360 -515 2420 -480
rect 2360 -545 2375 -515
rect 2405 -545 2420 -515
rect 2360 -575 2420 -545
rect 2360 -605 2375 -575
rect 2405 -605 2420 -575
rect 2360 -640 2420 -605
rect 2360 -670 2375 -640
rect 2405 -670 2420 -640
rect 2360 -710 2420 -670
rect 2360 -740 2375 -710
rect 2405 -740 2420 -710
rect 2360 -780 2420 -740
rect 2360 -810 2375 -780
rect 2405 -810 2420 -780
rect 2360 -850 2420 -810
rect 2360 -880 2375 -850
rect 2405 -880 2420 -850
rect 2360 -915 2420 -880
rect 2360 -945 2375 -915
rect 2405 -945 2420 -915
rect 2360 -975 2420 -945
rect 2360 -1005 2375 -975
rect 2405 -1005 2420 -975
rect 2360 -1040 2420 -1005
rect 2360 -1070 2375 -1040
rect 2405 -1070 2420 -1040
rect 2360 -1110 2420 -1070
rect 2360 -1140 2375 -1110
rect 2405 -1140 2420 -1110
rect 2360 -1180 2420 -1140
rect 2360 -1210 2375 -1180
rect 2405 -1210 2420 -1180
rect 2360 -1250 2420 -1210
rect 2360 -1280 2375 -1250
rect 2405 -1280 2420 -1250
rect 2360 -1315 2420 -1280
rect 2360 -1345 2375 -1315
rect 2405 -1345 2420 -1315
rect 2360 -1360 2420 -1345
rect 2710 225 2770 240
rect 2710 195 2725 225
rect 2755 195 2770 225
rect 2710 160 2770 195
rect 2710 130 2725 160
rect 2755 130 2770 160
rect 2710 90 2770 130
rect 2710 60 2725 90
rect 2755 60 2770 90
rect 2710 20 2770 60
rect 2710 -10 2725 20
rect 2755 -10 2770 20
rect 2710 -50 2770 -10
rect 2710 -80 2725 -50
rect 2755 -80 2770 -50
rect 2710 -115 2770 -80
rect 2710 -145 2725 -115
rect 2755 -145 2770 -115
rect 2710 -175 2770 -145
rect 2710 -205 2725 -175
rect 2755 -205 2770 -175
rect 2710 -240 2770 -205
rect 2710 -270 2725 -240
rect 2755 -270 2770 -240
rect 2710 -310 2770 -270
rect 2710 -340 2725 -310
rect 2755 -340 2770 -310
rect 2710 -380 2770 -340
rect 2710 -410 2725 -380
rect 2755 -410 2770 -380
rect 2710 -450 2770 -410
rect 2710 -480 2725 -450
rect 2755 -480 2770 -450
rect 2710 -515 2770 -480
rect 2710 -545 2725 -515
rect 2755 -545 2770 -515
rect 2710 -575 2770 -545
rect 2710 -605 2725 -575
rect 2755 -605 2770 -575
rect 2710 -640 2770 -605
rect 2710 -670 2725 -640
rect 2755 -670 2770 -640
rect 2710 -710 2770 -670
rect 2710 -740 2725 -710
rect 2755 -740 2770 -710
rect 2710 -780 2770 -740
rect 2710 -810 2725 -780
rect 2755 -810 2770 -780
rect 2710 -850 2770 -810
rect 2710 -880 2725 -850
rect 2755 -880 2770 -850
rect 2710 -915 2770 -880
rect 2710 -945 2725 -915
rect 2755 -945 2770 -915
rect 2710 -975 2770 -945
rect 2710 -1005 2725 -975
rect 2755 -1005 2770 -975
rect 2710 -1040 2770 -1005
rect 2710 -1070 2725 -1040
rect 2755 -1070 2770 -1040
rect 2710 -1110 2770 -1070
rect 2710 -1140 2725 -1110
rect 2755 -1140 2770 -1110
rect 2710 -1180 2770 -1140
rect 2710 -1210 2725 -1180
rect 2755 -1210 2770 -1180
rect 2710 -1250 2770 -1210
rect 2710 -1280 2725 -1250
rect 2755 -1280 2770 -1250
rect 2710 -1315 2770 -1280
rect 2710 -1345 2725 -1315
rect 2755 -1345 2770 -1315
rect 2710 -1360 2770 -1345
rect 3060 225 3120 240
rect 3060 195 3075 225
rect 3105 195 3120 225
rect 3060 160 3120 195
rect 3060 130 3075 160
rect 3105 130 3120 160
rect 3060 90 3120 130
rect 3060 60 3075 90
rect 3105 60 3120 90
rect 3060 20 3120 60
rect 3060 -10 3075 20
rect 3105 -10 3120 20
rect 3060 -50 3120 -10
rect 3060 -80 3075 -50
rect 3105 -80 3120 -50
rect 3060 -115 3120 -80
rect 3060 -145 3075 -115
rect 3105 -145 3120 -115
rect 3060 -175 3120 -145
rect 3060 -205 3075 -175
rect 3105 -205 3120 -175
rect 3060 -240 3120 -205
rect 3060 -270 3075 -240
rect 3105 -270 3120 -240
rect 3060 -310 3120 -270
rect 3060 -340 3075 -310
rect 3105 -340 3120 -310
rect 3060 -380 3120 -340
rect 3060 -410 3075 -380
rect 3105 -410 3120 -380
rect 3060 -450 3120 -410
rect 3060 -480 3075 -450
rect 3105 -480 3120 -450
rect 3060 -515 3120 -480
rect 3060 -545 3075 -515
rect 3105 -545 3120 -515
rect 3060 -575 3120 -545
rect 3060 -605 3075 -575
rect 3105 -605 3120 -575
rect 3060 -640 3120 -605
rect 3060 -670 3075 -640
rect 3105 -670 3120 -640
rect 3060 -710 3120 -670
rect 3060 -740 3075 -710
rect 3105 -740 3120 -710
rect 3060 -780 3120 -740
rect 3060 -810 3075 -780
rect 3105 -810 3120 -780
rect 3060 -850 3120 -810
rect 3060 -880 3075 -850
rect 3105 -880 3120 -850
rect 3060 -915 3120 -880
rect 3060 -945 3075 -915
rect 3105 -945 3120 -915
rect 3060 -975 3120 -945
rect 3060 -1005 3075 -975
rect 3105 -1005 3120 -975
rect 3060 -1040 3120 -1005
rect 3060 -1070 3075 -1040
rect 3105 -1070 3120 -1040
rect 3060 -1110 3120 -1070
rect 3060 -1140 3075 -1110
rect 3105 -1140 3120 -1110
rect 3060 -1180 3120 -1140
rect 3060 -1210 3075 -1180
rect 3105 -1210 3120 -1180
rect 3060 -1250 3120 -1210
rect 3060 -1280 3075 -1250
rect 3105 -1280 3120 -1250
rect 3060 -1315 3120 -1280
rect 3060 -1345 3075 -1315
rect 3105 -1345 3120 -1315
rect 3060 -1360 3120 -1345
rect 3410 225 3470 240
rect 3410 195 3425 225
rect 3455 195 3470 225
rect 3410 160 3470 195
rect 3410 130 3425 160
rect 3455 130 3470 160
rect 3410 90 3470 130
rect 3410 60 3425 90
rect 3455 60 3470 90
rect 3410 20 3470 60
rect 3410 -10 3425 20
rect 3455 -10 3470 20
rect 3410 -50 3470 -10
rect 3410 -80 3425 -50
rect 3455 -80 3470 -50
rect 3410 -115 3470 -80
rect 3410 -145 3425 -115
rect 3455 -145 3470 -115
rect 3410 -175 3470 -145
rect 3410 -205 3425 -175
rect 3455 -205 3470 -175
rect 3410 -240 3470 -205
rect 3410 -270 3425 -240
rect 3455 -270 3470 -240
rect 3410 -310 3470 -270
rect 3410 -340 3425 -310
rect 3455 -340 3470 -310
rect 3410 -380 3470 -340
rect 3410 -410 3425 -380
rect 3455 -410 3470 -380
rect 3410 -450 3470 -410
rect 3410 -480 3425 -450
rect 3455 -480 3470 -450
rect 3410 -515 3470 -480
rect 3410 -545 3425 -515
rect 3455 -545 3470 -515
rect 3410 -575 3470 -545
rect 3410 -605 3425 -575
rect 3455 -605 3470 -575
rect 3410 -640 3470 -605
rect 3410 -670 3425 -640
rect 3455 -670 3470 -640
rect 3410 -710 3470 -670
rect 3410 -740 3425 -710
rect 3455 -740 3470 -710
rect 3410 -780 3470 -740
rect 3410 -810 3425 -780
rect 3455 -810 3470 -780
rect 3410 -850 3470 -810
rect 3410 -880 3425 -850
rect 3455 -880 3470 -850
rect 3410 -915 3470 -880
rect 3410 -945 3425 -915
rect 3455 -945 3470 -915
rect 3410 -975 3470 -945
rect 3410 -1005 3425 -975
rect 3455 -1005 3470 -975
rect 3410 -1040 3470 -1005
rect 3410 -1070 3425 -1040
rect 3455 -1070 3470 -1040
rect 3410 -1110 3470 -1070
rect 3410 -1140 3425 -1110
rect 3455 -1140 3470 -1110
rect 3410 -1180 3470 -1140
rect 3410 -1210 3425 -1180
rect 3455 -1210 3470 -1180
rect 3410 -1250 3470 -1210
rect 3410 -1280 3425 -1250
rect 3455 -1280 3470 -1250
rect 3410 -1315 3470 -1280
rect 3410 -1345 3425 -1315
rect 3455 -1345 3470 -1315
rect 3410 -1360 3470 -1345
rect 3760 225 3820 240
rect 3760 195 3775 225
rect 3805 195 3820 225
rect 3760 160 3820 195
rect 3760 130 3775 160
rect 3805 130 3820 160
rect 3760 90 3820 130
rect 3760 60 3775 90
rect 3805 60 3820 90
rect 3760 20 3820 60
rect 3760 -10 3775 20
rect 3805 -10 3820 20
rect 3760 -50 3820 -10
rect 3760 -80 3775 -50
rect 3805 -80 3820 -50
rect 3760 -115 3820 -80
rect 3760 -145 3775 -115
rect 3805 -145 3820 -115
rect 3760 -175 3820 -145
rect 3760 -205 3775 -175
rect 3805 -205 3820 -175
rect 3760 -240 3820 -205
rect 3760 -270 3775 -240
rect 3805 -270 3820 -240
rect 3760 -310 3820 -270
rect 3760 -340 3775 -310
rect 3805 -340 3820 -310
rect 3760 -380 3820 -340
rect 3760 -410 3775 -380
rect 3805 -410 3820 -380
rect 3760 -450 3820 -410
rect 3760 -480 3775 -450
rect 3805 -480 3820 -450
rect 3760 -515 3820 -480
rect 3760 -545 3775 -515
rect 3805 -545 3820 -515
rect 3760 -575 3820 -545
rect 3760 -605 3775 -575
rect 3805 -605 3820 -575
rect 3760 -640 3820 -605
rect 3760 -670 3775 -640
rect 3805 -670 3820 -640
rect 3760 -710 3820 -670
rect 3760 -740 3775 -710
rect 3805 -740 3820 -710
rect 3760 -780 3820 -740
rect 3760 -810 3775 -780
rect 3805 -810 3820 -780
rect 3760 -850 3820 -810
rect 3760 -880 3775 -850
rect 3805 -880 3820 -850
rect 3760 -915 3820 -880
rect 3760 -945 3775 -915
rect 3805 -945 3820 -915
rect 3760 -975 3820 -945
rect 3760 -1005 3775 -975
rect 3805 -1005 3820 -975
rect 3760 -1040 3820 -1005
rect 3760 -1070 3775 -1040
rect 3805 -1070 3820 -1040
rect 3760 -1110 3820 -1070
rect 3760 -1140 3775 -1110
rect 3805 -1140 3820 -1110
rect 3760 -1180 3820 -1140
rect 3760 -1210 3775 -1180
rect 3805 -1210 3820 -1180
rect 3760 -1250 3820 -1210
rect 3760 -1280 3775 -1250
rect 3805 -1280 3820 -1250
rect 3760 -1315 3820 -1280
rect 3760 -1345 3775 -1315
rect 3805 -1345 3820 -1315
rect 3760 -1360 3820 -1345
rect 4110 225 4170 240
rect 4110 195 4125 225
rect 4155 195 4170 225
rect 4110 160 4170 195
rect 4110 130 4125 160
rect 4155 130 4170 160
rect 4110 90 4170 130
rect 4110 60 4125 90
rect 4155 60 4170 90
rect 4110 20 4170 60
rect 4110 -10 4125 20
rect 4155 -10 4170 20
rect 4110 -50 4170 -10
rect 4110 -80 4125 -50
rect 4155 -80 4170 -50
rect 4110 -115 4170 -80
rect 4110 -145 4125 -115
rect 4155 -145 4170 -115
rect 4110 -175 4170 -145
rect 4110 -205 4125 -175
rect 4155 -205 4170 -175
rect 4110 -240 4170 -205
rect 4110 -270 4125 -240
rect 4155 -270 4170 -240
rect 4110 -310 4170 -270
rect 4110 -340 4125 -310
rect 4155 -340 4170 -310
rect 4110 -380 4170 -340
rect 4110 -410 4125 -380
rect 4155 -410 4170 -380
rect 4110 -450 4170 -410
rect 4110 -480 4125 -450
rect 4155 -480 4170 -450
rect 4110 -515 4170 -480
rect 4110 -545 4125 -515
rect 4155 -545 4170 -515
rect 4110 -575 4170 -545
rect 4110 -605 4125 -575
rect 4155 -605 4170 -575
rect 4110 -640 4170 -605
rect 4110 -670 4125 -640
rect 4155 -670 4170 -640
rect 4110 -710 4170 -670
rect 4110 -740 4125 -710
rect 4155 -740 4170 -710
rect 4110 -780 4170 -740
rect 4110 -810 4125 -780
rect 4155 -810 4170 -780
rect 4110 -850 4170 -810
rect 4110 -880 4125 -850
rect 4155 -880 4170 -850
rect 4110 -915 4170 -880
rect 4110 -945 4125 -915
rect 4155 -945 4170 -915
rect 4110 -975 4170 -945
rect 4110 -1005 4125 -975
rect 4155 -1005 4170 -975
rect 4110 -1040 4170 -1005
rect 4110 -1070 4125 -1040
rect 4155 -1070 4170 -1040
rect 4110 -1110 4170 -1070
rect 4110 -1140 4125 -1110
rect 4155 -1140 4170 -1110
rect 4110 -1180 4170 -1140
rect 4110 -1210 4125 -1180
rect 4155 -1210 4170 -1180
rect 4110 -1250 4170 -1210
rect 4110 -1280 4125 -1250
rect 4155 -1280 4170 -1250
rect 4110 -1315 4170 -1280
rect 4110 -1345 4125 -1315
rect 4155 -1345 4170 -1315
rect 4110 -1360 4170 -1345
rect 4460 225 4520 240
rect 4460 195 4475 225
rect 4505 195 4520 225
rect 4460 160 4520 195
rect 4460 130 4475 160
rect 4505 130 4520 160
rect 4460 90 4520 130
rect 4460 60 4475 90
rect 4505 60 4520 90
rect 4460 20 4520 60
rect 4460 -10 4475 20
rect 4505 -10 4520 20
rect 4460 -50 4520 -10
rect 4460 -80 4475 -50
rect 4505 -80 4520 -50
rect 4460 -115 4520 -80
rect 4460 -145 4475 -115
rect 4505 -145 4520 -115
rect 4460 -175 4520 -145
rect 4460 -205 4475 -175
rect 4505 -205 4520 -175
rect 4460 -240 4520 -205
rect 4460 -270 4475 -240
rect 4505 -270 4520 -240
rect 4460 -310 4520 -270
rect 4460 -340 4475 -310
rect 4505 -340 4520 -310
rect 4460 -380 4520 -340
rect 4460 -410 4475 -380
rect 4505 -410 4520 -380
rect 4460 -450 4520 -410
rect 4460 -480 4475 -450
rect 4505 -480 4520 -450
rect 4460 -515 4520 -480
rect 4460 -545 4475 -515
rect 4505 -545 4520 -515
rect 4460 -575 4520 -545
rect 4460 -605 4475 -575
rect 4505 -605 4520 -575
rect 4460 -640 4520 -605
rect 4460 -670 4475 -640
rect 4505 -670 4520 -640
rect 4460 -710 4520 -670
rect 4460 -740 4475 -710
rect 4505 -740 4520 -710
rect 4460 -780 4520 -740
rect 4460 -810 4475 -780
rect 4505 -810 4520 -780
rect 4460 -850 4520 -810
rect 4460 -880 4475 -850
rect 4505 -880 4520 -850
rect 4460 -915 4520 -880
rect 4460 -945 4475 -915
rect 4505 -945 4520 -915
rect 4460 -975 4520 -945
rect 4460 -1005 4475 -975
rect 4505 -1005 4520 -975
rect 4460 -1040 4520 -1005
rect 4460 -1070 4475 -1040
rect 4505 -1070 4520 -1040
rect 4460 -1110 4520 -1070
rect 4460 -1140 4475 -1110
rect 4505 -1140 4520 -1110
rect 4460 -1180 4520 -1140
rect 4460 -1210 4475 -1180
rect 4505 -1210 4520 -1180
rect 4460 -1250 4520 -1210
rect 4460 -1280 4475 -1250
rect 4505 -1280 4520 -1250
rect 4460 -1315 4520 -1280
rect 4460 -1345 4475 -1315
rect 4505 -1345 4520 -1315
rect 4460 -1360 4520 -1345
rect 4810 225 4870 240
rect 4810 195 4825 225
rect 4855 195 4870 225
rect 4810 160 4870 195
rect 4810 130 4825 160
rect 4855 130 4870 160
rect 4810 90 4870 130
rect 4810 60 4825 90
rect 4855 60 4870 90
rect 4810 20 4870 60
rect 4810 -10 4825 20
rect 4855 -10 4870 20
rect 4810 -50 4870 -10
rect 4810 -80 4825 -50
rect 4855 -80 4870 -50
rect 4810 -115 4870 -80
rect 4810 -145 4825 -115
rect 4855 -145 4870 -115
rect 4810 -175 4870 -145
rect 4810 -205 4825 -175
rect 4855 -205 4870 -175
rect 4810 -240 4870 -205
rect 4810 -270 4825 -240
rect 4855 -270 4870 -240
rect 4810 -310 4870 -270
rect 4810 -340 4825 -310
rect 4855 -340 4870 -310
rect 4810 -380 4870 -340
rect 4810 -410 4825 -380
rect 4855 -410 4870 -380
rect 4810 -450 4870 -410
rect 4810 -480 4825 -450
rect 4855 -480 4870 -450
rect 4810 -515 4870 -480
rect 4810 -545 4825 -515
rect 4855 -545 4870 -515
rect 4810 -575 4870 -545
rect 4810 -605 4825 -575
rect 4855 -605 4870 -575
rect 4810 -640 4870 -605
rect 4810 -670 4825 -640
rect 4855 -670 4870 -640
rect 4810 -710 4870 -670
rect 4810 -740 4825 -710
rect 4855 -740 4870 -710
rect 4810 -780 4870 -740
rect 4810 -810 4825 -780
rect 4855 -810 4870 -780
rect 4810 -850 4870 -810
rect 4810 -880 4825 -850
rect 4855 -880 4870 -850
rect 4810 -915 4870 -880
rect 4810 -945 4825 -915
rect 4855 -945 4870 -915
rect 4810 -975 4870 -945
rect 4810 -1005 4825 -975
rect 4855 -1005 4870 -975
rect 4810 -1040 4870 -1005
rect 4810 -1070 4825 -1040
rect 4855 -1070 4870 -1040
rect 4810 -1110 4870 -1070
rect 4810 -1140 4825 -1110
rect 4855 -1140 4870 -1110
rect 4810 -1180 4870 -1140
rect 4810 -1210 4825 -1180
rect 4855 -1210 4870 -1180
rect 4810 -1250 4870 -1210
rect 4810 -1280 4825 -1250
rect 4855 -1280 4870 -1250
rect 4810 -1315 4870 -1280
rect 4810 -1345 4825 -1315
rect 4855 -1345 4870 -1315
rect 4810 -1360 4870 -1345
rect 5160 225 5220 240
rect 5160 195 5175 225
rect 5205 195 5220 225
rect 5160 160 5220 195
rect 5160 130 5175 160
rect 5205 130 5220 160
rect 5160 90 5220 130
rect 5160 60 5175 90
rect 5205 60 5220 90
rect 5160 20 5220 60
rect 5160 -10 5175 20
rect 5205 -10 5220 20
rect 5160 -50 5220 -10
rect 5160 -80 5175 -50
rect 5205 -80 5220 -50
rect 5160 -115 5220 -80
rect 5160 -145 5175 -115
rect 5205 -145 5220 -115
rect 5160 -175 5220 -145
rect 5160 -205 5175 -175
rect 5205 -205 5220 -175
rect 5160 -240 5220 -205
rect 5160 -270 5175 -240
rect 5205 -270 5220 -240
rect 5160 -310 5220 -270
rect 5160 -340 5175 -310
rect 5205 -340 5220 -310
rect 5160 -380 5220 -340
rect 5160 -410 5175 -380
rect 5205 -410 5220 -380
rect 5160 -450 5220 -410
rect 5160 -480 5175 -450
rect 5205 -480 5220 -450
rect 5160 -515 5220 -480
rect 5160 -545 5175 -515
rect 5205 -545 5220 -515
rect 5160 -575 5220 -545
rect 5160 -605 5175 -575
rect 5205 -605 5220 -575
rect 5160 -640 5220 -605
rect 5160 -670 5175 -640
rect 5205 -670 5220 -640
rect 5160 -710 5220 -670
rect 5160 -740 5175 -710
rect 5205 -740 5220 -710
rect 5160 -780 5220 -740
rect 5160 -810 5175 -780
rect 5205 -810 5220 -780
rect 5160 -850 5220 -810
rect 5160 -880 5175 -850
rect 5205 -880 5220 -850
rect 5160 -915 5220 -880
rect 5160 -945 5175 -915
rect 5205 -945 5220 -915
rect 5160 -975 5220 -945
rect 5160 -1005 5175 -975
rect 5205 -1005 5220 -975
rect 5160 -1040 5220 -1005
rect 5160 -1070 5175 -1040
rect 5205 -1070 5220 -1040
rect 5160 -1110 5220 -1070
rect 5160 -1140 5175 -1110
rect 5205 -1140 5220 -1110
rect 5160 -1180 5220 -1140
rect 5160 -1210 5175 -1180
rect 5205 -1210 5220 -1180
rect 5160 -1250 5220 -1210
rect 5160 -1280 5175 -1250
rect 5205 -1280 5220 -1250
rect 5160 -1315 5220 -1280
rect 5160 -1345 5175 -1315
rect 5205 -1345 5220 -1315
rect 5160 -1360 5220 -1345
rect 5510 225 5570 240
rect 5510 195 5525 225
rect 5555 195 5570 225
rect 5510 160 5570 195
rect 5510 130 5525 160
rect 5555 130 5570 160
rect 5510 90 5570 130
rect 5510 60 5525 90
rect 5555 60 5570 90
rect 5510 20 5570 60
rect 5510 -10 5525 20
rect 5555 -10 5570 20
rect 5510 -50 5570 -10
rect 5510 -80 5525 -50
rect 5555 -80 5570 -50
rect 5510 -115 5570 -80
rect 5510 -145 5525 -115
rect 5555 -145 5570 -115
rect 5510 -175 5570 -145
rect 5510 -205 5525 -175
rect 5555 -205 5570 -175
rect 5510 -240 5570 -205
rect 5510 -270 5525 -240
rect 5555 -270 5570 -240
rect 5510 -310 5570 -270
rect 5510 -340 5525 -310
rect 5555 -340 5570 -310
rect 5510 -380 5570 -340
rect 5510 -410 5525 -380
rect 5555 -410 5570 -380
rect 5510 -450 5570 -410
rect 5510 -480 5525 -450
rect 5555 -480 5570 -450
rect 5510 -515 5570 -480
rect 5510 -545 5525 -515
rect 5555 -545 5570 -515
rect 5510 -575 5570 -545
rect 5510 -605 5525 -575
rect 5555 -605 5570 -575
rect 5510 -640 5570 -605
rect 5510 -670 5525 -640
rect 5555 -670 5570 -640
rect 5510 -710 5570 -670
rect 5510 -740 5525 -710
rect 5555 -740 5570 -710
rect 5510 -780 5570 -740
rect 5510 -810 5525 -780
rect 5555 -810 5570 -780
rect 5510 -850 5570 -810
rect 5510 -880 5525 -850
rect 5555 -880 5570 -850
rect 5510 -915 5570 -880
rect 5510 -945 5525 -915
rect 5555 -945 5570 -915
rect 5510 -975 5570 -945
rect 5510 -1005 5525 -975
rect 5555 -1005 5570 -975
rect 5510 -1040 5570 -1005
rect 5510 -1070 5525 -1040
rect 5555 -1070 5570 -1040
rect 5510 -1110 5570 -1070
rect 5510 -1140 5525 -1110
rect 5555 -1140 5570 -1110
rect 5510 -1180 5570 -1140
rect 5510 -1210 5525 -1180
rect 5555 -1210 5570 -1180
rect 5510 -1250 5570 -1210
rect 5510 -1280 5525 -1250
rect 5555 -1280 5570 -1250
rect 5510 -1315 5570 -1280
rect 5510 -1345 5525 -1315
rect 5555 -1345 5570 -1315
rect 5510 -1360 5570 -1345
rect 5860 225 5920 240
rect 5860 195 5875 225
rect 5905 195 5920 225
rect 5860 160 5920 195
rect 5860 130 5875 160
rect 5905 130 5920 160
rect 5860 90 5920 130
rect 5860 60 5875 90
rect 5905 60 5920 90
rect 5860 20 5920 60
rect 5860 -10 5875 20
rect 5905 -10 5920 20
rect 5860 -50 5920 -10
rect 5860 -80 5875 -50
rect 5905 -80 5920 -50
rect 5860 -115 5920 -80
rect 5860 -145 5875 -115
rect 5905 -145 5920 -115
rect 5860 -175 5920 -145
rect 5860 -205 5875 -175
rect 5905 -205 5920 -175
rect 5860 -240 5920 -205
rect 5860 -270 5875 -240
rect 5905 -270 5920 -240
rect 5860 -310 5920 -270
rect 5860 -340 5875 -310
rect 5905 -340 5920 -310
rect 5860 -380 5920 -340
rect 5860 -410 5875 -380
rect 5905 -410 5920 -380
rect 5860 -450 5920 -410
rect 5860 -480 5875 -450
rect 5905 -480 5920 -450
rect 5860 -515 5920 -480
rect 5860 -545 5875 -515
rect 5905 -545 5920 -515
rect 5860 -575 5920 -545
rect 5860 -605 5875 -575
rect 5905 -605 5920 -575
rect 5860 -640 5920 -605
rect 5860 -670 5875 -640
rect 5905 -670 5920 -640
rect 5860 -710 5920 -670
rect 5860 -740 5875 -710
rect 5905 -740 5920 -710
rect 5860 -780 5920 -740
rect 5860 -810 5875 -780
rect 5905 -810 5920 -780
rect 5860 -850 5920 -810
rect 5860 -880 5875 -850
rect 5905 -880 5920 -850
rect 5860 -915 5920 -880
rect 5860 -945 5875 -915
rect 5905 -945 5920 -915
rect 5860 -975 5920 -945
rect 5860 -1005 5875 -975
rect 5905 -1005 5920 -975
rect 5860 -1040 5920 -1005
rect 5860 -1070 5875 -1040
rect 5905 -1070 5920 -1040
rect 5860 -1110 5920 -1070
rect 5860 -1140 5875 -1110
rect 5905 -1140 5920 -1110
rect 5860 -1180 5920 -1140
rect 5860 -1210 5875 -1180
rect 5905 -1210 5920 -1180
rect 5860 -1250 5920 -1210
rect 5860 -1280 5875 -1250
rect 5905 -1280 5920 -1250
rect 5860 -1315 5920 -1280
rect 5860 -1345 5875 -1315
rect 5905 -1345 5920 -1315
rect 5860 -1360 5920 -1345
rect 6210 225 6270 240
rect 6210 195 6225 225
rect 6255 195 6270 225
rect 6210 160 6270 195
rect 6210 130 6225 160
rect 6255 130 6270 160
rect 6210 90 6270 130
rect 6210 60 6225 90
rect 6255 60 6270 90
rect 6210 20 6270 60
rect 6210 -10 6225 20
rect 6255 -10 6270 20
rect 6210 -50 6270 -10
rect 6210 -80 6225 -50
rect 6255 -80 6270 -50
rect 6210 -115 6270 -80
rect 6210 -145 6225 -115
rect 6255 -145 6270 -115
rect 6210 -175 6270 -145
rect 6210 -205 6225 -175
rect 6255 -205 6270 -175
rect 6210 -240 6270 -205
rect 6210 -270 6225 -240
rect 6255 -270 6270 -240
rect 6210 -310 6270 -270
rect 6210 -340 6225 -310
rect 6255 -340 6270 -310
rect 6210 -380 6270 -340
rect 6210 -410 6225 -380
rect 6255 -410 6270 -380
rect 6210 -450 6270 -410
rect 6210 -480 6225 -450
rect 6255 -480 6270 -450
rect 6210 -515 6270 -480
rect 6210 -545 6225 -515
rect 6255 -545 6270 -515
rect 6210 -575 6270 -545
rect 6210 -605 6225 -575
rect 6255 -605 6270 -575
rect 6210 -640 6270 -605
rect 6210 -670 6225 -640
rect 6255 -670 6270 -640
rect 6210 -710 6270 -670
rect 6210 -740 6225 -710
rect 6255 -740 6270 -710
rect 6210 -780 6270 -740
rect 6210 -810 6225 -780
rect 6255 -810 6270 -780
rect 6210 -850 6270 -810
rect 6210 -880 6225 -850
rect 6255 -880 6270 -850
rect 6210 -915 6270 -880
rect 6210 -945 6225 -915
rect 6255 -945 6270 -915
rect 6210 -975 6270 -945
rect 6210 -1005 6225 -975
rect 6255 -1005 6270 -975
rect 6210 -1040 6270 -1005
rect 6210 -1070 6225 -1040
rect 6255 -1070 6270 -1040
rect 6210 -1110 6270 -1070
rect 6210 -1140 6225 -1110
rect 6255 -1140 6270 -1110
rect 6210 -1180 6270 -1140
rect 6210 -1210 6225 -1180
rect 6255 -1210 6270 -1180
rect 6210 -1250 6270 -1210
rect 6210 -1280 6225 -1250
rect 6255 -1280 6270 -1250
rect 6210 -1315 6270 -1280
rect 6210 -1345 6225 -1315
rect 6255 -1345 6270 -1315
rect 6210 -1360 6270 -1345
rect 6560 225 6620 240
rect 6560 195 6575 225
rect 6605 195 6620 225
rect 6560 160 6620 195
rect 6560 130 6575 160
rect 6605 130 6620 160
rect 6560 90 6620 130
rect 6560 60 6575 90
rect 6605 60 6620 90
rect 6560 20 6620 60
rect 6560 -10 6575 20
rect 6605 -10 6620 20
rect 6560 -50 6620 -10
rect 6560 -80 6575 -50
rect 6605 -80 6620 -50
rect 6560 -115 6620 -80
rect 6560 -145 6575 -115
rect 6605 -145 6620 -115
rect 6560 -175 6620 -145
rect 6560 -205 6575 -175
rect 6605 -205 6620 -175
rect 6560 -240 6620 -205
rect 6560 -270 6575 -240
rect 6605 -270 6620 -240
rect 6560 -310 6620 -270
rect 6560 -340 6575 -310
rect 6605 -340 6620 -310
rect 6560 -380 6620 -340
rect 6560 -410 6575 -380
rect 6605 -410 6620 -380
rect 6560 -450 6620 -410
rect 6560 -480 6575 -450
rect 6605 -480 6620 -450
rect 6560 -515 6620 -480
rect 6560 -545 6575 -515
rect 6605 -545 6620 -515
rect 6560 -575 6620 -545
rect 6560 -605 6575 -575
rect 6605 -605 6620 -575
rect 6560 -640 6620 -605
rect 6560 -670 6575 -640
rect 6605 -670 6620 -640
rect 6560 -710 6620 -670
rect 6560 -740 6575 -710
rect 6605 -740 6620 -710
rect 6560 -780 6620 -740
rect 6560 -810 6575 -780
rect 6605 -810 6620 -780
rect 6560 -850 6620 -810
rect 6560 -880 6575 -850
rect 6605 -880 6620 -850
rect 6560 -915 6620 -880
rect 6560 -945 6575 -915
rect 6605 -945 6620 -915
rect 6560 -975 6620 -945
rect 6560 -1005 6575 -975
rect 6605 -1005 6620 -975
rect 6560 -1040 6620 -1005
rect 6560 -1070 6575 -1040
rect 6605 -1070 6620 -1040
rect 6560 -1110 6620 -1070
rect 6560 -1140 6575 -1110
rect 6605 -1140 6620 -1110
rect 6560 -1180 6620 -1140
rect 6560 -1210 6575 -1180
rect 6605 -1210 6620 -1180
rect 6560 -1250 6620 -1210
rect 6560 -1280 6575 -1250
rect 6605 -1280 6620 -1250
rect 6560 -1315 6620 -1280
rect 6560 -1345 6575 -1315
rect 6605 -1345 6620 -1315
rect 6560 -1360 6620 -1345
rect 6910 225 6970 240
rect 6910 195 6925 225
rect 6955 195 6970 225
rect 6910 160 6970 195
rect 6910 130 6925 160
rect 6955 130 6970 160
rect 6910 90 6970 130
rect 6910 60 6925 90
rect 6955 60 6970 90
rect 6910 20 6970 60
rect 6910 -10 6925 20
rect 6955 -10 6970 20
rect 6910 -50 6970 -10
rect 6910 -80 6925 -50
rect 6955 -80 6970 -50
rect 6910 -115 6970 -80
rect 6910 -145 6925 -115
rect 6955 -145 6970 -115
rect 6910 -175 6970 -145
rect 6910 -205 6925 -175
rect 6955 -205 6970 -175
rect 6910 -240 6970 -205
rect 6910 -270 6925 -240
rect 6955 -270 6970 -240
rect 6910 -310 6970 -270
rect 6910 -340 6925 -310
rect 6955 -340 6970 -310
rect 6910 -380 6970 -340
rect 6910 -410 6925 -380
rect 6955 -410 6970 -380
rect 6910 -450 6970 -410
rect 6910 -480 6925 -450
rect 6955 -480 6970 -450
rect 6910 -515 6970 -480
rect 6910 -545 6925 -515
rect 6955 -545 6970 -515
rect 6910 -575 6970 -545
rect 6910 -605 6925 -575
rect 6955 -605 6970 -575
rect 6910 -640 6970 -605
rect 6910 -670 6925 -640
rect 6955 -670 6970 -640
rect 6910 -710 6970 -670
rect 6910 -740 6925 -710
rect 6955 -740 6970 -710
rect 6910 -780 6970 -740
rect 6910 -810 6925 -780
rect 6955 -810 6970 -780
rect 6910 -850 6970 -810
rect 6910 -880 6925 -850
rect 6955 -880 6970 -850
rect 6910 -915 6970 -880
rect 6910 -945 6925 -915
rect 6955 -945 6970 -915
rect 6910 -975 6970 -945
rect 6910 -1005 6925 -975
rect 6955 -1005 6970 -975
rect 6910 -1040 6970 -1005
rect 6910 -1070 6925 -1040
rect 6955 -1070 6970 -1040
rect 6910 -1110 6970 -1070
rect 6910 -1140 6925 -1110
rect 6955 -1140 6970 -1110
rect 6910 -1180 6970 -1140
rect 6910 -1210 6925 -1180
rect 6955 -1210 6970 -1180
rect 6910 -1250 6970 -1210
rect 6910 -1280 6925 -1250
rect 6955 -1280 6970 -1250
rect 6910 -1315 6970 -1280
rect 6910 -1345 6925 -1315
rect 6955 -1345 6970 -1315
rect 6910 -1360 6970 -1345
rect 7260 225 7320 240
rect 7260 195 7275 225
rect 7305 195 7320 225
rect 7260 160 7320 195
rect 7260 130 7275 160
rect 7305 130 7320 160
rect 7260 90 7320 130
rect 7260 60 7275 90
rect 7305 60 7320 90
rect 7260 20 7320 60
rect 7260 -10 7275 20
rect 7305 -10 7320 20
rect 7260 -50 7320 -10
rect 7260 -80 7275 -50
rect 7305 -80 7320 -50
rect 7260 -115 7320 -80
rect 7260 -145 7275 -115
rect 7305 -145 7320 -115
rect 7260 -175 7320 -145
rect 7260 -205 7275 -175
rect 7305 -205 7320 -175
rect 7260 -240 7320 -205
rect 7260 -270 7275 -240
rect 7305 -270 7320 -240
rect 7260 -310 7320 -270
rect 7260 -340 7275 -310
rect 7305 -340 7320 -310
rect 7260 -380 7320 -340
rect 7260 -410 7275 -380
rect 7305 -410 7320 -380
rect 7260 -450 7320 -410
rect 7260 -480 7275 -450
rect 7305 -480 7320 -450
rect 7260 -515 7320 -480
rect 7260 -545 7275 -515
rect 7305 -545 7320 -515
rect 7260 -575 7320 -545
rect 7260 -605 7275 -575
rect 7305 -605 7320 -575
rect 7260 -640 7320 -605
rect 7260 -670 7275 -640
rect 7305 -670 7320 -640
rect 7260 -710 7320 -670
rect 7260 -740 7275 -710
rect 7305 -740 7320 -710
rect 7260 -780 7320 -740
rect 7260 -810 7275 -780
rect 7305 -810 7320 -780
rect 7260 -850 7320 -810
rect 7260 -880 7275 -850
rect 7305 -880 7320 -850
rect 7260 -915 7320 -880
rect 7260 -945 7275 -915
rect 7305 -945 7320 -915
rect 7260 -975 7320 -945
rect 7260 -1005 7275 -975
rect 7305 -1005 7320 -975
rect 7260 -1040 7320 -1005
rect 7260 -1070 7275 -1040
rect 7305 -1070 7320 -1040
rect 7260 -1110 7320 -1070
rect 7260 -1140 7275 -1110
rect 7305 -1140 7320 -1110
rect 7260 -1180 7320 -1140
rect 7260 -1210 7275 -1180
rect 7305 -1210 7320 -1180
rect 7260 -1250 7320 -1210
rect 7260 -1280 7275 -1250
rect 7305 -1280 7320 -1250
rect 7260 -1315 7320 -1280
rect 7260 -1345 7275 -1315
rect 7305 -1345 7320 -1315
rect 7260 -1360 7320 -1345
rect 7610 225 7670 240
rect 7610 195 7625 225
rect 7655 195 7670 225
rect 7610 160 7670 195
rect 7610 130 7625 160
rect 7655 130 7670 160
rect 7610 90 7670 130
rect 7610 60 7625 90
rect 7655 60 7670 90
rect 7610 20 7670 60
rect 7610 -10 7625 20
rect 7655 -10 7670 20
rect 7610 -50 7670 -10
rect 7610 -80 7625 -50
rect 7655 -80 7670 -50
rect 7610 -115 7670 -80
rect 7610 -145 7625 -115
rect 7655 -145 7670 -115
rect 7610 -175 7670 -145
rect 7610 -205 7625 -175
rect 7655 -205 7670 -175
rect 7610 -240 7670 -205
rect 7610 -270 7625 -240
rect 7655 -270 7670 -240
rect 7610 -310 7670 -270
rect 7610 -340 7625 -310
rect 7655 -340 7670 -310
rect 7610 -380 7670 -340
rect 7610 -410 7625 -380
rect 7655 -410 7670 -380
rect 7610 -450 7670 -410
rect 7610 -480 7625 -450
rect 7655 -480 7670 -450
rect 7610 -515 7670 -480
rect 7610 -545 7625 -515
rect 7655 -545 7670 -515
rect 7610 -575 7670 -545
rect 7610 -605 7625 -575
rect 7655 -605 7670 -575
rect 7610 -640 7670 -605
rect 7610 -670 7625 -640
rect 7655 -670 7670 -640
rect 7610 -710 7670 -670
rect 7610 -740 7625 -710
rect 7655 -740 7670 -710
rect 7610 -780 7670 -740
rect 7610 -810 7625 -780
rect 7655 -810 7670 -780
rect 7610 -850 7670 -810
rect 7610 -880 7625 -850
rect 7655 -880 7670 -850
rect 7610 -915 7670 -880
rect 7610 -945 7625 -915
rect 7655 -945 7670 -915
rect 7610 -975 7670 -945
rect 7610 -1005 7625 -975
rect 7655 -1005 7670 -975
rect 7610 -1040 7670 -1005
rect 7610 -1070 7625 -1040
rect 7655 -1070 7670 -1040
rect 7610 -1110 7670 -1070
rect 7610 -1140 7625 -1110
rect 7655 -1140 7670 -1110
rect 7610 -1180 7670 -1140
rect 7610 -1210 7625 -1180
rect 7655 -1210 7670 -1180
rect 7610 -1250 7670 -1210
rect 7610 -1280 7625 -1250
rect 7655 -1280 7670 -1250
rect 7610 -1315 7670 -1280
rect 7610 -1345 7625 -1315
rect 7655 -1345 7670 -1315
rect 7610 -1360 7670 -1345
rect 7960 225 8020 240
rect 7960 195 7975 225
rect 8005 195 8020 225
rect 7960 160 8020 195
rect 7960 130 7975 160
rect 8005 130 8020 160
rect 7960 90 8020 130
rect 7960 60 7975 90
rect 8005 60 8020 90
rect 7960 20 8020 60
rect 7960 -10 7975 20
rect 8005 -10 8020 20
rect 7960 -50 8020 -10
rect 7960 -80 7975 -50
rect 8005 -80 8020 -50
rect 7960 -115 8020 -80
rect 7960 -145 7975 -115
rect 8005 -145 8020 -115
rect 7960 -175 8020 -145
rect 7960 -205 7975 -175
rect 8005 -205 8020 -175
rect 7960 -240 8020 -205
rect 7960 -270 7975 -240
rect 8005 -270 8020 -240
rect 7960 -310 8020 -270
rect 7960 -340 7975 -310
rect 8005 -340 8020 -310
rect 7960 -380 8020 -340
rect 7960 -410 7975 -380
rect 8005 -410 8020 -380
rect 7960 -450 8020 -410
rect 7960 -480 7975 -450
rect 8005 -480 8020 -450
rect 7960 -515 8020 -480
rect 7960 -545 7975 -515
rect 8005 -545 8020 -515
rect 7960 -575 8020 -545
rect 7960 -605 7975 -575
rect 8005 -605 8020 -575
rect 7960 -640 8020 -605
rect 7960 -670 7975 -640
rect 8005 -670 8020 -640
rect 7960 -710 8020 -670
rect 7960 -740 7975 -710
rect 8005 -740 8020 -710
rect 7960 -780 8020 -740
rect 7960 -810 7975 -780
rect 8005 -810 8020 -780
rect 7960 -850 8020 -810
rect 7960 -880 7975 -850
rect 8005 -880 8020 -850
rect 7960 -915 8020 -880
rect 7960 -945 7975 -915
rect 8005 -945 8020 -915
rect 7960 -975 8020 -945
rect 7960 -1005 7975 -975
rect 8005 -1005 8020 -975
rect 7960 -1040 8020 -1005
rect 7960 -1070 7975 -1040
rect 8005 -1070 8020 -1040
rect 7960 -1110 8020 -1070
rect 7960 -1140 7975 -1110
rect 8005 -1140 8020 -1110
rect 7960 -1180 8020 -1140
rect 7960 -1210 7975 -1180
rect 8005 -1210 8020 -1180
rect 7960 -1250 8020 -1210
rect 7960 -1280 7975 -1250
rect 8005 -1280 8020 -1250
rect 7960 -1315 8020 -1280
rect 7960 -1345 7975 -1315
rect 8005 -1345 8020 -1315
rect 7960 -1360 8020 -1345
rect 8310 225 8370 240
rect 8310 195 8325 225
rect 8355 195 8370 225
rect 8310 160 8370 195
rect 8310 130 8325 160
rect 8355 130 8370 160
rect 8310 90 8370 130
rect 8310 60 8325 90
rect 8355 60 8370 90
rect 8310 20 8370 60
rect 8310 -10 8325 20
rect 8355 -10 8370 20
rect 8310 -50 8370 -10
rect 8310 -80 8325 -50
rect 8355 -80 8370 -50
rect 8310 -115 8370 -80
rect 8310 -145 8325 -115
rect 8355 -145 8370 -115
rect 8310 -175 8370 -145
rect 8310 -205 8325 -175
rect 8355 -205 8370 -175
rect 8310 -240 8370 -205
rect 8310 -270 8325 -240
rect 8355 -270 8370 -240
rect 8310 -310 8370 -270
rect 8310 -340 8325 -310
rect 8355 -340 8370 -310
rect 8310 -380 8370 -340
rect 8310 -410 8325 -380
rect 8355 -410 8370 -380
rect 8310 -450 8370 -410
rect 8310 -480 8325 -450
rect 8355 -480 8370 -450
rect 8310 -515 8370 -480
rect 8310 -545 8325 -515
rect 8355 -545 8370 -515
rect 8310 -575 8370 -545
rect 8310 -605 8325 -575
rect 8355 -605 8370 -575
rect 8310 -640 8370 -605
rect 8310 -670 8325 -640
rect 8355 -670 8370 -640
rect 8310 -710 8370 -670
rect 8310 -740 8325 -710
rect 8355 -740 8370 -710
rect 8310 -780 8370 -740
rect 8310 -810 8325 -780
rect 8355 -810 8370 -780
rect 8310 -850 8370 -810
rect 8310 -880 8325 -850
rect 8355 -880 8370 -850
rect 8310 -915 8370 -880
rect 8310 -945 8325 -915
rect 8355 -945 8370 -915
rect 8310 -975 8370 -945
rect 8310 -1005 8325 -975
rect 8355 -1005 8370 -975
rect 8310 -1040 8370 -1005
rect 8310 -1070 8325 -1040
rect 8355 -1070 8370 -1040
rect 8310 -1110 8370 -1070
rect 8310 -1140 8325 -1110
rect 8355 -1140 8370 -1110
rect 8310 -1180 8370 -1140
rect 8310 -1210 8325 -1180
rect 8355 -1210 8370 -1180
rect 8310 -1250 8370 -1210
rect 8310 -1280 8325 -1250
rect 8355 -1280 8370 -1250
rect 8310 -1315 8370 -1280
rect 8310 -1345 8325 -1315
rect 8355 -1345 8370 -1315
rect 8310 -1360 8370 -1345
rect 8660 225 8720 240
rect 8660 195 8675 225
rect 8705 195 8720 225
rect 8660 160 8720 195
rect 8660 130 8675 160
rect 8705 130 8720 160
rect 8660 90 8720 130
rect 8660 60 8675 90
rect 8705 60 8720 90
rect 8660 20 8720 60
rect 8660 -10 8675 20
rect 8705 -10 8720 20
rect 8660 -50 8720 -10
rect 8660 -80 8675 -50
rect 8705 -80 8720 -50
rect 8660 -115 8720 -80
rect 8660 -145 8675 -115
rect 8705 -145 8720 -115
rect 8660 -175 8720 -145
rect 8660 -205 8675 -175
rect 8705 -205 8720 -175
rect 8660 -240 8720 -205
rect 8660 -270 8675 -240
rect 8705 -270 8720 -240
rect 8660 -310 8720 -270
rect 8660 -340 8675 -310
rect 8705 -340 8720 -310
rect 8660 -380 8720 -340
rect 8660 -410 8675 -380
rect 8705 -410 8720 -380
rect 8660 -450 8720 -410
rect 8660 -480 8675 -450
rect 8705 -480 8720 -450
rect 8660 -515 8720 -480
rect 8660 -545 8675 -515
rect 8705 -545 8720 -515
rect 8660 -575 8720 -545
rect 8660 -605 8675 -575
rect 8705 -605 8720 -575
rect 8660 -640 8720 -605
rect 8660 -670 8675 -640
rect 8705 -670 8720 -640
rect 8660 -710 8720 -670
rect 8660 -740 8675 -710
rect 8705 -740 8720 -710
rect 8660 -780 8720 -740
rect 8660 -810 8675 -780
rect 8705 -810 8720 -780
rect 8660 -850 8720 -810
rect 8660 -880 8675 -850
rect 8705 -880 8720 -850
rect 8660 -915 8720 -880
rect 8660 -945 8675 -915
rect 8705 -945 8720 -915
rect 8660 -975 8720 -945
rect 8660 -1005 8675 -975
rect 8705 -1005 8720 -975
rect 8660 -1040 8720 -1005
rect 8660 -1070 8675 -1040
rect 8705 -1070 8720 -1040
rect 8660 -1110 8720 -1070
rect 8660 -1140 8675 -1110
rect 8705 -1140 8720 -1110
rect 8660 -1180 8720 -1140
rect 8660 -1210 8675 -1180
rect 8705 -1210 8720 -1180
rect 8660 -1250 8720 -1210
rect 8660 -1280 8675 -1250
rect 8705 -1280 8720 -1250
rect 8660 -1315 8720 -1280
rect 8660 -1345 8675 -1315
rect 8705 -1345 8720 -1315
rect 8660 -1360 8720 -1345
rect 9010 225 9070 240
rect 9010 195 9025 225
rect 9055 195 9070 225
rect 9010 160 9070 195
rect 9010 130 9025 160
rect 9055 130 9070 160
rect 9010 90 9070 130
rect 9010 60 9025 90
rect 9055 60 9070 90
rect 9010 20 9070 60
rect 9010 -10 9025 20
rect 9055 -10 9070 20
rect 9010 -50 9070 -10
rect 9010 -80 9025 -50
rect 9055 -80 9070 -50
rect 9010 -115 9070 -80
rect 9010 -145 9025 -115
rect 9055 -145 9070 -115
rect 9010 -175 9070 -145
rect 9010 -205 9025 -175
rect 9055 -205 9070 -175
rect 9010 -240 9070 -205
rect 9010 -270 9025 -240
rect 9055 -270 9070 -240
rect 9010 -310 9070 -270
rect 9010 -340 9025 -310
rect 9055 -340 9070 -310
rect 9010 -380 9070 -340
rect 9010 -410 9025 -380
rect 9055 -410 9070 -380
rect 9010 -450 9070 -410
rect 9010 -480 9025 -450
rect 9055 -480 9070 -450
rect 9010 -515 9070 -480
rect 9010 -545 9025 -515
rect 9055 -545 9070 -515
rect 9010 -575 9070 -545
rect 9010 -605 9025 -575
rect 9055 -605 9070 -575
rect 9010 -640 9070 -605
rect 9010 -670 9025 -640
rect 9055 -670 9070 -640
rect 9010 -710 9070 -670
rect 9010 -740 9025 -710
rect 9055 -740 9070 -710
rect 9010 -780 9070 -740
rect 9010 -810 9025 -780
rect 9055 -810 9070 -780
rect 9010 -850 9070 -810
rect 9010 -880 9025 -850
rect 9055 -880 9070 -850
rect 9010 -915 9070 -880
rect 9010 -945 9025 -915
rect 9055 -945 9070 -915
rect 9010 -975 9070 -945
rect 9010 -1005 9025 -975
rect 9055 -1005 9070 -975
rect 9010 -1040 9070 -1005
rect 9010 -1070 9025 -1040
rect 9055 -1070 9070 -1040
rect 9010 -1110 9070 -1070
rect 9010 -1140 9025 -1110
rect 9055 -1140 9070 -1110
rect 9010 -1180 9070 -1140
rect 9010 -1210 9025 -1180
rect 9055 -1210 9070 -1180
rect 9010 -1250 9070 -1210
rect 9010 -1280 9025 -1250
rect 9055 -1280 9070 -1250
rect 9010 -1315 9070 -1280
rect 9010 -1345 9025 -1315
rect 9055 -1345 9070 -1315
rect 9010 -1360 9070 -1345
<< via2 >>
rect 2115 19280 2145 19310
rect 2115 19215 2145 19245
rect 2115 19145 2145 19175
rect 2115 19075 2145 19105
rect 2115 19005 2145 19035
rect 2115 18940 2145 18970
rect 2115 18880 2145 18910
rect 2115 18815 2145 18845
rect 2115 18745 2145 18775
rect 2115 18675 2145 18705
rect 2115 18605 2145 18635
rect 2115 18540 2145 18570
rect 2115 18480 2145 18510
rect 2115 18415 2145 18445
rect 2115 18345 2145 18375
rect 2115 18275 2145 18305
rect 2115 18205 2145 18235
rect 2115 18140 2145 18170
rect 2115 18080 2145 18110
rect 2115 18015 2145 18045
rect 2115 17945 2145 17975
rect 2115 17875 2145 17905
rect 2115 17805 2145 17835
rect 2115 17740 2145 17770
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 1325 9605 1355 9635
rect 1325 9540 1355 9570
rect 1325 9470 1355 9500
rect 1325 9400 1355 9430
rect 1325 9330 1355 9360
rect 1325 9265 1355 9295
rect 1325 9205 1355 9235
rect 1325 9140 1355 9170
rect 1325 9070 1355 9100
rect 1325 9000 1355 9030
rect 1325 8930 1355 8960
rect 1325 8865 1355 8895
rect 1325 8805 1355 8835
rect 1325 8740 1355 8770
rect 1325 8670 1355 8700
rect 1325 8600 1355 8630
rect 1325 8530 1355 8560
rect 1325 8465 1355 8495
rect 1325 8405 1355 8435
rect 1325 8340 1355 8370
rect 1325 8270 1355 8300
rect 1325 8200 1355 8230
rect 1325 8130 1355 8160
rect 2250 9605 2280 9635
rect 2250 9540 2280 9570
rect 2250 9470 2280 9500
rect 2250 9400 2280 9430
rect 2250 9330 2280 9360
rect 2250 9265 2280 9295
rect 2250 9205 2280 9235
rect 2250 9140 2280 9170
rect 2250 9070 2280 9100
rect 2250 9000 2280 9030
rect 2250 8930 2280 8960
rect 2250 8865 2280 8895
rect 2250 8805 2280 8835
rect 2250 8740 2280 8770
rect 2250 8670 2280 8700
rect 2250 8600 2280 8630
rect 2250 8530 2280 8560
rect 2250 8465 2280 8495
rect 2250 8405 2280 8435
rect 2250 8340 2280 8370
rect 2250 8270 2280 8300
rect 2250 8200 2280 8230
rect 2250 8130 2280 8160
rect 3180 9605 3210 9635
rect 3180 9540 3210 9570
rect 3180 9470 3210 9500
rect 3180 9400 3210 9430
rect 3180 9330 3210 9360
rect 3180 9265 3210 9295
rect 3180 9205 3210 9235
rect 3180 9140 3210 9170
rect 3180 9070 3210 9100
rect 3180 9000 3210 9030
rect 3180 8930 3210 8960
rect 3180 8865 3210 8895
rect 3180 8805 3210 8835
rect 3180 8740 3210 8770
rect 3180 8670 3210 8700
rect 3180 8600 3210 8630
rect 3180 8530 3210 8560
rect 3180 8465 3210 8495
rect 3180 8405 3210 8435
rect 3180 8340 3210 8370
rect 3180 8270 3210 8300
rect 3180 8200 3210 8230
rect 3180 8130 3210 8160
rect 6705 9605 6735 9635
rect 6705 9540 6735 9570
rect 6705 9470 6735 9500
rect 6705 9400 6735 9430
rect 6705 9330 6735 9360
rect 6705 9265 6735 9295
rect 6705 9205 6735 9235
rect 6705 9140 6735 9170
rect 6705 9070 6735 9100
rect 6705 9000 6735 9030
rect 6705 8930 6735 8960
rect 6705 8865 6735 8895
rect 6705 8805 6735 8835
rect 6705 8740 6735 8770
rect 6705 8670 6735 8700
rect 6705 8600 6735 8630
rect 6705 8530 6735 8560
rect 6705 8465 6735 8495
rect 6705 8405 6735 8435
rect 6705 8340 6735 8370
rect 6705 8270 6735 8300
rect 6705 8200 6735 8230
rect 6705 8130 6735 8160
rect 7625 9605 7655 9635
rect 7625 9540 7655 9570
rect 7625 9470 7655 9500
rect 7625 9400 7655 9430
rect 7625 9330 7655 9360
rect 7625 9265 7655 9295
rect 7625 9205 7655 9235
rect 7625 9140 7655 9170
rect 7625 9070 7655 9100
rect 7625 9000 7655 9030
rect 7625 8930 7655 8960
rect 7625 8865 7655 8895
rect 7625 8805 7655 8835
rect 7625 8740 7655 8770
rect 7625 8670 7655 8700
rect 7625 8600 7655 8630
rect 7625 8530 7655 8560
rect 7625 8465 7655 8495
rect 7625 8405 7655 8435
rect 7625 8340 7655 8370
rect 7625 8270 7655 8300
rect 7625 8200 7655 8230
rect 7625 8130 7655 8160
rect -75 195 -45 225
rect -75 130 -45 160
rect -75 60 -45 90
rect -75 -10 -45 20
rect -75 -80 -45 -50
rect -75 -145 -45 -115
rect -75 -205 -45 -175
rect -75 -270 -45 -240
rect -75 -340 -45 -310
rect -75 -410 -45 -380
rect -75 -480 -45 -450
rect -75 -545 -45 -515
rect -75 -605 -45 -575
rect -75 -670 -45 -640
rect -75 -740 -45 -710
rect -75 -810 -45 -780
rect -75 -880 -45 -850
rect -75 -945 -45 -915
rect -75 -1005 -45 -975
rect -75 -1070 -45 -1040
rect -75 -1140 -45 -1110
rect -75 -1210 -45 -1180
rect -75 -1280 -45 -1250
rect -75 -1345 -45 -1315
rect 275 195 305 225
rect 275 130 305 160
rect 275 60 305 90
rect 275 -10 305 20
rect 275 -80 305 -50
rect 275 -145 305 -115
rect 275 -205 305 -175
rect 275 -270 305 -240
rect 275 -340 305 -310
rect 275 -410 305 -380
rect 275 -480 305 -450
rect 275 -545 305 -515
rect 275 -605 305 -575
rect 275 -670 305 -640
rect 275 -740 305 -710
rect 275 -810 305 -780
rect 275 -880 305 -850
rect 275 -945 305 -915
rect 275 -1005 305 -975
rect 275 -1070 305 -1040
rect 275 -1140 305 -1110
rect 275 -1210 305 -1180
rect 275 -1280 305 -1250
rect 275 -1345 305 -1315
rect 625 195 655 225
rect 625 130 655 160
rect 625 60 655 90
rect 625 -10 655 20
rect 625 -80 655 -50
rect 625 -145 655 -115
rect 625 -205 655 -175
rect 625 -270 655 -240
rect 625 -340 655 -310
rect 625 -410 655 -380
rect 625 -480 655 -450
rect 625 -545 655 -515
rect 625 -605 655 -575
rect 625 -670 655 -640
rect 625 -740 655 -710
rect 625 -810 655 -780
rect 625 -880 655 -850
rect 625 -945 655 -915
rect 625 -1005 655 -975
rect 625 -1070 655 -1040
rect 625 -1140 655 -1110
rect 625 -1210 655 -1180
rect 625 -1280 655 -1250
rect 625 -1345 655 -1315
rect 975 195 1005 225
rect 975 130 1005 160
rect 975 60 1005 90
rect 975 -10 1005 20
rect 975 -80 1005 -50
rect 975 -145 1005 -115
rect 975 -205 1005 -175
rect 975 -270 1005 -240
rect 975 -340 1005 -310
rect 975 -410 1005 -380
rect 975 -480 1005 -450
rect 975 -545 1005 -515
rect 975 -605 1005 -575
rect 975 -670 1005 -640
rect 975 -740 1005 -710
rect 975 -810 1005 -780
rect 975 -880 1005 -850
rect 975 -945 1005 -915
rect 975 -1005 1005 -975
rect 975 -1070 1005 -1040
rect 975 -1140 1005 -1110
rect 975 -1210 1005 -1180
rect 975 -1280 1005 -1250
rect 975 -1345 1005 -1315
rect 1325 195 1355 225
rect 1325 130 1355 160
rect 1325 60 1355 90
rect 1325 -10 1355 20
rect 1325 -80 1355 -50
rect 1325 -145 1355 -115
rect 1325 -205 1355 -175
rect 1325 -270 1355 -240
rect 1325 -340 1355 -310
rect 1325 -410 1355 -380
rect 1325 -480 1355 -450
rect 1325 -545 1355 -515
rect 1325 -605 1355 -575
rect 1325 -670 1355 -640
rect 1325 -740 1355 -710
rect 1325 -810 1355 -780
rect 1325 -880 1355 -850
rect 1325 -945 1355 -915
rect 1325 -1005 1355 -975
rect 1325 -1070 1355 -1040
rect 1325 -1140 1355 -1110
rect 1325 -1210 1355 -1180
rect 1325 -1280 1355 -1250
rect 1325 -1345 1355 -1315
rect 1675 195 1705 225
rect 1675 130 1705 160
rect 1675 60 1705 90
rect 1675 -10 1705 20
rect 1675 -80 1705 -50
rect 1675 -145 1705 -115
rect 1675 -205 1705 -175
rect 1675 -270 1705 -240
rect 1675 -340 1705 -310
rect 1675 -410 1705 -380
rect 1675 -480 1705 -450
rect 1675 -545 1705 -515
rect 1675 -605 1705 -575
rect 1675 -670 1705 -640
rect 1675 -740 1705 -710
rect 1675 -810 1705 -780
rect 1675 -880 1705 -850
rect 1675 -945 1705 -915
rect 1675 -1005 1705 -975
rect 1675 -1070 1705 -1040
rect 1675 -1140 1705 -1110
rect 1675 -1210 1705 -1180
rect 1675 -1280 1705 -1250
rect 1675 -1345 1705 -1315
rect 2025 195 2055 225
rect 2025 130 2055 160
rect 2025 60 2055 90
rect 2025 -10 2055 20
rect 2025 -80 2055 -50
rect 2025 -145 2055 -115
rect 2025 -205 2055 -175
rect 2025 -270 2055 -240
rect 2025 -340 2055 -310
rect 2025 -410 2055 -380
rect 2025 -480 2055 -450
rect 2025 -545 2055 -515
rect 2025 -605 2055 -575
rect 2025 -670 2055 -640
rect 2025 -740 2055 -710
rect 2025 -810 2055 -780
rect 2025 -880 2055 -850
rect 2025 -945 2055 -915
rect 2025 -1005 2055 -975
rect 2025 -1070 2055 -1040
rect 2025 -1140 2055 -1110
rect 2025 -1210 2055 -1180
rect 2025 -1280 2055 -1250
rect 2025 -1345 2055 -1315
rect 2375 195 2405 225
rect 2375 130 2405 160
rect 2375 60 2405 90
rect 2375 -10 2405 20
rect 2375 -80 2405 -50
rect 2375 -145 2405 -115
rect 2375 -205 2405 -175
rect 2375 -270 2405 -240
rect 2375 -340 2405 -310
rect 2375 -410 2405 -380
rect 2375 -480 2405 -450
rect 2375 -545 2405 -515
rect 2375 -605 2405 -575
rect 2375 -670 2405 -640
rect 2375 -740 2405 -710
rect 2375 -810 2405 -780
rect 2375 -880 2405 -850
rect 2375 -945 2405 -915
rect 2375 -1005 2405 -975
rect 2375 -1070 2405 -1040
rect 2375 -1140 2405 -1110
rect 2375 -1210 2405 -1180
rect 2375 -1280 2405 -1250
rect 2375 -1345 2405 -1315
rect 2725 195 2755 225
rect 2725 130 2755 160
rect 2725 60 2755 90
rect 2725 -10 2755 20
rect 2725 -80 2755 -50
rect 2725 -145 2755 -115
rect 2725 -205 2755 -175
rect 2725 -270 2755 -240
rect 2725 -340 2755 -310
rect 2725 -410 2755 -380
rect 2725 -480 2755 -450
rect 2725 -545 2755 -515
rect 2725 -605 2755 -575
rect 2725 -670 2755 -640
rect 2725 -740 2755 -710
rect 2725 -810 2755 -780
rect 2725 -880 2755 -850
rect 2725 -945 2755 -915
rect 2725 -1005 2755 -975
rect 2725 -1070 2755 -1040
rect 2725 -1140 2755 -1110
rect 2725 -1210 2755 -1180
rect 2725 -1280 2755 -1250
rect 2725 -1345 2755 -1315
rect 3075 195 3105 225
rect 3075 130 3105 160
rect 3075 60 3105 90
rect 3075 -10 3105 20
rect 3075 -80 3105 -50
rect 3075 -145 3105 -115
rect 3075 -205 3105 -175
rect 3075 -270 3105 -240
rect 3075 -340 3105 -310
rect 3075 -410 3105 -380
rect 3075 -480 3105 -450
rect 3075 -545 3105 -515
rect 3075 -605 3105 -575
rect 3075 -670 3105 -640
rect 3075 -740 3105 -710
rect 3075 -810 3105 -780
rect 3075 -880 3105 -850
rect 3075 -945 3105 -915
rect 3075 -1005 3105 -975
rect 3075 -1070 3105 -1040
rect 3075 -1140 3105 -1110
rect 3075 -1210 3105 -1180
rect 3075 -1280 3105 -1250
rect 3075 -1345 3105 -1315
rect 3425 195 3455 225
rect 3425 130 3455 160
rect 3425 60 3455 90
rect 3425 -10 3455 20
rect 3425 -80 3455 -50
rect 3425 -145 3455 -115
rect 3425 -205 3455 -175
rect 3425 -270 3455 -240
rect 3425 -340 3455 -310
rect 3425 -410 3455 -380
rect 3425 -480 3455 -450
rect 3425 -545 3455 -515
rect 3425 -605 3455 -575
rect 3425 -670 3455 -640
rect 3425 -740 3455 -710
rect 3425 -810 3455 -780
rect 3425 -880 3455 -850
rect 3425 -945 3455 -915
rect 3425 -1005 3455 -975
rect 3425 -1070 3455 -1040
rect 3425 -1140 3455 -1110
rect 3425 -1210 3455 -1180
rect 3425 -1280 3455 -1250
rect 3425 -1345 3455 -1315
rect 3775 195 3805 225
rect 3775 130 3805 160
rect 3775 60 3805 90
rect 3775 -10 3805 20
rect 3775 -80 3805 -50
rect 3775 -145 3805 -115
rect 3775 -205 3805 -175
rect 3775 -270 3805 -240
rect 3775 -340 3805 -310
rect 3775 -410 3805 -380
rect 3775 -480 3805 -450
rect 3775 -545 3805 -515
rect 3775 -605 3805 -575
rect 3775 -670 3805 -640
rect 3775 -740 3805 -710
rect 3775 -810 3805 -780
rect 3775 -880 3805 -850
rect 3775 -945 3805 -915
rect 3775 -1005 3805 -975
rect 3775 -1070 3805 -1040
rect 3775 -1140 3805 -1110
rect 3775 -1210 3805 -1180
rect 3775 -1280 3805 -1250
rect 3775 -1345 3805 -1315
rect 4125 195 4155 225
rect 4125 130 4155 160
rect 4125 60 4155 90
rect 4125 -10 4155 20
rect 4125 -80 4155 -50
rect 4125 -145 4155 -115
rect 4125 -205 4155 -175
rect 4125 -270 4155 -240
rect 4125 -340 4155 -310
rect 4125 -410 4155 -380
rect 4125 -480 4155 -450
rect 4125 -545 4155 -515
rect 4125 -605 4155 -575
rect 4125 -670 4155 -640
rect 4125 -740 4155 -710
rect 4125 -810 4155 -780
rect 4125 -880 4155 -850
rect 4125 -945 4155 -915
rect 4125 -1005 4155 -975
rect 4125 -1070 4155 -1040
rect 4125 -1140 4155 -1110
rect 4125 -1210 4155 -1180
rect 4125 -1280 4155 -1250
rect 4125 -1345 4155 -1315
rect 4475 195 4505 225
rect 4475 130 4505 160
rect 4475 60 4505 90
rect 4475 -10 4505 20
rect 4475 -80 4505 -50
rect 4475 -145 4505 -115
rect 4475 -205 4505 -175
rect 4475 -270 4505 -240
rect 4475 -340 4505 -310
rect 4475 -410 4505 -380
rect 4475 -480 4505 -450
rect 4475 -545 4505 -515
rect 4475 -605 4505 -575
rect 4475 -670 4505 -640
rect 4475 -740 4505 -710
rect 4475 -810 4505 -780
rect 4475 -880 4505 -850
rect 4475 -945 4505 -915
rect 4475 -1005 4505 -975
rect 4475 -1070 4505 -1040
rect 4475 -1140 4505 -1110
rect 4475 -1210 4505 -1180
rect 4475 -1280 4505 -1250
rect 4475 -1345 4505 -1315
rect 4825 195 4855 225
rect 4825 130 4855 160
rect 4825 60 4855 90
rect 4825 -10 4855 20
rect 4825 -80 4855 -50
rect 4825 -145 4855 -115
rect 4825 -205 4855 -175
rect 4825 -270 4855 -240
rect 4825 -340 4855 -310
rect 4825 -410 4855 -380
rect 4825 -480 4855 -450
rect 4825 -545 4855 -515
rect 4825 -605 4855 -575
rect 4825 -670 4855 -640
rect 4825 -740 4855 -710
rect 4825 -810 4855 -780
rect 4825 -880 4855 -850
rect 4825 -945 4855 -915
rect 4825 -1005 4855 -975
rect 4825 -1070 4855 -1040
rect 4825 -1140 4855 -1110
rect 4825 -1210 4855 -1180
rect 4825 -1280 4855 -1250
rect 4825 -1345 4855 -1315
rect 5175 195 5205 225
rect 5175 130 5205 160
rect 5175 60 5205 90
rect 5175 -10 5205 20
rect 5175 -80 5205 -50
rect 5175 -145 5205 -115
rect 5175 -205 5205 -175
rect 5175 -270 5205 -240
rect 5175 -340 5205 -310
rect 5175 -410 5205 -380
rect 5175 -480 5205 -450
rect 5175 -545 5205 -515
rect 5175 -605 5205 -575
rect 5175 -670 5205 -640
rect 5175 -740 5205 -710
rect 5175 -810 5205 -780
rect 5175 -880 5205 -850
rect 5175 -945 5205 -915
rect 5175 -1005 5205 -975
rect 5175 -1070 5205 -1040
rect 5175 -1140 5205 -1110
rect 5175 -1210 5205 -1180
rect 5175 -1280 5205 -1250
rect 5175 -1345 5205 -1315
rect 5525 195 5555 225
rect 5525 130 5555 160
rect 5525 60 5555 90
rect 5525 -10 5555 20
rect 5525 -80 5555 -50
rect 5525 -145 5555 -115
rect 5525 -205 5555 -175
rect 5525 -270 5555 -240
rect 5525 -340 5555 -310
rect 5525 -410 5555 -380
rect 5525 -480 5555 -450
rect 5525 -545 5555 -515
rect 5525 -605 5555 -575
rect 5525 -670 5555 -640
rect 5525 -740 5555 -710
rect 5525 -810 5555 -780
rect 5525 -880 5555 -850
rect 5525 -945 5555 -915
rect 5525 -1005 5555 -975
rect 5525 -1070 5555 -1040
rect 5525 -1140 5555 -1110
rect 5525 -1210 5555 -1180
rect 5525 -1280 5555 -1250
rect 5525 -1345 5555 -1315
rect 5875 195 5905 225
rect 5875 130 5905 160
rect 5875 60 5905 90
rect 5875 -10 5905 20
rect 5875 -80 5905 -50
rect 5875 -145 5905 -115
rect 5875 -205 5905 -175
rect 5875 -270 5905 -240
rect 5875 -340 5905 -310
rect 5875 -410 5905 -380
rect 5875 -480 5905 -450
rect 5875 -545 5905 -515
rect 5875 -605 5905 -575
rect 5875 -670 5905 -640
rect 5875 -740 5905 -710
rect 5875 -810 5905 -780
rect 5875 -880 5905 -850
rect 5875 -945 5905 -915
rect 5875 -1005 5905 -975
rect 5875 -1070 5905 -1040
rect 5875 -1140 5905 -1110
rect 5875 -1210 5905 -1180
rect 5875 -1280 5905 -1250
rect 5875 -1345 5905 -1315
rect 6225 195 6255 225
rect 6225 130 6255 160
rect 6225 60 6255 90
rect 6225 -10 6255 20
rect 6225 -80 6255 -50
rect 6225 -145 6255 -115
rect 6225 -205 6255 -175
rect 6225 -270 6255 -240
rect 6225 -340 6255 -310
rect 6225 -410 6255 -380
rect 6225 -480 6255 -450
rect 6225 -545 6255 -515
rect 6225 -605 6255 -575
rect 6225 -670 6255 -640
rect 6225 -740 6255 -710
rect 6225 -810 6255 -780
rect 6225 -880 6255 -850
rect 6225 -945 6255 -915
rect 6225 -1005 6255 -975
rect 6225 -1070 6255 -1040
rect 6225 -1140 6255 -1110
rect 6225 -1210 6255 -1180
rect 6225 -1280 6255 -1250
rect 6225 -1345 6255 -1315
rect 6575 195 6605 225
rect 6575 130 6605 160
rect 6575 60 6605 90
rect 6575 -10 6605 20
rect 6575 -80 6605 -50
rect 6575 -145 6605 -115
rect 6575 -205 6605 -175
rect 6575 -270 6605 -240
rect 6575 -340 6605 -310
rect 6575 -410 6605 -380
rect 6575 -480 6605 -450
rect 6575 -545 6605 -515
rect 6575 -605 6605 -575
rect 6575 -670 6605 -640
rect 6575 -740 6605 -710
rect 6575 -810 6605 -780
rect 6575 -880 6605 -850
rect 6575 -945 6605 -915
rect 6575 -1005 6605 -975
rect 6575 -1070 6605 -1040
rect 6575 -1140 6605 -1110
rect 6575 -1210 6605 -1180
rect 6575 -1280 6605 -1250
rect 6575 -1345 6605 -1315
rect 6925 195 6955 225
rect 6925 130 6955 160
rect 6925 60 6955 90
rect 6925 -10 6955 20
rect 6925 -80 6955 -50
rect 6925 -145 6955 -115
rect 6925 -205 6955 -175
rect 6925 -270 6955 -240
rect 6925 -340 6955 -310
rect 6925 -410 6955 -380
rect 6925 -480 6955 -450
rect 6925 -545 6955 -515
rect 6925 -605 6955 -575
rect 6925 -670 6955 -640
rect 6925 -740 6955 -710
rect 6925 -810 6955 -780
rect 6925 -880 6955 -850
rect 6925 -945 6955 -915
rect 6925 -1005 6955 -975
rect 6925 -1070 6955 -1040
rect 6925 -1140 6955 -1110
rect 6925 -1210 6955 -1180
rect 6925 -1280 6955 -1250
rect 6925 -1345 6955 -1315
rect 7275 195 7305 225
rect 7275 130 7305 160
rect 7275 60 7305 90
rect 7275 -10 7305 20
rect 7275 -80 7305 -50
rect 7275 -145 7305 -115
rect 7275 -205 7305 -175
rect 7275 -270 7305 -240
rect 7275 -340 7305 -310
rect 7275 -410 7305 -380
rect 7275 -480 7305 -450
rect 7275 -545 7305 -515
rect 7275 -605 7305 -575
rect 7275 -670 7305 -640
rect 7275 -740 7305 -710
rect 7275 -810 7305 -780
rect 7275 -880 7305 -850
rect 7275 -945 7305 -915
rect 7275 -1005 7305 -975
rect 7275 -1070 7305 -1040
rect 7275 -1140 7305 -1110
rect 7275 -1210 7305 -1180
rect 7275 -1280 7305 -1250
rect 7275 -1345 7305 -1315
rect 7625 195 7655 225
rect 7625 130 7655 160
rect 7625 60 7655 90
rect 7625 -10 7655 20
rect 7625 -80 7655 -50
rect 7625 -145 7655 -115
rect 7625 -205 7655 -175
rect 7625 -270 7655 -240
rect 7625 -340 7655 -310
rect 7625 -410 7655 -380
rect 7625 -480 7655 -450
rect 7625 -545 7655 -515
rect 7625 -605 7655 -575
rect 7625 -670 7655 -640
rect 7625 -740 7655 -710
rect 7625 -810 7655 -780
rect 7625 -880 7655 -850
rect 7625 -945 7655 -915
rect 7625 -1005 7655 -975
rect 7625 -1070 7655 -1040
rect 7625 -1140 7655 -1110
rect 7625 -1210 7655 -1180
rect 7625 -1280 7655 -1250
rect 7625 -1345 7655 -1315
rect 7975 195 8005 225
rect 7975 130 8005 160
rect 7975 60 8005 90
rect 7975 -10 8005 20
rect 7975 -80 8005 -50
rect 7975 -145 8005 -115
rect 7975 -205 8005 -175
rect 7975 -270 8005 -240
rect 7975 -340 8005 -310
rect 7975 -410 8005 -380
rect 7975 -480 8005 -450
rect 7975 -545 8005 -515
rect 7975 -605 8005 -575
rect 7975 -670 8005 -640
rect 7975 -740 8005 -710
rect 7975 -810 8005 -780
rect 7975 -880 8005 -850
rect 7975 -945 8005 -915
rect 7975 -1005 8005 -975
rect 7975 -1070 8005 -1040
rect 7975 -1140 8005 -1110
rect 7975 -1210 8005 -1180
rect 7975 -1280 8005 -1250
rect 7975 -1345 8005 -1315
rect 8325 195 8355 225
rect 8325 130 8355 160
rect 8325 60 8355 90
rect 8325 -10 8355 20
rect 8325 -80 8355 -50
rect 8325 -145 8355 -115
rect 8325 -205 8355 -175
rect 8325 -270 8355 -240
rect 8325 -340 8355 -310
rect 8325 -410 8355 -380
rect 8325 -480 8355 -450
rect 8325 -545 8355 -515
rect 8325 -605 8355 -575
rect 8325 -670 8355 -640
rect 8325 -740 8355 -710
rect 8325 -810 8355 -780
rect 8325 -880 8355 -850
rect 8325 -945 8355 -915
rect 8325 -1005 8355 -975
rect 8325 -1070 8355 -1040
rect 8325 -1140 8355 -1110
rect 8325 -1210 8355 -1180
rect 8325 -1280 8355 -1250
rect 8325 -1345 8355 -1315
rect 8675 195 8705 225
rect 8675 130 8705 160
rect 8675 60 8705 90
rect 8675 -10 8705 20
rect 8675 -80 8705 -50
rect 8675 -145 8705 -115
rect 8675 -205 8705 -175
rect 8675 -270 8705 -240
rect 8675 -340 8705 -310
rect 8675 -410 8705 -380
rect 8675 -480 8705 -450
rect 8675 -545 8705 -515
rect 8675 -605 8705 -575
rect 8675 -670 8705 -640
rect 8675 -740 8705 -710
rect 8675 -810 8705 -780
rect 8675 -880 8705 -850
rect 8675 -945 8705 -915
rect 8675 -1005 8705 -975
rect 8675 -1070 8705 -1040
rect 8675 -1140 8705 -1110
rect 8675 -1210 8705 -1180
rect 8675 -1280 8705 -1250
rect 8675 -1345 8705 -1315
rect 9025 195 9055 225
rect 9025 130 9055 160
rect 9025 60 9055 90
rect 9025 -10 9055 20
rect 9025 -80 9055 -50
rect 9025 -145 9055 -115
rect 9025 -205 9055 -175
rect 9025 -270 9055 -240
rect 9025 -340 9055 -310
rect 9025 -410 9055 -380
rect 9025 -480 9055 -450
rect 9025 -545 9055 -515
rect 9025 -605 9055 -575
rect 9025 -670 9055 -640
rect 9025 -740 9055 -710
rect 9025 -810 9055 -780
rect 9025 -880 9055 -850
rect 9025 -945 9055 -915
rect 9025 -1005 9055 -975
rect 9025 -1070 9055 -1040
rect 9025 -1140 9055 -1110
rect 9025 -1210 9055 -1180
rect 9025 -1280 9055 -1250
rect 9025 -1345 9055 -1315
<< metal3 >>
rect 2100 19315 2160 19325
rect 2100 19275 2110 19315
rect 2150 19275 2160 19315
rect 2100 19250 2160 19275
rect 2100 19210 2110 19250
rect 2150 19210 2160 19250
rect 2100 19180 2160 19210
rect 2100 19140 2110 19180
rect 2150 19140 2160 19180
rect 2100 19110 2160 19140
rect 2100 19070 2110 19110
rect 2150 19070 2160 19110
rect 2100 19040 2160 19070
rect 2100 19000 2110 19040
rect 2150 19000 2160 19040
rect 2100 18975 2160 19000
rect 2100 18935 2110 18975
rect 2150 18935 2160 18975
rect 2100 18915 2160 18935
rect 2100 18875 2110 18915
rect 2150 18875 2160 18915
rect 2100 18850 2160 18875
rect 2100 18810 2110 18850
rect 2150 18810 2160 18850
rect 2100 18780 2160 18810
rect 2100 18740 2110 18780
rect 2150 18740 2160 18780
rect 2100 18710 2160 18740
rect 2100 18670 2110 18710
rect 2150 18670 2160 18710
rect 2100 18640 2160 18670
rect 2100 18600 2110 18640
rect 2150 18600 2160 18640
rect 2100 18575 2160 18600
rect 2100 18535 2110 18575
rect 2150 18535 2160 18575
rect 2100 18515 2160 18535
rect 2100 18475 2110 18515
rect 2150 18475 2160 18515
rect 2100 18450 2160 18475
rect 2100 18410 2110 18450
rect 2150 18410 2160 18450
rect 2100 18380 2160 18410
rect 2100 18340 2110 18380
rect 2150 18340 2160 18380
rect 2100 18310 2160 18340
rect 2100 18270 2110 18310
rect 2150 18270 2160 18310
rect 2100 18240 2160 18270
rect 2100 18200 2110 18240
rect 2150 18200 2160 18240
rect 2100 18175 2160 18200
rect 2100 18135 2110 18175
rect 2150 18135 2160 18175
rect 2100 18115 2160 18135
rect 2100 18075 2110 18115
rect 2150 18075 2160 18115
rect 2100 18050 2160 18075
rect 2100 18010 2110 18050
rect 2150 18010 2160 18050
rect 2100 17980 2160 18010
rect 2100 17940 2110 17980
rect 2150 17940 2160 17980
rect 2100 17910 2160 17940
rect 2100 17870 2110 17910
rect 2150 17870 2160 17910
rect 2100 17840 2160 17870
rect 2100 17800 2110 17840
rect 2150 17800 2160 17840
rect 2100 17775 2160 17800
rect 2100 17735 2110 17775
rect 2150 17735 2160 17775
rect 2100 17725 2160 17735
rect 6690 19315 6750 19325
rect 6690 19275 6700 19315
rect 6740 19275 6750 19315
rect 6690 19250 6750 19275
rect 6690 19210 6700 19250
rect 6740 19210 6750 19250
rect 6690 19180 6750 19210
rect 6690 19140 6700 19180
rect 6740 19140 6750 19180
rect 6690 19110 6750 19140
rect 6690 19070 6700 19110
rect 6740 19070 6750 19110
rect 6690 19040 6750 19070
rect 6690 19000 6700 19040
rect 6740 19000 6750 19040
rect 6690 18975 6750 19000
rect 6690 18935 6700 18975
rect 6740 18935 6750 18975
rect 6690 18915 6750 18935
rect 6690 18875 6700 18915
rect 6740 18875 6750 18915
rect 6690 18850 6750 18875
rect 6690 18810 6700 18850
rect 6740 18810 6750 18850
rect 6690 18780 6750 18810
rect 6690 18740 6700 18780
rect 6740 18740 6750 18780
rect 6690 18710 6750 18740
rect 6690 18670 6700 18710
rect 6740 18670 6750 18710
rect 6690 18640 6750 18670
rect 6690 18600 6700 18640
rect 6740 18600 6750 18640
rect 6690 18575 6750 18600
rect 6690 18535 6700 18575
rect 6740 18535 6750 18575
rect 6690 18515 6750 18535
rect 6690 18475 6700 18515
rect 6740 18475 6750 18515
rect 6690 18450 6750 18475
rect 6690 18410 6700 18450
rect 6740 18410 6750 18450
rect 6690 18380 6750 18410
rect 6690 18340 6700 18380
rect 6740 18340 6750 18380
rect 6690 18310 6750 18340
rect 6690 18270 6700 18310
rect 6740 18270 6750 18310
rect 6690 18240 6750 18270
rect 6690 18200 6700 18240
rect 6740 18200 6750 18240
rect 6690 18175 6750 18200
rect 6690 18135 6700 18175
rect 6740 18135 6750 18175
rect 6690 18115 6750 18135
rect 6690 18075 6700 18115
rect 6740 18075 6750 18115
rect 6690 18050 6750 18075
rect 6690 18010 6700 18050
rect 6740 18010 6750 18050
rect 6690 17980 6750 18010
rect 6690 17940 6700 17980
rect 6740 17940 6750 17980
rect 6690 17910 6750 17940
rect 6690 17870 6700 17910
rect 6740 17870 6750 17910
rect 6690 17840 6750 17870
rect 6690 17800 6700 17840
rect 6740 17800 6750 17840
rect 6690 17775 6750 17800
rect 6690 17735 6700 17775
rect 6740 17735 6750 17775
rect 6690 17725 6750 17735
rect 31290 19305 32890 19325
rect 31290 19270 31305 19305
rect 31340 19270 31350 19305
rect 31385 19270 31395 19305
rect 31430 19270 31440 19305
rect 31475 19270 31485 19305
rect 31520 19270 31530 19305
rect 31565 19270 31575 19305
rect 31610 19270 31620 19305
rect 31655 19270 31665 19305
rect 31700 19270 31710 19305
rect 31745 19270 31755 19305
rect 31790 19270 31800 19305
rect 31835 19270 31845 19305
rect 31880 19270 31890 19305
rect 31925 19270 31935 19305
rect 31970 19270 31980 19305
rect 32015 19270 32025 19305
rect 32060 19270 32070 19305
rect 32105 19270 32115 19305
rect 32150 19270 32160 19305
rect 32195 19270 32205 19305
rect 32240 19270 32250 19305
rect 32285 19270 32295 19305
rect 32330 19270 32340 19305
rect 32375 19270 32385 19305
rect 32420 19270 32430 19305
rect 32465 19270 32475 19305
rect 32510 19270 32520 19305
rect 32555 19270 32565 19305
rect 32600 19270 32610 19305
rect 32645 19270 32655 19305
rect 32690 19270 32700 19305
rect 32735 19270 32745 19305
rect 32780 19270 32790 19305
rect 32825 19270 32835 19305
rect 32870 19270 32890 19305
rect 31290 19260 32890 19270
rect 31290 19225 31305 19260
rect 31340 19225 31350 19260
rect 31385 19225 31395 19260
rect 31430 19225 31440 19260
rect 31475 19225 31485 19260
rect 31520 19225 31530 19260
rect 31565 19225 31575 19260
rect 31610 19225 31620 19260
rect 31655 19225 31665 19260
rect 31700 19225 31710 19260
rect 31745 19225 31755 19260
rect 31790 19225 31800 19260
rect 31835 19225 31845 19260
rect 31880 19225 31890 19260
rect 31925 19225 31935 19260
rect 31970 19225 31980 19260
rect 32015 19225 32025 19260
rect 32060 19225 32070 19260
rect 32105 19225 32115 19260
rect 32150 19225 32160 19260
rect 32195 19225 32205 19260
rect 32240 19225 32250 19260
rect 32285 19225 32295 19260
rect 32330 19225 32340 19260
rect 32375 19225 32385 19260
rect 32420 19225 32430 19260
rect 32465 19225 32475 19260
rect 32510 19225 32520 19260
rect 32555 19225 32565 19260
rect 32600 19225 32610 19260
rect 32645 19225 32655 19260
rect 32690 19225 32700 19260
rect 32735 19225 32745 19260
rect 32780 19225 32790 19260
rect 32825 19225 32835 19260
rect 32870 19225 32890 19260
rect 31290 19215 32890 19225
rect 31290 19180 31305 19215
rect 31340 19180 31350 19215
rect 31385 19180 31395 19215
rect 31430 19180 31440 19215
rect 31475 19180 31485 19215
rect 31520 19180 31530 19215
rect 31565 19180 31575 19215
rect 31610 19180 31620 19215
rect 31655 19180 31665 19215
rect 31700 19180 31710 19215
rect 31745 19180 31755 19215
rect 31790 19180 31800 19215
rect 31835 19180 31845 19215
rect 31880 19180 31890 19215
rect 31925 19180 31935 19215
rect 31970 19180 31980 19215
rect 32015 19180 32025 19215
rect 32060 19180 32070 19215
rect 32105 19180 32115 19215
rect 32150 19180 32160 19215
rect 32195 19180 32205 19215
rect 32240 19180 32250 19215
rect 32285 19180 32295 19215
rect 32330 19180 32340 19215
rect 32375 19180 32385 19215
rect 32420 19180 32430 19215
rect 32465 19180 32475 19215
rect 32510 19180 32520 19215
rect 32555 19180 32565 19215
rect 32600 19180 32610 19215
rect 32645 19180 32655 19215
rect 32690 19180 32700 19215
rect 32735 19180 32745 19215
rect 32780 19180 32790 19215
rect 32825 19180 32835 19215
rect 32870 19180 32890 19215
rect 31290 19170 32890 19180
rect 31290 19135 31305 19170
rect 31340 19135 31350 19170
rect 31385 19135 31395 19170
rect 31430 19135 31440 19170
rect 31475 19135 31485 19170
rect 31520 19135 31530 19170
rect 31565 19135 31575 19170
rect 31610 19135 31620 19170
rect 31655 19135 31665 19170
rect 31700 19135 31710 19170
rect 31745 19135 31755 19170
rect 31790 19135 31800 19170
rect 31835 19135 31845 19170
rect 31880 19135 31890 19170
rect 31925 19135 31935 19170
rect 31970 19135 31980 19170
rect 32015 19135 32025 19170
rect 32060 19135 32070 19170
rect 32105 19135 32115 19170
rect 32150 19135 32160 19170
rect 32195 19135 32205 19170
rect 32240 19135 32250 19170
rect 32285 19135 32295 19170
rect 32330 19135 32340 19170
rect 32375 19135 32385 19170
rect 32420 19135 32430 19170
rect 32465 19135 32475 19170
rect 32510 19135 32520 19170
rect 32555 19135 32565 19170
rect 32600 19135 32610 19170
rect 32645 19135 32655 19170
rect 32690 19135 32700 19170
rect 32735 19135 32745 19170
rect 32780 19135 32790 19170
rect 32825 19135 32835 19170
rect 32870 19135 32890 19170
rect 31290 19125 32890 19135
rect 31290 19090 31305 19125
rect 31340 19090 31350 19125
rect 31385 19090 31395 19125
rect 31430 19090 31440 19125
rect 31475 19090 31485 19125
rect 31520 19090 31530 19125
rect 31565 19090 31575 19125
rect 31610 19090 31620 19125
rect 31655 19090 31665 19125
rect 31700 19090 31710 19125
rect 31745 19090 31755 19125
rect 31790 19090 31800 19125
rect 31835 19090 31845 19125
rect 31880 19090 31890 19125
rect 31925 19090 31935 19125
rect 31970 19090 31980 19125
rect 32015 19090 32025 19125
rect 32060 19090 32070 19125
rect 32105 19090 32115 19125
rect 32150 19090 32160 19125
rect 32195 19090 32205 19125
rect 32240 19090 32250 19125
rect 32285 19090 32295 19125
rect 32330 19090 32340 19125
rect 32375 19090 32385 19125
rect 32420 19090 32430 19125
rect 32465 19090 32475 19125
rect 32510 19090 32520 19125
rect 32555 19090 32565 19125
rect 32600 19090 32610 19125
rect 32645 19090 32655 19125
rect 32690 19090 32700 19125
rect 32735 19090 32745 19125
rect 32780 19090 32790 19125
rect 32825 19090 32835 19125
rect 32870 19090 32890 19125
rect 31290 19080 32890 19090
rect 31290 19045 31305 19080
rect 31340 19045 31350 19080
rect 31385 19045 31395 19080
rect 31430 19045 31440 19080
rect 31475 19045 31485 19080
rect 31520 19045 31530 19080
rect 31565 19045 31575 19080
rect 31610 19045 31620 19080
rect 31655 19045 31665 19080
rect 31700 19045 31710 19080
rect 31745 19045 31755 19080
rect 31790 19045 31800 19080
rect 31835 19045 31845 19080
rect 31880 19045 31890 19080
rect 31925 19045 31935 19080
rect 31970 19045 31980 19080
rect 32015 19045 32025 19080
rect 32060 19045 32070 19080
rect 32105 19045 32115 19080
rect 32150 19045 32160 19080
rect 32195 19045 32205 19080
rect 32240 19045 32250 19080
rect 32285 19045 32295 19080
rect 32330 19045 32340 19080
rect 32375 19045 32385 19080
rect 32420 19045 32430 19080
rect 32465 19045 32475 19080
rect 32510 19045 32520 19080
rect 32555 19045 32565 19080
rect 32600 19045 32610 19080
rect 32645 19045 32655 19080
rect 32690 19045 32700 19080
rect 32735 19045 32745 19080
rect 32780 19045 32790 19080
rect 32825 19045 32835 19080
rect 32870 19045 32890 19080
rect 31290 19035 32890 19045
rect 31290 19000 31305 19035
rect 31340 19000 31350 19035
rect 31385 19000 31395 19035
rect 31430 19000 31440 19035
rect 31475 19000 31485 19035
rect 31520 19000 31530 19035
rect 31565 19000 31575 19035
rect 31610 19000 31620 19035
rect 31655 19000 31665 19035
rect 31700 19000 31710 19035
rect 31745 19000 31755 19035
rect 31790 19000 31800 19035
rect 31835 19000 31845 19035
rect 31880 19000 31890 19035
rect 31925 19000 31935 19035
rect 31970 19000 31980 19035
rect 32015 19000 32025 19035
rect 32060 19000 32070 19035
rect 32105 19000 32115 19035
rect 32150 19000 32160 19035
rect 32195 19000 32205 19035
rect 32240 19000 32250 19035
rect 32285 19000 32295 19035
rect 32330 19000 32340 19035
rect 32375 19000 32385 19035
rect 32420 19000 32430 19035
rect 32465 19000 32475 19035
rect 32510 19000 32520 19035
rect 32555 19000 32565 19035
rect 32600 19000 32610 19035
rect 32645 19000 32655 19035
rect 32690 19000 32700 19035
rect 32735 19000 32745 19035
rect 32780 19000 32790 19035
rect 32825 19000 32835 19035
rect 32870 19000 32890 19035
rect 31290 18990 32890 19000
rect 31290 18955 31305 18990
rect 31340 18955 31350 18990
rect 31385 18955 31395 18990
rect 31430 18955 31440 18990
rect 31475 18955 31485 18990
rect 31520 18955 31530 18990
rect 31565 18955 31575 18990
rect 31610 18955 31620 18990
rect 31655 18955 31665 18990
rect 31700 18955 31710 18990
rect 31745 18955 31755 18990
rect 31790 18955 31800 18990
rect 31835 18955 31845 18990
rect 31880 18955 31890 18990
rect 31925 18955 31935 18990
rect 31970 18955 31980 18990
rect 32015 18955 32025 18990
rect 32060 18955 32070 18990
rect 32105 18955 32115 18990
rect 32150 18955 32160 18990
rect 32195 18955 32205 18990
rect 32240 18955 32250 18990
rect 32285 18955 32295 18990
rect 32330 18955 32340 18990
rect 32375 18955 32385 18990
rect 32420 18955 32430 18990
rect 32465 18955 32475 18990
rect 32510 18955 32520 18990
rect 32555 18955 32565 18990
rect 32600 18955 32610 18990
rect 32645 18955 32655 18990
rect 32690 18955 32700 18990
rect 32735 18955 32745 18990
rect 32780 18955 32790 18990
rect 32825 18955 32835 18990
rect 32870 18955 32890 18990
rect 31290 18945 32890 18955
rect 31290 18910 31305 18945
rect 31340 18910 31350 18945
rect 31385 18910 31395 18945
rect 31430 18910 31440 18945
rect 31475 18910 31485 18945
rect 31520 18910 31530 18945
rect 31565 18910 31575 18945
rect 31610 18910 31620 18945
rect 31655 18910 31665 18945
rect 31700 18910 31710 18945
rect 31745 18910 31755 18945
rect 31790 18910 31800 18945
rect 31835 18910 31845 18945
rect 31880 18910 31890 18945
rect 31925 18910 31935 18945
rect 31970 18910 31980 18945
rect 32015 18910 32025 18945
rect 32060 18910 32070 18945
rect 32105 18910 32115 18945
rect 32150 18910 32160 18945
rect 32195 18910 32205 18945
rect 32240 18910 32250 18945
rect 32285 18910 32295 18945
rect 32330 18910 32340 18945
rect 32375 18910 32385 18945
rect 32420 18910 32430 18945
rect 32465 18910 32475 18945
rect 32510 18910 32520 18945
rect 32555 18910 32565 18945
rect 32600 18910 32610 18945
rect 32645 18910 32655 18945
rect 32690 18910 32700 18945
rect 32735 18910 32745 18945
rect 32780 18910 32790 18945
rect 32825 18910 32835 18945
rect 32870 18910 32890 18945
rect 31290 18900 32890 18910
rect 31290 18865 31305 18900
rect 31340 18865 31350 18900
rect 31385 18865 31395 18900
rect 31430 18865 31440 18900
rect 31475 18865 31485 18900
rect 31520 18865 31530 18900
rect 31565 18865 31575 18900
rect 31610 18865 31620 18900
rect 31655 18865 31665 18900
rect 31700 18865 31710 18900
rect 31745 18865 31755 18900
rect 31790 18865 31800 18900
rect 31835 18865 31845 18900
rect 31880 18865 31890 18900
rect 31925 18865 31935 18900
rect 31970 18865 31980 18900
rect 32015 18865 32025 18900
rect 32060 18865 32070 18900
rect 32105 18865 32115 18900
rect 32150 18865 32160 18900
rect 32195 18865 32205 18900
rect 32240 18865 32250 18900
rect 32285 18865 32295 18900
rect 32330 18865 32340 18900
rect 32375 18865 32385 18900
rect 32420 18865 32430 18900
rect 32465 18865 32475 18900
rect 32510 18865 32520 18900
rect 32555 18865 32565 18900
rect 32600 18865 32610 18900
rect 32645 18865 32655 18900
rect 32690 18865 32700 18900
rect 32735 18865 32745 18900
rect 32780 18865 32790 18900
rect 32825 18865 32835 18900
rect 32870 18865 32890 18900
rect 31290 18855 32890 18865
rect 31290 18820 31305 18855
rect 31340 18820 31350 18855
rect 31385 18820 31395 18855
rect 31430 18820 31440 18855
rect 31475 18820 31485 18855
rect 31520 18820 31530 18855
rect 31565 18820 31575 18855
rect 31610 18820 31620 18855
rect 31655 18820 31665 18855
rect 31700 18820 31710 18855
rect 31745 18820 31755 18855
rect 31790 18820 31800 18855
rect 31835 18820 31845 18855
rect 31880 18820 31890 18855
rect 31925 18820 31935 18855
rect 31970 18820 31980 18855
rect 32015 18820 32025 18855
rect 32060 18820 32070 18855
rect 32105 18820 32115 18855
rect 32150 18820 32160 18855
rect 32195 18820 32205 18855
rect 32240 18820 32250 18855
rect 32285 18820 32295 18855
rect 32330 18820 32340 18855
rect 32375 18820 32385 18855
rect 32420 18820 32430 18855
rect 32465 18820 32475 18855
rect 32510 18820 32520 18855
rect 32555 18820 32565 18855
rect 32600 18820 32610 18855
rect 32645 18820 32655 18855
rect 32690 18820 32700 18855
rect 32735 18820 32745 18855
rect 32780 18820 32790 18855
rect 32825 18820 32835 18855
rect 32870 18820 32890 18855
rect 31290 18810 32890 18820
rect 31290 18775 31305 18810
rect 31340 18775 31350 18810
rect 31385 18775 31395 18810
rect 31430 18775 31440 18810
rect 31475 18775 31485 18810
rect 31520 18775 31530 18810
rect 31565 18775 31575 18810
rect 31610 18775 31620 18810
rect 31655 18775 31665 18810
rect 31700 18775 31710 18810
rect 31745 18775 31755 18810
rect 31790 18775 31800 18810
rect 31835 18775 31845 18810
rect 31880 18775 31890 18810
rect 31925 18775 31935 18810
rect 31970 18775 31980 18810
rect 32015 18775 32025 18810
rect 32060 18775 32070 18810
rect 32105 18775 32115 18810
rect 32150 18775 32160 18810
rect 32195 18775 32205 18810
rect 32240 18775 32250 18810
rect 32285 18775 32295 18810
rect 32330 18775 32340 18810
rect 32375 18775 32385 18810
rect 32420 18775 32430 18810
rect 32465 18775 32475 18810
rect 32510 18775 32520 18810
rect 32555 18775 32565 18810
rect 32600 18775 32610 18810
rect 32645 18775 32655 18810
rect 32690 18775 32700 18810
rect 32735 18775 32745 18810
rect 32780 18775 32790 18810
rect 32825 18775 32835 18810
rect 32870 18775 32890 18810
rect 31290 18765 32890 18775
rect 31290 18730 31305 18765
rect 31340 18730 31350 18765
rect 31385 18730 31395 18765
rect 31430 18730 31440 18765
rect 31475 18730 31485 18765
rect 31520 18730 31530 18765
rect 31565 18730 31575 18765
rect 31610 18730 31620 18765
rect 31655 18730 31665 18765
rect 31700 18730 31710 18765
rect 31745 18730 31755 18765
rect 31790 18730 31800 18765
rect 31835 18730 31845 18765
rect 31880 18730 31890 18765
rect 31925 18730 31935 18765
rect 31970 18730 31980 18765
rect 32015 18730 32025 18765
rect 32060 18730 32070 18765
rect 32105 18730 32115 18765
rect 32150 18730 32160 18765
rect 32195 18730 32205 18765
rect 32240 18730 32250 18765
rect 32285 18730 32295 18765
rect 32330 18730 32340 18765
rect 32375 18730 32385 18765
rect 32420 18730 32430 18765
rect 32465 18730 32475 18765
rect 32510 18730 32520 18765
rect 32555 18730 32565 18765
rect 32600 18730 32610 18765
rect 32645 18730 32655 18765
rect 32690 18730 32700 18765
rect 32735 18730 32745 18765
rect 32780 18730 32790 18765
rect 32825 18730 32835 18765
rect 32870 18730 32890 18765
rect 31290 18720 32890 18730
rect 31290 18685 31305 18720
rect 31340 18685 31350 18720
rect 31385 18685 31395 18720
rect 31430 18685 31440 18720
rect 31475 18685 31485 18720
rect 31520 18685 31530 18720
rect 31565 18685 31575 18720
rect 31610 18685 31620 18720
rect 31655 18685 31665 18720
rect 31700 18685 31710 18720
rect 31745 18685 31755 18720
rect 31790 18685 31800 18720
rect 31835 18685 31845 18720
rect 31880 18685 31890 18720
rect 31925 18685 31935 18720
rect 31970 18685 31980 18720
rect 32015 18685 32025 18720
rect 32060 18685 32070 18720
rect 32105 18685 32115 18720
rect 32150 18685 32160 18720
rect 32195 18685 32205 18720
rect 32240 18685 32250 18720
rect 32285 18685 32295 18720
rect 32330 18685 32340 18720
rect 32375 18685 32385 18720
rect 32420 18685 32430 18720
rect 32465 18685 32475 18720
rect 32510 18685 32520 18720
rect 32555 18685 32565 18720
rect 32600 18685 32610 18720
rect 32645 18685 32655 18720
rect 32690 18685 32700 18720
rect 32735 18685 32745 18720
rect 32780 18685 32790 18720
rect 32825 18685 32835 18720
rect 32870 18685 32890 18720
rect 31290 18675 32890 18685
rect 31290 18640 31305 18675
rect 31340 18640 31350 18675
rect 31385 18640 31395 18675
rect 31430 18640 31440 18675
rect 31475 18640 31485 18675
rect 31520 18640 31530 18675
rect 31565 18640 31575 18675
rect 31610 18640 31620 18675
rect 31655 18640 31665 18675
rect 31700 18640 31710 18675
rect 31745 18640 31755 18675
rect 31790 18640 31800 18675
rect 31835 18640 31845 18675
rect 31880 18640 31890 18675
rect 31925 18640 31935 18675
rect 31970 18640 31980 18675
rect 32015 18640 32025 18675
rect 32060 18640 32070 18675
rect 32105 18640 32115 18675
rect 32150 18640 32160 18675
rect 32195 18640 32205 18675
rect 32240 18640 32250 18675
rect 32285 18640 32295 18675
rect 32330 18640 32340 18675
rect 32375 18640 32385 18675
rect 32420 18640 32430 18675
rect 32465 18640 32475 18675
rect 32510 18640 32520 18675
rect 32555 18640 32565 18675
rect 32600 18640 32610 18675
rect 32645 18640 32655 18675
rect 32690 18640 32700 18675
rect 32735 18640 32745 18675
rect 32780 18640 32790 18675
rect 32825 18640 32835 18675
rect 32870 18640 32890 18675
rect 31290 18630 32890 18640
rect 31290 18595 31305 18630
rect 31340 18595 31350 18630
rect 31385 18595 31395 18630
rect 31430 18595 31440 18630
rect 31475 18595 31485 18630
rect 31520 18595 31530 18630
rect 31565 18595 31575 18630
rect 31610 18595 31620 18630
rect 31655 18595 31665 18630
rect 31700 18595 31710 18630
rect 31745 18595 31755 18630
rect 31790 18595 31800 18630
rect 31835 18595 31845 18630
rect 31880 18595 31890 18630
rect 31925 18595 31935 18630
rect 31970 18595 31980 18630
rect 32015 18595 32025 18630
rect 32060 18595 32070 18630
rect 32105 18595 32115 18630
rect 32150 18595 32160 18630
rect 32195 18595 32205 18630
rect 32240 18595 32250 18630
rect 32285 18595 32295 18630
rect 32330 18595 32340 18630
rect 32375 18595 32385 18630
rect 32420 18595 32430 18630
rect 32465 18595 32475 18630
rect 32510 18595 32520 18630
rect 32555 18595 32565 18630
rect 32600 18595 32610 18630
rect 32645 18595 32655 18630
rect 32690 18595 32700 18630
rect 32735 18595 32745 18630
rect 32780 18595 32790 18630
rect 32825 18595 32835 18630
rect 32870 18595 32890 18630
rect 31290 18585 32890 18595
rect 31290 18550 31305 18585
rect 31340 18550 31350 18585
rect 31385 18550 31395 18585
rect 31430 18550 31440 18585
rect 31475 18550 31485 18585
rect 31520 18550 31530 18585
rect 31565 18550 31575 18585
rect 31610 18550 31620 18585
rect 31655 18550 31665 18585
rect 31700 18550 31710 18585
rect 31745 18550 31755 18585
rect 31790 18550 31800 18585
rect 31835 18550 31845 18585
rect 31880 18550 31890 18585
rect 31925 18550 31935 18585
rect 31970 18550 31980 18585
rect 32015 18550 32025 18585
rect 32060 18550 32070 18585
rect 32105 18550 32115 18585
rect 32150 18550 32160 18585
rect 32195 18550 32205 18585
rect 32240 18550 32250 18585
rect 32285 18550 32295 18585
rect 32330 18550 32340 18585
rect 32375 18550 32385 18585
rect 32420 18550 32430 18585
rect 32465 18550 32475 18585
rect 32510 18550 32520 18585
rect 32555 18550 32565 18585
rect 32600 18550 32610 18585
rect 32645 18550 32655 18585
rect 32690 18550 32700 18585
rect 32735 18550 32745 18585
rect 32780 18550 32790 18585
rect 32825 18550 32835 18585
rect 32870 18550 32890 18585
rect 31290 18540 32890 18550
rect 31290 18505 31305 18540
rect 31340 18505 31350 18540
rect 31385 18505 31395 18540
rect 31430 18505 31440 18540
rect 31475 18505 31485 18540
rect 31520 18505 31530 18540
rect 31565 18505 31575 18540
rect 31610 18505 31620 18540
rect 31655 18505 31665 18540
rect 31700 18505 31710 18540
rect 31745 18505 31755 18540
rect 31790 18505 31800 18540
rect 31835 18505 31845 18540
rect 31880 18505 31890 18540
rect 31925 18505 31935 18540
rect 31970 18505 31980 18540
rect 32015 18505 32025 18540
rect 32060 18505 32070 18540
rect 32105 18505 32115 18540
rect 32150 18505 32160 18540
rect 32195 18505 32205 18540
rect 32240 18505 32250 18540
rect 32285 18505 32295 18540
rect 32330 18505 32340 18540
rect 32375 18505 32385 18540
rect 32420 18505 32430 18540
rect 32465 18505 32475 18540
rect 32510 18505 32520 18540
rect 32555 18505 32565 18540
rect 32600 18505 32610 18540
rect 32645 18505 32655 18540
rect 32690 18505 32700 18540
rect 32735 18505 32745 18540
rect 32780 18505 32790 18540
rect 32825 18505 32835 18540
rect 32870 18505 32890 18540
rect 31290 18495 32890 18505
rect 31290 18460 31305 18495
rect 31340 18460 31350 18495
rect 31385 18460 31395 18495
rect 31430 18460 31440 18495
rect 31475 18460 31485 18495
rect 31520 18460 31530 18495
rect 31565 18460 31575 18495
rect 31610 18460 31620 18495
rect 31655 18460 31665 18495
rect 31700 18460 31710 18495
rect 31745 18460 31755 18495
rect 31790 18460 31800 18495
rect 31835 18460 31845 18495
rect 31880 18460 31890 18495
rect 31925 18460 31935 18495
rect 31970 18460 31980 18495
rect 32015 18460 32025 18495
rect 32060 18460 32070 18495
rect 32105 18460 32115 18495
rect 32150 18460 32160 18495
rect 32195 18460 32205 18495
rect 32240 18460 32250 18495
rect 32285 18460 32295 18495
rect 32330 18460 32340 18495
rect 32375 18460 32385 18495
rect 32420 18460 32430 18495
rect 32465 18460 32475 18495
rect 32510 18460 32520 18495
rect 32555 18460 32565 18495
rect 32600 18460 32610 18495
rect 32645 18460 32655 18495
rect 32690 18460 32700 18495
rect 32735 18460 32745 18495
rect 32780 18460 32790 18495
rect 32825 18460 32835 18495
rect 32870 18460 32890 18495
rect 31290 18450 32890 18460
rect 31290 18415 31305 18450
rect 31340 18415 31350 18450
rect 31385 18415 31395 18450
rect 31430 18415 31440 18450
rect 31475 18415 31485 18450
rect 31520 18415 31530 18450
rect 31565 18415 31575 18450
rect 31610 18415 31620 18450
rect 31655 18415 31665 18450
rect 31700 18415 31710 18450
rect 31745 18415 31755 18450
rect 31790 18415 31800 18450
rect 31835 18415 31845 18450
rect 31880 18415 31890 18450
rect 31925 18415 31935 18450
rect 31970 18415 31980 18450
rect 32015 18415 32025 18450
rect 32060 18415 32070 18450
rect 32105 18415 32115 18450
rect 32150 18415 32160 18450
rect 32195 18415 32205 18450
rect 32240 18415 32250 18450
rect 32285 18415 32295 18450
rect 32330 18415 32340 18450
rect 32375 18415 32385 18450
rect 32420 18415 32430 18450
rect 32465 18415 32475 18450
rect 32510 18415 32520 18450
rect 32555 18415 32565 18450
rect 32600 18415 32610 18450
rect 32645 18415 32655 18450
rect 32690 18415 32700 18450
rect 32735 18415 32745 18450
rect 32780 18415 32790 18450
rect 32825 18415 32835 18450
rect 32870 18415 32890 18450
rect 31290 18405 32890 18415
rect 31290 18370 31305 18405
rect 31340 18370 31350 18405
rect 31385 18370 31395 18405
rect 31430 18370 31440 18405
rect 31475 18370 31485 18405
rect 31520 18370 31530 18405
rect 31565 18370 31575 18405
rect 31610 18370 31620 18405
rect 31655 18370 31665 18405
rect 31700 18370 31710 18405
rect 31745 18370 31755 18405
rect 31790 18370 31800 18405
rect 31835 18370 31845 18405
rect 31880 18370 31890 18405
rect 31925 18370 31935 18405
rect 31970 18370 31980 18405
rect 32015 18370 32025 18405
rect 32060 18370 32070 18405
rect 32105 18370 32115 18405
rect 32150 18370 32160 18405
rect 32195 18370 32205 18405
rect 32240 18370 32250 18405
rect 32285 18370 32295 18405
rect 32330 18370 32340 18405
rect 32375 18370 32385 18405
rect 32420 18370 32430 18405
rect 32465 18370 32475 18405
rect 32510 18370 32520 18405
rect 32555 18370 32565 18405
rect 32600 18370 32610 18405
rect 32645 18370 32655 18405
rect 32690 18370 32700 18405
rect 32735 18370 32745 18405
rect 32780 18370 32790 18405
rect 32825 18370 32835 18405
rect 32870 18370 32890 18405
rect 31290 18360 32890 18370
rect 31290 18325 31305 18360
rect 31340 18325 31350 18360
rect 31385 18325 31395 18360
rect 31430 18325 31440 18360
rect 31475 18325 31485 18360
rect 31520 18325 31530 18360
rect 31565 18325 31575 18360
rect 31610 18325 31620 18360
rect 31655 18325 31665 18360
rect 31700 18325 31710 18360
rect 31745 18325 31755 18360
rect 31790 18325 31800 18360
rect 31835 18325 31845 18360
rect 31880 18325 31890 18360
rect 31925 18325 31935 18360
rect 31970 18325 31980 18360
rect 32015 18325 32025 18360
rect 32060 18325 32070 18360
rect 32105 18325 32115 18360
rect 32150 18325 32160 18360
rect 32195 18325 32205 18360
rect 32240 18325 32250 18360
rect 32285 18325 32295 18360
rect 32330 18325 32340 18360
rect 32375 18325 32385 18360
rect 32420 18325 32430 18360
rect 32465 18325 32475 18360
rect 32510 18325 32520 18360
rect 32555 18325 32565 18360
rect 32600 18325 32610 18360
rect 32645 18325 32655 18360
rect 32690 18325 32700 18360
rect 32735 18325 32745 18360
rect 32780 18325 32790 18360
rect 32825 18325 32835 18360
rect 32870 18325 32890 18360
rect 31290 18315 32890 18325
rect 31290 18280 31305 18315
rect 31340 18280 31350 18315
rect 31385 18280 31395 18315
rect 31430 18280 31440 18315
rect 31475 18280 31485 18315
rect 31520 18280 31530 18315
rect 31565 18280 31575 18315
rect 31610 18280 31620 18315
rect 31655 18280 31665 18315
rect 31700 18280 31710 18315
rect 31745 18280 31755 18315
rect 31790 18280 31800 18315
rect 31835 18280 31845 18315
rect 31880 18280 31890 18315
rect 31925 18280 31935 18315
rect 31970 18280 31980 18315
rect 32015 18280 32025 18315
rect 32060 18280 32070 18315
rect 32105 18280 32115 18315
rect 32150 18280 32160 18315
rect 32195 18280 32205 18315
rect 32240 18280 32250 18315
rect 32285 18280 32295 18315
rect 32330 18280 32340 18315
rect 32375 18280 32385 18315
rect 32420 18280 32430 18315
rect 32465 18280 32475 18315
rect 32510 18280 32520 18315
rect 32555 18280 32565 18315
rect 32600 18280 32610 18315
rect 32645 18280 32655 18315
rect 32690 18280 32700 18315
rect 32735 18280 32745 18315
rect 32780 18280 32790 18315
rect 32825 18280 32835 18315
rect 32870 18280 32890 18315
rect 31290 18270 32890 18280
rect 31290 18235 31305 18270
rect 31340 18235 31350 18270
rect 31385 18235 31395 18270
rect 31430 18235 31440 18270
rect 31475 18235 31485 18270
rect 31520 18235 31530 18270
rect 31565 18235 31575 18270
rect 31610 18235 31620 18270
rect 31655 18235 31665 18270
rect 31700 18235 31710 18270
rect 31745 18235 31755 18270
rect 31790 18235 31800 18270
rect 31835 18235 31845 18270
rect 31880 18235 31890 18270
rect 31925 18235 31935 18270
rect 31970 18235 31980 18270
rect 32015 18235 32025 18270
rect 32060 18235 32070 18270
rect 32105 18235 32115 18270
rect 32150 18235 32160 18270
rect 32195 18235 32205 18270
rect 32240 18235 32250 18270
rect 32285 18235 32295 18270
rect 32330 18235 32340 18270
rect 32375 18235 32385 18270
rect 32420 18235 32430 18270
rect 32465 18235 32475 18270
rect 32510 18235 32520 18270
rect 32555 18235 32565 18270
rect 32600 18235 32610 18270
rect 32645 18235 32655 18270
rect 32690 18235 32700 18270
rect 32735 18235 32745 18270
rect 32780 18235 32790 18270
rect 32825 18235 32835 18270
rect 32870 18235 32890 18270
rect 31290 18225 32890 18235
rect 31290 18190 31305 18225
rect 31340 18190 31350 18225
rect 31385 18190 31395 18225
rect 31430 18190 31440 18225
rect 31475 18190 31485 18225
rect 31520 18190 31530 18225
rect 31565 18190 31575 18225
rect 31610 18190 31620 18225
rect 31655 18190 31665 18225
rect 31700 18190 31710 18225
rect 31745 18190 31755 18225
rect 31790 18190 31800 18225
rect 31835 18190 31845 18225
rect 31880 18190 31890 18225
rect 31925 18190 31935 18225
rect 31970 18190 31980 18225
rect 32015 18190 32025 18225
rect 32060 18190 32070 18225
rect 32105 18190 32115 18225
rect 32150 18190 32160 18225
rect 32195 18190 32205 18225
rect 32240 18190 32250 18225
rect 32285 18190 32295 18225
rect 32330 18190 32340 18225
rect 32375 18190 32385 18225
rect 32420 18190 32430 18225
rect 32465 18190 32475 18225
rect 32510 18190 32520 18225
rect 32555 18190 32565 18225
rect 32600 18190 32610 18225
rect 32645 18190 32655 18225
rect 32690 18190 32700 18225
rect 32735 18190 32745 18225
rect 32780 18190 32790 18225
rect 32825 18190 32835 18225
rect 32870 18190 32890 18225
rect 31290 18180 32890 18190
rect 31290 18145 31305 18180
rect 31340 18145 31350 18180
rect 31385 18145 31395 18180
rect 31430 18145 31440 18180
rect 31475 18145 31485 18180
rect 31520 18145 31530 18180
rect 31565 18145 31575 18180
rect 31610 18145 31620 18180
rect 31655 18145 31665 18180
rect 31700 18145 31710 18180
rect 31745 18145 31755 18180
rect 31790 18145 31800 18180
rect 31835 18145 31845 18180
rect 31880 18145 31890 18180
rect 31925 18145 31935 18180
rect 31970 18145 31980 18180
rect 32015 18145 32025 18180
rect 32060 18145 32070 18180
rect 32105 18145 32115 18180
rect 32150 18145 32160 18180
rect 32195 18145 32205 18180
rect 32240 18145 32250 18180
rect 32285 18145 32295 18180
rect 32330 18145 32340 18180
rect 32375 18145 32385 18180
rect 32420 18145 32430 18180
rect 32465 18145 32475 18180
rect 32510 18145 32520 18180
rect 32555 18145 32565 18180
rect 32600 18145 32610 18180
rect 32645 18145 32655 18180
rect 32690 18145 32700 18180
rect 32735 18145 32745 18180
rect 32780 18145 32790 18180
rect 32825 18145 32835 18180
rect 32870 18145 32890 18180
rect 31290 18135 32890 18145
rect 31290 18100 31305 18135
rect 31340 18100 31350 18135
rect 31385 18100 31395 18135
rect 31430 18100 31440 18135
rect 31475 18100 31485 18135
rect 31520 18100 31530 18135
rect 31565 18100 31575 18135
rect 31610 18100 31620 18135
rect 31655 18100 31665 18135
rect 31700 18100 31710 18135
rect 31745 18100 31755 18135
rect 31790 18100 31800 18135
rect 31835 18100 31845 18135
rect 31880 18100 31890 18135
rect 31925 18100 31935 18135
rect 31970 18100 31980 18135
rect 32015 18100 32025 18135
rect 32060 18100 32070 18135
rect 32105 18100 32115 18135
rect 32150 18100 32160 18135
rect 32195 18100 32205 18135
rect 32240 18100 32250 18135
rect 32285 18100 32295 18135
rect 32330 18100 32340 18135
rect 32375 18100 32385 18135
rect 32420 18100 32430 18135
rect 32465 18100 32475 18135
rect 32510 18100 32520 18135
rect 32555 18100 32565 18135
rect 32600 18100 32610 18135
rect 32645 18100 32655 18135
rect 32690 18100 32700 18135
rect 32735 18100 32745 18135
rect 32780 18100 32790 18135
rect 32825 18100 32835 18135
rect 32870 18100 32890 18135
rect 31290 18090 32890 18100
rect 31290 18055 31305 18090
rect 31340 18055 31350 18090
rect 31385 18055 31395 18090
rect 31430 18055 31440 18090
rect 31475 18055 31485 18090
rect 31520 18055 31530 18090
rect 31565 18055 31575 18090
rect 31610 18055 31620 18090
rect 31655 18055 31665 18090
rect 31700 18055 31710 18090
rect 31745 18055 31755 18090
rect 31790 18055 31800 18090
rect 31835 18055 31845 18090
rect 31880 18055 31890 18090
rect 31925 18055 31935 18090
rect 31970 18055 31980 18090
rect 32015 18055 32025 18090
rect 32060 18055 32070 18090
rect 32105 18055 32115 18090
rect 32150 18055 32160 18090
rect 32195 18055 32205 18090
rect 32240 18055 32250 18090
rect 32285 18055 32295 18090
rect 32330 18055 32340 18090
rect 32375 18055 32385 18090
rect 32420 18055 32430 18090
rect 32465 18055 32475 18090
rect 32510 18055 32520 18090
rect 32555 18055 32565 18090
rect 32600 18055 32610 18090
rect 32645 18055 32655 18090
rect 32690 18055 32700 18090
rect 32735 18055 32745 18090
rect 32780 18055 32790 18090
rect 32825 18055 32835 18090
rect 32870 18055 32890 18090
rect 31290 18045 32890 18055
rect 31290 18010 31305 18045
rect 31340 18010 31350 18045
rect 31385 18010 31395 18045
rect 31430 18010 31440 18045
rect 31475 18010 31485 18045
rect 31520 18010 31530 18045
rect 31565 18010 31575 18045
rect 31610 18010 31620 18045
rect 31655 18010 31665 18045
rect 31700 18010 31710 18045
rect 31745 18010 31755 18045
rect 31790 18010 31800 18045
rect 31835 18010 31845 18045
rect 31880 18010 31890 18045
rect 31925 18010 31935 18045
rect 31970 18010 31980 18045
rect 32015 18010 32025 18045
rect 32060 18010 32070 18045
rect 32105 18010 32115 18045
rect 32150 18010 32160 18045
rect 32195 18010 32205 18045
rect 32240 18010 32250 18045
rect 32285 18010 32295 18045
rect 32330 18010 32340 18045
rect 32375 18010 32385 18045
rect 32420 18010 32430 18045
rect 32465 18010 32475 18045
rect 32510 18010 32520 18045
rect 32555 18010 32565 18045
rect 32600 18010 32610 18045
rect 32645 18010 32655 18045
rect 32690 18010 32700 18045
rect 32735 18010 32745 18045
rect 32780 18010 32790 18045
rect 32825 18010 32835 18045
rect 32870 18010 32890 18045
rect 31290 18000 32890 18010
rect 31290 17965 31305 18000
rect 31340 17965 31350 18000
rect 31385 17965 31395 18000
rect 31430 17965 31440 18000
rect 31475 17965 31485 18000
rect 31520 17965 31530 18000
rect 31565 17965 31575 18000
rect 31610 17965 31620 18000
rect 31655 17965 31665 18000
rect 31700 17965 31710 18000
rect 31745 17965 31755 18000
rect 31790 17965 31800 18000
rect 31835 17965 31845 18000
rect 31880 17965 31890 18000
rect 31925 17965 31935 18000
rect 31970 17965 31980 18000
rect 32015 17965 32025 18000
rect 32060 17965 32070 18000
rect 32105 17965 32115 18000
rect 32150 17965 32160 18000
rect 32195 17965 32205 18000
rect 32240 17965 32250 18000
rect 32285 17965 32295 18000
rect 32330 17965 32340 18000
rect 32375 17965 32385 18000
rect 32420 17965 32430 18000
rect 32465 17965 32475 18000
rect 32510 17965 32520 18000
rect 32555 17965 32565 18000
rect 32600 17965 32610 18000
rect 32645 17965 32655 18000
rect 32690 17965 32700 18000
rect 32735 17965 32745 18000
rect 32780 17965 32790 18000
rect 32825 17965 32835 18000
rect 32870 17965 32890 18000
rect 31290 17955 32890 17965
rect 31290 17920 31305 17955
rect 31340 17920 31350 17955
rect 31385 17920 31395 17955
rect 31430 17920 31440 17955
rect 31475 17920 31485 17955
rect 31520 17920 31530 17955
rect 31565 17920 31575 17955
rect 31610 17920 31620 17955
rect 31655 17920 31665 17955
rect 31700 17920 31710 17955
rect 31745 17920 31755 17955
rect 31790 17920 31800 17955
rect 31835 17920 31845 17955
rect 31880 17920 31890 17955
rect 31925 17920 31935 17955
rect 31970 17920 31980 17955
rect 32015 17920 32025 17955
rect 32060 17920 32070 17955
rect 32105 17920 32115 17955
rect 32150 17920 32160 17955
rect 32195 17920 32205 17955
rect 32240 17920 32250 17955
rect 32285 17920 32295 17955
rect 32330 17920 32340 17955
rect 32375 17920 32385 17955
rect 32420 17920 32430 17955
rect 32465 17920 32475 17955
rect 32510 17920 32520 17955
rect 32555 17920 32565 17955
rect 32600 17920 32610 17955
rect 32645 17920 32655 17955
rect 32690 17920 32700 17955
rect 32735 17920 32745 17955
rect 32780 17920 32790 17955
rect 32825 17920 32835 17955
rect 32870 17920 32890 17955
rect 31290 17910 32890 17920
rect 31290 17875 31305 17910
rect 31340 17875 31350 17910
rect 31385 17875 31395 17910
rect 31430 17875 31440 17910
rect 31475 17875 31485 17910
rect 31520 17875 31530 17910
rect 31565 17875 31575 17910
rect 31610 17875 31620 17910
rect 31655 17875 31665 17910
rect 31700 17875 31710 17910
rect 31745 17875 31755 17910
rect 31790 17875 31800 17910
rect 31835 17875 31845 17910
rect 31880 17875 31890 17910
rect 31925 17875 31935 17910
rect 31970 17875 31980 17910
rect 32015 17875 32025 17910
rect 32060 17875 32070 17910
rect 32105 17875 32115 17910
rect 32150 17875 32160 17910
rect 32195 17875 32205 17910
rect 32240 17875 32250 17910
rect 32285 17875 32295 17910
rect 32330 17875 32340 17910
rect 32375 17875 32385 17910
rect 32420 17875 32430 17910
rect 32465 17875 32475 17910
rect 32510 17875 32520 17910
rect 32555 17875 32565 17910
rect 32600 17875 32610 17910
rect 32645 17875 32655 17910
rect 32690 17875 32700 17910
rect 32735 17875 32745 17910
rect 32780 17875 32790 17910
rect 32825 17875 32835 17910
rect 32870 17875 32890 17910
rect 31290 17865 32890 17875
rect 31290 17830 31305 17865
rect 31340 17830 31350 17865
rect 31385 17830 31395 17865
rect 31430 17830 31440 17865
rect 31475 17830 31485 17865
rect 31520 17830 31530 17865
rect 31565 17830 31575 17865
rect 31610 17830 31620 17865
rect 31655 17830 31665 17865
rect 31700 17830 31710 17865
rect 31745 17830 31755 17865
rect 31790 17830 31800 17865
rect 31835 17830 31845 17865
rect 31880 17830 31890 17865
rect 31925 17830 31935 17865
rect 31970 17830 31980 17865
rect 32015 17830 32025 17865
rect 32060 17830 32070 17865
rect 32105 17830 32115 17865
rect 32150 17830 32160 17865
rect 32195 17830 32205 17865
rect 32240 17830 32250 17865
rect 32285 17830 32295 17865
rect 32330 17830 32340 17865
rect 32375 17830 32385 17865
rect 32420 17830 32430 17865
rect 32465 17830 32475 17865
rect 32510 17830 32520 17865
rect 32555 17830 32565 17865
rect 32600 17830 32610 17865
rect 32645 17830 32655 17865
rect 32690 17830 32700 17865
rect 32735 17830 32745 17865
rect 32780 17830 32790 17865
rect 32825 17830 32835 17865
rect 32870 17830 32890 17865
rect 31290 17820 32890 17830
rect 31290 17785 31305 17820
rect 31340 17785 31350 17820
rect 31385 17785 31395 17820
rect 31430 17785 31440 17820
rect 31475 17785 31485 17820
rect 31520 17785 31530 17820
rect 31565 17785 31575 17820
rect 31610 17785 31620 17820
rect 31655 17785 31665 17820
rect 31700 17785 31710 17820
rect 31745 17785 31755 17820
rect 31790 17785 31800 17820
rect 31835 17785 31845 17820
rect 31880 17785 31890 17820
rect 31925 17785 31935 17820
rect 31970 17785 31980 17820
rect 32015 17785 32025 17820
rect 32060 17785 32070 17820
rect 32105 17785 32115 17820
rect 32150 17785 32160 17820
rect 32195 17785 32205 17820
rect 32240 17785 32250 17820
rect 32285 17785 32295 17820
rect 32330 17785 32340 17820
rect 32375 17785 32385 17820
rect 32420 17785 32430 17820
rect 32465 17785 32475 17820
rect 32510 17785 32520 17820
rect 32555 17785 32565 17820
rect 32600 17785 32610 17820
rect 32645 17785 32655 17820
rect 32690 17785 32700 17820
rect 32735 17785 32745 17820
rect 32780 17785 32790 17820
rect 32825 17785 32835 17820
rect 32870 17785 32890 17820
rect 31290 17775 32890 17785
rect 31290 17740 31305 17775
rect 31340 17740 31350 17775
rect 31385 17740 31395 17775
rect 31430 17740 31440 17775
rect 31475 17740 31485 17775
rect 31520 17740 31530 17775
rect 31565 17740 31575 17775
rect 31610 17740 31620 17775
rect 31655 17740 31665 17775
rect 31700 17740 31710 17775
rect 31745 17740 31755 17775
rect 31790 17740 31800 17775
rect 31835 17740 31845 17775
rect 31880 17740 31890 17775
rect 31925 17740 31935 17775
rect 31970 17740 31980 17775
rect 32015 17740 32025 17775
rect 32060 17740 32070 17775
rect 32105 17740 32115 17775
rect 32150 17740 32160 17775
rect 32195 17740 32205 17775
rect 32240 17740 32250 17775
rect 32285 17740 32295 17775
rect 32330 17740 32340 17775
rect 32375 17740 32385 17775
rect 32420 17740 32430 17775
rect 32465 17740 32475 17775
rect 32510 17740 32520 17775
rect 32555 17740 32565 17775
rect 32600 17740 32610 17775
rect 32645 17740 32655 17775
rect 32690 17740 32700 17775
rect 32735 17740 32745 17775
rect 32780 17740 32790 17775
rect 32825 17740 32835 17775
rect 32870 17740 32890 17775
rect 31290 10530 32890 17740
rect 31290 10495 31305 10530
rect 31340 10495 31350 10530
rect 31385 10495 31395 10530
rect 31430 10495 31440 10530
rect 31475 10495 31485 10530
rect 31520 10495 31530 10530
rect 31565 10495 31575 10530
rect 31610 10495 31620 10530
rect 31655 10495 31665 10530
rect 31700 10495 31710 10530
rect 31745 10495 31755 10530
rect 31790 10495 31800 10530
rect 31835 10495 31845 10530
rect 31880 10495 31890 10530
rect 31925 10495 31935 10530
rect 31970 10495 31980 10530
rect 32015 10495 32025 10530
rect 32060 10495 32070 10530
rect 32105 10495 32115 10530
rect 32150 10495 32160 10530
rect 32195 10495 32205 10530
rect 32240 10495 32250 10530
rect 32285 10495 32295 10530
rect 32330 10495 32340 10530
rect 32375 10495 32385 10530
rect 32420 10495 32430 10530
rect 32465 10495 32475 10530
rect 32510 10495 32520 10530
rect 32555 10495 32565 10530
rect 32600 10495 32610 10530
rect 32645 10495 32655 10530
rect 32690 10495 32700 10530
rect 32735 10495 32745 10530
rect 32780 10495 32790 10530
rect 32825 10495 32835 10530
rect 32870 10495 32890 10530
rect 31290 10485 32890 10495
rect 31290 10450 31305 10485
rect 31340 10450 31350 10485
rect 31385 10450 31395 10485
rect 31430 10450 31440 10485
rect 31475 10450 31485 10485
rect 31520 10450 31530 10485
rect 31565 10450 31575 10485
rect 31610 10450 31620 10485
rect 31655 10450 31665 10485
rect 31700 10450 31710 10485
rect 31745 10450 31755 10485
rect 31790 10450 31800 10485
rect 31835 10450 31845 10485
rect 31880 10450 31890 10485
rect 31925 10450 31935 10485
rect 31970 10450 31980 10485
rect 32015 10450 32025 10485
rect 32060 10450 32070 10485
rect 32105 10450 32115 10485
rect 32150 10450 32160 10485
rect 32195 10450 32205 10485
rect 32240 10450 32250 10485
rect 32285 10450 32295 10485
rect 32330 10450 32340 10485
rect 32375 10450 32385 10485
rect 32420 10450 32430 10485
rect 32465 10450 32475 10485
rect 32510 10450 32520 10485
rect 32555 10450 32565 10485
rect 32600 10450 32610 10485
rect 32645 10450 32655 10485
rect 32690 10450 32700 10485
rect 32735 10450 32745 10485
rect 32780 10450 32790 10485
rect 32825 10450 32835 10485
rect 32870 10450 32890 10485
rect 31290 10440 32890 10450
rect 31290 10405 31305 10440
rect 31340 10405 31350 10440
rect 31385 10405 31395 10440
rect 31430 10405 31440 10440
rect 31475 10405 31485 10440
rect 31520 10405 31530 10440
rect 31565 10405 31575 10440
rect 31610 10405 31620 10440
rect 31655 10405 31665 10440
rect 31700 10405 31710 10440
rect 31745 10405 31755 10440
rect 31790 10405 31800 10440
rect 31835 10405 31845 10440
rect 31880 10405 31890 10440
rect 31925 10405 31935 10440
rect 31970 10405 31980 10440
rect 32015 10405 32025 10440
rect 32060 10405 32070 10440
rect 32105 10405 32115 10440
rect 32150 10405 32160 10440
rect 32195 10405 32205 10440
rect 32240 10405 32250 10440
rect 32285 10405 32295 10440
rect 32330 10405 32340 10440
rect 32375 10405 32385 10440
rect 32420 10405 32430 10440
rect 32465 10405 32475 10440
rect 32510 10405 32520 10440
rect 32555 10405 32565 10440
rect 32600 10405 32610 10440
rect 32645 10405 32655 10440
rect 32690 10405 32700 10440
rect 32735 10405 32745 10440
rect 32780 10405 32790 10440
rect 32825 10405 32835 10440
rect 32870 10405 32890 10440
rect 31290 10395 32890 10405
rect 31290 10360 31305 10395
rect 31340 10360 31350 10395
rect 31385 10360 31395 10395
rect 31430 10360 31440 10395
rect 31475 10360 31485 10395
rect 31520 10360 31530 10395
rect 31565 10360 31575 10395
rect 31610 10360 31620 10395
rect 31655 10360 31665 10395
rect 31700 10360 31710 10395
rect 31745 10360 31755 10395
rect 31790 10360 31800 10395
rect 31835 10360 31845 10395
rect 31880 10360 31890 10395
rect 31925 10360 31935 10395
rect 31970 10360 31980 10395
rect 32015 10360 32025 10395
rect 32060 10360 32070 10395
rect 32105 10360 32115 10395
rect 32150 10360 32160 10395
rect 32195 10360 32205 10395
rect 32240 10360 32250 10395
rect 32285 10360 32295 10395
rect 32330 10360 32340 10395
rect 32375 10360 32385 10395
rect 32420 10360 32430 10395
rect 32465 10360 32475 10395
rect 32510 10360 32520 10395
rect 32555 10360 32565 10395
rect 32600 10360 32610 10395
rect 32645 10360 32655 10395
rect 32690 10360 32700 10395
rect 32735 10360 32745 10395
rect 32780 10360 32790 10395
rect 32825 10360 32835 10395
rect 32870 10360 32890 10395
rect 31290 10350 32890 10360
rect 31290 10315 31305 10350
rect 31340 10315 31350 10350
rect 31385 10315 31395 10350
rect 31430 10315 31440 10350
rect 31475 10315 31485 10350
rect 31520 10315 31530 10350
rect 31565 10315 31575 10350
rect 31610 10315 31620 10350
rect 31655 10315 31665 10350
rect 31700 10315 31710 10350
rect 31745 10315 31755 10350
rect 31790 10315 31800 10350
rect 31835 10315 31845 10350
rect 31880 10315 31890 10350
rect 31925 10315 31935 10350
rect 31970 10315 31980 10350
rect 32015 10315 32025 10350
rect 32060 10315 32070 10350
rect 32105 10315 32115 10350
rect 32150 10315 32160 10350
rect 32195 10315 32205 10350
rect 32240 10315 32250 10350
rect 32285 10315 32295 10350
rect 32330 10315 32340 10350
rect 32375 10315 32385 10350
rect 32420 10315 32430 10350
rect 32465 10315 32475 10350
rect 32510 10315 32520 10350
rect 32555 10315 32565 10350
rect 32600 10315 32610 10350
rect 32645 10315 32655 10350
rect 32690 10315 32700 10350
rect 32735 10315 32745 10350
rect 32780 10315 32790 10350
rect 32825 10315 32835 10350
rect 32870 10315 32890 10350
rect 31290 10305 32890 10315
rect 31290 10270 31305 10305
rect 31340 10270 31350 10305
rect 31385 10270 31395 10305
rect 31430 10270 31440 10305
rect 31475 10270 31485 10305
rect 31520 10270 31530 10305
rect 31565 10270 31575 10305
rect 31610 10270 31620 10305
rect 31655 10270 31665 10305
rect 31700 10270 31710 10305
rect 31745 10270 31755 10305
rect 31790 10270 31800 10305
rect 31835 10270 31845 10305
rect 31880 10270 31890 10305
rect 31925 10270 31935 10305
rect 31970 10270 31980 10305
rect 32015 10270 32025 10305
rect 32060 10270 32070 10305
rect 32105 10270 32115 10305
rect 32150 10270 32160 10305
rect 32195 10270 32205 10305
rect 32240 10270 32250 10305
rect 32285 10270 32295 10305
rect 32330 10270 32340 10305
rect 32375 10270 32385 10305
rect 32420 10270 32430 10305
rect 32465 10270 32475 10305
rect 32510 10270 32520 10305
rect 32555 10270 32565 10305
rect 32600 10270 32610 10305
rect 32645 10270 32655 10305
rect 32690 10270 32700 10305
rect 32735 10270 32745 10305
rect 32780 10270 32790 10305
rect 32825 10270 32835 10305
rect 32870 10270 32890 10305
rect 31290 10260 32890 10270
rect 31290 10225 31305 10260
rect 31340 10225 31350 10260
rect 31385 10225 31395 10260
rect 31430 10225 31440 10260
rect 31475 10225 31485 10260
rect 31520 10225 31530 10260
rect 31565 10225 31575 10260
rect 31610 10225 31620 10260
rect 31655 10225 31665 10260
rect 31700 10225 31710 10260
rect 31745 10225 31755 10260
rect 31790 10225 31800 10260
rect 31835 10225 31845 10260
rect 31880 10225 31890 10260
rect 31925 10225 31935 10260
rect 31970 10225 31980 10260
rect 32015 10225 32025 10260
rect 32060 10225 32070 10260
rect 32105 10225 32115 10260
rect 32150 10225 32160 10260
rect 32195 10225 32205 10260
rect 32240 10225 32250 10260
rect 32285 10225 32295 10260
rect 32330 10225 32340 10260
rect 32375 10225 32385 10260
rect 32420 10225 32430 10260
rect 32465 10225 32475 10260
rect 32510 10225 32520 10260
rect 32555 10225 32565 10260
rect 32600 10225 32610 10260
rect 32645 10225 32655 10260
rect 32690 10225 32700 10260
rect 32735 10225 32745 10260
rect 32780 10225 32790 10260
rect 32825 10225 32835 10260
rect 32870 10225 32890 10260
rect 31290 10215 32890 10225
rect 31290 10180 31305 10215
rect 31340 10180 31350 10215
rect 31385 10180 31395 10215
rect 31430 10180 31440 10215
rect 31475 10180 31485 10215
rect 31520 10180 31530 10215
rect 31565 10180 31575 10215
rect 31610 10180 31620 10215
rect 31655 10180 31665 10215
rect 31700 10180 31710 10215
rect 31745 10180 31755 10215
rect 31790 10180 31800 10215
rect 31835 10180 31845 10215
rect 31880 10180 31890 10215
rect 31925 10180 31935 10215
rect 31970 10180 31980 10215
rect 32015 10180 32025 10215
rect 32060 10180 32070 10215
rect 32105 10180 32115 10215
rect 32150 10180 32160 10215
rect 32195 10180 32205 10215
rect 32240 10180 32250 10215
rect 32285 10180 32295 10215
rect 32330 10180 32340 10215
rect 32375 10180 32385 10215
rect 32420 10180 32430 10215
rect 32465 10180 32475 10215
rect 32510 10180 32520 10215
rect 32555 10180 32565 10215
rect 32600 10180 32610 10215
rect 32645 10180 32655 10215
rect 32690 10180 32700 10215
rect 32735 10180 32745 10215
rect 32780 10180 32790 10215
rect 32825 10180 32835 10215
rect 32870 10180 32890 10215
rect 31290 10170 32890 10180
rect -38770 9630 -37170 10155
rect 31290 10135 31305 10170
rect 31340 10135 31350 10170
rect 31385 10135 31395 10170
rect 31430 10135 31440 10170
rect 31475 10135 31485 10170
rect 31520 10135 31530 10170
rect 31565 10135 31575 10170
rect 31610 10135 31620 10170
rect 31655 10135 31665 10170
rect 31700 10135 31710 10170
rect 31745 10135 31755 10170
rect 31790 10135 31800 10170
rect 31835 10135 31845 10170
rect 31880 10135 31890 10170
rect 31925 10135 31935 10170
rect 31970 10135 31980 10170
rect 32015 10135 32025 10170
rect 32060 10135 32070 10170
rect 32105 10135 32115 10170
rect 32150 10135 32160 10170
rect 32195 10135 32205 10170
rect 32240 10135 32250 10170
rect 32285 10135 32295 10170
rect 32330 10135 32340 10170
rect 32375 10135 32385 10170
rect 32420 10135 32430 10170
rect 32465 10135 32475 10170
rect 32510 10135 32520 10170
rect 32555 10135 32565 10170
rect 32600 10135 32610 10170
rect 32645 10135 32655 10170
rect 32690 10135 32700 10170
rect 32735 10135 32745 10170
rect 32780 10135 32790 10170
rect 32825 10135 32835 10170
rect 32870 10135 32890 10170
rect 31290 10125 32890 10135
rect 31290 10090 31305 10125
rect 31340 10090 31350 10125
rect 31385 10090 31395 10125
rect 31430 10090 31440 10125
rect 31475 10090 31485 10125
rect 31520 10090 31530 10125
rect 31565 10090 31575 10125
rect 31610 10090 31620 10125
rect 31655 10090 31665 10125
rect 31700 10090 31710 10125
rect 31745 10090 31755 10125
rect 31790 10090 31800 10125
rect 31835 10090 31845 10125
rect 31880 10090 31890 10125
rect 31925 10090 31935 10125
rect 31970 10090 31980 10125
rect 32015 10090 32025 10125
rect 32060 10090 32070 10125
rect 32105 10090 32115 10125
rect 32150 10090 32160 10125
rect 32195 10090 32205 10125
rect 32240 10090 32250 10125
rect 32285 10090 32295 10125
rect 32330 10090 32340 10125
rect 32375 10090 32385 10125
rect 32420 10090 32430 10125
rect 32465 10090 32475 10125
rect 32510 10090 32520 10125
rect 32555 10090 32565 10125
rect 32600 10090 32610 10125
rect 32645 10090 32655 10125
rect 32690 10090 32700 10125
rect 32735 10090 32745 10125
rect 32780 10090 32790 10125
rect 32825 10090 32835 10125
rect 32870 10090 32890 10125
rect 31290 10080 32890 10090
rect 31290 10045 31305 10080
rect 31340 10045 31350 10080
rect 31385 10045 31395 10080
rect 31430 10045 31440 10080
rect 31475 10045 31485 10080
rect 31520 10045 31530 10080
rect 31565 10045 31575 10080
rect 31610 10045 31620 10080
rect 31655 10045 31665 10080
rect 31700 10045 31710 10080
rect 31745 10045 31755 10080
rect 31790 10045 31800 10080
rect 31835 10045 31845 10080
rect 31880 10045 31890 10080
rect 31925 10045 31935 10080
rect 31970 10045 31980 10080
rect 32015 10045 32025 10080
rect 32060 10045 32070 10080
rect 32105 10045 32115 10080
rect 32150 10045 32160 10080
rect 32195 10045 32205 10080
rect 32240 10045 32250 10080
rect 32285 10045 32295 10080
rect 32330 10045 32340 10080
rect 32375 10045 32385 10080
rect 32420 10045 32430 10080
rect 32465 10045 32475 10080
rect 32510 10045 32520 10080
rect 32555 10045 32565 10080
rect 32600 10045 32610 10080
rect 32645 10045 32655 10080
rect 32690 10045 32700 10080
rect 32735 10045 32745 10080
rect 32780 10045 32790 10080
rect 32825 10045 32835 10080
rect 32870 10045 32890 10080
rect 31290 10035 32890 10045
rect 31290 10000 31305 10035
rect 31340 10000 31350 10035
rect 31385 10000 31395 10035
rect 31430 10000 31440 10035
rect 31475 10000 31485 10035
rect 31520 10000 31530 10035
rect 31565 10000 31575 10035
rect 31610 10000 31620 10035
rect 31655 10000 31665 10035
rect 31700 10000 31710 10035
rect 31745 10000 31755 10035
rect 31790 10000 31800 10035
rect 31835 10000 31845 10035
rect 31880 10000 31890 10035
rect 31925 10000 31935 10035
rect 31970 10000 31980 10035
rect 32015 10000 32025 10035
rect 32060 10000 32070 10035
rect 32105 10000 32115 10035
rect 32150 10000 32160 10035
rect 32195 10000 32205 10035
rect 32240 10000 32250 10035
rect 32285 10000 32295 10035
rect 32330 10000 32340 10035
rect 32375 10000 32385 10035
rect 32420 10000 32430 10035
rect 32465 10000 32475 10035
rect 32510 10000 32520 10035
rect 32555 10000 32565 10035
rect 32600 10000 32610 10035
rect 32645 10000 32655 10035
rect 32690 10000 32700 10035
rect 32735 10000 32745 10035
rect 32780 10000 32790 10035
rect 32825 10000 32835 10035
rect 32870 10000 32890 10035
rect 31290 9990 32890 10000
rect 31290 9955 31305 9990
rect 31340 9955 31350 9990
rect 31385 9955 31395 9990
rect 31430 9955 31440 9990
rect 31475 9955 31485 9990
rect 31520 9955 31530 9990
rect 31565 9955 31575 9990
rect 31610 9955 31620 9990
rect 31655 9955 31665 9990
rect 31700 9955 31710 9990
rect 31745 9955 31755 9990
rect 31790 9955 31800 9990
rect 31835 9955 31845 9990
rect 31880 9955 31890 9990
rect 31925 9955 31935 9990
rect 31970 9955 31980 9990
rect 32015 9955 32025 9990
rect 32060 9955 32070 9990
rect 32105 9955 32115 9990
rect 32150 9955 32160 9990
rect 32195 9955 32205 9990
rect 32240 9955 32250 9990
rect 32285 9955 32295 9990
rect 32330 9955 32340 9990
rect 32375 9955 32385 9990
rect 32420 9955 32430 9990
rect 32465 9955 32475 9990
rect 32510 9955 32520 9990
rect 32555 9955 32565 9990
rect 32600 9955 32610 9990
rect 32645 9955 32655 9990
rect 32690 9955 32700 9990
rect 32735 9955 32745 9990
rect 32780 9955 32790 9990
rect 32825 9955 32835 9990
rect 32870 9955 32890 9990
rect 31290 9945 32890 9955
rect 31290 9910 31305 9945
rect 31340 9910 31350 9945
rect 31385 9910 31395 9945
rect 31430 9910 31440 9945
rect 31475 9910 31485 9945
rect 31520 9910 31530 9945
rect 31565 9910 31575 9945
rect 31610 9910 31620 9945
rect 31655 9910 31665 9945
rect 31700 9910 31710 9945
rect 31745 9910 31755 9945
rect 31790 9910 31800 9945
rect 31835 9910 31845 9945
rect 31880 9910 31890 9945
rect 31925 9910 31935 9945
rect 31970 9910 31980 9945
rect 32015 9910 32025 9945
rect 32060 9910 32070 9945
rect 32105 9910 32115 9945
rect 32150 9910 32160 9945
rect 32195 9910 32205 9945
rect 32240 9910 32250 9945
rect 32285 9910 32295 9945
rect 32330 9910 32340 9945
rect 32375 9910 32385 9945
rect 32420 9910 32430 9945
rect 32465 9910 32475 9945
rect 32510 9910 32520 9945
rect 32555 9910 32565 9945
rect 32600 9910 32610 9945
rect 32645 9910 32655 9945
rect 32690 9910 32700 9945
rect 32735 9910 32745 9945
rect 32780 9910 32790 9945
rect 32825 9910 32835 9945
rect 32870 9910 32890 9945
rect 31290 9900 32890 9910
rect 31290 9865 31305 9900
rect 31340 9865 31350 9900
rect 31385 9865 31395 9900
rect 31430 9865 31440 9900
rect 31475 9865 31485 9900
rect 31520 9865 31530 9900
rect 31565 9865 31575 9900
rect 31610 9865 31620 9900
rect 31655 9865 31665 9900
rect 31700 9865 31710 9900
rect 31745 9865 31755 9900
rect 31790 9865 31800 9900
rect 31835 9865 31845 9900
rect 31880 9865 31890 9900
rect 31925 9865 31935 9900
rect 31970 9865 31980 9900
rect 32015 9865 32025 9900
rect 32060 9865 32070 9900
rect 32105 9865 32115 9900
rect 32150 9865 32160 9900
rect 32195 9865 32205 9900
rect 32240 9865 32250 9900
rect 32285 9865 32295 9900
rect 32330 9865 32340 9900
rect 32375 9865 32385 9900
rect 32420 9865 32430 9900
rect 32465 9865 32475 9900
rect 32510 9865 32520 9900
rect 32555 9865 32565 9900
rect 32600 9865 32610 9900
rect 32645 9865 32655 9900
rect 32690 9865 32700 9900
rect 32735 9865 32745 9900
rect 32780 9865 32790 9900
rect 32825 9865 32835 9900
rect 32870 9865 32890 9900
rect 31290 9855 32890 9865
rect 31290 9820 31305 9855
rect 31340 9820 31350 9855
rect 31385 9820 31395 9855
rect 31430 9820 31440 9855
rect 31475 9820 31485 9855
rect 31520 9820 31530 9855
rect 31565 9820 31575 9855
rect 31610 9820 31620 9855
rect 31655 9820 31665 9855
rect 31700 9820 31710 9855
rect 31745 9820 31755 9855
rect 31790 9820 31800 9855
rect 31835 9820 31845 9855
rect 31880 9820 31890 9855
rect 31925 9820 31935 9855
rect 31970 9820 31980 9855
rect 32015 9820 32025 9855
rect 32060 9820 32070 9855
rect 32105 9820 32115 9855
rect 32150 9820 32160 9855
rect 32195 9820 32205 9855
rect 32240 9820 32250 9855
rect 32285 9820 32295 9855
rect 32330 9820 32340 9855
rect 32375 9820 32385 9855
rect 32420 9820 32430 9855
rect 32465 9820 32475 9855
rect 32510 9820 32520 9855
rect 32555 9820 32565 9855
rect 32600 9820 32610 9855
rect 32645 9820 32655 9855
rect 32690 9820 32700 9855
rect 32735 9820 32745 9855
rect 32780 9820 32790 9855
rect 32825 9820 32835 9855
rect 32870 9820 32890 9855
rect 31290 9810 32890 9820
rect 31290 9775 31305 9810
rect 31340 9775 31350 9810
rect 31385 9775 31395 9810
rect 31430 9775 31440 9810
rect 31475 9775 31485 9810
rect 31520 9775 31530 9810
rect 31565 9775 31575 9810
rect 31610 9775 31620 9810
rect 31655 9775 31665 9810
rect 31700 9775 31710 9810
rect 31745 9775 31755 9810
rect 31790 9775 31800 9810
rect 31835 9775 31845 9810
rect 31880 9775 31890 9810
rect 31925 9775 31935 9810
rect 31970 9775 31980 9810
rect 32015 9775 32025 9810
rect 32060 9775 32070 9810
rect 32105 9775 32115 9810
rect 32150 9775 32160 9810
rect 32195 9775 32205 9810
rect 32240 9775 32250 9810
rect 32285 9775 32295 9810
rect 32330 9775 32340 9810
rect 32375 9775 32385 9810
rect 32420 9775 32430 9810
rect 32465 9775 32475 9810
rect 32510 9775 32520 9810
rect 32555 9775 32565 9810
rect 32600 9775 32610 9810
rect 32645 9775 32655 9810
rect 32690 9775 32700 9810
rect 32735 9775 32745 9810
rect 32780 9775 32790 9810
rect 32825 9775 32835 9810
rect 32870 9775 32890 9810
rect 31290 9765 32890 9775
rect 31290 9730 31305 9765
rect 31340 9730 31350 9765
rect 31385 9730 31395 9765
rect 31430 9730 31440 9765
rect 31475 9730 31485 9765
rect 31520 9730 31530 9765
rect 31565 9730 31575 9765
rect 31610 9730 31620 9765
rect 31655 9730 31665 9765
rect 31700 9730 31710 9765
rect 31745 9730 31755 9765
rect 31790 9730 31800 9765
rect 31835 9730 31845 9765
rect 31880 9730 31890 9765
rect 31925 9730 31935 9765
rect 31970 9730 31980 9765
rect 32015 9730 32025 9765
rect 32060 9730 32070 9765
rect 32105 9730 32115 9765
rect 32150 9730 32160 9765
rect 32195 9730 32205 9765
rect 32240 9730 32250 9765
rect 32285 9730 32295 9765
rect 32330 9730 32340 9765
rect 32375 9730 32385 9765
rect 32420 9730 32430 9765
rect 32465 9730 32475 9765
rect 32510 9730 32520 9765
rect 32555 9730 32565 9765
rect 32600 9730 32610 9765
rect 32645 9730 32655 9765
rect 32690 9730 32700 9765
rect 32735 9730 32745 9765
rect 32780 9730 32790 9765
rect 32825 9730 32835 9765
rect 32870 9730 32890 9765
rect 31290 9720 32890 9730
rect 31290 9685 31305 9720
rect 31340 9685 31350 9720
rect 31385 9685 31395 9720
rect 31430 9685 31440 9720
rect 31475 9685 31485 9720
rect 31520 9685 31530 9720
rect 31565 9685 31575 9720
rect 31610 9685 31620 9720
rect 31655 9685 31665 9720
rect 31700 9685 31710 9720
rect 31745 9685 31755 9720
rect 31790 9685 31800 9720
rect 31835 9685 31845 9720
rect 31880 9685 31890 9720
rect 31925 9685 31935 9720
rect 31970 9685 31980 9720
rect 32015 9685 32025 9720
rect 32060 9685 32070 9720
rect 32105 9685 32115 9720
rect 32150 9685 32160 9720
rect 32195 9685 32205 9720
rect 32240 9685 32250 9720
rect 32285 9685 32295 9720
rect 32330 9685 32340 9720
rect 32375 9685 32385 9720
rect 32420 9685 32430 9720
rect 32465 9685 32475 9720
rect 32510 9685 32520 9720
rect 32555 9685 32565 9720
rect 32600 9685 32610 9720
rect 32645 9685 32655 9720
rect 32690 9685 32700 9720
rect 32735 9685 32745 9720
rect 32780 9685 32790 9720
rect 32825 9685 32835 9720
rect 32870 9685 32890 9720
rect 31290 9675 32890 9685
rect -38770 9595 -38755 9630
rect -38720 9595 -38710 9630
rect -38675 9595 -38665 9630
rect -38630 9595 -38620 9630
rect -38585 9595 -38575 9630
rect -38540 9595 -38530 9630
rect -38495 9595 -38485 9630
rect -38450 9595 -38440 9630
rect -38405 9595 -38395 9630
rect -38360 9595 -38350 9630
rect -38315 9595 -38305 9630
rect -38270 9595 -38260 9630
rect -38225 9595 -38215 9630
rect -38180 9595 -38170 9630
rect -38135 9595 -38125 9630
rect -38090 9595 -38080 9630
rect -38045 9595 -38035 9630
rect -38000 9595 -37990 9630
rect -37955 9595 -37945 9630
rect -37910 9595 -37900 9630
rect -37865 9595 -37855 9630
rect -37820 9595 -37810 9630
rect -37775 9595 -37765 9630
rect -37730 9595 -37720 9630
rect -37685 9595 -37675 9630
rect -37640 9595 -37630 9630
rect -37595 9595 -37585 9630
rect -37550 9595 -37540 9630
rect -37505 9595 -37495 9630
rect -37460 9595 -37450 9630
rect -37415 9595 -37405 9630
rect -37370 9595 -37360 9630
rect -37325 9595 -37315 9630
rect -37280 9595 -37270 9630
rect -37235 9595 -37225 9630
rect -37190 9595 -37170 9630
rect -38770 9585 -37170 9595
rect -38770 9550 -38755 9585
rect -38720 9550 -38710 9585
rect -38675 9550 -38665 9585
rect -38630 9550 -38620 9585
rect -38585 9550 -38575 9585
rect -38540 9550 -38530 9585
rect -38495 9550 -38485 9585
rect -38450 9550 -38440 9585
rect -38405 9550 -38395 9585
rect -38360 9550 -38350 9585
rect -38315 9550 -38305 9585
rect -38270 9550 -38260 9585
rect -38225 9550 -38215 9585
rect -38180 9550 -38170 9585
rect -38135 9550 -38125 9585
rect -38090 9550 -38080 9585
rect -38045 9550 -38035 9585
rect -38000 9550 -37990 9585
rect -37955 9550 -37945 9585
rect -37910 9550 -37900 9585
rect -37865 9550 -37855 9585
rect -37820 9550 -37810 9585
rect -37775 9550 -37765 9585
rect -37730 9550 -37720 9585
rect -37685 9550 -37675 9585
rect -37640 9550 -37630 9585
rect -37595 9550 -37585 9585
rect -37550 9550 -37540 9585
rect -37505 9550 -37495 9585
rect -37460 9550 -37450 9585
rect -37415 9550 -37405 9585
rect -37370 9550 -37360 9585
rect -37325 9550 -37315 9585
rect -37280 9550 -37270 9585
rect -37235 9550 -37225 9585
rect -37190 9550 -37170 9585
rect -38770 9540 -37170 9550
rect -38770 9505 -38755 9540
rect -38720 9505 -38710 9540
rect -38675 9505 -38665 9540
rect -38630 9505 -38620 9540
rect -38585 9505 -38575 9540
rect -38540 9505 -38530 9540
rect -38495 9505 -38485 9540
rect -38450 9505 -38440 9540
rect -38405 9505 -38395 9540
rect -38360 9505 -38350 9540
rect -38315 9505 -38305 9540
rect -38270 9505 -38260 9540
rect -38225 9505 -38215 9540
rect -38180 9505 -38170 9540
rect -38135 9505 -38125 9540
rect -38090 9505 -38080 9540
rect -38045 9505 -38035 9540
rect -38000 9505 -37990 9540
rect -37955 9505 -37945 9540
rect -37910 9505 -37900 9540
rect -37865 9505 -37855 9540
rect -37820 9505 -37810 9540
rect -37775 9505 -37765 9540
rect -37730 9505 -37720 9540
rect -37685 9505 -37675 9540
rect -37640 9505 -37630 9540
rect -37595 9505 -37585 9540
rect -37550 9505 -37540 9540
rect -37505 9505 -37495 9540
rect -37460 9505 -37450 9540
rect -37415 9505 -37405 9540
rect -37370 9505 -37360 9540
rect -37325 9505 -37315 9540
rect -37280 9505 -37270 9540
rect -37235 9505 -37225 9540
rect -37190 9505 -37170 9540
rect -38770 9495 -37170 9505
rect -38770 9460 -38755 9495
rect -38720 9460 -38710 9495
rect -38675 9460 -38665 9495
rect -38630 9460 -38620 9495
rect -38585 9460 -38575 9495
rect -38540 9460 -38530 9495
rect -38495 9460 -38485 9495
rect -38450 9460 -38440 9495
rect -38405 9460 -38395 9495
rect -38360 9460 -38350 9495
rect -38315 9460 -38305 9495
rect -38270 9460 -38260 9495
rect -38225 9460 -38215 9495
rect -38180 9460 -38170 9495
rect -38135 9460 -38125 9495
rect -38090 9460 -38080 9495
rect -38045 9460 -38035 9495
rect -38000 9460 -37990 9495
rect -37955 9460 -37945 9495
rect -37910 9460 -37900 9495
rect -37865 9460 -37855 9495
rect -37820 9460 -37810 9495
rect -37775 9460 -37765 9495
rect -37730 9460 -37720 9495
rect -37685 9460 -37675 9495
rect -37640 9460 -37630 9495
rect -37595 9460 -37585 9495
rect -37550 9460 -37540 9495
rect -37505 9460 -37495 9495
rect -37460 9460 -37450 9495
rect -37415 9460 -37405 9495
rect -37370 9460 -37360 9495
rect -37325 9460 -37315 9495
rect -37280 9460 -37270 9495
rect -37235 9460 -37225 9495
rect -37190 9460 -37170 9495
rect -38770 9450 -37170 9460
rect -38770 9415 -38755 9450
rect -38720 9415 -38710 9450
rect -38675 9415 -38665 9450
rect -38630 9415 -38620 9450
rect -38585 9415 -38575 9450
rect -38540 9415 -38530 9450
rect -38495 9415 -38485 9450
rect -38450 9415 -38440 9450
rect -38405 9415 -38395 9450
rect -38360 9415 -38350 9450
rect -38315 9415 -38305 9450
rect -38270 9415 -38260 9450
rect -38225 9415 -38215 9450
rect -38180 9415 -38170 9450
rect -38135 9415 -38125 9450
rect -38090 9415 -38080 9450
rect -38045 9415 -38035 9450
rect -38000 9415 -37990 9450
rect -37955 9415 -37945 9450
rect -37910 9415 -37900 9450
rect -37865 9415 -37855 9450
rect -37820 9415 -37810 9450
rect -37775 9415 -37765 9450
rect -37730 9415 -37720 9450
rect -37685 9415 -37675 9450
rect -37640 9415 -37630 9450
rect -37595 9415 -37585 9450
rect -37550 9415 -37540 9450
rect -37505 9415 -37495 9450
rect -37460 9415 -37450 9450
rect -37415 9415 -37405 9450
rect -37370 9415 -37360 9450
rect -37325 9415 -37315 9450
rect -37280 9415 -37270 9450
rect -37235 9415 -37225 9450
rect -37190 9415 -37170 9450
rect -38770 9405 -37170 9415
rect -38770 9370 -38755 9405
rect -38720 9370 -38710 9405
rect -38675 9370 -38665 9405
rect -38630 9370 -38620 9405
rect -38585 9370 -38575 9405
rect -38540 9370 -38530 9405
rect -38495 9370 -38485 9405
rect -38450 9370 -38440 9405
rect -38405 9370 -38395 9405
rect -38360 9370 -38350 9405
rect -38315 9370 -38305 9405
rect -38270 9370 -38260 9405
rect -38225 9370 -38215 9405
rect -38180 9370 -38170 9405
rect -38135 9370 -38125 9405
rect -38090 9370 -38080 9405
rect -38045 9370 -38035 9405
rect -38000 9370 -37990 9405
rect -37955 9370 -37945 9405
rect -37910 9370 -37900 9405
rect -37865 9370 -37855 9405
rect -37820 9370 -37810 9405
rect -37775 9370 -37765 9405
rect -37730 9370 -37720 9405
rect -37685 9370 -37675 9405
rect -37640 9370 -37630 9405
rect -37595 9370 -37585 9405
rect -37550 9370 -37540 9405
rect -37505 9370 -37495 9405
rect -37460 9370 -37450 9405
rect -37415 9370 -37405 9405
rect -37370 9370 -37360 9405
rect -37325 9370 -37315 9405
rect -37280 9370 -37270 9405
rect -37235 9370 -37225 9405
rect -37190 9370 -37170 9405
rect -38770 9360 -37170 9370
rect -38770 9325 -38755 9360
rect -38720 9325 -38710 9360
rect -38675 9325 -38665 9360
rect -38630 9325 -38620 9360
rect -38585 9325 -38575 9360
rect -38540 9325 -38530 9360
rect -38495 9325 -38485 9360
rect -38450 9325 -38440 9360
rect -38405 9325 -38395 9360
rect -38360 9325 -38350 9360
rect -38315 9325 -38305 9360
rect -38270 9325 -38260 9360
rect -38225 9325 -38215 9360
rect -38180 9325 -38170 9360
rect -38135 9325 -38125 9360
rect -38090 9325 -38080 9360
rect -38045 9325 -38035 9360
rect -38000 9325 -37990 9360
rect -37955 9325 -37945 9360
rect -37910 9325 -37900 9360
rect -37865 9325 -37855 9360
rect -37820 9325 -37810 9360
rect -37775 9325 -37765 9360
rect -37730 9325 -37720 9360
rect -37685 9325 -37675 9360
rect -37640 9325 -37630 9360
rect -37595 9325 -37585 9360
rect -37550 9325 -37540 9360
rect -37505 9325 -37495 9360
rect -37460 9325 -37450 9360
rect -37415 9325 -37405 9360
rect -37370 9325 -37360 9360
rect -37325 9325 -37315 9360
rect -37280 9325 -37270 9360
rect -37235 9325 -37225 9360
rect -37190 9325 -37170 9360
rect -38770 9315 -37170 9325
rect -38770 9280 -38755 9315
rect -38720 9280 -38710 9315
rect -38675 9280 -38665 9315
rect -38630 9280 -38620 9315
rect -38585 9280 -38575 9315
rect -38540 9280 -38530 9315
rect -38495 9280 -38485 9315
rect -38450 9280 -38440 9315
rect -38405 9280 -38395 9315
rect -38360 9280 -38350 9315
rect -38315 9280 -38305 9315
rect -38270 9280 -38260 9315
rect -38225 9280 -38215 9315
rect -38180 9280 -38170 9315
rect -38135 9280 -38125 9315
rect -38090 9280 -38080 9315
rect -38045 9280 -38035 9315
rect -38000 9280 -37990 9315
rect -37955 9280 -37945 9315
rect -37910 9280 -37900 9315
rect -37865 9280 -37855 9315
rect -37820 9280 -37810 9315
rect -37775 9280 -37765 9315
rect -37730 9280 -37720 9315
rect -37685 9280 -37675 9315
rect -37640 9280 -37630 9315
rect -37595 9280 -37585 9315
rect -37550 9280 -37540 9315
rect -37505 9280 -37495 9315
rect -37460 9280 -37450 9315
rect -37415 9280 -37405 9315
rect -37370 9280 -37360 9315
rect -37325 9280 -37315 9315
rect -37280 9280 -37270 9315
rect -37235 9280 -37225 9315
rect -37190 9280 -37170 9315
rect -38770 9270 -37170 9280
rect -38770 9235 -38755 9270
rect -38720 9235 -38710 9270
rect -38675 9235 -38665 9270
rect -38630 9235 -38620 9270
rect -38585 9235 -38575 9270
rect -38540 9235 -38530 9270
rect -38495 9235 -38485 9270
rect -38450 9235 -38440 9270
rect -38405 9235 -38395 9270
rect -38360 9235 -38350 9270
rect -38315 9235 -38305 9270
rect -38270 9235 -38260 9270
rect -38225 9235 -38215 9270
rect -38180 9235 -38170 9270
rect -38135 9235 -38125 9270
rect -38090 9235 -38080 9270
rect -38045 9235 -38035 9270
rect -38000 9235 -37990 9270
rect -37955 9235 -37945 9270
rect -37910 9235 -37900 9270
rect -37865 9235 -37855 9270
rect -37820 9235 -37810 9270
rect -37775 9235 -37765 9270
rect -37730 9235 -37720 9270
rect -37685 9235 -37675 9270
rect -37640 9235 -37630 9270
rect -37595 9235 -37585 9270
rect -37550 9235 -37540 9270
rect -37505 9235 -37495 9270
rect -37460 9235 -37450 9270
rect -37415 9235 -37405 9270
rect -37370 9235 -37360 9270
rect -37325 9235 -37315 9270
rect -37280 9235 -37270 9270
rect -37235 9235 -37225 9270
rect -37190 9235 -37170 9270
rect -38770 9225 -37170 9235
rect -38770 9190 -38755 9225
rect -38720 9190 -38710 9225
rect -38675 9190 -38665 9225
rect -38630 9190 -38620 9225
rect -38585 9190 -38575 9225
rect -38540 9190 -38530 9225
rect -38495 9190 -38485 9225
rect -38450 9190 -38440 9225
rect -38405 9190 -38395 9225
rect -38360 9190 -38350 9225
rect -38315 9190 -38305 9225
rect -38270 9190 -38260 9225
rect -38225 9190 -38215 9225
rect -38180 9190 -38170 9225
rect -38135 9190 -38125 9225
rect -38090 9190 -38080 9225
rect -38045 9190 -38035 9225
rect -38000 9190 -37990 9225
rect -37955 9190 -37945 9225
rect -37910 9190 -37900 9225
rect -37865 9190 -37855 9225
rect -37820 9190 -37810 9225
rect -37775 9190 -37765 9225
rect -37730 9190 -37720 9225
rect -37685 9190 -37675 9225
rect -37640 9190 -37630 9225
rect -37595 9190 -37585 9225
rect -37550 9190 -37540 9225
rect -37505 9190 -37495 9225
rect -37460 9190 -37450 9225
rect -37415 9190 -37405 9225
rect -37370 9190 -37360 9225
rect -37325 9190 -37315 9225
rect -37280 9190 -37270 9225
rect -37235 9190 -37225 9225
rect -37190 9190 -37170 9225
rect -38770 9180 -37170 9190
rect -38770 9145 -38755 9180
rect -38720 9145 -38710 9180
rect -38675 9145 -38665 9180
rect -38630 9145 -38620 9180
rect -38585 9145 -38575 9180
rect -38540 9145 -38530 9180
rect -38495 9145 -38485 9180
rect -38450 9145 -38440 9180
rect -38405 9145 -38395 9180
rect -38360 9145 -38350 9180
rect -38315 9145 -38305 9180
rect -38270 9145 -38260 9180
rect -38225 9145 -38215 9180
rect -38180 9145 -38170 9180
rect -38135 9145 -38125 9180
rect -38090 9145 -38080 9180
rect -38045 9145 -38035 9180
rect -38000 9145 -37990 9180
rect -37955 9145 -37945 9180
rect -37910 9145 -37900 9180
rect -37865 9145 -37855 9180
rect -37820 9145 -37810 9180
rect -37775 9145 -37765 9180
rect -37730 9145 -37720 9180
rect -37685 9145 -37675 9180
rect -37640 9145 -37630 9180
rect -37595 9145 -37585 9180
rect -37550 9145 -37540 9180
rect -37505 9145 -37495 9180
rect -37460 9145 -37450 9180
rect -37415 9145 -37405 9180
rect -37370 9145 -37360 9180
rect -37325 9145 -37315 9180
rect -37280 9145 -37270 9180
rect -37235 9145 -37225 9180
rect -37190 9145 -37170 9180
rect -38770 9135 -37170 9145
rect -38770 9100 -38755 9135
rect -38720 9100 -38710 9135
rect -38675 9100 -38665 9135
rect -38630 9100 -38620 9135
rect -38585 9100 -38575 9135
rect -38540 9100 -38530 9135
rect -38495 9100 -38485 9135
rect -38450 9100 -38440 9135
rect -38405 9100 -38395 9135
rect -38360 9100 -38350 9135
rect -38315 9100 -38305 9135
rect -38270 9100 -38260 9135
rect -38225 9100 -38215 9135
rect -38180 9100 -38170 9135
rect -38135 9100 -38125 9135
rect -38090 9100 -38080 9135
rect -38045 9100 -38035 9135
rect -38000 9100 -37990 9135
rect -37955 9100 -37945 9135
rect -37910 9100 -37900 9135
rect -37865 9100 -37855 9135
rect -37820 9100 -37810 9135
rect -37775 9100 -37765 9135
rect -37730 9100 -37720 9135
rect -37685 9100 -37675 9135
rect -37640 9100 -37630 9135
rect -37595 9100 -37585 9135
rect -37550 9100 -37540 9135
rect -37505 9100 -37495 9135
rect -37460 9100 -37450 9135
rect -37415 9100 -37405 9135
rect -37370 9100 -37360 9135
rect -37325 9100 -37315 9135
rect -37280 9100 -37270 9135
rect -37235 9100 -37225 9135
rect -37190 9100 -37170 9135
rect -38770 9090 -37170 9100
rect -38770 9055 -38755 9090
rect -38720 9055 -38710 9090
rect -38675 9055 -38665 9090
rect -38630 9055 -38620 9090
rect -38585 9055 -38575 9090
rect -38540 9055 -38530 9090
rect -38495 9055 -38485 9090
rect -38450 9055 -38440 9090
rect -38405 9055 -38395 9090
rect -38360 9055 -38350 9090
rect -38315 9055 -38305 9090
rect -38270 9055 -38260 9090
rect -38225 9055 -38215 9090
rect -38180 9055 -38170 9090
rect -38135 9055 -38125 9090
rect -38090 9055 -38080 9090
rect -38045 9055 -38035 9090
rect -38000 9055 -37990 9090
rect -37955 9055 -37945 9090
rect -37910 9055 -37900 9090
rect -37865 9055 -37855 9090
rect -37820 9055 -37810 9090
rect -37775 9055 -37765 9090
rect -37730 9055 -37720 9090
rect -37685 9055 -37675 9090
rect -37640 9055 -37630 9090
rect -37595 9055 -37585 9090
rect -37550 9055 -37540 9090
rect -37505 9055 -37495 9090
rect -37460 9055 -37450 9090
rect -37415 9055 -37405 9090
rect -37370 9055 -37360 9090
rect -37325 9055 -37315 9090
rect -37280 9055 -37270 9090
rect -37235 9055 -37225 9090
rect -37190 9055 -37170 9090
rect -38770 9045 -37170 9055
rect -38770 9010 -38755 9045
rect -38720 9010 -38710 9045
rect -38675 9010 -38665 9045
rect -38630 9010 -38620 9045
rect -38585 9010 -38575 9045
rect -38540 9010 -38530 9045
rect -38495 9010 -38485 9045
rect -38450 9010 -38440 9045
rect -38405 9010 -38395 9045
rect -38360 9010 -38350 9045
rect -38315 9010 -38305 9045
rect -38270 9010 -38260 9045
rect -38225 9010 -38215 9045
rect -38180 9010 -38170 9045
rect -38135 9010 -38125 9045
rect -38090 9010 -38080 9045
rect -38045 9010 -38035 9045
rect -38000 9010 -37990 9045
rect -37955 9010 -37945 9045
rect -37910 9010 -37900 9045
rect -37865 9010 -37855 9045
rect -37820 9010 -37810 9045
rect -37775 9010 -37765 9045
rect -37730 9010 -37720 9045
rect -37685 9010 -37675 9045
rect -37640 9010 -37630 9045
rect -37595 9010 -37585 9045
rect -37550 9010 -37540 9045
rect -37505 9010 -37495 9045
rect -37460 9010 -37450 9045
rect -37415 9010 -37405 9045
rect -37370 9010 -37360 9045
rect -37325 9010 -37315 9045
rect -37280 9010 -37270 9045
rect -37235 9010 -37225 9045
rect -37190 9010 -37170 9045
rect -38770 9000 -37170 9010
rect -38770 8965 -38755 9000
rect -38720 8965 -38710 9000
rect -38675 8965 -38665 9000
rect -38630 8965 -38620 9000
rect -38585 8965 -38575 9000
rect -38540 8965 -38530 9000
rect -38495 8965 -38485 9000
rect -38450 8965 -38440 9000
rect -38405 8965 -38395 9000
rect -38360 8965 -38350 9000
rect -38315 8965 -38305 9000
rect -38270 8965 -38260 9000
rect -38225 8965 -38215 9000
rect -38180 8965 -38170 9000
rect -38135 8965 -38125 9000
rect -38090 8965 -38080 9000
rect -38045 8965 -38035 9000
rect -38000 8965 -37990 9000
rect -37955 8965 -37945 9000
rect -37910 8965 -37900 9000
rect -37865 8965 -37855 9000
rect -37820 8965 -37810 9000
rect -37775 8965 -37765 9000
rect -37730 8965 -37720 9000
rect -37685 8965 -37675 9000
rect -37640 8965 -37630 9000
rect -37595 8965 -37585 9000
rect -37550 8965 -37540 9000
rect -37505 8965 -37495 9000
rect -37460 8965 -37450 9000
rect -37415 8965 -37405 9000
rect -37370 8965 -37360 9000
rect -37325 8965 -37315 9000
rect -37280 8965 -37270 9000
rect -37235 8965 -37225 9000
rect -37190 8965 -37170 9000
rect -38770 8955 -37170 8965
rect -38770 8920 -38755 8955
rect -38720 8920 -38710 8955
rect -38675 8920 -38665 8955
rect -38630 8920 -38620 8955
rect -38585 8920 -38575 8955
rect -38540 8920 -38530 8955
rect -38495 8920 -38485 8955
rect -38450 8920 -38440 8955
rect -38405 8920 -38395 8955
rect -38360 8920 -38350 8955
rect -38315 8920 -38305 8955
rect -38270 8920 -38260 8955
rect -38225 8920 -38215 8955
rect -38180 8920 -38170 8955
rect -38135 8920 -38125 8955
rect -38090 8920 -38080 8955
rect -38045 8920 -38035 8955
rect -38000 8920 -37990 8955
rect -37955 8920 -37945 8955
rect -37910 8920 -37900 8955
rect -37865 8920 -37855 8955
rect -37820 8920 -37810 8955
rect -37775 8920 -37765 8955
rect -37730 8920 -37720 8955
rect -37685 8920 -37675 8955
rect -37640 8920 -37630 8955
rect -37595 8920 -37585 8955
rect -37550 8920 -37540 8955
rect -37505 8920 -37495 8955
rect -37460 8920 -37450 8955
rect -37415 8920 -37405 8955
rect -37370 8920 -37360 8955
rect -37325 8920 -37315 8955
rect -37280 8920 -37270 8955
rect -37235 8920 -37225 8955
rect -37190 8920 -37170 8955
rect -38770 8910 -37170 8920
rect -38770 8875 -38755 8910
rect -38720 8875 -38710 8910
rect -38675 8875 -38665 8910
rect -38630 8875 -38620 8910
rect -38585 8875 -38575 8910
rect -38540 8875 -38530 8910
rect -38495 8875 -38485 8910
rect -38450 8875 -38440 8910
rect -38405 8875 -38395 8910
rect -38360 8875 -38350 8910
rect -38315 8875 -38305 8910
rect -38270 8875 -38260 8910
rect -38225 8875 -38215 8910
rect -38180 8875 -38170 8910
rect -38135 8875 -38125 8910
rect -38090 8875 -38080 8910
rect -38045 8875 -38035 8910
rect -38000 8875 -37990 8910
rect -37955 8875 -37945 8910
rect -37910 8875 -37900 8910
rect -37865 8875 -37855 8910
rect -37820 8875 -37810 8910
rect -37775 8875 -37765 8910
rect -37730 8875 -37720 8910
rect -37685 8875 -37675 8910
rect -37640 8875 -37630 8910
rect -37595 8875 -37585 8910
rect -37550 8875 -37540 8910
rect -37505 8875 -37495 8910
rect -37460 8875 -37450 8910
rect -37415 8875 -37405 8910
rect -37370 8875 -37360 8910
rect -37325 8875 -37315 8910
rect -37280 8875 -37270 8910
rect -37235 8875 -37225 8910
rect -37190 8875 -37170 8910
rect -38770 8865 -37170 8875
rect -38770 8830 -38755 8865
rect -38720 8830 -38710 8865
rect -38675 8830 -38665 8865
rect -38630 8830 -38620 8865
rect -38585 8830 -38575 8865
rect -38540 8830 -38530 8865
rect -38495 8830 -38485 8865
rect -38450 8830 -38440 8865
rect -38405 8830 -38395 8865
rect -38360 8830 -38350 8865
rect -38315 8830 -38305 8865
rect -38270 8830 -38260 8865
rect -38225 8830 -38215 8865
rect -38180 8830 -38170 8865
rect -38135 8830 -38125 8865
rect -38090 8830 -38080 8865
rect -38045 8830 -38035 8865
rect -38000 8830 -37990 8865
rect -37955 8830 -37945 8865
rect -37910 8830 -37900 8865
rect -37865 8830 -37855 8865
rect -37820 8830 -37810 8865
rect -37775 8830 -37765 8865
rect -37730 8830 -37720 8865
rect -37685 8830 -37675 8865
rect -37640 8830 -37630 8865
rect -37595 8830 -37585 8865
rect -37550 8830 -37540 8865
rect -37505 8830 -37495 8865
rect -37460 8830 -37450 8865
rect -37415 8830 -37405 8865
rect -37370 8830 -37360 8865
rect -37325 8830 -37315 8865
rect -37280 8830 -37270 8865
rect -37235 8830 -37225 8865
rect -37190 8830 -37170 8865
rect -38770 8820 -37170 8830
rect -38770 8785 -38755 8820
rect -38720 8785 -38710 8820
rect -38675 8785 -38665 8820
rect -38630 8785 -38620 8820
rect -38585 8785 -38575 8820
rect -38540 8785 -38530 8820
rect -38495 8785 -38485 8820
rect -38450 8785 -38440 8820
rect -38405 8785 -38395 8820
rect -38360 8785 -38350 8820
rect -38315 8785 -38305 8820
rect -38270 8785 -38260 8820
rect -38225 8785 -38215 8820
rect -38180 8785 -38170 8820
rect -38135 8785 -38125 8820
rect -38090 8785 -38080 8820
rect -38045 8785 -38035 8820
rect -38000 8785 -37990 8820
rect -37955 8785 -37945 8820
rect -37910 8785 -37900 8820
rect -37865 8785 -37855 8820
rect -37820 8785 -37810 8820
rect -37775 8785 -37765 8820
rect -37730 8785 -37720 8820
rect -37685 8785 -37675 8820
rect -37640 8785 -37630 8820
rect -37595 8785 -37585 8820
rect -37550 8785 -37540 8820
rect -37505 8785 -37495 8820
rect -37460 8785 -37450 8820
rect -37415 8785 -37405 8820
rect -37370 8785 -37360 8820
rect -37325 8785 -37315 8820
rect -37280 8785 -37270 8820
rect -37235 8785 -37225 8820
rect -37190 8785 -37170 8820
rect -38770 8775 -37170 8785
rect -38770 8740 -38755 8775
rect -38720 8740 -38710 8775
rect -38675 8740 -38665 8775
rect -38630 8740 -38620 8775
rect -38585 8740 -38575 8775
rect -38540 8740 -38530 8775
rect -38495 8740 -38485 8775
rect -38450 8740 -38440 8775
rect -38405 8740 -38395 8775
rect -38360 8740 -38350 8775
rect -38315 8740 -38305 8775
rect -38270 8740 -38260 8775
rect -38225 8740 -38215 8775
rect -38180 8740 -38170 8775
rect -38135 8740 -38125 8775
rect -38090 8740 -38080 8775
rect -38045 8740 -38035 8775
rect -38000 8740 -37990 8775
rect -37955 8740 -37945 8775
rect -37910 8740 -37900 8775
rect -37865 8740 -37855 8775
rect -37820 8740 -37810 8775
rect -37775 8740 -37765 8775
rect -37730 8740 -37720 8775
rect -37685 8740 -37675 8775
rect -37640 8740 -37630 8775
rect -37595 8740 -37585 8775
rect -37550 8740 -37540 8775
rect -37505 8740 -37495 8775
rect -37460 8740 -37450 8775
rect -37415 8740 -37405 8775
rect -37370 8740 -37360 8775
rect -37325 8740 -37315 8775
rect -37280 8740 -37270 8775
rect -37235 8740 -37225 8775
rect -37190 8740 -37170 8775
rect -38770 8730 -37170 8740
rect -38770 8695 -38755 8730
rect -38720 8695 -38710 8730
rect -38675 8695 -38665 8730
rect -38630 8695 -38620 8730
rect -38585 8695 -38575 8730
rect -38540 8695 -38530 8730
rect -38495 8695 -38485 8730
rect -38450 8695 -38440 8730
rect -38405 8695 -38395 8730
rect -38360 8695 -38350 8730
rect -38315 8695 -38305 8730
rect -38270 8695 -38260 8730
rect -38225 8695 -38215 8730
rect -38180 8695 -38170 8730
rect -38135 8695 -38125 8730
rect -38090 8695 -38080 8730
rect -38045 8695 -38035 8730
rect -38000 8695 -37990 8730
rect -37955 8695 -37945 8730
rect -37910 8695 -37900 8730
rect -37865 8695 -37855 8730
rect -37820 8695 -37810 8730
rect -37775 8695 -37765 8730
rect -37730 8695 -37720 8730
rect -37685 8695 -37675 8730
rect -37640 8695 -37630 8730
rect -37595 8695 -37585 8730
rect -37550 8695 -37540 8730
rect -37505 8695 -37495 8730
rect -37460 8695 -37450 8730
rect -37415 8695 -37405 8730
rect -37370 8695 -37360 8730
rect -37325 8695 -37315 8730
rect -37280 8695 -37270 8730
rect -37235 8695 -37225 8730
rect -37190 8695 -37170 8730
rect -38770 8685 -37170 8695
rect -38770 8650 -38755 8685
rect -38720 8650 -38710 8685
rect -38675 8650 -38665 8685
rect -38630 8650 -38620 8685
rect -38585 8650 -38575 8685
rect -38540 8650 -38530 8685
rect -38495 8650 -38485 8685
rect -38450 8650 -38440 8685
rect -38405 8650 -38395 8685
rect -38360 8650 -38350 8685
rect -38315 8650 -38305 8685
rect -38270 8650 -38260 8685
rect -38225 8650 -38215 8685
rect -38180 8650 -38170 8685
rect -38135 8650 -38125 8685
rect -38090 8650 -38080 8685
rect -38045 8650 -38035 8685
rect -38000 8650 -37990 8685
rect -37955 8650 -37945 8685
rect -37910 8650 -37900 8685
rect -37865 8650 -37855 8685
rect -37820 8650 -37810 8685
rect -37775 8650 -37765 8685
rect -37730 8650 -37720 8685
rect -37685 8650 -37675 8685
rect -37640 8650 -37630 8685
rect -37595 8650 -37585 8685
rect -37550 8650 -37540 8685
rect -37505 8650 -37495 8685
rect -37460 8650 -37450 8685
rect -37415 8650 -37405 8685
rect -37370 8650 -37360 8685
rect -37325 8650 -37315 8685
rect -37280 8650 -37270 8685
rect -37235 8650 -37225 8685
rect -37190 8650 -37170 8685
rect -38770 8640 -37170 8650
rect -38770 8605 -38755 8640
rect -38720 8605 -38710 8640
rect -38675 8605 -38665 8640
rect -38630 8605 -38620 8640
rect -38585 8605 -38575 8640
rect -38540 8605 -38530 8640
rect -38495 8605 -38485 8640
rect -38450 8605 -38440 8640
rect -38405 8605 -38395 8640
rect -38360 8605 -38350 8640
rect -38315 8605 -38305 8640
rect -38270 8605 -38260 8640
rect -38225 8605 -38215 8640
rect -38180 8605 -38170 8640
rect -38135 8605 -38125 8640
rect -38090 8605 -38080 8640
rect -38045 8605 -38035 8640
rect -38000 8605 -37990 8640
rect -37955 8605 -37945 8640
rect -37910 8605 -37900 8640
rect -37865 8605 -37855 8640
rect -37820 8605 -37810 8640
rect -37775 8605 -37765 8640
rect -37730 8605 -37720 8640
rect -37685 8605 -37675 8640
rect -37640 8605 -37630 8640
rect -37595 8605 -37585 8640
rect -37550 8605 -37540 8640
rect -37505 8605 -37495 8640
rect -37460 8605 -37450 8640
rect -37415 8605 -37405 8640
rect -37370 8605 -37360 8640
rect -37325 8605 -37315 8640
rect -37280 8605 -37270 8640
rect -37235 8605 -37225 8640
rect -37190 8605 -37170 8640
rect -38770 8595 -37170 8605
rect -38770 8560 -38755 8595
rect -38720 8560 -38710 8595
rect -38675 8560 -38665 8595
rect -38630 8560 -38620 8595
rect -38585 8560 -38575 8595
rect -38540 8560 -38530 8595
rect -38495 8560 -38485 8595
rect -38450 8560 -38440 8595
rect -38405 8560 -38395 8595
rect -38360 8560 -38350 8595
rect -38315 8560 -38305 8595
rect -38270 8560 -38260 8595
rect -38225 8560 -38215 8595
rect -38180 8560 -38170 8595
rect -38135 8560 -38125 8595
rect -38090 8560 -38080 8595
rect -38045 8560 -38035 8595
rect -38000 8560 -37990 8595
rect -37955 8560 -37945 8595
rect -37910 8560 -37900 8595
rect -37865 8560 -37855 8595
rect -37820 8560 -37810 8595
rect -37775 8560 -37765 8595
rect -37730 8560 -37720 8595
rect -37685 8560 -37675 8595
rect -37640 8560 -37630 8595
rect -37595 8560 -37585 8595
rect -37550 8560 -37540 8595
rect -37505 8560 -37495 8595
rect -37460 8560 -37450 8595
rect -37415 8560 -37405 8595
rect -37370 8560 -37360 8595
rect -37325 8560 -37315 8595
rect -37280 8560 -37270 8595
rect -37235 8560 -37225 8595
rect -37190 8560 -37170 8595
rect -38770 8550 -37170 8560
rect -38770 8515 -38755 8550
rect -38720 8515 -38710 8550
rect -38675 8515 -38665 8550
rect -38630 8515 -38620 8550
rect -38585 8515 -38575 8550
rect -38540 8515 -38530 8550
rect -38495 8515 -38485 8550
rect -38450 8515 -38440 8550
rect -38405 8515 -38395 8550
rect -38360 8515 -38350 8550
rect -38315 8515 -38305 8550
rect -38270 8515 -38260 8550
rect -38225 8515 -38215 8550
rect -38180 8515 -38170 8550
rect -38135 8515 -38125 8550
rect -38090 8515 -38080 8550
rect -38045 8515 -38035 8550
rect -38000 8515 -37990 8550
rect -37955 8515 -37945 8550
rect -37910 8515 -37900 8550
rect -37865 8515 -37855 8550
rect -37820 8515 -37810 8550
rect -37775 8515 -37765 8550
rect -37730 8515 -37720 8550
rect -37685 8515 -37675 8550
rect -37640 8515 -37630 8550
rect -37595 8515 -37585 8550
rect -37550 8515 -37540 8550
rect -37505 8515 -37495 8550
rect -37460 8515 -37450 8550
rect -37415 8515 -37405 8550
rect -37370 8515 -37360 8550
rect -37325 8515 -37315 8550
rect -37280 8515 -37270 8550
rect -37235 8515 -37225 8550
rect -37190 8515 -37170 8550
rect -38770 8505 -37170 8515
rect -38770 8470 -38755 8505
rect -38720 8470 -38710 8505
rect -38675 8470 -38665 8505
rect -38630 8470 -38620 8505
rect -38585 8470 -38575 8505
rect -38540 8470 -38530 8505
rect -38495 8470 -38485 8505
rect -38450 8470 -38440 8505
rect -38405 8470 -38395 8505
rect -38360 8470 -38350 8505
rect -38315 8470 -38305 8505
rect -38270 8470 -38260 8505
rect -38225 8470 -38215 8505
rect -38180 8470 -38170 8505
rect -38135 8470 -38125 8505
rect -38090 8470 -38080 8505
rect -38045 8470 -38035 8505
rect -38000 8470 -37990 8505
rect -37955 8470 -37945 8505
rect -37910 8470 -37900 8505
rect -37865 8470 -37855 8505
rect -37820 8470 -37810 8505
rect -37775 8470 -37765 8505
rect -37730 8470 -37720 8505
rect -37685 8470 -37675 8505
rect -37640 8470 -37630 8505
rect -37595 8470 -37585 8505
rect -37550 8470 -37540 8505
rect -37505 8470 -37495 8505
rect -37460 8470 -37450 8505
rect -37415 8470 -37405 8505
rect -37370 8470 -37360 8505
rect -37325 8470 -37315 8505
rect -37280 8470 -37270 8505
rect -37235 8470 -37225 8505
rect -37190 8470 -37170 8505
rect -38770 8460 -37170 8470
rect -38770 8425 -38755 8460
rect -38720 8425 -38710 8460
rect -38675 8425 -38665 8460
rect -38630 8425 -38620 8460
rect -38585 8425 -38575 8460
rect -38540 8425 -38530 8460
rect -38495 8425 -38485 8460
rect -38450 8425 -38440 8460
rect -38405 8425 -38395 8460
rect -38360 8425 -38350 8460
rect -38315 8425 -38305 8460
rect -38270 8425 -38260 8460
rect -38225 8425 -38215 8460
rect -38180 8425 -38170 8460
rect -38135 8425 -38125 8460
rect -38090 8425 -38080 8460
rect -38045 8425 -38035 8460
rect -38000 8425 -37990 8460
rect -37955 8425 -37945 8460
rect -37910 8425 -37900 8460
rect -37865 8425 -37855 8460
rect -37820 8425 -37810 8460
rect -37775 8425 -37765 8460
rect -37730 8425 -37720 8460
rect -37685 8425 -37675 8460
rect -37640 8425 -37630 8460
rect -37595 8425 -37585 8460
rect -37550 8425 -37540 8460
rect -37505 8425 -37495 8460
rect -37460 8425 -37450 8460
rect -37415 8425 -37405 8460
rect -37370 8425 -37360 8460
rect -37325 8425 -37315 8460
rect -37280 8425 -37270 8460
rect -37235 8425 -37225 8460
rect -37190 8425 -37170 8460
rect -38770 8415 -37170 8425
rect -38770 8380 -38755 8415
rect -38720 8380 -38710 8415
rect -38675 8380 -38665 8415
rect -38630 8380 -38620 8415
rect -38585 8380 -38575 8415
rect -38540 8380 -38530 8415
rect -38495 8380 -38485 8415
rect -38450 8380 -38440 8415
rect -38405 8380 -38395 8415
rect -38360 8380 -38350 8415
rect -38315 8380 -38305 8415
rect -38270 8380 -38260 8415
rect -38225 8380 -38215 8415
rect -38180 8380 -38170 8415
rect -38135 8380 -38125 8415
rect -38090 8380 -38080 8415
rect -38045 8380 -38035 8415
rect -38000 8380 -37990 8415
rect -37955 8380 -37945 8415
rect -37910 8380 -37900 8415
rect -37865 8380 -37855 8415
rect -37820 8380 -37810 8415
rect -37775 8380 -37765 8415
rect -37730 8380 -37720 8415
rect -37685 8380 -37675 8415
rect -37640 8380 -37630 8415
rect -37595 8380 -37585 8415
rect -37550 8380 -37540 8415
rect -37505 8380 -37495 8415
rect -37460 8380 -37450 8415
rect -37415 8380 -37405 8415
rect -37370 8380 -37360 8415
rect -37325 8380 -37315 8415
rect -37280 8380 -37270 8415
rect -37235 8380 -37225 8415
rect -37190 8380 -37170 8415
rect -38770 8370 -37170 8380
rect -38770 8335 -38755 8370
rect -38720 8335 -38710 8370
rect -38675 8335 -38665 8370
rect -38630 8335 -38620 8370
rect -38585 8335 -38575 8370
rect -38540 8335 -38530 8370
rect -38495 8335 -38485 8370
rect -38450 8335 -38440 8370
rect -38405 8335 -38395 8370
rect -38360 8335 -38350 8370
rect -38315 8335 -38305 8370
rect -38270 8335 -38260 8370
rect -38225 8335 -38215 8370
rect -38180 8335 -38170 8370
rect -38135 8335 -38125 8370
rect -38090 8335 -38080 8370
rect -38045 8335 -38035 8370
rect -38000 8335 -37990 8370
rect -37955 8335 -37945 8370
rect -37910 8335 -37900 8370
rect -37865 8335 -37855 8370
rect -37820 8335 -37810 8370
rect -37775 8335 -37765 8370
rect -37730 8335 -37720 8370
rect -37685 8335 -37675 8370
rect -37640 8335 -37630 8370
rect -37595 8335 -37585 8370
rect -37550 8335 -37540 8370
rect -37505 8335 -37495 8370
rect -37460 8335 -37450 8370
rect -37415 8335 -37405 8370
rect -37370 8335 -37360 8370
rect -37325 8335 -37315 8370
rect -37280 8335 -37270 8370
rect -37235 8335 -37225 8370
rect -37190 8335 -37170 8370
rect -38770 8325 -37170 8335
rect -38770 8290 -38755 8325
rect -38720 8290 -38710 8325
rect -38675 8290 -38665 8325
rect -38630 8290 -38620 8325
rect -38585 8290 -38575 8325
rect -38540 8290 -38530 8325
rect -38495 8290 -38485 8325
rect -38450 8290 -38440 8325
rect -38405 8290 -38395 8325
rect -38360 8290 -38350 8325
rect -38315 8290 -38305 8325
rect -38270 8290 -38260 8325
rect -38225 8290 -38215 8325
rect -38180 8290 -38170 8325
rect -38135 8290 -38125 8325
rect -38090 8290 -38080 8325
rect -38045 8290 -38035 8325
rect -38000 8290 -37990 8325
rect -37955 8290 -37945 8325
rect -37910 8290 -37900 8325
rect -37865 8290 -37855 8325
rect -37820 8290 -37810 8325
rect -37775 8290 -37765 8325
rect -37730 8290 -37720 8325
rect -37685 8290 -37675 8325
rect -37640 8290 -37630 8325
rect -37595 8290 -37585 8325
rect -37550 8290 -37540 8325
rect -37505 8290 -37495 8325
rect -37460 8290 -37450 8325
rect -37415 8290 -37405 8325
rect -37370 8290 -37360 8325
rect -37325 8290 -37315 8325
rect -37280 8290 -37270 8325
rect -37235 8290 -37225 8325
rect -37190 8290 -37170 8325
rect -38770 8280 -37170 8290
rect -38770 8245 -38755 8280
rect -38720 8245 -38710 8280
rect -38675 8245 -38665 8280
rect -38630 8245 -38620 8280
rect -38585 8245 -38575 8280
rect -38540 8245 -38530 8280
rect -38495 8245 -38485 8280
rect -38450 8245 -38440 8280
rect -38405 8245 -38395 8280
rect -38360 8245 -38350 8280
rect -38315 8245 -38305 8280
rect -38270 8245 -38260 8280
rect -38225 8245 -38215 8280
rect -38180 8245 -38170 8280
rect -38135 8245 -38125 8280
rect -38090 8245 -38080 8280
rect -38045 8245 -38035 8280
rect -38000 8245 -37990 8280
rect -37955 8245 -37945 8280
rect -37910 8245 -37900 8280
rect -37865 8245 -37855 8280
rect -37820 8245 -37810 8280
rect -37775 8245 -37765 8280
rect -37730 8245 -37720 8280
rect -37685 8245 -37675 8280
rect -37640 8245 -37630 8280
rect -37595 8245 -37585 8280
rect -37550 8245 -37540 8280
rect -37505 8245 -37495 8280
rect -37460 8245 -37450 8280
rect -37415 8245 -37405 8280
rect -37370 8245 -37360 8280
rect -37325 8245 -37315 8280
rect -37280 8245 -37270 8280
rect -37235 8245 -37225 8280
rect -37190 8245 -37170 8280
rect -38770 8235 -37170 8245
rect -38770 8200 -38755 8235
rect -38720 8200 -38710 8235
rect -38675 8200 -38665 8235
rect -38630 8200 -38620 8235
rect -38585 8200 -38575 8235
rect -38540 8200 -38530 8235
rect -38495 8200 -38485 8235
rect -38450 8200 -38440 8235
rect -38405 8200 -38395 8235
rect -38360 8200 -38350 8235
rect -38315 8200 -38305 8235
rect -38270 8200 -38260 8235
rect -38225 8200 -38215 8235
rect -38180 8200 -38170 8235
rect -38135 8200 -38125 8235
rect -38090 8200 -38080 8235
rect -38045 8200 -38035 8235
rect -38000 8200 -37990 8235
rect -37955 8200 -37945 8235
rect -37910 8200 -37900 8235
rect -37865 8200 -37855 8235
rect -37820 8200 -37810 8235
rect -37775 8200 -37765 8235
rect -37730 8200 -37720 8235
rect -37685 8200 -37675 8235
rect -37640 8200 -37630 8235
rect -37595 8200 -37585 8235
rect -37550 8200 -37540 8235
rect -37505 8200 -37495 8235
rect -37460 8200 -37450 8235
rect -37415 8200 -37405 8235
rect -37370 8200 -37360 8235
rect -37325 8200 -37315 8235
rect -37280 8200 -37270 8235
rect -37235 8200 -37225 8235
rect -37190 8200 -37170 8235
rect -38770 8190 -37170 8200
rect -38770 8155 -38755 8190
rect -38720 8155 -38710 8190
rect -38675 8155 -38665 8190
rect -38630 8155 -38620 8190
rect -38585 8155 -38575 8190
rect -38540 8155 -38530 8190
rect -38495 8155 -38485 8190
rect -38450 8155 -38440 8190
rect -38405 8155 -38395 8190
rect -38360 8155 -38350 8190
rect -38315 8155 -38305 8190
rect -38270 8155 -38260 8190
rect -38225 8155 -38215 8190
rect -38180 8155 -38170 8190
rect -38135 8155 -38125 8190
rect -38090 8155 -38080 8190
rect -38045 8155 -38035 8190
rect -38000 8155 -37990 8190
rect -37955 8155 -37945 8190
rect -37910 8155 -37900 8190
rect -37865 8155 -37855 8190
rect -37820 8155 -37810 8190
rect -37775 8155 -37765 8190
rect -37730 8155 -37720 8190
rect -37685 8155 -37675 8190
rect -37640 8155 -37630 8190
rect -37595 8155 -37585 8190
rect -37550 8155 -37540 8190
rect -37505 8155 -37495 8190
rect -37460 8155 -37450 8190
rect -37415 8155 -37405 8190
rect -37370 8155 -37360 8190
rect -37325 8155 -37315 8190
rect -37280 8155 -37270 8190
rect -37235 8155 -37225 8190
rect -37190 8155 -37170 8190
rect -38770 8145 -37170 8155
rect -38770 8110 -38755 8145
rect -38720 8110 -38710 8145
rect -38675 8110 -38665 8145
rect -38630 8110 -38620 8145
rect -38585 8110 -38575 8145
rect -38540 8110 -38530 8145
rect -38495 8110 -38485 8145
rect -38450 8110 -38440 8145
rect -38405 8110 -38395 8145
rect -38360 8110 -38350 8145
rect -38315 8110 -38305 8145
rect -38270 8110 -38260 8145
rect -38225 8110 -38215 8145
rect -38180 8110 -38170 8145
rect -38135 8110 -38125 8145
rect -38090 8110 -38080 8145
rect -38045 8110 -38035 8145
rect -38000 8110 -37990 8145
rect -37955 8110 -37945 8145
rect -37910 8110 -37900 8145
rect -37865 8110 -37855 8145
rect -37820 8110 -37810 8145
rect -37775 8110 -37765 8145
rect -37730 8110 -37720 8145
rect -37685 8110 -37675 8145
rect -37640 8110 -37630 8145
rect -37595 8110 -37585 8145
rect -37550 8110 -37540 8145
rect -37505 8110 -37495 8145
rect -37460 8110 -37450 8145
rect -37415 8110 -37405 8145
rect -37370 8110 -37360 8145
rect -37325 8110 -37315 8145
rect -37280 8110 -37270 8145
rect -37235 8110 -37225 8145
rect -37190 8110 -37170 8145
rect -38770 8105 -37170 8110
rect 1310 9640 1370 9650
rect 1310 9600 1320 9640
rect 1360 9600 1370 9640
rect 1310 9575 1370 9600
rect 1310 9535 1320 9575
rect 1360 9535 1370 9575
rect 1310 9505 1370 9535
rect 1310 9465 1320 9505
rect 1360 9465 1370 9505
rect 1310 9435 1370 9465
rect 1310 9395 1320 9435
rect 1360 9395 1370 9435
rect 1310 9365 1370 9395
rect 1310 9325 1320 9365
rect 1360 9325 1370 9365
rect 1310 9300 1370 9325
rect 1310 9260 1320 9300
rect 1360 9260 1370 9300
rect 1310 9240 1370 9260
rect 1310 9200 1320 9240
rect 1360 9200 1370 9240
rect 1310 9175 1370 9200
rect 1310 9135 1320 9175
rect 1360 9135 1370 9175
rect 1310 9105 1370 9135
rect 1310 9065 1320 9105
rect 1360 9065 1370 9105
rect 1310 9035 1370 9065
rect 1310 8995 1320 9035
rect 1360 8995 1370 9035
rect 1310 8965 1370 8995
rect 1310 8925 1320 8965
rect 1360 8925 1370 8965
rect 1310 8900 1370 8925
rect 1310 8860 1320 8900
rect 1360 8860 1370 8900
rect 1310 8840 1370 8860
rect 1310 8800 1320 8840
rect 1360 8800 1370 8840
rect 1310 8775 1370 8800
rect 1310 8735 1320 8775
rect 1360 8735 1370 8775
rect 1310 8705 1370 8735
rect 1310 8665 1320 8705
rect 1360 8665 1370 8705
rect 1310 8635 1370 8665
rect 1310 8595 1320 8635
rect 1360 8595 1370 8635
rect 1310 8565 1370 8595
rect 1310 8525 1320 8565
rect 1360 8525 1370 8565
rect 1310 8500 1370 8525
rect 1310 8460 1320 8500
rect 1360 8460 1370 8500
rect 1310 8440 1370 8460
rect 1310 8400 1320 8440
rect 1360 8400 1370 8440
rect 1310 8375 1370 8400
rect 1310 8335 1320 8375
rect 1360 8335 1370 8375
rect 1310 8305 1370 8335
rect 1310 8265 1320 8305
rect 1360 8265 1370 8305
rect 1310 8235 1370 8265
rect 1310 8195 1320 8235
rect 1360 8195 1370 8235
rect 1310 8165 1370 8195
rect 1310 8125 1320 8165
rect 1360 8125 1370 8165
rect 1310 8105 1370 8125
rect 2235 9640 2295 9650
rect 2235 9600 2245 9640
rect 2285 9600 2295 9640
rect 2235 9575 2295 9600
rect 2235 9535 2245 9575
rect 2285 9535 2295 9575
rect 2235 9505 2295 9535
rect 2235 9465 2245 9505
rect 2285 9465 2295 9505
rect 2235 9435 2295 9465
rect 2235 9395 2245 9435
rect 2285 9395 2295 9435
rect 2235 9365 2295 9395
rect 2235 9325 2245 9365
rect 2285 9325 2295 9365
rect 2235 9300 2295 9325
rect 2235 9260 2245 9300
rect 2285 9260 2295 9300
rect 2235 9240 2295 9260
rect 2235 9200 2245 9240
rect 2285 9200 2295 9240
rect 2235 9175 2295 9200
rect 2235 9135 2245 9175
rect 2285 9135 2295 9175
rect 2235 9105 2295 9135
rect 2235 9065 2245 9105
rect 2285 9065 2295 9105
rect 2235 9035 2295 9065
rect 2235 8995 2245 9035
rect 2285 8995 2295 9035
rect 2235 8965 2295 8995
rect 2235 8925 2245 8965
rect 2285 8925 2295 8965
rect 2235 8900 2295 8925
rect 2235 8860 2245 8900
rect 2285 8860 2295 8900
rect 2235 8840 2295 8860
rect 2235 8800 2245 8840
rect 2285 8800 2295 8840
rect 2235 8775 2295 8800
rect 2235 8735 2245 8775
rect 2285 8735 2295 8775
rect 2235 8705 2295 8735
rect 2235 8665 2245 8705
rect 2285 8665 2295 8705
rect 2235 8635 2295 8665
rect 2235 8595 2245 8635
rect 2285 8595 2295 8635
rect 2235 8565 2295 8595
rect 2235 8525 2245 8565
rect 2285 8525 2295 8565
rect 2235 8500 2295 8525
rect 2235 8460 2245 8500
rect 2285 8460 2295 8500
rect 2235 8440 2295 8460
rect 2235 8400 2245 8440
rect 2285 8400 2295 8440
rect 2235 8375 2295 8400
rect 2235 8335 2245 8375
rect 2285 8335 2295 8375
rect 2235 8305 2295 8335
rect 2235 8265 2245 8305
rect 2285 8265 2295 8305
rect 2235 8235 2295 8265
rect 2235 8195 2245 8235
rect 2285 8195 2295 8235
rect 2235 8165 2295 8195
rect 2235 8125 2245 8165
rect 2285 8125 2295 8165
rect 2235 8105 2295 8125
rect 3165 9640 3225 9650
rect 3165 9600 3175 9640
rect 3215 9600 3225 9640
rect 3165 9575 3225 9600
rect 3165 9535 3175 9575
rect 3215 9535 3225 9575
rect 3165 9505 3225 9535
rect 3165 9465 3175 9505
rect 3215 9465 3225 9505
rect 3165 9435 3225 9465
rect 3165 9395 3175 9435
rect 3215 9395 3225 9435
rect 3165 9365 3225 9395
rect 3165 9325 3175 9365
rect 3215 9325 3225 9365
rect 3165 9300 3225 9325
rect 3165 9260 3175 9300
rect 3215 9260 3225 9300
rect 3165 9240 3225 9260
rect 3165 9200 3175 9240
rect 3215 9200 3225 9240
rect 3165 9175 3225 9200
rect 3165 9135 3175 9175
rect 3215 9135 3225 9175
rect 3165 9105 3225 9135
rect 3165 9065 3175 9105
rect 3215 9065 3225 9105
rect 3165 9035 3225 9065
rect 3165 8995 3175 9035
rect 3215 8995 3225 9035
rect 3165 8965 3225 8995
rect 3165 8925 3175 8965
rect 3215 8925 3225 8965
rect 3165 8900 3225 8925
rect 3165 8860 3175 8900
rect 3215 8860 3225 8900
rect 3165 8840 3225 8860
rect 3165 8800 3175 8840
rect 3215 8800 3225 8840
rect 3165 8775 3225 8800
rect 3165 8735 3175 8775
rect 3215 8735 3225 8775
rect 3165 8705 3225 8735
rect 3165 8665 3175 8705
rect 3215 8665 3225 8705
rect 3165 8635 3225 8665
rect 3165 8595 3175 8635
rect 3215 8595 3225 8635
rect 3165 8565 3225 8595
rect 3165 8525 3175 8565
rect 3215 8525 3225 8565
rect 3165 8500 3225 8525
rect 3165 8460 3175 8500
rect 3215 8460 3225 8500
rect 3165 8440 3225 8460
rect 3165 8400 3175 8440
rect 3215 8400 3225 8440
rect 3165 8375 3225 8400
rect 3165 8335 3175 8375
rect 3215 8335 3225 8375
rect 3165 8305 3225 8335
rect 3165 8265 3175 8305
rect 3215 8265 3225 8305
rect 3165 8235 3225 8265
rect 3165 8195 3175 8235
rect 3215 8195 3225 8235
rect 3165 8165 3225 8195
rect 3165 8125 3175 8165
rect 3215 8125 3225 8165
rect 3165 8105 3225 8125
rect 6690 9640 6750 9650
rect 6690 9600 6700 9640
rect 6740 9600 6750 9640
rect 6690 9575 6750 9600
rect 6690 9535 6700 9575
rect 6740 9535 6750 9575
rect 6690 9505 6750 9535
rect 6690 9465 6700 9505
rect 6740 9465 6750 9505
rect 6690 9435 6750 9465
rect 6690 9395 6700 9435
rect 6740 9395 6750 9435
rect 6690 9365 6750 9395
rect 6690 9325 6700 9365
rect 6740 9325 6750 9365
rect 6690 9300 6750 9325
rect 6690 9260 6700 9300
rect 6740 9260 6750 9300
rect 6690 9240 6750 9260
rect 6690 9200 6700 9240
rect 6740 9200 6750 9240
rect 6690 9175 6750 9200
rect 6690 9135 6700 9175
rect 6740 9135 6750 9175
rect 6690 9105 6750 9135
rect 6690 9065 6700 9105
rect 6740 9065 6750 9105
rect 6690 9035 6750 9065
rect 6690 8995 6700 9035
rect 6740 8995 6750 9035
rect 6690 8965 6750 8995
rect 6690 8925 6700 8965
rect 6740 8925 6750 8965
rect 6690 8900 6750 8925
rect 6690 8860 6700 8900
rect 6740 8860 6750 8900
rect 6690 8840 6750 8860
rect 6690 8800 6700 8840
rect 6740 8800 6750 8840
rect 6690 8775 6750 8800
rect 6690 8735 6700 8775
rect 6740 8735 6750 8775
rect 6690 8705 6750 8735
rect 6690 8665 6700 8705
rect 6740 8665 6750 8705
rect 6690 8635 6750 8665
rect 6690 8595 6700 8635
rect 6740 8595 6750 8635
rect 6690 8565 6750 8595
rect 6690 8525 6700 8565
rect 6740 8525 6750 8565
rect 6690 8500 6750 8525
rect 6690 8460 6700 8500
rect 6740 8460 6750 8500
rect 6690 8440 6750 8460
rect 6690 8400 6700 8440
rect 6740 8400 6750 8440
rect 6690 8375 6750 8400
rect 6690 8335 6700 8375
rect 6740 8335 6750 8375
rect 6690 8305 6750 8335
rect 6690 8265 6700 8305
rect 6740 8265 6750 8305
rect 6690 8235 6750 8265
rect 6690 8195 6700 8235
rect 6740 8195 6750 8235
rect 6690 8165 6750 8195
rect 6690 8125 6700 8165
rect 6740 8125 6750 8165
rect 6690 8105 6750 8125
rect 7610 9640 7670 9650
rect 7610 9600 7620 9640
rect 7660 9600 7670 9640
rect 7610 9575 7670 9600
rect 7610 9535 7620 9575
rect 7660 9535 7670 9575
rect 7610 9505 7670 9535
rect 7610 9465 7620 9505
rect 7660 9465 7670 9505
rect 7610 9435 7670 9465
rect 7610 9395 7620 9435
rect 7660 9395 7670 9435
rect 7610 9365 7670 9395
rect 7610 9325 7620 9365
rect 7660 9325 7670 9365
rect 7610 9300 7670 9325
rect 7610 9260 7620 9300
rect 7660 9260 7670 9300
rect 7610 9240 7670 9260
rect 7610 9200 7620 9240
rect 7660 9200 7670 9240
rect 7610 9175 7670 9200
rect 7610 9135 7620 9175
rect 7660 9135 7670 9175
rect 7610 9105 7670 9135
rect 7610 9065 7620 9105
rect 7660 9065 7670 9105
rect 7610 9035 7670 9065
rect 7610 8995 7620 9035
rect 7660 8995 7670 9035
rect 7610 8965 7670 8995
rect 7610 8925 7620 8965
rect 7660 8925 7670 8965
rect 7610 8900 7670 8925
rect 7610 8860 7620 8900
rect 7660 8860 7670 8900
rect 7610 8840 7670 8860
rect 7610 8800 7620 8840
rect 7660 8800 7670 8840
rect 7610 8775 7670 8800
rect 7610 8735 7620 8775
rect 7660 8735 7670 8775
rect 7610 8705 7670 8735
rect 7610 8665 7620 8705
rect 7660 8665 7670 8705
rect 7610 8635 7670 8665
rect 7610 8595 7620 8635
rect 7660 8595 7670 8635
rect 7610 8565 7670 8595
rect 7610 8525 7620 8565
rect 7660 8525 7670 8565
rect 7610 8500 7670 8525
rect 7610 8460 7620 8500
rect 7660 8460 7670 8500
rect 7610 8440 7670 8460
rect 7610 8400 7620 8440
rect 7660 8400 7670 8440
rect 7610 8375 7670 8400
rect 7610 8335 7620 8375
rect 7660 8335 7670 8375
rect 7610 8305 7670 8335
rect 7610 8265 7620 8305
rect 7660 8265 7670 8305
rect 7610 8235 7670 8265
rect 7610 8195 7620 8235
rect 7660 8195 7670 8235
rect 7610 8165 7670 8195
rect 7610 8125 7620 8165
rect 7660 8125 7670 8165
rect 7610 8105 7670 8125
rect 31290 9640 31305 9675
rect 31340 9640 31350 9675
rect 31385 9640 31395 9675
rect 31430 9640 31440 9675
rect 31475 9640 31485 9675
rect 31520 9640 31530 9675
rect 31565 9640 31575 9675
rect 31610 9640 31620 9675
rect 31655 9640 31665 9675
rect 31700 9640 31710 9675
rect 31745 9640 31755 9675
rect 31790 9640 31800 9675
rect 31835 9640 31845 9675
rect 31880 9640 31890 9675
rect 31925 9640 31935 9675
rect 31970 9640 31980 9675
rect 32015 9640 32025 9675
rect 32060 9640 32070 9675
rect 32105 9640 32115 9675
rect 32150 9640 32160 9675
rect 32195 9640 32205 9675
rect 32240 9640 32250 9675
rect 32285 9640 32295 9675
rect 32330 9640 32340 9675
rect 32375 9640 32385 9675
rect 32420 9640 32430 9675
rect 32465 9640 32475 9675
rect 32510 9640 32520 9675
rect 32555 9640 32565 9675
rect 32600 9640 32610 9675
rect 32645 9640 32655 9675
rect 32690 9640 32700 9675
rect 32735 9640 32745 9675
rect 32780 9640 32790 9675
rect 32825 9640 32835 9675
rect 32870 9640 32890 9675
rect 31290 9630 32890 9640
rect 31290 9595 31305 9630
rect 31340 9595 31350 9630
rect 31385 9595 31395 9630
rect 31430 9595 31440 9630
rect 31475 9595 31485 9630
rect 31520 9595 31530 9630
rect 31565 9595 31575 9630
rect 31610 9595 31620 9630
rect 31655 9595 31665 9630
rect 31700 9595 31710 9630
rect 31745 9595 31755 9630
rect 31790 9595 31800 9630
rect 31835 9595 31845 9630
rect 31880 9595 31890 9630
rect 31925 9595 31935 9630
rect 31970 9595 31980 9630
rect 32015 9595 32025 9630
rect 32060 9595 32070 9630
rect 32105 9595 32115 9630
rect 32150 9595 32160 9630
rect 32195 9595 32205 9630
rect 32240 9595 32250 9630
rect 32285 9595 32295 9630
rect 32330 9595 32340 9630
rect 32375 9595 32385 9630
rect 32420 9595 32430 9630
rect 32465 9595 32475 9630
rect 32510 9595 32520 9630
rect 32555 9595 32565 9630
rect 32600 9595 32610 9630
rect 32645 9595 32655 9630
rect 32690 9595 32700 9630
rect 32735 9595 32745 9630
rect 32780 9595 32790 9630
rect 32825 9595 32835 9630
rect 32870 9595 32890 9630
rect 31290 9585 32890 9595
rect 31290 9550 31305 9585
rect 31340 9550 31350 9585
rect 31385 9550 31395 9585
rect 31430 9550 31440 9585
rect 31475 9550 31485 9585
rect 31520 9550 31530 9585
rect 31565 9550 31575 9585
rect 31610 9550 31620 9585
rect 31655 9550 31665 9585
rect 31700 9550 31710 9585
rect 31745 9550 31755 9585
rect 31790 9550 31800 9585
rect 31835 9550 31845 9585
rect 31880 9550 31890 9585
rect 31925 9550 31935 9585
rect 31970 9550 31980 9585
rect 32015 9550 32025 9585
rect 32060 9550 32070 9585
rect 32105 9550 32115 9585
rect 32150 9550 32160 9585
rect 32195 9550 32205 9585
rect 32240 9550 32250 9585
rect 32285 9550 32295 9585
rect 32330 9550 32340 9585
rect 32375 9550 32385 9585
rect 32420 9550 32430 9585
rect 32465 9550 32475 9585
rect 32510 9550 32520 9585
rect 32555 9550 32565 9585
rect 32600 9550 32610 9585
rect 32645 9550 32655 9585
rect 32690 9550 32700 9585
rect 32735 9550 32745 9585
rect 32780 9550 32790 9585
rect 32825 9550 32835 9585
rect 32870 9550 32890 9585
rect 31290 9540 32890 9550
rect 31290 9505 31305 9540
rect 31340 9505 31350 9540
rect 31385 9505 31395 9540
rect 31430 9505 31440 9540
rect 31475 9505 31485 9540
rect 31520 9505 31530 9540
rect 31565 9505 31575 9540
rect 31610 9505 31620 9540
rect 31655 9505 31665 9540
rect 31700 9505 31710 9540
rect 31745 9505 31755 9540
rect 31790 9505 31800 9540
rect 31835 9505 31845 9540
rect 31880 9505 31890 9540
rect 31925 9505 31935 9540
rect 31970 9505 31980 9540
rect 32015 9505 32025 9540
rect 32060 9505 32070 9540
rect 32105 9505 32115 9540
rect 32150 9505 32160 9540
rect 32195 9505 32205 9540
rect 32240 9505 32250 9540
rect 32285 9505 32295 9540
rect 32330 9505 32340 9540
rect 32375 9505 32385 9540
rect 32420 9505 32430 9540
rect 32465 9505 32475 9540
rect 32510 9505 32520 9540
rect 32555 9505 32565 9540
rect 32600 9505 32610 9540
rect 32645 9505 32655 9540
rect 32690 9505 32700 9540
rect 32735 9505 32745 9540
rect 32780 9505 32790 9540
rect 32825 9505 32835 9540
rect 32870 9505 32890 9540
rect 31290 9495 32890 9505
rect 31290 9460 31305 9495
rect 31340 9460 31350 9495
rect 31385 9460 31395 9495
rect 31430 9460 31440 9495
rect 31475 9460 31485 9495
rect 31520 9460 31530 9495
rect 31565 9460 31575 9495
rect 31610 9460 31620 9495
rect 31655 9460 31665 9495
rect 31700 9460 31710 9495
rect 31745 9460 31755 9495
rect 31790 9460 31800 9495
rect 31835 9460 31845 9495
rect 31880 9460 31890 9495
rect 31925 9460 31935 9495
rect 31970 9460 31980 9495
rect 32015 9460 32025 9495
rect 32060 9460 32070 9495
rect 32105 9460 32115 9495
rect 32150 9460 32160 9495
rect 32195 9460 32205 9495
rect 32240 9460 32250 9495
rect 32285 9460 32295 9495
rect 32330 9460 32340 9495
rect 32375 9460 32385 9495
rect 32420 9460 32430 9495
rect 32465 9460 32475 9495
rect 32510 9460 32520 9495
rect 32555 9460 32565 9495
rect 32600 9460 32610 9495
rect 32645 9460 32655 9495
rect 32690 9460 32700 9495
rect 32735 9460 32745 9495
rect 32780 9460 32790 9495
rect 32825 9460 32835 9495
rect 32870 9460 32890 9495
rect 31290 9450 32890 9460
rect 31290 9415 31305 9450
rect 31340 9415 31350 9450
rect 31385 9415 31395 9450
rect 31430 9415 31440 9450
rect 31475 9415 31485 9450
rect 31520 9415 31530 9450
rect 31565 9415 31575 9450
rect 31610 9415 31620 9450
rect 31655 9415 31665 9450
rect 31700 9415 31710 9450
rect 31745 9415 31755 9450
rect 31790 9415 31800 9450
rect 31835 9415 31845 9450
rect 31880 9415 31890 9450
rect 31925 9415 31935 9450
rect 31970 9415 31980 9450
rect 32015 9415 32025 9450
rect 32060 9415 32070 9450
rect 32105 9415 32115 9450
rect 32150 9415 32160 9450
rect 32195 9415 32205 9450
rect 32240 9415 32250 9450
rect 32285 9415 32295 9450
rect 32330 9415 32340 9450
rect 32375 9415 32385 9450
rect 32420 9415 32430 9450
rect 32465 9415 32475 9450
rect 32510 9415 32520 9450
rect 32555 9415 32565 9450
rect 32600 9415 32610 9450
rect 32645 9415 32655 9450
rect 32690 9415 32700 9450
rect 32735 9415 32745 9450
rect 32780 9415 32790 9450
rect 32825 9415 32835 9450
rect 32870 9415 32890 9450
rect 31290 9405 32890 9415
rect 31290 9370 31305 9405
rect 31340 9370 31350 9405
rect 31385 9370 31395 9405
rect 31430 9370 31440 9405
rect 31475 9370 31485 9405
rect 31520 9370 31530 9405
rect 31565 9370 31575 9405
rect 31610 9370 31620 9405
rect 31655 9370 31665 9405
rect 31700 9370 31710 9405
rect 31745 9370 31755 9405
rect 31790 9370 31800 9405
rect 31835 9370 31845 9405
rect 31880 9370 31890 9405
rect 31925 9370 31935 9405
rect 31970 9370 31980 9405
rect 32015 9370 32025 9405
rect 32060 9370 32070 9405
rect 32105 9370 32115 9405
rect 32150 9370 32160 9405
rect 32195 9370 32205 9405
rect 32240 9370 32250 9405
rect 32285 9370 32295 9405
rect 32330 9370 32340 9405
rect 32375 9370 32385 9405
rect 32420 9370 32430 9405
rect 32465 9370 32475 9405
rect 32510 9370 32520 9405
rect 32555 9370 32565 9405
rect 32600 9370 32610 9405
rect 32645 9370 32655 9405
rect 32690 9370 32700 9405
rect 32735 9370 32745 9405
rect 32780 9370 32790 9405
rect 32825 9370 32835 9405
rect 32870 9370 32890 9405
rect 31290 9360 32890 9370
rect 31290 9325 31305 9360
rect 31340 9325 31350 9360
rect 31385 9325 31395 9360
rect 31430 9325 31440 9360
rect 31475 9325 31485 9360
rect 31520 9325 31530 9360
rect 31565 9325 31575 9360
rect 31610 9325 31620 9360
rect 31655 9325 31665 9360
rect 31700 9325 31710 9360
rect 31745 9325 31755 9360
rect 31790 9325 31800 9360
rect 31835 9325 31845 9360
rect 31880 9325 31890 9360
rect 31925 9325 31935 9360
rect 31970 9325 31980 9360
rect 32015 9325 32025 9360
rect 32060 9325 32070 9360
rect 32105 9325 32115 9360
rect 32150 9325 32160 9360
rect 32195 9325 32205 9360
rect 32240 9325 32250 9360
rect 32285 9325 32295 9360
rect 32330 9325 32340 9360
rect 32375 9325 32385 9360
rect 32420 9325 32430 9360
rect 32465 9325 32475 9360
rect 32510 9325 32520 9360
rect 32555 9325 32565 9360
rect 32600 9325 32610 9360
rect 32645 9325 32655 9360
rect 32690 9325 32700 9360
rect 32735 9325 32745 9360
rect 32780 9325 32790 9360
rect 32825 9325 32835 9360
rect 32870 9325 32890 9360
rect 31290 9315 32890 9325
rect 31290 9280 31305 9315
rect 31340 9280 31350 9315
rect 31385 9280 31395 9315
rect 31430 9280 31440 9315
rect 31475 9280 31485 9315
rect 31520 9280 31530 9315
rect 31565 9280 31575 9315
rect 31610 9280 31620 9315
rect 31655 9280 31665 9315
rect 31700 9280 31710 9315
rect 31745 9280 31755 9315
rect 31790 9280 31800 9315
rect 31835 9280 31845 9315
rect 31880 9280 31890 9315
rect 31925 9280 31935 9315
rect 31970 9280 31980 9315
rect 32015 9280 32025 9315
rect 32060 9280 32070 9315
rect 32105 9280 32115 9315
rect 32150 9280 32160 9315
rect 32195 9280 32205 9315
rect 32240 9280 32250 9315
rect 32285 9280 32295 9315
rect 32330 9280 32340 9315
rect 32375 9280 32385 9315
rect 32420 9280 32430 9315
rect 32465 9280 32475 9315
rect 32510 9280 32520 9315
rect 32555 9280 32565 9315
rect 32600 9280 32610 9315
rect 32645 9280 32655 9315
rect 32690 9280 32700 9315
rect 32735 9280 32745 9315
rect 32780 9280 32790 9315
rect 32825 9280 32835 9315
rect 32870 9280 32890 9315
rect 31290 9270 32890 9280
rect 31290 9235 31305 9270
rect 31340 9235 31350 9270
rect 31385 9235 31395 9270
rect 31430 9235 31440 9270
rect 31475 9235 31485 9270
rect 31520 9235 31530 9270
rect 31565 9235 31575 9270
rect 31610 9235 31620 9270
rect 31655 9235 31665 9270
rect 31700 9235 31710 9270
rect 31745 9235 31755 9270
rect 31790 9235 31800 9270
rect 31835 9235 31845 9270
rect 31880 9235 31890 9270
rect 31925 9235 31935 9270
rect 31970 9235 31980 9270
rect 32015 9235 32025 9270
rect 32060 9235 32070 9270
rect 32105 9235 32115 9270
rect 32150 9235 32160 9270
rect 32195 9235 32205 9270
rect 32240 9235 32250 9270
rect 32285 9235 32295 9270
rect 32330 9235 32340 9270
rect 32375 9235 32385 9270
rect 32420 9235 32430 9270
rect 32465 9235 32475 9270
rect 32510 9235 32520 9270
rect 32555 9235 32565 9270
rect 32600 9235 32610 9270
rect 32645 9235 32655 9270
rect 32690 9235 32700 9270
rect 32735 9235 32745 9270
rect 32780 9235 32790 9270
rect 32825 9235 32835 9270
rect 32870 9235 32890 9270
rect 31290 9225 32890 9235
rect 31290 9190 31305 9225
rect 31340 9190 31350 9225
rect 31385 9190 31395 9225
rect 31430 9190 31440 9225
rect 31475 9190 31485 9225
rect 31520 9190 31530 9225
rect 31565 9190 31575 9225
rect 31610 9190 31620 9225
rect 31655 9190 31665 9225
rect 31700 9190 31710 9225
rect 31745 9190 31755 9225
rect 31790 9190 31800 9225
rect 31835 9190 31845 9225
rect 31880 9190 31890 9225
rect 31925 9190 31935 9225
rect 31970 9190 31980 9225
rect 32015 9190 32025 9225
rect 32060 9190 32070 9225
rect 32105 9190 32115 9225
rect 32150 9190 32160 9225
rect 32195 9190 32205 9225
rect 32240 9190 32250 9225
rect 32285 9190 32295 9225
rect 32330 9190 32340 9225
rect 32375 9190 32385 9225
rect 32420 9190 32430 9225
rect 32465 9190 32475 9225
rect 32510 9190 32520 9225
rect 32555 9190 32565 9225
rect 32600 9190 32610 9225
rect 32645 9190 32655 9225
rect 32690 9190 32700 9225
rect 32735 9190 32745 9225
rect 32780 9190 32790 9225
rect 32825 9190 32835 9225
rect 32870 9190 32890 9225
rect 31290 9180 32890 9190
rect 31290 9145 31305 9180
rect 31340 9145 31350 9180
rect 31385 9145 31395 9180
rect 31430 9145 31440 9180
rect 31475 9145 31485 9180
rect 31520 9145 31530 9180
rect 31565 9145 31575 9180
rect 31610 9145 31620 9180
rect 31655 9145 31665 9180
rect 31700 9145 31710 9180
rect 31745 9145 31755 9180
rect 31790 9145 31800 9180
rect 31835 9145 31845 9180
rect 31880 9145 31890 9180
rect 31925 9145 31935 9180
rect 31970 9145 31980 9180
rect 32015 9145 32025 9180
rect 32060 9145 32070 9180
rect 32105 9145 32115 9180
rect 32150 9145 32160 9180
rect 32195 9145 32205 9180
rect 32240 9145 32250 9180
rect 32285 9145 32295 9180
rect 32330 9145 32340 9180
rect 32375 9145 32385 9180
rect 32420 9145 32430 9180
rect 32465 9145 32475 9180
rect 32510 9145 32520 9180
rect 32555 9145 32565 9180
rect 32600 9145 32610 9180
rect 32645 9145 32655 9180
rect 32690 9145 32700 9180
rect 32735 9145 32745 9180
rect 32780 9145 32790 9180
rect 32825 9145 32835 9180
rect 32870 9145 32890 9180
rect 31290 9135 32890 9145
rect 31290 9100 31305 9135
rect 31340 9100 31350 9135
rect 31385 9100 31395 9135
rect 31430 9100 31440 9135
rect 31475 9100 31485 9135
rect 31520 9100 31530 9135
rect 31565 9100 31575 9135
rect 31610 9100 31620 9135
rect 31655 9100 31665 9135
rect 31700 9100 31710 9135
rect 31745 9100 31755 9135
rect 31790 9100 31800 9135
rect 31835 9100 31845 9135
rect 31880 9100 31890 9135
rect 31925 9100 31935 9135
rect 31970 9100 31980 9135
rect 32015 9100 32025 9135
rect 32060 9100 32070 9135
rect 32105 9100 32115 9135
rect 32150 9100 32160 9135
rect 32195 9100 32205 9135
rect 32240 9100 32250 9135
rect 32285 9100 32295 9135
rect 32330 9100 32340 9135
rect 32375 9100 32385 9135
rect 32420 9100 32430 9135
rect 32465 9100 32475 9135
rect 32510 9100 32520 9135
rect 32555 9100 32565 9135
rect 32600 9100 32610 9135
rect 32645 9100 32655 9135
rect 32690 9100 32700 9135
rect 32735 9100 32745 9135
rect 32780 9100 32790 9135
rect 32825 9100 32835 9135
rect 32870 9100 32890 9135
rect 31290 9090 32890 9100
rect 31290 9055 31305 9090
rect 31340 9055 31350 9090
rect 31385 9055 31395 9090
rect 31430 9055 31440 9090
rect 31475 9055 31485 9090
rect 31520 9055 31530 9090
rect 31565 9055 31575 9090
rect 31610 9055 31620 9090
rect 31655 9055 31665 9090
rect 31700 9055 31710 9090
rect 31745 9055 31755 9090
rect 31790 9055 31800 9090
rect 31835 9055 31845 9090
rect 31880 9055 31890 9090
rect 31925 9055 31935 9090
rect 31970 9055 31980 9090
rect 32015 9055 32025 9090
rect 32060 9055 32070 9090
rect 32105 9055 32115 9090
rect 32150 9055 32160 9090
rect 32195 9055 32205 9090
rect 32240 9055 32250 9090
rect 32285 9055 32295 9090
rect 32330 9055 32340 9090
rect 32375 9055 32385 9090
rect 32420 9055 32430 9090
rect 32465 9055 32475 9090
rect 32510 9055 32520 9090
rect 32555 9055 32565 9090
rect 32600 9055 32610 9090
rect 32645 9055 32655 9090
rect 32690 9055 32700 9090
rect 32735 9055 32745 9090
rect 32780 9055 32790 9090
rect 32825 9055 32835 9090
rect 32870 9055 32890 9090
rect 31290 9045 32890 9055
rect 31290 9010 31305 9045
rect 31340 9010 31350 9045
rect 31385 9010 31395 9045
rect 31430 9010 31440 9045
rect 31475 9010 31485 9045
rect 31520 9010 31530 9045
rect 31565 9010 31575 9045
rect 31610 9010 31620 9045
rect 31655 9010 31665 9045
rect 31700 9010 31710 9045
rect 31745 9010 31755 9045
rect 31790 9010 31800 9045
rect 31835 9010 31845 9045
rect 31880 9010 31890 9045
rect 31925 9010 31935 9045
rect 31970 9010 31980 9045
rect 32015 9010 32025 9045
rect 32060 9010 32070 9045
rect 32105 9010 32115 9045
rect 32150 9010 32160 9045
rect 32195 9010 32205 9045
rect 32240 9010 32250 9045
rect 32285 9010 32295 9045
rect 32330 9010 32340 9045
rect 32375 9010 32385 9045
rect 32420 9010 32430 9045
rect 32465 9010 32475 9045
rect 32510 9010 32520 9045
rect 32555 9010 32565 9045
rect 32600 9010 32610 9045
rect 32645 9010 32655 9045
rect 32690 9010 32700 9045
rect 32735 9010 32745 9045
rect 32780 9010 32790 9045
rect 32825 9010 32835 9045
rect 32870 9010 32890 9045
rect 31290 9000 32890 9010
rect 31290 8965 31305 9000
rect 31340 8965 31350 9000
rect 31385 8965 31395 9000
rect 31430 8965 31440 9000
rect 31475 8965 31485 9000
rect 31520 8965 31530 9000
rect 31565 8965 31575 9000
rect 31610 8965 31620 9000
rect 31655 8965 31665 9000
rect 31700 8965 31710 9000
rect 31745 8965 31755 9000
rect 31790 8965 31800 9000
rect 31835 8965 31845 9000
rect 31880 8965 31890 9000
rect 31925 8965 31935 9000
rect 31970 8965 31980 9000
rect 32015 8965 32025 9000
rect 32060 8965 32070 9000
rect 32105 8965 32115 9000
rect 32150 8965 32160 9000
rect 32195 8965 32205 9000
rect 32240 8965 32250 9000
rect 32285 8965 32295 9000
rect 32330 8965 32340 9000
rect 32375 8965 32385 9000
rect 32420 8965 32430 9000
rect 32465 8965 32475 9000
rect 32510 8965 32520 9000
rect 32555 8965 32565 9000
rect 32600 8965 32610 9000
rect 32645 8965 32655 9000
rect 32690 8965 32700 9000
rect 32735 8965 32745 9000
rect 32780 8965 32790 9000
rect 32825 8965 32835 9000
rect 32870 8965 32890 9000
rect -90 230 -30 240
rect -90 190 -80 230
rect -40 190 -30 230
rect -90 165 -30 190
rect -90 125 -80 165
rect -40 125 -30 165
rect -90 95 -30 125
rect -90 55 -80 95
rect -40 55 -30 95
rect -90 25 -30 55
rect -90 -15 -80 25
rect -40 -15 -30 25
rect -90 -45 -30 -15
rect -90 -85 -80 -45
rect -40 -85 -30 -45
rect -90 -110 -30 -85
rect -90 -150 -80 -110
rect -40 -150 -30 -110
rect -90 -170 -30 -150
rect -90 -210 -80 -170
rect -40 -210 -30 -170
rect -90 -235 -30 -210
rect -90 -275 -80 -235
rect -40 -275 -30 -235
rect -90 -305 -30 -275
rect -90 -345 -80 -305
rect -40 -345 -30 -305
rect -90 -375 -30 -345
rect -90 -415 -80 -375
rect -40 -415 -30 -375
rect -90 -445 -30 -415
rect -90 -485 -80 -445
rect -40 -485 -30 -445
rect -90 -510 -30 -485
rect -90 -550 -80 -510
rect -40 -550 -30 -510
rect -90 -570 -30 -550
rect -90 -610 -80 -570
rect -40 -610 -30 -570
rect -90 -635 -30 -610
rect -90 -675 -80 -635
rect -40 -675 -30 -635
rect -90 -705 -30 -675
rect -90 -745 -80 -705
rect -40 -745 -30 -705
rect -90 -775 -30 -745
rect -90 -815 -80 -775
rect -40 -815 -30 -775
rect -90 -845 -30 -815
rect -90 -885 -80 -845
rect -40 -885 -30 -845
rect -90 -910 -30 -885
rect -90 -950 -80 -910
rect -40 -950 -30 -910
rect -90 -970 -30 -950
rect -90 -1010 -80 -970
rect -40 -1010 -30 -970
rect -90 -1035 -30 -1010
rect -90 -1075 -80 -1035
rect -40 -1075 -30 -1035
rect -90 -1105 -30 -1075
rect -90 -1145 -80 -1105
rect -40 -1145 -30 -1105
rect -90 -1175 -30 -1145
rect -90 -1215 -80 -1175
rect -40 -1215 -30 -1175
rect -90 -1245 -30 -1215
rect -90 -1285 -80 -1245
rect -40 -1285 -30 -1245
rect -90 -1310 -30 -1285
rect -90 -1350 -80 -1310
rect -40 -1350 -30 -1310
rect -90 -1360 -30 -1350
rect 260 230 320 240
rect 260 190 270 230
rect 310 190 320 230
rect 260 165 320 190
rect 260 125 270 165
rect 310 125 320 165
rect 260 95 320 125
rect 260 55 270 95
rect 310 55 320 95
rect 260 25 320 55
rect 260 -15 270 25
rect 310 -15 320 25
rect 260 -45 320 -15
rect 260 -85 270 -45
rect 310 -85 320 -45
rect 260 -110 320 -85
rect 260 -150 270 -110
rect 310 -150 320 -110
rect 260 -170 320 -150
rect 260 -210 270 -170
rect 310 -210 320 -170
rect 260 -235 320 -210
rect 260 -275 270 -235
rect 310 -275 320 -235
rect 260 -305 320 -275
rect 260 -345 270 -305
rect 310 -345 320 -305
rect 260 -375 320 -345
rect 260 -415 270 -375
rect 310 -415 320 -375
rect 260 -445 320 -415
rect 260 -485 270 -445
rect 310 -485 320 -445
rect 260 -510 320 -485
rect 260 -550 270 -510
rect 310 -550 320 -510
rect 260 -570 320 -550
rect 260 -610 270 -570
rect 310 -610 320 -570
rect 260 -635 320 -610
rect 260 -675 270 -635
rect 310 -675 320 -635
rect 260 -705 320 -675
rect 260 -745 270 -705
rect 310 -745 320 -705
rect 260 -775 320 -745
rect 260 -815 270 -775
rect 310 -815 320 -775
rect 260 -845 320 -815
rect 260 -885 270 -845
rect 310 -885 320 -845
rect 260 -910 320 -885
rect 260 -950 270 -910
rect 310 -950 320 -910
rect 260 -970 320 -950
rect 260 -1010 270 -970
rect 310 -1010 320 -970
rect 260 -1035 320 -1010
rect 260 -1075 270 -1035
rect 310 -1075 320 -1035
rect 260 -1105 320 -1075
rect 260 -1145 270 -1105
rect 310 -1145 320 -1105
rect 260 -1175 320 -1145
rect 260 -1215 270 -1175
rect 310 -1215 320 -1175
rect 260 -1245 320 -1215
rect 260 -1285 270 -1245
rect 310 -1285 320 -1245
rect 260 -1310 320 -1285
rect 260 -1350 270 -1310
rect 310 -1350 320 -1310
rect 260 -1360 320 -1350
rect 610 230 670 240
rect 610 190 620 230
rect 660 190 670 230
rect 610 165 670 190
rect 610 125 620 165
rect 660 125 670 165
rect 610 95 670 125
rect 610 55 620 95
rect 660 55 670 95
rect 610 25 670 55
rect 610 -15 620 25
rect 660 -15 670 25
rect 610 -45 670 -15
rect 610 -85 620 -45
rect 660 -85 670 -45
rect 610 -110 670 -85
rect 610 -150 620 -110
rect 660 -150 670 -110
rect 610 -170 670 -150
rect 610 -210 620 -170
rect 660 -210 670 -170
rect 610 -235 670 -210
rect 610 -275 620 -235
rect 660 -275 670 -235
rect 610 -305 670 -275
rect 610 -345 620 -305
rect 660 -345 670 -305
rect 610 -375 670 -345
rect 610 -415 620 -375
rect 660 -415 670 -375
rect 610 -445 670 -415
rect 610 -485 620 -445
rect 660 -485 670 -445
rect 610 -510 670 -485
rect 610 -550 620 -510
rect 660 -550 670 -510
rect 610 -570 670 -550
rect 610 -610 620 -570
rect 660 -610 670 -570
rect 610 -635 670 -610
rect 610 -675 620 -635
rect 660 -675 670 -635
rect 610 -705 670 -675
rect 610 -745 620 -705
rect 660 -745 670 -705
rect 610 -775 670 -745
rect 610 -815 620 -775
rect 660 -815 670 -775
rect 610 -845 670 -815
rect 610 -885 620 -845
rect 660 -885 670 -845
rect 610 -910 670 -885
rect 610 -950 620 -910
rect 660 -950 670 -910
rect 610 -970 670 -950
rect 610 -1010 620 -970
rect 660 -1010 670 -970
rect 610 -1035 670 -1010
rect 610 -1075 620 -1035
rect 660 -1075 670 -1035
rect 610 -1105 670 -1075
rect 610 -1145 620 -1105
rect 660 -1145 670 -1105
rect 610 -1175 670 -1145
rect 610 -1215 620 -1175
rect 660 -1215 670 -1175
rect 610 -1245 670 -1215
rect 610 -1285 620 -1245
rect 660 -1285 670 -1245
rect 610 -1310 670 -1285
rect 610 -1350 620 -1310
rect 660 -1350 670 -1310
rect 610 -1360 670 -1350
rect 960 230 1020 240
rect 960 190 970 230
rect 1010 190 1020 230
rect 960 165 1020 190
rect 960 125 970 165
rect 1010 125 1020 165
rect 960 95 1020 125
rect 960 55 970 95
rect 1010 55 1020 95
rect 960 25 1020 55
rect 960 -15 970 25
rect 1010 -15 1020 25
rect 960 -45 1020 -15
rect 960 -85 970 -45
rect 1010 -85 1020 -45
rect 960 -110 1020 -85
rect 960 -150 970 -110
rect 1010 -150 1020 -110
rect 960 -170 1020 -150
rect 960 -210 970 -170
rect 1010 -210 1020 -170
rect 960 -235 1020 -210
rect 960 -275 970 -235
rect 1010 -275 1020 -235
rect 960 -305 1020 -275
rect 960 -345 970 -305
rect 1010 -345 1020 -305
rect 960 -375 1020 -345
rect 960 -415 970 -375
rect 1010 -415 1020 -375
rect 960 -445 1020 -415
rect 960 -485 970 -445
rect 1010 -485 1020 -445
rect 960 -510 1020 -485
rect 960 -550 970 -510
rect 1010 -550 1020 -510
rect 960 -570 1020 -550
rect 960 -610 970 -570
rect 1010 -610 1020 -570
rect 960 -635 1020 -610
rect 960 -675 970 -635
rect 1010 -675 1020 -635
rect 960 -705 1020 -675
rect 960 -745 970 -705
rect 1010 -745 1020 -705
rect 960 -775 1020 -745
rect 960 -815 970 -775
rect 1010 -815 1020 -775
rect 960 -845 1020 -815
rect 960 -885 970 -845
rect 1010 -885 1020 -845
rect 960 -910 1020 -885
rect 960 -950 970 -910
rect 1010 -950 1020 -910
rect 960 -970 1020 -950
rect 960 -1010 970 -970
rect 1010 -1010 1020 -970
rect 960 -1035 1020 -1010
rect 960 -1075 970 -1035
rect 1010 -1075 1020 -1035
rect 960 -1105 1020 -1075
rect 960 -1145 970 -1105
rect 1010 -1145 1020 -1105
rect 960 -1175 1020 -1145
rect 960 -1215 970 -1175
rect 1010 -1215 1020 -1175
rect 960 -1245 1020 -1215
rect 960 -1285 970 -1245
rect 1010 -1285 1020 -1245
rect 960 -1310 1020 -1285
rect 960 -1350 970 -1310
rect 1010 -1350 1020 -1310
rect 960 -1360 1020 -1350
rect 1310 230 1370 240
rect 1310 190 1320 230
rect 1360 190 1370 230
rect 1310 165 1370 190
rect 1310 125 1320 165
rect 1360 125 1370 165
rect 1310 95 1370 125
rect 1310 55 1320 95
rect 1360 55 1370 95
rect 1310 25 1370 55
rect 1310 -15 1320 25
rect 1360 -15 1370 25
rect 1310 -45 1370 -15
rect 1310 -85 1320 -45
rect 1360 -85 1370 -45
rect 1310 -110 1370 -85
rect 1310 -150 1320 -110
rect 1360 -150 1370 -110
rect 1310 -170 1370 -150
rect 1310 -210 1320 -170
rect 1360 -210 1370 -170
rect 1310 -235 1370 -210
rect 1310 -275 1320 -235
rect 1360 -275 1370 -235
rect 1310 -305 1370 -275
rect 1310 -345 1320 -305
rect 1360 -345 1370 -305
rect 1310 -375 1370 -345
rect 1310 -415 1320 -375
rect 1360 -415 1370 -375
rect 1310 -445 1370 -415
rect 1310 -485 1320 -445
rect 1360 -485 1370 -445
rect 1310 -510 1370 -485
rect 1310 -550 1320 -510
rect 1360 -550 1370 -510
rect 1310 -570 1370 -550
rect 1310 -610 1320 -570
rect 1360 -610 1370 -570
rect 1310 -635 1370 -610
rect 1310 -675 1320 -635
rect 1360 -675 1370 -635
rect 1310 -705 1370 -675
rect 1310 -745 1320 -705
rect 1360 -745 1370 -705
rect 1310 -775 1370 -745
rect 1310 -815 1320 -775
rect 1360 -815 1370 -775
rect 1310 -845 1370 -815
rect 1310 -885 1320 -845
rect 1360 -885 1370 -845
rect 1310 -910 1370 -885
rect 1310 -950 1320 -910
rect 1360 -950 1370 -910
rect 1310 -970 1370 -950
rect 1310 -1010 1320 -970
rect 1360 -1010 1370 -970
rect 1310 -1035 1370 -1010
rect 1310 -1075 1320 -1035
rect 1360 -1075 1370 -1035
rect 1310 -1105 1370 -1075
rect 1310 -1145 1320 -1105
rect 1360 -1145 1370 -1105
rect 1310 -1175 1370 -1145
rect 1310 -1215 1320 -1175
rect 1360 -1215 1370 -1175
rect 1310 -1245 1370 -1215
rect 1310 -1285 1320 -1245
rect 1360 -1285 1370 -1245
rect 1310 -1310 1370 -1285
rect 1310 -1350 1320 -1310
rect 1360 -1350 1370 -1310
rect 1310 -1360 1370 -1350
rect 1660 230 1720 240
rect 1660 190 1670 230
rect 1710 190 1720 230
rect 1660 165 1720 190
rect 1660 125 1670 165
rect 1710 125 1720 165
rect 1660 95 1720 125
rect 1660 55 1670 95
rect 1710 55 1720 95
rect 1660 25 1720 55
rect 1660 -15 1670 25
rect 1710 -15 1720 25
rect 1660 -45 1720 -15
rect 1660 -85 1670 -45
rect 1710 -85 1720 -45
rect 1660 -110 1720 -85
rect 1660 -150 1670 -110
rect 1710 -150 1720 -110
rect 1660 -170 1720 -150
rect 1660 -210 1670 -170
rect 1710 -210 1720 -170
rect 1660 -235 1720 -210
rect 1660 -275 1670 -235
rect 1710 -275 1720 -235
rect 1660 -305 1720 -275
rect 1660 -345 1670 -305
rect 1710 -345 1720 -305
rect 1660 -375 1720 -345
rect 1660 -415 1670 -375
rect 1710 -415 1720 -375
rect 1660 -445 1720 -415
rect 1660 -485 1670 -445
rect 1710 -485 1720 -445
rect 1660 -510 1720 -485
rect 1660 -550 1670 -510
rect 1710 -550 1720 -510
rect 1660 -570 1720 -550
rect 1660 -610 1670 -570
rect 1710 -610 1720 -570
rect 1660 -635 1720 -610
rect 1660 -675 1670 -635
rect 1710 -675 1720 -635
rect 1660 -705 1720 -675
rect 1660 -745 1670 -705
rect 1710 -745 1720 -705
rect 1660 -775 1720 -745
rect 1660 -815 1670 -775
rect 1710 -815 1720 -775
rect 1660 -845 1720 -815
rect 1660 -885 1670 -845
rect 1710 -885 1720 -845
rect 1660 -910 1720 -885
rect 1660 -950 1670 -910
rect 1710 -950 1720 -910
rect 1660 -970 1720 -950
rect 1660 -1010 1670 -970
rect 1710 -1010 1720 -970
rect 1660 -1035 1720 -1010
rect 1660 -1075 1670 -1035
rect 1710 -1075 1720 -1035
rect 1660 -1105 1720 -1075
rect 1660 -1145 1670 -1105
rect 1710 -1145 1720 -1105
rect 1660 -1175 1720 -1145
rect 1660 -1215 1670 -1175
rect 1710 -1215 1720 -1175
rect 1660 -1245 1720 -1215
rect 1660 -1285 1670 -1245
rect 1710 -1285 1720 -1245
rect 1660 -1310 1720 -1285
rect 1660 -1350 1670 -1310
rect 1710 -1350 1720 -1310
rect 1660 -1360 1720 -1350
rect 2010 230 2070 240
rect 2010 190 2020 230
rect 2060 190 2070 230
rect 2010 165 2070 190
rect 2010 125 2020 165
rect 2060 125 2070 165
rect 2010 95 2070 125
rect 2010 55 2020 95
rect 2060 55 2070 95
rect 2010 25 2070 55
rect 2010 -15 2020 25
rect 2060 -15 2070 25
rect 2010 -45 2070 -15
rect 2010 -85 2020 -45
rect 2060 -85 2070 -45
rect 2010 -110 2070 -85
rect 2010 -150 2020 -110
rect 2060 -150 2070 -110
rect 2010 -170 2070 -150
rect 2010 -210 2020 -170
rect 2060 -210 2070 -170
rect 2010 -235 2070 -210
rect 2010 -275 2020 -235
rect 2060 -275 2070 -235
rect 2010 -305 2070 -275
rect 2010 -345 2020 -305
rect 2060 -345 2070 -305
rect 2010 -375 2070 -345
rect 2010 -415 2020 -375
rect 2060 -415 2070 -375
rect 2010 -445 2070 -415
rect 2010 -485 2020 -445
rect 2060 -485 2070 -445
rect 2010 -510 2070 -485
rect 2010 -550 2020 -510
rect 2060 -550 2070 -510
rect 2010 -570 2070 -550
rect 2010 -610 2020 -570
rect 2060 -610 2070 -570
rect 2010 -635 2070 -610
rect 2010 -675 2020 -635
rect 2060 -675 2070 -635
rect 2010 -705 2070 -675
rect 2010 -745 2020 -705
rect 2060 -745 2070 -705
rect 2010 -775 2070 -745
rect 2010 -815 2020 -775
rect 2060 -815 2070 -775
rect 2010 -845 2070 -815
rect 2010 -885 2020 -845
rect 2060 -885 2070 -845
rect 2010 -910 2070 -885
rect 2010 -950 2020 -910
rect 2060 -950 2070 -910
rect 2010 -970 2070 -950
rect 2010 -1010 2020 -970
rect 2060 -1010 2070 -970
rect 2010 -1035 2070 -1010
rect 2010 -1075 2020 -1035
rect 2060 -1075 2070 -1035
rect 2010 -1105 2070 -1075
rect 2010 -1145 2020 -1105
rect 2060 -1145 2070 -1105
rect 2010 -1175 2070 -1145
rect 2010 -1215 2020 -1175
rect 2060 -1215 2070 -1175
rect 2010 -1245 2070 -1215
rect 2010 -1285 2020 -1245
rect 2060 -1285 2070 -1245
rect 2010 -1310 2070 -1285
rect 2010 -1350 2020 -1310
rect 2060 -1350 2070 -1310
rect 2010 -1360 2070 -1350
rect 2360 230 2420 240
rect 2360 190 2370 230
rect 2410 190 2420 230
rect 2360 165 2420 190
rect 2360 125 2370 165
rect 2410 125 2420 165
rect 2360 95 2420 125
rect 2360 55 2370 95
rect 2410 55 2420 95
rect 2360 25 2420 55
rect 2360 -15 2370 25
rect 2410 -15 2420 25
rect 2360 -45 2420 -15
rect 2360 -85 2370 -45
rect 2410 -85 2420 -45
rect 2360 -110 2420 -85
rect 2360 -150 2370 -110
rect 2410 -150 2420 -110
rect 2360 -170 2420 -150
rect 2360 -210 2370 -170
rect 2410 -210 2420 -170
rect 2360 -235 2420 -210
rect 2360 -275 2370 -235
rect 2410 -275 2420 -235
rect 2360 -305 2420 -275
rect 2360 -345 2370 -305
rect 2410 -345 2420 -305
rect 2360 -375 2420 -345
rect 2360 -415 2370 -375
rect 2410 -415 2420 -375
rect 2360 -445 2420 -415
rect 2360 -485 2370 -445
rect 2410 -485 2420 -445
rect 2360 -510 2420 -485
rect 2360 -550 2370 -510
rect 2410 -550 2420 -510
rect 2360 -570 2420 -550
rect 2360 -610 2370 -570
rect 2410 -610 2420 -570
rect 2360 -635 2420 -610
rect 2360 -675 2370 -635
rect 2410 -675 2420 -635
rect 2360 -705 2420 -675
rect 2360 -745 2370 -705
rect 2410 -745 2420 -705
rect 2360 -775 2420 -745
rect 2360 -815 2370 -775
rect 2410 -815 2420 -775
rect 2360 -845 2420 -815
rect 2360 -885 2370 -845
rect 2410 -885 2420 -845
rect 2360 -910 2420 -885
rect 2360 -950 2370 -910
rect 2410 -950 2420 -910
rect 2360 -970 2420 -950
rect 2360 -1010 2370 -970
rect 2410 -1010 2420 -970
rect 2360 -1035 2420 -1010
rect 2360 -1075 2370 -1035
rect 2410 -1075 2420 -1035
rect 2360 -1105 2420 -1075
rect 2360 -1145 2370 -1105
rect 2410 -1145 2420 -1105
rect 2360 -1175 2420 -1145
rect 2360 -1215 2370 -1175
rect 2410 -1215 2420 -1175
rect 2360 -1245 2420 -1215
rect 2360 -1285 2370 -1245
rect 2410 -1285 2420 -1245
rect 2360 -1310 2420 -1285
rect 2360 -1350 2370 -1310
rect 2410 -1350 2420 -1310
rect 2360 -1360 2420 -1350
rect 2710 230 2770 240
rect 2710 190 2720 230
rect 2760 190 2770 230
rect 2710 165 2770 190
rect 2710 125 2720 165
rect 2760 125 2770 165
rect 2710 95 2770 125
rect 2710 55 2720 95
rect 2760 55 2770 95
rect 2710 25 2770 55
rect 2710 -15 2720 25
rect 2760 -15 2770 25
rect 2710 -45 2770 -15
rect 2710 -85 2720 -45
rect 2760 -85 2770 -45
rect 2710 -110 2770 -85
rect 2710 -150 2720 -110
rect 2760 -150 2770 -110
rect 2710 -170 2770 -150
rect 2710 -210 2720 -170
rect 2760 -210 2770 -170
rect 2710 -235 2770 -210
rect 2710 -275 2720 -235
rect 2760 -275 2770 -235
rect 2710 -305 2770 -275
rect 2710 -345 2720 -305
rect 2760 -345 2770 -305
rect 2710 -375 2770 -345
rect 2710 -415 2720 -375
rect 2760 -415 2770 -375
rect 2710 -445 2770 -415
rect 2710 -485 2720 -445
rect 2760 -485 2770 -445
rect 2710 -510 2770 -485
rect 2710 -550 2720 -510
rect 2760 -550 2770 -510
rect 2710 -570 2770 -550
rect 2710 -610 2720 -570
rect 2760 -610 2770 -570
rect 2710 -635 2770 -610
rect 2710 -675 2720 -635
rect 2760 -675 2770 -635
rect 2710 -705 2770 -675
rect 2710 -745 2720 -705
rect 2760 -745 2770 -705
rect 2710 -775 2770 -745
rect 2710 -815 2720 -775
rect 2760 -815 2770 -775
rect 2710 -845 2770 -815
rect 2710 -885 2720 -845
rect 2760 -885 2770 -845
rect 2710 -910 2770 -885
rect 2710 -950 2720 -910
rect 2760 -950 2770 -910
rect 2710 -970 2770 -950
rect 2710 -1010 2720 -970
rect 2760 -1010 2770 -970
rect 2710 -1035 2770 -1010
rect 2710 -1075 2720 -1035
rect 2760 -1075 2770 -1035
rect 2710 -1105 2770 -1075
rect 2710 -1145 2720 -1105
rect 2760 -1145 2770 -1105
rect 2710 -1175 2770 -1145
rect 2710 -1215 2720 -1175
rect 2760 -1215 2770 -1175
rect 2710 -1245 2770 -1215
rect 2710 -1285 2720 -1245
rect 2760 -1285 2770 -1245
rect 2710 -1310 2770 -1285
rect 2710 -1350 2720 -1310
rect 2760 -1350 2770 -1310
rect 2710 -1360 2770 -1350
rect 3060 230 3120 240
rect 3060 190 3070 230
rect 3110 190 3120 230
rect 3060 165 3120 190
rect 3060 125 3070 165
rect 3110 125 3120 165
rect 3060 95 3120 125
rect 3060 55 3070 95
rect 3110 55 3120 95
rect 3060 25 3120 55
rect 3060 -15 3070 25
rect 3110 -15 3120 25
rect 3060 -45 3120 -15
rect 3060 -85 3070 -45
rect 3110 -85 3120 -45
rect 3060 -110 3120 -85
rect 3060 -150 3070 -110
rect 3110 -150 3120 -110
rect 3060 -170 3120 -150
rect 3060 -210 3070 -170
rect 3110 -210 3120 -170
rect 3060 -235 3120 -210
rect 3060 -275 3070 -235
rect 3110 -275 3120 -235
rect 3060 -305 3120 -275
rect 3060 -345 3070 -305
rect 3110 -345 3120 -305
rect 3060 -375 3120 -345
rect 3060 -415 3070 -375
rect 3110 -415 3120 -375
rect 3060 -445 3120 -415
rect 3060 -485 3070 -445
rect 3110 -485 3120 -445
rect 3060 -510 3120 -485
rect 3060 -550 3070 -510
rect 3110 -550 3120 -510
rect 3060 -570 3120 -550
rect 3060 -610 3070 -570
rect 3110 -610 3120 -570
rect 3060 -635 3120 -610
rect 3060 -675 3070 -635
rect 3110 -675 3120 -635
rect 3060 -705 3120 -675
rect 3060 -745 3070 -705
rect 3110 -745 3120 -705
rect 3060 -775 3120 -745
rect 3060 -815 3070 -775
rect 3110 -815 3120 -775
rect 3060 -845 3120 -815
rect 3060 -885 3070 -845
rect 3110 -885 3120 -845
rect 3060 -910 3120 -885
rect 3060 -950 3070 -910
rect 3110 -950 3120 -910
rect 3060 -970 3120 -950
rect 3060 -1010 3070 -970
rect 3110 -1010 3120 -970
rect 3060 -1035 3120 -1010
rect 3060 -1075 3070 -1035
rect 3110 -1075 3120 -1035
rect 3060 -1105 3120 -1075
rect 3060 -1145 3070 -1105
rect 3110 -1145 3120 -1105
rect 3060 -1175 3120 -1145
rect 3060 -1215 3070 -1175
rect 3110 -1215 3120 -1175
rect 3060 -1245 3120 -1215
rect 3060 -1285 3070 -1245
rect 3110 -1285 3120 -1245
rect 3060 -1310 3120 -1285
rect 3060 -1350 3070 -1310
rect 3110 -1350 3120 -1310
rect 3060 -1360 3120 -1350
rect 3410 230 3470 240
rect 3410 190 3420 230
rect 3460 190 3470 230
rect 3410 165 3470 190
rect 3410 125 3420 165
rect 3460 125 3470 165
rect 3410 95 3470 125
rect 3410 55 3420 95
rect 3460 55 3470 95
rect 3410 25 3470 55
rect 3410 -15 3420 25
rect 3460 -15 3470 25
rect 3410 -45 3470 -15
rect 3410 -85 3420 -45
rect 3460 -85 3470 -45
rect 3410 -110 3470 -85
rect 3410 -150 3420 -110
rect 3460 -150 3470 -110
rect 3410 -170 3470 -150
rect 3410 -210 3420 -170
rect 3460 -210 3470 -170
rect 3410 -235 3470 -210
rect 3410 -275 3420 -235
rect 3460 -275 3470 -235
rect 3410 -305 3470 -275
rect 3410 -345 3420 -305
rect 3460 -345 3470 -305
rect 3410 -375 3470 -345
rect 3410 -415 3420 -375
rect 3460 -415 3470 -375
rect 3410 -445 3470 -415
rect 3410 -485 3420 -445
rect 3460 -485 3470 -445
rect 3410 -510 3470 -485
rect 3410 -550 3420 -510
rect 3460 -550 3470 -510
rect 3410 -570 3470 -550
rect 3410 -610 3420 -570
rect 3460 -610 3470 -570
rect 3410 -635 3470 -610
rect 3410 -675 3420 -635
rect 3460 -675 3470 -635
rect 3410 -705 3470 -675
rect 3410 -745 3420 -705
rect 3460 -745 3470 -705
rect 3410 -775 3470 -745
rect 3410 -815 3420 -775
rect 3460 -815 3470 -775
rect 3410 -845 3470 -815
rect 3410 -885 3420 -845
rect 3460 -885 3470 -845
rect 3410 -910 3470 -885
rect 3410 -950 3420 -910
rect 3460 -950 3470 -910
rect 3410 -970 3470 -950
rect 3410 -1010 3420 -970
rect 3460 -1010 3470 -970
rect 3410 -1035 3470 -1010
rect 3410 -1075 3420 -1035
rect 3460 -1075 3470 -1035
rect 3410 -1105 3470 -1075
rect 3410 -1145 3420 -1105
rect 3460 -1145 3470 -1105
rect 3410 -1175 3470 -1145
rect 3410 -1215 3420 -1175
rect 3460 -1215 3470 -1175
rect 3410 -1245 3470 -1215
rect 3410 -1285 3420 -1245
rect 3460 -1285 3470 -1245
rect 3410 -1310 3470 -1285
rect 3410 -1350 3420 -1310
rect 3460 -1350 3470 -1310
rect 3410 -1360 3470 -1350
rect 3760 230 3820 240
rect 3760 190 3770 230
rect 3810 190 3820 230
rect 3760 165 3820 190
rect 3760 125 3770 165
rect 3810 125 3820 165
rect 3760 95 3820 125
rect 3760 55 3770 95
rect 3810 55 3820 95
rect 3760 25 3820 55
rect 3760 -15 3770 25
rect 3810 -15 3820 25
rect 3760 -45 3820 -15
rect 3760 -85 3770 -45
rect 3810 -85 3820 -45
rect 3760 -110 3820 -85
rect 3760 -150 3770 -110
rect 3810 -150 3820 -110
rect 3760 -170 3820 -150
rect 3760 -210 3770 -170
rect 3810 -210 3820 -170
rect 3760 -235 3820 -210
rect 3760 -275 3770 -235
rect 3810 -275 3820 -235
rect 3760 -305 3820 -275
rect 3760 -345 3770 -305
rect 3810 -345 3820 -305
rect 3760 -375 3820 -345
rect 3760 -415 3770 -375
rect 3810 -415 3820 -375
rect 3760 -445 3820 -415
rect 3760 -485 3770 -445
rect 3810 -485 3820 -445
rect 3760 -510 3820 -485
rect 3760 -550 3770 -510
rect 3810 -550 3820 -510
rect 3760 -570 3820 -550
rect 3760 -610 3770 -570
rect 3810 -610 3820 -570
rect 3760 -635 3820 -610
rect 3760 -675 3770 -635
rect 3810 -675 3820 -635
rect 3760 -705 3820 -675
rect 3760 -745 3770 -705
rect 3810 -745 3820 -705
rect 3760 -775 3820 -745
rect 3760 -815 3770 -775
rect 3810 -815 3820 -775
rect 3760 -845 3820 -815
rect 3760 -885 3770 -845
rect 3810 -885 3820 -845
rect 3760 -910 3820 -885
rect 3760 -950 3770 -910
rect 3810 -950 3820 -910
rect 3760 -970 3820 -950
rect 3760 -1010 3770 -970
rect 3810 -1010 3820 -970
rect 3760 -1035 3820 -1010
rect 3760 -1075 3770 -1035
rect 3810 -1075 3820 -1035
rect 3760 -1105 3820 -1075
rect 3760 -1145 3770 -1105
rect 3810 -1145 3820 -1105
rect 3760 -1175 3820 -1145
rect 3760 -1215 3770 -1175
rect 3810 -1215 3820 -1175
rect 3760 -1245 3820 -1215
rect 3760 -1285 3770 -1245
rect 3810 -1285 3820 -1245
rect 3760 -1310 3820 -1285
rect 3760 -1350 3770 -1310
rect 3810 -1350 3820 -1310
rect 3760 -1360 3820 -1350
rect 4110 230 4170 240
rect 4110 190 4120 230
rect 4160 190 4170 230
rect 4110 165 4170 190
rect 4110 125 4120 165
rect 4160 125 4170 165
rect 4110 95 4170 125
rect 4110 55 4120 95
rect 4160 55 4170 95
rect 4110 25 4170 55
rect 4110 -15 4120 25
rect 4160 -15 4170 25
rect 4110 -45 4170 -15
rect 4110 -85 4120 -45
rect 4160 -85 4170 -45
rect 4110 -110 4170 -85
rect 4110 -150 4120 -110
rect 4160 -150 4170 -110
rect 4110 -170 4170 -150
rect 4110 -210 4120 -170
rect 4160 -210 4170 -170
rect 4110 -235 4170 -210
rect 4110 -275 4120 -235
rect 4160 -275 4170 -235
rect 4110 -305 4170 -275
rect 4110 -345 4120 -305
rect 4160 -345 4170 -305
rect 4110 -375 4170 -345
rect 4110 -415 4120 -375
rect 4160 -415 4170 -375
rect 4110 -445 4170 -415
rect 4110 -485 4120 -445
rect 4160 -485 4170 -445
rect 4110 -510 4170 -485
rect 4110 -550 4120 -510
rect 4160 -550 4170 -510
rect 4110 -570 4170 -550
rect 4110 -610 4120 -570
rect 4160 -610 4170 -570
rect 4110 -635 4170 -610
rect 4110 -675 4120 -635
rect 4160 -675 4170 -635
rect 4110 -705 4170 -675
rect 4110 -745 4120 -705
rect 4160 -745 4170 -705
rect 4110 -775 4170 -745
rect 4110 -815 4120 -775
rect 4160 -815 4170 -775
rect 4110 -845 4170 -815
rect 4110 -885 4120 -845
rect 4160 -885 4170 -845
rect 4110 -910 4170 -885
rect 4110 -950 4120 -910
rect 4160 -950 4170 -910
rect 4110 -970 4170 -950
rect 4110 -1010 4120 -970
rect 4160 -1010 4170 -970
rect 4110 -1035 4170 -1010
rect 4110 -1075 4120 -1035
rect 4160 -1075 4170 -1035
rect 4110 -1105 4170 -1075
rect 4110 -1145 4120 -1105
rect 4160 -1145 4170 -1105
rect 4110 -1175 4170 -1145
rect 4110 -1215 4120 -1175
rect 4160 -1215 4170 -1175
rect 4110 -1245 4170 -1215
rect 4110 -1285 4120 -1245
rect 4160 -1285 4170 -1245
rect 4110 -1310 4170 -1285
rect 4110 -1350 4120 -1310
rect 4160 -1350 4170 -1310
rect 4110 -1360 4170 -1350
rect 4460 230 4520 240
rect 4460 190 4470 230
rect 4510 190 4520 230
rect 4460 165 4520 190
rect 4460 125 4470 165
rect 4510 125 4520 165
rect 4460 95 4520 125
rect 4460 55 4470 95
rect 4510 55 4520 95
rect 4460 25 4520 55
rect 4460 -15 4470 25
rect 4510 -15 4520 25
rect 4460 -45 4520 -15
rect 4460 -85 4470 -45
rect 4510 -85 4520 -45
rect 4460 -110 4520 -85
rect 4460 -150 4470 -110
rect 4510 -150 4520 -110
rect 4460 -170 4520 -150
rect 4460 -210 4470 -170
rect 4510 -210 4520 -170
rect 4460 -235 4520 -210
rect 4460 -275 4470 -235
rect 4510 -275 4520 -235
rect 4460 -305 4520 -275
rect 4460 -345 4470 -305
rect 4510 -345 4520 -305
rect 4460 -375 4520 -345
rect 4460 -415 4470 -375
rect 4510 -415 4520 -375
rect 4460 -445 4520 -415
rect 4460 -485 4470 -445
rect 4510 -485 4520 -445
rect 4460 -510 4520 -485
rect 4460 -550 4470 -510
rect 4510 -550 4520 -510
rect 4460 -570 4520 -550
rect 4460 -610 4470 -570
rect 4510 -610 4520 -570
rect 4460 -635 4520 -610
rect 4460 -675 4470 -635
rect 4510 -675 4520 -635
rect 4460 -705 4520 -675
rect 4460 -745 4470 -705
rect 4510 -745 4520 -705
rect 4460 -775 4520 -745
rect 4460 -815 4470 -775
rect 4510 -815 4520 -775
rect 4460 -845 4520 -815
rect 4460 -885 4470 -845
rect 4510 -885 4520 -845
rect 4460 -910 4520 -885
rect 4460 -950 4470 -910
rect 4510 -950 4520 -910
rect 4460 -970 4520 -950
rect 4460 -1010 4470 -970
rect 4510 -1010 4520 -970
rect 4460 -1035 4520 -1010
rect 4460 -1075 4470 -1035
rect 4510 -1075 4520 -1035
rect 4460 -1105 4520 -1075
rect 4460 -1145 4470 -1105
rect 4510 -1145 4520 -1105
rect 4460 -1175 4520 -1145
rect 4460 -1215 4470 -1175
rect 4510 -1215 4520 -1175
rect 4460 -1245 4520 -1215
rect 4460 -1285 4470 -1245
rect 4510 -1285 4520 -1245
rect 4460 -1310 4520 -1285
rect 4460 -1350 4470 -1310
rect 4510 -1350 4520 -1310
rect 4460 -1360 4520 -1350
rect 4810 230 4870 240
rect 4810 190 4820 230
rect 4860 190 4870 230
rect 4810 165 4870 190
rect 4810 125 4820 165
rect 4860 125 4870 165
rect 4810 95 4870 125
rect 4810 55 4820 95
rect 4860 55 4870 95
rect 4810 25 4870 55
rect 4810 -15 4820 25
rect 4860 -15 4870 25
rect 4810 -45 4870 -15
rect 4810 -85 4820 -45
rect 4860 -85 4870 -45
rect 4810 -110 4870 -85
rect 4810 -150 4820 -110
rect 4860 -150 4870 -110
rect 4810 -170 4870 -150
rect 4810 -210 4820 -170
rect 4860 -210 4870 -170
rect 4810 -235 4870 -210
rect 4810 -275 4820 -235
rect 4860 -275 4870 -235
rect 4810 -305 4870 -275
rect 4810 -345 4820 -305
rect 4860 -345 4870 -305
rect 4810 -375 4870 -345
rect 4810 -415 4820 -375
rect 4860 -415 4870 -375
rect 4810 -445 4870 -415
rect 4810 -485 4820 -445
rect 4860 -485 4870 -445
rect 4810 -510 4870 -485
rect 4810 -550 4820 -510
rect 4860 -550 4870 -510
rect 4810 -570 4870 -550
rect 4810 -610 4820 -570
rect 4860 -610 4870 -570
rect 4810 -635 4870 -610
rect 4810 -675 4820 -635
rect 4860 -675 4870 -635
rect 4810 -705 4870 -675
rect 4810 -745 4820 -705
rect 4860 -745 4870 -705
rect 4810 -775 4870 -745
rect 4810 -815 4820 -775
rect 4860 -815 4870 -775
rect 4810 -845 4870 -815
rect 4810 -885 4820 -845
rect 4860 -885 4870 -845
rect 4810 -910 4870 -885
rect 4810 -950 4820 -910
rect 4860 -950 4870 -910
rect 4810 -970 4870 -950
rect 4810 -1010 4820 -970
rect 4860 -1010 4870 -970
rect 4810 -1035 4870 -1010
rect 4810 -1075 4820 -1035
rect 4860 -1075 4870 -1035
rect 4810 -1105 4870 -1075
rect 4810 -1145 4820 -1105
rect 4860 -1145 4870 -1105
rect 4810 -1175 4870 -1145
rect 4810 -1215 4820 -1175
rect 4860 -1215 4870 -1175
rect 4810 -1245 4870 -1215
rect 4810 -1285 4820 -1245
rect 4860 -1285 4870 -1245
rect 4810 -1310 4870 -1285
rect 4810 -1350 4820 -1310
rect 4860 -1350 4870 -1310
rect 4810 -1360 4870 -1350
rect 5160 230 5220 240
rect 5160 190 5170 230
rect 5210 190 5220 230
rect 5160 165 5220 190
rect 5160 125 5170 165
rect 5210 125 5220 165
rect 5160 95 5220 125
rect 5160 55 5170 95
rect 5210 55 5220 95
rect 5160 25 5220 55
rect 5160 -15 5170 25
rect 5210 -15 5220 25
rect 5160 -45 5220 -15
rect 5160 -85 5170 -45
rect 5210 -85 5220 -45
rect 5160 -110 5220 -85
rect 5160 -150 5170 -110
rect 5210 -150 5220 -110
rect 5160 -170 5220 -150
rect 5160 -210 5170 -170
rect 5210 -210 5220 -170
rect 5160 -235 5220 -210
rect 5160 -275 5170 -235
rect 5210 -275 5220 -235
rect 5160 -305 5220 -275
rect 5160 -345 5170 -305
rect 5210 -345 5220 -305
rect 5160 -375 5220 -345
rect 5160 -415 5170 -375
rect 5210 -415 5220 -375
rect 5160 -445 5220 -415
rect 5160 -485 5170 -445
rect 5210 -485 5220 -445
rect 5160 -510 5220 -485
rect 5160 -550 5170 -510
rect 5210 -550 5220 -510
rect 5160 -570 5220 -550
rect 5160 -610 5170 -570
rect 5210 -610 5220 -570
rect 5160 -635 5220 -610
rect 5160 -675 5170 -635
rect 5210 -675 5220 -635
rect 5160 -705 5220 -675
rect 5160 -745 5170 -705
rect 5210 -745 5220 -705
rect 5160 -775 5220 -745
rect 5160 -815 5170 -775
rect 5210 -815 5220 -775
rect 5160 -845 5220 -815
rect 5160 -885 5170 -845
rect 5210 -885 5220 -845
rect 5160 -910 5220 -885
rect 5160 -950 5170 -910
rect 5210 -950 5220 -910
rect 5160 -970 5220 -950
rect 5160 -1010 5170 -970
rect 5210 -1010 5220 -970
rect 5160 -1035 5220 -1010
rect 5160 -1075 5170 -1035
rect 5210 -1075 5220 -1035
rect 5160 -1105 5220 -1075
rect 5160 -1145 5170 -1105
rect 5210 -1145 5220 -1105
rect 5160 -1175 5220 -1145
rect 5160 -1215 5170 -1175
rect 5210 -1215 5220 -1175
rect 5160 -1245 5220 -1215
rect 5160 -1285 5170 -1245
rect 5210 -1285 5220 -1245
rect 5160 -1310 5220 -1285
rect 5160 -1350 5170 -1310
rect 5210 -1350 5220 -1310
rect 5160 -1360 5220 -1350
rect 5510 230 5570 240
rect 5510 190 5520 230
rect 5560 190 5570 230
rect 5510 165 5570 190
rect 5510 125 5520 165
rect 5560 125 5570 165
rect 5510 95 5570 125
rect 5510 55 5520 95
rect 5560 55 5570 95
rect 5510 25 5570 55
rect 5510 -15 5520 25
rect 5560 -15 5570 25
rect 5510 -45 5570 -15
rect 5510 -85 5520 -45
rect 5560 -85 5570 -45
rect 5510 -110 5570 -85
rect 5510 -150 5520 -110
rect 5560 -150 5570 -110
rect 5510 -170 5570 -150
rect 5510 -210 5520 -170
rect 5560 -210 5570 -170
rect 5510 -235 5570 -210
rect 5510 -275 5520 -235
rect 5560 -275 5570 -235
rect 5510 -305 5570 -275
rect 5510 -345 5520 -305
rect 5560 -345 5570 -305
rect 5510 -375 5570 -345
rect 5510 -415 5520 -375
rect 5560 -415 5570 -375
rect 5510 -445 5570 -415
rect 5510 -485 5520 -445
rect 5560 -485 5570 -445
rect 5510 -510 5570 -485
rect 5510 -550 5520 -510
rect 5560 -550 5570 -510
rect 5510 -570 5570 -550
rect 5510 -610 5520 -570
rect 5560 -610 5570 -570
rect 5510 -635 5570 -610
rect 5510 -675 5520 -635
rect 5560 -675 5570 -635
rect 5510 -705 5570 -675
rect 5510 -745 5520 -705
rect 5560 -745 5570 -705
rect 5510 -775 5570 -745
rect 5510 -815 5520 -775
rect 5560 -815 5570 -775
rect 5510 -845 5570 -815
rect 5510 -885 5520 -845
rect 5560 -885 5570 -845
rect 5510 -910 5570 -885
rect 5510 -950 5520 -910
rect 5560 -950 5570 -910
rect 5510 -970 5570 -950
rect 5510 -1010 5520 -970
rect 5560 -1010 5570 -970
rect 5510 -1035 5570 -1010
rect 5510 -1075 5520 -1035
rect 5560 -1075 5570 -1035
rect 5510 -1105 5570 -1075
rect 5510 -1145 5520 -1105
rect 5560 -1145 5570 -1105
rect 5510 -1175 5570 -1145
rect 5510 -1215 5520 -1175
rect 5560 -1215 5570 -1175
rect 5510 -1245 5570 -1215
rect 5510 -1285 5520 -1245
rect 5560 -1285 5570 -1245
rect 5510 -1310 5570 -1285
rect 5510 -1350 5520 -1310
rect 5560 -1350 5570 -1310
rect 5510 -1360 5570 -1350
rect 5860 230 5920 240
rect 5860 190 5870 230
rect 5910 190 5920 230
rect 5860 165 5920 190
rect 5860 125 5870 165
rect 5910 125 5920 165
rect 5860 95 5920 125
rect 5860 55 5870 95
rect 5910 55 5920 95
rect 5860 25 5920 55
rect 5860 -15 5870 25
rect 5910 -15 5920 25
rect 5860 -45 5920 -15
rect 5860 -85 5870 -45
rect 5910 -85 5920 -45
rect 5860 -110 5920 -85
rect 5860 -150 5870 -110
rect 5910 -150 5920 -110
rect 5860 -170 5920 -150
rect 5860 -210 5870 -170
rect 5910 -210 5920 -170
rect 5860 -235 5920 -210
rect 5860 -275 5870 -235
rect 5910 -275 5920 -235
rect 5860 -305 5920 -275
rect 5860 -345 5870 -305
rect 5910 -345 5920 -305
rect 5860 -375 5920 -345
rect 5860 -415 5870 -375
rect 5910 -415 5920 -375
rect 5860 -445 5920 -415
rect 5860 -485 5870 -445
rect 5910 -485 5920 -445
rect 5860 -510 5920 -485
rect 5860 -550 5870 -510
rect 5910 -550 5920 -510
rect 5860 -570 5920 -550
rect 5860 -610 5870 -570
rect 5910 -610 5920 -570
rect 5860 -635 5920 -610
rect 5860 -675 5870 -635
rect 5910 -675 5920 -635
rect 5860 -705 5920 -675
rect 5860 -745 5870 -705
rect 5910 -745 5920 -705
rect 5860 -775 5920 -745
rect 5860 -815 5870 -775
rect 5910 -815 5920 -775
rect 5860 -845 5920 -815
rect 5860 -885 5870 -845
rect 5910 -885 5920 -845
rect 5860 -910 5920 -885
rect 5860 -950 5870 -910
rect 5910 -950 5920 -910
rect 5860 -970 5920 -950
rect 5860 -1010 5870 -970
rect 5910 -1010 5920 -970
rect 5860 -1035 5920 -1010
rect 5860 -1075 5870 -1035
rect 5910 -1075 5920 -1035
rect 5860 -1105 5920 -1075
rect 5860 -1145 5870 -1105
rect 5910 -1145 5920 -1105
rect 5860 -1175 5920 -1145
rect 5860 -1215 5870 -1175
rect 5910 -1215 5920 -1175
rect 5860 -1245 5920 -1215
rect 5860 -1285 5870 -1245
rect 5910 -1285 5920 -1245
rect 5860 -1310 5920 -1285
rect 5860 -1350 5870 -1310
rect 5910 -1350 5920 -1310
rect 5860 -1360 5920 -1350
rect 6210 230 6270 240
rect 6210 190 6220 230
rect 6260 190 6270 230
rect 6210 165 6270 190
rect 6210 125 6220 165
rect 6260 125 6270 165
rect 6210 95 6270 125
rect 6210 55 6220 95
rect 6260 55 6270 95
rect 6210 25 6270 55
rect 6210 -15 6220 25
rect 6260 -15 6270 25
rect 6210 -45 6270 -15
rect 6210 -85 6220 -45
rect 6260 -85 6270 -45
rect 6210 -110 6270 -85
rect 6210 -150 6220 -110
rect 6260 -150 6270 -110
rect 6210 -170 6270 -150
rect 6210 -210 6220 -170
rect 6260 -210 6270 -170
rect 6210 -235 6270 -210
rect 6210 -275 6220 -235
rect 6260 -275 6270 -235
rect 6210 -305 6270 -275
rect 6210 -345 6220 -305
rect 6260 -345 6270 -305
rect 6210 -375 6270 -345
rect 6210 -415 6220 -375
rect 6260 -415 6270 -375
rect 6210 -445 6270 -415
rect 6210 -485 6220 -445
rect 6260 -485 6270 -445
rect 6210 -510 6270 -485
rect 6210 -550 6220 -510
rect 6260 -550 6270 -510
rect 6210 -570 6270 -550
rect 6210 -610 6220 -570
rect 6260 -610 6270 -570
rect 6210 -635 6270 -610
rect 6210 -675 6220 -635
rect 6260 -675 6270 -635
rect 6210 -705 6270 -675
rect 6210 -745 6220 -705
rect 6260 -745 6270 -705
rect 6210 -775 6270 -745
rect 6210 -815 6220 -775
rect 6260 -815 6270 -775
rect 6210 -845 6270 -815
rect 6210 -885 6220 -845
rect 6260 -885 6270 -845
rect 6210 -910 6270 -885
rect 6210 -950 6220 -910
rect 6260 -950 6270 -910
rect 6210 -970 6270 -950
rect 6210 -1010 6220 -970
rect 6260 -1010 6270 -970
rect 6210 -1035 6270 -1010
rect 6210 -1075 6220 -1035
rect 6260 -1075 6270 -1035
rect 6210 -1105 6270 -1075
rect 6210 -1145 6220 -1105
rect 6260 -1145 6270 -1105
rect 6210 -1175 6270 -1145
rect 6210 -1215 6220 -1175
rect 6260 -1215 6270 -1175
rect 6210 -1245 6270 -1215
rect 6210 -1285 6220 -1245
rect 6260 -1285 6270 -1245
rect 6210 -1310 6270 -1285
rect 6210 -1350 6220 -1310
rect 6260 -1350 6270 -1310
rect 6210 -1360 6270 -1350
rect 6560 230 6620 240
rect 6560 190 6570 230
rect 6610 190 6620 230
rect 6560 165 6620 190
rect 6560 125 6570 165
rect 6610 125 6620 165
rect 6560 95 6620 125
rect 6560 55 6570 95
rect 6610 55 6620 95
rect 6560 25 6620 55
rect 6560 -15 6570 25
rect 6610 -15 6620 25
rect 6560 -45 6620 -15
rect 6560 -85 6570 -45
rect 6610 -85 6620 -45
rect 6560 -110 6620 -85
rect 6560 -150 6570 -110
rect 6610 -150 6620 -110
rect 6560 -170 6620 -150
rect 6560 -210 6570 -170
rect 6610 -210 6620 -170
rect 6560 -235 6620 -210
rect 6560 -275 6570 -235
rect 6610 -275 6620 -235
rect 6560 -305 6620 -275
rect 6560 -345 6570 -305
rect 6610 -345 6620 -305
rect 6560 -375 6620 -345
rect 6560 -415 6570 -375
rect 6610 -415 6620 -375
rect 6560 -445 6620 -415
rect 6560 -485 6570 -445
rect 6610 -485 6620 -445
rect 6560 -510 6620 -485
rect 6560 -550 6570 -510
rect 6610 -550 6620 -510
rect 6560 -570 6620 -550
rect 6560 -610 6570 -570
rect 6610 -610 6620 -570
rect 6560 -635 6620 -610
rect 6560 -675 6570 -635
rect 6610 -675 6620 -635
rect 6560 -705 6620 -675
rect 6560 -745 6570 -705
rect 6610 -745 6620 -705
rect 6560 -775 6620 -745
rect 6560 -815 6570 -775
rect 6610 -815 6620 -775
rect 6560 -845 6620 -815
rect 6560 -885 6570 -845
rect 6610 -885 6620 -845
rect 6560 -910 6620 -885
rect 6560 -950 6570 -910
rect 6610 -950 6620 -910
rect 6560 -970 6620 -950
rect 6560 -1010 6570 -970
rect 6610 -1010 6620 -970
rect 6560 -1035 6620 -1010
rect 6560 -1075 6570 -1035
rect 6610 -1075 6620 -1035
rect 6560 -1105 6620 -1075
rect 6560 -1145 6570 -1105
rect 6610 -1145 6620 -1105
rect 6560 -1175 6620 -1145
rect 6560 -1215 6570 -1175
rect 6610 -1215 6620 -1175
rect 6560 -1245 6620 -1215
rect 6560 -1285 6570 -1245
rect 6610 -1285 6620 -1245
rect 6560 -1310 6620 -1285
rect 6560 -1350 6570 -1310
rect 6610 -1350 6620 -1310
rect 6560 -1360 6620 -1350
rect 6910 230 6970 240
rect 6910 190 6920 230
rect 6960 190 6970 230
rect 6910 165 6970 190
rect 6910 125 6920 165
rect 6960 125 6970 165
rect 6910 95 6970 125
rect 6910 55 6920 95
rect 6960 55 6970 95
rect 6910 25 6970 55
rect 6910 -15 6920 25
rect 6960 -15 6970 25
rect 6910 -45 6970 -15
rect 6910 -85 6920 -45
rect 6960 -85 6970 -45
rect 6910 -110 6970 -85
rect 6910 -150 6920 -110
rect 6960 -150 6970 -110
rect 6910 -170 6970 -150
rect 6910 -210 6920 -170
rect 6960 -210 6970 -170
rect 6910 -235 6970 -210
rect 6910 -275 6920 -235
rect 6960 -275 6970 -235
rect 6910 -305 6970 -275
rect 6910 -345 6920 -305
rect 6960 -345 6970 -305
rect 6910 -375 6970 -345
rect 6910 -415 6920 -375
rect 6960 -415 6970 -375
rect 6910 -445 6970 -415
rect 6910 -485 6920 -445
rect 6960 -485 6970 -445
rect 6910 -510 6970 -485
rect 6910 -550 6920 -510
rect 6960 -550 6970 -510
rect 6910 -570 6970 -550
rect 6910 -610 6920 -570
rect 6960 -610 6970 -570
rect 6910 -635 6970 -610
rect 6910 -675 6920 -635
rect 6960 -675 6970 -635
rect 6910 -705 6970 -675
rect 6910 -745 6920 -705
rect 6960 -745 6970 -705
rect 6910 -775 6970 -745
rect 6910 -815 6920 -775
rect 6960 -815 6970 -775
rect 6910 -845 6970 -815
rect 6910 -885 6920 -845
rect 6960 -885 6970 -845
rect 6910 -910 6970 -885
rect 6910 -950 6920 -910
rect 6960 -950 6970 -910
rect 6910 -970 6970 -950
rect 6910 -1010 6920 -970
rect 6960 -1010 6970 -970
rect 6910 -1035 6970 -1010
rect 6910 -1075 6920 -1035
rect 6960 -1075 6970 -1035
rect 6910 -1105 6970 -1075
rect 6910 -1145 6920 -1105
rect 6960 -1145 6970 -1105
rect 6910 -1175 6970 -1145
rect 6910 -1215 6920 -1175
rect 6960 -1215 6970 -1175
rect 6910 -1245 6970 -1215
rect 6910 -1285 6920 -1245
rect 6960 -1285 6970 -1245
rect 6910 -1310 6970 -1285
rect 6910 -1350 6920 -1310
rect 6960 -1350 6970 -1310
rect 6910 -1360 6970 -1350
rect 7260 230 7320 240
rect 7260 190 7270 230
rect 7310 190 7320 230
rect 7260 165 7320 190
rect 7260 125 7270 165
rect 7310 125 7320 165
rect 7260 95 7320 125
rect 7260 55 7270 95
rect 7310 55 7320 95
rect 7260 25 7320 55
rect 7260 -15 7270 25
rect 7310 -15 7320 25
rect 7260 -45 7320 -15
rect 7260 -85 7270 -45
rect 7310 -85 7320 -45
rect 7260 -110 7320 -85
rect 7260 -150 7270 -110
rect 7310 -150 7320 -110
rect 7260 -170 7320 -150
rect 7260 -210 7270 -170
rect 7310 -210 7320 -170
rect 7260 -235 7320 -210
rect 7260 -275 7270 -235
rect 7310 -275 7320 -235
rect 7260 -305 7320 -275
rect 7260 -345 7270 -305
rect 7310 -345 7320 -305
rect 7260 -375 7320 -345
rect 7260 -415 7270 -375
rect 7310 -415 7320 -375
rect 7260 -445 7320 -415
rect 7260 -485 7270 -445
rect 7310 -485 7320 -445
rect 7260 -510 7320 -485
rect 7260 -550 7270 -510
rect 7310 -550 7320 -510
rect 7260 -570 7320 -550
rect 7260 -610 7270 -570
rect 7310 -610 7320 -570
rect 7260 -635 7320 -610
rect 7260 -675 7270 -635
rect 7310 -675 7320 -635
rect 7260 -705 7320 -675
rect 7260 -745 7270 -705
rect 7310 -745 7320 -705
rect 7260 -775 7320 -745
rect 7260 -815 7270 -775
rect 7310 -815 7320 -775
rect 7260 -845 7320 -815
rect 7260 -885 7270 -845
rect 7310 -885 7320 -845
rect 7260 -910 7320 -885
rect 7260 -950 7270 -910
rect 7310 -950 7320 -910
rect 7260 -970 7320 -950
rect 7260 -1010 7270 -970
rect 7310 -1010 7320 -970
rect 7260 -1035 7320 -1010
rect 7260 -1075 7270 -1035
rect 7310 -1075 7320 -1035
rect 7260 -1105 7320 -1075
rect 7260 -1145 7270 -1105
rect 7310 -1145 7320 -1105
rect 7260 -1175 7320 -1145
rect 7260 -1215 7270 -1175
rect 7310 -1215 7320 -1175
rect 7260 -1245 7320 -1215
rect 7260 -1285 7270 -1245
rect 7310 -1285 7320 -1245
rect 7260 -1310 7320 -1285
rect 7260 -1350 7270 -1310
rect 7310 -1350 7320 -1310
rect 7260 -1360 7320 -1350
rect 7610 230 7670 240
rect 7610 190 7620 230
rect 7660 190 7670 230
rect 7610 165 7670 190
rect 7610 125 7620 165
rect 7660 125 7670 165
rect 7610 95 7670 125
rect 7610 55 7620 95
rect 7660 55 7670 95
rect 7610 25 7670 55
rect 7610 -15 7620 25
rect 7660 -15 7670 25
rect 7610 -45 7670 -15
rect 7610 -85 7620 -45
rect 7660 -85 7670 -45
rect 7610 -110 7670 -85
rect 7610 -150 7620 -110
rect 7660 -150 7670 -110
rect 7610 -170 7670 -150
rect 7610 -210 7620 -170
rect 7660 -210 7670 -170
rect 7610 -235 7670 -210
rect 7610 -275 7620 -235
rect 7660 -275 7670 -235
rect 7610 -305 7670 -275
rect 7610 -345 7620 -305
rect 7660 -345 7670 -305
rect 7610 -375 7670 -345
rect 7610 -415 7620 -375
rect 7660 -415 7670 -375
rect 7610 -445 7670 -415
rect 7610 -485 7620 -445
rect 7660 -485 7670 -445
rect 7610 -510 7670 -485
rect 7610 -550 7620 -510
rect 7660 -550 7670 -510
rect 7610 -570 7670 -550
rect 7610 -610 7620 -570
rect 7660 -610 7670 -570
rect 7610 -635 7670 -610
rect 7610 -675 7620 -635
rect 7660 -675 7670 -635
rect 7610 -705 7670 -675
rect 7610 -745 7620 -705
rect 7660 -745 7670 -705
rect 7610 -775 7670 -745
rect 7610 -815 7620 -775
rect 7660 -815 7670 -775
rect 7610 -845 7670 -815
rect 7610 -885 7620 -845
rect 7660 -885 7670 -845
rect 7610 -910 7670 -885
rect 7610 -950 7620 -910
rect 7660 -950 7670 -910
rect 7610 -970 7670 -950
rect 7610 -1010 7620 -970
rect 7660 -1010 7670 -970
rect 7610 -1035 7670 -1010
rect 7610 -1075 7620 -1035
rect 7660 -1075 7670 -1035
rect 7610 -1105 7670 -1075
rect 7610 -1145 7620 -1105
rect 7660 -1145 7670 -1105
rect 7610 -1175 7670 -1145
rect 7610 -1215 7620 -1175
rect 7660 -1215 7670 -1175
rect 7610 -1245 7670 -1215
rect 7610 -1285 7620 -1245
rect 7660 -1285 7670 -1245
rect 7610 -1310 7670 -1285
rect 7610 -1350 7620 -1310
rect 7660 -1350 7670 -1310
rect 7610 -1360 7670 -1350
rect 7960 230 8020 240
rect 7960 190 7970 230
rect 8010 190 8020 230
rect 7960 165 8020 190
rect 7960 125 7970 165
rect 8010 125 8020 165
rect 7960 95 8020 125
rect 7960 55 7970 95
rect 8010 55 8020 95
rect 7960 25 8020 55
rect 7960 -15 7970 25
rect 8010 -15 8020 25
rect 7960 -45 8020 -15
rect 7960 -85 7970 -45
rect 8010 -85 8020 -45
rect 7960 -110 8020 -85
rect 7960 -150 7970 -110
rect 8010 -150 8020 -110
rect 7960 -170 8020 -150
rect 7960 -210 7970 -170
rect 8010 -210 8020 -170
rect 7960 -235 8020 -210
rect 7960 -275 7970 -235
rect 8010 -275 8020 -235
rect 7960 -305 8020 -275
rect 7960 -345 7970 -305
rect 8010 -345 8020 -305
rect 7960 -375 8020 -345
rect 7960 -415 7970 -375
rect 8010 -415 8020 -375
rect 7960 -445 8020 -415
rect 7960 -485 7970 -445
rect 8010 -485 8020 -445
rect 7960 -510 8020 -485
rect 7960 -550 7970 -510
rect 8010 -550 8020 -510
rect 7960 -570 8020 -550
rect 7960 -610 7970 -570
rect 8010 -610 8020 -570
rect 7960 -635 8020 -610
rect 7960 -675 7970 -635
rect 8010 -675 8020 -635
rect 7960 -705 8020 -675
rect 7960 -745 7970 -705
rect 8010 -745 8020 -705
rect 7960 -775 8020 -745
rect 7960 -815 7970 -775
rect 8010 -815 8020 -775
rect 7960 -845 8020 -815
rect 7960 -885 7970 -845
rect 8010 -885 8020 -845
rect 7960 -910 8020 -885
rect 7960 -950 7970 -910
rect 8010 -950 8020 -910
rect 7960 -970 8020 -950
rect 7960 -1010 7970 -970
rect 8010 -1010 8020 -970
rect 7960 -1035 8020 -1010
rect 7960 -1075 7970 -1035
rect 8010 -1075 8020 -1035
rect 7960 -1105 8020 -1075
rect 7960 -1145 7970 -1105
rect 8010 -1145 8020 -1105
rect 7960 -1175 8020 -1145
rect 7960 -1215 7970 -1175
rect 8010 -1215 8020 -1175
rect 7960 -1245 8020 -1215
rect 7960 -1285 7970 -1245
rect 8010 -1285 8020 -1245
rect 7960 -1310 8020 -1285
rect 7960 -1350 7970 -1310
rect 8010 -1350 8020 -1310
rect 7960 -1360 8020 -1350
rect 8310 230 8370 240
rect 8310 190 8320 230
rect 8360 190 8370 230
rect 8310 165 8370 190
rect 8310 125 8320 165
rect 8360 125 8370 165
rect 8310 95 8370 125
rect 8310 55 8320 95
rect 8360 55 8370 95
rect 8310 25 8370 55
rect 8310 -15 8320 25
rect 8360 -15 8370 25
rect 8310 -45 8370 -15
rect 8310 -85 8320 -45
rect 8360 -85 8370 -45
rect 8310 -110 8370 -85
rect 8310 -150 8320 -110
rect 8360 -150 8370 -110
rect 8310 -170 8370 -150
rect 8310 -210 8320 -170
rect 8360 -210 8370 -170
rect 8310 -235 8370 -210
rect 8310 -275 8320 -235
rect 8360 -275 8370 -235
rect 8310 -305 8370 -275
rect 8310 -345 8320 -305
rect 8360 -345 8370 -305
rect 8310 -375 8370 -345
rect 8310 -415 8320 -375
rect 8360 -415 8370 -375
rect 8310 -445 8370 -415
rect 8310 -485 8320 -445
rect 8360 -485 8370 -445
rect 8310 -510 8370 -485
rect 8310 -550 8320 -510
rect 8360 -550 8370 -510
rect 8310 -570 8370 -550
rect 8310 -610 8320 -570
rect 8360 -610 8370 -570
rect 8310 -635 8370 -610
rect 8310 -675 8320 -635
rect 8360 -675 8370 -635
rect 8310 -705 8370 -675
rect 8310 -745 8320 -705
rect 8360 -745 8370 -705
rect 8310 -775 8370 -745
rect 8310 -815 8320 -775
rect 8360 -815 8370 -775
rect 8310 -845 8370 -815
rect 8310 -885 8320 -845
rect 8360 -885 8370 -845
rect 8310 -910 8370 -885
rect 8310 -950 8320 -910
rect 8360 -950 8370 -910
rect 8310 -970 8370 -950
rect 8310 -1010 8320 -970
rect 8360 -1010 8370 -970
rect 8310 -1035 8370 -1010
rect 8310 -1075 8320 -1035
rect 8360 -1075 8370 -1035
rect 8310 -1105 8370 -1075
rect 8310 -1145 8320 -1105
rect 8360 -1145 8370 -1105
rect 8310 -1175 8370 -1145
rect 8310 -1215 8320 -1175
rect 8360 -1215 8370 -1175
rect 8310 -1245 8370 -1215
rect 8310 -1285 8320 -1245
rect 8360 -1285 8370 -1245
rect 8310 -1310 8370 -1285
rect 8310 -1350 8320 -1310
rect 8360 -1350 8370 -1310
rect 8310 -1360 8370 -1350
rect 8660 230 8720 240
rect 8660 190 8670 230
rect 8710 190 8720 230
rect 8660 165 8720 190
rect 8660 125 8670 165
rect 8710 125 8720 165
rect 8660 95 8720 125
rect 8660 55 8670 95
rect 8710 55 8720 95
rect 8660 25 8720 55
rect 8660 -15 8670 25
rect 8710 -15 8720 25
rect 8660 -45 8720 -15
rect 8660 -85 8670 -45
rect 8710 -85 8720 -45
rect 8660 -110 8720 -85
rect 8660 -150 8670 -110
rect 8710 -150 8720 -110
rect 8660 -170 8720 -150
rect 8660 -210 8670 -170
rect 8710 -210 8720 -170
rect 8660 -235 8720 -210
rect 8660 -275 8670 -235
rect 8710 -275 8720 -235
rect 8660 -305 8720 -275
rect 8660 -345 8670 -305
rect 8710 -345 8720 -305
rect 8660 -375 8720 -345
rect 8660 -415 8670 -375
rect 8710 -415 8720 -375
rect 8660 -445 8720 -415
rect 8660 -485 8670 -445
rect 8710 -485 8720 -445
rect 8660 -510 8720 -485
rect 8660 -550 8670 -510
rect 8710 -550 8720 -510
rect 8660 -570 8720 -550
rect 8660 -610 8670 -570
rect 8710 -610 8720 -570
rect 8660 -635 8720 -610
rect 8660 -675 8670 -635
rect 8710 -675 8720 -635
rect 8660 -705 8720 -675
rect 8660 -745 8670 -705
rect 8710 -745 8720 -705
rect 8660 -775 8720 -745
rect 8660 -815 8670 -775
rect 8710 -815 8720 -775
rect 8660 -845 8720 -815
rect 8660 -885 8670 -845
rect 8710 -885 8720 -845
rect 8660 -910 8720 -885
rect 8660 -950 8670 -910
rect 8710 -950 8720 -910
rect 8660 -970 8720 -950
rect 8660 -1010 8670 -970
rect 8710 -1010 8720 -970
rect 8660 -1035 8720 -1010
rect 8660 -1075 8670 -1035
rect 8710 -1075 8720 -1035
rect 8660 -1105 8720 -1075
rect 8660 -1145 8670 -1105
rect 8710 -1145 8720 -1105
rect 8660 -1175 8720 -1145
rect 8660 -1215 8670 -1175
rect 8710 -1215 8720 -1175
rect 8660 -1245 8720 -1215
rect 8660 -1285 8670 -1245
rect 8710 -1285 8720 -1245
rect 8660 -1310 8720 -1285
rect 8660 -1350 8670 -1310
rect 8710 -1350 8720 -1310
rect 8660 -1360 8720 -1350
rect 9010 230 9070 240
rect 9010 190 9020 230
rect 9060 190 9070 230
rect 9010 165 9070 190
rect 9010 125 9020 165
rect 9060 125 9070 165
rect 9010 95 9070 125
rect 9010 55 9020 95
rect 9060 55 9070 95
rect 9010 25 9070 55
rect 9010 -15 9020 25
rect 9060 -15 9070 25
rect 9010 -45 9070 -15
rect 9010 -85 9020 -45
rect 9060 -85 9070 -45
rect 9010 -110 9070 -85
rect 9010 -150 9020 -110
rect 9060 -150 9070 -110
rect 9010 -170 9070 -150
rect 9010 -210 9020 -170
rect 9060 -210 9070 -170
rect 9010 -235 9070 -210
rect 9010 -275 9020 -235
rect 9060 -275 9070 -235
rect 9010 -305 9070 -275
rect 9010 -345 9020 -305
rect 9060 -345 9070 -305
rect 9010 -375 9070 -345
rect 9010 -415 9020 -375
rect 9060 -415 9070 -375
rect 9010 -445 9070 -415
rect 9010 -485 9020 -445
rect 9060 -485 9070 -445
rect 9010 -510 9070 -485
rect 9010 -550 9020 -510
rect 9060 -550 9070 -510
rect 9010 -570 9070 -550
rect 9010 -610 9020 -570
rect 9060 -610 9070 -570
rect 9010 -635 9070 -610
rect 9010 -675 9020 -635
rect 9060 -675 9070 -635
rect 9010 -705 9070 -675
rect 9010 -745 9020 -705
rect 9060 -745 9070 -705
rect 9010 -775 9070 -745
rect 9010 -815 9020 -775
rect 9060 -815 9070 -775
rect 9010 -845 9070 -815
rect 9010 -885 9020 -845
rect 9060 -885 9070 -845
rect 9010 -910 9070 -885
rect 9010 -950 9020 -910
rect 9060 -950 9070 -910
rect 9010 -970 9070 -950
rect 9010 -1010 9020 -970
rect 9060 -1010 9070 -970
rect 9010 -1035 9070 -1010
rect 9010 -1075 9020 -1035
rect 9060 -1075 9070 -1035
rect 9010 -1105 9070 -1075
rect 9010 -1145 9020 -1105
rect 9060 -1145 9070 -1105
rect 9010 -1175 9070 -1145
rect 9010 -1215 9020 -1175
rect 9060 -1215 9070 -1175
rect 9010 -1245 9070 -1215
rect 9010 -1285 9020 -1245
rect 9060 -1285 9070 -1245
rect 9010 -1310 9070 -1285
rect 9010 -1350 9020 -1310
rect 9060 -1350 9070 -1310
rect 9010 -1360 9070 -1350
rect 31290 220 32890 8965
rect 31290 185 31305 220
rect 31340 185 31350 220
rect 31385 185 31395 220
rect 31430 185 31440 220
rect 31475 185 31485 220
rect 31520 185 31530 220
rect 31565 185 31575 220
rect 31610 185 31620 220
rect 31655 185 31665 220
rect 31700 185 31710 220
rect 31745 185 31755 220
rect 31790 185 31800 220
rect 31835 185 31845 220
rect 31880 185 31890 220
rect 31925 185 31935 220
rect 31970 185 31980 220
rect 32015 185 32025 220
rect 32060 185 32070 220
rect 32105 185 32115 220
rect 32150 185 32160 220
rect 32195 185 32205 220
rect 32240 185 32250 220
rect 32285 185 32295 220
rect 32330 185 32340 220
rect 32375 185 32385 220
rect 32420 185 32430 220
rect 32465 185 32475 220
rect 32510 185 32520 220
rect 32555 185 32565 220
rect 32600 185 32610 220
rect 32645 185 32655 220
rect 32690 185 32700 220
rect 32735 185 32745 220
rect 32780 185 32790 220
rect 32825 185 32835 220
rect 32870 185 32890 220
rect 31290 175 32890 185
rect 31290 140 31305 175
rect 31340 140 31350 175
rect 31385 140 31395 175
rect 31430 140 31440 175
rect 31475 140 31485 175
rect 31520 140 31530 175
rect 31565 140 31575 175
rect 31610 140 31620 175
rect 31655 140 31665 175
rect 31700 140 31710 175
rect 31745 140 31755 175
rect 31790 140 31800 175
rect 31835 140 31845 175
rect 31880 140 31890 175
rect 31925 140 31935 175
rect 31970 140 31980 175
rect 32015 140 32025 175
rect 32060 140 32070 175
rect 32105 140 32115 175
rect 32150 140 32160 175
rect 32195 140 32205 175
rect 32240 140 32250 175
rect 32285 140 32295 175
rect 32330 140 32340 175
rect 32375 140 32385 175
rect 32420 140 32430 175
rect 32465 140 32475 175
rect 32510 140 32520 175
rect 32555 140 32565 175
rect 32600 140 32610 175
rect 32645 140 32655 175
rect 32690 140 32700 175
rect 32735 140 32745 175
rect 32780 140 32790 175
rect 32825 140 32835 175
rect 32870 140 32890 175
rect 31290 130 32890 140
rect 31290 95 31305 130
rect 31340 95 31350 130
rect 31385 95 31395 130
rect 31430 95 31440 130
rect 31475 95 31485 130
rect 31520 95 31530 130
rect 31565 95 31575 130
rect 31610 95 31620 130
rect 31655 95 31665 130
rect 31700 95 31710 130
rect 31745 95 31755 130
rect 31790 95 31800 130
rect 31835 95 31845 130
rect 31880 95 31890 130
rect 31925 95 31935 130
rect 31970 95 31980 130
rect 32015 95 32025 130
rect 32060 95 32070 130
rect 32105 95 32115 130
rect 32150 95 32160 130
rect 32195 95 32205 130
rect 32240 95 32250 130
rect 32285 95 32295 130
rect 32330 95 32340 130
rect 32375 95 32385 130
rect 32420 95 32430 130
rect 32465 95 32475 130
rect 32510 95 32520 130
rect 32555 95 32565 130
rect 32600 95 32610 130
rect 32645 95 32655 130
rect 32690 95 32700 130
rect 32735 95 32745 130
rect 32780 95 32790 130
rect 32825 95 32835 130
rect 32870 95 32890 130
rect 31290 85 32890 95
rect 31290 50 31305 85
rect 31340 50 31350 85
rect 31385 50 31395 85
rect 31430 50 31440 85
rect 31475 50 31485 85
rect 31520 50 31530 85
rect 31565 50 31575 85
rect 31610 50 31620 85
rect 31655 50 31665 85
rect 31700 50 31710 85
rect 31745 50 31755 85
rect 31790 50 31800 85
rect 31835 50 31845 85
rect 31880 50 31890 85
rect 31925 50 31935 85
rect 31970 50 31980 85
rect 32015 50 32025 85
rect 32060 50 32070 85
rect 32105 50 32115 85
rect 32150 50 32160 85
rect 32195 50 32205 85
rect 32240 50 32250 85
rect 32285 50 32295 85
rect 32330 50 32340 85
rect 32375 50 32385 85
rect 32420 50 32430 85
rect 32465 50 32475 85
rect 32510 50 32520 85
rect 32555 50 32565 85
rect 32600 50 32610 85
rect 32645 50 32655 85
rect 32690 50 32700 85
rect 32735 50 32745 85
rect 32780 50 32790 85
rect 32825 50 32835 85
rect 32870 50 32890 85
rect 31290 40 32890 50
rect 31290 5 31305 40
rect 31340 5 31350 40
rect 31385 5 31395 40
rect 31430 5 31440 40
rect 31475 5 31485 40
rect 31520 5 31530 40
rect 31565 5 31575 40
rect 31610 5 31620 40
rect 31655 5 31665 40
rect 31700 5 31710 40
rect 31745 5 31755 40
rect 31790 5 31800 40
rect 31835 5 31845 40
rect 31880 5 31890 40
rect 31925 5 31935 40
rect 31970 5 31980 40
rect 32015 5 32025 40
rect 32060 5 32070 40
rect 32105 5 32115 40
rect 32150 5 32160 40
rect 32195 5 32205 40
rect 32240 5 32250 40
rect 32285 5 32295 40
rect 32330 5 32340 40
rect 32375 5 32385 40
rect 32420 5 32430 40
rect 32465 5 32475 40
rect 32510 5 32520 40
rect 32555 5 32565 40
rect 32600 5 32610 40
rect 32645 5 32655 40
rect 32690 5 32700 40
rect 32735 5 32745 40
rect 32780 5 32790 40
rect 32825 5 32835 40
rect 32870 5 32890 40
rect 31290 -5 32890 5
rect 31290 -40 31305 -5
rect 31340 -40 31350 -5
rect 31385 -40 31395 -5
rect 31430 -40 31440 -5
rect 31475 -40 31485 -5
rect 31520 -40 31530 -5
rect 31565 -40 31575 -5
rect 31610 -40 31620 -5
rect 31655 -40 31665 -5
rect 31700 -40 31710 -5
rect 31745 -40 31755 -5
rect 31790 -40 31800 -5
rect 31835 -40 31845 -5
rect 31880 -40 31890 -5
rect 31925 -40 31935 -5
rect 31970 -40 31980 -5
rect 32015 -40 32025 -5
rect 32060 -40 32070 -5
rect 32105 -40 32115 -5
rect 32150 -40 32160 -5
rect 32195 -40 32205 -5
rect 32240 -40 32250 -5
rect 32285 -40 32295 -5
rect 32330 -40 32340 -5
rect 32375 -40 32385 -5
rect 32420 -40 32430 -5
rect 32465 -40 32475 -5
rect 32510 -40 32520 -5
rect 32555 -40 32565 -5
rect 32600 -40 32610 -5
rect 32645 -40 32655 -5
rect 32690 -40 32700 -5
rect 32735 -40 32745 -5
rect 32780 -40 32790 -5
rect 32825 -40 32835 -5
rect 32870 -40 32890 -5
rect 31290 -50 32890 -40
rect 31290 -85 31305 -50
rect 31340 -85 31350 -50
rect 31385 -85 31395 -50
rect 31430 -85 31440 -50
rect 31475 -85 31485 -50
rect 31520 -85 31530 -50
rect 31565 -85 31575 -50
rect 31610 -85 31620 -50
rect 31655 -85 31665 -50
rect 31700 -85 31710 -50
rect 31745 -85 31755 -50
rect 31790 -85 31800 -50
rect 31835 -85 31845 -50
rect 31880 -85 31890 -50
rect 31925 -85 31935 -50
rect 31970 -85 31980 -50
rect 32015 -85 32025 -50
rect 32060 -85 32070 -50
rect 32105 -85 32115 -50
rect 32150 -85 32160 -50
rect 32195 -85 32205 -50
rect 32240 -85 32250 -50
rect 32285 -85 32295 -50
rect 32330 -85 32340 -50
rect 32375 -85 32385 -50
rect 32420 -85 32430 -50
rect 32465 -85 32475 -50
rect 32510 -85 32520 -50
rect 32555 -85 32565 -50
rect 32600 -85 32610 -50
rect 32645 -85 32655 -50
rect 32690 -85 32700 -50
rect 32735 -85 32745 -50
rect 32780 -85 32790 -50
rect 32825 -85 32835 -50
rect 32870 -85 32890 -50
rect 31290 -95 32890 -85
rect 31290 -130 31305 -95
rect 31340 -130 31350 -95
rect 31385 -130 31395 -95
rect 31430 -130 31440 -95
rect 31475 -130 31485 -95
rect 31520 -130 31530 -95
rect 31565 -130 31575 -95
rect 31610 -130 31620 -95
rect 31655 -130 31665 -95
rect 31700 -130 31710 -95
rect 31745 -130 31755 -95
rect 31790 -130 31800 -95
rect 31835 -130 31845 -95
rect 31880 -130 31890 -95
rect 31925 -130 31935 -95
rect 31970 -130 31980 -95
rect 32015 -130 32025 -95
rect 32060 -130 32070 -95
rect 32105 -130 32115 -95
rect 32150 -130 32160 -95
rect 32195 -130 32205 -95
rect 32240 -130 32250 -95
rect 32285 -130 32295 -95
rect 32330 -130 32340 -95
rect 32375 -130 32385 -95
rect 32420 -130 32430 -95
rect 32465 -130 32475 -95
rect 32510 -130 32520 -95
rect 32555 -130 32565 -95
rect 32600 -130 32610 -95
rect 32645 -130 32655 -95
rect 32690 -130 32700 -95
rect 32735 -130 32745 -95
rect 32780 -130 32790 -95
rect 32825 -130 32835 -95
rect 32870 -130 32890 -95
rect 31290 -140 32890 -130
rect 31290 -175 31305 -140
rect 31340 -175 31350 -140
rect 31385 -175 31395 -140
rect 31430 -175 31440 -140
rect 31475 -175 31485 -140
rect 31520 -175 31530 -140
rect 31565 -175 31575 -140
rect 31610 -175 31620 -140
rect 31655 -175 31665 -140
rect 31700 -175 31710 -140
rect 31745 -175 31755 -140
rect 31790 -175 31800 -140
rect 31835 -175 31845 -140
rect 31880 -175 31890 -140
rect 31925 -175 31935 -140
rect 31970 -175 31980 -140
rect 32015 -175 32025 -140
rect 32060 -175 32070 -140
rect 32105 -175 32115 -140
rect 32150 -175 32160 -140
rect 32195 -175 32205 -140
rect 32240 -175 32250 -140
rect 32285 -175 32295 -140
rect 32330 -175 32340 -140
rect 32375 -175 32385 -140
rect 32420 -175 32430 -140
rect 32465 -175 32475 -140
rect 32510 -175 32520 -140
rect 32555 -175 32565 -140
rect 32600 -175 32610 -140
rect 32645 -175 32655 -140
rect 32690 -175 32700 -140
rect 32735 -175 32745 -140
rect 32780 -175 32790 -140
rect 32825 -175 32835 -140
rect 32870 -175 32890 -140
rect 31290 -185 32890 -175
rect 31290 -220 31305 -185
rect 31340 -220 31350 -185
rect 31385 -220 31395 -185
rect 31430 -220 31440 -185
rect 31475 -220 31485 -185
rect 31520 -220 31530 -185
rect 31565 -220 31575 -185
rect 31610 -220 31620 -185
rect 31655 -220 31665 -185
rect 31700 -220 31710 -185
rect 31745 -220 31755 -185
rect 31790 -220 31800 -185
rect 31835 -220 31845 -185
rect 31880 -220 31890 -185
rect 31925 -220 31935 -185
rect 31970 -220 31980 -185
rect 32015 -220 32025 -185
rect 32060 -220 32070 -185
rect 32105 -220 32115 -185
rect 32150 -220 32160 -185
rect 32195 -220 32205 -185
rect 32240 -220 32250 -185
rect 32285 -220 32295 -185
rect 32330 -220 32340 -185
rect 32375 -220 32385 -185
rect 32420 -220 32430 -185
rect 32465 -220 32475 -185
rect 32510 -220 32520 -185
rect 32555 -220 32565 -185
rect 32600 -220 32610 -185
rect 32645 -220 32655 -185
rect 32690 -220 32700 -185
rect 32735 -220 32745 -185
rect 32780 -220 32790 -185
rect 32825 -220 32835 -185
rect 32870 -220 32890 -185
rect 31290 -230 32890 -220
rect 31290 -265 31305 -230
rect 31340 -265 31350 -230
rect 31385 -265 31395 -230
rect 31430 -265 31440 -230
rect 31475 -265 31485 -230
rect 31520 -265 31530 -230
rect 31565 -265 31575 -230
rect 31610 -265 31620 -230
rect 31655 -265 31665 -230
rect 31700 -265 31710 -230
rect 31745 -265 31755 -230
rect 31790 -265 31800 -230
rect 31835 -265 31845 -230
rect 31880 -265 31890 -230
rect 31925 -265 31935 -230
rect 31970 -265 31980 -230
rect 32015 -265 32025 -230
rect 32060 -265 32070 -230
rect 32105 -265 32115 -230
rect 32150 -265 32160 -230
rect 32195 -265 32205 -230
rect 32240 -265 32250 -230
rect 32285 -265 32295 -230
rect 32330 -265 32340 -230
rect 32375 -265 32385 -230
rect 32420 -265 32430 -230
rect 32465 -265 32475 -230
rect 32510 -265 32520 -230
rect 32555 -265 32565 -230
rect 32600 -265 32610 -230
rect 32645 -265 32655 -230
rect 32690 -265 32700 -230
rect 32735 -265 32745 -230
rect 32780 -265 32790 -230
rect 32825 -265 32835 -230
rect 32870 -265 32890 -230
rect 31290 -275 32890 -265
rect 31290 -310 31305 -275
rect 31340 -310 31350 -275
rect 31385 -310 31395 -275
rect 31430 -310 31440 -275
rect 31475 -310 31485 -275
rect 31520 -310 31530 -275
rect 31565 -310 31575 -275
rect 31610 -310 31620 -275
rect 31655 -310 31665 -275
rect 31700 -310 31710 -275
rect 31745 -310 31755 -275
rect 31790 -310 31800 -275
rect 31835 -310 31845 -275
rect 31880 -310 31890 -275
rect 31925 -310 31935 -275
rect 31970 -310 31980 -275
rect 32015 -310 32025 -275
rect 32060 -310 32070 -275
rect 32105 -310 32115 -275
rect 32150 -310 32160 -275
rect 32195 -310 32205 -275
rect 32240 -310 32250 -275
rect 32285 -310 32295 -275
rect 32330 -310 32340 -275
rect 32375 -310 32385 -275
rect 32420 -310 32430 -275
rect 32465 -310 32475 -275
rect 32510 -310 32520 -275
rect 32555 -310 32565 -275
rect 32600 -310 32610 -275
rect 32645 -310 32655 -275
rect 32690 -310 32700 -275
rect 32735 -310 32745 -275
rect 32780 -310 32790 -275
rect 32825 -310 32835 -275
rect 32870 -310 32890 -275
rect 31290 -320 32890 -310
rect 31290 -355 31305 -320
rect 31340 -355 31350 -320
rect 31385 -355 31395 -320
rect 31430 -355 31440 -320
rect 31475 -355 31485 -320
rect 31520 -355 31530 -320
rect 31565 -355 31575 -320
rect 31610 -355 31620 -320
rect 31655 -355 31665 -320
rect 31700 -355 31710 -320
rect 31745 -355 31755 -320
rect 31790 -355 31800 -320
rect 31835 -355 31845 -320
rect 31880 -355 31890 -320
rect 31925 -355 31935 -320
rect 31970 -355 31980 -320
rect 32015 -355 32025 -320
rect 32060 -355 32070 -320
rect 32105 -355 32115 -320
rect 32150 -355 32160 -320
rect 32195 -355 32205 -320
rect 32240 -355 32250 -320
rect 32285 -355 32295 -320
rect 32330 -355 32340 -320
rect 32375 -355 32385 -320
rect 32420 -355 32430 -320
rect 32465 -355 32475 -320
rect 32510 -355 32520 -320
rect 32555 -355 32565 -320
rect 32600 -355 32610 -320
rect 32645 -355 32655 -320
rect 32690 -355 32700 -320
rect 32735 -355 32745 -320
rect 32780 -355 32790 -320
rect 32825 -355 32835 -320
rect 32870 -355 32890 -320
rect 31290 -365 32890 -355
rect 31290 -400 31305 -365
rect 31340 -400 31350 -365
rect 31385 -400 31395 -365
rect 31430 -400 31440 -365
rect 31475 -400 31485 -365
rect 31520 -400 31530 -365
rect 31565 -400 31575 -365
rect 31610 -400 31620 -365
rect 31655 -400 31665 -365
rect 31700 -400 31710 -365
rect 31745 -400 31755 -365
rect 31790 -400 31800 -365
rect 31835 -400 31845 -365
rect 31880 -400 31890 -365
rect 31925 -400 31935 -365
rect 31970 -400 31980 -365
rect 32015 -400 32025 -365
rect 32060 -400 32070 -365
rect 32105 -400 32115 -365
rect 32150 -400 32160 -365
rect 32195 -400 32205 -365
rect 32240 -400 32250 -365
rect 32285 -400 32295 -365
rect 32330 -400 32340 -365
rect 32375 -400 32385 -365
rect 32420 -400 32430 -365
rect 32465 -400 32475 -365
rect 32510 -400 32520 -365
rect 32555 -400 32565 -365
rect 32600 -400 32610 -365
rect 32645 -400 32655 -365
rect 32690 -400 32700 -365
rect 32735 -400 32745 -365
rect 32780 -400 32790 -365
rect 32825 -400 32835 -365
rect 32870 -400 32890 -365
rect 31290 -410 32890 -400
rect 31290 -445 31305 -410
rect 31340 -445 31350 -410
rect 31385 -445 31395 -410
rect 31430 -445 31440 -410
rect 31475 -445 31485 -410
rect 31520 -445 31530 -410
rect 31565 -445 31575 -410
rect 31610 -445 31620 -410
rect 31655 -445 31665 -410
rect 31700 -445 31710 -410
rect 31745 -445 31755 -410
rect 31790 -445 31800 -410
rect 31835 -445 31845 -410
rect 31880 -445 31890 -410
rect 31925 -445 31935 -410
rect 31970 -445 31980 -410
rect 32015 -445 32025 -410
rect 32060 -445 32070 -410
rect 32105 -445 32115 -410
rect 32150 -445 32160 -410
rect 32195 -445 32205 -410
rect 32240 -445 32250 -410
rect 32285 -445 32295 -410
rect 32330 -445 32340 -410
rect 32375 -445 32385 -410
rect 32420 -445 32430 -410
rect 32465 -445 32475 -410
rect 32510 -445 32520 -410
rect 32555 -445 32565 -410
rect 32600 -445 32610 -410
rect 32645 -445 32655 -410
rect 32690 -445 32700 -410
rect 32735 -445 32745 -410
rect 32780 -445 32790 -410
rect 32825 -445 32835 -410
rect 32870 -445 32890 -410
rect 31290 -455 32890 -445
rect 31290 -490 31305 -455
rect 31340 -490 31350 -455
rect 31385 -490 31395 -455
rect 31430 -490 31440 -455
rect 31475 -490 31485 -455
rect 31520 -490 31530 -455
rect 31565 -490 31575 -455
rect 31610 -490 31620 -455
rect 31655 -490 31665 -455
rect 31700 -490 31710 -455
rect 31745 -490 31755 -455
rect 31790 -490 31800 -455
rect 31835 -490 31845 -455
rect 31880 -490 31890 -455
rect 31925 -490 31935 -455
rect 31970 -490 31980 -455
rect 32015 -490 32025 -455
rect 32060 -490 32070 -455
rect 32105 -490 32115 -455
rect 32150 -490 32160 -455
rect 32195 -490 32205 -455
rect 32240 -490 32250 -455
rect 32285 -490 32295 -455
rect 32330 -490 32340 -455
rect 32375 -490 32385 -455
rect 32420 -490 32430 -455
rect 32465 -490 32475 -455
rect 32510 -490 32520 -455
rect 32555 -490 32565 -455
rect 32600 -490 32610 -455
rect 32645 -490 32655 -455
rect 32690 -490 32700 -455
rect 32735 -490 32745 -455
rect 32780 -490 32790 -455
rect 32825 -490 32835 -455
rect 32870 -490 32890 -455
rect 31290 -500 32890 -490
rect 31290 -535 31305 -500
rect 31340 -535 31350 -500
rect 31385 -535 31395 -500
rect 31430 -535 31440 -500
rect 31475 -535 31485 -500
rect 31520 -535 31530 -500
rect 31565 -535 31575 -500
rect 31610 -535 31620 -500
rect 31655 -535 31665 -500
rect 31700 -535 31710 -500
rect 31745 -535 31755 -500
rect 31790 -535 31800 -500
rect 31835 -535 31845 -500
rect 31880 -535 31890 -500
rect 31925 -535 31935 -500
rect 31970 -535 31980 -500
rect 32015 -535 32025 -500
rect 32060 -535 32070 -500
rect 32105 -535 32115 -500
rect 32150 -535 32160 -500
rect 32195 -535 32205 -500
rect 32240 -535 32250 -500
rect 32285 -535 32295 -500
rect 32330 -535 32340 -500
rect 32375 -535 32385 -500
rect 32420 -535 32430 -500
rect 32465 -535 32475 -500
rect 32510 -535 32520 -500
rect 32555 -535 32565 -500
rect 32600 -535 32610 -500
rect 32645 -535 32655 -500
rect 32690 -535 32700 -500
rect 32735 -535 32745 -500
rect 32780 -535 32790 -500
rect 32825 -535 32835 -500
rect 32870 -535 32890 -500
rect 31290 -545 32890 -535
rect 31290 -580 31305 -545
rect 31340 -580 31350 -545
rect 31385 -580 31395 -545
rect 31430 -580 31440 -545
rect 31475 -580 31485 -545
rect 31520 -580 31530 -545
rect 31565 -580 31575 -545
rect 31610 -580 31620 -545
rect 31655 -580 31665 -545
rect 31700 -580 31710 -545
rect 31745 -580 31755 -545
rect 31790 -580 31800 -545
rect 31835 -580 31845 -545
rect 31880 -580 31890 -545
rect 31925 -580 31935 -545
rect 31970 -580 31980 -545
rect 32015 -580 32025 -545
rect 32060 -580 32070 -545
rect 32105 -580 32115 -545
rect 32150 -580 32160 -545
rect 32195 -580 32205 -545
rect 32240 -580 32250 -545
rect 32285 -580 32295 -545
rect 32330 -580 32340 -545
rect 32375 -580 32385 -545
rect 32420 -580 32430 -545
rect 32465 -580 32475 -545
rect 32510 -580 32520 -545
rect 32555 -580 32565 -545
rect 32600 -580 32610 -545
rect 32645 -580 32655 -545
rect 32690 -580 32700 -545
rect 32735 -580 32745 -545
rect 32780 -580 32790 -545
rect 32825 -580 32835 -545
rect 32870 -580 32890 -545
rect 31290 -590 32890 -580
rect 31290 -625 31305 -590
rect 31340 -625 31350 -590
rect 31385 -625 31395 -590
rect 31430 -625 31440 -590
rect 31475 -625 31485 -590
rect 31520 -625 31530 -590
rect 31565 -625 31575 -590
rect 31610 -625 31620 -590
rect 31655 -625 31665 -590
rect 31700 -625 31710 -590
rect 31745 -625 31755 -590
rect 31790 -625 31800 -590
rect 31835 -625 31845 -590
rect 31880 -625 31890 -590
rect 31925 -625 31935 -590
rect 31970 -625 31980 -590
rect 32015 -625 32025 -590
rect 32060 -625 32070 -590
rect 32105 -625 32115 -590
rect 32150 -625 32160 -590
rect 32195 -625 32205 -590
rect 32240 -625 32250 -590
rect 32285 -625 32295 -590
rect 32330 -625 32340 -590
rect 32375 -625 32385 -590
rect 32420 -625 32430 -590
rect 32465 -625 32475 -590
rect 32510 -625 32520 -590
rect 32555 -625 32565 -590
rect 32600 -625 32610 -590
rect 32645 -625 32655 -590
rect 32690 -625 32700 -590
rect 32735 -625 32745 -590
rect 32780 -625 32790 -590
rect 32825 -625 32835 -590
rect 32870 -625 32890 -590
rect 31290 -635 32890 -625
rect 31290 -670 31305 -635
rect 31340 -670 31350 -635
rect 31385 -670 31395 -635
rect 31430 -670 31440 -635
rect 31475 -670 31485 -635
rect 31520 -670 31530 -635
rect 31565 -670 31575 -635
rect 31610 -670 31620 -635
rect 31655 -670 31665 -635
rect 31700 -670 31710 -635
rect 31745 -670 31755 -635
rect 31790 -670 31800 -635
rect 31835 -670 31845 -635
rect 31880 -670 31890 -635
rect 31925 -670 31935 -635
rect 31970 -670 31980 -635
rect 32015 -670 32025 -635
rect 32060 -670 32070 -635
rect 32105 -670 32115 -635
rect 32150 -670 32160 -635
rect 32195 -670 32205 -635
rect 32240 -670 32250 -635
rect 32285 -670 32295 -635
rect 32330 -670 32340 -635
rect 32375 -670 32385 -635
rect 32420 -670 32430 -635
rect 32465 -670 32475 -635
rect 32510 -670 32520 -635
rect 32555 -670 32565 -635
rect 32600 -670 32610 -635
rect 32645 -670 32655 -635
rect 32690 -670 32700 -635
rect 32735 -670 32745 -635
rect 32780 -670 32790 -635
rect 32825 -670 32835 -635
rect 32870 -670 32890 -635
rect 31290 -680 32890 -670
rect 31290 -715 31305 -680
rect 31340 -715 31350 -680
rect 31385 -715 31395 -680
rect 31430 -715 31440 -680
rect 31475 -715 31485 -680
rect 31520 -715 31530 -680
rect 31565 -715 31575 -680
rect 31610 -715 31620 -680
rect 31655 -715 31665 -680
rect 31700 -715 31710 -680
rect 31745 -715 31755 -680
rect 31790 -715 31800 -680
rect 31835 -715 31845 -680
rect 31880 -715 31890 -680
rect 31925 -715 31935 -680
rect 31970 -715 31980 -680
rect 32015 -715 32025 -680
rect 32060 -715 32070 -680
rect 32105 -715 32115 -680
rect 32150 -715 32160 -680
rect 32195 -715 32205 -680
rect 32240 -715 32250 -680
rect 32285 -715 32295 -680
rect 32330 -715 32340 -680
rect 32375 -715 32385 -680
rect 32420 -715 32430 -680
rect 32465 -715 32475 -680
rect 32510 -715 32520 -680
rect 32555 -715 32565 -680
rect 32600 -715 32610 -680
rect 32645 -715 32655 -680
rect 32690 -715 32700 -680
rect 32735 -715 32745 -680
rect 32780 -715 32790 -680
rect 32825 -715 32835 -680
rect 32870 -715 32890 -680
rect 31290 -725 32890 -715
rect 31290 -760 31305 -725
rect 31340 -760 31350 -725
rect 31385 -760 31395 -725
rect 31430 -760 31440 -725
rect 31475 -760 31485 -725
rect 31520 -760 31530 -725
rect 31565 -760 31575 -725
rect 31610 -760 31620 -725
rect 31655 -760 31665 -725
rect 31700 -760 31710 -725
rect 31745 -760 31755 -725
rect 31790 -760 31800 -725
rect 31835 -760 31845 -725
rect 31880 -760 31890 -725
rect 31925 -760 31935 -725
rect 31970 -760 31980 -725
rect 32015 -760 32025 -725
rect 32060 -760 32070 -725
rect 32105 -760 32115 -725
rect 32150 -760 32160 -725
rect 32195 -760 32205 -725
rect 32240 -760 32250 -725
rect 32285 -760 32295 -725
rect 32330 -760 32340 -725
rect 32375 -760 32385 -725
rect 32420 -760 32430 -725
rect 32465 -760 32475 -725
rect 32510 -760 32520 -725
rect 32555 -760 32565 -725
rect 32600 -760 32610 -725
rect 32645 -760 32655 -725
rect 32690 -760 32700 -725
rect 32735 -760 32745 -725
rect 32780 -760 32790 -725
rect 32825 -760 32835 -725
rect 32870 -760 32890 -725
rect 31290 -770 32890 -760
rect 31290 -805 31305 -770
rect 31340 -805 31350 -770
rect 31385 -805 31395 -770
rect 31430 -805 31440 -770
rect 31475 -805 31485 -770
rect 31520 -805 31530 -770
rect 31565 -805 31575 -770
rect 31610 -805 31620 -770
rect 31655 -805 31665 -770
rect 31700 -805 31710 -770
rect 31745 -805 31755 -770
rect 31790 -805 31800 -770
rect 31835 -805 31845 -770
rect 31880 -805 31890 -770
rect 31925 -805 31935 -770
rect 31970 -805 31980 -770
rect 32015 -805 32025 -770
rect 32060 -805 32070 -770
rect 32105 -805 32115 -770
rect 32150 -805 32160 -770
rect 32195 -805 32205 -770
rect 32240 -805 32250 -770
rect 32285 -805 32295 -770
rect 32330 -805 32340 -770
rect 32375 -805 32385 -770
rect 32420 -805 32430 -770
rect 32465 -805 32475 -770
rect 32510 -805 32520 -770
rect 32555 -805 32565 -770
rect 32600 -805 32610 -770
rect 32645 -805 32655 -770
rect 32690 -805 32700 -770
rect 32735 -805 32745 -770
rect 32780 -805 32790 -770
rect 32825 -805 32835 -770
rect 32870 -805 32890 -770
rect 31290 -815 32890 -805
rect 31290 -850 31305 -815
rect 31340 -850 31350 -815
rect 31385 -850 31395 -815
rect 31430 -850 31440 -815
rect 31475 -850 31485 -815
rect 31520 -850 31530 -815
rect 31565 -850 31575 -815
rect 31610 -850 31620 -815
rect 31655 -850 31665 -815
rect 31700 -850 31710 -815
rect 31745 -850 31755 -815
rect 31790 -850 31800 -815
rect 31835 -850 31845 -815
rect 31880 -850 31890 -815
rect 31925 -850 31935 -815
rect 31970 -850 31980 -815
rect 32015 -850 32025 -815
rect 32060 -850 32070 -815
rect 32105 -850 32115 -815
rect 32150 -850 32160 -815
rect 32195 -850 32205 -815
rect 32240 -850 32250 -815
rect 32285 -850 32295 -815
rect 32330 -850 32340 -815
rect 32375 -850 32385 -815
rect 32420 -850 32430 -815
rect 32465 -850 32475 -815
rect 32510 -850 32520 -815
rect 32555 -850 32565 -815
rect 32600 -850 32610 -815
rect 32645 -850 32655 -815
rect 32690 -850 32700 -815
rect 32735 -850 32745 -815
rect 32780 -850 32790 -815
rect 32825 -850 32835 -815
rect 32870 -850 32890 -815
rect 31290 -860 32890 -850
rect 31290 -895 31305 -860
rect 31340 -895 31350 -860
rect 31385 -895 31395 -860
rect 31430 -895 31440 -860
rect 31475 -895 31485 -860
rect 31520 -895 31530 -860
rect 31565 -895 31575 -860
rect 31610 -895 31620 -860
rect 31655 -895 31665 -860
rect 31700 -895 31710 -860
rect 31745 -895 31755 -860
rect 31790 -895 31800 -860
rect 31835 -895 31845 -860
rect 31880 -895 31890 -860
rect 31925 -895 31935 -860
rect 31970 -895 31980 -860
rect 32015 -895 32025 -860
rect 32060 -895 32070 -860
rect 32105 -895 32115 -860
rect 32150 -895 32160 -860
rect 32195 -895 32205 -860
rect 32240 -895 32250 -860
rect 32285 -895 32295 -860
rect 32330 -895 32340 -860
rect 32375 -895 32385 -860
rect 32420 -895 32430 -860
rect 32465 -895 32475 -860
rect 32510 -895 32520 -860
rect 32555 -895 32565 -860
rect 32600 -895 32610 -860
rect 32645 -895 32655 -860
rect 32690 -895 32700 -860
rect 32735 -895 32745 -860
rect 32780 -895 32790 -860
rect 32825 -895 32835 -860
rect 32870 -895 32890 -860
rect 31290 -905 32890 -895
rect 31290 -940 31305 -905
rect 31340 -940 31350 -905
rect 31385 -940 31395 -905
rect 31430 -940 31440 -905
rect 31475 -940 31485 -905
rect 31520 -940 31530 -905
rect 31565 -940 31575 -905
rect 31610 -940 31620 -905
rect 31655 -940 31665 -905
rect 31700 -940 31710 -905
rect 31745 -940 31755 -905
rect 31790 -940 31800 -905
rect 31835 -940 31845 -905
rect 31880 -940 31890 -905
rect 31925 -940 31935 -905
rect 31970 -940 31980 -905
rect 32015 -940 32025 -905
rect 32060 -940 32070 -905
rect 32105 -940 32115 -905
rect 32150 -940 32160 -905
rect 32195 -940 32205 -905
rect 32240 -940 32250 -905
rect 32285 -940 32295 -905
rect 32330 -940 32340 -905
rect 32375 -940 32385 -905
rect 32420 -940 32430 -905
rect 32465 -940 32475 -905
rect 32510 -940 32520 -905
rect 32555 -940 32565 -905
rect 32600 -940 32610 -905
rect 32645 -940 32655 -905
rect 32690 -940 32700 -905
rect 32735 -940 32745 -905
rect 32780 -940 32790 -905
rect 32825 -940 32835 -905
rect 32870 -940 32890 -905
rect 31290 -950 32890 -940
rect 31290 -985 31305 -950
rect 31340 -985 31350 -950
rect 31385 -985 31395 -950
rect 31430 -985 31440 -950
rect 31475 -985 31485 -950
rect 31520 -985 31530 -950
rect 31565 -985 31575 -950
rect 31610 -985 31620 -950
rect 31655 -985 31665 -950
rect 31700 -985 31710 -950
rect 31745 -985 31755 -950
rect 31790 -985 31800 -950
rect 31835 -985 31845 -950
rect 31880 -985 31890 -950
rect 31925 -985 31935 -950
rect 31970 -985 31980 -950
rect 32015 -985 32025 -950
rect 32060 -985 32070 -950
rect 32105 -985 32115 -950
rect 32150 -985 32160 -950
rect 32195 -985 32205 -950
rect 32240 -985 32250 -950
rect 32285 -985 32295 -950
rect 32330 -985 32340 -950
rect 32375 -985 32385 -950
rect 32420 -985 32430 -950
rect 32465 -985 32475 -950
rect 32510 -985 32520 -950
rect 32555 -985 32565 -950
rect 32600 -985 32610 -950
rect 32645 -985 32655 -950
rect 32690 -985 32700 -950
rect 32735 -985 32745 -950
rect 32780 -985 32790 -950
rect 32825 -985 32835 -950
rect 32870 -985 32890 -950
rect 31290 -995 32890 -985
rect 31290 -1030 31305 -995
rect 31340 -1030 31350 -995
rect 31385 -1030 31395 -995
rect 31430 -1030 31440 -995
rect 31475 -1030 31485 -995
rect 31520 -1030 31530 -995
rect 31565 -1030 31575 -995
rect 31610 -1030 31620 -995
rect 31655 -1030 31665 -995
rect 31700 -1030 31710 -995
rect 31745 -1030 31755 -995
rect 31790 -1030 31800 -995
rect 31835 -1030 31845 -995
rect 31880 -1030 31890 -995
rect 31925 -1030 31935 -995
rect 31970 -1030 31980 -995
rect 32015 -1030 32025 -995
rect 32060 -1030 32070 -995
rect 32105 -1030 32115 -995
rect 32150 -1030 32160 -995
rect 32195 -1030 32205 -995
rect 32240 -1030 32250 -995
rect 32285 -1030 32295 -995
rect 32330 -1030 32340 -995
rect 32375 -1030 32385 -995
rect 32420 -1030 32430 -995
rect 32465 -1030 32475 -995
rect 32510 -1030 32520 -995
rect 32555 -1030 32565 -995
rect 32600 -1030 32610 -995
rect 32645 -1030 32655 -995
rect 32690 -1030 32700 -995
rect 32735 -1030 32745 -995
rect 32780 -1030 32790 -995
rect 32825 -1030 32835 -995
rect 32870 -1030 32890 -995
rect 31290 -1040 32890 -1030
rect 31290 -1075 31305 -1040
rect 31340 -1075 31350 -1040
rect 31385 -1075 31395 -1040
rect 31430 -1075 31440 -1040
rect 31475 -1075 31485 -1040
rect 31520 -1075 31530 -1040
rect 31565 -1075 31575 -1040
rect 31610 -1075 31620 -1040
rect 31655 -1075 31665 -1040
rect 31700 -1075 31710 -1040
rect 31745 -1075 31755 -1040
rect 31790 -1075 31800 -1040
rect 31835 -1075 31845 -1040
rect 31880 -1075 31890 -1040
rect 31925 -1075 31935 -1040
rect 31970 -1075 31980 -1040
rect 32015 -1075 32025 -1040
rect 32060 -1075 32070 -1040
rect 32105 -1075 32115 -1040
rect 32150 -1075 32160 -1040
rect 32195 -1075 32205 -1040
rect 32240 -1075 32250 -1040
rect 32285 -1075 32295 -1040
rect 32330 -1075 32340 -1040
rect 32375 -1075 32385 -1040
rect 32420 -1075 32430 -1040
rect 32465 -1075 32475 -1040
rect 32510 -1075 32520 -1040
rect 32555 -1075 32565 -1040
rect 32600 -1075 32610 -1040
rect 32645 -1075 32655 -1040
rect 32690 -1075 32700 -1040
rect 32735 -1075 32745 -1040
rect 32780 -1075 32790 -1040
rect 32825 -1075 32835 -1040
rect 32870 -1075 32890 -1040
rect 31290 -1085 32890 -1075
rect 31290 -1120 31305 -1085
rect 31340 -1120 31350 -1085
rect 31385 -1120 31395 -1085
rect 31430 -1120 31440 -1085
rect 31475 -1120 31485 -1085
rect 31520 -1120 31530 -1085
rect 31565 -1120 31575 -1085
rect 31610 -1120 31620 -1085
rect 31655 -1120 31665 -1085
rect 31700 -1120 31710 -1085
rect 31745 -1120 31755 -1085
rect 31790 -1120 31800 -1085
rect 31835 -1120 31845 -1085
rect 31880 -1120 31890 -1085
rect 31925 -1120 31935 -1085
rect 31970 -1120 31980 -1085
rect 32015 -1120 32025 -1085
rect 32060 -1120 32070 -1085
rect 32105 -1120 32115 -1085
rect 32150 -1120 32160 -1085
rect 32195 -1120 32205 -1085
rect 32240 -1120 32250 -1085
rect 32285 -1120 32295 -1085
rect 32330 -1120 32340 -1085
rect 32375 -1120 32385 -1085
rect 32420 -1120 32430 -1085
rect 32465 -1120 32475 -1085
rect 32510 -1120 32520 -1085
rect 32555 -1120 32565 -1085
rect 32600 -1120 32610 -1085
rect 32645 -1120 32655 -1085
rect 32690 -1120 32700 -1085
rect 32735 -1120 32745 -1085
rect 32780 -1120 32790 -1085
rect 32825 -1120 32835 -1085
rect 32870 -1120 32890 -1085
rect 31290 -1130 32890 -1120
rect 31290 -1165 31305 -1130
rect 31340 -1165 31350 -1130
rect 31385 -1165 31395 -1130
rect 31430 -1165 31440 -1130
rect 31475 -1165 31485 -1130
rect 31520 -1165 31530 -1130
rect 31565 -1165 31575 -1130
rect 31610 -1165 31620 -1130
rect 31655 -1165 31665 -1130
rect 31700 -1165 31710 -1130
rect 31745 -1165 31755 -1130
rect 31790 -1165 31800 -1130
rect 31835 -1165 31845 -1130
rect 31880 -1165 31890 -1130
rect 31925 -1165 31935 -1130
rect 31970 -1165 31980 -1130
rect 32015 -1165 32025 -1130
rect 32060 -1165 32070 -1130
rect 32105 -1165 32115 -1130
rect 32150 -1165 32160 -1130
rect 32195 -1165 32205 -1130
rect 32240 -1165 32250 -1130
rect 32285 -1165 32295 -1130
rect 32330 -1165 32340 -1130
rect 32375 -1165 32385 -1130
rect 32420 -1165 32430 -1130
rect 32465 -1165 32475 -1130
rect 32510 -1165 32520 -1130
rect 32555 -1165 32565 -1130
rect 32600 -1165 32610 -1130
rect 32645 -1165 32655 -1130
rect 32690 -1165 32700 -1130
rect 32735 -1165 32745 -1130
rect 32780 -1165 32790 -1130
rect 32825 -1165 32835 -1130
rect 32870 -1165 32890 -1130
rect 31290 -1175 32890 -1165
rect 31290 -1210 31305 -1175
rect 31340 -1210 31350 -1175
rect 31385 -1210 31395 -1175
rect 31430 -1210 31440 -1175
rect 31475 -1210 31485 -1175
rect 31520 -1210 31530 -1175
rect 31565 -1210 31575 -1175
rect 31610 -1210 31620 -1175
rect 31655 -1210 31665 -1175
rect 31700 -1210 31710 -1175
rect 31745 -1210 31755 -1175
rect 31790 -1210 31800 -1175
rect 31835 -1210 31845 -1175
rect 31880 -1210 31890 -1175
rect 31925 -1210 31935 -1175
rect 31970 -1210 31980 -1175
rect 32015 -1210 32025 -1175
rect 32060 -1210 32070 -1175
rect 32105 -1210 32115 -1175
rect 32150 -1210 32160 -1175
rect 32195 -1210 32205 -1175
rect 32240 -1210 32250 -1175
rect 32285 -1210 32295 -1175
rect 32330 -1210 32340 -1175
rect 32375 -1210 32385 -1175
rect 32420 -1210 32430 -1175
rect 32465 -1210 32475 -1175
rect 32510 -1210 32520 -1175
rect 32555 -1210 32565 -1175
rect 32600 -1210 32610 -1175
rect 32645 -1210 32655 -1175
rect 32690 -1210 32700 -1175
rect 32735 -1210 32745 -1175
rect 32780 -1210 32790 -1175
rect 32825 -1210 32835 -1175
rect 32870 -1210 32890 -1175
rect 31290 -1220 32890 -1210
rect 31290 -1255 31305 -1220
rect 31340 -1255 31350 -1220
rect 31385 -1255 31395 -1220
rect 31430 -1255 31440 -1220
rect 31475 -1255 31485 -1220
rect 31520 -1255 31530 -1220
rect 31565 -1255 31575 -1220
rect 31610 -1255 31620 -1220
rect 31655 -1255 31665 -1220
rect 31700 -1255 31710 -1220
rect 31745 -1255 31755 -1220
rect 31790 -1255 31800 -1220
rect 31835 -1255 31845 -1220
rect 31880 -1255 31890 -1220
rect 31925 -1255 31935 -1220
rect 31970 -1255 31980 -1220
rect 32015 -1255 32025 -1220
rect 32060 -1255 32070 -1220
rect 32105 -1255 32115 -1220
rect 32150 -1255 32160 -1220
rect 32195 -1255 32205 -1220
rect 32240 -1255 32250 -1220
rect 32285 -1255 32295 -1220
rect 32330 -1255 32340 -1220
rect 32375 -1255 32385 -1220
rect 32420 -1255 32430 -1220
rect 32465 -1255 32475 -1220
rect 32510 -1255 32520 -1220
rect 32555 -1255 32565 -1220
rect 32600 -1255 32610 -1220
rect 32645 -1255 32655 -1220
rect 32690 -1255 32700 -1220
rect 32735 -1255 32745 -1220
rect 32780 -1255 32790 -1220
rect 32825 -1255 32835 -1220
rect 32870 -1255 32890 -1220
rect 31290 -1265 32890 -1255
rect 31290 -1300 31305 -1265
rect 31340 -1300 31350 -1265
rect 31385 -1300 31395 -1265
rect 31430 -1300 31440 -1265
rect 31475 -1300 31485 -1265
rect 31520 -1300 31530 -1265
rect 31565 -1300 31575 -1265
rect 31610 -1300 31620 -1265
rect 31655 -1300 31665 -1265
rect 31700 -1300 31710 -1265
rect 31745 -1300 31755 -1265
rect 31790 -1300 31800 -1265
rect 31835 -1300 31845 -1265
rect 31880 -1300 31890 -1265
rect 31925 -1300 31935 -1265
rect 31970 -1300 31980 -1265
rect 32015 -1300 32025 -1265
rect 32060 -1300 32070 -1265
rect 32105 -1300 32115 -1265
rect 32150 -1300 32160 -1265
rect 32195 -1300 32205 -1265
rect 32240 -1300 32250 -1265
rect 32285 -1300 32295 -1265
rect 32330 -1300 32340 -1265
rect 32375 -1300 32385 -1265
rect 32420 -1300 32430 -1265
rect 32465 -1300 32475 -1265
rect 32510 -1300 32520 -1265
rect 32555 -1300 32565 -1265
rect 32600 -1300 32610 -1265
rect 32645 -1300 32655 -1265
rect 32690 -1300 32700 -1265
rect 32735 -1300 32745 -1265
rect 32780 -1300 32790 -1265
rect 32825 -1300 32835 -1265
rect 32870 -1300 32890 -1265
rect 31290 -1310 32890 -1300
rect 31290 -1345 31305 -1310
rect 31340 -1345 31350 -1310
rect 31385 -1345 31395 -1310
rect 31430 -1345 31440 -1310
rect 31475 -1345 31485 -1310
rect 31520 -1345 31530 -1310
rect 31565 -1345 31575 -1310
rect 31610 -1345 31620 -1310
rect 31655 -1345 31665 -1310
rect 31700 -1345 31710 -1310
rect 31745 -1345 31755 -1310
rect 31790 -1345 31800 -1310
rect 31835 -1345 31845 -1310
rect 31880 -1345 31890 -1310
rect 31925 -1345 31935 -1310
rect 31970 -1345 31980 -1310
rect 32015 -1345 32025 -1310
rect 32060 -1345 32070 -1310
rect 32105 -1345 32115 -1310
rect 32150 -1345 32160 -1310
rect 32195 -1345 32205 -1310
rect 32240 -1345 32250 -1310
rect 32285 -1345 32295 -1310
rect 32330 -1345 32340 -1310
rect 32375 -1345 32385 -1310
rect 32420 -1345 32430 -1310
rect 32465 -1345 32475 -1310
rect 32510 -1345 32520 -1310
rect 32555 -1345 32565 -1310
rect 32600 -1345 32610 -1310
rect 32645 -1345 32655 -1310
rect 32690 -1345 32700 -1310
rect 32735 -1345 32745 -1310
rect 32780 -1345 32790 -1310
rect 32825 -1345 32835 -1310
rect 32870 -1345 32890 -1310
rect 31290 -1360 32890 -1345
<< via3 >>
rect 2110 19310 2150 19315
rect 2110 19280 2115 19310
rect 2115 19280 2145 19310
rect 2145 19280 2150 19310
rect 2110 19275 2150 19280
rect 2110 19245 2150 19250
rect 2110 19215 2115 19245
rect 2115 19215 2145 19245
rect 2145 19215 2150 19245
rect 2110 19210 2150 19215
rect 2110 19175 2150 19180
rect 2110 19145 2115 19175
rect 2115 19145 2145 19175
rect 2145 19145 2150 19175
rect 2110 19140 2150 19145
rect 2110 19105 2150 19110
rect 2110 19075 2115 19105
rect 2115 19075 2145 19105
rect 2145 19075 2150 19105
rect 2110 19070 2150 19075
rect 2110 19035 2150 19040
rect 2110 19005 2115 19035
rect 2115 19005 2145 19035
rect 2145 19005 2150 19035
rect 2110 19000 2150 19005
rect 2110 18970 2150 18975
rect 2110 18940 2115 18970
rect 2115 18940 2145 18970
rect 2145 18940 2150 18970
rect 2110 18935 2150 18940
rect 2110 18910 2150 18915
rect 2110 18880 2115 18910
rect 2115 18880 2145 18910
rect 2145 18880 2150 18910
rect 2110 18875 2150 18880
rect 2110 18845 2150 18850
rect 2110 18815 2115 18845
rect 2115 18815 2145 18845
rect 2145 18815 2150 18845
rect 2110 18810 2150 18815
rect 2110 18775 2150 18780
rect 2110 18745 2115 18775
rect 2115 18745 2145 18775
rect 2145 18745 2150 18775
rect 2110 18740 2150 18745
rect 2110 18705 2150 18710
rect 2110 18675 2115 18705
rect 2115 18675 2145 18705
rect 2145 18675 2150 18705
rect 2110 18670 2150 18675
rect 2110 18635 2150 18640
rect 2110 18605 2115 18635
rect 2115 18605 2145 18635
rect 2145 18605 2150 18635
rect 2110 18600 2150 18605
rect 2110 18570 2150 18575
rect 2110 18540 2115 18570
rect 2115 18540 2145 18570
rect 2145 18540 2150 18570
rect 2110 18535 2150 18540
rect 2110 18510 2150 18515
rect 2110 18480 2115 18510
rect 2115 18480 2145 18510
rect 2145 18480 2150 18510
rect 2110 18475 2150 18480
rect 2110 18445 2150 18450
rect 2110 18415 2115 18445
rect 2115 18415 2145 18445
rect 2145 18415 2150 18445
rect 2110 18410 2150 18415
rect 2110 18375 2150 18380
rect 2110 18345 2115 18375
rect 2115 18345 2145 18375
rect 2145 18345 2150 18375
rect 2110 18340 2150 18345
rect 2110 18305 2150 18310
rect 2110 18275 2115 18305
rect 2115 18275 2145 18305
rect 2145 18275 2150 18305
rect 2110 18270 2150 18275
rect 2110 18235 2150 18240
rect 2110 18205 2115 18235
rect 2115 18205 2145 18235
rect 2145 18205 2150 18235
rect 2110 18200 2150 18205
rect 2110 18170 2150 18175
rect 2110 18140 2115 18170
rect 2115 18140 2145 18170
rect 2145 18140 2150 18170
rect 2110 18135 2150 18140
rect 2110 18110 2150 18115
rect 2110 18080 2115 18110
rect 2115 18080 2145 18110
rect 2145 18080 2150 18110
rect 2110 18075 2150 18080
rect 2110 18045 2150 18050
rect 2110 18015 2115 18045
rect 2115 18015 2145 18045
rect 2145 18015 2150 18045
rect 2110 18010 2150 18015
rect 2110 17975 2150 17980
rect 2110 17945 2115 17975
rect 2115 17945 2145 17975
rect 2145 17945 2150 17975
rect 2110 17940 2150 17945
rect 2110 17905 2150 17910
rect 2110 17875 2115 17905
rect 2115 17875 2145 17905
rect 2145 17875 2150 17905
rect 2110 17870 2150 17875
rect 2110 17835 2150 17840
rect 2110 17805 2115 17835
rect 2115 17805 2145 17835
rect 2145 17805 2150 17835
rect 2110 17800 2150 17805
rect 2110 17770 2150 17775
rect 2110 17740 2115 17770
rect 2115 17740 2145 17770
rect 2145 17740 2150 17770
rect 2110 17735 2150 17740
rect 6700 19310 6740 19315
rect 6700 19280 6705 19310
rect 6705 19280 6735 19310
rect 6735 19280 6740 19310
rect 6700 19275 6740 19280
rect 6700 19245 6740 19250
rect 6700 19215 6705 19245
rect 6705 19215 6735 19245
rect 6735 19215 6740 19245
rect 6700 19210 6740 19215
rect 6700 19175 6740 19180
rect 6700 19145 6705 19175
rect 6705 19145 6735 19175
rect 6735 19145 6740 19175
rect 6700 19140 6740 19145
rect 6700 19105 6740 19110
rect 6700 19075 6705 19105
rect 6705 19075 6735 19105
rect 6735 19075 6740 19105
rect 6700 19070 6740 19075
rect 6700 19035 6740 19040
rect 6700 19005 6705 19035
rect 6705 19005 6735 19035
rect 6735 19005 6740 19035
rect 6700 19000 6740 19005
rect 6700 18970 6740 18975
rect 6700 18940 6705 18970
rect 6705 18940 6735 18970
rect 6735 18940 6740 18970
rect 6700 18935 6740 18940
rect 6700 18910 6740 18915
rect 6700 18880 6705 18910
rect 6705 18880 6735 18910
rect 6735 18880 6740 18910
rect 6700 18875 6740 18880
rect 6700 18845 6740 18850
rect 6700 18815 6705 18845
rect 6705 18815 6735 18845
rect 6735 18815 6740 18845
rect 6700 18810 6740 18815
rect 6700 18775 6740 18780
rect 6700 18745 6705 18775
rect 6705 18745 6735 18775
rect 6735 18745 6740 18775
rect 6700 18740 6740 18745
rect 6700 18705 6740 18710
rect 6700 18675 6705 18705
rect 6705 18675 6735 18705
rect 6735 18675 6740 18705
rect 6700 18670 6740 18675
rect 6700 18635 6740 18640
rect 6700 18605 6705 18635
rect 6705 18605 6735 18635
rect 6735 18605 6740 18635
rect 6700 18600 6740 18605
rect 6700 18570 6740 18575
rect 6700 18540 6705 18570
rect 6705 18540 6735 18570
rect 6735 18540 6740 18570
rect 6700 18535 6740 18540
rect 6700 18510 6740 18515
rect 6700 18480 6705 18510
rect 6705 18480 6735 18510
rect 6735 18480 6740 18510
rect 6700 18475 6740 18480
rect 6700 18445 6740 18450
rect 6700 18415 6705 18445
rect 6705 18415 6735 18445
rect 6735 18415 6740 18445
rect 6700 18410 6740 18415
rect 6700 18375 6740 18380
rect 6700 18345 6705 18375
rect 6705 18345 6735 18375
rect 6735 18345 6740 18375
rect 6700 18340 6740 18345
rect 6700 18305 6740 18310
rect 6700 18275 6705 18305
rect 6705 18275 6735 18305
rect 6735 18275 6740 18305
rect 6700 18270 6740 18275
rect 6700 18235 6740 18240
rect 6700 18205 6705 18235
rect 6705 18205 6735 18235
rect 6735 18205 6740 18235
rect 6700 18200 6740 18205
rect 6700 18170 6740 18175
rect 6700 18140 6705 18170
rect 6705 18140 6735 18170
rect 6735 18140 6740 18170
rect 6700 18135 6740 18140
rect 6700 18110 6740 18115
rect 6700 18080 6705 18110
rect 6705 18080 6735 18110
rect 6735 18080 6740 18110
rect 6700 18075 6740 18080
rect 6700 18045 6740 18050
rect 6700 18015 6705 18045
rect 6705 18015 6735 18045
rect 6735 18015 6740 18045
rect 6700 18010 6740 18015
rect 6700 17975 6740 17980
rect 6700 17945 6705 17975
rect 6705 17945 6735 17975
rect 6735 17945 6740 17975
rect 6700 17940 6740 17945
rect 6700 17905 6740 17910
rect 6700 17875 6705 17905
rect 6705 17875 6735 17905
rect 6735 17875 6740 17905
rect 6700 17870 6740 17875
rect 6700 17835 6740 17840
rect 6700 17805 6705 17835
rect 6705 17805 6735 17835
rect 6735 17805 6740 17835
rect 6700 17800 6740 17805
rect 6700 17770 6740 17775
rect 6700 17740 6705 17770
rect 6705 17740 6735 17770
rect 6735 17740 6740 17770
rect 6700 17735 6740 17740
rect 31305 19270 31340 19305
rect 31350 19270 31385 19305
rect 31395 19270 31430 19305
rect 31440 19270 31475 19305
rect 31485 19270 31520 19305
rect 31530 19270 31565 19305
rect 31575 19270 31610 19305
rect 31620 19270 31655 19305
rect 31665 19270 31700 19305
rect 31710 19270 31745 19305
rect 31755 19270 31790 19305
rect 31800 19270 31835 19305
rect 31845 19270 31880 19305
rect 31890 19270 31925 19305
rect 31935 19270 31970 19305
rect 31980 19270 32015 19305
rect 32025 19270 32060 19305
rect 32070 19270 32105 19305
rect 32115 19270 32150 19305
rect 32160 19270 32195 19305
rect 32205 19270 32240 19305
rect 32250 19270 32285 19305
rect 32295 19270 32330 19305
rect 32340 19270 32375 19305
rect 32385 19270 32420 19305
rect 32430 19270 32465 19305
rect 32475 19270 32510 19305
rect 32520 19270 32555 19305
rect 32565 19270 32600 19305
rect 32610 19270 32645 19305
rect 32655 19270 32690 19305
rect 32700 19270 32735 19305
rect 32745 19270 32780 19305
rect 32790 19270 32825 19305
rect 32835 19270 32870 19305
rect 31305 19225 31340 19260
rect 31350 19225 31385 19260
rect 31395 19225 31430 19260
rect 31440 19225 31475 19260
rect 31485 19225 31520 19260
rect 31530 19225 31565 19260
rect 31575 19225 31610 19260
rect 31620 19225 31655 19260
rect 31665 19225 31700 19260
rect 31710 19225 31745 19260
rect 31755 19225 31790 19260
rect 31800 19225 31835 19260
rect 31845 19225 31880 19260
rect 31890 19225 31925 19260
rect 31935 19225 31970 19260
rect 31980 19225 32015 19260
rect 32025 19225 32060 19260
rect 32070 19225 32105 19260
rect 32115 19225 32150 19260
rect 32160 19225 32195 19260
rect 32205 19225 32240 19260
rect 32250 19225 32285 19260
rect 32295 19225 32330 19260
rect 32340 19225 32375 19260
rect 32385 19225 32420 19260
rect 32430 19225 32465 19260
rect 32475 19225 32510 19260
rect 32520 19225 32555 19260
rect 32565 19225 32600 19260
rect 32610 19225 32645 19260
rect 32655 19225 32690 19260
rect 32700 19225 32735 19260
rect 32745 19225 32780 19260
rect 32790 19225 32825 19260
rect 32835 19225 32870 19260
rect 31305 19180 31340 19215
rect 31350 19180 31385 19215
rect 31395 19180 31430 19215
rect 31440 19180 31475 19215
rect 31485 19180 31520 19215
rect 31530 19180 31565 19215
rect 31575 19180 31610 19215
rect 31620 19180 31655 19215
rect 31665 19180 31700 19215
rect 31710 19180 31745 19215
rect 31755 19180 31790 19215
rect 31800 19180 31835 19215
rect 31845 19180 31880 19215
rect 31890 19180 31925 19215
rect 31935 19180 31970 19215
rect 31980 19180 32015 19215
rect 32025 19180 32060 19215
rect 32070 19180 32105 19215
rect 32115 19180 32150 19215
rect 32160 19180 32195 19215
rect 32205 19180 32240 19215
rect 32250 19180 32285 19215
rect 32295 19180 32330 19215
rect 32340 19180 32375 19215
rect 32385 19180 32420 19215
rect 32430 19180 32465 19215
rect 32475 19180 32510 19215
rect 32520 19180 32555 19215
rect 32565 19180 32600 19215
rect 32610 19180 32645 19215
rect 32655 19180 32690 19215
rect 32700 19180 32735 19215
rect 32745 19180 32780 19215
rect 32790 19180 32825 19215
rect 32835 19180 32870 19215
rect 31305 19135 31340 19170
rect 31350 19135 31385 19170
rect 31395 19135 31430 19170
rect 31440 19135 31475 19170
rect 31485 19135 31520 19170
rect 31530 19135 31565 19170
rect 31575 19135 31610 19170
rect 31620 19135 31655 19170
rect 31665 19135 31700 19170
rect 31710 19135 31745 19170
rect 31755 19135 31790 19170
rect 31800 19135 31835 19170
rect 31845 19135 31880 19170
rect 31890 19135 31925 19170
rect 31935 19135 31970 19170
rect 31980 19135 32015 19170
rect 32025 19135 32060 19170
rect 32070 19135 32105 19170
rect 32115 19135 32150 19170
rect 32160 19135 32195 19170
rect 32205 19135 32240 19170
rect 32250 19135 32285 19170
rect 32295 19135 32330 19170
rect 32340 19135 32375 19170
rect 32385 19135 32420 19170
rect 32430 19135 32465 19170
rect 32475 19135 32510 19170
rect 32520 19135 32555 19170
rect 32565 19135 32600 19170
rect 32610 19135 32645 19170
rect 32655 19135 32690 19170
rect 32700 19135 32735 19170
rect 32745 19135 32780 19170
rect 32790 19135 32825 19170
rect 32835 19135 32870 19170
rect 31305 19090 31340 19125
rect 31350 19090 31385 19125
rect 31395 19090 31430 19125
rect 31440 19090 31475 19125
rect 31485 19090 31520 19125
rect 31530 19090 31565 19125
rect 31575 19090 31610 19125
rect 31620 19090 31655 19125
rect 31665 19090 31700 19125
rect 31710 19090 31745 19125
rect 31755 19090 31790 19125
rect 31800 19090 31835 19125
rect 31845 19090 31880 19125
rect 31890 19090 31925 19125
rect 31935 19090 31970 19125
rect 31980 19090 32015 19125
rect 32025 19090 32060 19125
rect 32070 19090 32105 19125
rect 32115 19090 32150 19125
rect 32160 19090 32195 19125
rect 32205 19090 32240 19125
rect 32250 19090 32285 19125
rect 32295 19090 32330 19125
rect 32340 19090 32375 19125
rect 32385 19090 32420 19125
rect 32430 19090 32465 19125
rect 32475 19090 32510 19125
rect 32520 19090 32555 19125
rect 32565 19090 32600 19125
rect 32610 19090 32645 19125
rect 32655 19090 32690 19125
rect 32700 19090 32735 19125
rect 32745 19090 32780 19125
rect 32790 19090 32825 19125
rect 32835 19090 32870 19125
rect 31305 19045 31340 19080
rect 31350 19045 31385 19080
rect 31395 19045 31430 19080
rect 31440 19045 31475 19080
rect 31485 19045 31520 19080
rect 31530 19045 31565 19080
rect 31575 19045 31610 19080
rect 31620 19045 31655 19080
rect 31665 19045 31700 19080
rect 31710 19045 31745 19080
rect 31755 19045 31790 19080
rect 31800 19045 31835 19080
rect 31845 19045 31880 19080
rect 31890 19045 31925 19080
rect 31935 19045 31970 19080
rect 31980 19045 32015 19080
rect 32025 19045 32060 19080
rect 32070 19045 32105 19080
rect 32115 19045 32150 19080
rect 32160 19045 32195 19080
rect 32205 19045 32240 19080
rect 32250 19045 32285 19080
rect 32295 19045 32330 19080
rect 32340 19045 32375 19080
rect 32385 19045 32420 19080
rect 32430 19045 32465 19080
rect 32475 19045 32510 19080
rect 32520 19045 32555 19080
rect 32565 19045 32600 19080
rect 32610 19045 32645 19080
rect 32655 19045 32690 19080
rect 32700 19045 32735 19080
rect 32745 19045 32780 19080
rect 32790 19045 32825 19080
rect 32835 19045 32870 19080
rect 31305 19000 31340 19035
rect 31350 19000 31385 19035
rect 31395 19000 31430 19035
rect 31440 19000 31475 19035
rect 31485 19000 31520 19035
rect 31530 19000 31565 19035
rect 31575 19000 31610 19035
rect 31620 19000 31655 19035
rect 31665 19000 31700 19035
rect 31710 19000 31745 19035
rect 31755 19000 31790 19035
rect 31800 19000 31835 19035
rect 31845 19000 31880 19035
rect 31890 19000 31925 19035
rect 31935 19000 31970 19035
rect 31980 19000 32015 19035
rect 32025 19000 32060 19035
rect 32070 19000 32105 19035
rect 32115 19000 32150 19035
rect 32160 19000 32195 19035
rect 32205 19000 32240 19035
rect 32250 19000 32285 19035
rect 32295 19000 32330 19035
rect 32340 19000 32375 19035
rect 32385 19000 32420 19035
rect 32430 19000 32465 19035
rect 32475 19000 32510 19035
rect 32520 19000 32555 19035
rect 32565 19000 32600 19035
rect 32610 19000 32645 19035
rect 32655 19000 32690 19035
rect 32700 19000 32735 19035
rect 32745 19000 32780 19035
rect 32790 19000 32825 19035
rect 32835 19000 32870 19035
rect 31305 18955 31340 18990
rect 31350 18955 31385 18990
rect 31395 18955 31430 18990
rect 31440 18955 31475 18990
rect 31485 18955 31520 18990
rect 31530 18955 31565 18990
rect 31575 18955 31610 18990
rect 31620 18955 31655 18990
rect 31665 18955 31700 18990
rect 31710 18955 31745 18990
rect 31755 18955 31790 18990
rect 31800 18955 31835 18990
rect 31845 18955 31880 18990
rect 31890 18955 31925 18990
rect 31935 18955 31970 18990
rect 31980 18955 32015 18990
rect 32025 18955 32060 18990
rect 32070 18955 32105 18990
rect 32115 18955 32150 18990
rect 32160 18955 32195 18990
rect 32205 18955 32240 18990
rect 32250 18955 32285 18990
rect 32295 18955 32330 18990
rect 32340 18955 32375 18990
rect 32385 18955 32420 18990
rect 32430 18955 32465 18990
rect 32475 18955 32510 18990
rect 32520 18955 32555 18990
rect 32565 18955 32600 18990
rect 32610 18955 32645 18990
rect 32655 18955 32690 18990
rect 32700 18955 32735 18990
rect 32745 18955 32780 18990
rect 32790 18955 32825 18990
rect 32835 18955 32870 18990
rect 31305 18910 31340 18945
rect 31350 18910 31385 18945
rect 31395 18910 31430 18945
rect 31440 18910 31475 18945
rect 31485 18910 31520 18945
rect 31530 18910 31565 18945
rect 31575 18910 31610 18945
rect 31620 18910 31655 18945
rect 31665 18910 31700 18945
rect 31710 18910 31745 18945
rect 31755 18910 31790 18945
rect 31800 18910 31835 18945
rect 31845 18910 31880 18945
rect 31890 18910 31925 18945
rect 31935 18910 31970 18945
rect 31980 18910 32015 18945
rect 32025 18910 32060 18945
rect 32070 18910 32105 18945
rect 32115 18910 32150 18945
rect 32160 18910 32195 18945
rect 32205 18910 32240 18945
rect 32250 18910 32285 18945
rect 32295 18910 32330 18945
rect 32340 18910 32375 18945
rect 32385 18910 32420 18945
rect 32430 18910 32465 18945
rect 32475 18910 32510 18945
rect 32520 18910 32555 18945
rect 32565 18910 32600 18945
rect 32610 18910 32645 18945
rect 32655 18910 32690 18945
rect 32700 18910 32735 18945
rect 32745 18910 32780 18945
rect 32790 18910 32825 18945
rect 32835 18910 32870 18945
rect 31305 18865 31340 18900
rect 31350 18865 31385 18900
rect 31395 18865 31430 18900
rect 31440 18865 31475 18900
rect 31485 18865 31520 18900
rect 31530 18865 31565 18900
rect 31575 18865 31610 18900
rect 31620 18865 31655 18900
rect 31665 18865 31700 18900
rect 31710 18865 31745 18900
rect 31755 18865 31790 18900
rect 31800 18865 31835 18900
rect 31845 18865 31880 18900
rect 31890 18865 31925 18900
rect 31935 18865 31970 18900
rect 31980 18865 32015 18900
rect 32025 18865 32060 18900
rect 32070 18865 32105 18900
rect 32115 18865 32150 18900
rect 32160 18865 32195 18900
rect 32205 18865 32240 18900
rect 32250 18865 32285 18900
rect 32295 18865 32330 18900
rect 32340 18865 32375 18900
rect 32385 18865 32420 18900
rect 32430 18865 32465 18900
rect 32475 18865 32510 18900
rect 32520 18865 32555 18900
rect 32565 18865 32600 18900
rect 32610 18865 32645 18900
rect 32655 18865 32690 18900
rect 32700 18865 32735 18900
rect 32745 18865 32780 18900
rect 32790 18865 32825 18900
rect 32835 18865 32870 18900
rect 31305 18820 31340 18855
rect 31350 18820 31385 18855
rect 31395 18820 31430 18855
rect 31440 18820 31475 18855
rect 31485 18820 31520 18855
rect 31530 18820 31565 18855
rect 31575 18820 31610 18855
rect 31620 18820 31655 18855
rect 31665 18820 31700 18855
rect 31710 18820 31745 18855
rect 31755 18820 31790 18855
rect 31800 18820 31835 18855
rect 31845 18820 31880 18855
rect 31890 18820 31925 18855
rect 31935 18820 31970 18855
rect 31980 18820 32015 18855
rect 32025 18820 32060 18855
rect 32070 18820 32105 18855
rect 32115 18820 32150 18855
rect 32160 18820 32195 18855
rect 32205 18820 32240 18855
rect 32250 18820 32285 18855
rect 32295 18820 32330 18855
rect 32340 18820 32375 18855
rect 32385 18820 32420 18855
rect 32430 18820 32465 18855
rect 32475 18820 32510 18855
rect 32520 18820 32555 18855
rect 32565 18820 32600 18855
rect 32610 18820 32645 18855
rect 32655 18820 32690 18855
rect 32700 18820 32735 18855
rect 32745 18820 32780 18855
rect 32790 18820 32825 18855
rect 32835 18820 32870 18855
rect 31305 18775 31340 18810
rect 31350 18775 31385 18810
rect 31395 18775 31430 18810
rect 31440 18775 31475 18810
rect 31485 18775 31520 18810
rect 31530 18775 31565 18810
rect 31575 18775 31610 18810
rect 31620 18775 31655 18810
rect 31665 18775 31700 18810
rect 31710 18775 31745 18810
rect 31755 18775 31790 18810
rect 31800 18775 31835 18810
rect 31845 18775 31880 18810
rect 31890 18775 31925 18810
rect 31935 18775 31970 18810
rect 31980 18775 32015 18810
rect 32025 18775 32060 18810
rect 32070 18775 32105 18810
rect 32115 18775 32150 18810
rect 32160 18775 32195 18810
rect 32205 18775 32240 18810
rect 32250 18775 32285 18810
rect 32295 18775 32330 18810
rect 32340 18775 32375 18810
rect 32385 18775 32420 18810
rect 32430 18775 32465 18810
rect 32475 18775 32510 18810
rect 32520 18775 32555 18810
rect 32565 18775 32600 18810
rect 32610 18775 32645 18810
rect 32655 18775 32690 18810
rect 32700 18775 32735 18810
rect 32745 18775 32780 18810
rect 32790 18775 32825 18810
rect 32835 18775 32870 18810
rect 31305 18730 31340 18765
rect 31350 18730 31385 18765
rect 31395 18730 31430 18765
rect 31440 18730 31475 18765
rect 31485 18730 31520 18765
rect 31530 18730 31565 18765
rect 31575 18730 31610 18765
rect 31620 18730 31655 18765
rect 31665 18730 31700 18765
rect 31710 18730 31745 18765
rect 31755 18730 31790 18765
rect 31800 18730 31835 18765
rect 31845 18730 31880 18765
rect 31890 18730 31925 18765
rect 31935 18730 31970 18765
rect 31980 18730 32015 18765
rect 32025 18730 32060 18765
rect 32070 18730 32105 18765
rect 32115 18730 32150 18765
rect 32160 18730 32195 18765
rect 32205 18730 32240 18765
rect 32250 18730 32285 18765
rect 32295 18730 32330 18765
rect 32340 18730 32375 18765
rect 32385 18730 32420 18765
rect 32430 18730 32465 18765
rect 32475 18730 32510 18765
rect 32520 18730 32555 18765
rect 32565 18730 32600 18765
rect 32610 18730 32645 18765
rect 32655 18730 32690 18765
rect 32700 18730 32735 18765
rect 32745 18730 32780 18765
rect 32790 18730 32825 18765
rect 32835 18730 32870 18765
rect 31305 18685 31340 18720
rect 31350 18685 31385 18720
rect 31395 18685 31430 18720
rect 31440 18685 31475 18720
rect 31485 18685 31520 18720
rect 31530 18685 31565 18720
rect 31575 18685 31610 18720
rect 31620 18685 31655 18720
rect 31665 18685 31700 18720
rect 31710 18685 31745 18720
rect 31755 18685 31790 18720
rect 31800 18685 31835 18720
rect 31845 18685 31880 18720
rect 31890 18685 31925 18720
rect 31935 18685 31970 18720
rect 31980 18685 32015 18720
rect 32025 18685 32060 18720
rect 32070 18685 32105 18720
rect 32115 18685 32150 18720
rect 32160 18685 32195 18720
rect 32205 18685 32240 18720
rect 32250 18685 32285 18720
rect 32295 18685 32330 18720
rect 32340 18685 32375 18720
rect 32385 18685 32420 18720
rect 32430 18685 32465 18720
rect 32475 18685 32510 18720
rect 32520 18685 32555 18720
rect 32565 18685 32600 18720
rect 32610 18685 32645 18720
rect 32655 18685 32690 18720
rect 32700 18685 32735 18720
rect 32745 18685 32780 18720
rect 32790 18685 32825 18720
rect 32835 18685 32870 18720
rect 31305 18640 31340 18675
rect 31350 18640 31385 18675
rect 31395 18640 31430 18675
rect 31440 18640 31475 18675
rect 31485 18640 31520 18675
rect 31530 18640 31565 18675
rect 31575 18640 31610 18675
rect 31620 18640 31655 18675
rect 31665 18640 31700 18675
rect 31710 18640 31745 18675
rect 31755 18640 31790 18675
rect 31800 18640 31835 18675
rect 31845 18640 31880 18675
rect 31890 18640 31925 18675
rect 31935 18640 31970 18675
rect 31980 18640 32015 18675
rect 32025 18640 32060 18675
rect 32070 18640 32105 18675
rect 32115 18640 32150 18675
rect 32160 18640 32195 18675
rect 32205 18640 32240 18675
rect 32250 18640 32285 18675
rect 32295 18640 32330 18675
rect 32340 18640 32375 18675
rect 32385 18640 32420 18675
rect 32430 18640 32465 18675
rect 32475 18640 32510 18675
rect 32520 18640 32555 18675
rect 32565 18640 32600 18675
rect 32610 18640 32645 18675
rect 32655 18640 32690 18675
rect 32700 18640 32735 18675
rect 32745 18640 32780 18675
rect 32790 18640 32825 18675
rect 32835 18640 32870 18675
rect 31305 18595 31340 18630
rect 31350 18595 31385 18630
rect 31395 18595 31430 18630
rect 31440 18595 31475 18630
rect 31485 18595 31520 18630
rect 31530 18595 31565 18630
rect 31575 18595 31610 18630
rect 31620 18595 31655 18630
rect 31665 18595 31700 18630
rect 31710 18595 31745 18630
rect 31755 18595 31790 18630
rect 31800 18595 31835 18630
rect 31845 18595 31880 18630
rect 31890 18595 31925 18630
rect 31935 18595 31970 18630
rect 31980 18595 32015 18630
rect 32025 18595 32060 18630
rect 32070 18595 32105 18630
rect 32115 18595 32150 18630
rect 32160 18595 32195 18630
rect 32205 18595 32240 18630
rect 32250 18595 32285 18630
rect 32295 18595 32330 18630
rect 32340 18595 32375 18630
rect 32385 18595 32420 18630
rect 32430 18595 32465 18630
rect 32475 18595 32510 18630
rect 32520 18595 32555 18630
rect 32565 18595 32600 18630
rect 32610 18595 32645 18630
rect 32655 18595 32690 18630
rect 32700 18595 32735 18630
rect 32745 18595 32780 18630
rect 32790 18595 32825 18630
rect 32835 18595 32870 18630
rect 31305 18550 31340 18585
rect 31350 18550 31385 18585
rect 31395 18550 31430 18585
rect 31440 18550 31475 18585
rect 31485 18550 31520 18585
rect 31530 18550 31565 18585
rect 31575 18550 31610 18585
rect 31620 18550 31655 18585
rect 31665 18550 31700 18585
rect 31710 18550 31745 18585
rect 31755 18550 31790 18585
rect 31800 18550 31835 18585
rect 31845 18550 31880 18585
rect 31890 18550 31925 18585
rect 31935 18550 31970 18585
rect 31980 18550 32015 18585
rect 32025 18550 32060 18585
rect 32070 18550 32105 18585
rect 32115 18550 32150 18585
rect 32160 18550 32195 18585
rect 32205 18550 32240 18585
rect 32250 18550 32285 18585
rect 32295 18550 32330 18585
rect 32340 18550 32375 18585
rect 32385 18550 32420 18585
rect 32430 18550 32465 18585
rect 32475 18550 32510 18585
rect 32520 18550 32555 18585
rect 32565 18550 32600 18585
rect 32610 18550 32645 18585
rect 32655 18550 32690 18585
rect 32700 18550 32735 18585
rect 32745 18550 32780 18585
rect 32790 18550 32825 18585
rect 32835 18550 32870 18585
rect 31305 18505 31340 18540
rect 31350 18505 31385 18540
rect 31395 18505 31430 18540
rect 31440 18505 31475 18540
rect 31485 18505 31520 18540
rect 31530 18505 31565 18540
rect 31575 18505 31610 18540
rect 31620 18505 31655 18540
rect 31665 18505 31700 18540
rect 31710 18505 31745 18540
rect 31755 18505 31790 18540
rect 31800 18505 31835 18540
rect 31845 18505 31880 18540
rect 31890 18505 31925 18540
rect 31935 18505 31970 18540
rect 31980 18505 32015 18540
rect 32025 18505 32060 18540
rect 32070 18505 32105 18540
rect 32115 18505 32150 18540
rect 32160 18505 32195 18540
rect 32205 18505 32240 18540
rect 32250 18505 32285 18540
rect 32295 18505 32330 18540
rect 32340 18505 32375 18540
rect 32385 18505 32420 18540
rect 32430 18505 32465 18540
rect 32475 18505 32510 18540
rect 32520 18505 32555 18540
rect 32565 18505 32600 18540
rect 32610 18505 32645 18540
rect 32655 18505 32690 18540
rect 32700 18505 32735 18540
rect 32745 18505 32780 18540
rect 32790 18505 32825 18540
rect 32835 18505 32870 18540
rect 31305 18460 31340 18495
rect 31350 18460 31385 18495
rect 31395 18460 31430 18495
rect 31440 18460 31475 18495
rect 31485 18460 31520 18495
rect 31530 18460 31565 18495
rect 31575 18460 31610 18495
rect 31620 18460 31655 18495
rect 31665 18460 31700 18495
rect 31710 18460 31745 18495
rect 31755 18460 31790 18495
rect 31800 18460 31835 18495
rect 31845 18460 31880 18495
rect 31890 18460 31925 18495
rect 31935 18460 31970 18495
rect 31980 18460 32015 18495
rect 32025 18460 32060 18495
rect 32070 18460 32105 18495
rect 32115 18460 32150 18495
rect 32160 18460 32195 18495
rect 32205 18460 32240 18495
rect 32250 18460 32285 18495
rect 32295 18460 32330 18495
rect 32340 18460 32375 18495
rect 32385 18460 32420 18495
rect 32430 18460 32465 18495
rect 32475 18460 32510 18495
rect 32520 18460 32555 18495
rect 32565 18460 32600 18495
rect 32610 18460 32645 18495
rect 32655 18460 32690 18495
rect 32700 18460 32735 18495
rect 32745 18460 32780 18495
rect 32790 18460 32825 18495
rect 32835 18460 32870 18495
rect 31305 18415 31340 18450
rect 31350 18415 31385 18450
rect 31395 18415 31430 18450
rect 31440 18415 31475 18450
rect 31485 18415 31520 18450
rect 31530 18415 31565 18450
rect 31575 18415 31610 18450
rect 31620 18415 31655 18450
rect 31665 18415 31700 18450
rect 31710 18415 31745 18450
rect 31755 18415 31790 18450
rect 31800 18415 31835 18450
rect 31845 18415 31880 18450
rect 31890 18415 31925 18450
rect 31935 18415 31970 18450
rect 31980 18415 32015 18450
rect 32025 18415 32060 18450
rect 32070 18415 32105 18450
rect 32115 18415 32150 18450
rect 32160 18415 32195 18450
rect 32205 18415 32240 18450
rect 32250 18415 32285 18450
rect 32295 18415 32330 18450
rect 32340 18415 32375 18450
rect 32385 18415 32420 18450
rect 32430 18415 32465 18450
rect 32475 18415 32510 18450
rect 32520 18415 32555 18450
rect 32565 18415 32600 18450
rect 32610 18415 32645 18450
rect 32655 18415 32690 18450
rect 32700 18415 32735 18450
rect 32745 18415 32780 18450
rect 32790 18415 32825 18450
rect 32835 18415 32870 18450
rect 31305 18370 31340 18405
rect 31350 18370 31385 18405
rect 31395 18370 31430 18405
rect 31440 18370 31475 18405
rect 31485 18370 31520 18405
rect 31530 18370 31565 18405
rect 31575 18370 31610 18405
rect 31620 18370 31655 18405
rect 31665 18370 31700 18405
rect 31710 18370 31745 18405
rect 31755 18370 31790 18405
rect 31800 18370 31835 18405
rect 31845 18370 31880 18405
rect 31890 18370 31925 18405
rect 31935 18370 31970 18405
rect 31980 18370 32015 18405
rect 32025 18370 32060 18405
rect 32070 18370 32105 18405
rect 32115 18370 32150 18405
rect 32160 18370 32195 18405
rect 32205 18370 32240 18405
rect 32250 18370 32285 18405
rect 32295 18370 32330 18405
rect 32340 18370 32375 18405
rect 32385 18370 32420 18405
rect 32430 18370 32465 18405
rect 32475 18370 32510 18405
rect 32520 18370 32555 18405
rect 32565 18370 32600 18405
rect 32610 18370 32645 18405
rect 32655 18370 32690 18405
rect 32700 18370 32735 18405
rect 32745 18370 32780 18405
rect 32790 18370 32825 18405
rect 32835 18370 32870 18405
rect 31305 18325 31340 18360
rect 31350 18325 31385 18360
rect 31395 18325 31430 18360
rect 31440 18325 31475 18360
rect 31485 18325 31520 18360
rect 31530 18325 31565 18360
rect 31575 18325 31610 18360
rect 31620 18325 31655 18360
rect 31665 18325 31700 18360
rect 31710 18325 31745 18360
rect 31755 18325 31790 18360
rect 31800 18325 31835 18360
rect 31845 18325 31880 18360
rect 31890 18325 31925 18360
rect 31935 18325 31970 18360
rect 31980 18325 32015 18360
rect 32025 18325 32060 18360
rect 32070 18325 32105 18360
rect 32115 18325 32150 18360
rect 32160 18325 32195 18360
rect 32205 18325 32240 18360
rect 32250 18325 32285 18360
rect 32295 18325 32330 18360
rect 32340 18325 32375 18360
rect 32385 18325 32420 18360
rect 32430 18325 32465 18360
rect 32475 18325 32510 18360
rect 32520 18325 32555 18360
rect 32565 18325 32600 18360
rect 32610 18325 32645 18360
rect 32655 18325 32690 18360
rect 32700 18325 32735 18360
rect 32745 18325 32780 18360
rect 32790 18325 32825 18360
rect 32835 18325 32870 18360
rect 31305 18280 31340 18315
rect 31350 18280 31385 18315
rect 31395 18280 31430 18315
rect 31440 18280 31475 18315
rect 31485 18280 31520 18315
rect 31530 18280 31565 18315
rect 31575 18280 31610 18315
rect 31620 18280 31655 18315
rect 31665 18280 31700 18315
rect 31710 18280 31745 18315
rect 31755 18280 31790 18315
rect 31800 18280 31835 18315
rect 31845 18280 31880 18315
rect 31890 18280 31925 18315
rect 31935 18280 31970 18315
rect 31980 18280 32015 18315
rect 32025 18280 32060 18315
rect 32070 18280 32105 18315
rect 32115 18280 32150 18315
rect 32160 18280 32195 18315
rect 32205 18280 32240 18315
rect 32250 18280 32285 18315
rect 32295 18280 32330 18315
rect 32340 18280 32375 18315
rect 32385 18280 32420 18315
rect 32430 18280 32465 18315
rect 32475 18280 32510 18315
rect 32520 18280 32555 18315
rect 32565 18280 32600 18315
rect 32610 18280 32645 18315
rect 32655 18280 32690 18315
rect 32700 18280 32735 18315
rect 32745 18280 32780 18315
rect 32790 18280 32825 18315
rect 32835 18280 32870 18315
rect 31305 18235 31340 18270
rect 31350 18235 31385 18270
rect 31395 18235 31430 18270
rect 31440 18235 31475 18270
rect 31485 18235 31520 18270
rect 31530 18235 31565 18270
rect 31575 18235 31610 18270
rect 31620 18235 31655 18270
rect 31665 18235 31700 18270
rect 31710 18235 31745 18270
rect 31755 18235 31790 18270
rect 31800 18235 31835 18270
rect 31845 18235 31880 18270
rect 31890 18235 31925 18270
rect 31935 18235 31970 18270
rect 31980 18235 32015 18270
rect 32025 18235 32060 18270
rect 32070 18235 32105 18270
rect 32115 18235 32150 18270
rect 32160 18235 32195 18270
rect 32205 18235 32240 18270
rect 32250 18235 32285 18270
rect 32295 18235 32330 18270
rect 32340 18235 32375 18270
rect 32385 18235 32420 18270
rect 32430 18235 32465 18270
rect 32475 18235 32510 18270
rect 32520 18235 32555 18270
rect 32565 18235 32600 18270
rect 32610 18235 32645 18270
rect 32655 18235 32690 18270
rect 32700 18235 32735 18270
rect 32745 18235 32780 18270
rect 32790 18235 32825 18270
rect 32835 18235 32870 18270
rect 31305 18190 31340 18225
rect 31350 18190 31385 18225
rect 31395 18190 31430 18225
rect 31440 18190 31475 18225
rect 31485 18190 31520 18225
rect 31530 18190 31565 18225
rect 31575 18190 31610 18225
rect 31620 18190 31655 18225
rect 31665 18190 31700 18225
rect 31710 18190 31745 18225
rect 31755 18190 31790 18225
rect 31800 18190 31835 18225
rect 31845 18190 31880 18225
rect 31890 18190 31925 18225
rect 31935 18190 31970 18225
rect 31980 18190 32015 18225
rect 32025 18190 32060 18225
rect 32070 18190 32105 18225
rect 32115 18190 32150 18225
rect 32160 18190 32195 18225
rect 32205 18190 32240 18225
rect 32250 18190 32285 18225
rect 32295 18190 32330 18225
rect 32340 18190 32375 18225
rect 32385 18190 32420 18225
rect 32430 18190 32465 18225
rect 32475 18190 32510 18225
rect 32520 18190 32555 18225
rect 32565 18190 32600 18225
rect 32610 18190 32645 18225
rect 32655 18190 32690 18225
rect 32700 18190 32735 18225
rect 32745 18190 32780 18225
rect 32790 18190 32825 18225
rect 32835 18190 32870 18225
rect 31305 18145 31340 18180
rect 31350 18145 31385 18180
rect 31395 18145 31430 18180
rect 31440 18145 31475 18180
rect 31485 18145 31520 18180
rect 31530 18145 31565 18180
rect 31575 18145 31610 18180
rect 31620 18145 31655 18180
rect 31665 18145 31700 18180
rect 31710 18145 31745 18180
rect 31755 18145 31790 18180
rect 31800 18145 31835 18180
rect 31845 18145 31880 18180
rect 31890 18145 31925 18180
rect 31935 18145 31970 18180
rect 31980 18145 32015 18180
rect 32025 18145 32060 18180
rect 32070 18145 32105 18180
rect 32115 18145 32150 18180
rect 32160 18145 32195 18180
rect 32205 18145 32240 18180
rect 32250 18145 32285 18180
rect 32295 18145 32330 18180
rect 32340 18145 32375 18180
rect 32385 18145 32420 18180
rect 32430 18145 32465 18180
rect 32475 18145 32510 18180
rect 32520 18145 32555 18180
rect 32565 18145 32600 18180
rect 32610 18145 32645 18180
rect 32655 18145 32690 18180
rect 32700 18145 32735 18180
rect 32745 18145 32780 18180
rect 32790 18145 32825 18180
rect 32835 18145 32870 18180
rect 31305 18100 31340 18135
rect 31350 18100 31385 18135
rect 31395 18100 31430 18135
rect 31440 18100 31475 18135
rect 31485 18100 31520 18135
rect 31530 18100 31565 18135
rect 31575 18100 31610 18135
rect 31620 18100 31655 18135
rect 31665 18100 31700 18135
rect 31710 18100 31745 18135
rect 31755 18100 31790 18135
rect 31800 18100 31835 18135
rect 31845 18100 31880 18135
rect 31890 18100 31925 18135
rect 31935 18100 31970 18135
rect 31980 18100 32015 18135
rect 32025 18100 32060 18135
rect 32070 18100 32105 18135
rect 32115 18100 32150 18135
rect 32160 18100 32195 18135
rect 32205 18100 32240 18135
rect 32250 18100 32285 18135
rect 32295 18100 32330 18135
rect 32340 18100 32375 18135
rect 32385 18100 32420 18135
rect 32430 18100 32465 18135
rect 32475 18100 32510 18135
rect 32520 18100 32555 18135
rect 32565 18100 32600 18135
rect 32610 18100 32645 18135
rect 32655 18100 32690 18135
rect 32700 18100 32735 18135
rect 32745 18100 32780 18135
rect 32790 18100 32825 18135
rect 32835 18100 32870 18135
rect 31305 18055 31340 18090
rect 31350 18055 31385 18090
rect 31395 18055 31430 18090
rect 31440 18055 31475 18090
rect 31485 18055 31520 18090
rect 31530 18055 31565 18090
rect 31575 18055 31610 18090
rect 31620 18055 31655 18090
rect 31665 18055 31700 18090
rect 31710 18055 31745 18090
rect 31755 18055 31790 18090
rect 31800 18055 31835 18090
rect 31845 18055 31880 18090
rect 31890 18055 31925 18090
rect 31935 18055 31970 18090
rect 31980 18055 32015 18090
rect 32025 18055 32060 18090
rect 32070 18055 32105 18090
rect 32115 18055 32150 18090
rect 32160 18055 32195 18090
rect 32205 18055 32240 18090
rect 32250 18055 32285 18090
rect 32295 18055 32330 18090
rect 32340 18055 32375 18090
rect 32385 18055 32420 18090
rect 32430 18055 32465 18090
rect 32475 18055 32510 18090
rect 32520 18055 32555 18090
rect 32565 18055 32600 18090
rect 32610 18055 32645 18090
rect 32655 18055 32690 18090
rect 32700 18055 32735 18090
rect 32745 18055 32780 18090
rect 32790 18055 32825 18090
rect 32835 18055 32870 18090
rect 31305 18010 31340 18045
rect 31350 18010 31385 18045
rect 31395 18010 31430 18045
rect 31440 18010 31475 18045
rect 31485 18010 31520 18045
rect 31530 18010 31565 18045
rect 31575 18010 31610 18045
rect 31620 18010 31655 18045
rect 31665 18010 31700 18045
rect 31710 18010 31745 18045
rect 31755 18010 31790 18045
rect 31800 18010 31835 18045
rect 31845 18010 31880 18045
rect 31890 18010 31925 18045
rect 31935 18010 31970 18045
rect 31980 18010 32015 18045
rect 32025 18010 32060 18045
rect 32070 18010 32105 18045
rect 32115 18010 32150 18045
rect 32160 18010 32195 18045
rect 32205 18010 32240 18045
rect 32250 18010 32285 18045
rect 32295 18010 32330 18045
rect 32340 18010 32375 18045
rect 32385 18010 32420 18045
rect 32430 18010 32465 18045
rect 32475 18010 32510 18045
rect 32520 18010 32555 18045
rect 32565 18010 32600 18045
rect 32610 18010 32645 18045
rect 32655 18010 32690 18045
rect 32700 18010 32735 18045
rect 32745 18010 32780 18045
rect 32790 18010 32825 18045
rect 32835 18010 32870 18045
rect 31305 17965 31340 18000
rect 31350 17965 31385 18000
rect 31395 17965 31430 18000
rect 31440 17965 31475 18000
rect 31485 17965 31520 18000
rect 31530 17965 31565 18000
rect 31575 17965 31610 18000
rect 31620 17965 31655 18000
rect 31665 17965 31700 18000
rect 31710 17965 31745 18000
rect 31755 17965 31790 18000
rect 31800 17965 31835 18000
rect 31845 17965 31880 18000
rect 31890 17965 31925 18000
rect 31935 17965 31970 18000
rect 31980 17965 32015 18000
rect 32025 17965 32060 18000
rect 32070 17965 32105 18000
rect 32115 17965 32150 18000
rect 32160 17965 32195 18000
rect 32205 17965 32240 18000
rect 32250 17965 32285 18000
rect 32295 17965 32330 18000
rect 32340 17965 32375 18000
rect 32385 17965 32420 18000
rect 32430 17965 32465 18000
rect 32475 17965 32510 18000
rect 32520 17965 32555 18000
rect 32565 17965 32600 18000
rect 32610 17965 32645 18000
rect 32655 17965 32690 18000
rect 32700 17965 32735 18000
rect 32745 17965 32780 18000
rect 32790 17965 32825 18000
rect 32835 17965 32870 18000
rect 31305 17920 31340 17955
rect 31350 17920 31385 17955
rect 31395 17920 31430 17955
rect 31440 17920 31475 17955
rect 31485 17920 31520 17955
rect 31530 17920 31565 17955
rect 31575 17920 31610 17955
rect 31620 17920 31655 17955
rect 31665 17920 31700 17955
rect 31710 17920 31745 17955
rect 31755 17920 31790 17955
rect 31800 17920 31835 17955
rect 31845 17920 31880 17955
rect 31890 17920 31925 17955
rect 31935 17920 31970 17955
rect 31980 17920 32015 17955
rect 32025 17920 32060 17955
rect 32070 17920 32105 17955
rect 32115 17920 32150 17955
rect 32160 17920 32195 17955
rect 32205 17920 32240 17955
rect 32250 17920 32285 17955
rect 32295 17920 32330 17955
rect 32340 17920 32375 17955
rect 32385 17920 32420 17955
rect 32430 17920 32465 17955
rect 32475 17920 32510 17955
rect 32520 17920 32555 17955
rect 32565 17920 32600 17955
rect 32610 17920 32645 17955
rect 32655 17920 32690 17955
rect 32700 17920 32735 17955
rect 32745 17920 32780 17955
rect 32790 17920 32825 17955
rect 32835 17920 32870 17955
rect 31305 17875 31340 17910
rect 31350 17875 31385 17910
rect 31395 17875 31430 17910
rect 31440 17875 31475 17910
rect 31485 17875 31520 17910
rect 31530 17875 31565 17910
rect 31575 17875 31610 17910
rect 31620 17875 31655 17910
rect 31665 17875 31700 17910
rect 31710 17875 31745 17910
rect 31755 17875 31790 17910
rect 31800 17875 31835 17910
rect 31845 17875 31880 17910
rect 31890 17875 31925 17910
rect 31935 17875 31970 17910
rect 31980 17875 32015 17910
rect 32025 17875 32060 17910
rect 32070 17875 32105 17910
rect 32115 17875 32150 17910
rect 32160 17875 32195 17910
rect 32205 17875 32240 17910
rect 32250 17875 32285 17910
rect 32295 17875 32330 17910
rect 32340 17875 32375 17910
rect 32385 17875 32420 17910
rect 32430 17875 32465 17910
rect 32475 17875 32510 17910
rect 32520 17875 32555 17910
rect 32565 17875 32600 17910
rect 32610 17875 32645 17910
rect 32655 17875 32690 17910
rect 32700 17875 32735 17910
rect 32745 17875 32780 17910
rect 32790 17875 32825 17910
rect 32835 17875 32870 17910
rect 31305 17830 31340 17865
rect 31350 17830 31385 17865
rect 31395 17830 31430 17865
rect 31440 17830 31475 17865
rect 31485 17830 31520 17865
rect 31530 17830 31565 17865
rect 31575 17830 31610 17865
rect 31620 17830 31655 17865
rect 31665 17830 31700 17865
rect 31710 17830 31745 17865
rect 31755 17830 31790 17865
rect 31800 17830 31835 17865
rect 31845 17830 31880 17865
rect 31890 17830 31925 17865
rect 31935 17830 31970 17865
rect 31980 17830 32015 17865
rect 32025 17830 32060 17865
rect 32070 17830 32105 17865
rect 32115 17830 32150 17865
rect 32160 17830 32195 17865
rect 32205 17830 32240 17865
rect 32250 17830 32285 17865
rect 32295 17830 32330 17865
rect 32340 17830 32375 17865
rect 32385 17830 32420 17865
rect 32430 17830 32465 17865
rect 32475 17830 32510 17865
rect 32520 17830 32555 17865
rect 32565 17830 32600 17865
rect 32610 17830 32645 17865
rect 32655 17830 32690 17865
rect 32700 17830 32735 17865
rect 32745 17830 32780 17865
rect 32790 17830 32825 17865
rect 32835 17830 32870 17865
rect 31305 17785 31340 17820
rect 31350 17785 31385 17820
rect 31395 17785 31430 17820
rect 31440 17785 31475 17820
rect 31485 17785 31520 17820
rect 31530 17785 31565 17820
rect 31575 17785 31610 17820
rect 31620 17785 31655 17820
rect 31665 17785 31700 17820
rect 31710 17785 31745 17820
rect 31755 17785 31790 17820
rect 31800 17785 31835 17820
rect 31845 17785 31880 17820
rect 31890 17785 31925 17820
rect 31935 17785 31970 17820
rect 31980 17785 32015 17820
rect 32025 17785 32060 17820
rect 32070 17785 32105 17820
rect 32115 17785 32150 17820
rect 32160 17785 32195 17820
rect 32205 17785 32240 17820
rect 32250 17785 32285 17820
rect 32295 17785 32330 17820
rect 32340 17785 32375 17820
rect 32385 17785 32420 17820
rect 32430 17785 32465 17820
rect 32475 17785 32510 17820
rect 32520 17785 32555 17820
rect 32565 17785 32600 17820
rect 32610 17785 32645 17820
rect 32655 17785 32690 17820
rect 32700 17785 32735 17820
rect 32745 17785 32780 17820
rect 32790 17785 32825 17820
rect 32835 17785 32870 17820
rect 31305 17740 31340 17775
rect 31350 17740 31385 17775
rect 31395 17740 31430 17775
rect 31440 17740 31475 17775
rect 31485 17740 31520 17775
rect 31530 17740 31565 17775
rect 31575 17740 31610 17775
rect 31620 17740 31655 17775
rect 31665 17740 31700 17775
rect 31710 17740 31745 17775
rect 31755 17740 31790 17775
rect 31800 17740 31835 17775
rect 31845 17740 31880 17775
rect 31890 17740 31925 17775
rect 31935 17740 31970 17775
rect 31980 17740 32015 17775
rect 32025 17740 32060 17775
rect 32070 17740 32105 17775
rect 32115 17740 32150 17775
rect 32160 17740 32195 17775
rect 32205 17740 32240 17775
rect 32250 17740 32285 17775
rect 32295 17740 32330 17775
rect 32340 17740 32375 17775
rect 32385 17740 32420 17775
rect 32430 17740 32465 17775
rect 32475 17740 32510 17775
rect 32520 17740 32555 17775
rect 32565 17740 32600 17775
rect 32610 17740 32645 17775
rect 32655 17740 32690 17775
rect 32700 17740 32735 17775
rect 32745 17740 32780 17775
rect 32790 17740 32825 17775
rect 32835 17740 32870 17775
rect 31305 10495 31340 10530
rect 31350 10495 31385 10530
rect 31395 10495 31430 10530
rect 31440 10495 31475 10530
rect 31485 10495 31520 10530
rect 31530 10495 31565 10530
rect 31575 10495 31610 10530
rect 31620 10495 31655 10530
rect 31665 10495 31700 10530
rect 31710 10495 31745 10530
rect 31755 10495 31790 10530
rect 31800 10495 31835 10530
rect 31845 10495 31880 10530
rect 31890 10495 31925 10530
rect 31935 10495 31970 10530
rect 31980 10495 32015 10530
rect 32025 10495 32060 10530
rect 32070 10495 32105 10530
rect 32115 10495 32150 10530
rect 32160 10495 32195 10530
rect 32205 10495 32240 10530
rect 32250 10495 32285 10530
rect 32295 10495 32330 10530
rect 32340 10495 32375 10530
rect 32385 10495 32420 10530
rect 32430 10495 32465 10530
rect 32475 10495 32510 10530
rect 32520 10495 32555 10530
rect 32565 10495 32600 10530
rect 32610 10495 32645 10530
rect 32655 10495 32690 10530
rect 32700 10495 32735 10530
rect 32745 10495 32780 10530
rect 32790 10495 32825 10530
rect 32835 10495 32870 10530
rect 31305 10450 31340 10485
rect 31350 10450 31385 10485
rect 31395 10450 31430 10485
rect 31440 10450 31475 10485
rect 31485 10450 31520 10485
rect 31530 10450 31565 10485
rect 31575 10450 31610 10485
rect 31620 10450 31655 10485
rect 31665 10450 31700 10485
rect 31710 10450 31745 10485
rect 31755 10450 31790 10485
rect 31800 10450 31835 10485
rect 31845 10450 31880 10485
rect 31890 10450 31925 10485
rect 31935 10450 31970 10485
rect 31980 10450 32015 10485
rect 32025 10450 32060 10485
rect 32070 10450 32105 10485
rect 32115 10450 32150 10485
rect 32160 10450 32195 10485
rect 32205 10450 32240 10485
rect 32250 10450 32285 10485
rect 32295 10450 32330 10485
rect 32340 10450 32375 10485
rect 32385 10450 32420 10485
rect 32430 10450 32465 10485
rect 32475 10450 32510 10485
rect 32520 10450 32555 10485
rect 32565 10450 32600 10485
rect 32610 10450 32645 10485
rect 32655 10450 32690 10485
rect 32700 10450 32735 10485
rect 32745 10450 32780 10485
rect 32790 10450 32825 10485
rect 32835 10450 32870 10485
rect 31305 10405 31340 10440
rect 31350 10405 31385 10440
rect 31395 10405 31430 10440
rect 31440 10405 31475 10440
rect 31485 10405 31520 10440
rect 31530 10405 31565 10440
rect 31575 10405 31610 10440
rect 31620 10405 31655 10440
rect 31665 10405 31700 10440
rect 31710 10405 31745 10440
rect 31755 10405 31790 10440
rect 31800 10405 31835 10440
rect 31845 10405 31880 10440
rect 31890 10405 31925 10440
rect 31935 10405 31970 10440
rect 31980 10405 32015 10440
rect 32025 10405 32060 10440
rect 32070 10405 32105 10440
rect 32115 10405 32150 10440
rect 32160 10405 32195 10440
rect 32205 10405 32240 10440
rect 32250 10405 32285 10440
rect 32295 10405 32330 10440
rect 32340 10405 32375 10440
rect 32385 10405 32420 10440
rect 32430 10405 32465 10440
rect 32475 10405 32510 10440
rect 32520 10405 32555 10440
rect 32565 10405 32600 10440
rect 32610 10405 32645 10440
rect 32655 10405 32690 10440
rect 32700 10405 32735 10440
rect 32745 10405 32780 10440
rect 32790 10405 32825 10440
rect 32835 10405 32870 10440
rect 31305 10360 31340 10395
rect 31350 10360 31385 10395
rect 31395 10360 31430 10395
rect 31440 10360 31475 10395
rect 31485 10360 31520 10395
rect 31530 10360 31565 10395
rect 31575 10360 31610 10395
rect 31620 10360 31655 10395
rect 31665 10360 31700 10395
rect 31710 10360 31745 10395
rect 31755 10360 31790 10395
rect 31800 10360 31835 10395
rect 31845 10360 31880 10395
rect 31890 10360 31925 10395
rect 31935 10360 31970 10395
rect 31980 10360 32015 10395
rect 32025 10360 32060 10395
rect 32070 10360 32105 10395
rect 32115 10360 32150 10395
rect 32160 10360 32195 10395
rect 32205 10360 32240 10395
rect 32250 10360 32285 10395
rect 32295 10360 32330 10395
rect 32340 10360 32375 10395
rect 32385 10360 32420 10395
rect 32430 10360 32465 10395
rect 32475 10360 32510 10395
rect 32520 10360 32555 10395
rect 32565 10360 32600 10395
rect 32610 10360 32645 10395
rect 32655 10360 32690 10395
rect 32700 10360 32735 10395
rect 32745 10360 32780 10395
rect 32790 10360 32825 10395
rect 32835 10360 32870 10395
rect 31305 10315 31340 10350
rect 31350 10315 31385 10350
rect 31395 10315 31430 10350
rect 31440 10315 31475 10350
rect 31485 10315 31520 10350
rect 31530 10315 31565 10350
rect 31575 10315 31610 10350
rect 31620 10315 31655 10350
rect 31665 10315 31700 10350
rect 31710 10315 31745 10350
rect 31755 10315 31790 10350
rect 31800 10315 31835 10350
rect 31845 10315 31880 10350
rect 31890 10315 31925 10350
rect 31935 10315 31970 10350
rect 31980 10315 32015 10350
rect 32025 10315 32060 10350
rect 32070 10315 32105 10350
rect 32115 10315 32150 10350
rect 32160 10315 32195 10350
rect 32205 10315 32240 10350
rect 32250 10315 32285 10350
rect 32295 10315 32330 10350
rect 32340 10315 32375 10350
rect 32385 10315 32420 10350
rect 32430 10315 32465 10350
rect 32475 10315 32510 10350
rect 32520 10315 32555 10350
rect 32565 10315 32600 10350
rect 32610 10315 32645 10350
rect 32655 10315 32690 10350
rect 32700 10315 32735 10350
rect 32745 10315 32780 10350
rect 32790 10315 32825 10350
rect 32835 10315 32870 10350
rect 31305 10270 31340 10305
rect 31350 10270 31385 10305
rect 31395 10270 31430 10305
rect 31440 10270 31475 10305
rect 31485 10270 31520 10305
rect 31530 10270 31565 10305
rect 31575 10270 31610 10305
rect 31620 10270 31655 10305
rect 31665 10270 31700 10305
rect 31710 10270 31745 10305
rect 31755 10270 31790 10305
rect 31800 10270 31835 10305
rect 31845 10270 31880 10305
rect 31890 10270 31925 10305
rect 31935 10270 31970 10305
rect 31980 10270 32015 10305
rect 32025 10270 32060 10305
rect 32070 10270 32105 10305
rect 32115 10270 32150 10305
rect 32160 10270 32195 10305
rect 32205 10270 32240 10305
rect 32250 10270 32285 10305
rect 32295 10270 32330 10305
rect 32340 10270 32375 10305
rect 32385 10270 32420 10305
rect 32430 10270 32465 10305
rect 32475 10270 32510 10305
rect 32520 10270 32555 10305
rect 32565 10270 32600 10305
rect 32610 10270 32645 10305
rect 32655 10270 32690 10305
rect 32700 10270 32735 10305
rect 32745 10270 32780 10305
rect 32790 10270 32825 10305
rect 32835 10270 32870 10305
rect 31305 10225 31340 10260
rect 31350 10225 31385 10260
rect 31395 10225 31430 10260
rect 31440 10225 31475 10260
rect 31485 10225 31520 10260
rect 31530 10225 31565 10260
rect 31575 10225 31610 10260
rect 31620 10225 31655 10260
rect 31665 10225 31700 10260
rect 31710 10225 31745 10260
rect 31755 10225 31790 10260
rect 31800 10225 31835 10260
rect 31845 10225 31880 10260
rect 31890 10225 31925 10260
rect 31935 10225 31970 10260
rect 31980 10225 32015 10260
rect 32025 10225 32060 10260
rect 32070 10225 32105 10260
rect 32115 10225 32150 10260
rect 32160 10225 32195 10260
rect 32205 10225 32240 10260
rect 32250 10225 32285 10260
rect 32295 10225 32330 10260
rect 32340 10225 32375 10260
rect 32385 10225 32420 10260
rect 32430 10225 32465 10260
rect 32475 10225 32510 10260
rect 32520 10225 32555 10260
rect 32565 10225 32600 10260
rect 32610 10225 32645 10260
rect 32655 10225 32690 10260
rect 32700 10225 32735 10260
rect 32745 10225 32780 10260
rect 32790 10225 32825 10260
rect 32835 10225 32870 10260
rect 31305 10180 31340 10215
rect 31350 10180 31385 10215
rect 31395 10180 31430 10215
rect 31440 10180 31475 10215
rect 31485 10180 31520 10215
rect 31530 10180 31565 10215
rect 31575 10180 31610 10215
rect 31620 10180 31655 10215
rect 31665 10180 31700 10215
rect 31710 10180 31745 10215
rect 31755 10180 31790 10215
rect 31800 10180 31835 10215
rect 31845 10180 31880 10215
rect 31890 10180 31925 10215
rect 31935 10180 31970 10215
rect 31980 10180 32015 10215
rect 32025 10180 32060 10215
rect 32070 10180 32105 10215
rect 32115 10180 32150 10215
rect 32160 10180 32195 10215
rect 32205 10180 32240 10215
rect 32250 10180 32285 10215
rect 32295 10180 32330 10215
rect 32340 10180 32375 10215
rect 32385 10180 32420 10215
rect 32430 10180 32465 10215
rect 32475 10180 32510 10215
rect 32520 10180 32555 10215
rect 32565 10180 32600 10215
rect 32610 10180 32645 10215
rect 32655 10180 32690 10215
rect 32700 10180 32735 10215
rect 32745 10180 32780 10215
rect 32790 10180 32825 10215
rect 32835 10180 32870 10215
rect 31305 10135 31340 10170
rect 31350 10135 31385 10170
rect 31395 10135 31430 10170
rect 31440 10135 31475 10170
rect 31485 10135 31520 10170
rect 31530 10135 31565 10170
rect 31575 10135 31610 10170
rect 31620 10135 31655 10170
rect 31665 10135 31700 10170
rect 31710 10135 31745 10170
rect 31755 10135 31790 10170
rect 31800 10135 31835 10170
rect 31845 10135 31880 10170
rect 31890 10135 31925 10170
rect 31935 10135 31970 10170
rect 31980 10135 32015 10170
rect 32025 10135 32060 10170
rect 32070 10135 32105 10170
rect 32115 10135 32150 10170
rect 32160 10135 32195 10170
rect 32205 10135 32240 10170
rect 32250 10135 32285 10170
rect 32295 10135 32330 10170
rect 32340 10135 32375 10170
rect 32385 10135 32420 10170
rect 32430 10135 32465 10170
rect 32475 10135 32510 10170
rect 32520 10135 32555 10170
rect 32565 10135 32600 10170
rect 32610 10135 32645 10170
rect 32655 10135 32690 10170
rect 32700 10135 32735 10170
rect 32745 10135 32780 10170
rect 32790 10135 32825 10170
rect 32835 10135 32870 10170
rect 31305 10090 31340 10125
rect 31350 10090 31385 10125
rect 31395 10090 31430 10125
rect 31440 10090 31475 10125
rect 31485 10090 31520 10125
rect 31530 10090 31565 10125
rect 31575 10090 31610 10125
rect 31620 10090 31655 10125
rect 31665 10090 31700 10125
rect 31710 10090 31745 10125
rect 31755 10090 31790 10125
rect 31800 10090 31835 10125
rect 31845 10090 31880 10125
rect 31890 10090 31925 10125
rect 31935 10090 31970 10125
rect 31980 10090 32015 10125
rect 32025 10090 32060 10125
rect 32070 10090 32105 10125
rect 32115 10090 32150 10125
rect 32160 10090 32195 10125
rect 32205 10090 32240 10125
rect 32250 10090 32285 10125
rect 32295 10090 32330 10125
rect 32340 10090 32375 10125
rect 32385 10090 32420 10125
rect 32430 10090 32465 10125
rect 32475 10090 32510 10125
rect 32520 10090 32555 10125
rect 32565 10090 32600 10125
rect 32610 10090 32645 10125
rect 32655 10090 32690 10125
rect 32700 10090 32735 10125
rect 32745 10090 32780 10125
rect 32790 10090 32825 10125
rect 32835 10090 32870 10125
rect 31305 10045 31340 10080
rect 31350 10045 31385 10080
rect 31395 10045 31430 10080
rect 31440 10045 31475 10080
rect 31485 10045 31520 10080
rect 31530 10045 31565 10080
rect 31575 10045 31610 10080
rect 31620 10045 31655 10080
rect 31665 10045 31700 10080
rect 31710 10045 31745 10080
rect 31755 10045 31790 10080
rect 31800 10045 31835 10080
rect 31845 10045 31880 10080
rect 31890 10045 31925 10080
rect 31935 10045 31970 10080
rect 31980 10045 32015 10080
rect 32025 10045 32060 10080
rect 32070 10045 32105 10080
rect 32115 10045 32150 10080
rect 32160 10045 32195 10080
rect 32205 10045 32240 10080
rect 32250 10045 32285 10080
rect 32295 10045 32330 10080
rect 32340 10045 32375 10080
rect 32385 10045 32420 10080
rect 32430 10045 32465 10080
rect 32475 10045 32510 10080
rect 32520 10045 32555 10080
rect 32565 10045 32600 10080
rect 32610 10045 32645 10080
rect 32655 10045 32690 10080
rect 32700 10045 32735 10080
rect 32745 10045 32780 10080
rect 32790 10045 32825 10080
rect 32835 10045 32870 10080
rect 31305 10000 31340 10035
rect 31350 10000 31385 10035
rect 31395 10000 31430 10035
rect 31440 10000 31475 10035
rect 31485 10000 31520 10035
rect 31530 10000 31565 10035
rect 31575 10000 31610 10035
rect 31620 10000 31655 10035
rect 31665 10000 31700 10035
rect 31710 10000 31745 10035
rect 31755 10000 31790 10035
rect 31800 10000 31835 10035
rect 31845 10000 31880 10035
rect 31890 10000 31925 10035
rect 31935 10000 31970 10035
rect 31980 10000 32015 10035
rect 32025 10000 32060 10035
rect 32070 10000 32105 10035
rect 32115 10000 32150 10035
rect 32160 10000 32195 10035
rect 32205 10000 32240 10035
rect 32250 10000 32285 10035
rect 32295 10000 32330 10035
rect 32340 10000 32375 10035
rect 32385 10000 32420 10035
rect 32430 10000 32465 10035
rect 32475 10000 32510 10035
rect 32520 10000 32555 10035
rect 32565 10000 32600 10035
rect 32610 10000 32645 10035
rect 32655 10000 32690 10035
rect 32700 10000 32735 10035
rect 32745 10000 32780 10035
rect 32790 10000 32825 10035
rect 32835 10000 32870 10035
rect 31305 9955 31340 9990
rect 31350 9955 31385 9990
rect 31395 9955 31430 9990
rect 31440 9955 31475 9990
rect 31485 9955 31520 9990
rect 31530 9955 31565 9990
rect 31575 9955 31610 9990
rect 31620 9955 31655 9990
rect 31665 9955 31700 9990
rect 31710 9955 31745 9990
rect 31755 9955 31790 9990
rect 31800 9955 31835 9990
rect 31845 9955 31880 9990
rect 31890 9955 31925 9990
rect 31935 9955 31970 9990
rect 31980 9955 32015 9990
rect 32025 9955 32060 9990
rect 32070 9955 32105 9990
rect 32115 9955 32150 9990
rect 32160 9955 32195 9990
rect 32205 9955 32240 9990
rect 32250 9955 32285 9990
rect 32295 9955 32330 9990
rect 32340 9955 32375 9990
rect 32385 9955 32420 9990
rect 32430 9955 32465 9990
rect 32475 9955 32510 9990
rect 32520 9955 32555 9990
rect 32565 9955 32600 9990
rect 32610 9955 32645 9990
rect 32655 9955 32690 9990
rect 32700 9955 32735 9990
rect 32745 9955 32780 9990
rect 32790 9955 32825 9990
rect 32835 9955 32870 9990
rect 31305 9910 31340 9945
rect 31350 9910 31385 9945
rect 31395 9910 31430 9945
rect 31440 9910 31475 9945
rect 31485 9910 31520 9945
rect 31530 9910 31565 9945
rect 31575 9910 31610 9945
rect 31620 9910 31655 9945
rect 31665 9910 31700 9945
rect 31710 9910 31745 9945
rect 31755 9910 31790 9945
rect 31800 9910 31835 9945
rect 31845 9910 31880 9945
rect 31890 9910 31925 9945
rect 31935 9910 31970 9945
rect 31980 9910 32015 9945
rect 32025 9910 32060 9945
rect 32070 9910 32105 9945
rect 32115 9910 32150 9945
rect 32160 9910 32195 9945
rect 32205 9910 32240 9945
rect 32250 9910 32285 9945
rect 32295 9910 32330 9945
rect 32340 9910 32375 9945
rect 32385 9910 32420 9945
rect 32430 9910 32465 9945
rect 32475 9910 32510 9945
rect 32520 9910 32555 9945
rect 32565 9910 32600 9945
rect 32610 9910 32645 9945
rect 32655 9910 32690 9945
rect 32700 9910 32735 9945
rect 32745 9910 32780 9945
rect 32790 9910 32825 9945
rect 32835 9910 32870 9945
rect 31305 9865 31340 9900
rect 31350 9865 31385 9900
rect 31395 9865 31430 9900
rect 31440 9865 31475 9900
rect 31485 9865 31520 9900
rect 31530 9865 31565 9900
rect 31575 9865 31610 9900
rect 31620 9865 31655 9900
rect 31665 9865 31700 9900
rect 31710 9865 31745 9900
rect 31755 9865 31790 9900
rect 31800 9865 31835 9900
rect 31845 9865 31880 9900
rect 31890 9865 31925 9900
rect 31935 9865 31970 9900
rect 31980 9865 32015 9900
rect 32025 9865 32060 9900
rect 32070 9865 32105 9900
rect 32115 9865 32150 9900
rect 32160 9865 32195 9900
rect 32205 9865 32240 9900
rect 32250 9865 32285 9900
rect 32295 9865 32330 9900
rect 32340 9865 32375 9900
rect 32385 9865 32420 9900
rect 32430 9865 32465 9900
rect 32475 9865 32510 9900
rect 32520 9865 32555 9900
rect 32565 9865 32600 9900
rect 32610 9865 32645 9900
rect 32655 9865 32690 9900
rect 32700 9865 32735 9900
rect 32745 9865 32780 9900
rect 32790 9865 32825 9900
rect 32835 9865 32870 9900
rect 31305 9820 31340 9855
rect 31350 9820 31385 9855
rect 31395 9820 31430 9855
rect 31440 9820 31475 9855
rect 31485 9820 31520 9855
rect 31530 9820 31565 9855
rect 31575 9820 31610 9855
rect 31620 9820 31655 9855
rect 31665 9820 31700 9855
rect 31710 9820 31745 9855
rect 31755 9820 31790 9855
rect 31800 9820 31835 9855
rect 31845 9820 31880 9855
rect 31890 9820 31925 9855
rect 31935 9820 31970 9855
rect 31980 9820 32015 9855
rect 32025 9820 32060 9855
rect 32070 9820 32105 9855
rect 32115 9820 32150 9855
rect 32160 9820 32195 9855
rect 32205 9820 32240 9855
rect 32250 9820 32285 9855
rect 32295 9820 32330 9855
rect 32340 9820 32375 9855
rect 32385 9820 32420 9855
rect 32430 9820 32465 9855
rect 32475 9820 32510 9855
rect 32520 9820 32555 9855
rect 32565 9820 32600 9855
rect 32610 9820 32645 9855
rect 32655 9820 32690 9855
rect 32700 9820 32735 9855
rect 32745 9820 32780 9855
rect 32790 9820 32825 9855
rect 32835 9820 32870 9855
rect 31305 9775 31340 9810
rect 31350 9775 31385 9810
rect 31395 9775 31430 9810
rect 31440 9775 31475 9810
rect 31485 9775 31520 9810
rect 31530 9775 31565 9810
rect 31575 9775 31610 9810
rect 31620 9775 31655 9810
rect 31665 9775 31700 9810
rect 31710 9775 31745 9810
rect 31755 9775 31790 9810
rect 31800 9775 31835 9810
rect 31845 9775 31880 9810
rect 31890 9775 31925 9810
rect 31935 9775 31970 9810
rect 31980 9775 32015 9810
rect 32025 9775 32060 9810
rect 32070 9775 32105 9810
rect 32115 9775 32150 9810
rect 32160 9775 32195 9810
rect 32205 9775 32240 9810
rect 32250 9775 32285 9810
rect 32295 9775 32330 9810
rect 32340 9775 32375 9810
rect 32385 9775 32420 9810
rect 32430 9775 32465 9810
rect 32475 9775 32510 9810
rect 32520 9775 32555 9810
rect 32565 9775 32600 9810
rect 32610 9775 32645 9810
rect 32655 9775 32690 9810
rect 32700 9775 32735 9810
rect 32745 9775 32780 9810
rect 32790 9775 32825 9810
rect 32835 9775 32870 9810
rect 31305 9730 31340 9765
rect 31350 9730 31385 9765
rect 31395 9730 31430 9765
rect 31440 9730 31475 9765
rect 31485 9730 31520 9765
rect 31530 9730 31565 9765
rect 31575 9730 31610 9765
rect 31620 9730 31655 9765
rect 31665 9730 31700 9765
rect 31710 9730 31745 9765
rect 31755 9730 31790 9765
rect 31800 9730 31835 9765
rect 31845 9730 31880 9765
rect 31890 9730 31925 9765
rect 31935 9730 31970 9765
rect 31980 9730 32015 9765
rect 32025 9730 32060 9765
rect 32070 9730 32105 9765
rect 32115 9730 32150 9765
rect 32160 9730 32195 9765
rect 32205 9730 32240 9765
rect 32250 9730 32285 9765
rect 32295 9730 32330 9765
rect 32340 9730 32375 9765
rect 32385 9730 32420 9765
rect 32430 9730 32465 9765
rect 32475 9730 32510 9765
rect 32520 9730 32555 9765
rect 32565 9730 32600 9765
rect 32610 9730 32645 9765
rect 32655 9730 32690 9765
rect 32700 9730 32735 9765
rect 32745 9730 32780 9765
rect 32790 9730 32825 9765
rect 32835 9730 32870 9765
rect 31305 9685 31340 9720
rect 31350 9685 31385 9720
rect 31395 9685 31430 9720
rect 31440 9685 31475 9720
rect 31485 9685 31520 9720
rect 31530 9685 31565 9720
rect 31575 9685 31610 9720
rect 31620 9685 31655 9720
rect 31665 9685 31700 9720
rect 31710 9685 31745 9720
rect 31755 9685 31790 9720
rect 31800 9685 31835 9720
rect 31845 9685 31880 9720
rect 31890 9685 31925 9720
rect 31935 9685 31970 9720
rect 31980 9685 32015 9720
rect 32025 9685 32060 9720
rect 32070 9685 32105 9720
rect 32115 9685 32150 9720
rect 32160 9685 32195 9720
rect 32205 9685 32240 9720
rect 32250 9685 32285 9720
rect 32295 9685 32330 9720
rect 32340 9685 32375 9720
rect 32385 9685 32420 9720
rect 32430 9685 32465 9720
rect 32475 9685 32510 9720
rect 32520 9685 32555 9720
rect 32565 9685 32600 9720
rect 32610 9685 32645 9720
rect 32655 9685 32690 9720
rect 32700 9685 32735 9720
rect 32745 9685 32780 9720
rect 32790 9685 32825 9720
rect 32835 9685 32870 9720
rect -38755 9595 -38720 9630
rect -38710 9595 -38675 9630
rect -38665 9595 -38630 9630
rect -38620 9595 -38585 9630
rect -38575 9595 -38540 9630
rect -38530 9595 -38495 9630
rect -38485 9595 -38450 9630
rect -38440 9595 -38405 9630
rect -38395 9595 -38360 9630
rect -38350 9595 -38315 9630
rect -38305 9595 -38270 9630
rect -38260 9595 -38225 9630
rect -38215 9595 -38180 9630
rect -38170 9595 -38135 9630
rect -38125 9595 -38090 9630
rect -38080 9595 -38045 9630
rect -38035 9595 -38000 9630
rect -37990 9595 -37955 9630
rect -37945 9595 -37910 9630
rect -37900 9595 -37865 9630
rect -37855 9595 -37820 9630
rect -37810 9595 -37775 9630
rect -37765 9595 -37730 9630
rect -37720 9595 -37685 9630
rect -37675 9595 -37640 9630
rect -37630 9595 -37595 9630
rect -37585 9595 -37550 9630
rect -37540 9595 -37505 9630
rect -37495 9595 -37460 9630
rect -37450 9595 -37415 9630
rect -37405 9595 -37370 9630
rect -37360 9595 -37325 9630
rect -37315 9595 -37280 9630
rect -37270 9595 -37235 9630
rect -37225 9595 -37190 9630
rect -38755 9550 -38720 9585
rect -38710 9550 -38675 9585
rect -38665 9550 -38630 9585
rect -38620 9550 -38585 9585
rect -38575 9550 -38540 9585
rect -38530 9550 -38495 9585
rect -38485 9550 -38450 9585
rect -38440 9550 -38405 9585
rect -38395 9550 -38360 9585
rect -38350 9550 -38315 9585
rect -38305 9550 -38270 9585
rect -38260 9550 -38225 9585
rect -38215 9550 -38180 9585
rect -38170 9550 -38135 9585
rect -38125 9550 -38090 9585
rect -38080 9550 -38045 9585
rect -38035 9550 -38000 9585
rect -37990 9550 -37955 9585
rect -37945 9550 -37910 9585
rect -37900 9550 -37865 9585
rect -37855 9550 -37820 9585
rect -37810 9550 -37775 9585
rect -37765 9550 -37730 9585
rect -37720 9550 -37685 9585
rect -37675 9550 -37640 9585
rect -37630 9550 -37595 9585
rect -37585 9550 -37550 9585
rect -37540 9550 -37505 9585
rect -37495 9550 -37460 9585
rect -37450 9550 -37415 9585
rect -37405 9550 -37370 9585
rect -37360 9550 -37325 9585
rect -37315 9550 -37280 9585
rect -37270 9550 -37235 9585
rect -37225 9550 -37190 9585
rect -38755 9505 -38720 9540
rect -38710 9505 -38675 9540
rect -38665 9505 -38630 9540
rect -38620 9505 -38585 9540
rect -38575 9505 -38540 9540
rect -38530 9505 -38495 9540
rect -38485 9505 -38450 9540
rect -38440 9505 -38405 9540
rect -38395 9505 -38360 9540
rect -38350 9505 -38315 9540
rect -38305 9505 -38270 9540
rect -38260 9505 -38225 9540
rect -38215 9505 -38180 9540
rect -38170 9505 -38135 9540
rect -38125 9505 -38090 9540
rect -38080 9505 -38045 9540
rect -38035 9505 -38000 9540
rect -37990 9505 -37955 9540
rect -37945 9505 -37910 9540
rect -37900 9505 -37865 9540
rect -37855 9505 -37820 9540
rect -37810 9505 -37775 9540
rect -37765 9505 -37730 9540
rect -37720 9505 -37685 9540
rect -37675 9505 -37640 9540
rect -37630 9505 -37595 9540
rect -37585 9505 -37550 9540
rect -37540 9505 -37505 9540
rect -37495 9505 -37460 9540
rect -37450 9505 -37415 9540
rect -37405 9505 -37370 9540
rect -37360 9505 -37325 9540
rect -37315 9505 -37280 9540
rect -37270 9505 -37235 9540
rect -37225 9505 -37190 9540
rect -38755 9460 -38720 9495
rect -38710 9460 -38675 9495
rect -38665 9460 -38630 9495
rect -38620 9460 -38585 9495
rect -38575 9460 -38540 9495
rect -38530 9460 -38495 9495
rect -38485 9460 -38450 9495
rect -38440 9460 -38405 9495
rect -38395 9460 -38360 9495
rect -38350 9460 -38315 9495
rect -38305 9460 -38270 9495
rect -38260 9460 -38225 9495
rect -38215 9460 -38180 9495
rect -38170 9460 -38135 9495
rect -38125 9460 -38090 9495
rect -38080 9460 -38045 9495
rect -38035 9460 -38000 9495
rect -37990 9460 -37955 9495
rect -37945 9460 -37910 9495
rect -37900 9460 -37865 9495
rect -37855 9460 -37820 9495
rect -37810 9460 -37775 9495
rect -37765 9460 -37730 9495
rect -37720 9460 -37685 9495
rect -37675 9460 -37640 9495
rect -37630 9460 -37595 9495
rect -37585 9460 -37550 9495
rect -37540 9460 -37505 9495
rect -37495 9460 -37460 9495
rect -37450 9460 -37415 9495
rect -37405 9460 -37370 9495
rect -37360 9460 -37325 9495
rect -37315 9460 -37280 9495
rect -37270 9460 -37235 9495
rect -37225 9460 -37190 9495
rect -38755 9415 -38720 9450
rect -38710 9415 -38675 9450
rect -38665 9415 -38630 9450
rect -38620 9415 -38585 9450
rect -38575 9415 -38540 9450
rect -38530 9415 -38495 9450
rect -38485 9415 -38450 9450
rect -38440 9415 -38405 9450
rect -38395 9415 -38360 9450
rect -38350 9415 -38315 9450
rect -38305 9415 -38270 9450
rect -38260 9415 -38225 9450
rect -38215 9415 -38180 9450
rect -38170 9415 -38135 9450
rect -38125 9415 -38090 9450
rect -38080 9415 -38045 9450
rect -38035 9415 -38000 9450
rect -37990 9415 -37955 9450
rect -37945 9415 -37910 9450
rect -37900 9415 -37865 9450
rect -37855 9415 -37820 9450
rect -37810 9415 -37775 9450
rect -37765 9415 -37730 9450
rect -37720 9415 -37685 9450
rect -37675 9415 -37640 9450
rect -37630 9415 -37595 9450
rect -37585 9415 -37550 9450
rect -37540 9415 -37505 9450
rect -37495 9415 -37460 9450
rect -37450 9415 -37415 9450
rect -37405 9415 -37370 9450
rect -37360 9415 -37325 9450
rect -37315 9415 -37280 9450
rect -37270 9415 -37235 9450
rect -37225 9415 -37190 9450
rect -38755 9370 -38720 9405
rect -38710 9370 -38675 9405
rect -38665 9370 -38630 9405
rect -38620 9370 -38585 9405
rect -38575 9370 -38540 9405
rect -38530 9370 -38495 9405
rect -38485 9370 -38450 9405
rect -38440 9370 -38405 9405
rect -38395 9370 -38360 9405
rect -38350 9370 -38315 9405
rect -38305 9370 -38270 9405
rect -38260 9370 -38225 9405
rect -38215 9370 -38180 9405
rect -38170 9370 -38135 9405
rect -38125 9370 -38090 9405
rect -38080 9370 -38045 9405
rect -38035 9370 -38000 9405
rect -37990 9370 -37955 9405
rect -37945 9370 -37910 9405
rect -37900 9370 -37865 9405
rect -37855 9370 -37820 9405
rect -37810 9370 -37775 9405
rect -37765 9370 -37730 9405
rect -37720 9370 -37685 9405
rect -37675 9370 -37640 9405
rect -37630 9370 -37595 9405
rect -37585 9370 -37550 9405
rect -37540 9370 -37505 9405
rect -37495 9370 -37460 9405
rect -37450 9370 -37415 9405
rect -37405 9370 -37370 9405
rect -37360 9370 -37325 9405
rect -37315 9370 -37280 9405
rect -37270 9370 -37235 9405
rect -37225 9370 -37190 9405
rect -38755 9325 -38720 9360
rect -38710 9325 -38675 9360
rect -38665 9325 -38630 9360
rect -38620 9325 -38585 9360
rect -38575 9325 -38540 9360
rect -38530 9325 -38495 9360
rect -38485 9325 -38450 9360
rect -38440 9325 -38405 9360
rect -38395 9325 -38360 9360
rect -38350 9325 -38315 9360
rect -38305 9325 -38270 9360
rect -38260 9325 -38225 9360
rect -38215 9325 -38180 9360
rect -38170 9325 -38135 9360
rect -38125 9325 -38090 9360
rect -38080 9325 -38045 9360
rect -38035 9325 -38000 9360
rect -37990 9325 -37955 9360
rect -37945 9325 -37910 9360
rect -37900 9325 -37865 9360
rect -37855 9325 -37820 9360
rect -37810 9325 -37775 9360
rect -37765 9325 -37730 9360
rect -37720 9325 -37685 9360
rect -37675 9325 -37640 9360
rect -37630 9325 -37595 9360
rect -37585 9325 -37550 9360
rect -37540 9325 -37505 9360
rect -37495 9325 -37460 9360
rect -37450 9325 -37415 9360
rect -37405 9325 -37370 9360
rect -37360 9325 -37325 9360
rect -37315 9325 -37280 9360
rect -37270 9325 -37235 9360
rect -37225 9325 -37190 9360
rect -38755 9280 -38720 9315
rect -38710 9280 -38675 9315
rect -38665 9280 -38630 9315
rect -38620 9280 -38585 9315
rect -38575 9280 -38540 9315
rect -38530 9280 -38495 9315
rect -38485 9280 -38450 9315
rect -38440 9280 -38405 9315
rect -38395 9280 -38360 9315
rect -38350 9280 -38315 9315
rect -38305 9280 -38270 9315
rect -38260 9280 -38225 9315
rect -38215 9280 -38180 9315
rect -38170 9280 -38135 9315
rect -38125 9280 -38090 9315
rect -38080 9280 -38045 9315
rect -38035 9280 -38000 9315
rect -37990 9280 -37955 9315
rect -37945 9280 -37910 9315
rect -37900 9280 -37865 9315
rect -37855 9280 -37820 9315
rect -37810 9280 -37775 9315
rect -37765 9280 -37730 9315
rect -37720 9280 -37685 9315
rect -37675 9280 -37640 9315
rect -37630 9280 -37595 9315
rect -37585 9280 -37550 9315
rect -37540 9280 -37505 9315
rect -37495 9280 -37460 9315
rect -37450 9280 -37415 9315
rect -37405 9280 -37370 9315
rect -37360 9280 -37325 9315
rect -37315 9280 -37280 9315
rect -37270 9280 -37235 9315
rect -37225 9280 -37190 9315
rect -38755 9235 -38720 9270
rect -38710 9235 -38675 9270
rect -38665 9235 -38630 9270
rect -38620 9235 -38585 9270
rect -38575 9235 -38540 9270
rect -38530 9235 -38495 9270
rect -38485 9235 -38450 9270
rect -38440 9235 -38405 9270
rect -38395 9235 -38360 9270
rect -38350 9235 -38315 9270
rect -38305 9235 -38270 9270
rect -38260 9235 -38225 9270
rect -38215 9235 -38180 9270
rect -38170 9235 -38135 9270
rect -38125 9235 -38090 9270
rect -38080 9235 -38045 9270
rect -38035 9235 -38000 9270
rect -37990 9235 -37955 9270
rect -37945 9235 -37910 9270
rect -37900 9235 -37865 9270
rect -37855 9235 -37820 9270
rect -37810 9235 -37775 9270
rect -37765 9235 -37730 9270
rect -37720 9235 -37685 9270
rect -37675 9235 -37640 9270
rect -37630 9235 -37595 9270
rect -37585 9235 -37550 9270
rect -37540 9235 -37505 9270
rect -37495 9235 -37460 9270
rect -37450 9235 -37415 9270
rect -37405 9235 -37370 9270
rect -37360 9235 -37325 9270
rect -37315 9235 -37280 9270
rect -37270 9235 -37235 9270
rect -37225 9235 -37190 9270
rect -38755 9190 -38720 9225
rect -38710 9190 -38675 9225
rect -38665 9190 -38630 9225
rect -38620 9190 -38585 9225
rect -38575 9190 -38540 9225
rect -38530 9190 -38495 9225
rect -38485 9190 -38450 9225
rect -38440 9190 -38405 9225
rect -38395 9190 -38360 9225
rect -38350 9190 -38315 9225
rect -38305 9190 -38270 9225
rect -38260 9190 -38225 9225
rect -38215 9190 -38180 9225
rect -38170 9190 -38135 9225
rect -38125 9190 -38090 9225
rect -38080 9190 -38045 9225
rect -38035 9190 -38000 9225
rect -37990 9190 -37955 9225
rect -37945 9190 -37910 9225
rect -37900 9190 -37865 9225
rect -37855 9190 -37820 9225
rect -37810 9190 -37775 9225
rect -37765 9190 -37730 9225
rect -37720 9190 -37685 9225
rect -37675 9190 -37640 9225
rect -37630 9190 -37595 9225
rect -37585 9190 -37550 9225
rect -37540 9190 -37505 9225
rect -37495 9190 -37460 9225
rect -37450 9190 -37415 9225
rect -37405 9190 -37370 9225
rect -37360 9190 -37325 9225
rect -37315 9190 -37280 9225
rect -37270 9190 -37235 9225
rect -37225 9190 -37190 9225
rect -38755 9145 -38720 9180
rect -38710 9145 -38675 9180
rect -38665 9145 -38630 9180
rect -38620 9145 -38585 9180
rect -38575 9145 -38540 9180
rect -38530 9145 -38495 9180
rect -38485 9145 -38450 9180
rect -38440 9145 -38405 9180
rect -38395 9145 -38360 9180
rect -38350 9145 -38315 9180
rect -38305 9145 -38270 9180
rect -38260 9145 -38225 9180
rect -38215 9145 -38180 9180
rect -38170 9145 -38135 9180
rect -38125 9145 -38090 9180
rect -38080 9145 -38045 9180
rect -38035 9145 -38000 9180
rect -37990 9145 -37955 9180
rect -37945 9145 -37910 9180
rect -37900 9145 -37865 9180
rect -37855 9145 -37820 9180
rect -37810 9145 -37775 9180
rect -37765 9145 -37730 9180
rect -37720 9145 -37685 9180
rect -37675 9145 -37640 9180
rect -37630 9145 -37595 9180
rect -37585 9145 -37550 9180
rect -37540 9145 -37505 9180
rect -37495 9145 -37460 9180
rect -37450 9145 -37415 9180
rect -37405 9145 -37370 9180
rect -37360 9145 -37325 9180
rect -37315 9145 -37280 9180
rect -37270 9145 -37235 9180
rect -37225 9145 -37190 9180
rect -38755 9100 -38720 9135
rect -38710 9100 -38675 9135
rect -38665 9100 -38630 9135
rect -38620 9100 -38585 9135
rect -38575 9100 -38540 9135
rect -38530 9100 -38495 9135
rect -38485 9100 -38450 9135
rect -38440 9100 -38405 9135
rect -38395 9100 -38360 9135
rect -38350 9100 -38315 9135
rect -38305 9100 -38270 9135
rect -38260 9100 -38225 9135
rect -38215 9100 -38180 9135
rect -38170 9100 -38135 9135
rect -38125 9100 -38090 9135
rect -38080 9100 -38045 9135
rect -38035 9100 -38000 9135
rect -37990 9100 -37955 9135
rect -37945 9100 -37910 9135
rect -37900 9100 -37865 9135
rect -37855 9100 -37820 9135
rect -37810 9100 -37775 9135
rect -37765 9100 -37730 9135
rect -37720 9100 -37685 9135
rect -37675 9100 -37640 9135
rect -37630 9100 -37595 9135
rect -37585 9100 -37550 9135
rect -37540 9100 -37505 9135
rect -37495 9100 -37460 9135
rect -37450 9100 -37415 9135
rect -37405 9100 -37370 9135
rect -37360 9100 -37325 9135
rect -37315 9100 -37280 9135
rect -37270 9100 -37235 9135
rect -37225 9100 -37190 9135
rect -38755 9055 -38720 9090
rect -38710 9055 -38675 9090
rect -38665 9055 -38630 9090
rect -38620 9055 -38585 9090
rect -38575 9055 -38540 9090
rect -38530 9055 -38495 9090
rect -38485 9055 -38450 9090
rect -38440 9055 -38405 9090
rect -38395 9055 -38360 9090
rect -38350 9055 -38315 9090
rect -38305 9055 -38270 9090
rect -38260 9055 -38225 9090
rect -38215 9055 -38180 9090
rect -38170 9055 -38135 9090
rect -38125 9055 -38090 9090
rect -38080 9055 -38045 9090
rect -38035 9055 -38000 9090
rect -37990 9055 -37955 9090
rect -37945 9055 -37910 9090
rect -37900 9055 -37865 9090
rect -37855 9055 -37820 9090
rect -37810 9055 -37775 9090
rect -37765 9055 -37730 9090
rect -37720 9055 -37685 9090
rect -37675 9055 -37640 9090
rect -37630 9055 -37595 9090
rect -37585 9055 -37550 9090
rect -37540 9055 -37505 9090
rect -37495 9055 -37460 9090
rect -37450 9055 -37415 9090
rect -37405 9055 -37370 9090
rect -37360 9055 -37325 9090
rect -37315 9055 -37280 9090
rect -37270 9055 -37235 9090
rect -37225 9055 -37190 9090
rect -38755 9010 -38720 9045
rect -38710 9010 -38675 9045
rect -38665 9010 -38630 9045
rect -38620 9010 -38585 9045
rect -38575 9010 -38540 9045
rect -38530 9010 -38495 9045
rect -38485 9010 -38450 9045
rect -38440 9010 -38405 9045
rect -38395 9010 -38360 9045
rect -38350 9010 -38315 9045
rect -38305 9010 -38270 9045
rect -38260 9010 -38225 9045
rect -38215 9010 -38180 9045
rect -38170 9010 -38135 9045
rect -38125 9010 -38090 9045
rect -38080 9010 -38045 9045
rect -38035 9010 -38000 9045
rect -37990 9010 -37955 9045
rect -37945 9010 -37910 9045
rect -37900 9010 -37865 9045
rect -37855 9010 -37820 9045
rect -37810 9010 -37775 9045
rect -37765 9010 -37730 9045
rect -37720 9010 -37685 9045
rect -37675 9010 -37640 9045
rect -37630 9010 -37595 9045
rect -37585 9010 -37550 9045
rect -37540 9010 -37505 9045
rect -37495 9010 -37460 9045
rect -37450 9010 -37415 9045
rect -37405 9010 -37370 9045
rect -37360 9010 -37325 9045
rect -37315 9010 -37280 9045
rect -37270 9010 -37235 9045
rect -37225 9010 -37190 9045
rect -38755 8965 -38720 9000
rect -38710 8965 -38675 9000
rect -38665 8965 -38630 9000
rect -38620 8965 -38585 9000
rect -38575 8965 -38540 9000
rect -38530 8965 -38495 9000
rect -38485 8965 -38450 9000
rect -38440 8965 -38405 9000
rect -38395 8965 -38360 9000
rect -38350 8965 -38315 9000
rect -38305 8965 -38270 9000
rect -38260 8965 -38225 9000
rect -38215 8965 -38180 9000
rect -38170 8965 -38135 9000
rect -38125 8965 -38090 9000
rect -38080 8965 -38045 9000
rect -38035 8965 -38000 9000
rect -37990 8965 -37955 9000
rect -37945 8965 -37910 9000
rect -37900 8965 -37865 9000
rect -37855 8965 -37820 9000
rect -37810 8965 -37775 9000
rect -37765 8965 -37730 9000
rect -37720 8965 -37685 9000
rect -37675 8965 -37640 9000
rect -37630 8965 -37595 9000
rect -37585 8965 -37550 9000
rect -37540 8965 -37505 9000
rect -37495 8965 -37460 9000
rect -37450 8965 -37415 9000
rect -37405 8965 -37370 9000
rect -37360 8965 -37325 9000
rect -37315 8965 -37280 9000
rect -37270 8965 -37235 9000
rect -37225 8965 -37190 9000
rect -38755 8920 -38720 8955
rect -38710 8920 -38675 8955
rect -38665 8920 -38630 8955
rect -38620 8920 -38585 8955
rect -38575 8920 -38540 8955
rect -38530 8920 -38495 8955
rect -38485 8920 -38450 8955
rect -38440 8920 -38405 8955
rect -38395 8920 -38360 8955
rect -38350 8920 -38315 8955
rect -38305 8920 -38270 8955
rect -38260 8920 -38225 8955
rect -38215 8920 -38180 8955
rect -38170 8920 -38135 8955
rect -38125 8920 -38090 8955
rect -38080 8920 -38045 8955
rect -38035 8920 -38000 8955
rect -37990 8920 -37955 8955
rect -37945 8920 -37910 8955
rect -37900 8920 -37865 8955
rect -37855 8920 -37820 8955
rect -37810 8920 -37775 8955
rect -37765 8920 -37730 8955
rect -37720 8920 -37685 8955
rect -37675 8920 -37640 8955
rect -37630 8920 -37595 8955
rect -37585 8920 -37550 8955
rect -37540 8920 -37505 8955
rect -37495 8920 -37460 8955
rect -37450 8920 -37415 8955
rect -37405 8920 -37370 8955
rect -37360 8920 -37325 8955
rect -37315 8920 -37280 8955
rect -37270 8920 -37235 8955
rect -37225 8920 -37190 8955
rect -38755 8875 -38720 8910
rect -38710 8875 -38675 8910
rect -38665 8875 -38630 8910
rect -38620 8875 -38585 8910
rect -38575 8875 -38540 8910
rect -38530 8875 -38495 8910
rect -38485 8875 -38450 8910
rect -38440 8875 -38405 8910
rect -38395 8875 -38360 8910
rect -38350 8875 -38315 8910
rect -38305 8875 -38270 8910
rect -38260 8875 -38225 8910
rect -38215 8875 -38180 8910
rect -38170 8875 -38135 8910
rect -38125 8875 -38090 8910
rect -38080 8875 -38045 8910
rect -38035 8875 -38000 8910
rect -37990 8875 -37955 8910
rect -37945 8875 -37910 8910
rect -37900 8875 -37865 8910
rect -37855 8875 -37820 8910
rect -37810 8875 -37775 8910
rect -37765 8875 -37730 8910
rect -37720 8875 -37685 8910
rect -37675 8875 -37640 8910
rect -37630 8875 -37595 8910
rect -37585 8875 -37550 8910
rect -37540 8875 -37505 8910
rect -37495 8875 -37460 8910
rect -37450 8875 -37415 8910
rect -37405 8875 -37370 8910
rect -37360 8875 -37325 8910
rect -37315 8875 -37280 8910
rect -37270 8875 -37235 8910
rect -37225 8875 -37190 8910
rect -38755 8830 -38720 8865
rect -38710 8830 -38675 8865
rect -38665 8830 -38630 8865
rect -38620 8830 -38585 8865
rect -38575 8830 -38540 8865
rect -38530 8830 -38495 8865
rect -38485 8830 -38450 8865
rect -38440 8830 -38405 8865
rect -38395 8830 -38360 8865
rect -38350 8830 -38315 8865
rect -38305 8830 -38270 8865
rect -38260 8830 -38225 8865
rect -38215 8830 -38180 8865
rect -38170 8830 -38135 8865
rect -38125 8830 -38090 8865
rect -38080 8830 -38045 8865
rect -38035 8830 -38000 8865
rect -37990 8830 -37955 8865
rect -37945 8830 -37910 8865
rect -37900 8830 -37865 8865
rect -37855 8830 -37820 8865
rect -37810 8830 -37775 8865
rect -37765 8830 -37730 8865
rect -37720 8830 -37685 8865
rect -37675 8830 -37640 8865
rect -37630 8830 -37595 8865
rect -37585 8830 -37550 8865
rect -37540 8830 -37505 8865
rect -37495 8830 -37460 8865
rect -37450 8830 -37415 8865
rect -37405 8830 -37370 8865
rect -37360 8830 -37325 8865
rect -37315 8830 -37280 8865
rect -37270 8830 -37235 8865
rect -37225 8830 -37190 8865
rect -38755 8785 -38720 8820
rect -38710 8785 -38675 8820
rect -38665 8785 -38630 8820
rect -38620 8785 -38585 8820
rect -38575 8785 -38540 8820
rect -38530 8785 -38495 8820
rect -38485 8785 -38450 8820
rect -38440 8785 -38405 8820
rect -38395 8785 -38360 8820
rect -38350 8785 -38315 8820
rect -38305 8785 -38270 8820
rect -38260 8785 -38225 8820
rect -38215 8785 -38180 8820
rect -38170 8785 -38135 8820
rect -38125 8785 -38090 8820
rect -38080 8785 -38045 8820
rect -38035 8785 -38000 8820
rect -37990 8785 -37955 8820
rect -37945 8785 -37910 8820
rect -37900 8785 -37865 8820
rect -37855 8785 -37820 8820
rect -37810 8785 -37775 8820
rect -37765 8785 -37730 8820
rect -37720 8785 -37685 8820
rect -37675 8785 -37640 8820
rect -37630 8785 -37595 8820
rect -37585 8785 -37550 8820
rect -37540 8785 -37505 8820
rect -37495 8785 -37460 8820
rect -37450 8785 -37415 8820
rect -37405 8785 -37370 8820
rect -37360 8785 -37325 8820
rect -37315 8785 -37280 8820
rect -37270 8785 -37235 8820
rect -37225 8785 -37190 8820
rect -38755 8740 -38720 8775
rect -38710 8740 -38675 8775
rect -38665 8740 -38630 8775
rect -38620 8740 -38585 8775
rect -38575 8740 -38540 8775
rect -38530 8740 -38495 8775
rect -38485 8740 -38450 8775
rect -38440 8740 -38405 8775
rect -38395 8740 -38360 8775
rect -38350 8740 -38315 8775
rect -38305 8740 -38270 8775
rect -38260 8740 -38225 8775
rect -38215 8740 -38180 8775
rect -38170 8740 -38135 8775
rect -38125 8740 -38090 8775
rect -38080 8740 -38045 8775
rect -38035 8740 -38000 8775
rect -37990 8740 -37955 8775
rect -37945 8740 -37910 8775
rect -37900 8740 -37865 8775
rect -37855 8740 -37820 8775
rect -37810 8740 -37775 8775
rect -37765 8740 -37730 8775
rect -37720 8740 -37685 8775
rect -37675 8740 -37640 8775
rect -37630 8740 -37595 8775
rect -37585 8740 -37550 8775
rect -37540 8740 -37505 8775
rect -37495 8740 -37460 8775
rect -37450 8740 -37415 8775
rect -37405 8740 -37370 8775
rect -37360 8740 -37325 8775
rect -37315 8740 -37280 8775
rect -37270 8740 -37235 8775
rect -37225 8740 -37190 8775
rect -38755 8695 -38720 8730
rect -38710 8695 -38675 8730
rect -38665 8695 -38630 8730
rect -38620 8695 -38585 8730
rect -38575 8695 -38540 8730
rect -38530 8695 -38495 8730
rect -38485 8695 -38450 8730
rect -38440 8695 -38405 8730
rect -38395 8695 -38360 8730
rect -38350 8695 -38315 8730
rect -38305 8695 -38270 8730
rect -38260 8695 -38225 8730
rect -38215 8695 -38180 8730
rect -38170 8695 -38135 8730
rect -38125 8695 -38090 8730
rect -38080 8695 -38045 8730
rect -38035 8695 -38000 8730
rect -37990 8695 -37955 8730
rect -37945 8695 -37910 8730
rect -37900 8695 -37865 8730
rect -37855 8695 -37820 8730
rect -37810 8695 -37775 8730
rect -37765 8695 -37730 8730
rect -37720 8695 -37685 8730
rect -37675 8695 -37640 8730
rect -37630 8695 -37595 8730
rect -37585 8695 -37550 8730
rect -37540 8695 -37505 8730
rect -37495 8695 -37460 8730
rect -37450 8695 -37415 8730
rect -37405 8695 -37370 8730
rect -37360 8695 -37325 8730
rect -37315 8695 -37280 8730
rect -37270 8695 -37235 8730
rect -37225 8695 -37190 8730
rect -38755 8650 -38720 8685
rect -38710 8650 -38675 8685
rect -38665 8650 -38630 8685
rect -38620 8650 -38585 8685
rect -38575 8650 -38540 8685
rect -38530 8650 -38495 8685
rect -38485 8650 -38450 8685
rect -38440 8650 -38405 8685
rect -38395 8650 -38360 8685
rect -38350 8650 -38315 8685
rect -38305 8650 -38270 8685
rect -38260 8650 -38225 8685
rect -38215 8650 -38180 8685
rect -38170 8650 -38135 8685
rect -38125 8650 -38090 8685
rect -38080 8650 -38045 8685
rect -38035 8650 -38000 8685
rect -37990 8650 -37955 8685
rect -37945 8650 -37910 8685
rect -37900 8650 -37865 8685
rect -37855 8650 -37820 8685
rect -37810 8650 -37775 8685
rect -37765 8650 -37730 8685
rect -37720 8650 -37685 8685
rect -37675 8650 -37640 8685
rect -37630 8650 -37595 8685
rect -37585 8650 -37550 8685
rect -37540 8650 -37505 8685
rect -37495 8650 -37460 8685
rect -37450 8650 -37415 8685
rect -37405 8650 -37370 8685
rect -37360 8650 -37325 8685
rect -37315 8650 -37280 8685
rect -37270 8650 -37235 8685
rect -37225 8650 -37190 8685
rect -38755 8605 -38720 8640
rect -38710 8605 -38675 8640
rect -38665 8605 -38630 8640
rect -38620 8605 -38585 8640
rect -38575 8605 -38540 8640
rect -38530 8605 -38495 8640
rect -38485 8605 -38450 8640
rect -38440 8605 -38405 8640
rect -38395 8605 -38360 8640
rect -38350 8605 -38315 8640
rect -38305 8605 -38270 8640
rect -38260 8605 -38225 8640
rect -38215 8605 -38180 8640
rect -38170 8605 -38135 8640
rect -38125 8605 -38090 8640
rect -38080 8605 -38045 8640
rect -38035 8605 -38000 8640
rect -37990 8605 -37955 8640
rect -37945 8605 -37910 8640
rect -37900 8605 -37865 8640
rect -37855 8605 -37820 8640
rect -37810 8605 -37775 8640
rect -37765 8605 -37730 8640
rect -37720 8605 -37685 8640
rect -37675 8605 -37640 8640
rect -37630 8605 -37595 8640
rect -37585 8605 -37550 8640
rect -37540 8605 -37505 8640
rect -37495 8605 -37460 8640
rect -37450 8605 -37415 8640
rect -37405 8605 -37370 8640
rect -37360 8605 -37325 8640
rect -37315 8605 -37280 8640
rect -37270 8605 -37235 8640
rect -37225 8605 -37190 8640
rect -38755 8560 -38720 8595
rect -38710 8560 -38675 8595
rect -38665 8560 -38630 8595
rect -38620 8560 -38585 8595
rect -38575 8560 -38540 8595
rect -38530 8560 -38495 8595
rect -38485 8560 -38450 8595
rect -38440 8560 -38405 8595
rect -38395 8560 -38360 8595
rect -38350 8560 -38315 8595
rect -38305 8560 -38270 8595
rect -38260 8560 -38225 8595
rect -38215 8560 -38180 8595
rect -38170 8560 -38135 8595
rect -38125 8560 -38090 8595
rect -38080 8560 -38045 8595
rect -38035 8560 -38000 8595
rect -37990 8560 -37955 8595
rect -37945 8560 -37910 8595
rect -37900 8560 -37865 8595
rect -37855 8560 -37820 8595
rect -37810 8560 -37775 8595
rect -37765 8560 -37730 8595
rect -37720 8560 -37685 8595
rect -37675 8560 -37640 8595
rect -37630 8560 -37595 8595
rect -37585 8560 -37550 8595
rect -37540 8560 -37505 8595
rect -37495 8560 -37460 8595
rect -37450 8560 -37415 8595
rect -37405 8560 -37370 8595
rect -37360 8560 -37325 8595
rect -37315 8560 -37280 8595
rect -37270 8560 -37235 8595
rect -37225 8560 -37190 8595
rect -38755 8515 -38720 8550
rect -38710 8515 -38675 8550
rect -38665 8515 -38630 8550
rect -38620 8515 -38585 8550
rect -38575 8515 -38540 8550
rect -38530 8515 -38495 8550
rect -38485 8515 -38450 8550
rect -38440 8515 -38405 8550
rect -38395 8515 -38360 8550
rect -38350 8515 -38315 8550
rect -38305 8515 -38270 8550
rect -38260 8515 -38225 8550
rect -38215 8515 -38180 8550
rect -38170 8515 -38135 8550
rect -38125 8515 -38090 8550
rect -38080 8515 -38045 8550
rect -38035 8515 -38000 8550
rect -37990 8515 -37955 8550
rect -37945 8515 -37910 8550
rect -37900 8515 -37865 8550
rect -37855 8515 -37820 8550
rect -37810 8515 -37775 8550
rect -37765 8515 -37730 8550
rect -37720 8515 -37685 8550
rect -37675 8515 -37640 8550
rect -37630 8515 -37595 8550
rect -37585 8515 -37550 8550
rect -37540 8515 -37505 8550
rect -37495 8515 -37460 8550
rect -37450 8515 -37415 8550
rect -37405 8515 -37370 8550
rect -37360 8515 -37325 8550
rect -37315 8515 -37280 8550
rect -37270 8515 -37235 8550
rect -37225 8515 -37190 8550
rect -38755 8470 -38720 8505
rect -38710 8470 -38675 8505
rect -38665 8470 -38630 8505
rect -38620 8470 -38585 8505
rect -38575 8470 -38540 8505
rect -38530 8470 -38495 8505
rect -38485 8470 -38450 8505
rect -38440 8470 -38405 8505
rect -38395 8470 -38360 8505
rect -38350 8470 -38315 8505
rect -38305 8470 -38270 8505
rect -38260 8470 -38225 8505
rect -38215 8470 -38180 8505
rect -38170 8470 -38135 8505
rect -38125 8470 -38090 8505
rect -38080 8470 -38045 8505
rect -38035 8470 -38000 8505
rect -37990 8470 -37955 8505
rect -37945 8470 -37910 8505
rect -37900 8470 -37865 8505
rect -37855 8470 -37820 8505
rect -37810 8470 -37775 8505
rect -37765 8470 -37730 8505
rect -37720 8470 -37685 8505
rect -37675 8470 -37640 8505
rect -37630 8470 -37595 8505
rect -37585 8470 -37550 8505
rect -37540 8470 -37505 8505
rect -37495 8470 -37460 8505
rect -37450 8470 -37415 8505
rect -37405 8470 -37370 8505
rect -37360 8470 -37325 8505
rect -37315 8470 -37280 8505
rect -37270 8470 -37235 8505
rect -37225 8470 -37190 8505
rect -38755 8425 -38720 8460
rect -38710 8425 -38675 8460
rect -38665 8425 -38630 8460
rect -38620 8425 -38585 8460
rect -38575 8425 -38540 8460
rect -38530 8425 -38495 8460
rect -38485 8425 -38450 8460
rect -38440 8425 -38405 8460
rect -38395 8425 -38360 8460
rect -38350 8425 -38315 8460
rect -38305 8425 -38270 8460
rect -38260 8425 -38225 8460
rect -38215 8425 -38180 8460
rect -38170 8425 -38135 8460
rect -38125 8425 -38090 8460
rect -38080 8425 -38045 8460
rect -38035 8425 -38000 8460
rect -37990 8425 -37955 8460
rect -37945 8425 -37910 8460
rect -37900 8425 -37865 8460
rect -37855 8425 -37820 8460
rect -37810 8425 -37775 8460
rect -37765 8425 -37730 8460
rect -37720 8425 -37685 8460
rect -37675 8425 -37640 8460
rect -37630 8425 -37595 8460
rect -37585 8425 -37550 8460
rect -37540 8425 -37505 8460
rect -37495 8425 -37460 8460
rect -37450 8425 -37415 8460
rect -37405 8425 -37370 8460
rect -37360 8425 -37325 8460
rect -37315 8425 -37280 8460
rect -37270 8425 -37235 8460
rect -37225 8425 -37190 8460
rect -38755 8380 -38720 8415
rect -38710 8380 -38675 8415
rect -38665 8380 -38630 8415
rect -38620 8380 -38585 8415
rect -38575 8380 -38540 8415
rect -38530 8380 -38495 8415
rect -38485 8380 -38450 8415
rect -38440 8380 -38405 8415
rect -38395 8380 -38360 8415
rect -38350 8380 -38315 8415
rect -38305 8380 -38270 8415
rect -38260 8380 -38225 8415
rect -38215 8380 -38180 8415
rect -38170 8380 -38135 8415
rect -38125 8380 -38090 8415
rect -38080 8380 -38045 8415
rect -38035 8380 -38000 8415
rect -37990 8380 -37955 8415
rect -37945 8380 -37910 8415
rect -37900 8380 -37865 8415
rect -37855 8380 -37820 8415
rect -37810 8380 -37775 8415
rect -37765 8380 -37730 8415
rect -37720 8380 -37685 8415
rect -37675 8380 -37640 8415
rect -37630 8380 -37595 8415
rect -37585 8380 -37550 8415
rect -37540 8380 -37505 8415
rect -37495 8380 -37460 8415
rect -37450 8380 -37415 8415
rect -37405 8380 -37370 8415
rect -37360 8380 -37325 8415
rect -37315 8380 -37280 8415
rect -37270 8380 -37235 8415
rect -37225 8380 -37190 8415
rect -38755 8335 -38720 8370
rect -38710 8335 -38675 8370
rect -38665 8335 -38630 8370
rect -38620 8335 -38585 8370
rect -38575 8335 -38540 8370
rect -38530 8335 -38495 8370
rect -38485 8335 -38450 8370
rect -38440 8335 -38405 8370
rect -38395 8335 -38360 8370
rect -38350 8335 -38315 8370
rect -38305 8335 -38270 8370
rect -38260 8335 -38225 8370
rect -38215 8335 -38180 8370
rect -38170 8335 -38135 8370
rect -38125 8335 -38090 8370
rect -38080 8335 -38045 8370
rect -38035 8335 -38000 8370
rect -37990 8335 -37955 8370
rect -37945 8335 -37910 8370
rect -37900 8335 -37865 8370
rect -37855 8335 -37820 8370
rect -37810 8335 -37775 8370
rect -37765 8335 -37730 8370
rect -37720 8335 -37685 8370
rect -37675 8335 -37640 8370
rect -37630 8335 -37595 8370
rect -37585 8335 -37550 8370
rect -37540 8335 -37505 8370
rect -37495 8335 -37460 8370
rect -37450 8335 -37415 8370
rect -37405 8335 -37370 8370
rect -37360 8335 -37325 8370
rect -37315 8335 -37280 8370
rect -37270 8335 -37235 8370
rect -37225 8335 -37190 8370
rect -38755 8290 -38720 8325
rect -38710 8290 -38675 8325
rect -38665 8290 -38630 8325
rect -38620 8290 -38585 8325
rect -38575 8290 -38540 8325
rect -38530 8290 -38495 8325
rect -38485 8290 -38450 8325
rect -38440 8290 -38405 8325
rect -38395 8290 -38360 8325
rect -38350 8290 -38315 8325
rect -38305 8290 -38270 8325
rect -38260 8290 -38225 8325
rect -38215 8290 -38180 8325
rect -38170 8290 -38135 8325
rect -38125 8290 -38090 8325
rect -38080 8290 -38045 8325
rect -38035 8290 -38000 8325
rect -37990 8290 -37955 8325
rect -37945 8290 -37910 8325
rect -37900 8290 -37865 8325
rect -37855 8290 -37820 8325
rect -37810 8290 -37775 8325
rect -37765 8290 -37730 8325
rect -37720 8290 -37685 8325
rect -37675 8290 -37640 8325
rect -37630 8290 -37595 8325
rect -37585 8290 -37550 8325
rect -37540 8290 -37505 8325
rect -37495 8290 -37460 8325
rect -37450 8290 -37415 8325
rect -37405 8290 -37370 8325
rect -37360 8290 -37325 8325
rect -37315 8290 -37280 8325
rect -37270 8290 -37235 8325
rect -37225 8290 -37190 8325
rect -38755 8245 -38720 8280
rect -38710 8245 -38675 8280
rect -38665 8245 -38630 8280
rect -38620 8245 -38585 8280
rect -38575 8245 -38540 8280
rect -38530 8245 -38495 8280
rect -38485 8245 -38450 8280
rect -38440 8245 -38405 8280
rect -38395 8245 -38360 8280
rect -38350 8245 -38315 8280
rect -38305 8245 -38270 8280
rect -38260 8245 -38225 8280
rect -38215 8245 -38180 8280
rect -38170 8245 -38135 8280
rect -38125 8245 -38090 8280
rect -38080 8245 -38045 8280
rect -38035 8245 -38000 8280
rect -37990 8245 -37955 8280
rect -37945 8245 -37910 8280
rect -37900 8245 -37865 8280
rect -37855 8245 -37820 8280
rect -37810 8245 -37775 8280
rect -37765 8245 -37730 8280
rect -37720 8245 -37685 8280
rect -37675 8245 -37640 8280
rect -37630 8245 -37595 8280
rect -37585 8245 -37550 8280
rect -37540 8245 -37505 8280
rect -37495 8245 -37460 8280
rect -37450 8245 -37415 8280
rect -37405 8245 -37370 8280
rect -37360 8245 -37325 8280
rect -37315 8245 -37280 8280
rect -37270 8245 -37235 8280
rect -37225 8245 -37190 8280
rect -38755 8200 -38720 8235
rect -38710 8200 -38675 8235
rect -38665 8200 -38630 8235
rect -38620 8200 -38585 8235
rect -38575 8200 -38540 8235
rect -38530 8200 -38495 8235
rect -38485 8200 -38450 8235
rect -38440 8200 -38405 8235
rect -38395 8200 -38360 8235
rect -38350 8200 -38315 8235
rect -38305 8200 -38270 8235
rect -38260 8200 -38225 8235
rect -38215 8200 -38180 8235
rect -38170 8200 -38135 8235
rect -38125 8200 -38090 8235
rect -38080 8200 -38045 8235
rect -38035 8200 -38000 8235
rect -37990 8200 -37955 8235
rect -37945 8200 -37910 8235
rect -37900 8200 -37865 8235
rect -37855 8200 -37820 8235
rect -37810 8200 -37775 8235
rect -37765 8200 -37730 8235
rect -37720 8200 -37685 8235
rect -37675 8200 -37640 8235
rect -37630 8200 -37595 8235
rect -37585 8200 -37550 8235
rect -37540 8200 -37505 8235
rect -37495 8200 -37460 8235
rect -37450 8200 -37415 8235
rect -37405 8200 -37370 8235
rect -37360 8200 -37325 8235
rect -37315 8200 -37280 8235
rect -37270 8200 -37235 8235
rect -37225 8200 -37190 8235
rect -38755 8155 -38720 8190
rect -38710 8155 -38675 8190
rect -38665 8155 -38630 8190
rect -38620 8155 -38585 8190
rect -38575 8155 -38540 8190
rect -38530 8155 -38495 8190
rect -38485 8155 -38450 8190
rect -38440 8155 -38405 8190
rect -38395 8155 -38360 8190
rect -38350 8155 -38315 8190
rect -38305 8155 -38270 8190
rect -38260 8155 -38225 8190
rect -38215 8155 -38180 8190
rect -38170 8155 -38135 8190
rect -38125 8155 -38090 8190
rect -38080 8155 -38045 8190
rect -38035 8155 -38000 8190
rect -37990 8155 -37955 8190
rect -37945 8155 -37910 8190
rect -37900 8155 -37865 8190
rect -37855 8155 -37820 8190
rect -37810 8155 -37775 8190
rect -37765 8155 -37730 8190
rect -37720 8155 -37685 8190
rect -37675 8155 -37640 8190
rect -37630 8155 -37595 8190
rect -37585 8155 -37550 8190
rect -37540 8155 -37505 8190
rect -37495 8155 -37460 8190
rect -37450 8155 -37415 8190
rect -37405 8155 -37370 8190
rect -37360 8155 -37325 8190
rect -37315 8155 -37280 8190
rect -37270 8155 -37235 8190
rect -37225 8155 -37190 8190
rect -38755 8110 -38720 8145
rect -38710 8110 -38675 8145
rect -38665 8110 -38630 8145
rect -38620 8110 -38585 8145
rect -38575 8110 -38540 8145
rect -38530 8110 -38495 8145
rect -38485 8110 -38450 8145
rect -38440 8110 -38405 8145
rect -38395 8110 -38360 8145
rect -38350 8110 -38315 8145
rect -38305 8110 -38270 8145
rect -38260 8110 -38225 8145
rect -38215 8110 -38180 8145
rect -38170 8110 -38135 8145
rect -38125 8110 -38090 8145
rect -38080 8110 -38045 8145
rect -38035 8110 -38000 8145
rect -37990 8110 -37955 8145
rect -37945 8110 -37910 8145
rect -37900 8110 -37865 8145
rect -37855 8110 -37820 8145
rect -37810 8110 -37775 8145
rect -37765 8110 -37730 8145
rect -37720 8110 -37685 8145
rect -37675 8110 -37640 8145
rect -37630 8110 -37595 8145
rect -37585 8110 -37550 8145
rect -37540 8110 -37505 8145
rect -37495 8110 -37460 8145
rect -37450 8110 -37415 8145
rect -37405 8110 -37370 8145
rect -37360 8110 -37325 8145
rect -37315 8110 -37280 8145
rect -37270 8110 -37235 8145
rect -37225 8110 -37190 8145
rect 1320 9635 1360 9640
rect 1320 9605 1325 9635
rect 1325 9605 1355 9635
rect 1355 9605 1360 9635
rect 1320 9600 1360 9605
rect 1320 9570 1360 9575
rect 1320 9540 1325 9570
rect 1325 9540 1355 9570
rect 1355 9540 1360 9570
rect 1320 9535 1360 9540
rect 1320 9500 1360 9505
rect 1320 9470 1325 9500
rect 1325 9470 1355 9500
rect 1355 9470 1360 9500
rect 1320 9465 1360 9470
rect 1320 9430 1360 9435
rect 1320 9400 1325 9430
rect 1325 9400 1355 9430
rect 1355 9400 1360 9430
rect 1320 9395 1360 9400
rect 1320 9360 1360 9365
rect 1320 9330 1325 9360
rect 1325 9330 1355 9360
rect 1355 9330 1360 9360
rect 1320 9325 1360 9330
rect 1320 9295 1360 9300
rect 1320 9265 1325 9295
rect 1325 9265 1355 9295
rect 1355 9265 1360 9295
rect 1320 9260 1360 9265
rect 1320 9235 1360 9240
rect 1320 9205 1325 9235
rect 1325 9205 1355 9235
rect 1355 9205 1360 9235
rect 1320 9200 1360 9205
rect 1320 9170 1360 9175
rect 1320 9140 1325 9170
rect 1325 9140 1355 9170
rect 1355 9140 1360 9170
rect 1320 9135 1360 9140
rect 1320 9100 1360 9105
rect 1320 9070 1325 9100
rect 1325 9070 1355 9100
rect 1355 9070 1360 9100
rect 1320 9065 1360 9070
rect 1320 9030 1360 9035
rect 1320 9000 1325 9030
rect 1325 9000 1355 9030
rect 1355 9000 1360 9030
rect 1320 8995 1360 9000
rect 1320 8960 1360 8965
rect 1320 8930 1325 8960
rect 1325 8930 1355 8960
rect 1355 8930 1360 8960
rect 1320 8925 1360 8930
rect 1320 8895 1360 8900
rect 1320 8865 1325 8895
rect 1325 8865 1355 8895
rect 1355 8865 1360 8895
rect 1320 8860 1360 8865
rect 1320 8835 1360 8840
rect 1320 8805 1325 8835
rect 1325 8805 1355 8835
rect 1355 8805 1360 8835
rect 1320 8800 1360 8805
rect 1320 8770 1360 8775
rect 1320 8740 1325 8770
rect 1325 8740 1355 8770
rect 1355 8740 1360 8770
rect 1320 8735 1360 8740
rect 1320 8700 1360 8705
rect 1320 8670 1325 8700
rect 1325 8670 1355 8700
rect 1355 8670 1360 8700
rect 1320 8665 1360 8670
rect 1320 8630 1360 8635
rect 1320 8600 1325 8630
rect 1325 8600 1355 8630
rect 1355 8600 1360 8630
rect 1320 8595 1360 8600
rect 1320 8560 1360 8565
rect 1320 8530 1325 8560
rect 1325 8530 1355 8560
rect 1355 8530 1360 8560
rect 1320 8525 1360 8530
rect 1320 8495 1360 8500
rect 1320 8465 1325 8495
rect 1325 8465 1355 8495
rect 1355 8465 1360 8495
rect 1320 8460 1360 8465
rect 1320 8435 1360 8440
rect 1320 8405 1325 8435
rect 1325 8405 1355 8435
rect 1355 8405 1360 8435
rect 1320 8400 1360 8405
rect 1320 8370 1360 8375
rect 1320 8340 1325 8370
rect 1325 8340 1355 8370
rect 1355 8340 1360 8370
rect 1320 8335 1360 8340
rect 1320 8300 1360 8305
rect 1320 8270 1325 8300
rect 1325 8270 1355 8300
rect 1355 8270 1360 8300
rect 1320 8265 1360 8270
rect 1320 8230 1360 8235
rect 1320 8200 1325 8230
rect 1325 8200 1355 8230
rect 1355 8200 1360 8230
rect 1320 8195 1360 8200
rect 1320 8160 1360 8165
rect 1320 8130 1325 8160
rect 1325 8130 1355 8160
rect 1355 8130 1360 8160
rect 1320 8125 1360 8130
rect 2245 9635 2285 9640
rect 2245 9605 2250 9635
rect 2250 9605 2280 9635
rect 2280 9605 2285 9635
rect 2245 9600 2285 9605
rect 2245 9570 2285 9575
rect 2245 9540 2250 9570
rect 2250 9540 2280 9570
rect 2280 9540 2285 9570
rect 2245 9535 2285 9540
rect 2245 9500 2285 9505
rect 2245 9470 2250 9500
rect 2250 9470 2280 9500
rect 2280 9470 2285 9500
rect 2245 9465 2285 9470
rect 2245 9430 2285 9435
rect 2245 9400 2250 9430
rect 2250 9400 2280 9430
rect 2280 9400 2285 9430
rect 2245 9395 2285 9400
rect 2245 9360 2285 9365
rect 2245 9330 2250 9360
rect 2250 9330 2280 9360
rect 2280 9330 2285 9360
rect 2245 9325 2285 9330
rect 2245 9295 2285 9300
rect 2245 9265 2250 9295
rect 2250 9265 2280 9295
rect 2280 9265 2285 9295
rect 2245 9260 2285 9265
rect 2245 9235 2285 9240
rect 2245 9205 2250 9235
rect 2250 9205 2280 9235
rect 2280 9205 2285 9235
rect 2245 9200 2285 9205
rect 2245 9170 2285 9175
rect 2245 9140 2250 9170
rect 2250 9140 2280 9170
rect 2280 9140 2285 9170
rect 2245 9135 2285 9140
rect 2245 9100 2285 9105
rect 2245 9070 2250 9100
rect 2250 9070 2280 9100
rect 2280 9070 2285 9100
rect 2245 9065 2285 9070
rect 2245 9030 2285 9035
rect 2245 9000 2250 9030
rect 2250 9000 2280 9030
rect 2280 9000 2285 9030
rect 2245 8995 2285 9000
rect 2245 8960 2285 8965
rect 2245 8930 2250 8960
rect 2250 8930 2280 8960
rect 2280 8930 2285 8960
rect 2245 8925 2285 8930
rect 2245 8895 2285 8900
rect 2245 8865 2250 8895
rect 2250 8865 2280 8895
rect 2280 8865 2285 8895
rect 2245 8860 2285 8865
rect 2245 8835 2285 8840
rect 2245 8805 2250 8835
rect 2250 8805 2280 8835
rect 2280 8805 2285 8835
rect 2245 8800 2285 8805
rect 2245 8770 2285 8775
rect 2245 8740 2250 8770
rect 2250 8740 2280 8770
rect 2280 8740 2285 8770
rect 2245 8735 2285 8740
rect 2245 8700 2285 8705
rect 2245 8670 2250 8700
rect 2250 8670 2280 8700
rect 2280 8670 2285 8700
rect 2245 8665 2285 8670
rect 2245 8630 2285 8635
rect 2245 8600 2250 8630
rect 2250 8600 2280 8630
rect 2280 8600 2285 8630
rect 2245 8595 2285 8600
rect 2245 8560 2285 8565
rect 2245 8530 2250 8560
rect 2250 8530 2280 8560
rect 2280 8530 2285 8560
rect 2245 8525 2285 8530
rect 2245 8495 2285 8500
rect 2245 8465 2250 8495
rect 2250 8465 2280 8495
rect 2280 8465 2285 8495
rect 2245 8460 2285 8465
rect 2245 8435 2285 8440
rect 2245 8405 2250 8435
rect 2250 8405 2280 8435
rect 2280 8405 2285 8435
rect 2245 8400 2285 8405
rect 2245 8370 2285 8375
rect 2245 8340 2250 8370
rect 2250 8340 2280 8370
rect 2280 8340 2285 8370
rect 2245 8335 2285 8340
rect 2245 8300 2285 8305
rect 2245 8270 2250 8300
rect 2250 8270 2280 8300
rect 2280 8270 2285 8300
rect 2245 8265 2285 8270
rect 2245 8230 2285 8235
rect 2245 8200 2250 8230
rect 2250 8200 2280 8230
rect 2280 8200 2285 8230
rect 2245 8195 2285 8200
rect 2245 8160 2285 8165
rect 2245 8130 2250 8160
rect 2250 8130 2280 8160
rect 2280 8130 2285 8160
rect 2245 8125 2285 8130
rect 3175 9635 3215 9640
rect 3175 9605 3180 9635
rect 3180 9605 3210 9635
rect 3210 9605 3215 9635
rect 3175 9600 3215 9605
rect 3175 9570 3215 9575
rect 3175 9540 3180 9570
rect 3180 9540 3210 9570
rect 3210 9540 3215 9570
rect 3175 9535 3215 9540
rect 3175 9500 3215 9505
rect 3175 9470 3180 9500
rect 3180 9470 3210 9500
rect 3210 9470 3215 9500
rect 3175 9465 3215 9470
rect 3175 9430 3215 9435
rect 3175 9400 3180 9430
rect 3180 9400 3210 9430
rect 3210 9400 3215 9430
rect 3175 9395 3215 9400
rect 3175 9360 3215 9365
rect 3175 9330 3180 9360
rect 3180 9330 3210 9360
rect 3210 9330 3215 9360
rect 3175 9325 3215 9330
rect 3175 9295 3215 9300
rect 3175 9265 3180 9295
rect 3180 9265 3210 9295
rect 3210 9265 3215 9295
rect 3175 9260 3215 9265
rect 3175 9235 3215 9240
rect 3175 9205 3180 9235
rect 3180 9205 3210 9235
rect 3210 9205 3215 9235
rect 3175 9200 3215 9205
rect 3175 9170 3215 9175
rect 3175 9140 3180 9170
rect 3180 9140 3210 9170
rect 3210 9140 3215 9170
rect 3175 9135 3215 9140
rect 3175 9100 3215 9105
rect 3175 9070 3180 9100
rect 3180 9070 3210 9100
rect 3210 9070 3215 9100
rect 3175 9065 3215 9070
rect 3175 9030 3215 9035
rect 3175 9000 3180 9030
rect 3180 9000 3210 9030
rect 3210 9000 3215 9030
rect 3175 8995 3215 9000
rect 3175 8960 3215 8965
rect 3175 8930 3180 8960
rect 3180 8930 3210 8960
rect 3210 8930 3215 8960
rect 3175 8925 3215 8930
rect 3175 8895 3215 8900
rect 3175 8865 3180 8895
rect 3180 8865 3210 8895
rect 3210 8865 3215 8895
rect 3175 8860 3215 8865
rect 3175 8835 3215 8840
rect 3175 8805 3180 8835
rect 3180 8805 3210 8835
rect 3210 8805 3215 8835
rect 3175 8800 3215 8805
rect 3175 8770 3215 8775
rect 3175 8740 3180 8770
rect 3180 8740 3210 8770
rect 3210 8740 3215 8770
rect 3175 8735 3215 8740
rect 3175 8700 3215 8705
rect 3175 8670 3180 8700
rect 3180 8670 3210 8700
rect 3210 8670 3215 8700
rect 3175 8665 3215 8670
rect 3175 8630 3215 8635
rect 3175 8600 3180 8630
rect 3180 8600 3210 8630
rect 3210 8600 3215 8630
rect 3175 8595 3215 8600
rect 3175 8560 3215 8565
rect 3175 8530 3180 8560
rect 3180 8530 3210 8560
rect 3210 8530 3215 8560
rect 3175 8525 3215 8530
rect 3175 8495 3215 8500
rect 3175 8465 3180 8495
rect 3180 8465 3210 8495
rect 3210 8465 3215 8495
rect 3175 8460 3215 8465
rect 3175 8435 3215 8440
rect 3175 8405 3180 8435
rect 3180 8405 3210 8435
rect 3210 8405 3215 8435
rect 3175 8400 3215 8405
rect 3175 8370 3215 8375
rect 3175 8340 3180 8370
rect 3180 8340 3210 8370
rect 3210 8340 3215 8370
rect 3175 8335 3215 8340
rect 3175 8300 3215 8305
rect 3175 8270 3180 8300
rect 3180 8270 3210 8300
rect 3210 8270 3215 8300
rect 3175 8265 3215 8270
rect 3175 8230 3215 8235
rect 3175 8200 3180 8230
rect 3180 8200 3210 8230
rect 3210 8200 3215 8230
rect 3175 8195 3215 8200
rect 3175 8160 3215 8165
rect 3175 8130 3180 8160
rect 3180 8130 3210 8160
rect 3210 8130 3215 8160
rect 3175 8125 3215 8130
rect 6700 9635 6740 9640
rect 6700 9605 6705 9635
rect 6705 9605 6735 9635
rect 6735 9605 6740 9635
rect 6700 9600 6740 9605
rect 6700 9570 6740 9575
rect 6700 9540 6705 9570
rect 6705 9540 6735 9570
rect 6735 9540 6740 9570
rect 6700 9535 6740 9540
rect 6700 9500 6740 9505
rect 6700 9470 6705 9500
rect 6705 9470 6735 9500
rect 6735 9470 6740 9500
rect 6700 9465 6740 9470
rect 6700 9430 6740 9435
rect 6700 9400 6705 9430
rect 6705 9400 6735 9430
rect 6735 9400 6740 9430
rect 6700 9395 6740 9400
rect 6700 9360 6740 9365
rect 6700 9330 6705 9360
rect 6705 9330 6735 9360
rect 6735 9330 6740 9360
rect 6700 9325 6740 9330
rect 6700 9295 6740 9300
rect 6700 9265 6705 9295
rect 6705 9265 6735 9295
rect 6735 9265 6740 9295
rect 6700 9260 6740 9265
rect 6700 9235 6740 9240
rect 6700 9205 6705 9235
rect 6705 9205 6735 9235
rect 6735 9205 6740 9235
rect 6700 9200 6740 9205
rect 6700 9170 6740 9175
rect 6700 9140 6705 9170
rect 6705 9140 6735 9170
rect 6735 9140 6740 9170
rect 6700 9135 6740 9140
rect 6700 9100 6740 9105
rect 6700 9070 6705 9100
rect 6705 9070 6735 9100
rect 6735 9070 6740 9100
rect 6700 9065 6740 9070
rect 6700 9030 6740 9035
rect 6700 9000 6705 9030
rect 6705 9000 6735 9030
rect 6735 9000 6740 9030
rect 6700 8995 6740 9000
rect 6700 8960 6740 8965
rect 6700 8930 6705 8960
rect 6705 8930 6735 8960
rect 6735 8930 6740 8960
rect 6700 8925 6740 8930
rect 6700 8895 6740 8900
rect 6700 8865 6705 8895
rect 6705 8865 6735 8895
rect 6735 8865 6740 8895
rect 6700 8860 6740 8865
rect 6700 8835 6740 8840
rect 6700 8805 6705 8835
rect 6705 8805 6735 8835
rect 6735 8805 6740 8835
rect 6700 8800 6740 8805
rect 6700 8770 6740 8775
rect 6700 8740 6705 8770
rect 6705 8740 6735 8770
rect 6735 8740 6740 8770
rect 6700 8735 6740 8740
rect 6700 8700 6740 8705
rect 6700 8670 6705 8700
rect 6705 8670 6735 8700
rect 6735 8670 6740 8700
rect 6700 8665 6740 8670
rect 6700 8630 6740 8635
rect 6700 8600 6705 8630
rect 6705 8600 6735 8630
rect 6735 8600 6740 8630
rect 6700 8595 6740 8600
rect 6700 8560 6740 8565
rect 6700 8530 6705 8560
rect 6705 8530 6735 8560
rect 6735 8530 6740 8560
rect 6700 8525 6740 8530
rect 6700 8495 6740 8500
rect 6700 8465 6705 8495
rect 6705 8465 6735 8495
rect 6735 8465 6740 8495
rect 6700 8460 6740 8465
rect 6700 8435 6740 8440
rect 6700 8405 6705 8435
rect 6705 8405 6735 8435
rect 6735 8405 6740 8435
rect 6700 8400 6740 8405
rect 6700 8370 6740 8375
rect 6700 8340 6705 8370
rect 6705 8340 6735 8370
rect 6735 8340 6740 8370
rect 6700 8335 6740 8340
rect 6700 8300 6740 8305
rect 6700 8270 6705 8300
rect 6705 8270 6735 8300
rect 6735 8270 6740 8300
rect 6700 8265 6740 8270
rect 6700 8230 6740 8235
rect 6700 8200 6705 8230
rect 6705 8200 6735 8230
rect 6735 8200 6740 8230
rect 6700 8195 6740 8200
rect 6700 8160 6740 8165
rect 6700 8130 6705 8160
rect 6705 8130 6735 8160
rect 6735 8130 6740 8160
rect 6700 8125 6740 8130
rect 7620 9635 7660 9640
rect 7620 9605 7625 9635
rect 7625 9605 7655 9635
rect 7655 9605 7660 9635
rect 7620 9600 7660 9605
rect 7620 9570 7660 9575
rect 7620 9540 7625 9570
rect 7625 9540 7655 9570
rect 7655 9540 7660 9570
rect 7620 9535 7660 9540
rect 7620 9500 7660 9505
rect 7620 9470 7625 9500
rect 7625 9470 7655 9500
rect 7655 9470 7660 9500
rect 7620 9465 7660 9470
rect 7620 9430 7660 9435
rect 7620 9400 7625 9430
rect 7625 9400 7655 9430
rect 7655 9400 7660 9430
rect 7620 9395 7660 9400
rect 7620 9360 7660 9365
rect 7620 9330 7625 9360
rect 7625 9330 7655 9360
rect 7655 9330 7660 9360
rect 7620 9325 7660 9330
rect 7620 9295 7660 9300
rect 7620 9265 7625 9295
rect 7625 9265 7655 9295
rect 7655 9265 7660 9295
rect 7620 9260 7660 9265
rect 7620 9235 7660 9240
rect 7620 9205 7625 9235
rect 7625 9205 7655 9235
rect 7655 9205 7660 9235
rect 7620 9200 7660 9205
rect 7620 9170 7660 9175
rect 7620 9140 7625 9170
rect 7625 9140 7655 9170
rect 7655 9140 7660 9170
rect 7620 9135 7660 9140
rect 7620 9100 7660 9105
rect 7620 9070 7625 9100
rect 7625 9070 7655 9100
rect 7655 9070 7660 9100
rect 7620 9065 7660 9070
rect 7620 9030 7660 9035
rect 7620 9000 7625 9030
rect 7625 9000 7655 9030
rect 7655 9000 7660 9030
rect 7620 8995 7660 9000
rect 7620 8960 7660 8965
rect 7620 8930 7625 8960
rect 7625 8930 7655 8960
rect 7655 8930 7660 8960
rect 7620 8925 7660 8930
rect 7620 8895 7660 8900
rect 7620 8865 7625 8895
rect 7625 8865 7655 8895
rect 7655 8865 7660 8895
rect 7620 8860 7660 8865
rect 7620 8835 7660 8840
rect 7620 8805 7625 8835
rect 7625 8805 7655 8835
rect 7655 8805 7660 8835
rect 7620 8800 7660 8805
rect 7620 8770 7660 8775
rect 7620 8740 7625 8770
rect 7625 8740 7655 8770
rect 7655 8740 7660 8770
rect 7620 8735 7660 8740
rect 7620 8700 7660 8705
rect 7620 8670 7625 8700
rect 7625 8670 7655 8700
rect 7655 8670 7660 8700
rect 7620 8665 7660 8670
rect 7620 8630 7660 8635
rect 7620 8600 7625 8630
rect 7625 8600 7655 8630
rect 7655 8600 7660 8630
rect 7620 8595 7660 8600
rect 7620 8560 7660 8565
rect 7620 8530 7625 8560
rect 7625 8530 7655 8560
rect 7655 8530 7660 8560
rect 7620 8525 7660 8530
rect 7620 8495 7660 8500
rect 7620 8465 7625 8495
rect 7625 8465 7655 8495
rect 7655 8465 7660 8495
rect 7620 8460 7660 8465
rect 7620 8435 7660 8440
rect 7620 8405 7625 8435
rect 7625 8405 7655 8435
rect 7655 8405 7660 8435
rect 7620 8400 7660 8405
rect 7620 8370 7660 8375
rect 7620 8340 7625 8370
rect 7625 8340 7655 8370
rect 7655 8340 7660 8370
rect 7620 8335 7660 8340
rect 7620 8300 7660 8305
rect 7620 8270 7625 8300
rect 7625 8270 7655 8300
rect 7655 8270 7660 8300
rect 7620 8265 7660 8270
rect 7620 8230 7660 8235
rect 7620 8200 7625 8230
rect 7625 8200 7655 8230
rect 7655 8200 7660 8230
rect 7620 8195 7660 8200
rect 7620 8160 7660 8165
rect 7620 8130 7625 8160
rect 7625 8130 7655 8160
rect 7655 8130 7660 8160
rect 7620 8125 7660 8130
rect 31305 9640 31340 9675
rect 31350 9640 31385 9675
rect 31395 9640 31430 9675
rect 31440 9640 31475 9675
rect 31485 9640 31520 9675
rect 31530 9640 31565 9675
rect 31575 9640 31610 9675
rect 31620 9640 31655 9675
rect 31665 9640 31700 9675
rect 31710 9640 31745 9675
rect 31755 9640 31790 9675
rect 31800 9640 31835 9675
rect 31845 9640 31880 9675
rect 31890 9640 31925 9675
rect 31935 9640 31970 9675
rect 31980 9640 32015 9675
rect 32025 9640 32060 9675
rect 32070 9640 32105 9675
rect 32115 9640 32150 9675
rect 32160 9640 32195 9675
rect 32205 9640 32240 9675
rect 32250 9640 32285 9675
rect 32295 9640 32330 9675
rect 32340 9640 32375 9675
rect 32385 9640 32420 9675
rect 32430 9640 32465 9675
rect 32475 9640 32510 9675
rect 32520 9640 32555 9675
rect 32565 9640 32600 9675
rect 32610 9640 32645 9675
rect 32655 9640 32690 9675
rect 32700 9640 32735 9675
rect 32745 9640 32780 9675
rect 32790 9640 32825 9675
rect 32835 9640 32870 9675
rect 31305 9595 31340 9630
rect 31350 9595 31385 9630
rect 31395 9595 31430 9630
rect 31440 9595 31475 9630
rect 31485 9595 31520 9630
rect 31530 9595 31565 9630
rect 31575 9595 31610 9630
rect 31620 9595 31655 9630
rect 31665 9595 31700 9630
rect 31710 9595 31745 9630
rect 31755 9595 31790 9630
rect 31800 9595 31835 9630
rect 31845 9595 31880 9630
rect 31890 9595 31925 9630
rect 31935 9595 31970 9630
rect 31980 9595 32015 9630
rect 32025 9595 32060 9630
rect 32070 9595 32105 9630
rect 32115 9595 32150 9630
rect 32160 9595 32195 9630
rect 32205 9595 32240 9630
rect 32250 9595 32285 9630
rect 32295 9595 32330 9630
rect 32340 9595 32375 9630
rect 32385 9595 32420 9630
rect 32430 9595 32465 9630
rect 32475 9595 32510 9630
rect 32520 9595 32555 9630
rect 32565 9595 32600 9630
rect 32610 9595 32645 9630
rect 32655 9595 32690 9630
rect 32700 9595 32735 9630
rect 32745 9595 32780 9630
rect 32790 9595 32825 9630
rect 32835 9595 32870 9630
rect 31305 9550 31340 9585
rect 31350 9550 31385 9585
rect 31395 9550 31430 9585
rect 31440 9550 31475 9585
rect 31485 9550 31520 9585
rect 31530 9550 31565 9585
rect 31575 9550 31610 9585
rect 31620 9550 31655 9585
rect 31665 9550 31700 9585
rect 31710 9550 31745 9585
rect 31755 9550 31790 9585
rect 31800 9550 31835 9585
rect 31845 9550 31880 9585
rect 31890 9550 31925 9585
rect 31935 9550 31970 9585
rect 31980 9550 32015 9585
rect 32025 9550 32060 9585
rect 32070 9550 32105 9585
rect 32115 9550 32150 9585
rect 32160 9550 32195 9585
rect 32205 9550 32240 9585
rect 32250 9550 32285 9585
rect 32295 9550 32330 9585
rect 32340 9550 32375 9585
rect 32385 9550 32420 9585
rect 32430 9550 32465 9585
rect 32475 9550 32510 9585
rect 32520 9550 32555 9585
rect 32565 9550 32600 9585
rect 32610 9550 32645 9585
rect 32655 9550 32690 9585
rect 32700 9550 32735 9585
rect 32745 9550 32780 9585
rect 32790 9550 32825 9585
rect 32835 9550 32870 9585
rect 31305 9505 31340 9540
rect 31350 9505 31385 9540
rect 31395 9505 31430 9540
rect 31440 9505 31475 9540
rect 31485 9505 31520 9540
rect 31530 9505 31565 9540
rect 31575 9505 31610 9540
rect 31620 9505 31655 9540
rect 31665 9505 31700 9540
rect 31710 9505 31745 9540
rect 31755 9505 31790 9540
rect 31800 9505 31835 9540
rect 31845 9505 31880 9540
rect 31890 9505 31925 9540
rect 31935 9505 31970 9540
rect 31980 9505 32015 9540
rect 32025 9505 32060 9540
rect 32070 9505 32105 9540
rect 32115 9505 32150 9540
rect 32160 9505 32195 9540
rect 32205 9505 32240 9540
rect 32250 9505 32285 9540
rect 32295 9505 32330 9540
rect 32340 9505 32375 9540
rect 32385 9505 32420 9540
rect 32430 9505 32465 9540
rect 32475 9505 32510 9540
rect 32520 9505 32555 9540
rect 32565 9505 32600 9540
rect 32610 9505 32645 9540
rect 32655 9505 32690 9540
rect 32700 9505 32735 9540
rect 32745 9505 32780 9540
rect 32790 9505 32825 9540
rect 32835 9505 32870 9540
rect 31305 9460 31340 9495
rect 31350 9460 31385 9495
rect 31395 9460 31430 9495
rect 31440 9460 31475 9495
rect 31485 9460 31520 9495
rect 31530 9460 31565 9495
rect 31575 9460 31610 9495
rect 31620 9460 31655 9495
rect 31665 9460 31700 9495
rect 31710 9460 31745 9495
rect 31755 9460 31790 9495
rect 31800 9460 31835 9495
rect 31845 9460 31880 9495
rect 31890 9460 31925 9495
rect 31935 9460 31970 9495
rect 31980 9460 32015 9495
rect 32025 9460 32060 9495
rect 32070 9460 32105 9495
rect 32115 9460 32150 9495
rect 32160 9460 32195 9495
rect 32205 9460 32240 9495
rect 32250 9460 32285 9495
rect 32295 9460 32330 9495
rect 32340 9460 32375 9495
rect 32385 9460 32420 9495
rect 32430 9460 32465 9495
rect 32475 9460 32510 9495
rect 32520 9460 32555 9495
rect 32565 9460 32600 9495
rect 32610 9460 32645 9495
rect 32655 9460 32690 9495
rect 32700 9460 32735 9495
rect 32745 9460 32780 9495
rect 32790 9460 32825 9495
rect 32835 9460 32870 9495
rect 31305 9415 31340 9450
rect 31350 9415 31385 9450
rect 31395 9415 31430 9450
rect 31440 9415 31475 9450
rect 31485 9415 31520 9450
rect 31530 9415 31565 9450
rect 31575 9415 31610 9450
rect 31620 9415 31655 9450
rect 31665 9415 31700 9450
rect 31710 9415 31745 9450
rect 31755 9415 31790 9450
rect 31800 9415 31835 9450
rect 31845 9415 31880 9450
rect 31890 9415 31925 9450
rect 31935 9415 31970 9450
rect 31980 9415 32015 9450
rect 32025 9415 32060 9450
rect 32070 9415 32105 9450
rect 32115 9415 32150 9450
rect 32160 9415 32195 9450
rect 32205 9415 32240 9450
rect 32250 9415 32285 9450
rect 32295 9415 32330 9450
rect 32340 9415 32375 9450
rect 32385 9415 32420 9450
rect 32430 9415 32465 9450
rect 32475 9415 32510 9450
rect 32520 9415 32555 9450
rect 32565 9415 32600 9450
rect 32610 9415 32645 9450
rect 32655 9415 32690 9450
rect 32700 9415 32735 9450
rect 32745 9415 32780 9450
rect 32790 9415 32825 9450
rect 32835 9415 32870 9450
rect 31305 9370 31340 9405
rect 31350 9370 31385 9405
rect 31395 9370 31430 9405
rect 31440 9370 31475 9405
rect 31485 9370 31520 9405
rect 31530 9370 31565 9405
rect 31575 9370 31610 9405
rect 31620 9370 31655 9405
rect 31665 9370 31700 9405
rect 31710 9370 31745 9405
rect 31755 9370 31790 9405
rect 31800 9370 31835 9405
rect 31845 9370 31880 9405
rect 31890 9370 31925 9405
rect 31935 9370 31970 9405
rect 31980 9370 32015 9405
rect 32025 9370 32060 9405
rect 32070 9370 32105 9405
rect 32115 9370 32150 9405
rect 32160 9370 32195 9405
rect 32205 9370 32240 9405
rect 32250 9370 32285 9405
rect 32295 9370 32330 9405
rect 32340 9370 32375 9405
rect 32385 9370 32420 9405
rect 32430 9370 32465 9405
rect 32475 9370 32510 9405
rect 32520 9370 32555 9405
rect 32565 9370 32600 9405
rect 32610 9370 32645 9405
rect 32655 9370 32690 9405
rect 32700 9370 32735 9405
rect 32745 9370 32780 9405
rect 32790 9370 32825 9405
rect 32835 9370 32870 9405
rect 31305 9325 31340 9360
rect 31350 9325 31385 9360
rect 31395 9325 31430 9360
rect 31440 9325 31475 9360
rect 31485 9325 31520 9360
rect 31530 9325 31565 9360
rect 31575 9325 31610 9360
rect 31620 9325 31655 9360
rect 31665 9325 31700 9360
rect 31710 9325 31745 9360
rect 31755 9325 31790 9360
rect 31800 9325 31835 9360
rect 31845 9325 31880 9360
rect 31890 9325 31925 9360
rect 31935 9325 31970 9360
rect 31980 9325 32015 9360
rect 32025 9325 32060 9360
rect 32070 9325 32105 9360
rect 32115 9325 32150 9360
rect 32160 9325 32195 9360
rect 32205 9325 32240 9360
rect 32250 9325 32285 9360
rect 32295 9325 32330 9360
rect 32340 9325 32375 9360
rect 32385 9325 32420 9360
rect 32430 9325 32465 9360
rect 32475 9325 32510 9360
rect 32520 9325 32555 9360
rect 32565 9325 32600 9360
rect 32610 9325 32645 9360
rect 32655 9325 32690 9360
rect 32700 9325 32735 9360
rect 32745 9325 32780 9360
rect 32790 9325 32825 9360
rect 32835 9325 32870 9360
rect 31305 9280 31340 9315
rect 31350 9280 31385 9315
rect 31395 9280 31430 9315
rect 31440 9280 31475 9315
rect 31485 9280 31520 9315
rect 31530 9280 31565 9315
rect 31575 9280 31610 9315
rect 31620 9280 31655 9315
rect 31665 9280 31700 9315
rect 31710 9280 31745 9315
rect 31755 9280 31790 9315
rect 31800 9280 31835 9315
rect 31845 9280 31880 9315
rect 31890 9280 31925 9315
rect 31935 9280 31970 9315
rect 31980 9280 32015 9315
rect 32025 9280 32060 9315
rect 32070 9280 32105 9315
rect 32115 9280 32150 9315
rect 32160 9280 32195 9315
rect 32205 9280 32240 9315
rect 32250 9280 32285 9315
rect 32295 9280 32330 9315
rect 32340 9280 32375 9315
rect 32385 9280 32420 9315
rect 32430 9280 32465 9315
rect 32475 9280 32510 9315
rect 32520 9280 32555 9315
rect 32565 9280 32600 9315
rect 32610 9280 32645 9315
rect 32655 9280 32690 9315
rect 32700 9280 32735 9315
rect 32745 9280 32780 9315
rect 32790 9280 32825 9315
rect 32835 9280 32870 9315
rect 31305 9235 31340 9270
rect 31350 9235 31385 9270
rect 31395 9235 31430 9270
rect 31440 9235 31475 9270
rect 31485 9235 31520 9270
rect 31530 9235 31565 9270
rect 31575 9235 31610 9270
rect 31620 9235 31655 9270
rect 31665 9235 31700 9270
rect 31710 9235 31745 9270
rect 31755 9235 31790 9270
rect 31800 9235 31835 9270
rect 31845 9235 31880 9270
rect 31890 9235 31925 9270
rect 31935 9235 31970 9270
rect 31980 9235 32015 9270
rect 32025 9235 32060 9270
rect 32070 9235 32105 9270
rect 32115 9235 32150 9270
rect 32160 9235 32195 9270
rect 32205 9235 32240 9270
rect 32250 9235 32285 9270
rect 32295 9235 32330 9270
rect 32340 9235 32375 9270
rect 32385 9235 32420 9270
rect 32430 9235 32465 9270
rect 32475 9235 32510 9270
rect 32520 9235 32555 9270
rect 32565 9235 32600 9270
rect 32610 9235 32645 9270
rect 32655 9235 32690 9270
rect 32700 9235 32735 9270
rect 32745 9235 32780 9270
rect 32790 9235 32825 9270
rect 32835 9235 32870 9270
rect 31305 9190 31340 9225
rect 31350 9190 31385 9225
rect 31395 9190 31430 9225
rect 31440 9190 31475 9225
rect 31485 9190 31520 9225
rect 31530 9190 31565 9225
rect 31575 9190 31610 9225
rect 31620 9190 31655 9225
rect 31665 9190 31700 9225
rect 31710 9190 31745 9225
rect 31755 9190 31790 9225
rect 31800 9190 31835 9225
rect 31845 9190 31880 9225
rect 31890 9190 31925 9225
rect 31935 9190 31970 9225
rect 31980 9190 32015 9225
rect 32025 9190 32060 9225
rect 32070 9190 32105 9225
rect 32115 9190 32150 9225
rect 32160 9190 32195 9225
rect 32205 9190 32240 9225
rect 32250 9190 32285 9225
rect 32295 9190 32330 9225
rect 32340 9190 32375 9225
rect 32385 9190 32420 9225
rect 32430 9190 32465 9225
rect 32475 9190 32510 9225
rect 32520 9190 32555 9225
rect 32565 9190 32600 9225
rect 32610 9190 32645 9225
rect 32655 9190 32690 9225
rect 32700 9190 32735 9225
rect 32745 9190 32780 9225
rect 32790 9190 32825 9225
rect 32835 9190 32870 9225
rect 31305 9145 31340 9180
rect 31350 9145 31385 9180
rect 31395 9145 31430 9180
rect 31440 9145 31475 9180
rect 31485 9145 31520 9180
rect 31530 9145 31565 9180
rect 31575 9145 31610 9180
rect 31620 9145 31655 9180
rect 31665 9145 31700 9180
rect 31710 9145 31745 9180
rect 31755 9145 31790 9180
rect 31800 9145 31835 9180
rect 31845 9145 31880 9180
rect 31890 9145 31925 9180
rect 31935 9145 31970 9180
rect 31980 9145 32015 9180
rect 32025 9145 32060 9180
rect 32070 9145 32105 9180
rect 32115 9145 32150 9180
rect 32160 9145 32195 9180
rect 32205 9145 32240 9180
rect 32250 9145 32285 9180
rect 32295 9145 32330 9180
rect 32340 9145 32375 9180
rect 32385 9145 32420 9180
rect 32430 9145 32465 9180
rect 32475 9145 32510 9180
rect 32520 9145 32555 9180
rect 32565 9145 32600 9180
rect 32610 9145 32645 9180
rect 32655 9145 32690 9180
rect 32700 9145 32735 9180
rect 32745 9145 32780 9180
rect 32790 9145 32825 9180
rect 32835 9145 32870 9180
rect 31305 9100 31340 9135
rect 31350 9100 31385 9135
rect 31395 9100 31430 9135
rect 31440 9100 31475 9135
rect 31485 9100 31520 9135
rect 31530 9100 31565 9135
rect 31575 9100 31610 9135
rect 31620 9100 31655 9135
rect 31665 9100 31700 9135
rect 31710 9100 31745 9135
rect 31755 9100 31790 9135
rect 31800 9100 31835 9135
rect 31845 9100 31880 9135
rect 31890 9100 31925 9135
rect 31935 9100 31970 9135
rect 31980 9100 32015 9135
rect 32025 9100 32060 9135
rect 32070 9100 32105 9135
rect 32115 9100 32150 9135
rect 32160 9100 32195 9135
rect 32205 9100 32240 9135
rect 32250 9100 32285 9135
rect 32295 9100 32330 9135
rect 32340 9100 32375 9135
rect 32385 9100 32420 9135
rect 32430 9100 32465 9135
rect 32475 9100 32510 9135
rect 32520 9100 32555 9135
rect 32565 9100 32600 9135
rect 32610 9100 32645 9135
rect 32655 9100 32690 9135
rect 32700 9100 32735 9135
rect 32745 9100 32780 9135
rect 32790 9100 32825 9135
rect 32835 9100 32870 9135
rect 31305 9055 31340 9090
rect 31350 9055 31385 9090
rect 31395 9055 31430 9090
rect 31440 9055 31475 9090
rect 31485 9055 31520 9090
rect 31530 9055 31565 9090
rect 31575 9055 31610 9090
rect 31620 9055 31655 9090
rect 31665 9055 31700 9090
rect 31710 9055 31745 9090
rect 31755 9055 31790 9090
rect 31800 9055 31835 9090
rect 31845 9055 31880 9090
rect 31890 9055 31925 9090
rect 31935 9055 31970 9090
rect 31980 9055 32015 9090
rect 32025 9055 32060 9090
rect 32070 9055 32105 9090
rect 32115 9055 32150 9090
rect 32160 9055 32195 9090
rect 32205 9055 32240 9090
rect 32250 9055 32285 9090
rect 32295 9055 32330 9090
rect 32340 9055 32375 9090
rect 32385 9055 32420 9090
rect 32430 9055 32465 9090
rect 32475 9055 32510 9090
rect 32520 9055 32555 9090
rect 32565 9055 32600 9090
rect 32610 9055 32645 9090
rect 32655 9055 32690 9090
rect 32700 9055 32735 9090
rect 32745 9055 32780 9090
rect 32790 9055 32825 9090
rect 32835 9055 32870 9090
rect 31305 9010 31340 9045
rect 31350 9010 31385 9045
rect 31395 9010 31430 9045
rect 31440 9010 31475 9045
rect 31485 9010 31520 9045
rect 31530 9010 31565 9045
rect 31575 9010 31610 9045
rect 31620 9010 31655 9045
rect 31665 9010 31700 9045
rect 31710 9010 31745 9045
rect 31755 9010 31790 9045
rect 31800 9010 31835 9045
rect 31845 9010 31880 9045
rect 31890 9010 31925 9045
rect 31935 9010 31970 9045
rect 31980 9010 32015 9045
rect 32025 9010 32060 9045
rect 32070 9010 32105 9045
rect 32115 9010 32150 9045
rect 32160 9010 32195 9045
rect 32205 9010 32240 9045
rect 32250 9010 32285 9045
rect 32295 9010 32330 9045
rect 32340 9010 32375 9045
rect 32385 9010 32420 9045
rect 32430 9010 32465 9045
rect 32475 9010 32510 9045
rect 32520 9010 32555 9045
rect 32565 9010 32600 9045
rect 32610 9010 32645 9045
rect 32655 9010 32690 9045
rect 32700 9010 32735 9045
rect 32745 9010 32780 9045
rect 32790 9010 32825 9045
rect 32835 9010 32870 9045
rect 31305 8965 31340 9000
rect 31350 8965 31385 9000
rect 31395 8965 31430 9000
rect 31440 8965 31475 9000
rect 31485 8965 31520 9000
rect 31530 8965 31565 9000
rect 31575 8965 31610 9000
rect 31620 8965 31655 9000
rect 31665 8965 31700 9000
rect 31710 8965 31745 9000
rect 31755 8965 31790 9000
rect 31800 8965 31835 9000
rect 31845 8965 31880 9000
rect 31890 8965 31925 9000
rect 31935 8965 31970 9000
rect 31980 8965 32015 9000
rect 32025 8965 32060 9000
rect 32070 8965 32105 9000
rect 32115 8965 32150 9000
rect 32160 8965 32195 9000
rect 32205 8965 32240 9000
rect 32250 8965 32285 9000
rect 32295 8965 32330 9000
rect 32340 8965 32375 9000
rect 32385 8965 32420 9000
rect 32430 8965 32465 9000
rect 32475 8965 32510 9000
rect 32520 8965 32555 9000
rect 32565 8965 32600 9000
rect 32610 8965 32645 9000
rect 32655 8965 32690 9000
rect 32700 8965 32735 9000
rect 32745 8965 32780 9000
rect 32790 8965 32825 9000
rect 32835 8965 32870 9000
rect -80 225 -40 230
rect -80 195 -75 225
rect -75 195 -45 225
rect -45 195 -40 225
rect -80 190 -40 195
rect -80 160 -40 165
rect -80 130 -75 160
rect -75 130 -45 160
rect -45 130 -40 160
rect -80 125 -40 130
rect -80 90 -40 95
rect -80 60 -75 90
rect -75 60 -45 90
rect -45 60 -40 90
rect -80 55 -40 60
rect -80 20 -40 25
rect -80 -10 -75 20
rect -75 -10 -45 20
rect -45 -10 -40 20
rect -80 -15 -40 -10
rect -80 -50 -40 -45
rect -80 -80 -75 -50
rect -75 -80 -45 -50
rect -45 -80 -40 -50
rect -80 -85 -40 -80
rect -80 -115 -40 -110
rect -80 -145 -75 -115
rect -75 -145 -45 -115
rect -45 -145 -40 -115
rect -80 -150 -40 -145
rect -80 -175 -40 -170
rect -80 -205 -75 -175
rect -75 -205 -45 -175
rect -45 -205 -40 -175
rect -80 -210 -40 -205
rect -80 -240 -40 -235
rect -80 -270 -75 -240
rect -75 -270 -45 -240
rect -45 -270 -40 -240
rect -80 -275 -40 -270
rect -80 -310 -40 -305
rect -80 -340 -75 -310
rect -75 -340 -45 -310
rect -45 -340 -40 -310
rect -80 -345 -40 -340
rect -80 -380 -40 -375
rect -80 -410 -75 -380
rect -75 -410 -45 -380
rect -45 -410 -40 -380
rect -80 -415 -40 -410
rect -80 -450 -40 -445
rect -80 -480 -75 -450
rect -75 -480 -45 -450
rect -45 -480 -40 -450
rect -80 -485 -40 -480
rect -80 -515 -40 -510
rect -80 -545 -75 -515
rect -75 -545 -45 -515
rect -45 -545 -40 -515
rect -80 -550 -40 -545
rect -80 -575 -40 -570
rect -80 -605 -75 -575
rect -75 -605 -45 -575
rect -45 -605 -40 -575
rect -80 -610 -40 -605
rect -80 -640 -40 -635
rect -80 -670 -75 -640
rect -75 -670 -45 -640
rect -45 -670 -40 -640
rect -80 -675 -40 -670
rect -80 -710 -40 -705
rect -80 -740 -75 -710
rect -75 -740 -45 -710
rect -45 -740 -40 -710
rect -80 -745 -40 -740
rect -80 -780 -40 -775
rect -80 -810 -75 -780
rect -75 -810 -45 -780
rect -45 -810 -40 -780
rect -80 -815 -40 -810
rect -80 -850 -40 -845
rect -80 -880 -75 -850
rect -75 -880 -45 -850
rect -45 -880 -40 -850
rect -80 -885 -40 -880
rect -80 -915 -40 -910
rect -80 -945 -75 -915
rect -75 -945 -45 -915
rect -45 -945 -40 -915
rect -80 -950 -40 -945
rect -80 -975 -40 -970
rect -80 -1005 -75 -975
rect -75 -1005 -45 -975
rect -45 -1005 -40 -975
rect -80 -1010 -40 -1005
rect -80 -1040 -40 -1035
rect -80 -1070 -75 -1040
rect -75 -1070 -45 -1040
rect -45 -1070 -40 -1040
rect -80 -1075 -40 -1070
rect -80 -1110 -40 -1105
rect -80 -1140 -75 -1110
rect -75 -1140 -45 -1110
rect -45 -1140 -40 -1110
rect -80 -1145 -40 -1140
rect -80 -1180 -40 -1175
rect -80 -1210 -75 -1180
rect -75 -1210 -45 -1180
rect -45 -1210 -40 -1180
rect -80 -1215 -40 -1210
rect -80 -1250 -40 -1245
rect -80 -1280 -75 -1250
rect -75 -1280 -45 -1250
rect -45 -1280 -40 -1250
rect -80 -1285 -40 -1280
rect -80 -1315 -40 -1310
rect -80 -1345 -75 -1315
rect -75 -1345 -45 -1315
rect -45 -1345 -40 -1315
rect -80 -1350 -40 -1345
rect 270 225 310 230
rect 270 195 275 225
rect 275 195 305 225
rect 305 195 310 225
rect 270 190 310 195
rect 270 160 310 165
rect 270 130 275 160
rect 275 130 305 160
rect 305 130 310 160
rect 270 125 310 130
rect 270 90 310 95
rect 270 60 275 90
rect 275 60 305 90
rect 305 60 310 90
rect 270 55 310 60
rect 270 20 310 25
rect 270 -10 275 20
rect 275 -10 305 20
rect 305 -10 310 20
rect 270 -15 310 -10
rect 270 -50 310 -45
rect 270 -80 275 -50
rect 275 -80 305 -50
rect 305 -80 310 -50
rect 270 -85 310 -80
rect 270 -115 310 -110
rect 270 -145 275 -115
rect 275 -145 305 -115
rect 305 -145 310 -115
rect 270 -150 310 -145
rect 270 -175 310 -170
rect 270 -205 275 -175
rect 275 -205 305 -175
rect 305 -205 310 -175
rect 270 -210 310 -205
rect 270 -240 310 -235
rect 270 -270 275 -240
rect 275 -270 305 -240
rect 305 -270 310 -240
rect 270 -275 310 -270
rect 270 -310 310 -305
rect 270 -340 275 -310
rect 275 -340 305 -310
rect 305 -340 310 -310
rect 270 -345 310 -340
rect 270 -380 310 -375
rect 270 -410 275 -380
rect 275 -410 305 -380
rect 305 -410 310 -380
rect 270 -415 310 -410
rect 270 -450 310 -445
rect 270 -480 275 -450
rect 275 -480 305 -450
rect 305 -480 310 -450
rect 270 -485 310 -480
rect 270 -515 310 -510
rect 270 -545 275 -515
rect 275 -545 305 -515
rect 305 -545 310 -515
rect 270 -550 310 -545
rect 270 -575 310 -570
rect 270 -605 275 -575
rect 275 -605 305 -575
rect 305 -605 310 -575
rect 270 -610 310 -605
rect 270 -640 310 -635
rect 270 -670 275 -640
rect 275 -670 305 -640
rect 305 -670 310 -640
rect 270 -675 310 -670
rect 270 -710 310 -705
rect 270 -740 275 -710
rect 275 -740 305 -710
rect 305 -740 310 -710
rect 270 -745 310 -740
rect 270 -780 310 -775
rect 270 -810 275 -780
rect 275 -810 305 -780
rect 305 -810 310 -780
rect 270 -815 310 -810
rect 270 -850 310 -845
rect 270 -880 275 -850
rect 275 -880 305 -850
rect 305 -880 310 -850
rect 270 -885 310 -880
rect 270 -915 310 -910
rect 270 -945 275 -915
rect 275 -945 305 -915
rect 305 -945 310 -915
rect 270 -950 310 -945
rect 270 -975 310 -970
rect 270 -1005 275 -975
rect 275 -1005 305 -975
rect 305 -1005 310 -975
rect 270 -1010 310 -1005
rect 270 -1040 310 -1035
rect 270 -1070 275 -1040
rect 275 -1070 305 -1040
rect 305 -1070 310 -1040
rect 270 -1075 310 -1070
rect 270 -1110 310 -1105
rect 270 -1140 275 -1110
rect 275 -1140 305 -1110
rect 305 -1140 310 -1110
rect 270 -1145 310 -1140
rect 270 -1180 310 -1175
rect 270 -1210 275 -1180
rect 275 -1210 305 -1180
rect 305 -1210 310 -1180
rect 270 -1215 310 -1210
rect 270 -1250 310 -1245
rect 270 -1280 275 -1250
rect 275 -1280 305 -1250
rect 305 -1280 310 -1250
rect 270 -1285 310 -1280
rect 270 -1315 310 -1310
rect 270 -1345 275 -1315
rect 275 -1345 305 -1315
rect 305 -1345 310 -1315
rect 270 -1350 310 -1345
rect 620 225 660 230
rect 620 195 625 225
rect 625 195 655 225
rect 655 195 660 225
rect 620 190 660 195
rect 620 160 660 165
rect 620 130 625 160
rect 625 130 655 160
rect 655 130 660 160
rect 620 125 660 130
rect 620 90 660 95
rect 620 60 625 90
rect 625 60 655 90
rect 655 60 660 90
rect 620 55 660 60
rect 620 20 660 25
rect 620 -10 625 20
rect 625 -10 655 20
rect 655 -10 660 20
rect 620 -15 660 -10
rect 620 -50 660 -45
rect 620 -80 625 -50
rect 625 -80 655 -50
rect 655 -80 660 -50
rect 620 -85 660 -80
rect 620 -115 660 -110
rect 620 -145 625 -115
rect 625 -145 655 -115
rect 655 -145 660 -115
rect 620 -150 660 -145
rect 620 -175 660 -170
rect 620 -205 625 -175
rect 625 -205 655 -175
rect 655 -205 660 -175
rect 620 -210 660 -205
rect 620 -240 660 -235
rect 620 -270 625 -240
rect 625 -270 655 -240
rect 655 -270 660 -240
rect 620 -275 660 -270
rect 620 -310 660 -305
rect 620 -340 625 -310
rect 625 -340 655 -310
rect 655 -340 660 -310
rect 620 -345 660 -340
rect 620 -380 660 -375
rect 620 -410 625 -380
rect 625 -410 655 -380
rect 655 -410 660 -380
rect 620 -415 660 -410
rect 620 -450 660 -445
rect 620 -480 625 -450
rect 625 -480 655 -450
rect 655 -480 660 -450
rect 620 -485 660 -480
rect 620 -515 660 -510
rect 620 -545 625 -515
rect 625 -545 655 -515
rect 655 -545 660 -515
rect 620 -550 660 -545
rect 620 -575 660 -570
rect 620 -605 625 -575
rect 625 -605 655 -575
rect 655 -605 660 -575
rect 620 -610 660 -605
rect 620 -640 660 -635
rect 620 -670 625 -640
rect 625 -670 655 -640
rect 655 -670 660 -640
rect 620 -675 660 -670
rect 620 -710 660 -705
rect 620 -740 625 -710
rect 625 -740 655 -710
rect 655 -740 660 -710
rect 620 -745 660 -740
rect 620 -780 660 -775
rect 620 -810 625 -780
rect 625 -810 655 -780
rect 655 -810 660 -780
rect 620 -815 660 -810
rect 620 -850 660 -845
rect 620 -880 625 -850
rect 625 -880 655 -850
rect 655 -880 660 -850
rect 620 -885 660 -880
rect 620 -915 660 -910
rect 620 -945 625 -915
rect 625 -945 655 -915
rect 655 -945 660 -915
rect 620 -950 660 -945
rect 620 -975 660 -970
rect 620 -1005 625 -975
rect 625 -1005 655 -975
rect 655 -1005 660 -975
rect 620 -1010 660 -1005
rect 620 -1040 660 -1035
rect 620 -1070 625 -1040
rect 625 -1070 655 -1040
rect 655 -1070 660 -1040
rect 620 -1075 660 -1070
rect 620 -1110 660 -1105
rect 620 -1140 625 -1110
rect 625 -1140 655 -1110
rect 655 -1140 660 -1110
rect 620 -1145 660 -1140
rect 620 -1180 660 -1175
rect 620 -1210 625 -1180
rect 625 -1210 655 -1180
rect 655 -1210 660 -1180
rect 620 -1215 660 -1210
rect 620 -1250 660 -1245
rect 620 -1280 625 -1250
rect 625 -1280 655 -1250
rect 655 -1280 660 -1250
rect 620 -1285 660 -1280
rect 620 -1315 660 -1310
rect 620 -1345 625 -1315
rect 625 -1345 655 -1315
rect 655 -1345 660 -1315
rect 620 -1350 660 -1345
rect 970 225 1010 230
rect 970 195 975 225
rect 975 195 1005 225
rect 1005 195 1010 225
rect 970 190 1010 195
rect 970 160 1010 165
rect 970 130 975 160
rect 975 130 1005 160
rect 1005 130 1010 160
rect 970 125 1010 130
rect 970 90 1010 95
rect 970 60 975 90
rect 975 60 1005 90
rect 1005 60 1010 90
rect 970 55 1010 60
rect 970 20 1010 25
rect 970 -10 975 20
rect 975 -10 1005 20
rect 1005 -10 1010 20
rect 970 -15 1010 -10
rect 970 -50 1010 -45
rect 970 -80 975 -50
rect 975 -80 1005 -50
rect 1005 -80 1010 -50
rect 970 -85 1010 -80
rect 970 -115 1010 -110
rect 970 -145 975 -115
rect 975 -145 1005 -115
rect 1005 -145 1010 -115
rect 970 -150 1010 -145
rect 970 -175 1010 -170
rect 970 -205 975 -175
rect 975 -205 1005 -175
rect 1005 -205 1010 -175
rect 970 -210 1010 -205
rect 970 -240 1010 -235
rect 970 -270 975 -240
rect 975 -270 1005 -240
rect 1005 -270 1010 -240
rect 970 -275 1010 -270
rect 970 -310 1010 -305
rect 970 -340 975 -310
rect 975 -340 1005 -310
rect 1005 -340 1010 -310
rect 970 -345 1010 -340
rect 970 -380 1010 -375
rect 970 -410 975 -380
rect 975 -410 1005 -380
rect 1005 -410 1010 -380
rect 970 -415 1010 -410
rect 970 -450 1010 -445
rect 970 -480 975 -450
rect 975 -480 1005 -450
rect 1005 -480 1010 -450
rect 970 -485 1010 -480
rect 970 -515 1010 -510
rect 970 -545 975 -515
rect 975 -545 1005 -515
rect 1005 -545 1010 -515
rect 970 -550 1010 -545
rect 970 -575 1010 -570
rect 970 -605 975 -575
rect 975 -605 1005 -575
rect 1005 -605 1010 -575
rect 970 -610 1010 -605
rect 970 -640 1010 -635
rect 970 -670 975 -640
rect 975 -670 1005 -640
rect 1005 -670 1010 -640
rect 970 -675 1010 -670
rect 970 -710 1010 -705
rect 970 -740 975 -710
rect 975 -740 1005 -710
rect 1005 -740 1010 -710
rect 970 -745 1010 -740
rect 970 -780 1010 -775
rect 970 -810 975 -780
rect 975 -810 1005 -780
rect 1005 -810 1010 -780
rect 970 -815 1010 -810
rect 970 -850 1010 -845
rect 970 -880 975 -850
rect 975 -880 1005 -850
rect 1005 -880 1010 -850
rect 970 -885 1010 -880
rect 970 -915 1010 -910
rect 970 -945 975 -915
rect 975 -945 1005 -915
rect 1005 -945 1010 -915
rect 970 -950 1010 -945
rect 970 -975 1010 -970
rect 970 -1005 975 -975
rect 975 -1005 1005 -975
rect 1005 -1005 1010 -975
rect 970 -1010 1010 -1005
rect 970 -1040 1010 -1035
rect 970 -1070 975 -1040
rect 975 -1070 1005 -1040
rect 1005 -1070 1010 -1040
rect 970 -1075 1010 -1070
rect 970 -1110 1010 -1105
rect 970 -1140 975 -1110
rect 975 -1140 1005 -1110
rect 1005 -1140 1010 -1110
rect 970 -1145 1010 -1140
rect 970 -1180 1010 -1175
rect 970 -1210 975 -1180
rect 975 -1210 1005 -1180
rect 1005 -1210 1010 -1180
rect 970 -1215 1010 -1210
rect 970 -1250 1010 -1245
rect 970 -1280 975 -1250
rect 975 -1280 1005 -1250
rect 1005 -1280 1010 -1250
rect 970 -1285 1010 -1280
rect 970 -1315 1010 -1310
rect 970 -1345 975 -1315
rect 975 -1345 1005 -1315
rect 1005 -1345 1010 -1315
rect 970 -1350 1010 -1345
rect 1320 225 1360 230
rect 1320 195 1325 225
rect 1325 195 1355 225
rect 1355 195 1360 225
rect 1320 190 1360 195
rect 1320 160 1360 165
rect 1320 130 1325 160
rect 1325 130 1355 160
rect 1355 130 1360 160
rect 1320 125 1360 130
rect 1320 90 1360 95
rect 1320 60 1325 90
rect 1325 60 1355 90
rect 1355 60 1360 90
rect 1320 55 1360 60
rect 1320 20 1360 25
rect 1320 -10 1325 20
rect 1325 -10 1355 20
rect 1355 -10 1360 20
rect 1320 -15 1360 -10
rect 1320 -50 1360 -45
rect 1320 -80 1325 -50
rect 1325 -80 1355 -50
rect 1355 -80 1360 -50
rect 1320 -85 1360 -80
rect 1320 -115 1360 -110
rect 1320 -145 1325 -115
rect 1325 -145 1355 -115
rect 1355 -145 1360 -115
rect 1320 -150 1360 -145
rect 1320 -175 1360 -170
rect 1320 -205 1325 -175
rect 1325 -205 1355 -175
rect 1355 -205 1360 -175
rect 1320 -210 1360 -205
rect 1320 -240 1360 -235
rect 1320 -270 1325 -240
rect 1325 -270 1355 -240
rect 1355 -270 1360 -240
rect 1320 -275 1360 -270
rect 1320 -310 1360 -305
rect 1320 -340 1325 -310
rect 1325 -340 1355 -310
rect 1355 -340 1360 -310
rect 1320 -345 1360 -340
rect 1320 -380 1360 -375
rect 1320 -410 1325 -380
rect 1325 -410 1355 -380
rect 1355 -410 1360 -380
rect 1320 -415 1360 -410
rect 1320 -450 1360 -445
rect 1320 -480 1325 -450
rect 1325 -480 1355 -450
rect 1355 -480 1360 -450
rect 1320 -485 1360 -480
rect 1320 -515 1360 -510
rect 1320 -545 1325 -515
rect 1325 -545 1355 -515
rect 1355 -545 1360 -515
rect 1320 -550 1360 -545
rect 1320 -575 1360 -570
rect 1320 -605 1325 -575
rect 1325 -605 1355 -575
rect 1355 -605 1360 -575
rect 1320 -610 1360 -605
rect 1320 -640 1360 -635
rect 1320 -670 1325 -640
rect 1325 -670 1355 -640
rect 1355 -670 1360 -640
rect 1320 -675 1360 -670
rect 1320 -710 1360 -705
rect 1320 -740 1325 -710
rect 1325 -740 1355 -710
rect 1355 -740 1360 -710
rect 1320 -745 1360 -740
rect 1320 -780 1360 -775
rect 1320 -810 1325 -780
rect 1325 -810 1355 -780
rect 1355 -810 1360 -780
rect 1320 -815 1360 -810
rect 1320 -850 1360 -845
rect 1320 -880 1325 -850
rect 1325 -880 1355 -850
rect 1355 -880 1360 -850
rect 1320 -885 1360 -880
rect 1320 -915 1360 -910
rect 1320 -945 1325 -915
rect 1325 -945 1355 -915
rect 1355 -945 1360 -915
rect 1320 -950 1360 -945
rect 1320 -975 1360 -970
rect 1320 -1005 1325 -975
rect 1325 -1005 1355 -975
rect 1355 -1005 1360 -975
rect 1320 -1010 1360 -1005
rect 1320 -1040 1360 -1035
rect 1320 -1070 1325 -1040
rect 1325 -1070 1355 -1040
rect 1355 -1070 1360 -1040
rect 1320 -1075 1360 -1070
rect 1320 -1110 1360 -1105
rect 1320 -1140 1325 -1110
rect 1325 -1140 1355 -1110
rect 1355 -1140 1360 -1110
rect 1320 -1145 1360 -1140
rect 1320 -1180 1360 -1175
rect 1320 -1210 1325 -1180
rect 1325 -1210 1355 -1180
rect 1355 -1210 1360 -1180
rect 1320 -1215 1360 -1210
rect 1320 -1250 1360 -1245
rect 1320 -1280 1325 -1250
rect 1325 -1280 1355 -1250
rect 1355 -1280 1360 -1250
rect 1320 -1285 1360 -1280
rect 1320 -1315 1360 -1310
rect 1320 -1345 1325 -1315
rect 1325 -1345 1355 -1315
rect 1355 -1345 1360 -1315
rect 1320 -1350 1360 -1345
rect 1670 225 1710 230
rect 1670 195 1675 225
rect 1675 195 1705 225
rect 1705 195 1710 225
rect 1670 190 1710 195
rect 1670 160 1710 165
rect 1670 130 1675 160
rect 1675 130 1705 160
rect 1705 130 1710 160
rect 1670 125 1710 130
rect 1670 90 1710 95
rect 1670 60 1675 90
rect 1675 60 1705 90
rect 1705 60 1710 90
rect 1670 55 1710 60
rect 1670 20 1710 25
rect 1670 -10 1675 20
rect 1675 -10 1705 20
rect 1705 -10 1710 20
rect 1670 -15 1710 -10
rect 1670 -50 1710 -45
rect 1670 -80 1675 -50
rect 1675 -80 1705 -50
rect 1705 -80 1710 -50
rect 1670 -85 1710 -80
rect 1670 -115 1710 -110
rect 1670 -145 1675 -115
rect 1675 -145 1705 -115
rect 1705 -145 1710 -115
rect 1670 -150 1710 -145
rect 1670 -175 1710 -170
rect 1670 -205 1675 -175
rect 1675 -205 1705 -175
rect 1705 -205 1710 -175
rect 1670 -210 1710 -205
rect 1670 -240 1710 -235
rect 1670 -270 1675 -240
rect 1675 -270 1705 -240
rect 1705 -270 1710 -240
rect 1670 -275 1710 -270
rect 1670 -310 1710 -305
rect 1670 -340 1675 -310
rect 1675 -340 1705 -310
rect 1705 -340 1710 -310
rect 1670 -345 1710 -340
rect 1670 -380 1710 -375
rect 1670 -410 1675 -380
rect 1675 -410 1705 -380
rect 1705 -410 1710 -380
rect 1670 -415 1710 -410
rect 1670 -450 1710 -445
rect 1670 -480 1675 -450
rect 1675 -480 1705 -450
rect 1705 -480 1710 -450
rect 1670 -485 1710 -480
rect 1670 -515 1710 -510
rect 1670 -545 1675 -515
rect 1675 -545 1705 -515
rect 1705 -545 1710 -515
rect 1670 -550 1710 -545
rect 1670 -575 1710 -570
rect 1670 -605 1675 -575
rect 1675 -605 1705 -575
rect 1705 -605 1710 -575
rect 1670 -610 1710 -605
rect 1670 -640 1710 -635
rect 1670 -670 1675 -640
rect 1675 -670 1705 -640
rect 1705 -670 1710 -640
rect 1670 -675 1710 -670
rect 1670 -710 1710 -705
rect 1670 -740 1675 -710
rect 1675 -740 1705 -710
rect 1705 -740 1710 -710
rect 1670 -745 1710 -740
rect 1670 -780 1710 -775
rect 1670 -810 1675 -780
rect 1675 -810 1705 -780
rect 1705 -810 1710 -780
rect 1670 -815 1710 -810
rect 1670 -850 1710 -845
rect 1670 -880 1675 -850
rect 1675 -880 1705 -850
rect 1705 -880 1710 -850
rect 1670 -885 1710 -880
rect 1670 -915 1710 -910
rect 1670 -945 1675 -915
rect 1675 -945 1705 -915
rect 1705 -945 1710 -915
rect 1670 -950 1710 -945
rect 1670 -975 1710 -970
rect 1670 -1005 1675 -975
rect 1675 -1005 1705 -975
rect 1705 -1005 1710 -975
rect 1670 -1010 1710 -1005
rect 1670 -1040 1710 -1035
rect 1670 -1070 1675 -1040
rect 1675 -1070 1705 -1040
rect 1705 -1070 1710 -1040
rect 1670 -1075 1710 -1070
rect 1670 -1110 1710 -1105
rect 1670 -1140 1675 -1110
rect 1675 -1140 1705 -1110
rect 1705 -1140 1710 -1110
rect 1670 -1145 1710 -1140
rect 1670 -1180 1710 -1175
rect 1670 -1210 1675 -1180
rect 1675 -1210 1705 -1180
rect 1705 -1210 1710 -1180
rect 1670 -1215 1710 -1210
rect 1670 -1250 1710 -1245
rect 1670 -1280 1675 -1250
rect 1675 -1280 1705 -1250
rect 1705 -1280 1710 -1250
rect 1670 -1285 1710 -1280
rect 1670 -1315 1710 -1310
rect 1670 -1345 1675 -1315
rect 1675 -1345 1705 -1315
rect 1705 -1345 1710 -1315
rect 1670 -1350 1710 -1345
rect 2020 225 2060 230
rect 2020 195 2025 225
rect 2025 195 2055 225
rect 2055 195 2060 225
rect 2020 190 2060 195
rect 2020 160 2060 165
rect 2020 130 2025 160
rect 2025 130 2055 160
rect 2055 130 2060 160
rect 2020 125 2060 130
rect 2020 90 2060 95
rect 2020 60 2025 90
rect 2025 60 2055 90
rect 2055 60 2060 90
rect 2020 55 2060 60
rect 2020 20 2060 25
rect 2020 -10 2025 20
rect 2025 -10 2055 20
rect 2055 -10 2060 20
rect 2020 -15 2060 -10
rect 2020 -50 2060 -45
rect 2020 -80 2025 -50
rect 2025 -80 2055 -50
rect 2055 -80 2060 -50
rect 2020 -85 2060 -80
rect 2020 -115 2060 -110
rect 2020 -145 2025 -115
rect 2025 -145 2055 -115
rect 2055 -145 2060 -115
rect 2020 -150 2060 -145
rect 2020 -175 2060 -170
rect 2020 -205 2025 -175
rect 2025 -205 2055 -175
rect 2055 -205 2060 -175
rect 2020 -210 2060 -205
rect 2020 -240 2060 -235
rect 2020 -270 2025 -240
rect 2025 -270 2055 -240
rect 2055 -270 2060 -240
rect 2020 -275 2060 -270
rect 2020 -310 2060 -305
rect 2020 -340 2025 -310
rect 2025 -340 2055 -310
rect 2055 -340 2060 -310
rect 2020 -345 2060 -340
rect 2020 -380 2060 -375
rect 2020 -410 2025 -380
rect 2025 -410 2055 -380
rect 2055 -410 2060 -380
rect 2020 -415 2060 -410
rect 2020 -450 2060 -445
rect 2020 -480 2025 -450
rect 2025 -480 2055 -450
rect 2055 -480 2060 -450
rect 2020 -485 2060 -480
rect 2020 -515 2060 -510
rect 2020 -545 2025 -515
rect 2025 -545 2055 -515
rect 2055 -545 2060 -515
rect 2020 -550 2060 -545
rect 2020 -575 2060 -570
rect 2020 -605 2025 -575
rect 2025 -605 2055 -575
rect 2055 -605 2060 -575
rect 2020 -610 2060 -605
rect 2020 -640 2060 -635
rect 2020 -670 2025 -640
rect 2025 -670 2055 -640
rect 2055 -670 2060 -640
rect 2020 -675 2060 -670
rect 2020 -710 2060 -705
rect 2020 -740 2025 -710
rect 2025 -740 2055 -710
rect 2055 -740 2060 -710
rect 2020 -745 2060 -740
rect 2020 -780 2060 -775
rect 2020 -810 2025 -780
rect 2025 -810 2055 -780
rect 2055 -810 2060 -780
rect 2020 -815 2060 -810
rect 2020 -850 2060 -845
rect 2020 -880 2025 -850
rect 2025 -880 2055 -850
rect 2055 -880 2060 -850
rect 2020 -885 2060 -880
rect 2020 -915 2060 -910
rect 2020 -945 2025 -915
rect 2025 -945 2055 -915
rect 2055 -945 2060 -915
rect 2020 -950 2060 -945
rect 2020 -975 2060 -970
rect 2020 -1005 2025 -975
rect 2025 -1005 2055 -975
rect 2055 -1005 2060 -975
rect 2020 -1010 2060 -1005
rect 2020 -1040 2060 -1035
rect 2020 -1070 2025 -1040
rect 2025 -1070 2055 -1040
rect 2055 -1070 2060 -1040
rect 2020 -1075 2060 -1070
rect 2020 -1110 2060 -1105
rect 2020 -1140 2025 -1110
rect 2025 -1140 2055 -1110
rect 2055 -1140 2060 -1110
rect 2020 -1145 2060 -1140
rect 2020 -1180 2060 -1175
rect 2020 -1210 2025 -1180
rect 2025 -1210 2055 -1180
rect 2055 -1210 2060 -1180
rect 2020 -1215 2060 -1210
rect 2020 -1250 2060 -1245
rect 2020 -1280 2025 -1250
rect 2025 -1280 2055 -1250
rect 2055 -1280 2060 -1250
rect 2020 -1285 2060 -1280
rect 2020 -1315 2060 -1310
rect 2020 -1345 2025 -1315
rect 2025 -1345 2055 -1315
rect 2055 -1345 2060 -1315
rect 2020 -1350 2060 -1345
rect 2370 225 2410 230
rect 2370 195 2375 225
rect 2375 195 2405 225
rect 2405 195 2410 225
rect 2370 190 2410 195
rect 2370 160 2410 165
rect 2370 130 2375 160
rect 2375 130 2405 160
rect 2405 130 2410 160
rect 2370 125 2410 130
rect 2370 90 2410 95
rect 2370 60 2375 90
rect 2375 60 2405 90
rect 2405 60 2410 90
rect 2370 55 2410 60
rect 2370 20 2410 25
rect 2370 -10 2375 20
rect 2375 -10 2405 20
rect 2405 -10 2410 20
rect 2370 -15 2410 -10
rect 2370 -50 2410 -45
rect 2370 -80 2375 -50
rect 2375 -80 2405 -50
rect 2405 -80 2410 -50
rect 2370 -85 2410 -80
rect 2370 -115 2410 -110
rect 2370 -145 2375 -115
rect 2375 -145 2405 -115
rect 2405 -145 2410 -115
rect 2370 -150 2410 -145
rect 2370 -175 2410 -170
rect 2370 -205 2375 -175
rect 2375 -205 2405 -175
rect 2405 -205 2410 -175
rect 2370 -210 2410 -205
rect 2370 -240 2410 -235
rect 2370 -270 2375 -240
rect 2375 -270 2405 -240
rect 2405 -270 2410 -240
rect 2370 -275 2410 -270
rect 2370 -310 2410 -305
rect 2370 -340 2375 -310
rect 2375 -340 2405 -310
rect 2405 -340 2410 -310
rect 2370 -345 2410 -340
rect 2370 -380 2410 -375
rect 2370 -410 2375 -380
rect 2375 -410 2405 -380
rect 2405 -410 2410 -380
rect 2370 -415 2410 -410
rect 2370 -450 2410 -445
rect 2370 -480 2375 -450
rect 2375 -480 2405 -450
rect 2405 -480 2410 -450
rect 2370 -485 2410 -480
rect 2370 -515 2410 -510
rect 2370 -545 2375 -515
rect 2375 -545 2405 -515
rect 2405 -545 2410 -515
rect 2370 -550 2410 -545
rect 2370 -575 2410 -570
rect 2370 -605 2375 -575
rect 2375 -605 2405 -575
rect 2405 -605 2410 -575
rect 2370 -610 2410 -605
rect 2370 -640 2410 -635
rect 2370 -670 2375 -640
rect 2375 -670 2405 -640
rect 2405 -670 2410 -640
rect 2370 -675 2410 -670
rect 2370 -710 2410 -705
rect 2370 -740 2375 -710
rect 2375 -740 2405 -710
rect 2405 -740 2410 -710
rect 2370 -745 2410 -740
rect 2370 -780 2410 -775
rect 2370 -810 2375 -780
rect 2375 -810 2405 -780
rect 2405 -810 2410 -780
rect 2370 -815 2410 -810
rect 2370 -850 2410 -845
rect 2370 -880 2375 -850
rect 2375 -880 2405 -850
rect 2405 -880 2410 -850
rect 2370 -885 2410 -880
rect 2370 -915 2410 -910
rect 2370 -945 2375 -915
rect 2375 -945 2405 -915
rect 2405 -945 2410 -915
rect 2370 -950 2410 -945
rect 2370 -975 2410 -970
rect 2370 -1005 2375 -975
rect 2375 -1005 2405 -975
rect 2405 -1005 2410 -975
rect 2370 -1010 2410 -1005
rect 2370 -1040 2410 -1035
rect 2370 -1070 2375 -1040
rect 2375 -1070 2405 -1040
rect 2405 -1070 2410 -1040
rect 2370 -1075 2410 -1070
rect 2370 -1110 2410 -1105
rect 2370 -1140 2375 -1110
rect 2375 -1140 2405 -1110
rect 2405 -1140 2410 -1110
rect 2370 -1145 2410 -1140
rect 2370 -1180 2410 -1175
rect 2370 -1210 2375 -1180
rect 2375 -1210 2405 -1180
rect 2405 -1210 2410 -1180
rect 2370 -1215 2410 -1210
rect 2370 -1250 2410 -1245
rect 2370 -1280 2375 -1250
rect 2375 -1280 2405 -1250
rect 2405 -1280 2410 -1250
rect 2370 -1285 2410 -1280
rect 2370 -1315 2410 -1310
rect 2370 -1345 2375 -1315
rect 2375 -1345 2405 -1315
rect 2405 -1345 2410 -1315
rect 2370 -1350 2410 -1345
rect 2720 225 2760 230
rect 2720 195 2725 225
rect 2725 195 2755 225
rect 2755 195 2760 225
rect 2720 190 2760 195
rect 2720 160 2760 165
rect 2720 130 2725 160
rect 2725 130 2755 160
rect 2755 130 2760 160
rect 2720 125 2760 130
rect 2720 90 2760 95
rect 2720 60 2725 90
rect 2725 60 2755 90
rect 2755 60 2760 90
rect 2720 55 2760 60
rect 2720 20 2760 25
rect 2720 -10 2725 20
rect 2725 -10 2755 20
rect 2755 -10 2760 20
rect 2720 -15 2760 -10
rect 2720 -50 2760 -45
rect 2720 -80 2725 -50
rect 2725 -80 2755 -50
rect 2755 -80 2760 -50
rect 2720 -85 2760 -80
rect 2720 -115 2760 -110
rect 2720 -145 2725 -115
rect 2725 -145 2755 -115
rect 2755 -145 2760 -115
rect 2720 -150 2760 -145
rect 2720 -175 2760 -170
rect 2720 -205 2725 -175
rect 2725 -205 2755 -175
rect 2755 -205 2760 -175
rect 2720 -210 2760 -205
rect 2720 -240 2760 -235
rect 2720 -270 2725 -240
rect 2725 -270 2755 -240
rect 2755 -270 2760 -240
rect 2720 -275 2760 -270
rect 2720 -310 2760 -305
rect 2720 -340 2725 -310
rect 2725 -340 2755 -310
rect 2755 -340 2760 -310
rect 2720 -345 2760 -340
rect 2720 -380 2760 -375
rect 2720 -410 2725 -380
rect 2725 -410 2755 -380
rect 2755 -410 2760 -380
rect 2720 -415 2760 -410
rect 2720 -450 2760 -445
rect 2720 -480 2725 -450
rect 2725 -480 2755 -450
rect 2755 -480 2760 -450
rect 2720 -485 2760 -480
rect 2720 -515 2760 -510
rect 2720 -545 2725 -515
rect 2725 -545 2755 -515
rect 2755 -545 2760 -515
rect 2720 -550 2760 -545
rect 2720 -575 2760 -570
rect 2720 -605 2725 -575
rect 2725 -605 2755 -575
rect 2755 -605 2760 -575
rect 2720 -610 2760 -605
rect 2720 -640 2760 -635
rect 2720 -670 2725 -640
rect 2725 -670 2755 -640
rect 2755 -670 2760 -640
rect 2720 -675 2760 -670
rect 2720 -710 2760 -705
rect 2720 -740 2725 -710
rect 2725 -740 2755 -710
rect 2755 -740 2760 -710
rect 2720 -745 2760 -740
rect 2720 -780 2760 -775
rect 2720 -810 2725 -780
rect 2725 -810 2755 -780
rect 2755 -810 2760 -780
rect 2720 -815 2760 -810
rect 2720 -850 2760 -845
rect 2720 -880 2725 -850
rect 2725 -880 2755 -850
rect 2755 -880 2760 -850
rect 2720 -885 2760 -880
rect 2720 -915 2760 -910
rect 2720 -945 2725 -915
rect 2725 -945 2755 -915
rect 2755 -945 2760 -915
rect 2720 -950 2760 -945
rect 2720 -975 2760 -970
rect 2720 -1005 2725 -975
rect 2725 -1005 2755 -975
rect 2755 -1005 2760 -975
rect 2720 -1010 2760 -1005
rect 2720 -1040 2760 -1035
rect 2720 -1070 2725 -1040
rect 2725 -1070 2755 -1040
rect 2755 -1070 2760 -1040
rect 2720 -1075 2760 -1070
rect 2720 -1110 2760 -1105
rect 2720 -1140 2725 -1110
rect 2725 -1140 2755 -1110
rect 2755 -1140 2760 -1110
rect 2720 -1145 2760 -1140
rect 2720 -1180 2760 -1175
rect 2720 -1210 2725 -1180
rect 2725 -1210 2755 -1180
rect 2755 -1210 2760 -1180
rect 2720 -1215 2760 -1210
rect 2720 -1250 2760 -1245
rect 2720 -1280 2725 -1250
rect 2725 -1280 2755 -1250
rect 2755 -1280 2760 -1250
rect 2720 -1285 2760 -1280
rect 2720 -1315 2760 -1310
rect 2720 -1345 2725 -1315
rect 2725 -1345 2755 -1315
rect 2755 -1345 2760 -1315
rect 2720 -1350 2760 -1345
rect 3070 225 3110 230
rect 3070 195 3075 225
rect 3075 195 3105 225
rect 3105 195 3110 225
rect 3070 190 3110 195
rect 3070 160 3110 165
rect 3070 130 3075 160
rect 3075 130 3105 160
rect 3105 130 3110 160
rect 3070 125 3110 130
rect 3070 90 3110 95
rect 3070 60 3075 90
rect 3075 60 3105 90
rect 3105 60 3110 90
rect 3070 55 3110 60
rect 3070 20 3110 25
rect 3070 -10 3075 20
rect 3075 -10 3105 20
rect 3105 -10 3110 20
rect 3070 -15 3110 -10
rect 3070 -50 3110 -45
rect 3070 -80 3075 -50
rect 3075 -80 3105 -50
rect 3105 -80 3110 -50
rect 3070 -85 3110 -80
rect 3070 -115 3110 -110
rect 3070 -145 3075 -115
rect 3075 -145 3105 -115
rect 3105 -145 3110 -115
rect 3070 -150 3110 -145
rect 3070 -175 3110 -170
rect 3070 -205 3075 -175
rect 3075 -205 3105 -175
rect 3105 -205 3110 -175
rect 3070 -210 3110 -205
rect 3070 -240 3110 -235
rect 3070 -270 3075 -240
rect 3075 -270 3105 -240
rect 3105 -270 3110 -240
rect 3070 -275 3110 -270
rect 3070 -310 3110 -305
rect 3070 -340 3075 -310
rect 3075 -340 3105 -310
rect 3105 -340 3110 -310
rect 3070 -345 3110 -340
rect 3070 -380 3110 -375
rect 3070 -410 3075 -380
rect 3075 -410 3105 -380
rect 3105 -410 3110 -380
rect 3070 -415 3110 -410
rect 3070 -450 3110 -445
rect 3070 -480 3075 -450
rect 3075 -480 3105 -450
rect 3105 -480 3110 -450
rect 3070 -485 3110 -480
rect 3070 -515 3110 -510
rect 3070 -545 3075 -515
rect 3075 -545 3105 -515
rect 3105 -545 3110 -515
rect 3070 -550 3110 -545
rect 3070 -575 3110 -570
rect 3070 -605 3075 -575
rect 3075 -605 3105 -575
rect 3105 -605 3110 -575
rect 3070 -610 3110 -605
rect 3070 -640 3110 -635
rect 3070 -670 3075 -640
rect 3075 -670 3105 -640
rect 3105 -670 3110 -640
rect 3070 -675 3110 -670
rect 3070 -710 3110 -705
rect 3070 -740 3075 -710
rect 3075 -740 3105 -710
rect 3105 -740 3110 -710
rect 3070 -745 3110 -740
rect 3070 -780 3110 -775
rect 3070 -810 3075 -780
rect 3075 -810 3105 -780
rect 3105 -810 3110 -780
rect 3070 -815 3110 -810
rect 3070 -850 3110 -845
rect 3070 -880 3075 -850
rect 3075 -880 3105 -850
rect 3105 -880 3110 -850
rect 3070 -885 3110 -880
rect 3070 -915 3110 -910
rect 3070 -945 3075 -915
rect 3075 -945 3105 -915
rect 3105 -945 3110 -915
rect 3070 -950 3110 -945
rect 3070 -975 3110 -970
rect 3070 -1005 3075 -975
rect 3075 -1005 3105 -975
rect 3105 -1005 3110 -975
rect 3070 -1010 3110 -1005
rect 3070 -1040 3110 -1035
rect 3070 -1070 3075 -1040
rect 3075 -1070 3105 -1040
rect 3105 -1070 3110 -1040
rect 3070 -1075 3110 -1070
rect 3070 -1110 3110 -1105
rect 3070 -1140 3075 -1110
rect 3075 -1140 3105 -1110
rect 3105 -1140 3110 -1110
rect 3070 -1145 3110 -1140
rect 3070 -1180 3110 -1175
rect 3070 -1210 3075 -1180
rect 3075 -1210 3105 -1180
rect 3105 -1210 3110 -1180
rect 3070 -1215 3110 -1210
rect 3070 -1250 3110 -1245
rect 3070 -1280 3075 -1250
rect 3075 -1280 3105 -1250
rect 3105 -1280 3110 -1250
rect 3070 -1285 3110 -1280
rect 3070 -1315 3110 -1310
rect 3070 -1345 3075 -1315
rect 3075 -1345 3105 -1315
rect 3105 -1345 3110 -1315
rect 3070 -1350 3110 -1345
rect 3420 225 3460 230
rect 3420 195 3425 225
rect 3425 195 3455 225
rect 3455 195 3460 225
rect 3420 190 3460 195
rect 3420 160 3460 165
rect 3420 130 3425 160
rect 3425 130 3455 160
rect 3455 130 3460 160
rect 3420 125 3460 130
rect 3420 90 3460 95
rect 3420 60 3425 90
rect 3425 60 3455 90
rect 3455 60 3460 90
rect 3420 55 3460 60
rect 3420 20 3460 25
rect 3420 -10 3425 20
rect 3425 -10 3455 20
rect 3455 -10 3460 20
rect 3420 -15 3460 -10
rect 3420 -50 3460 -45
rect 3420 -80 3425 -50
rect 3425 -80 3455 -50
rect 3455 -80 3460 -50
rect 3420 -85 3460 -80
rect 3420 -115 3460 -110
rect 3420 -145 3425 -115
rect 3425 -145 3455 -115
rect 3455 -145 3460 -115
rect 3420 -150 3460 -145
rect 3420 -175 3460 -170
rect 3420 -205 3425 -175
rect 3425 -205 3455 -175
rect 3455 -205 3460 -175
rect 3420 -210 3460 -205
rect 3420 -240 3460 -235
rect 3420 -270 3425 -240
rect 3425 -270 3455 -240
rect 3455 -270 3460 -240
rect 3420 -275 3460 -270
rect 3420 -310 3460 -305
rect 3420 -340 3425 -310
rect 3425 -340 3455 -310
rect 3455 -340 3460 -310
rect 3420 -345 3460 -340
rect 3420 -380 3460 -375
rect 3420 -410 3425 -380
rect 3425 -410 3455 -380
rect 3455 -410 3460 -380
rect 3420 -415 3460 -410
rect 3420 -450 3460 -445
rect 3420 -480 3425 -450
rect 3425 -480 3455 -450
rect 3455 -480 3460 -450
rect 3420 -485 3460 -480
rect 3420 -515 3460 -510
rect 3420 -545 3425 -515
rect 3425 -545 3455 -515
rect 3455 -545 3460 -515
rect 3420 -550 3460 -545
rect 3420 -575 3460 -570
rect 3420 -605 3425 -575
rect 3425 -605 3455 -575
rect 3455 -605 3460 -575
rect 3420 -610 3460 -605
rect 3420 -640 3460 -635
rect 3420 -670 3425 -640
rect 3425 -670 3455 -640
rect 3455 -670 3460 -640
rect 3420 -675 3460 -670
rect 3420 -710 3460 -705
rect 3420 -740 3425 -710
rect 3425 -740 3455 -710
rect 3455 -740 3460 -710
rect 3420 -745 3460 -740
rect 3420 -780 3460 -775
rect 3420 -810 3425 -780
rect 3425 -810 3455 -780
rect 3455 -810 3460 -780
rect 3420 -815 3460 -810
rect 3420 -850 3460 -845
rect 3420 -880 3425 -850
rect 3425 -880 3455 -850
rect 3455 -880 3460 -850
rect 3420 -885 3460 -880
rect 3420 -915 3460 -910
rect 3420 -945 3425 -915
rect 3425 -945 3455 -915
rect 3455 -945 3460 -915
rect 3420 -950 3460 -945
rect 3420 -975 3460 -970
rect 3420 -1005 3425 -975
rect 3425 -1005 3455 -975
rect 3455 -1005 3460 -975
rect 3420 -1010 3460 -1005
rect 3420 -1040 3460 -1035
rect 3420 -1070 3425 -1040
rect 3425 -1070 3455 -1040
rect 3455 -1070 3460 -1040
rect 3420 -1075 3460 -1070
rect 3420 -1110 3460 -1105
rect 3420 -1140 3425 -1110
rect 3425 -1140 3455 -1110
rect 3455 -1140 3460 -1110
rect 3420 -1145 3460 -1140
rect 3420 -1180 3460 -1175
rect 3420 -1210 3425 -1180
rect 3425 -1210 3455 -1180
rect 3455 -1210 3460 -1180
rect 3420 -1215 3460 -1210
rect 3420 -1250 3460 -1245
rect 3420 -1280 3425 -1250
rect 3425 -1280 3455 -1250
rect 3455 -1280 3460 -1250
rect 3420 -1285 3460 -1280
rect 3420 -1315 3460 -1310
rect 3420 -1345 3425 -1315
rect 3425 -1345 3455 -1315
rect 3455 -1345 3460 -1315
rect 3420 -1350 3460 -1345
rect 3770 225 3810 230
rect 3770 195 3775 225
rect 3775 195 3805 225
rect 3805 195 3810 225
rect 3770 190 3810 195
rect 3770 160 3810 165
rect 3770 130 3775 160
rect 3775 130 3805 160
rect 3805 130 3810 160
rect 3770 125 3810 130
rect 3770 90 3810 95
rect 3770 60 3775 90
rect 3775 60 3805 90
rect 3805 60 3810 90
rect 3770 55 3810 60
rect 3770 20 3810 25
rect 3770 -10 3775 20
rect 3775 -10 3805 20
rect 3805 -10 3810 20
rect 3770 -15 3810 -10
rect 3770 -50 3810 -45
rect 3770 -80 3775 -50
rect 3775 -80 3805 -50
rect 3805 -80 3810 -50
rect 3770 -85 3810 -80
rect 3770 -115 3810 -110
rect 3770 -145 3775 -115
rect 3775 -145 3805 -115
rect 3805 -145 3810 -115
rect 3770 -150 3810 -145
rect 3770 -175 3810 -170
rect 3770 -205 3775 -175
rect 3775 -205 3805 -175
rect 3805 -205 3810 -175
rect 3770 -210 3810 -205
rect 3770 -240 3810 -235
rect 3770 -270 3775 -240
rect 3775 -270 3805 -240
rect 3805 -270 3810 -240
rect 3770 -275 3810 -270
rect 3770 -310 3810 -305
rect 3770 -340 3775 -310
rect 3775 -340 3805 -310
rect 3805 -340 3810 -310
rect 3770 -345 3810 -340
rect 3770 -380 3810 -375
rect 3770 -410 3775 -380
rect 3775 -410 3805 -380
rect 3805 -410 3810 -380
rect 3770 -415 3810 -410
rect 3770 -450 3810 -445
rect 3770 -480 3775 -450
rect 3775 -480 3805 -450
rect 3805 -480 3810 -450
rect 3770 -485 3810 -480
rect 3770 -515 3810 -510
rect 3770 -545 3775 -515
rect 3775 -545 3805 -515
rect 3805 -545 3810 -515
rect 3770 -550 3810 -545
rect 3770 -575 3810 -570
rect 3770 -605 3775 -575
rect 3775 -605 3805 -575
rect 3805 -605 3810 -575
rect 3770 -610 3810 -605
rect 3770 -640 3810 -635
rect 3770 -670 3775 -640
rect 3775 -670 3805 -640
rect 3805 -670 3810 -640
rect 3770 -675 3810 -670
rect 3770 -710 3810 -705
rect 3770 -740 3775 -710
rect 3775 -740 3805 -710
rect 3805 -740 3810 -710
rect 3770 -745 3810 -740
rect 3770 -780 3810 -775
rect 3770 -810 3775 -780
rect 3775 -810 3805 -780
rect 3805 -810 3810 -780
rect 3770 -815 3810 -810
rect 3770 -850 3810 -845
rect 3770 -880 3775 -850
rect 3775 -880 3805 -850
rect 3805 -880 3810 -850
rect 3770 -885 3810 -880
rect 3770 -915 3810 -910
rect 3770 -945 3775 -915
rect 3775 -945 3805 -915
rect 3805 -945 3810 -915
rect 3770 -950 3810 -945
rect 3770 -975 3810 -970
rect 3770 -1005 3775 -975
rect 3775 -1005 3805 -975
rect 3805 -1005 3810 -975
rect 3770 -1010 3810 -1005
rect 3770 -1040 3810 -1035
rect 3770 -1070 3775 -1040
rect 3775 -1070 3805 -1040
rect 3805 -1070 3810 -1040
rect 3770 -1075 3810 -1070
rect 3770 -1110 3810 -1105
rect 3770 -1140 3775 -1110
rect 3775 -1140 3805 -1110
rect 3805 -1140 3810 -1110
rect 3770 -1145 3810 -1140
rect 3770 -1180 3810 -1175
rect 3770 -1210 3775 -1180
rect 3775 -1210 3805 -1180
rect 3805 -1210 3810 -1180
rect 3770 -1215 3810 -1210
rect 3770 -1250 3810 -1245
rect 3770 -1280 3775 -1250
rect 3775 -1280 3805 -1250
rect 3805 -1280 3810 -1250
rect 3770 -1285 3810 -1280
rect 3770 -1315 3810 -1310
rect 3770 -1345 3775 -1315
rect 3775 -1345 3805 -1315
rect 3805 -1345 3810 -1315
rect 3770 -1350 3810 -1345
rect 4120 225 4160 230
rect 4120 195 4125 225
rect 4125 195 4155 225
rect 4155 195 4160 225
rect 4120 190 4160 195
rect 4120 160 4160 165
rect 4120 130 4125 160
rect 4125 130 4155 160
rect 4155 130 4160 160
rect 4120 125 4160 130
rect 4120 90 4160 95
rect 4120 60 4125 90
rect 4125 60 4155 90
rect 4155 60 4160 90
rect 4120 55 4160 60
rect 4120 20 4160 25
rect 4120 -10 4125 20
rect 4125 -10 4155 20
rect 4155 -10 4160 20
rect 4120 -15 4160 -10
rect 4120 -50 4160 -45
rect 4120 -80 4125 -50
rect 4125 -80 4155 -50
rect 4155 -80 4160 -50
rect 4120 -85 4160 -80
rect 4120 -115 4160 -110
rect 4120 -145 4125 -115
rect 4125 -145 4155 -115
rect 4155 -145 4160 -115
rect 4120 -150 4160 -145
rect 4120 -175 4160 -170
rect 4120 -205 4125 -175
rect 4125 -205 4155 -175
rect 4155 -205 4160 -175
rect 4120 -210 4160 -205
rect 4120 -240 4160 -235
rect 4120 -270 4125 -240
rect 4125 -270 4155 -240
rect 4155 -270 4160 -240
rect 4120 -275 4160 -270
rect 4120 -310 4160 -305
rect 4120 -340 4125 -310
rect 4125 -340 4155 -310
rect 4155 -340 4160 -310
rect 4120 -345 4160 -340
rect 4120 -380 4160 -375
rect 4120 -410 4125 -380
rect 4125 -410 4155 -380
rect 4155 -410 4160 -380
rect 4120 -415 4160 -410
rect 4120 -450 4160 -445
rect 4120 -480 4125 -450
rect 4125 -480 4155 -450
rect 4155 -480 4160 -450
rect 4120 -485 4160 -480
rect 4120 -515 4160 -510
rect 4120 -545 4125 -515
rect 4125 -545 4155 -515
rect 4155 -545 4160 -515
rect 4120 -550 4160 -545
rect 4120 -575 4160 -570
rect 4120 -605 4125 -575
rect 4125 -605 4155 -575
rect 4155 -605 4160 -575
rect 4120 -610 4160 -605
rect 4120 -640 4160 -635
rect 4120 -670 4125 -640
rect 4125 -670 4155 -640
rect 4155 -670 4160 -640
rect 4120 -675 4160 -670
rect 4120 -710 4160 -705
rect 4120 -740 4125 -710
rect 4125 -740 4155 -710
rect 4155 -740 4160 -710
rect 4120 -745 4160 -740
rect 4120 -780 4160 -775
rect 4120 -810 4125 -780
rect 4125 -810 4155 -780
rect 4155 -810 4160 -780
rect 4120 -815 4160 -810
rect 4120 -850 4160 -845
rect 4120 -880 4125 -850
rect 4125 -880 4155 -850
rect 4155 -880 4160 -850
rect 4120 -885 4160 -880
rect 4120 -915 4160 -910
rect 4120 -945 4125 -915
rect 4125 -945 4155 -915
rect 4155 -945 4160 -915
rect 4120 -950 4160 -945
rect 4120 -975 4160 -970
rect 4120 -1005 4125 -975
rect 4125 -1005 4155 -975
rect 4155 -1005 4160 -975
rect 4120 -1010 4160 -1005
rect 4120 -1040 4160 -1035
rect 4120 -1070 4125 -1040
rect 4125 -1070 4155 -1040
rect 4155 -1070 4160 -1040
rect 4120 -1075 4160 -1070
rect 4120 -1110 4160 -1105
rect 4120 -1140 4125 -1110
rect 4125 -1140 4155 -1110
rect 4155 -1140 4160 -1110
rect 4120 -1145 4160 -1140
rect 4120 -1180 4160 -1175
rect 4120 -1210 4125 -1180
rect 4125 -1210 4155 -1180
rect 4155 -1210 4160 -1180
rect 4120 -1215 4160 -1210
rect 4120 -1250 4160 -1245
rect 4120 -1280 4125 -1250
rect 4125 -1280 4155 -1250
rect 4155 -1280 4160 -1250
rect 4120 -1285 4160 -1280
rect 4120 -1315 4160 -1310
rect 4120 -1345 4125 -1315
rect 4125 -1345 4155 -1315
rect 4155 -1345 4160 -1315
rect 4120 -1350 4160 -1345
rect 4470 225 4510 230
rect 4470 195 4475 225
rect 4475 195 4505 225
rect 4505 195 4510 225
rect 4470 190 4510 195
rect 4470 160 4510 165
rect 4470 130 4475 160
rect 4475 130 4505 160
rect 4505 130 4510 160
rect 4470 125 4510 130
rect 4470 90 4510 95
rect 4470 60 4475 90
rect 4475 60 4505 90
rect 4505 60 4510 90
rect 4470 55 4510 60
rect 4470 20 4510 25
rect 4470 -10 4475 20
rect 4475 -10 4505 20
rect 4505 -10 4510 20
rect 4470 -15 4510 -10
rect 4470 -50 4510 -45
rect 4470 -80 4475 -50
rect 4475 -80 4505 -50
rect 4505 -80 4510 -50
rect 4470 -85 4510 -80
rect 4470 -115 4510 -110
rect 4470 -145 4475 -115
rect 4475 -145 4505 -115
rect 4505 -145 4510 -115
rect 4470 -150 4510 -145
rect 4470 -175 4510 -170
rect 4470 -205 4475 -175
rect 4475 -205 4505 -175
rect 4505 -205 4510 -175
rect 4470 -210 4510 -205
rect 4470 -240 4510 -235
rect 4470 -270 4475 -240
rect 4475 -270 4505 -240
rect 4505 -270 4510 -240
rect 4470 -275 4510 -270
rect 4470 -310 4510 -305
rect 4470 -340 4475 -310
rect 4475 -340 4505 -310
rect 4505 -340 4510 -310
rect 4470 -345 4510 -340
rect 4470 -380 4510 -375
rect 4470 -410 4475 -380
rect 4475 -410 4505 -380
rect 4505 -410 4510 -380
rect 4470 -415 4510 -410
rect 4470 -450 4510 -445
rect 4470 -480 4475 -450
rect 4475 -480 4505 -450
rect 4505 -480 4510 -450
rect 4470 -485 4510 -480
rect 4470 -515 4510 -510
rect 4470 -545 4475 -515
rect 4475 -545 4505 -515
rect 4505 -545 4510 -515
rect 4470 -550 4510 -545
rect 4470 -575 4510 -570
rect 4470 -605 4475 -575
rect 4475 -605 4505 -575
rect 4505 -605 4510 -575
rect 4470 -610 4510 -605
rect 4470 -640 4510 -635
rect 4470 -670 4475 -640
rect 4475 -670 4505 -640
rect 4505 -670 4510 -640
rect 4470 -675 4510 -670
rect 4470 -710 4510 -705
rect 4470 -740 4475 -710
rect 4475 -740 4505 -710
rect 4505 -740 4510 -710
rect 4470 -745 4510 -740
rect 4470 -780 4510 -775
rect 4470 -810 4475 -780
rect 4475 -810 4505 -780
rect 4505 -810 4510 -780
rect 4470 -815 4510 -810
rect 4470 -850 4510 -845
rect 4470 -880 4475 -850
rect 4475 -880 4505 -850
rect 4505 -880 4510 -850
rect 4470 -885 4510 -880
rect 4470 -915 4510 -910
rect 4470 -945 4475 -915
rect 4475 -945 4505 -915
rect 4505 -945 4510 -915
rect 4470 -950 4510 -945
rect 4470 -975 4510 -970
rect 4470 -1005 4475 -975
rect 4475 -1005 4505 -975
rect 4505 -1005 4510 -975
rect 4470 -1010 4510 -1005
rect 4470 -1040 4510 -1035
rect 4470 -1070 4475 -1040
rect 4475 -1070 4505 -1040
rect 4505 -1070 4510 -1040
rect 4470 -1075 4510 -1070
rect 4470 -1110 4510 -1105
rect 4470 -1140 4475 -1110
rect 4475 -1140 4505 -1110
rect 4505 -1140 4510 -1110
rect 4470 -1145 4510 -1140
rect 4470 -1180 4510 -1175
rect 4470 -1210 4475 -1180
rect 4475 -1210 4505 -1180
rect 4505 -1210 4510 -1180
rect 4470 -1215 4510 -1210
rect 4470 -1250 4510 -1245
rect 4470 -1280 4475 -1250
rect 4475 -1280 4505 -1250
rect 4505 -1280 4510 -1250
rect 4470 -1285 4510 -1280
rect 4470 -1315 4510 -1310
rect 4470 -1345 4475 -1315
rect 4475 -1345 4505 -1315
rect 4505 -1345 4510 -1315
rect 4470 -1350 4510 -1345
rect 4820 225 4860 230
rect 4820 195 4825 225
rect 4825 195 4855 225
rect 4855 195 4860 225
rect 4820 190 4860 195
rect 4820 160 4860 165
rect 4820 130 4825 160
rect 4825 130 4855 160
rect 4855 130 4860 160
rect 4820 125 4860 130
rect 4820 90 4860 95
rect 4820 60 4825 90
rect 4825 60 4855 90
rect 4855 60 4860 90
rect 4820 55 4860 60
rect 4820 20 4860 25
rect 4820 -10 4825 20
rect 4825 -10 4855 20
rect 4855 -10 4860 20
rect 4820 -15 4860 -10
rect 4820 -50 4860 -45
rect 4820 -80 4825 -50
rect 4825 -80 4855 -50
rect 4855 -80 4860 -50
rect 4820 -85 4860 -80
rect 4820 -115 4860 -110
rect 4820 -145 4825 -115
rect 4825 -145 4855 -115
rect 4855 -145 4860 -115
rect 4820 -150 4860 -145
rect 4820 -175 4860 -170
rect 4820 -205 4825 -175
rect 4825 -205 4855 -175
rect 4855 -205 4860 -175
rect 4820 -210 4860 -205
rect 4820 -240 4860 -235
rect 4820 -270 4825 -240
rect 4825 -270 4855 -240
rect 4855 -270 4860 -240
rect 4820 -275 4860 -270
rect 4820 -310 4860 -305
rect 4820 -340 4825 -310
rect 4825 -340 4855 -310
rect 4855 -340 4860 -310
rect 4820 -345 4860 -340
rect 4820 -380 4860 -375
rect 4820 -410 4825 -380
rect 4825 -410 4855 -380
rect 4855 -410 4860 -380
rect 4820 -415 4860 -410
rect 4820 -450 4860 -445
rect 4820 -480 4825 -450
rect 4825 -480 4855 -450
rect 4855 -480 4860 -450
rect 4820 -485 4860 -480
rect 4820 -515 4860 -510
rect 4820 -545 4825 -515
rect 4825 -545 4855 -515
rect 4855 -545 4860 -515
rect 4820 -550 4860 -545
rect 4820 -575 4860 -570
rect 4820 -605 4825 -575
rect 4825 -605 4855 -575
rect 4855 -605 4860 -575
rect 4820 -610 4860 -605
rect 4820 -640 4860 -635
rect 4820 -670 4825 -640
rect 4825 -670 4855 -640
rect 4855 -670 4860 -640
rect 4820 -675 4860 -670
rect 4820 -710 4860 -705
rect 4820 -740 4825 -710
rect 4825 -740 4855 -710
rect 4855 -740 4860 -710
rect 4820 -745 4860 -740
rect 4820 -780 4860 -775
rect 4820 -810 4825 -780
rect 4825 -810 4855 -780
rect 4855 -810 4860 -780
rect 4820 -815 4860 -810
rect 4820 -850 4860 -845
rect 4820 -880 4825 -850
rect 4825 -880 4855 -850
rect 4855 -880 4860 -850
rect 4820 -885 4860 -880
rect 4820 -915 4860 -910
rect 4820 -945 4825 -915
rect 4825 -945 4855 -915
rect 4855 -945 4860 -915
rect 4820 -950 4860 -945
rect 4820 -975 4860 -970
rect 4820 -1005 4825 -975
rect 4825 -1005 4855 -975
rect 4855 -1005 4860 -975
rect 4820 -1010 4860 -1005
rect 4820 -1040 4860 -1035
rect 4820 -1070 4825 -1040
rect 4825 -1070 4855 -1040
rect 4855 -1070 4860 -1040
rect 4820 -1075 4860 -1070
rect 4820 -1110 4860 -1105
rect 4820 -1140 4825 -1110
rect 4825 -1140 4855 -1110
rect 4855 -1140 4860 -1110
rect 4820 -1145 4860 -1140
rect 4820 -1180 4860 -1175
rect 4820 -1210 4825 -1180
rect 4825 -1210 4855 -1180
rect 4855 -1210 4860 -1180
rect 4820 -1215 4860 -1210
rect 4820 -1250 4860 -1245
rect 4820 -1280 4825 -1250
rect 4825 -1280 4855 -1250
rect 4855 -1280 4860 -1250
rect 4820 -1285 4860 -1280
rect 4820 -1315 4860 -1310
rect 4820 -1345 4825 -1315
rect 4825 -1345 4855 -1315
rect 4855 -1345 4860 -1315
rect 4820 -1350 4860 -1345
rect 5170 225 5210 230
rect 5170 195 5175 225
rect 5175 195 5205 225
rect 5205 195 5210 225
rect 5170 190 5210 195
rect 5170 160 5210 165
rect 5170 130 5175 160
rect 5175 130 5205 160
rect 5205 130 5210 160
rect 5170 125 5210 130
rect 5170 90 5210 95
rect 5170 60 5175 90
rect 5175 60 5205 90
rect 5205 60 5210 90
rect 5170 55 5210 60
rect 5170 20 5210 25
rect 5170 -10 5175 20
rect 5175 -10 5205 20
rect 5205 -10 5210 20
rect 5170 -15 5210 -10
rect 5170 -50 5210 -45
rect 5170 -80 5175 -50
rect 5175 -80 5205 -50
rect 5205 -80 5210 -50
rect 5170 -85 5210 -80
rect 5170 -115 5210 -110
rect 5170 -145 5175 -115
rect 5175 -145 5205 -115
rect 5205 -145 5210 -115
rect 5170 -150 5210 -145
rect 5170 -175 5210 -170
rect 5170 -205 5175 -175
rect 5175 -205 5205 -175
rect 5205 -205 5210 -175
rect 5170 -210 5210 -205
rect 5170 -240 5210 -235
rect 5170 -270 5175 -240
rect 5175 -270 5205 -240
rect 5205 -270 5210 -240
rect 5170 -275 5210 -270
rect 5170 -310 5210 -305
rect 5170 -340 5175 -310
rect 5175 -340 5205 -310
rect 5205 -340 5210 -310
rect 5170 -345 5210 -340
rect 5170 -380 5210 -375
rect 5170 -410 5175 -380
rect 5175 -410 5205 -380
rect 5205 -410 5210 -380
rect 5170 -415 5210 -410
rect 5170 -450 5210 -445
rect 5170 -480 5175 -450
rect 5175 -480 5205 -450
rect 5205 -480 5210 -450
rect 5170 -485 5210 -480
rect 5170 -515 5210 -510
rect 5170 -545 5175 -515
rect 5175 -545 5205 -515
rect 5205 -545 5210 -515
rect 5170 -550 5210 -545
rect 5170 -575 5210 -570
rect 5170 -605 5175 -575
rect 5175 -605 5205 -575
rect 5205 -605 5210 -575
rect 5170 -610 5210 -605
rect 5170 -640 5210 -635
rect 5170 -670 5175 -640
rect 5175 -670 5205 -640
rect 5205 -670 5210 -640
rect 5170 -675 5210 -670
rect 5170 -710 5210 -705
rect 5170 -740 5175 -710
rect 5175 -740 5205 -710
rect 5205 -740 5210 -710
rect 5170 -745 5210 -740
rect 5170 -780 5210 -775
rect 5170 -810 5175 -780
rect 5175 -810 5205 -780
rect 5205 -810 5210 -780
rect 5170 -815 5210 -810
rect 5170 -850 5210 -845
rect 5170 -880 5175 -850
rect 5175 -880 5205 -850
rect 5205 -880 5210 -850
rect 5170 -885 5210 -880
rect 5170 -915 5210 -910
rect 5170 -945 5175 -915
rect 5175 -945 5205 -915
rect 5205 -945 5210 -915
rect 5170 -950 5210 -945
rect 5170 -975 5210 -970
rect 5170 -1005 5175 -975
rect 5175 -1005 5205 -975
rect 5205 -1005 5210 -975
rect 5170 -1010 5210 -1005
rect 5170 -1040 5210 -1035
rect 5170 -1070 5175 -1040
rect 5175 -1070 5205 -1040
rect 5205 -1070 5210 -1040
rect 5170 -1075 5210 -1070
rect 5170 -1110 5210 -1105
rect 5170 -1140 5175 -1110
rect 5175 -1140 5205 -1110
rect 5205 -1140 5210 -1110
rect 5170 -1145 5210 -1140
rect 5170 -1180 5210 -1175
rect 5170 -1210 5175 -1180
rect 5175 -1210 5205 -1180
rect 5205 -1210 5210 -1180
rect 5170 -1215 5210 -1210
rect 5170 -1250 5210 -1245
rect 5170 -1280 5175 -1250
rect 5175 -1280 5205 -1250
rect 5205 -1280 5210 -1250
rect 5170 -1285 5210 -1280
rect 5170 -1315 5210 -1310
rect 5170 -1345 5175 -1315
rect 5175 -1345 5205 -1315
rect 5205 -1345 5210 -1315
rect 5170 -1350 5210 -1345
rect 5520 225 5560 230
rect 5520 195 5525 225
rect 5525 195 5555 225
rect 5555 195 5560 225
rect 5520 190 5560 195
rect 5520 160 5560 165
rect 5520 130 5525 160
rect 5525 130 5555 160
rect 5555 130 5560 160
rect 5520 125 5560 130
rect 5520 90 5560 95
rect 5520 60 5525 90
rect 5525 60 5555 90
rect 5555 60 5560 90
rect 5520 55 5560 60
rect 5520 20 5560 25
rect 5520 -10 5525 20
rect 5525 -10 5555 20
rect 5555 -10 5560 20
rect 5520 -15 5560 -10
rect 5520 -50 5560 -45
rect 5520 -80 5525 -50
rect 5525 -80 5555 -50
rect 5555 -80 5560 -50
rect 5520 -85 5560 -80
rect 5520 -115 5560 -110
rect 5520 -145 5525 -115
rect 5525 -145 5555 -115
rect 5555 -145 5560 -115
rect 5520 -150 5560 -145
rect 5520 -175 5560 -170
rect 5520 -205 5525 -175
rect 5525 -205 5555 -175
rect 5555 -205 5560 -175
rect 5520 -210 5560 -205
rect 5520 -240 5560 -235
rect 5520 -270 5525 -240
rect 5525 -270 5555 -240
rect 5555 -270 5560 -240
rect 5520 -275 5560 -270
rect 5520 -310 5560 -305
rect 5520 -340 5525 -310
rect 5525 -340 5555 -310
rect 5555 -340 5560 -310
rect 5520 -345 5560 -340
rect 5520 -380 5560 -375
rect 5520 -410 5525 -380
rect 5525 -410 5555 -380
rect 5555 -410 5560 -380
rect 5520 -415 5560 -410
rect 5520 -450 5560 -445
rect 5520 -480 5525 -450
rect 5525 -480 5555 -450
rect 5555 -480 5560 -450
rect 5520 -485 5560 -480
rect 5520 -515 5560 -510
rect 5520 -545 5525 -515
rect 5525 -545 5555 -515
rect 5555 -545 5560 -515
rect 5520 -550 5560 -545
rect 5520 -575 5560 -570
rect 5520 -605 5525 -575
rect 5525 -605 5555 -575
rect 5555 -605 5560 -575
rect 5520 -610 5560 -605
rect 5520 -640 5560 -635
rect 5520 -670 5525 -640
rect 5525 -670 5555 -640
rect 5555 -670 5560 -640
rect 5520 -675 5560 -670
rect 5520 -710 5560 -705
rect 5520 -740 5525 -710
rect 5525 -740 5555 -710
rect 5555 -740 5560 -710
rect 5520 -745 5560 -740
rect 5520 -780 5560 -775
rect 5520 -810 5525 -780
rect 5525 -810 5555 -780
rect 5555 -810 5560 -780
rect 5520 -815 5560 -810
rect 5520 -850 5560 -845
rect 5520 -880 5525 -850
rect 5525 -880 5555 -850
rect 5555 -880 5560 -850
rect 5520 -885 5560 -880
rect 5520 -915 5560 -910
rect 5520 -945 5525 -915
rect 5525 -945 5555 -915
rect 5555 -945 5560 -915
rect 5520 -950 5560 -945
rect 5520 -975 5560 -970
rect 5520 -1005 5525 -975
rect 5525 -1005 5555 -975
rect 5555 -1005 5560 -975
rect 5520 -1010 5560 -1005
rect 5520 -1040 5560 -1035
rect 5520 -1070 5525 -1040
rect 5525 -1070 5555 -1040
rect 5555 -1070 5560 -1040
rect 5520 -1075 5560 -1070
rect 5520 -1110 5560 -1105
rect 5520 -1140 5525 -1110
rect 5525 -1140 5555 -1110
rect 5555 -1140 5560 -1110
rect 5520 -1145 5560 -1140
rect 5520 -1180 5560 -1175
rect 5520 -1210 5525 -1180
rect 5525 -1210 5555 -1180
rect 5555 -1210 5560 -1180
rect 5520 -1215 5560 -1210
rect 5520 -1250 5560 -1245
rect 5520 -1280 5525 -1250
rect 5525 -1280 5555 -1250
rect 5555 -1280 5560 -1250
rect 5520 -1285 5560 -1280
rect 5520 -1315 5560 -1310
rect 5520 -1345 5525 -1315
rect 5525 -1345 5555 -1315
rect 5555 -1345 5560 -1315
rect 5520 -1350 5560 -1345
rect 5870 225 5910 230
rect 5870 195 5875 225
rect 5875 195 5905 225
rect 5905 195 5910 225
rect 5870 190 5910 195
rect 5870 160 5910 165
rect 5870 130 5875 160
rect 5875 130 5905 160
rect 5905 130 5910 160
rect 5870 125 5910 130
rect 5870 90 5910 95
rect 5870 60 5875 90
rect 5875 60 5905 90
rect 5905 60 5910 90
rect 5870 55 5910 60
rect 5870 20 5910 25
rect 5870 -10 5875 20
rect 5875 -10 5905 20
rect 5905 -10 5910 20
rect 5870 -15 5910 -10
rect 5870 -50 5910 -45
rect 5870 -80 5875 -50
rect 5875 -80 5905 -50
rect 5905 -80 5910 -50
rect 5870 -85 5910 -80
rect 5870 -115 5910 -110
rect 5870 -145 5875 -115
rect 5875 -145 5905 -115
rect 5905 -145 5910 -115
rect 5870 -150 5910 -145
rect 5870 -175 5910 -170
rect 5870 -205 5875 -175
rect 5875 -205 5905 -175
rect 5905 -205 5910 -175
rect 5870 -210 5910 -205
rect 5870 -240 5910 -235
rect 5870 -270 5875 -240
rect 5875 -270 5905 -240
rect 5905 -270 5910 -240
rect 5870 -275 5910 -270
rect 5870 -310 5910 -305
rect 5870 -340 5875 -310
rect 5875 -340 5905 -310
rect 5905 -340 5910 -310
rect 5870 -345 5910 -340
rect 5870 -380 5910 -375
rect 5870 -410 5875 -380
rect 5875 -410 5905 -380
rect 5905 -410 5910 -380
rect 5870 -415 5910 -410
rect 5870 -450 5910 -445
rect 5870 -480 5875 -450
rect 5875 -480 5905 -450
rect 5905 -480 5910 -450
rect 5870 -485 5910 -480
rect 5870 -515 5910 -510
rect 5870 -545 5875 -515
rect 5875 -545 5905 -515
rect 5905 -545 5910 -515
rect 5870 -550 5910 -545
rect 5870 -575 5910 -570
rect 5870 -605 5875 -575
rect 5875 -605 5905 -575
rect 5905 -605 5910 -575
rect 5870 -610 5910 -605
rect 5870 -640 5910 -635
rect 5870 -670 5875 -640
rect 5875 -670 5905 -640
rect 5905 -670 5910 -640
rect 5870 -675 5910 -670
rect 5870 -710 5910 -705
rect 5870 -740 5875 -710
rect 5875 -740 5905 -710
rect 5905 -740 5910 -710
rect 5870 -745 5910 -740
rect 5870 -780 5910 -775
rect 5870 -810 5875 -780
rect 5875 -810 5905 -780
rect 5905 -810 5910 -780
rect 5870 -815 5910 -810
rect 5870 -850 5910 -845
rect 5870 -880 5875 -850
rect 5875 -880 5905 -850
rect 5905 -880 5910 -850
rect 5870 -885 5910 -880
rect 5870 -915 5910 -910
rect 5870 -945 5875 -915
rect 5875 -945 5905 -915
rect 5905 -945 5910 -915
rect 5870 -950 5910 -945
rect 5870 -975 5910 -970
rect 5870 -1005 5875 -975
rect 5875 -1005 5905 -975
rect 5905 -1005 5910 -975
rect 5870 -1010 5910 -1005
rect 5870 -1040 5910 -1035
rect 5870 -1070 5875 -1040
rect 5875 -1070 5905 -1040
rect 5905 -1070 5910 -1040
rect 5870 -1075 5910 -1070
rect 5870 -1110 5910 -1105
rect 5870 -1140 5875 -1110
rect 5875 -1140 5905 -1110
rect 5905 -1140 5910 -1110
rect 5870 -1145 5910 -1140
rect 5870 -1180 5910 -1175
rect 5870 -1210 5875 -1180
rect 5875 -1210 5905 -1180
rect 5905 -1210 5910 -1180
rect 5870 -1215 5910 -1210
rect 5870 -1250 5910 -1245
rect 5870 -1280 5875 -1250
rect 5875 -1280 5905 -1250
rect 5905 -1280 5910 -1250
rect 5870 -1285 5910 -1280
rect 5870 -1315 5910 -1310
rect 5870 -1345 5875 -1315
rect 5875 -1345 5905 -1315
rect 5905 -1345 5910 -1315
rect 5870 -1350 5910 -1345
rect 6220 225 6260 230
rect 6220 195 6225 225
rect 6225 195 6255 225
rect 6255 195 6260 225
rect 6220 190 6260 195
rect 6220 160 6260 165
rect 6220 130 6225 160
rect 6225 130 6255 160
rect 6255 130 6260 160
rect 6220 125 6260 130
rect 6220 90 6260 95
rect 6220 60 6225 90
rect 6225 60 6255 90
rect 6255 60 6260 90
rect 6220 55 6260 60
rect 6220 20 6260 25
rect 6220 -10 6225 20
rect 6225 -10 6255 20
rect 6255 -10 6260 20
rect 6220 -15 6260 -10
rect 6220 -50 6260 -45
rect 6220 -80 6225 -50
rect 6225 -80 6255 -50
rect 6255 -80 6260 -50
rect 6220 -85 6260 -80
rect 6220 -115 6260 -110
rect 6220 -145 6225 -115
rect 6225 -145 6255 -115
rect 6255 -145 6260 -115
rect 6220 -150 6260 -145
rect 6220 -175 6260 -170
rect 6220 -205 6225 -175
rect 6225 -205 6255 -175
rect 6255 -205 6260 -175
rect 6220 -210 6260 -205
rect 6220 -240 6260 -235
rect 6220 -270 6225 -240
rect 6225 -270 6255 -240
rect 6255 -270 6260 -240
rect 6220 -275 6260 -270
rect 6220 -310 6260 -305
rect 6220 -340 6225 -310
rect 6225 -340 6255 -310
rect 6255 -340 6260 -310
rect 6220 -345 6260 -340
rect 6220 -380 6260 -375
rect 6220 -410 6225 -380
rect 6225 -410 6255 -380
rect 6255 -410 6260 -380
rect 6220 -415 6260 -410
rect 6220 -450 6260 -445
rect 6220 -480 6225 -450
rect 6225 -480 6255 -450
rect 6255 -480 6260 -450
rect 6220 -485 6260 -480
rect 6220 -515 6260 -510
rect 6220 -545 6225 -515
rect 6225 -545 6255 -515
rect 6255 -545 6260 -515
rect 6220 -550 6260 -545
rect 6220 -575 6260 -570
rect 6220 -605 6225 -575
rect 6225 -605 6255 -575
rect 6255 -605 6260 -575
rect 6220 -610 6260 -605
rect 6220 -640 6260 -635
rect 6220 -670 6225 -640
rect 6225 -670 6255 -640
rect 6255 -670 6260 -640
rect 6220 -675 6260 -670
rect 6220 -710 6260 -705
rect 6220 -740 6225 -710
rect 6225 -740 6255 -710
rect 6255 -740 6260 -710
rect 6220 -745 6260 -740
rect 6220 -780 6260 -775
rect 6220 -810 6225 -780
rect 6225 -810 6255 -780
rect 6255 -810 6260 -780
rect 6220 -815 6260 -810
rect 6220 -850 6260 -845
rect 6220 -880 6225 -850
rect 6225 -880 6255 -850
rect 6255 -880 6260 -850
rect 6220 -885 6260 -880
rect 6220 -915 6260 -910
rect 6220 -945 6225 -915
rect 6225 -945 6255 -915
rect 6255 -945 6260 -915
rect 6220 -950 6260 -945
rect 6220 -975 6260 -970
rect 6220 -1005 6225 -975
rect 6225 -1005 6255 -975
rect 6255 -1005 6260 -975
rect 6220 -1010 6260 -1005
rect 6220 -1040 6260 -1035
rect 6220 -1070 6225 -1040
rect 6225 -1070 6255 -1040
rect 6255 -1070 6260 -1040
rect 6220 -1075 6260 -1070
rect 6220 -1110 6260 -1105
rect 6220 -1140 6225 -1110
rect 6225 -1140 6255 -1110
rect 6255 -1140 6260 -1110
rect 6220 -1145 6260 -1140
rect 6220 -1180 6260 -1175
rect 6220 -1210 6225 -1180
rect 6225 -1210 6255 -1180
rect 6255 -1210 6260 -1180
rect 6220 -1215 6260 -1210
rect 6220 -1250 6260 -1245
rect 6220 -1280 6225 -1250
rect 6225 -1280 6255 -1250
rect 6255 -1280 6260 -1250
rect 6220 -1285 6260 -1280
rect 6220 -1315 6260 -1310
rect 6220 -1345 6225 -1315
rect 6225 -1345 6255 -1315
rect 6255 -1345 6260 -1315
rect 6220 -1350 6260 -1345
rect 6570 225 6610 230
rect 6570 195 6575 225
rect 6575 195 6605 225
rect 6605 195 6610 225
rect 6570 190 6610 195
rect 6570 160 6610 165
rect 6570 130 6575 160
rect 6575 130 6605 160
rect 6605 130 6610 160
rect 6570 125 6610 130
rect 6570 90 6610 95
rect 6570 60 6575 90
rect 6575 60 6605 90
rect 6605 60 6610 90
rect 6570 55 6610 60
rect 6570 20 6610 25
rect 6570 -10 6575 20
rect 6575 -10 6605 20
rect 6605 -10 6610 20
rect 6570 -15 6610 -10
rect 6570 -50 6610 -45
rect 6570 -80 6575 -50
rect 6575 -80 6605 -50
rect 6605 -80 6610 -50
rect 6570 -85 6610 -80
rect 6570 -115 6610 -110
rect 6570 -145 6575 -115
rect 6575 -145 6605 -115
rect 6605 -145 6610 -115
rect 6570 -150 6610 -145
rect 6570 -175 6610 -170
rect 6570 -205 6575 -175
rect 6575 -205 6605 -175
rect 6605 -205 6610 -175
rect 6570 -210 6610 -205
rect 6570 -240 6610 -235
rect 6570 -270 6575 -240
rect 6575 -270 6605 -240
rect 6605 -270 6610 -240
rect 6570 -275 6610 -270
rect 6570 -310 6610 -305
rect 6570 -340 6575 -310
rect 6575 -340 6605 -310
rect 6605 -340 6610 -310
rect 6570 -345 6610 -340
rect 6570 -380 6610 -375
rect 6570 -410 6575 -380
rect 6575 -410 6605 -380
rect 6605 -410 6610 -380
rect 6570 -415 6610 -410
rect 6570 -450 6610 -445
rect 6570 -480 6575 -450
rect 6575 -480 6605 -450
rect 6605 -480 6610 -450
rect 6570 -485 6610 -480
rect 6570 -515 6610 -510
rect 6570 -545 6575 -515
rect 6575 -545 6605 -515
rect 6605 -545 6610 -515
rect 6570 -550 6610 -545
rect 6570 -575 6610 -570
rect 6570 -605 6575 -575
rect 6575 -605 6605 -575
rect 6605 -605 6610 -575
rect 6570 -610 6610 -605
rect 6570 -640 6610 -635
rect 6570 -670 6575 -640
rect 6575 -670 6605 -640
rect 6605 -670 6610 -640
rect 6570 -675 6610 -670
rect 6570 -710 6610 -705
rect 6570 -740 6575 -710
rect 6575 -740 6605 -710
rect 6605 -740 6610 -710
rect 6570 -745 6610 -740
rect 6570 -780 6610 -775
rect 6570 -810 6575 -780
rect 6575 -810 6605 -780
rect 6605 -810 6610 -780
rect 6570 -815 6610 -810
rect 6570 -850 6610 -845
rect 6570 -880 6575 -850
rect 6575 -880 6605 -850
rect 6605 -880 6610 -850
rect 6570 -885 6610 -880
rect 6570 -915 6610 -910
rect 6570 -945 6575 -915
rect 6575 -945 6605 -915
rect 6605 -945 6610 -915
rect 6570 -950 6610 -945
rect 6570 -975 6610 -970
rect 6570 -1005 6575 -975
rect 6575 -1005 6605 -975
rect 6605 -1005 6610 -975
rect 6570 -1010 6610 -1005
rect 6570 -1040 6610 -1035
rect 6570 -1070 6575 -1040
rect 6575 -1070 6605 -1040
rect 6605 -1070 6610 -1040
rect 6570 -1075 6610 -1070
rect 6570 -1110 6610 -1105
rect 6570 -1140 6575 -1110
rect 6575 -1140 6605 -1110
rect 6605 -1140 6610 -1110
rect 6570 -1145 6610 -1140
rect 6570 -1180 6610 -1175
rect 6570 -1210 6575 -1180
rect 6575 -1210 6605 -1180
rect 6605 -1210 6610 -1180
rect 6570 -1215 6610 -1210
rect 6570 -1250 6610 -1245
rect 6570 -1280 6575 -1250
rect 6575 -1280 6605 -1250
rect 6605 -1280 6610 -1250
rect 6570 -1285 6610 -1280
rect 6570 -1315 6610 -1310
rect 6570 -1345 6575 -1315
rect 6575 -1345 6605 -1315
rect 6605 -1345 6610 -1315
rect 6570 -1350 6610 -1345
rect 6920 225 6960 230
rect 6920 195 6925 225
rect 6925 195 6955 225
rect 6955 195 6960 225
rect 6920 190 6960 195
rect 6920 160 6960 165
rect 6920 130 6925 160
rect 6925 130 6955 160
rect 6955 130 6960 160
rect 6920 125 6960 130
rect 6920 90 6960 95
rect 6920 60 6925 90
rect 6925 60 6955 90
rect 6955 60 6960 90
rect 6920 55 6960 60
rect 6920 20 6960 25
rect 6920 -10 6925 20
rect 6925 -10 6955 20
rect 6955 -10 6960 20
rect 6920 -15 6960 -10
rect 6920 -50 6960 -45
rect 6920 -80 6925 -50
rect 6925 -80 6955 -50
rect 6955 -80 6960 -50
rect 6920 -85 6960 -80
rect 6920 -115 6960 -110
rect 6920 -145 6925 -115
rect 6925 -145 6955 -115
rect 6955 -145 6960 -115
rect 6920 -150 6960 -145
rect 6920 -175 6960 -170
rect 6920 -205 6925 -175
rect 6925 -205 6955 -175
rect 6955 -205 6960 -175
rect 6920 -210 6960 -205
rect 6920 -240 6960 -235
rect 6920 -270 6925 -240
rect 6925 -270 6955 -240
rect 6955 -270 6960 -240
rect 6920 -275 6960 -270
rect 6920 -310 6960 -305
rect 6920 -340 6925 -310
rect 6925 -340 6955 -310
rect 6955 -340 6960 -310
rect 6920 -345 6960 -340
rect 6920 -380 6960 -375
rect 6920 -410 6925 -380
rect 6925 -410 6955 -380
rect 6955 -410 6960 -380
rect 6920 -415 6960 -410
rect 6920 -450 6960 -445
rect 6920 -480 6925 -450
rect 6925 -480 6955 -450
rect 6955 -480 6960 -450
rect 6920 -485 6960 -480
rect 6920 -515 6960 -510
rect 6920 -545 6925 -515
rect 6925 -545 6955 -515
rect 6955 -545 6960 -515
rect 6920 -550 6960 -545
rect 6920 -575 6960 -570
rect 6920 -605 6925 -575
rect 6925 -605 6955 -575
rect 6955 -605 6960 -575
rect 6920 -610 6960 -605
rect 6920 -640 6960 -635
rect 6920 -670 6925 -640
rect 6925 -670 6955 -640
rect 6955 -670 6960 -640
rect 6920 -675 6960 -670
rect 6920 -710 6960 -705
rect 6920 -740 6925 -710
rect 6925 -740 6955 -710
rect 6955 -740 6960 -710
rect 6920 -745 6960 -740
rect 6920 -780 6960 -775
rect 6920 -810 6925 -780
rect 6925 -810 6955 -780
rect 6955 -810 6960 -780
rect 6920 -815 6960 -810
rect 6920 -850 6960 -845
rect 6920 -880 6925 -850
rect 6925 -880 6955 -850
rect 6955 -880 6960 -850
rect 6920 -885 6960 -880
rect 6920 -915 6960 -910
rect 6920 -945 6925 -915
rect 6925 -945 6955 -915
rect 6955 -945 6960 -915
rect 6920 -950 6960 -945
rect 6920 -975 6960 -970
rect 6920 -1005 6925 -975
rect 6925 -1005 6955 -975
rect 6955 -1005 6960 -975
rect 6920 -1010 6960 -1005
rect 6920 -1040 6960 -1035
rect 6920 -1070 6925 -1040
rect 6925 -1070 6955 -1040
rect 6955 -1070 6960 -1040
rect 6920 -1075 6960 -1070
rect 6920 -1110 6960 -1105
rect 6920 -1140 6925 -1110
rect 6925 -1140 6955 -1110
rect 6955 -1140 6960 -1110
rect 6920 -1145 6960 -1140
rect 6920 -1180 6960 -1175
rect 6920 -1210 6925 -1180
rect 6925 -1210 6955 -1180
rect 6955 -1210 6960 -1180
rect 6920 -1215 6960 -1210
rect 6920 -1250 6960 -1245
rect 6920 -1280 6925 -1250
rect 6925 -1280 6955 -1250
rect 6955 -1280 6960 -1250
rect 6920 -1285 6960 -1280
rect 6920 -1315 6960 -1310
rect 6920 -1345 6925 -1315
rect 6925 -1345 6955 -1315
rect 6955 -1345 6960 -1315
rect 6920 -1350 6960 -1345
rect 7270 225 7310 230
rect 7270 195 7275 225
rect 7275 195 7305 225
rect 7305 195 7310 225
rect 7270 190 7310 195
rect 7270 160 7310 165
rect 7270 130 7275 160
rect 7275 130 7305 160
rect 7305 130 7310 160
rect 7270 125 7310 130
rect 7270 90 7310 95
rect 7270 60 7275 90
rect 7275 60 7305 90
rect 7305 60 7310 90
rect 7270 55 7310 60
rect 7270 20 7310 25
rect 7270 -10 7275 20
rect 7275 -10 7305 20
rect 7305 -10 7310 20
rect 7270 -15 7310 -10
rect 7270 -50 7310 -45
rect 7270 -80 7275 -50
rect 7275 -80 7305 -50
rect 7305 -80 7310 -50
rect 7270 -85 7310 -80
rect 7270 -115 7310 -110
rect 7270 -145 7275 -115
rect 7275 -145 7305 -115
rect 7305 -145 7310 -115
rect 7270 -150 7310 -145
rect 7270 -175 7310 -170
rect 7270 -205 7275 -175
rect 7275 -205 7305 -175
rect 7305 -205 7310 -175
rect 7270 -210 7310 -205
rect 7270 -240 7310 -235
rect 7270 -270 7275 -240
rect 7275 -270 7305 -240
rect 7305 -270 7310 -240
rect 7270 -275 7310 -270
rect 7270 -310 7310 -305
rect 7270 -340 7275 -310
rect 7275 -340 7305 -310
rect 7305 -340 7310 -310
rect 7270 -345 7310 -340
rect 7270 -380 7310 -375
rect 7270 -410 7275 -380
rect 7275 -410 7305 -380
rect 7305 -410 7310 -380
rect 7270 -415 7310 -410
rect 7270 -450 7310 -445
rect 7270 -480 7275 -450
rect 7275 -480 7305 -450
rect 7305 -480 7310 -450
rect 7270 -485 7310 -480
rect 7270 -515 7310 -510
rect 7270 -545 7275 -515
rect 7275 -545 7305 -515
rect 7305 -545 7310 -515
rect 7270 -550 7310 -545
rect 7270 -575 7310 -570
rect 7270 -605 7275 -575
rect 7275 -605 7305 -575
rect 7305 -605 7310 -575
rect 7270 -610 7310 -605
rect 7270 -640 7310 -635
rect 7270 -670 7275 -640
rect 7275 -670 7305 -640
rect 7305 -670 7310 -640
rect 7270 -675 7310 -670
rect 7270 -710 7310 -705
rect 7270 -740 7275 -710
rect 7275 -740 7305 -710
rect 7305 -740 7310 -710
rect 7270 -745 7310 -740
rect 7270 -780 7310 -775
rect 7270 -810 7275 -780
rect 7275 -810 7305 -780
rect 7305 -810 7310 -780
rect 7270 -815 7310 -810
rect 7270 -850 7310 -845
rect 7270 -880 7275 -850
rect 7275 -880 7305 -850
rect 7305 -880 7310 -850
rect 7270 -885 7310 -880
rect 7270 -915 7310 -910
rect 7270 -945 7275 -915
rect 7275 -945 7305 -915
rect 7305 -945 7310 -915
rect 7270 -950 7310 -945
rect 7270 -975 7310 -970
rect 7270 -1005 7275 -975
rect 7275 -1005 7305 -975
rect 7305 -1005 7310 -975
rect 7270 -1010 7310 -1005
rect 7270 -1040 7310 -1035
rect 7270 -1070 7275 -1040
rect 7275 -1070 7305 -1040
rect 7305 -1070 7310 -1040
rect 7270 -1075 7310 -1070
rect 7270 -1110 7310 -1105
rect 7270 -1140 7275 -1110
rect 7275 -1140 7305 -1110
rect 7305 -1140 7310 -1110
rect 7270 -1145 7310 -1140
rect 7270 -1180 7310 -1175
rect 7270 -1210 7275 -1180
rect 7275 -1210 7305 -1180
rect 7305 -1210 7310 -1180
rect 7270 -1215 7310 -1210
rect 7270 -1250 7310 -1245
rect 7270 -1280 7275 -1250
rect 7275 -1280 7305 -1250
rect 7305 -1280 7310 -1250
rect 7270 -1285 7310 -1280
rect 7270 -1315 7310 -1310
rect 7270 -1345 7275 -1315
rect 7275 -1345 7305 -1315
rect 7305 -1345 7310 -1315
rect 7270 -1350 7310 -1345
rect 7620 225 7660 230
rect 7620 195 7625 225
rect 7625 195 7655 225
rect 7655 195 7660 225
rect 7620 190 7660 195
rect 7620 160 7660 165
rect 7620 130 7625 160
rect 7625 130 7655 160
rect 7655 130 7660 160
rect 7620 125 7660 130
rect 7620 90 7660 95
rect 7620 60 7625 90
rect 7625 60 7655 90
rect 7655 60 7660 90
rect 7620 55 7660 60
rect 7620 20 7660 25
rect 7620 -10 7625 20
rect 7625 -10 7655 20
rect 7655 -10 7660 20
rect 7620 -15 7660 -10
rect 7620 -50 7660 -45
rect 7620 -80 7625 -50
rect 7625 -80 7655 -50
rect 7655 -80 7660 -50
rect 7620 -85 7660 -80
rect 7620 -115 7660 -110
rect 7620 -145 7625 -115
rect 7625 -145 7655 -115
rect 7655 -145 7660 -115
rect 7620 -150 7660 -145
rect 7620 -175 7660 -170
rect 7620 -205 7625 -175
rect 7625 -205 7655 -175
rect 7655 -205 7660 -175
rect 7620 -210 7660 -205
rect 7620 -240 7660 -235
rect 7620 -270 7625 -240
rect 7625 -270 7655 -240
rect 7655 -270 7660 -240
rect 7620 -275 7660 -270
rect 7620 -310 7660 -305
rect 7620 -340 7625 -310
rect 7625 -340 7655 -310
rect 7655 -340 7660 -310
rect 7620 -345 7660 -340
rect 7620 -380 7660 -375
rect 7620 -410 7625 -380
rect 7625 -410 7655 -380
rect 7655 -410 7660 -380
rect 7620 -415 7660 -410
rect 7620 -450 7660 -445
rect 7620 -480 7625 -450
rect 7625 -480 7655 -450
rect 7655 -480 7660 -450
rect 7620 -485 7660 -480
rect 7620 -515 7660 -510
rect 7620 -545 7625 -515
rect 7625 -545 7655 -515
rect 7655 -545 7660 -515
rect 7620 -550 7660 -545
rect 7620 -575 7660 -570
rect 7620 -605 7625 -575
rect 7625 -605 7655 -575
rect 7655 -605 7660 -575
rect 7620 -610 7660 -605
rect 7620 -640 7660 -635
rect 7620 -670 7625 -640
rect 7625 -670 7655 -640
rect 7655 -670 7660 -640
rect 7620 -675 7660 -670
rect 7620 -710 7660 -705
rect 7620 -740 7625 -710
rect 7625 -740 7655 -710
rect 7655 -740 7660 -710
rect 7620 -745 7660 -740
rect 7620 -780 7660 -775
rect 7620 -810 7625 -780
rect 7625 -810 7655 -780
rect 7655 -810 7660 -780
rect 7620 -815 7660 -810
rect 7620 -850 7660 -845
rect 7620 -880 7625 -850
rect 7625 -880 7655 -850
rect 7655 -880 7660 -850
rect 7620 -885 7660 -880
rect 7620 -915 7660 -910
rect 7620 -945 7625 -915
rect 7625 -945 7655 -915
rect 7655 -945 7660 -915
rect 7620 -950 7660 -945
rect 7620 -975 7660 -970
rect 7620 -1005 7625 -975
rect 7625 -1005 7655 -975
rect 7655 -1005 7660 -975
rect 7620 -1010 7660 -1005
rect 7620 -1040 7660 -1035
rect 7620 -1070 7625 -1040
rect 7625 -1070 7655 -1040
rect 7655 -1070 7660 -1040
rect 7620 -1075 7660 -1070
rect 7620 -1110 7660 -1105
rect 7620 -1140 7625 -1110
rect 7625 -1140 7655 -1110
rect 7655 -1140 7660 -1110
rect 7620 -1145 7660 -1140
rect 7620 -1180 7660 -1175
rect 7620 -1210 7625 -1180
rect 7625 -1210 7655 -1180
rect 7655 -1210 7660 -1180
rect 7620 -1215 7660 -1210
rect 7620 -1250 7660 -1245
rect 7620 -1280 7625 -1250
rect 7625 -1280 7655 -1250
rect 7655 -1280 7660 -1250
rect 7620 -1285 7660 -1280
rect 7620 -1315 7660 -1310
rect 7620 -1345 7625 -1315
rect 7625 -1345 7655 -1315
rect 7655 -1345 7660 -1315
rect 7620 -1350 7660 -1345
rect 7970 225 8010 230
rect 7970 195 7975 225
rect 7975 195 8005 225
rect 8005 195 8010 225
rect 7970 190 8010 195
rect 7970 160 8010 165
rect 7970 130 7975 160
rect 7975 130 8005 160
rect 8005 130 8010 160
rect 7970 125 8010 130
rect 7970 90 8010 95
rect 7970 60 7975 90
rect 7975 60 8005 90
rect 8005 60 8010 90
rect 7970 55 8010 60
rect 7970 20 8010 25
rect 7970 -10 7975 20
rect 7975 -10 8005 20
rect 8005 -10 8010 20
rect 7970 -15 8010 -10
rect 7970 -50 8010 -45
rect 7970 -80 7975 -50
rect 7975 -80 8005 -50
rect 8005 -80 8010 -50
rect 7970 -85 8010 -80
rect 7970 -115 8010 -110
rect 7970 -145 7975 -115
rect 7975 -145 8005 -115
rect 8005 -145 8010 -115
rect 7970 -150 8010 -145
rect 7970 -175 8010 -170
rect 7970 -205 7975 -175
rect 7975 -205 8005 -175
rect 8005 -205 8010 -175
rect 7970 -210 8010 -205
rect 7970 -240 8010 -235
rect 7970 -270 7975 -240
rect 7975 -270 8005 -240
rect 8005 -270 8010 -240
rect 7970 -275 8010 -270
rect 7970 -310 8010 -305
rect 7970 -340 7975 -310
rect 7975 -340 8005 -310
rect 8005 -340 8010 -310
rect 7970 -345 8010 -340
rect 7970 -380 8010 -375
rect 7970 -410 7975 -380
rect 7975 -410 8005 -380
rect 8005 -410 8010 -380
rect 7970 -415 8010 -410
rect 7970 -450 8010 -445
rect 7970 -480 7975 -450
rect 7975 -480 8005 -450
rect 8005 -480 8010 -450
rect 7970 -485 8010 -480
rect 7970 -515 8010 -510
rect 7970 -545 7975 -515
rect 7975 -545 8005 -515
rect 8005 -545 8010 -515
rect 7970 -550 8010 -545
rect 7970 -575 8010 -570
rect 7970 -605 7975 -575
rect 7975 -605 8005 -575
rect 8005 -605 8010 -575
rect 7970 -610 8010 -605
rect 7970 -640 8010 -635
rect 7970 -670 7975 -640
rect 7975 -670 8005 -640
rect 8005 -670 8010 -640
rect 7970 -675 8010 -670
rect 7970 -710 8010 -705
rect 7970 -740 7975 -710
rect 7975 -740 8005 -710
rect 8005 -740 8010 -710
rect 7970 -745 8010 -740
rect 7970 -780 8010 -775
rect 7970 -810 7975 -780
rect 7975 -810 8005 -780
rect 8005 -810 8010 -780
rect 7970 -815 8010 -810
rect 7970 -850 8010 -845
rect 7970 -880 7975 -850
rect 7975 -880 8005 -850
rect 8005 -880 8010 -850
rect 7970 -885 8010 -880
rect 7970 -915 8010 -910
rect 7970 -945 7975 -915
rect 7975 -945 8005 -915
rect 8005 -945 8010 -915
rect 7970 -950 8010 -945
rect 7970 -975 8010 -970
rect 7970 -1005 7975 -975
rect 7975 -1005 8005 -975
rect 8005 -1005 8010 -975
rect 7970 -1010 8010 -1005
rect 7970 -1040 8010 -1035
rect 7970 -1070 7975 -1040
rect 7975 -1070 8005 -1040
rect 8005 -1070 8010 -1040
rect 7970 -1075 8010 -1070
rect 7970 -1110 8010 -1105
rect 7970 -1140 7975 -1110
rect 7975 -1140 8005 -1110
rect 8005 -1140 8010 -1110
rect 7970 -1145 8010 -1140
rect 7970 -1180 8010 -1175
rect 7970 -1210 7975 -1180
rect 7975 -1210 8005 -1180
rect 8005 -1210 8010 -1180
rect 7970 -1215 8010 -1210
rect 7970 -1250 8010 -1245
rect 7970 -1280 7975 -1250
rect 7975 -1280 8005 -1250
rect 8005 -1280 8010 -1250
rect 7970 -1285 8010 -1280
rect 7970 -1315 8010 -1310
rect 7970 -1345 7975 -1315
rect 7975 -1345 8005 -1315
rect 8005 -1345 8010 -1315
rect 7970 -1350 8010 -1345
rect 8320 225 8360 230
rect 8320 195 8325 225
rect 8325 195 8355 225
rect 8355 195 8360 225
rect 8320 190 8360 195
rect 8320 160 8360 165
rect 8320 130 8325 160
rect 8325 130 8355 160
rect 8355 130 8360 160
rect 8320 125 8360 130
rect 8320 90 8360 95
rect 8320 60 8325 90
rect 8325 60 8355 90
rect 8355 60 8360 90
rect 8320 55 8360 60
rect 8320 20 8360 25
rect 8320 -10 8325 20
rect 8325 -10 8355 20
rect 8355 -10 8360 20
rect 8320 -15 8360 -10
rect 8320 -50 8360 -45
rect 8320 -80 8325 -50
rect 8325 -80 8355 -50
rect 8355 -80 8360 -50
rect 8320 -85 8360 -80
rect 8320 -115 8360 -110
rect 8320 -145 8325 -115
rect 8325 -145 8355 -115
rect 8355 -145 8360 -115
rect 8320 -150 8360 -145
rect 8320 -175 8360 -170
rect 8320 -205 8325 -175
rect 8325 -205 8355 -175
rect 8355 -205 8360 -175
rect 8320 -210 8360 -205
rect 8320 -240 8360 -235
rect 8320 -270 8325 -240
rect 8325 -270 8355 -240
rect 8355 -270 8360 -240
rect 8320 -275 8360 -270
rect 8320 -310 8360 -305
rect 8320 -340 8325 -310
rect 8325 -340 8355 -310
rect 8355 -340 8360 -310
rect 8320 -345 8360 -340
rect 8320 -380 8360 -375
rect 8320 -410 8325 -380
rect 8325 -410 8355 -380
rect 8355 -410 8360 -380
rect 8320 -415 8360 -410
rect 8320 -450 8360 -445
rect 8320 -480 8325 -450
rect 8325 -480 8355 -450
rect 8355 -480 8360 -450
rect 8320 -485 8360 -480
rect 8320 -515 8360 -510
rect 8320 -545 8325 -515
rect 8325 -545 8355 -515
rect 8355 -545 8360 -515
rect 8320 -550 8360 -545
rect 8320 -575 8360 -570
rect 8320 -605 8325 -575
rect 8325 -605 8355 -575
rect 8355 -605 8360 -575
rect 8320 -610 8360 -605
rect 8320 -640 8360 -635
rect 8320 -670 8325 -640
rect 8325 -670 8355 -640
rect 8355 -670 8360 -640
rect 8320 -675 8360 -670
rect 8320 -710 8360 -705
rect 8320 -740 8325 -710
rect 8325 -740 8355 -710
rect 8355 -740 8360 -710
rect 8320 -745 8360 -740
rect 8320 -780 8360 -775
rect 8320 -810 8325 -780
rect 8325 -810 8355 -780
rect 8355 -810 8360 -780
rect 8320 -815 8360 -810
rect 8320 -850 8360 -845
rect 8320 -880 8325 -850
rect 8325 -880 8355 -850
rect 8355 -880 8360 -850
rect 8320 -885 8360 -880
rect 8320 -915 8360 -910
rect 8320 -945 8325 -915
rect 8325 -945 8355 -915
rect 8355 -945 8360 -915
rect 8320 -950 8360 -945
rect 8320 -975 8360 -970
rect 8320 -1005 8325 -975
rect 8325 -1005 8355 -975
rect 8355 -1005 8360 -975
rect 8320 -1010 8360 -1005
rect 8320 -1040 8360 -1035
rect 8320 -1070 8325 -1040
rect 8325 -1070 8355 -1040
rect 8355 -1070 8360 -1040
rect 8320 -1075 8360 -1070
rect 8320 -1110 8360 -1105
rect 8320 -1140 8325 -1110
rect 8325 -1140 8355 -1110
rect 8355 -1140 8360 -1110
rect 8320 -1145 8360 -1140
rect 8320 -1180 8360 -1175
rect 8320 -1210 8325 -1180
rect 8325 -1210 8355 -1180
rect 8355 -1210 8360 -1180
rect 8320 -1215 8360 -1210
rect 8320 -1250 8360 -1245
rect 8320 -1280 8325 -1250
rect 8325 -1280 8355 -1250
rect 8355 -1280 8360 -1250
rect 8320 -1285 8360 -1280
rect 8320 -1315 8360 -1310
rect 8320 -1345 8325 -1315
rect 8325 -1345 8355 -1315
rect 8355 -1345 8360 -1315
rect 8320 -1350 8360 -1345
rect 8670 225 8710 230
rect 8670 195 8675 225
rect 8675 195 8705 225
rect 8705 195 8710 225
rect 8670 190 8710 195
rect 8670 160 8710 165
rect 8670 130 8675 160
rect 8675 130 8705 160
rect 8705 130 8710 160
rect 8670 125 8710 130
rect 8670 90 8710 95
rect 8670 60 8675 90
rect 8675 60 8705 90
rect 8705 60 8710 90
rect 8670 55 8710 60
rect 8670 20 8710 25
rect 8670 -10 8675 20
rect 8675 -10 8705 20
rect 8705 -10 8710 20
rect 8670 -15 8710 -10
rect 8670 -50 8710 -45
rect 8670 -80 8675 -50
rect 8675 -80 8705 -50
rect 8705 -80 8710 -50
rect 8670 -85 8710 -80
rect 8670 -115 8710 -110
rect 8670 -145 8675 -115
rect 8675 -145 8705 -115
rect 8705 -145 8710 -115
rect 8670 -150 8710 -145
rect 8670 -175 8710 -170
rect 8670 -205 8675 -175
rect 8675 -205 8705 -175
rect 8705 -205 8710 -175
rect 8670 -210 8710 -205
rect 8670 -240 8710 -235
rect 8670 -270 8675 -240
rect 8675 -270 8705 -240
rect 8705 -270 8710 -240
rect 8670 -275 8710 -270
rect 8670 -310 8710 -305
rect 8670 -340 8675 -310
rect 8675 -340 8705 -310
rect 8705 -340 8710 -310
rect 8670 -345 8710 -340
rect 8670 -380 8710 -375
rect 8670 -410 8675 -380
rect 8675 -410 8705 -380
rect 8705 -410 8710 -380
rect 8670 -415 8710 -410
rect 8670 -450 8710 -445
rect 8670 -480 8675 -450
rect 8675 -480 8705 -450
rect 8705 -480 8710 -450
rect 8670 -485 8710 -480
rect 8670 -515 8710 -510
rect 8670 -545 8675 -515
rect 8675 -545 8705 -515
rect 8705 -545 8710 -515
rect 8670 -550 8710 -545
rect 8670 -575 8710 -570
rect 8670 -605 8675 -575
rect 8675 -605 8705 -575
rect 8705 -605 8710 -575
rect 8670 -610 8710 -605
rect 8670 -640 8710 -635
rect 8670 -670 8675 -640
rect 8675 -670 8705 -640
rect 8705 -670 8710 -640
rect 8670 -675 8710 -670
rect 8670 -710 8710 -705
rect 8670 -740 8675 -710
rect 8675 -740 8705 -710
rect 8705 -740 8710 -710
rect 8670 -745 8710 -740
rect 8670 -780 8710 -775
rect 8670 -810 8675 -780
rect 8675 -810 8705 -780
rect 8705 -810 8710 -780
rect 8670 -815 8710 -810
rect 8670 -850 8710 -845
rect 8670 -880 8675 -850
rect 8675 -880 8705 -850
rect 8705 -880 8710 -850
rect 8670 -885 8710 -880
rect 8670 -915 8710 -910
rect 8670 -945 8675 -915
rect 8675 -945 8705 -915
rect 8705 -945 8710 -915
rect 8670 -950 8710 -945
rect 8670 -975 8710 -970
rect 8670 -1005 8675 -975
rect 8675 -1005 8705 -975
rect 8705 -1005 8710 -975
rect 8670 -1010 8710 -1005
rect 8670 -1040 8710 -1035
rect 8670 -1070 8675 -1040
rect 8675 -1070 8705 -1040
rect 8705 -1070 8710 -1040
rect 8670 -1075 8710 -1070
rect 8670 -1110 8710 -1105
rect 8670 -1140 8675 -1110
rect 8675 -1140 8705 -1110
rect 8705 -1140 8710 -1110
rect 8670 -1145 8710 -1140
rect 8670 -1180 8710 -1175
rect 8670 -1210 8675 -1180
rect 8675 -1210 8705 -1180
rect 8705 -1210 8710 -1180
rect 8670 -1215 8710 -1210
rect 8670 -1250 8710 -1245
rect 8670 -1280 8675 -1250
rect 8675 -1280 8705 -1250
rect 8705 -1280 8710 -1250
rect 8670 -1285 8710 -1280
rect 8670 -1315 8710 -1310
rect 8670 -1345 8675 -1315
rect 8675 -1345 8705 -1315
rect 8705 -1345 8710 -1315
rect 8670 -1350 8710 -1345
rect 9020 225 9060 230
rect 9020 195 9025 225
rect 9025 195 9055 225
rect 9055 195 9060 225
rect 9020 190 9060 195
rect 9020 160 9060 165
rect 9020 130 9025 160
rect 9025 130 9055 160
rect 9055 130 9060 160
rect 9020 125 9060 130
rect 9020 90 9060 95
rect 9020 60 9025 90
rect 9025 60 9055 90
rect 9055 60 9060 90
rect 9020 55 9060 60
rect 9020 20 9060 25
rect 9020 -10 9025 20
rect 9025 -10 9055 20
rect 9055 -10 9060 20
rect 9020 -15 9060 -10
rect 9020 -50 9060 -45
rect 9020 -80 9025 -50
rect 9025 -80 9055 -50
rect 9055 -80 9060 -50
rect 9020 -85 9060 -80
rect 9020 -115 9060 -110
rect 9020 -145 9025 -115
rect 9025 -145 9055 -115
rect 9055 -145 9060 -115
rect 9020 -150 9060 -145
rect 9020 -175 9060 -170
rect 9020 -205 9025 -175
rect 9025 -205 9055 -175
rect 9055 -205 9060 -175
rect 9020 -210 9060 -205
rect 9020 -240 9060 -235
rect 9020 -270 9025 -240
rect 9025 -270 9055 -240
rect 9055 -270 9060 -240
rect 9020 -275 9060 -270
rect 9020 -310 9060 -305
rect 9020 -340 9025 -310
rect 9025 -340 9055 -310
rect 9055 -340 9060 -310
rect 9020 -345 9060 -340
rect 9020 -380 9060 -375
rect 9020 -410 9025 -380
rect 9025 -410 9055 -380
rect 9055 -410 9060 -380
rect 9020 -415 9060 -410
rect 9020 -450 9060 -445
rect 9020 -480 9025 -450
rect 9025 -480 9055 -450
rect 9055 -480 9060 -450
rect 9020 -485 9060 -480
rect 9020 -515 9060 -510
rect 9020 -545 9025 -515
rect 9025 -545 9055 -515
rect 9055 -545 9060 -515
rect 9020 -550 9060 -545
rect 9020 -575 9060 -570
rect 9020 -605 9025 -575
rect 9025 -605 9055 -575
rect 9055 -605 9060 -575
rect 9020 -610 9060 -605
rect 9020 -640 9060 -635
rect 9020 -670 9025 -640
rect 9025 -670 9055 -640
rect 9055 -670 9060 -640
rect 9020 -675 9060 -670
rect 9020 -710 9060 -705
rect 9020 -740 9025 -710
rect 9025 -740 9055 -710
rect 9055 -740 9060 -710
rect 9020 -745 9060 -740
rect 9020 -780 9060 -775
rect 9020 -810 9025 -780
rect 9025 -810 9055 -780
rect 9055 -810 9060 -780
rect 9020 -815 9060 -810
rect 9020 -850 9060 -845
rect 9020 -880 9025 -850
rect 9025 -880 9055 -850
rect 9055 -880 9060 -850
rect 9020 -885 9060 -880
rect 9020 -915 9060 -910
rect 9020 -945 9025 -915
rect 9025 -945 9055 -915
rect 9055 -945 9060 -915
rect 9020 -950 9060 -945
rect 9020 -975 9060 -970
rect 9020 -1005 9025 -975
rect 9025 -1005 9055 -975
rect 9055 -1005 9060 -975
rect 9020 -1010 9060 -1005
rect 9020 -1040 9060 -1035
rect 9020 -1070 9025 -1040
rect 9025 -1070 9055 -1040
rect 9055 -1070 9060 -1040
rect 9020 -1075 9060 -1070
rect 9020 -1110 9060 -1105
rect 9020 -1140 9025 -1110
rect 9025 -1140 9055 -1110
rect 9055 -1140 9060 -1110
rect 9020 -1145 9060 -1140
rect 9020 -1180 9060 -1175
rect 9020 -1210 9025 -1180
rect 9025 -1210 9055 -1180
rect 9055 -1210 9060 -1180
rect 9020 -1215 9060 -1210
rect 9020 -1250 9060 -1245
rect 9020 -1280 9025 -1250
rect 9025 -1280 9055 -1250
rect 9055 -1280 9060 -1250
rect 9020 -1285 9060 -1280
rect 9020 -1315 9060 -1310
rect 9020 -1345 9025 -1315
rect 9025 -1345 9055 -1315
rect 9055 -1345 9060 -1315
rect 9020 -1350 9060 -1345
rect 31305 185 31340 220
rect 31350 185 31385 220
rect 31395 185 31430 220
rect 31440 185 31475 220
rect 31485 185 31520 220
rect 31530 185 31565 220
rect 31575 185 31610 220
rect 31620 185 31655 220
rect 31665 185 31700 220
rect 31710 185 31745 220
rect 31755 185 31790 220
rect 31800 185 31835 220
rect 31845 185 31880 220
rect 31890 185 31925 220
rect 31935 185 31970 220
rect 31980 185 32015 220
rect 32025 185 32060 220
rect 32070 185 32105 220
rect 32115 185 32150 220
rect 32160 185 32195 220
rect 32205 185 32240 220
rect 32250 185 32285 220
rect 32295 185 32330 220
rect 32340 185 32375 220
rect 32385 185 32420 220
rect 32430 185 32465 220
rect 32475 185 32510 220
rect 32520 185 32555 220
rect 32565 185 32600 220
rect 32610 185 32645 220
rect 32655 185 32690 220
rect 32700 185 32735 220
rect 32745 185 32780 220
rect 32790 185 32825 220
rect 32835 185 32870 220
rect 31305 140 31340 175
rect 31350 140 31385 175
rect 31395 140 31430 175
rect 31440 140 31475 175
rect 31485 140 31520 175
rect 31530 140 31565 175
rect 31575 140 31610 175
rect 31620 140 31655 175
rect 31665 140 31700 175
rect 31710 140 31745 175
rect 31755 140 31790 175
rect 31800 140 31835 175
rect 31845 140 31880 175
rect 31890 140 31925 175
rect 31935 140 31970 175
rect 31980 140 32015 175
rect 32025 140 32060 175
rect 32070 140 32105 175
rect 32115 140 32150 175
rect 32160 140 32195 175
rect 32205 140 32240 175
rect 32250 140 32285 175
rect 32295 140 32330 175
rect 32340 140 32375 175
rect 32385 140 32420 175
rect 32430 140 32465 175
rect 32475 140 32510 175
rect 32520 140 32555 175
rect 32565 140 32600 175
rect 32610 140 32645 175
rect 32655 140 32690 175
rect 32700 140 32735 175
rect 32745 140 32780 175
rect 32790 140 32825 175
rect 32835 140 32870 175
rect 31305 95 31340 130
rect 31350 95 31385 130
rect 31395 95 31430 130
rect 31440 95 31475 130
rect 31485 95 31520 130
rect 31530 95 31565 130
rect 31575 95 31610 130
rect 31620 95 31655 130
rect 31665 95 31700 130
rect 31710 95 31745 130
rect 31755 95 31790 130
rect 31800 95 31835 130
rect 31845 95 31880 130
rect 31890 95 31925 130
rect 31935 95 31970 130
rect 31980 95 32015 130
rect 32025 95 32060 130
rect 32070 95 32105 130
rect 32115 95 32150 130
rect 32160 95 32195 130
rect 32205 95 32240 130
rect 32250 95 32285 130
rect 32295 95 32330 130
rect 32340 95 32375 130
rect 32385 95 32420 130
rect 32430 95 32465 130
rect 32475 95 32510 130
rect 32520 95 32555 130
rect 32565 95 32600 130
rect 32610 95 32645 130
rect 32655 95 32690 130
rect 32700 95 32735 130
rect 32745 95 32780 130
rect 32790 95 32825 130
rect 32835 95 32870 130
rect 31305 50 31340 85
rect 31350 50 31385 85
rect 31395 50 31430 85
rect 31440 50 31475 85
rect 31485 50 31520 85
rect 31530 50 31565 85
rect 31575 50 31610 85
rect 31620 50 31655 85
rect 31665 50 31700 85
rect 31710 50 31745 85
rect 31755 50 31790 85
rect 31800 50 31835 85
rect 31845 50 31880 85
rect 31890 50 31925 85
rect 31935 50 31970 85
rect 31980 50 32015 85
rect 32025 50 32060 85
rect 32070 50 32105 85
rect 32115 50 32150 85
rect 32160 50 32195 85
rect 32205 50 32240 85
rect 32250 50 32285 85
rect 32295 50 32330 85
rect 32340 50 32375 85
rect 32385 50 32420 85
rect 32430 50 32465 85
rect 32475 50 32510 85
rect 32520 50 32555 85
rect 32565 50 32600 85
rect 32610 50 32645 85
rect 32655 50 32690 85
rect 32700 50 32735 85
rect 32745 50 32780 85
rect 32790 50 32825 85
rect 32835 50 32870 85
rect 31305 5 31340 40
rect 31350 5 31385 40
rect 31395 5 31430 40
rect 31440 5 31475 40
rect 31485 5 31520 40
rect 31530 5 31565 40
rect 31575 5 31610 40
rect 31620 5 31655 40
rect 31665 5 31700 40
rect 31710 5 31745 40
rect 31755 5 31790 40
rect 31800 5 31835 40
rect 31845 5 31880 40
rect 31890 5 31925 40
rect 31935 5 31970 40
rect 31980 5 32015 40
rect 32025 5 32060 40
rect 32070 5 32105 40
rect 32115 5 32150 40
rect 32160 5 32195 40
rect 32205 5 32240 40
rect 32250 5 32285 40
rect 32295 5 32330 40
rect 32340 5 32375 40
rect 32385 5 32420 40
rect 32430 5 32465 40
rect 32475 5 32510 40
rect 32520 5 32555 40
rect 32565 5 32600 40
rect 32610 5 32645 40
rect 32655 5 32690 40
rect 32700 5 32735 40
rect 32745 5 32780 40
rect 32790 5 32825 40
rect 32835 5 32870 40
rect 31305 -40 31340 -5
rect 31350 -40 31385 -5
rect 31395 -40 31430 -5
rect 31440 -40 31475 -5
rect 31485 -40 31520 -5
rect 31530 -40 31565 -5
rect 31575 -40 31610 -5
rect 31620 -40 31655 -5
rect 31665 -40 31700 -5
rect 31710 -40 31745 -5
rect 31755 -40 31790 -5
rect 31800 -40 31835 -5
rect 31845 -40 31880 -5
rect 31890 -40 31925 -5
rect 31935 -40 31970 -5
rect 31980 -40 32015 -5
rect 32025 -40 32060 -5
rect 32070 -40 32105 -5
rect 32115 -40 32150 -5
rect 32160 -40 32195 -5
rect 32205 -40 32240 -5
rect 32250 -40 32285 -5
rect 32295 -40 32330 -5
rect 32340 -40 32375 -5
rect 32385 -40 32420 -5
rect 32430 -40 32465 -5
rect 32475 -40 32510 -5
rect 32520 -40 32555 -5
rect 32565 -40 32600 -5
rect 32610 -40 32645 -5
rect 32655 -40 32690 -5
rect 32700 -40 32735 -5
rect 32745 -40 32780 -5
rect 32790 -40 32825 -5
rect 32835 -40 32870 -5
rect 31305 -85 31340 -50
rect 31350 -85 31385 -50
rect 31395 -85 31430 -50
rect 31440 -85 31475 -50
rect 31485 -85 31520 -50
rect 31530 -85 31565 -50
rect 31575 -85 31610 -50
rect 31620 -85 31655 -50
rect 31665 -85 31700 -50
rect 31710 -85 31745 -50
rect 31755 -85 31790 -50
rect 31800 -85 31835 -50
rect 31845 -85 31880 -50
rect 31890 -85 31925 -50
rect 31935 -85 31970 -50
rect 31980 -85 32015 -50
rect 32025 -85 32060 -50
rect 32070 -85 32105 -50
rect 32115 -85 32150 -50
rect 32160 -85 32195 -50
rect 32205 -85 32240 -50
rect 32250 -85 32285 -50
rect 32295 -85 32330 -50
rect 32340 -85 32375 -50
rect 32385 -85 32420 -50
rect 32430 -85 32465 -50
rect 32475 -85 32510 -50
rect 32520 -85 32555 -50
rect 32565 -85 32600 -50
rect 32610 -85 32645 -50
rect 32655 -85 32690 -50
rect 32700 -85 32735 -50
rect 32745 -85 32780 -50
rect 32790 -85 32825 -50
rect 32835 -85 32870 -50
rect 31305 -130 31340 -95
rect 31350 -130 31385 -95
rect 31395 -130 31430 -95
rect 31440 -130 31475 -95
rect 31485 -130 31520 -95
rect 31530 -130 31565 -95
rect 31575 -130 31610 -95
rect 31620 -130 31655 -95
rect 31665 -130 31700 -95
rect 31710 -130 31745 -95
rect 31755 -130 31790 -95
rect 31800 -130 31835 -95
rect 31845 -130 31880 -95
rect 31890 -130 31925 -95
rect 31935 -130 31970 -95
rect 31980 -130 32015 -95
rect 32025 -130 32060 -95
rect 32070 -130 32105 -95
rect 32115 -130 32150 -95
rect 32160 -130 32195 -95
rect 32205 -130 32240 -95
rect 32250 -130 32285 -95
rect 32295 -130 32330 -95
rect 32340 -130 32375 -95
rect 32385 -130 32420 -95
rect 32430 -130 32465 -95
rect 32475 -130 32510 -95
rect 32520 -130 32555 -95
rect 32565 -130 32600 -95
rect 32610 -130 32645 -95
rect 32655 -130 32690 -95
rect 32700 -130 32735 -95
rect 32745 -130 32780 -95
rect 32790 -130 32825 -95
rect 32835 -130 32870 -95
rect 31305 -175 31340 -140
rect 31350 -175 31385 -140
rect 31395 -175 31430 -140
rect 31440 -175 31475 -140
rect 31485 -175 31520 -140
rect 31530 -175 31565 -140
rect 31575 -175 31610 -140
rect 31620 -175 31655 -140
rect 31665 -175 31700 -140
rect 31710 -175 31745 -140
rect 31755 -175 31790 -140
rect 31800 -175 31835 -140
rect 31845 -175 31880 -140
rect 31890 -175 31925 -140
rect 31935 -175 31970 -140
rect 31980 -175 32015 -140
rect 32025 -175 32060 -140
rect 32070 -175 32105 -140
rect 32115 -175 32150 -140
rect 32160 -175 32195 -140
rect 32205 -175 32240 -140
rect 32250 -175 32285 -140
rect 32295 -175 32330 -140
rect 32340 -175 32375 -140
rect 32385 -175 32420 -140
rect 32430 -175 32465 -140
rect 32475 -175 32510 -140
rect 32520 -175 32555 -140
rect 32565 -175 32600 -140
rect 32610 -175 32645 -140
rect 32655 -175 32690 -140
rect 32700 -175 32735 -140
rect 32745 -175 32780 -140
rect 32790 -175 32825 -140
rect 32835 -175 32870 -140
rect 31305 -220 31340 -185
rect 31350 -220 31385 -185
rect 31395 -220 31430 -185
rect 31440 -220 31475 -185
rect 31485 -220 31520 -185
rect 31530 -220 31565 -185
rect 31575 -220 31610 -185
rect 31620 -220 31655 -185
rect 31665 -220 31700 -185
rect 31710 -220 31745 -185
rect 31755 -220 31790 -185
rect 31800 -220 31835 -185
rect 31845 -220 31880 -185
rect 31890 -220 31925 -185
rect 31935 -220 31970 -185
rect 31980 -220 32015 -185
rect 32025 -220 32060 -185
rect 32070 -220 32105 -185
rect 32115 -220 32150 -185
rect 32160 -220 32195 -185
rect 32205 -220 32240 -185
rect 32250 -220 32285 -185
rect 32295 -220 32330 -185
rect 32340 -220 32375 -185
rect 32385 -220 32420 -185
rect 32430 -220 32465 -185
rect 32475 -220 32510 -185
rect 32520 -220 32555 -185
rect 32565 -220 32600 -185
rect 32610 -220 32645 -185
rect 32655 -220 32690 -185
rect 32700 -220 32735 -185
rect 32745 -220 32780 -185
rect 32790 -220 32825 -185
rect 32835 -220 32870 -185
rect 31305 -265 31340 -230
rect 31350 -265 31385 -230
rect 31395 -265 31430 -230
rect 31440 -265 31475 -230
rect 31485 -265 31520 -230
rect 31530 -265 31565 -230
rect 31575 -265 31610 -230
rect 31620 -265 31655 -230
rect 31665 -265 31700 -230
rect 31710 -265 31745 -230
rect 31755 -265 31790 -230
rect 31800 -265 31835 -230
rect 31845 -265 31880 -230
rect 31890 -265 31925 -230
rect 31935 -265 31970 -230
rect 31980 -265 32015 -230
rect 32025 -265 32060 -230
rect 32070 -265 32105 -230
rect 32115 -265 32150 -230
rect 32160 -265 32195 -230
rect 32205 -265 32240 -230
rect 32250 -265 32285 -230
rect 32295 -265 32330 -230
rect 32340 -265 32375 -230
rect 32385 -265 32420 -230
rect 32430 -265 32465 -230
rect 32475 -265 32510 -230
rect 32520 -265 32555 -230
rect 32565 -265 32600 -230
rect 32610 -265 32645 -230
rect 32655 -265 32690 -230
rect 32700 -265 32735 -230
rect 32745 -265 32780 -230
rect 32790 -265 32825 -230
rect 32835 -265 32870 -230
rect 31305 -310 31340 -275
rect 31350 -310 31385 -275
rect 31395 -310 31430 -275
rect 31440 -310 31475 -275
rect 31485 -310 31520 -275
rect 31530 -310 31565 -275
rect 31575 -310 31610 -275
rect 31620 -310 31655 -275
rect 31665 -310 31700 -275
rect 31710 -310 31745 -275
rect 31755 -310 31790 -275
rect 31800 -310 31835 -275
rect 31845 -310 31880 -275
rect 31890 -310 31925 -275
rect 31935 -310 31970 -275
rect 31980 -310 32015 -275
rect 32025 -310 32060 -275
rect 32070 -310 32105 -275
rect 32115 -310 32150 -275
rect 32160 -310 32195 -275
rect 32205 -310 32240 -275
rect 32250 -310 32285 -275
rect 32295 -310 32330 -275
rect 32340 -310 32375 -275
rect 32385 -310 32420 -275
rect 32430 -310 32465 -275
rect 32475 -310 32510 -275
rect 32520 -310 32555 -275
rect 32565 -310 32600 -275
rect 32610 -310 32645 -275
rect 32655 -310 32690 -275
rect 32700 -310 32735 -275
rect 32745 -310 32780 -275
rect 32790 -310 32825 -275
rect 32835 -310 32870 -275
rect 31305 -355 31340 -320
rect 31350 -355 31385 -320
rect 31395 -355 31430 -320
rect 31440 -355 31475 -320
rect 31485 -355 31520 -320
rect 31530 -355 31565 -320
rect 31575 -355 31610 -320
rect 31620 -355 31655 -320
rect 31665 -355 31700 -320
rect 31710 -355 31745 -320
rect 31755 -355 31790 -320
rect 31800 -355 31835 -320
rect 31845 -355 31880 -320
rect 31890 -355 31925 -320
rect 31935 -355 31970 -320
rect 31980 -355 32015 -320
rect 32025 -355 32060 -320
rect 32070 -355 32105 -320
rect 32115 -355 32150 -320
rect 32160 -355 32195 -320
rect 32205 -355 32240 -320
rect 32250 -355 32285 -320
rect 32295 -355 32330 -320
rect 32340 -355 32375 -320
rect 32385 -355 32420 -320
rect 32430 -355 32465 -320
rect 32475 -355 32510 -320
rect 32520 -355 32555 -320
rect 32565 -355 32600 -320
rect 32610 -355 32645 -320
rect 32655 -355 32690 -320
rect 32700 -355 32735 -320
rect 32745 -355 32780 -320
rect 32790 -355 32825 -320
rect 32835 -355 32870 -320
rect 31305 -400 31340 -365
rect 31350 -400 31385 -365
rect 31395 -400 31430 -365
rect 31440 -400 31475 -365
rect 31485 -400 31520 -365
rect 31530 -400 31565 -365
rect 31575 -400 31610 -365
rect 31620 -400 31655 -365
rect 31665 -400 31700 -365
rect 31710 -400 31745 -365
rect 31755 -400 31790 -365
rect 31800 -400 31835 -365
rect 31845 -400 31880 -365
rect 31890 -400 31925 -365
rect 31935 -400 31970 -365
rect 31980 -400 32015 -365
rect 32025 -400 32060 -365
rect 32070 -400 32105 -365
rect 32115 -400 32150 -365
rect 32160 -400 32195 -365
rect 32205 -400 32240 -365
rect 32250 -400 32285 -365
rect 32295 -400 32330 -365
rect 32340 -400 32375 -365
rect 32385 -400 32420 -365
rect 32430 -400 32465 -365
rect 32475 -400 32510 -365
rect 32520 -400 32555 -365
rect 32565 -400 32600 -365
rect 32610 -400 32645 -365
rect 32655 -400 32690 -365
rect 32700 -400 32735 -365
rect 32745 -400 32780 -365
rect 32790 -400 32825 -365
rect 32835 -400 32870 -365
rect 31305 -445 31340 -410
rect 31350 -445 31385 -410
rect 31395 -445 31430 -410
rect 31440 -445 31475 -410
rect 31485 -445 31520 -410
rect 31530 -445 31565 -410
rect 31575 -445 31610 -410
rect 31620 -445 31655 -410
rect 31665 -445 31700 -410
rect 31710 -445 31745 -410
rect 31755 -445 31790 -410
rect 31800 -445 31835 -410
rect 31845 -445 31880 -410
rect 31890 -445 31925 -410
rect 31935 -445 31970 -410
rect 31980 -445 32015 -410
rect 32025 -445 32060 -410
rect 32070 -445 32105 -410
rect 32115 -445 32150 -410
rect 32160 -445 32195 -410
rect 32205 -445 32240 -410
rect 32250 -445 32285 -410
rect 32295 -445 32330 -410
rect 32340 -445 32375 -410
rect 32385 -445 32420 -410
rect 32430 -445 32465 -410
rect 32475 -445 32510 -410
rect 32520 -445 32555 -410
rect 32565 -445 32600 -410
rect 32610 -445 32645 -410
rect 32655 -445 32690 -410
rect 32700 -445 32735 -410
rect 32745 -445 32780 -410
rect 32790 -445 32825 -410
rect 32835 -445 32870 -410
rect 31305 -490 31340 -455
rect 31350 -490 31385 -455
rect 31395 -490 31430 -455
rect 31440 -490 31475 -455
rect 31485 -490 31520 -455
rect 31530 -490 31565 -455
rect 31575 -490 31610 -455
rect 31620 -490 31655 -455
rect 31665 -490 31700 -455
rect 31710 -490 31745 -455
rect 31755 -490 31790 -455
rect 31800 -490 31835 -455
rect 31845 -490 31880 -455
rect 31890 -490 31925 -455
rect 31935 -490 31970 -455
rect 31980 -490 32015 -455
rect 32025 -490 32060 -455
rect 32070 -490 32105 -455
rect 32115 -490 32150 -455
rect 32160 -490 32195 -455
rect 32205 -490 32240 -455
rect 32250 -490 32285 -455
rect 32295 -490 32330 -455
rect 32340 -490 32375 -455
rect 32385 -490 32420 -455
rect 32430 -490 32465 -455
rect 32475 -490 32510 -455
rect 32520 -490 32555 -455
rect 32565 -490 32600 -455
rect 32610 -490 32645 -455
rect 32655 -490 32690 -455
rect 32700 -490 32735 -455
rect 32745 -490 32780 -455
rect 32790 -490 32825 -455
rect 32835 -490 32870 -455
rect 31305 -535 31340 -500
rect 31350 -535 31385 -500
rect 31395 -535 31430 -500
rect 31440 -535 31475 -500
rect 31485 -535 31520 -500
rect 31530 -535 31565 -500
rect 31575 -535 31610 -500
rect 31620 -535 31655 -500
rect 31665 -535 31700 -500
rect 31710 -535 31745 -500
rect 31755 -535 31790 -500
rect 31800 -535 31835 -500
rect 31845 -535 31880 -500
rect 31890 -535 31925 -500
rect 31935 -535 31970 -500
rect 31980 -535 32015 -500
rect 32025 -535 32060 -500
rect 32070 -535 32105 -500
rect 32115 -535 32150 -500
rect 32160 -535 32195 -500
rect 32205 -535 32240 -500
rect 32250 -535 32285 -500
rect 32295 -535 32330 -500
rect 32340 -535 32375 -500
rect 32385 -535 32420 -500
rect 32430 -535 32465 -500
rect 32475 -535 32510 -500
rect 32520 -535 32555 -500
rect 32565 -535 32600 -500
rect 32610 -535 32645 -500
rect 32655 -535 32690 -500
rect 32700 -535 32735 -500
rect 32745 -535 32780 -500
rect 32790 -535 32825 -500
rect 32835 -535 32870 -500
rect 31305 -580 31340 -545
rect 31350 -580 31385 -545
rect 31395 -580 31430 -545
rect 31440 -580 31475 -545
rect 31485 -580 31520 -545
rect 31530 -580 31565 -545
rect 31575 -580 31610 -545
rect 31620 -580 31655 -545
rect 31665 -580 31700 -545
rect 31710 -580 31745 -545
rect 31755 -580 31790 -545
rect 31800 -580 31835 -545
rect 31845 -580 31880 -545
rect 31890 -580 31925 -545
rect 31935 -580 31970 -545
rect 31980 -580 32015 -545
rect 32025 -580 32060 -545
rect 32070 -580 32105 -545
rect 32115 -580 32150 -545
rect 32160 -580 32195 -545
rect 32205 -580 32240 -545
rect 32250 -580 32285 -545
rect 32295 -580 32330 -545
rect 32340 -580 32375 -545
rect 32385 -580 32420 -545
rect 32430 -580 32465 -545
rect 32475 -580 32510 -545
rect 32520 -580 32555 -545
rect 32565 -580 32600 -545
rect 32610 -580 32645 -545
rect 32655 -580 32690 -545
rect 32700 -580 32735 -545
rect 32745 -580 32780 -545
rect 32790 -580 32825 -545
rect 32835 -580 32870 -545
rect 31305 -625 31340 -590
rect 31350 -625 31385 -590
rect 31395 -625 31430 -590
rect 31440 -625 31475 -590
rect 31485 -625 31520 -590
rect 31530 -625 31565 -590
rect 31575 -625 31610 -590
rect 31620 -625 31655 -590
rect 31665 -625 31700 -590
rect 31710 -625 31745 -590
rect 31755 -625 31790 -590
rect 31800 -625 31835 -590
rect 31845 -625 31880 -590
rect 31890 -625 31925 -590
rect 31935 -625 31970 -590
rect 31980 -625 32015 -590
rect 32025 -625 32060 -590
rect 32070 -625 32105 -590
rect 32115 -625 32150 -590
rect 32160 -625 32195 -590
rect 32205 -625 32240 -590
rect 32250 -625 32285 -590
rect 32295 -625 32330 -590
rect 32340 -625 32375 -590
rect 32385 -625 32420 -590
rect 32430 -625 32465 -590
rect 32475 -625 32510 -590
rect 32520 -625 32555 -590
rect 32565 -625 32600 -590
rect 32610 -625 32645 -590
rect 32655 -625 32690 -590
rect 32700 -625 32735 -590
rect 32745 -625 32780 -590
rect 32790 -625 32825 -590
rect 32835 -625 32870 -590
rect 31305 -670 31340 -635
rect 31350 -670 31385 -635
rect 31395 -670 31430 -635
rect 31440 -670 31475 -635
rect 31485 -670 31520 -635
rect 31530 -670 31565 -635
rect 31575 -670 31610 -635
rect 31620 -670 31655 -635
rect 31665 -670 31700 -635
rect 31710 -670 31745 -635
rect 31755 -670 31790 -635
rect 31800 -670 31835 -635
rect 31845 -670 31880 -635
rect 31890 -670 31925 -635
rect 31935 -670 31970 -635
rect 31980 -670 32015 -635
rect 32025 -670 32060 -635
rect 32070 -670 32105 -635
rect 32115 -670 32150 -635
rect 32160 -670 32195 -635
rect 32205 -670 32240 -635
rect 32250 -670 32285 -635
rect 32295 -670 32330 -635
rect 32340 -670 32375 -635
rect 32385 -670 32420 -635
rect 32430 -670 32465 -635
rect 32475 -670 32510 -635
rect 32520 -670 32555 -635
rect 32565 -670 32600 -635
rect 32610 -670 32645 -635
rect 32655 -670 32690 -635
rect 32700 -670 32735 -635
rect 32745 -670 32780 -635
rect 32790 -670 32825 -635
rect 32835 -670 32870 -635
rect 31305 -715 31340 -680
rect 31350 -715 31385 -680
rect 31395 -715 31430 -680
rect 31440 -715 31475 -680
rect 31485 -715 31520 -680
rect 31530 -715 31565 -680
rect 31575 -715 31610 -680
rect 31620 -715 31655 -680
rect 31665 -715 31700 -680
rect 31710 -715 31745 -680
rect 31755 -715 31790 -680
rect 31800 -715 31835 -680
rect 31845 -715 31880 -680
rect 31890 -715 31925 -680
rect 31935 -715 31970 -680
rect 31980 -715 32015 -680
rect 32025 -715 32060 -680
rect 32070 -715 32105 -680
rect 32115 -715 32150 -680
rect 32160 -715 32195 -680
rect 32205 -715 32240 -680
rect 32250 -715 32285 -680
rect 32295 -715 32330 -680
rect 32340 -715 32375 -680
rect 32385 -715 32420 -680
rect 32430 -715 32465 -680
rect 32475 -715 32510 -680
rect 32520 -715 32555 -680
rect 32565 -715 32600 -680
rect 32610 -715 32645 -680
rect 32655 -715 32690 -680
rect 32700 -715 32735 -680
rect 32745 -715 32780 -680
rect 32790 -715 32825 -680
rect 32835 -715 32870 -680
rect 31305 -760 31340 -725
rect 31350 -760 31385 -725
rect 31395 -760 31430 -725
rect 31440 -760 31475 -725
rect 31485 -760 31520 -725
rect 31530 -760 31565 -725
rect 31575 -760 31610 -725
rect 31620 -760 31655 -725
rect 31665 -760 31700 -725
rect 31710 -760 31745 -725
rect 31755 -760 31790 -725
rect 31800 -760 31835 -725
rect 31845 -760 31880 -725
rect 31890 -760 31925 -725
rect 31935 -760 31970 -725
rect 31980 -760 32015 -725
rect 32025 -760 32060 -725
rect 32070 -760 32105 -725
rect 32115 -760 32150 -725
rect 32160 -760 32195 -725
rect 32205 -760 32240 -725
rect 32250 -760 32285 -725
rect 32295 -760 32330 -725
rect 32340 -760 32375 -725
rect 32385 -760 32420 -725
rect 32430 -760 32465 -725
rect 32475 -760 32510 -725
rect 32520 -760 32555 -725
rect 32565 -760 32600 -725
rect 32610 -760 32645 -725
rect 32655 -760 32690 -725
rect 32700 -760 32735 -725
rect 32745 -760 32780 -725
rect 32790 -760 32825 -725
rect 32835 -760 32870 -725
rect 31305 -805 31340 -770
rect 31350 -805 31385 -770
rect 31395 -805 31430 -770
rect 31440 -805 31475 -770
rect 31485 -805 31520 -770
rect 31530 -805 31565 -770
rect 31575 -805 31610 -770
rect 31620 -805 31655 -770
rect 31665 -805 31700 -770
rect 31710 -805 31745 -770
rect 31755 -805 31790 -770
rect 31800 -805 31835 -770
rect 31845 -805 31880 -770
rect 31890 -805 31925 -770
rect 31935 -805 31970 -770
rect 31980 -805 32015 -770
rect 32025 -805 32060 -770
rect 32070 -805 32105 -770
rect 32115 -805 32150 -770
rect 32160 -805 32195 -770
rect 32205 -805 32240 -770
rect 32250 -805 32285 -770
rect 32295 -805 32330 -770
rect 32340 -805 32375 -770
rect 32385 -805 32420 -770
rect 32430 -805 32465 -770
rect 32475 -805 32510 -770
rect 32520 -805 32555 -770
rect 32565 -805 32600 -770
rect 32610 -805 32645 -770
rect 32655 -805 32690 -770
rect 32700 -805 32735 -770
rect 32745 -805 32780 -770
rect 32790 -805 32825 -770
rect 32835 -805 32870 -770
rect 31305 -850 31340 -815
rect 31350 -850 31385 -815
rect 31395 -850 31430 -815
rect 31440 -850 31475 -815
rect 31485 -850 31520 -815
rect 31530 -850 31565 -815
rect 31575 -850 31610 -815
rect 31620 -850 31655 -815
rect 31665 -850 31700 -815
rect 31710 -850 31745 -815
rect 31755 -850 31790 -815
rect 31800 -850 31835 -815
rect 31845 -850 31880 -815
rect 31890 -850 31925 -815
rect 31935 -850 31970 -815
rect 31980 -850 32015 -815
rect 32025 -850 32060 -815
rect 32070 -850 32105 -815
rect 32115 -850 32150 -815
rect 32160 -850 32195 -815
rect 32205 -850 32240 -815
rect 32250 -850 32285 -815
rect 32295 -850 32330 -815
rect 32340 -850 32375 -815
rect 32385 -850 32420 -815
rect 32430 -850 32465 -815
rect 32475 -850 32510 -815
rect 32520 -850 32555 -815
rect 32565 -850 32600 -815
rect 32610 -850 32645 -815
rect 32655 -850 32690 -815
rect 32700 -850 32735 -815
rect 32745 -850 32780 -815
rect 32790 -850 32825 -815
rect 32835 -850 32870 -815
rect 31305 -895 31340 -860
rect 31350 -895 31385 -860
rect 31395 -895 31430 -860
rect 31440 -895 31475 -860
rect 31485 -895 31520 -860
rect 31530 -895 31565 -860
rect 31575 -895 31610 -860
rect 31620 -895 31655 -860
rect 31665 -895 31700 -860
rect 31710 -895 31745 -860
rect 31755 -895 31790 -860
rect 31800 -895 31835 -860
rect 31845 -895 31880 -860
rect 31890 -895 31925 -860
rect 31935 -895 31970 -860
rect 31980 -895 32015 -860
rect 32025 -895 32060 -860
rect 32070 -895 32105 -860
rect 32115 -895 32150 -860
rect 32160 -895 32195 -860
rect 32205 -895 32240 -860
rect 32250 -895 32285 -860
rect 32295 -895 32330 -860
rect 32340 -895 32375 -860
rect 32385 -895 32420 -860
rect 32430 -895 32465 -860
rect 32475 -895 32510 -860
rect 32520 -895 32555 -860
rect 32565 -895 32600 -860
rect 32610 -895 32645 -860
rect 32655 -895 32690 -860
rect 32700 -895 32735 -860
rect 32745 -895 32780 -860
rect 32790 -895 32825 -860
rect 32835 -895 32870 -860
rect 31305 -940 31340 -905
rect 31350 -940 31385 -905
rect 31395 -940 31430 -905
rect 31440 -940 31475 -905
rect 31485 -940 31520 -905
rect 31530 -940 31565 -905
rect 31575 -940 31610 -905
rect 31620 -940 31655 -905
rect 31665 -940 31700 -905
rect 31710 -940 31745 -905
rect 31755 -940 31790 -905
rect 31800 -940 31835 -905
rect 31845 -940 31880 -905
rect 31890 -940 31925 -905
rect 31935 -940 31970 -905
rect 31980 -940 32015 -905
rect 32025 -940 32060 -905
rect 32070 -940 32105 -905
rect 32115 -940 32150 -905
rect 32160 -940 32195 -905
rect 32205 -940 32240 -905
rect 32250 -940 32285 -905
rect 32295 -940 32330 -905
rect 32340 -940 32375 -905
rect 32385 -940 32420 -905
rect 32430 -940 32465 -905
rect 32475 -940 32510 -905
rect 32520 -940 32555 -905
rect 32565 -940 32600 -905
rect 32610 -940 32645 -905
rect 32655 -940 32690 -905
rect 32700 -940 32735 -905
rect 32745 -940 32780 -905
rect 32790 -940 32825 -905
rect 32835 -940 32870 -905
rect 31305 -985 31340 -950
rect 31350 -985 31385 -950
rect 31395 -985 31430 -950
rect 31440 -985 31475 -950
rect 31485 -985 31520 -950
rect 31530 -985 31565 -950
rect 31575 -985 31610 -950
rect 31620 -985 31655 -950
rect 31665 -985 31700 -950
rect 31710 -985 31745 -950
rect 31755 -985 31790 -950
rect 31800 -985 31835 -950
rect 31845 -985 31880 -950
rect 31890 -985 31925 -950
rect 31935 -985 31970 -950
rect 31980 -985 32015 -950
rect 32025 -985 32060 -950
rect 32070 -985 32105 -950
rect 32115 -985 32150 -950
rect 32160 -985 32195 -950
rect 32205 -985 32240 -950
rect 32250 -985 32285 -950
rect 32295 -985 32330 -950
rect 32340 -985 32375 -950
rect 32385 -985 32420 -950
rect 32430 -985 32465 -950
rect 32475 -985 32510 -950
rect 32520 -985 32555 -950
rect 32565 -985 32600 -950
rect 32610 -985 32645 -950
rect 32655 -985 32690 -950
rect 32700 -985 32735 -950
rect 32745 -985 32780 -950
rect 32790 -985 32825 -950
rect 32835 -985 32870 -950
rect 31305 -1030 31340 -995
rect 31350 -1030 31385 -995
rect 31395 -1030 31430 -995
rect 31440 -1030 31475 -995
rect 31485 -1030 31520 -995
rect 31530 -1030 31565 -995
rect 31575 -1030 31610 -995
rect 31620 -1030 31655 -995
rect 31665 -1030 31700 -995
rect 31710 -1030 31745 -995
rect 31755 -1030 31790 -995
rect 31800 -1030 31835 -995
rect 31845 -1030 31880 -995
rect 31890 -1030 31925 -995
rect 31935 -1030 31970 -995
rect 31980 -1030 32015 -995
rect 32025 -1030 32060 -995
rect 32070 -1030 32105 -995
rect 32115 -1030 32150 -995
rect 32160 -1030 32195 -995
rect 32205 -1030 32240 -995
rect 32250 -1030 32285 -995
rect 32295 -1030 32330 -995
rect 32340 -1030 32375 -995
rect 32385 -1030 32420 -995
rect 32430 -1030 32465 -995
rect 32475 -1030 32510 -995
rect 32520 -1030 32555 -995
rect 32565 -1030 32600 -995
rect 32610 -1030 32645 -995
rect 32655 -1030 32690 -995
rect 32700 -1030 32735 -995
rect 32745 -1030 32780 -995
rect 32790 -1030 32825 -995
rect 32835 -1030 32870 -995
rect 31305 -1075 31340 -1040
rect 31350 -1075 31385 -1040
rect 31395 -1075 31430 -1040
rect 31440 -1075 31475 -1040
rect 31485 -1075 31520 -1040
rect 31530 -1075 31565 -1040
rect 31575 -1075 31610 -1040
rect 31620 -1075 31655 -1040
rect 31665 -1075 31700 -1040
rect 31710 -1075 31745 -1040
rect 31755 -1075 31790 -1040
rect 31800 -1075 31835 -1040
rect 31845 -1075 31880 -1040
rect 31890 -1075 31925 -1040
rect 31935 -1075 31970 -1040
rect 31980 -1075 32015 -1040
rect 32025 -1075 32060 -1040
rect 32070 -1075 32105 -1040
rect 32115 -1075 32150 -1040
rect 32160 -1075 32195 -1040
rect 32205 -1075 32240 -1040
rect 32250 -1075 32285 -1040
rect 32295 -1075 32330 -1040
rect 32340 -1075 32375 -1040
rect 32385 -1075 32420 -1040
rect 32430 -1075 32465 -1040
rect 32475 -1075 32510 -1040
rect 32520 -1075 32555 -1040
rect 32565 -1075 32600 -1040
rect 32610 -1075 32645 -1040
rect 32655 -1075 32690 -1040
rect 32700 -1075 32735 -1040
rect 32745 -1075 32780 -1040
rect 32790 -1075 32825 -1040
rect 32835 -1075 32870 -1040
rect 31305 -1120 31340 -1085
rect 31350 -1120 31385 -1085
rect 31395 -1120 31430 -1085
rect 31440 -1120 31475 -1085
rect 31485 -1120 31520 -1085
rect 31530 -1120 31565 -1085
rect 31575 -1120 31610 -1085
rect 31620 -1120 31655 -1085
rect 31665 -1120 31700 -1085
rect 31710 -1120 31745 -1085
rect 31755 -1120 31790 -1085
rect 31800 -1120 31835 -1085
rect 31845 -1120 31880 -1085
rect 31890 -1120 31925 -1085
rect 31935 -1120 31970 -1085
rect 31980 -1120 32015 -1085
rect 32025 -1120 32060 -1085
rect 32070 -1120 32105 -1085
rect 32115 -1120 32150 -1085
rect 32160 -1120 32195 -1085
rect 32205 -1120 32240 -1085
rect 32250 -1120 32285 -1085
rect 32295 -1120 32330 -1085
rect 32340 -1120 32375 -1085
rect 32385 -1120 32420 -1085
rect 32430 -1120 32465 -1085
rect 32475 -1120 32510 -1085
rect 32520 -1120 32555 -1085
rect 32565 -1120 32600 -1085
rect 32610 -1120 32645 -1085
rect 32655 -1120 32690 -1085
rect 32700 -1120 32735 -1085
rect 32745 -1120 32780 -1085
rect 32790 -1120 32825 -1085
rect 32835 -1120 32870 -1085
rect 31305 -1165 31340 -1130
rect 31350 -1165 31385 -1130
rect 31395 -1165 31430 -1130
rect 31440 -1165 31475 -1130
rect 31485 -1165 31520 -1130
rect 31530 -1165 31565 -1130
rect 31575 -1165 31610 -1130
rect 31620 -1165 31655 -1130
rect 31665 -1165 31700 -1130
rect 31710 -1165 31745 -1130
rect 31755 -1165 31790 -1130
rect 31800 -1165 31835 -1130
rect 31845 -1165 31880 -1130
rect 31890 -1165 31925 -1130
rect 31935 -1165 31970 -1130
rect 31980 -1165 32015 -1130
rect 32025 -1165 32060 -1130
rect 32070 -1165 32105 -1130
rect 32115 -1165 32150 -1130
rect 32160 -1165 32195 -1130
rect 32205 -1165 32240 -1130
rect 32250 -1165 32285 -1130
rect 32295 -1165 32330 -1130
rect 32340 -1165 32375 -1130
rect 32385 -1165 32420 -1130
rect 32430 -1165 32465 -1130
rect 32475 -1165 32510 -1130
rect 32520 -1165 32555 -1130
rect 32565 -1165 32600 -1130
rect 32610 -1165 32645 -1130
rect 32655 -1165 32690 -1130
rect 32700 -1165 32735 -1130
rect 32745 -1165 32780 -1130
rect 32790 -1165 32825 -1130
rect 32835 -1165 32870 -1130
rect 31305 -1210 31340 -1175
rect 31350 -1210 31385 -1175
rect 31395 -1210 31430 -1175
rect 31440 -1210 31475 -1175
rect 31485 -1210 31520 -1175
rect 31530 -1210 31565 -1175
rect 31575 -1210 31610 -1175
rect 31620 -1210 31655 -1175
rect 31665 -1210 31700 -1175
rect 31710 -1210 31745 -1175
rect 31755 -1210 31790 -1175
rect 31800 -1210 31835 -1175
rect 31845 -1210 31880 -1175
rect 31890 -1210 31925 -1175
rect 31935 -1210 31970 -1175
rect 31980 -1210 32015 -1175
rect 32025 -1210 32060 -1175
rect 32070 -1210 32105 -1175
rect 32115 -1210 32150 -1175
rect 32160 -1210 32195 -1175
rect 32205 -1210 32240 -1175
rect 32250 -1210 32285 -1175
rect 32295 -1210 32330 -1175
rect 32340 -1210 32375 -1175
rect 32385 -1210 32420 -1175
rect 32430 -1210 32465 -1175
rect 32475 -1210 32510 -1175
rect 32520 -1210 32555 -1175
rect 32565 -1210 32600 -1175
rect 32610 -1210 32645 -1175
rect 32655 -1210 32690 -1175
rect 32700 -1210 32735 -1175
rect 32745 -1210 32780 -1175
rect 32790 -1210 32825 -1175
rect 32835 -1210 32870 -1175
rect 31305 -1255 31340 -1220
rect 31350 -1255 31385 -1220
rect 31395 -1255 31430 -1220
rect 31440 -1255 31475 -1220
rect 31485 -1255 31520 -1220
rect 31530 -1255 31565 -1220
rect 31575 -1255 31610 -1220
rect 31620 -1255 31655 -1220
rect 31665 -1255 31700 -1220
rect 31710 -1255 31745 -1220
rect 31755 -1255 31790 -1220
rect 31800 -1255 31835 -1220
rect 31845 -1255 31880 -1220
rect 31890 -1255 31925 -1220
rect 31935 -1255 31970 -1220
rect 31980 -1255 32015 -1220
rect 32025 -1255 32060 -1220
rect 32070 -1255 32105 -1220
rect 32115 -1255 32150 -1220
rect 32160 -1255 32195 -1220
rect 32205 -1255 32240 -1220
rect 32250 -1255 32285 -1220
rect 32295 -1255 32330 -1220
rect 32340 -1255 32375 -1220
rect 32385 -1255 32420 -1220
rect 32430 -1255 32465 -1220
rect 32475 -1255 32510 -1220
rect 32520 -1255 32555 -1220
rect 32565 -1255 32600 -1220
rect 32610 -1255 32645 -1220
rect 32655 -1255 32690 -1220
rect 32700 -1255 32735 -1220
rect 32745 -1255 32780 -1220
rect 32790 -1255 32825 -1220
rect 32835 -1255 32870 -1220
rect 31305 -1300 31340 -1265
rect 31350 -1300 31385 -1265
rect 31395 -1300 31430 -1265
rect 31440 -1300 31475 -1265
rect 31485 -1300 31520 -1265
rect 31530 -1300 31565 -1265
rect 31575 -1300 31610 -1265
rect 31620 -1300 31655 -1265
rect 31665 -1300 31700 -1265
rect 31710 -1300 31745 -1265
rect 31755 -1300 31790 -1265
rect 31800 -1300 31835 -1265
rect 31845 -1300 31880 -1265
rect 31890 -1300 31925 -1265
rect 31935 -1300 31970 -1265
rect 31980 -1300 32015 -1265
rect 32025 -1300 32060 -1265
rect 32070 -1300 32105 -1265
rect 32115 -1300 32150 -1265
rect 32160 -1300 32195 -1265
rect 32205 -1300 32240 -1265
rect 32250 -1300 32285 -1265
rect 32295 -1300 32330 -1265
rect 32340 -1300 32375 -1265
rect 32385 -1300 32420 -1265
rect 32430 -1300 32465 -1265
rect 32475 -1300 32510 -1265
rect 32520 -1300 32555 -1265
rect 32565 -1300 32600 -1265
rect 32610 -1300 32645 -1265
rect 32655 -1300 32690 -1265
rect 32700 -1300 32735 -1265
rect 32745 -1300 32780 -1265
rect 32790 -1300 32825 -1265
rect 32835 -1300 32870 -1265
rect 31305 -1345 31340 -1310
rect 31350 -1345 31385 -1310
rect 31395 -1345 31430 -1310
rect 31440 -1345 31475 -1310
rect 31485 -1345 31520 -1310
rect 31530 -1345 31565 -1310
rect 31575 -1345 31610 -1310
rect 31620 -1345 31655 -1310
rect 31665 -1345 31700 -1310
rect 31710 -1345 31745 -1310
rect 31755 -1345 31790 -1310
rect 31800 -1345 31835 -1310
rect 31845 -1345 31880 -1310
rect 31890 -1345 31925 -1310
rect 31935 -1345 31970 -1310
rect 31980 -1345 32015 -1310
rect 32025 -1345 32060 -1310
rect 32070 -1345 32105 -1310
rect 32115 -1345 32150 -1310
rect 32160 -1345 32195 -1310
rect 32205 -1345 32240 -1310
rect 32250 -1345 32285 -1310
rect 32295 -1345 32330 -1310
rect 32340 -1345 32375 -1310
rect 32385 -1345 32420 -1310
rect 32430 -1345 32465 -1310
rect 32475 -1345 32510 -1310
rect 32520 -1345 32555 -1310
rect 32565 -1345 32600 -1310
rect 32610 -1345 32645 -1310
rect 32655 -1345 32690 -1310
rect 32700 -1345 32735 -1310
rect 32745 -1345 32780 -1310
rect 32790 -1345 32825 -1310
rect 32835 -1345 32870 -1310
<< metal4 >>
rect 2070 19315 32890 19325
rect 2070 19275 2110 19315
rect 2150 19275 6700 19315
rect 6740 19305 32890 19315
rect 6740 19275 31305 19305
rect 2070 19270 31305 19275
rect 31340 19270 31350 19305
rect 31385 19270 31395 19305
rect 31430 19270 31440 19305
rect 31475 19270 31485 19305
rect 31520 19270 31530 19305
rect 31565 19270 31575 19305
rect 31610 19270 31620 19305
rect 31655 19270 31665 19305
rect 31700 19270 31710 19305
rect 31745 19270 31755 19305
rect 31790 19270 31800 19305
rect 31835 19270 31845 19305
rect 31880 19270 31890 19305
rect 31925 19270 31935 19305
rect 31970 19270 31980 19305
rect 32015 19270 32025 19305
rect 32060 19270 32070 19305
rect 32105 19270 32115 19305
rect 32150 19270 32160 19305
rect 32195 19270 32205 19305
rect 32240 19270 32250 19305
rect 32285 19270 32295 19305
rect 32330 19270 32340 19305
rect 32375 19270 32385 19305
rect 32420 19270 32430 19305
rect 32465 19270 32475 19305
rect 32510 19270 32520 19305
rect 32555 19270 32565 19305
rect 32600 19270 32610 19305
rect 32645 19270 32655 19305
rect 32690 19270 32700 19305
rect 32735 19270 32745 19305
rect 32780 19270 32790 19305
rect 32825 19270 32835 19305
rect 32870 19270 32890 19305
rect 2070 19260 32890 19270
rect 2070 19250 31305 19260
rect 2070 19210 2110 19250
rect 2150 19210 6700 19250
rect 6740 19225 31305 19250
rect 31340 19225 31350 19260
rect 31385 19225 31395 19260
rect 31430 19225 31440 19260
rect 31475 19225 31485 19260
rect 31520 19225 31530 19260
rect 31565 19225 31575 19260
rect 31610 19225 31620 19260
rect 31655 19225 31665 19260
rect 31700 19225 31710 19260
rect 31745 19225 31755 19260
rect 31790 19225 31800 19260
rect 31835 19225 31845 19260
rect 31880 19225 31890 19260
rect 31925 19225 31935 19260
rect 31970 19225 31980 19260
rect 32015 19225 32025 19260
rect 32060 19225 32070 19260
rect 32105 19225 32115 19260
rect 32150 19225 32160 19260
rect 32195 19225 32205 19260
rect 32240 19225 32250 19260
rect 32285 19225 32295 19260
rect 32330 19225 32340 19260
rect 32375 19225 32385 19260
rect 32420 19225 32430 19260
rect 32465 19225 32475 19260
rect 32510 19225 32520 19260
rect 32555 19225 32565 19260
rect 32600 19225 32610 19260
rect 32645 19225 32655 19260
rect 32690 19225 32700 19260
rect 32735 19225 32745 19260
rect 32780 19225 32790 19260
rect 32825 19225 32835 19260
rect 32870 19225 32890 19260
rect 6740 19215 32890 19225
rect 6740 19210 31305 19215
rect 2070 19180 31305 19210
rect 31340 19180 31350 19215
rect 31385 19180 31395 19215
rect 31430 19180 31440 19215
rect 31475 19180 31485 19215
rect 31520 19180 31530 19215
rect 31565 19180 31575 19215
rect 31610 19180 31620 19215
rect 31655 19180 31665 19215
rect 31700 19180 31710 19215
rect 31745 19180 31755 19215
rect 31790 19180 31800 19215
rect 31835 19180 31845 19215
rect 31880 19180 31890 19215
rect 31925 19180 31935 19215
rect 31970 19180 31980 19215
rect 32015 19180 32025 19215
rect 32060 19180 32070 19215
rect 32105 19180 32115 19215
rect 32150 19180 32160 19215
rect 32195 19180 32205 19215
rect 32240 19180 32250 19215
rect 32285 19180 32295 19215
rect 32330 19180 32340 19215
rect 32375 19180 32385 19215
rect 32420 19180 32430 19215
rect 32465 19180 32475 19215
rect 32510 19180 32520 19215
rect 32555 19180 32565 19215
rect 32600 19180 32610 19215
rect 32645 19180 32655 19215
rect 32690 19180 32700 19215
rect 32735 19180 32745 19215
rect 32780 19180 32790 19215
rect 32825 19180 32835 19215
rect 32870 19180 32890 19215
rect 2070 19140 2110 19180
rect 2150 19140 6700 19180
rect 6740 19170 32890 19180
rect 6740 19140 31305 19170
rect 2070 19135 31305 19140
rect 31340 19135 31350 19170
rect 31385 19135 31395 19170
rect 31430 19135 31440 19170
rect 31475 19135 31485 19170
rect 31520 19135 31530 19170
rect 31565 19135 31575 19170
rect 31610 19135 31620 19170
rect 31655 19135 31665 19170
rect 31700 19135 31710 19170
rect 31745 19135 31755 19170
rect 31790 19135 31800 19170
rect 31835 19135 31845 19170
rect 31880 19135 31890 19170
rect 31925 19135 31935 19170
rect 31970 19135 31980 19170
rect 32015 19135 32025 19170
rect 32060 19135 32070 19170
rect 32105 19135 32115 19170
rect 32150 19135 32160 19170
rect 32195 19135 32205 19170
rect 32240 19135 32250 19170
rect 32285 19135 32295 19170
rect 32330 19135 32340 19170
rect 32375 19135 32385 19170
rect 32420 19135 32430 19170
rect 32465 19135 32475 19170
rect 32510 19135 32520 19170
rect 32555 19135 32565 19170
rect 32600 19135 32610 19170
rect 32645 19135 32655 19170
rect 32690 19135 32700 19170
rect 32735 19135 32745 19170
rect 32780 19135 32790 19170
rect 32825 19135 32835 19170
rect 32870 19135 32890 19170
rect 2070 19125 32890 19135
rect 2070 19110 31305 19125
rect 2070 19070 2110 19110
rect 2150 19070 6700 19110
rect 6740 19090 31305 19110
rect 31340 19090 31350 19125
rect 31385 19090 31395 19125
rect 31430 19090 31440 19125
rect 31475 19090 31485 19125
rect 31520 19090 31530 19125
rect 31565 19090 31575 19125
rect 31610 19090 31620 19125
rect 31655 19090 31665 19125
rect 31700 19090 31710 19125
rect 31745 19090 31755 19125
rect 31790 19090 31800 19125
rect 31835 19090 31845 19125
rect 31880 19090 31890 19125
rect 31925 19090 31935 19125
rect 31970 19090 31980 19125
rect 32015 19090 32025 19125
rect 32060 19090 32070 19125
rect 32105 19090 32115 19125
rect 32150 19090 32160 19125
rect 32195 19090 32205 19125
rect 32240 19090 32250 19125
rect 32285 19090 32295 19125
rect 32330 19090 32340 19125
rect 32375 19090 32385 19125
rect 32420 19090 32430 19125
rect 32465 19090 32475 19125
rect 32510 19090 32520 19125
rect 32555 19090 32565 19125
rect 32600 19090 32610 19125
rect 32645 19090 32655 19125
rect 32690 19090 32700 19125
rect 32735 19090 32745 19125
rect 32780 19090 32790 19125
rect 32825 19090 32835 19125
rect 32870 19090 32890 19125
rect 6740 19080 32890 19090
rect 6740 19070 31305 19080
rect 2070 19045 31305 19070
rect 31340 19045 31350 19080
rect 31385 19045 31395 19080
rect 31430 19045 31440 19080
rect 31475 19045 31485 19080
rect 31520 19045 31530 19080
rect 31565 19045 31575 19080
rect 31610 19045 31620 19080
rect 31655 19045 31665 19080
rect 31700 19045 31710 19080
rect 31745 19045 31755 19080
rect 31790 19045 31800 19080
rect 31835 19045 31845 19080
rect 31880 19045 31890 19080
rect 31925 19045 31935 19080
rect 31970 19045 31980 19080
rect 32015 19045 32025 19080
rect 32060 19045 32070 19080
rect 32105 19045 32115 19080
rect 32150 19045 32160 19080
rect 32195 19045 32205 19080
rect 32240 19045 32250 19080
rect 32285 19045 32295 19080
rect 32330 19045 32340 19080
rect 32375 19045 32385 19080
rect 32420 19045 32430 19080
rect 32465 19045 32475 19080
rect 32510 19045 32520 19080
rect 32555 19045 32565 19080
rect 32600 19045 32610 19080
rect 32645 19045 32655 19080
rect 32690 19045 32700 19080
rect 32735 19045 32745 19080
rect 32780 19045 32790 19080
rect 32825 19045 32835 19080
rect 32870 19045 32890 19080
rect 2070 19040 32890 19045
rect 2070 19000 2110 19040
rect 2150 19000 6700 19040
rect 6740 19035 32890 19040
rect 6740 19000 31305 19035
rect 31340 19000 31350 19035
rect 31385 19000 31395 19035
rect 31430 19000 31440 19035
rect 31475 19000 31485 19035
rect 31520 19000 31530 19035
rect 31565 19000 31575 19035
rect 31610 19000 31620 19035
rect 31655 19000 31665 19035
rect 31700 19000 31710 19035
rect 31745 19000 31755 19035
rect 31790 19000 31800 19035
rect 31835 19000 31845 19035
rect 31880 19000 31890 19035
rect 31925 19000 31935 19035
rect 31970 19000 31980 19035
rect 32015 19000 32025 19035
rect 32060 19000 32070 19035
rect 32105 19000 32115 19035
rect 32150 19000 32160 19035
rect 32195 19000 32205 19035
rect 32240 19000 32250 19035
rect 32285 19000 32295 19035
rect 32330 19000 32340 19035
rect 32375 19000 32385 19035
rect 32420 19000 32430 19035
rect 32465 19000 32475 19035
rect 32510 19000 32520 19035
rect 32555 19000 32565 19035
rect 32600 19000 32610 19035
rect 32645 19000 32655 19035
rect 32690 19000 32700 19035
rect 32735 19000 32745 19035
rect 32780 19000 32790 19035
rect 32825 19000 32835 19035
rect 32870 19000 32890 19035
rect 2070 18990 32890 19000
rect 2070 18975 31305 18990
rect 2070 18935 2110 18975
rect 2150 18935 6700 18975
rect 6740 18955 31305 18975
rect 31340 18955 31350 18990
rect 31385 18955 31395 18990
rect 31430 18955 31440 18990
rect 31475 18955 31485 18990
rect 31520 18955 31530 18990
rect 31565 18955 31575 18990
rect 31610 18955 31620 18990
rect 31655 18955 31665 18990
rect 31700 18955 31710 18990
rect 31745 18955 31755 18990
rect 31790 18955 31800 18990
rect 31835 18955 31845 18990
rect 31880 18955 31890 18990
rect 31925 18955 31935 18990
rect 31970 18955 31980 18990
rect 32015 18955 32025 18990
rect 32060 18955 32070 18990
rect 32105 18955 32115 18990
rect 32150 18955 32160 18990
rect 32195 18955 32205 18990
rect 32240 18955 32250 18990
rect 32285 18955 32295 18990
rect 32330 18955 32340 18990
rect 32375 18955 32385 18990
rect 32420 18955 32430 18990
rect 32465 18955 32475 18990
rect 32510 18955 32520 18990
rect 32555 18955 32565 18990
rect 32600 18955 32610 18990
rect 32645 18955 32655 18990
rect 32690 18955 32700 18990
rect 32735 18955 32745 18990
rect 32780 18955 32790 18990
rect 32825 18955 32835 18990
rect 32870 18955 32890 18990
rect 6740 18945 32890 18955
rect 6740 18935 31305 18945
rect 2070 18915 31305 18935
rect 2070 18875 2110 18915
rect 2150 18875 6700 18915
rect 6740 18910 31305 18915
rect 31340 18910 31350 18945
rect 31385 18910 31395 18945
rect 31430 18910 31440 18945
rect 31475 18910 31485 18945
rect 31520 18910 31530 18945
rect 31565 18910 31575 18945
rect 31610 18910 31620 18945
rect 31655 18910 31665 18945
rect 31700 18910 31710 18945
rect 31745 18910 31755 18945
rect 31790 18910 31800 18945
rect 31835 18910 31845 18945
rect 31880 18910 31890 18945
rect 31925 18910 31935 18945
rect 31970 18910 31980 18945
rect 32015 18910 32025 18945
rect 32060 18910 32070 18945
rect 32105 18910 32115 18945
rect 32150 18910 32160 18945
rect 32195 18910 32205 18945
rect 32240 18910 32250 18945
rect 32285 18910 32295 18945
rect 32330 18910 32340 18945
rect 32375 18910 32385 18945
rect 32420 18910 32430 18945
rect 32465 18910 32475 18945
rect 32510 18910 32520 18945
rect 32555 18910 32565 18945
rect 32600 18910 32610 18945
rect 32645 18910 32655 18945
rect 32690 18910 32700 18945
rect 32735 18910 32745 18945
rect 32780 18910 32790 18945
rect 32825 18910 32835 18945
rect 32870 18910 32890 18945
rect 6740 18900 32890 18910
rect 6740 18875 31305 18900
rect 2070 18865 31305 18875
rect 31340 18865 31350 18900
rect 31385 18865 31395 18900
rect 31430 18865 31440 18900
rect 31475 18865 31485 18900
rect 31520 18865 31530 18900
rect 31565 18865 31575 18900
rect 31610 18865 31620 18900
rect 31655 18865 31665 18900
rect 31700 18865 31710 18900
rect 31745 18865 31755 18900
rect 31790 18865 31800 18900
rect 31835 18865 31845 18900
rect 31880 18865 31890 18900
rect 31925 18865 31935 18900
rect 31970 18865 31980 18900
rect 32015 18865 32025 18900
rect 32060 18865 32070 18900
rect 32105 18865 32115 18900
rect 32150 18865 32160 18900
rect 32195 18865 32205 18900
rect 32240 18865 32250 18900
rect 32285 18865 32295 18900
rect 32330 18865 32340 18900
rect 32375 18865 32385 18900
rect 32420 18865 32430 18900
rect 32465 18865 32475 18900
rect 32510 18865 32520 18900
rect 32555 18865 32565 18900
rect 32600 18865 32610 18900
rect 32645 18865 32655 18900
rect 32690 18865 32700 18900
rect 32735 18865 32745 18900
rect 32780 18865 32790 18900
rect 32825 18865 32835 18900
rect 32870 18865 32890 18900
rect 2070 18855 32890 18865
rect 2070 18850 31305 18855
rect 2070 18810 2110 18850
rect 2150 18810 6700 18850
rect 6740 18820 31305 18850
rect 31340 18820 31350 18855
rect 31385 18820 31395 18855
rect 31430 18820 31440 18855
rect 31475 18820 31485 18855
rect 31520 18820 31530 18855
rect 31565 18820 31575 18855
rect 31610 18820 31620 18855
rect 31655 18820 31665 18855
rect 31700 18820 31710 18855
rect 31745 18820 31755 18855
rect 31790 18820 31800 18855
rect 31835 18820 31845 18855
rect 31880 18820 31890 18855
rect 31925 18820 31935 18855
rect 31970 18820 31980 18855
rect 32015 18820 32025 18855
rect 32060 18820 32070 18855
rect 32105 18820 32115 18855
rect 32150 18820 32160 18855
rect 32195 18820 32205 18855
rect 32240 18820 32250 18855
rect 32285 18820 32295 18855
rect 32330 18820 32340 18855
rect 32375 18820 32385 18855
rect 32420 18820 32430 18855
rect 32465 18820 32475 18855
rect 32510 18820 32520 18855
rect 32555 18820 32565 18855
rect 32600 18820 32610 18855
rect 32645 18820 32655 18855
rect 32690 18820 32700 18855
rect 32735 18820 32745 18855
rect 32780 18820 32790 18855
rect 32825 18820 32835 18855
rect 32870 18820 32890 18855
rect 6740 18810 32890 18820
rect 2070 18780 31305 18810
rect 2070 18740 2110 18780
rect 2150 18740 6700 18780
rect 6740 18775 31305 18780
rect 31340 18775 31350 18810
rect 31385 18775 31395 18810
rect 31430 18775 31440 18810
rect 31475 18775 31485 18810
rect 31520 18775 31530 18810
rect 31565 18775 31575 18810
rect 31610 18775 31620 18810
rect 31655 18775 31665 18810
rect 31700 18775 31710 18810
rect 31745 18775 31755 18810
rect 31790 18775 31800 18810
rect 31835 18775 31845 18810
rect 31880 18775 31890 18810
rect 31925 18775 31935 18810
rect 31970 18775 31980 18810
rect 32015 18775 32025 18810
rect 32060 18775 32070 18810
rect 32105 18775 32115 18810
rect 32150 18775 32160 18810
rect 32195 18775 32205 18810
rect 32240 18775 32250 18810
rect 32285 18775 32295 18810
rect 32330 18775 32340 18810
rect 32375 18775 32385 18810
rect 32420 18775 32430 18810
rect 32465 18775 32475 18810
rect 32510 18775 32520 18810
rect 32555 18775 32565 18810
rect 32600 18775 32610 18810
rect 32645 18775 32655 18810
rect 32690 18775 32700 18810
rect 32735 18775 32745 18810
rect 32780 18775 32790 18810
rect 32825 18775 32835 18810
rect 32870 18775 32890 18810
rect 6740 18765 32890 18775
rect 6740 18740 31305 18765
rect 2070 18730 31305 18740
rect 31340 18730 31350 18765
rect 31385 18730 31395 18765
rect 31430 18730 31440 18765
rect 31475 18730 31485 18765
rect 31520 18730 31530 18765
rect 31565 18730 31575 18765
rect 31610 18730 31620 18765
rect 31655 18730 31665 18765
rect 31700 18730 31710 18765
rect 31745 18730 31755 18765
rect 31790 18730 31800 18765
rect 31835 18730 31845 18765
rect 31880 18730 31890 18765
rect 31925 18730 31935 18765
rect 31970 18730 31980 18765
rect 32015 18730 32025 18765
rect 32060 18730 32070 18765
rect 32105 18730 32115 18765
rect 32150 18730 32160 18765
rect 32195 18730 32205 18765
rect 32240 18730 32250 18765
rect 32285 18730 32295 18765
rect 32330 18730 32340 18765
rect 32375 18730 32385 18765
rect 32420 18730 32430 18765
rect 32465 18730 32475 18765
rect 32510 18730 32520 18765
rect 32555 18730 32565 18765
rect 32600 18730 32610 18765
rect 32645 18730 32655 18765
rect 32690 18730 32700 18765
rect 32735 18730 32745 18765
rect 32780 18730 32790 18765
rect 32825 18730 32835 18765
rect 32870 18730 32890 18765
rect 2070 18720 32890 18730
rect 2070 18710 31305 18720
rect 2070 18670 2110 18710
rect 2150 18670 6700 18710
rect 6740 18685 31305 18710
rect 31340 18685 31350 18720
rect 31385 18685 31395 18720
rect 31430 18685 31440 18720
rect 31475 18685 31485 18720
rect 31520 18685 31530 18720
rect 31565 18685 31575 18720
rect 31610 18685 31620 18720
rect 31655 18685 31665 18720
rect 31700 18685 31710 18720
rect 31745 18685 31755 18720
rect 31790 18685 31800 18720
rect 31835 18685 31845 18720
rect 31880 18685 31890 18720
rect 31925 18685 31935 18720
rect 31970 18685 31980 18720
rect 32015 18685 32025 18720
rect 32060 18685 32070 18720
rect 32105 18685 32115 18720
rect 32150 18685 32160 18720
rect 32195 18685 32205 18720
rect 32240 18685 32250 18720
rect 32285 18685 32295 18720
rect 32330 18685 32340 18720
rect 32375 18685 32385 18720
rect 32420 18685 32430 18720
rect 32465 18685 32475 18720
rect 32510 18685 32520 18720
rect 32555 18685 32565 18720
rect 32600 18685 32610 18720
rect 32645 18685 32655 18720
rect 32690 18685 32700 18720
rect 32735 18685 32745 18720
rect 32780 18685 32790 18720
rect 32825 18685 32835 18720
rect 32870 18685 32890 18720
rect 6740 18675 32890 18685
rect 6740 18670 31305 18675
rect 2070 18640 31305 18670
rect 31340 18640 31350 18675
rect 31385 18640 31395 18675
rect 31430 18640 31440 18675
rect 31475 18640 31485 18675
rect 31520 18640 31530 18675
rect 31565 18640 31575 18675
rect 31610 18640 31620 18675
rect 31655 18640 31665 18675
rect 31700 18640 31710 18675
rect 31745 18640 31755 18675
rect 31790 18640 31800 18675
rect 31835 18640 31845 18675
rect 31880 18640 31890 18675
rect 31925 18640 31935 18675
rect 31970 18640 31980 18675
rect 32015 18640 32025 18675
rect 32060 18640 32070 18675
rect 32105 18640 32115 18675
rect 32150 18640 32160 18675
rect 32195 18640 32205 18675
rect 32240 18640 32250 18675
rect 32285 18640 32295 18675
rect 32330 18640 32340 18675
rect 32375 18640 32385 18675
rect 32420 18640 32430 18675
rect 32465 18640 32475 18675
rect 32510 18640 32520 18675
rect 32555 18640 32565 18675
rect 32600 18640 32610 18675
rect 32645 18640 32655 18675
rect 32690 18640 32700 18675
rect 32735 18640 32745 18675
rect 32780 18640 32790 18675
rect 32825 18640 32835 18675
rect 32870 18640 32890 18675
rect 2070 18600 2110 18640
rect 2150 18600 6700 18640
rect 6740 18630 32890 18640
rect 6740 18600 31305 18630
rect 2070 18595 31305 18600
rect 31340 18595 31350 18630
rect 31385 18595 31395 18630
rect 31430 18595 31440 18630
rect 31475 18595 31485 18630
rect 31520 18595 31530 18630
rect 31565 18595 31575 18630
rect 31610 18595 31620 18630
rect 31655 18595 31665 18630
rect 31700 18595 31710 18630
rect 31745 18595 31755 18630
rect 31790 18595 31800 18630
rect 31835 18595 31845 18630
rect 31880 18595 31890 18630
rect 31925 18595 31935 18630
rect 31970 18595 31980 18630
rect 32015 18595 32025 18630
rect 32060 18595 32070 18630
rect 32105 18595 32115 18630
rect 32150 18595 32160 18630
rect 32195 18595 32205 18630
rect 32240 18595 32250 18630
rect 32285 18595 32295 18630
rect 32330 18595 32340 18630
rect 32375 18595 32385 18630
rect 32420 18595 32430 18630
rect 32465 18595 32475 18630
rect 32510 18595 32520 18630
rect 32555 18595 32565 18630
rect 32600 18595 32610 18630
rect 32645 18595 32655 18630
rect 32690 18595 32700 18630
rect 32735 18595 32745 18630
rect 32780 18595 32790 18630
rect 32825 18595 32835 18630
rect 32870 18595 32890 18630
rect 2070 18585 32890 18595
rect 2070 18575 31305 18585
rect 2070 18535 2110 18575
rect 2150 18535 6700 18575
rect 6740 18550 31305 18575
rect 31340 18550 31350 18585
rect 31385 18550 31395 18585
rect 31430 18550 31440 18585
rect 31475 18550 31485 18585
rect 31520 18550 31530 18585
rect 31565 18550 31575 18585
rect 31610 18550 31620 18585
rect 31655 18550 31665 18585
rect 31700 18550 31710 18585
rect 31745 18550 31755 18585
rect 31790 18550 31800 18585
rect 31835 18550 31845 18585
rect 31880 18550 31890 18585
rect 31925 18550 31935 18585
rect 31970 18550 31980 18585
rect 32015 18550 32025 18585
rect 32060 18550 32070 18585
rect 32105 18550 32115 18585
rect 32150 18550 32160 18585
rect 32195 18550 32205 18585
rect 32240 18550 32250 18585
rect 32285 18550 32295 18585
rect 32330 18550 32340 18585
rect 32375 18550 32385 18585
rect 32420 18550 32430 18585
rect 32465 18550 32475 18585
rect 32510 18550 32520 18585
rect 32555 18550 32565 18585
rect 32600 18550 32610 18585
rect 32645 18550 32655 18585
rect 32690 18550 32700 18585
rect 32735 18550 32745 18585
rect 32780 18550 32790 18585
rect 32825 18550 32835 18585
rect 32870 18550 32890 18585
rect 6740 18540 32890 18550
rect 6740 18535 31305 18540
rect 2070 18515 31305 18535
rect 2070 18475 2110 18515
rect 2150 18475 6700 18515
rect 6740 18505 31305 18515
rect 31340 18505 31350 18540
rect 31385 18505 31395 18540
rect 31430 18505 31440 18540
rect 31475 18505 31485 18540
rect 31520 18505 31530 18540
rect 31565 18505 31575 18540
rect 31610 18505 31620 18540
rect 31655 18505 31665 18540
rect 31700 18505 31710 18540
rect 31745 18505 31755 18540
rect 31790 18505 31800 18540
rect 31835 18505 31845 18540
rect 31880 18505 31890 18540
rect 31925 18505 31935 18540
rect 31970 18505 31980 18540
rect 32015 18505 32025 18540
rect 32060 18505 32070 18540
rect 32105 18505 32115 18540
rect 32150 18505 32160 18540
rect 32195 18505 32205 18540
rect 32240 18505 32250 18540
rect 32285 18505 32295 18540
rect 32330 18505 32340 18540
rect 32375 18505 32385 18540
rect 32420 18505 32430 18540
rect 32465 18505 32475 18540
rect 32510 18505 32520 18540
rect 32555 18505 32565 18540
rect 32600 18505 32610 18540
rect 32645 18505 32655 18540
rect 32690 18505 32700 18540
rect 32735 18505 32745 18540
rect 32780 18505 32790 18540
rect 32825 18505 32835 18540
rect 32870 18505 32890 18540
rect 6740 18495 32890 18505
rect 6740 18475 31305 18495
rect 2070 18460 31305 18475
rect 31340 18460 31350 18495
rect 31385 18460 31395 18495
rect 31430 18460 31440 18495
rect 31475 18460 31485 18495
rect 31520 18460 31530 18495
rect 31565 18460 31575 18495
rect 31610 18460 31620 18495
rect 31655 18460 31665 18495
rect 31700 18460 31710 18495
rect 31745 18460 31755 18495
rect 31790 18460 31800 18495
rect 31835 18460 31845 18495
rect 31880 18460 31890 18495
rect 31925 18460 31935 18495
rect 31970 18460 31980 18495
rect 32015 18460 32025 18495
rect 32060 18460 32070 18495
rect 32105 18460 32115 18495
rect 32150 18460 32160 18495
rect 32195 18460 32205 18495
rect 32240 18460 32250 18495
rect 32285 18460 32295 18495
rect 32330 18460 32340 18495
rect 32375 18460 32385 18495
rect 32420 18460 32430 18495
rect 32465 18460 32475 18495
rect 32510 18460 32520 18495
rect 32555 18460 32565 18495
rect 32600 18460 32610 18495
rect 32645 18460 32655 18495
rect 32690 18460 32700 18495
rect 32735 18460 32745 18495
rect 32780 18460 32790 18495
rect 32825 18460 32835 18495
rect 32870 18460 32890 18495
rect 2070 18450 32890 18460
rect 2070 18410 2110 18450
rect 2150 18410 6700 18450
rect 6740 18415 31305 18450
rect 31340 18415 31350 18450
rect 31385 18415 31395 18450
rect 31430 18415 31440 18450
rect 31475 18415 31485 18450
rect 31520 18415 31530 18450
rect 31565 18415 31575 18450
rect 31610 18415 31620 18450
rect 31655 18415 31665 18450
rect 31700 18415 31710 18450
rect 31745 18415 31755 18450
rect 31790 18415 31800 18450
rect 31835 18415 31845 18450
rect 31880 18415 31890 18450
rect 31925 18415 31935 18450
rect 31970 18415 31980 18450
rect 32015 18415 32025 18450
rect 32060 18415 32070 18450
rect 32105 18415 32115 18450
rect 32150 18415 32160 18450
rect 32195 18415 32205 18450
rect 32240 18415 32250 18450
rect 32285 18415 32295 18450
rect 32330 18415 32340 18450
rect 32375 18415 32385 18450
rect 32420 18415 32430 18450
rect 32465 18415 32475 18450
rect 32510 18415 32520 18450
rect 32555 18415 32565 18450
rect 32600 18415 32610 18450
rect 32645 18415 32655 18450
rect 32690 18415 32700 18450
rect 32735 18415 32745 18450
rect 32780 18415 32790 18450
rect 32825 18415 32835 18450
rect 32870 18415 32890 18450
rect 6740 18410 32890 18415
rect 2070 18405 32890 18410
rect 2070 18380 31305 18405
rect 2070 18340 2110 18380
rect 2150 18340 6700 18380
rect 6740 18370 31305 18380
rect 31340 18370 31350 18405
rect 31385 18370 31395 18405
rect 31430 18370 31440 18405
rect 31475 18370 31485 18405
rect 31520 18370 31530 18405
rect 31565 18370 31575 18405
rect 31610 18370 31620 18405
rect 31655 18370 31665 18405
rect 31700 18370 31710 18405
rect 31745 18370 31755 18405
rect 31790 18370 31800 18405
rect 31835 18370 31845 18405
rect 31880 18370 31890 18405
rect 31925 18370 31935 18405
rect 31970 18370 31980 18405
rect 32015 18370 32025 18405
rect 32060 18370 32070 18405
rect 32105 18370 32115 18405
rect 32150 18370 32160 18405
rect 32195 18370 32205 18405
rect 32240 18370 32250 18405
rect 32285 18370 32295 18405
rect 32330 18370 32340 18405
rect 32375 18370 32385 18405
rect 32420 18370 32430 18405
rect 32465 18370 32475 18405
rect 32510 18370 32520 18405
rect 32555 18370 32565 18405
rect 32600 18370 32610 18405
rect 32645 18370 32655 18405
rect 32690 18370 32700 18405
rect 32735 18370 32745 18405
rect 32780 18370 32790 18405
rect 32825 18370 32835 18405
rect 32870 18370 32890 18405
rect 6740 18360 32890 18370
rect 6740 18340 31305 18360
rect 2070 18325 31305 18340
rect 31340 18325 31350 18360
rect 31385 18325 31395 18360
rect 31430 18325 31440 18360
rect 31475 18325 31485 18360
rect 31520 18325 31530 18360
rect 31565 18325 31575 18360
rect 31610 18325 31620 18360
rect 31655 18325 31665 18360
rect 31700 18325 31710 18360
rect 31745 18325 31755 18360
rect 31790 18325 31800 18360
rect 31835 18325 31845 18360
rect 31880 18325 31890 18360
rect 31925 18325 31935 18360
rect 31970 18325 31980 18360
rect 32015 18325 32025 18360
rect 32060 18325 32070 18360
rect 32105 18325 32115 18360
rect 32150 18325 32160 18360
rect 32195 18325 32205 18360
rect 32240 18325 32250 18360
rect 32285 18325 32295 18360
rect 32330 18325 32340 18360
rect 32375 18325 32385 18360
rect 32420 18325 32430 18360
rect 32465 18325 32475 18360
rect 32510 18325 32520 18360
rect 32555 18325 32565 18360
rect 32600 18325 32610 18360
rect 32645 18325 32655 18360
rect 32690 18325 32700 18360
rect 32735 18325 32745 18360
rect 32780 18325 32790 18360
rect 32825 18325 32835 18360
rect 32870 18325 32890 18360
rect 2070 18315 32890 18325
rect 2070 18310 31305 18315
rect 2070 18270 2110 18310
rect 2150 18270 6700 18310
rect 6740 18280 31305 18310
rect 31340 18280 31350 18315
rect 31385 18280 31395 18315
rect 31430 18280 31440 18315
rect 31475 18280 31485 18315
rect 31520 18280 31530 18315
rect 31565 18280 31575 18315
rect 31610 18280 31620 18315
rect 31655 18280 31665 18315
rect 31700 18280 31710 18315
rect 31745 18280 31755 18315
rect 31790 18280 31800 18315
rect 31835 18280 31845 18315
rect 31880 18280 31890 18315
rect 31925 18280 31935 18315
rect 31970 18280 31980 18315
rect 32015 18280 32025 18315
rect 32060 18280 32070 18315
rect 32105 18280 32115 18315
rect 32150 18280 32160 18315
rect 32195 18280 32205 18315
rect 32240 18280 32250 18315
rect 32285 18280 32295 18315
rect 32330 18280 32340 18315
rect 32375 18280 32385 18315
rect 32420 18280 32430 18315
rect 32465 18280 32475 18315
rect 32510 18280 32520 18315
rect 32555 18280 32565 18315
rect 32600 18280 32610 18315
rect 32645 18280 32655 18315
rect 32690 18280 32700 18315
rect 32735 18280 32745 18315
rect 32780 18280 32790 18315
rect 32825 18280 32835 18315
rect 32870 18280 32890 18315
rect 6740 18270 32890 18280
rect 2070 18240 31305 18270
rect 2070 18200 2110 18240
rect 2150 18200 6700 18240
rect 6740 18235 31305 18240
rect 31340 18235 31350 18270
rect 31385 18235 31395 18270
rect 31430 18235 31440 18270
rect 31475 18235 31485 18270
rect 31520 18235 31530 18270
rect 31565 18235 31575 18270
rect 31610 18235 31620 18270
rect 31655 18235 31665 18270
rect 31700 18235 31710 18270
rect 31745 18235 31755 18270
rect 31790 18235 31800 18270
rect 31835 18235 31845 18270
rect 31880 18235 31890 18270
rect 31925 18235 31935 18270
rect 31970 18235 31980 18270
rect 32015 18235 32025 18270
rect 32060 18235 32070 18270
rect 32105 18235 32115 18270
rect 32150 18235 32160 18270
rect 32195 18235 32205 18270
rect 32240 18235 32250 18270
rect 32285 18235 32295 18270
rect 32330 18235 32340 18270
rect 32375 18235 32385 18270
rect 32420 18235 32430 18270
rect 32465 18235 32475 18270
rect 32510 18235 32520 18270
rect 32555 18235 32565 18270
rect 32600 18235 32610 18270
rect 32645 18235 32655 18270
rect 32690 18235 32700 18270
rect 32735 18235 32745 18270
rect 32780 18235 32790 18270
rect 32825 18235 32835 18270
rect 32870 18235 32890 18270
rect 6740 18225 32890 18235
rect 6740 18200 31305 18225
rect 2070 18190 31305 18200
rect 31340 18190 31350 18225
rect 31385 18190 31395 18225
rect 31430 18190 31440 18225
rect 31475 18190 31485 18225
rect 31520 18190 31530 18225
rect 31565 18190 31575 18225
rect 31610 18190 31620 18225
rect 31655 18190 31665 18225
rect 31700 18190 31710 18225
rect 31745 18190 31755 18225
rect 31790 18190 31800 18225
rect 31835 18190 31845 18225
rect 31880 18190 31890 18225
rect 31925 18190 31935 18225
rect 31970 18190 31980 18225
rect 32015 18190 32025 18225
rect 32060 18190 32070 18225
rect 32105 18190 32115 18225
rect 32150 18190 32160 18225
rect 32195 18190 32205 18225
rect 32240 18190 32250 18225
rect 32285 18190 32295 18225
rect 32330 18190 32340 18225
rect 32375 18190 32385 18225
rect 32420 18190 32430 18225
rect 32465 18190 32475 18225
rect 32510 18190 32520 18225
rect 32555 18190 32565 18225
rect 32600 18190 32610 18225
rect 32645 18190 32655 18225
rect 32690 18190 32700 18225
rect 32735 18190 32745 18225
rect 32780 18190 32790 18225
rect 32825 18190 32835 18225
rect 32870 18190 32890 18225
rect 2070 18180 32890 18190
rect 2070 18175 31305 18180
rect 2070 18135 2110 18175
rect 2150 18135 6700 18175
rect 6740 18145 31305 18175
rect 31340 18145 31350 18180
rect 31385 18145 31395 18180
rect 31430 18145 31440 18180
rect 31475 18145 31485 18180
rect 31520 18145 31530 18180
rect 31565 18145 31575 18180
rect 31610 18145 31620 18180
rect 31655 18145 31665 18180
rect 31700 18145 31710 18180
rect 31745 18145 31755 18180
rect 31790 18145 31800 18180
rect 31835 18145 31845 18180
rect 31880 18145 31890 18180
rect 31925 18145 31935 18180
rect 31970 18145 31980 18180
rect 32015 18145 32025 18180
rect 32060 18145 32070 18180
rect 32105 18145 32115 18180
rect 32150 18145 32160 18180
rect 32195 18145 32205 18180
rect 32240 18145 32250 18180
rect 32285 18145 32295 18180
rect 32330 18145 32340 18180
rect 32375 18145 32385 18180
rect 32420 18145 32430 18180
rect 32465 18145 32475 18180
rect 32510 18145 32520 18180
rect 32555 18145 32565 18180
rect 32600 18145 32610 18180
rect 32645 18145 32655 18180
rect 32690 18145 32700 18180
rect 32735 18145 32745 18180
rect 32780 18145 32790 18180
rect 32825 18145 32835 18180
rect 32870 18145 32890 18180
rect 6740 18135 32890 18145
rect 2070 18115 31305 18135
rect 2070 18075 2110 18115
rect 2150 18075 6700 18115
rect 6740 18100 31305 18115
rect 31340 18100 31350 18135
rect 31385 18100 31395 18135
rect 31430 18100 31440 18135
rect 31475 18100 31485 18135
rect 31520 18100 31530 18135
rect 31565 18100 31575 18135
rect 31610 18100 31620 18135
rect 31655 18100 31665 18135
rect 31700 18100 31710 18135
rect 31745 18100 31755 18135
rect 31790 18100 31800 18135
rect 31835 18100 31845 18135
rect 31880 18100 31890 18135
rect 31925 18100 31935 18135
rect 31970 18100 31980 18135
rect 32015 18100 32025 18135
rect 32060 18100 32070 18135
rect 32105 18100 32115 18135
rect 32150 18100 32160 18135
rect 32195 18100 32205 18135
rect 32240 18100 32250 18135
rect 32285 18100 32295 18135
rect 32330 18100 32340 18135
rect 32375 18100 32385 18135
rect 32420 18100 32430 18135
rect 32465 18100 32475 18135
rect 32510 18100 32520 18135
rect 32555 18100 32565 18135
rect 32600 18100 32610 18135
rect 32645 18100 32655 18135
rect 32690 18100 32700 18135
rect 32735 18100 32745 18135
rect 32780 18100 32790 18135
rect 32825 18100 32835 18135
rect 32870 18100 32890 18135
rect 6740 18090 32890 18100
rect 6740 18075 31305 18090
rect 2070 18055 31305 18075
rect 31340 18055 31350 18090
rect 31385 18055 31395 18090
rect 31430 18055 31440 18090
rect 31475 18055 31485 18090
rect 31520 18055 31530 18090
rect 31565 18055 31575 18090
rect 31610 18055 31620 18090
rect 31655 18055 31665 18090
rect 31700 18055 31710 18090
rect 31745 18055 31755 18090
rect 31790 18055 31800 18090
rect 31835 18055 31845 18090
rect 31880 18055 31890 18090
rect 31925 18055 31935 18090
rect 31970 18055 31980 18090
rect 32015 18055 32025 18090
rect 32060 18055 32070 18090
rect 32105 18055 32115 18090
rect 32150 18055 32160 18090
rect 32195 18055 32205 18090
rect 32240 18055 32250 18090
rect 32285 18055 32295 18090
rect 32330 18055 32340 18090
rect 32375 18055 32385 18090
rect 32420 18055 32430 18090
rect 32465 18055 32475 18090
rect 32510 18055 32520 18090
rect 32555 18055 32565 18090
rect 32600 18055 32610 18090
rect 32645 18055 32655 18090
rect 32690 18055 32700 18090
rect 32735 18055 32745 18090
rect 32780 18055 32790 18090
rect 32825 18055 32835 18090
rect 32870 18055 32890 18090
rect 2070 18050 32890 18055
rect 2070 18010 2110 18050
rect 2150 18010 6700 18050
rect 6740 18045 32890 18050
rect 6740 18010 31305 18045
rect 31340 18010 31350 18045
rect 31385 18010 31395 18045
rect 31430 18010 31440 18045
rect 31475 18010 31485 18045
rect 31520 18010 31530 18045
rect 31565 18010 31575 18045
rect 31610 18010 31620 18045
rect 31655 18010 31665 18045
rect 31700 18010 31710 18045
rect 31745 18010 31755 18045
rect 31790 18010 31800 18045
rect 31835 18010 31845 18045
rect 31880 18010 31890 18045
rect 31925 18010 31935 18045
rect 31970 18010 31980 18045
rect 32015 18010 32025 18045
rect 32060 18010 32070 18045
rect 32105 18010 32115 18045
rect 32150 18010 32160 18045
rect 32195 18010 32205 18045
rect 32240 18010 32250 18045
rect 32285 18010 32295 18045
rect 32330 18010 32340 18045
rect 32375 18010 32385 18045
rect 32420 18010 32430 18045
rect 32465 18010 32475 18045
rect 32510 18010 32520 18045
rect 32555 18010 32565 18045
rect 32600 18010 32610 18045
rect 32645 18010 32655 18045
rect 32690 18010 32700 18045
rect 32735 18010 32745 18045
rect 32780 18010 32790 18045
rect 32825 18010 32835 18045
rect 32870 18010 32890 18045
rect 2070 18000 32890 18010
rect 2070 17980 31305 18000
rect 2070 17940 2110 17980
rect 2150 17940 6700 17980
rect 6740 17965 31305 17980
rect 31340 17965 31350 18000
rect 31385 17965 31395 18000
rect 31430 17965 31440 18000
rect 31475 17965 31485 18000
rect 31520 17965 31530 18000
rect 31565 17965 31575 18000
rect 31610 17965 31620 18000
rect 31655 17965 31665 18000
rect 31700 17965 31710 18000
rect 31745 17965 31755 18000
rect 31790 17965 31800 18000
rect 31835 17965 31845 18000
rect 31880 17965 31890 18000
rect 31925 17965 31935 18000
rect 31970 17965 31980 18000
rect 32015 17965 32025 18000
rect 32060 17965 32070 18000
rect 32105 17965 32115 18000
rect 32150 17965 32160 18000
rect 32195 17965 32205 18000
rect 32240 17965 32250 18000
rect 32285 17965 32295 18000
rect 32330 17965 32340 18000
rect 32375 17965 32385 18000
rect 32420 17965 32430 18000
rect 32465 17965 32475 18000
rect 32510 17965 32520 18000
rect 32555 17965 32565 18000
rect 32600 17965 32610 18000
rect 32645 17965 32655 18000
rect 32690 17965 32700 18000
rect 32735 17965 32745 18000
rect 32780 17965 32790 18000
rect 32825 17965 32835 18000
rect 32870 17965 32890 18000
rect 6740 17955 32890 17965
rect 6740 17940 31305 17955
rect 2070 17920 31305 17940
rect 31340 17920 31350 17955
rect 31385 17920 31395 17955
rect 31430 17920 31440 17955
rect 31475 17920 31485 17955
rect 31520 17920 31530 17955
rect 31565 17920 31575 17955
rect 31610 17920 31620 17955
rect 31655 17920 31665 17955
rect 31700 17920 31710 17955
rect 31745 17920 31755 17955
rect 31790 17920 31800 17955
rect 31835 17920 31845 17955
rect 31880 17920 31890 17955
rect 31925 17920 31935 17955
rect 31970 17920 31980 17955
rect 32015 17920 32025 17955
rect 32060 17920 32070 17955
rect 32105 17920 32115 17955
rect 32150 17920 32160 17955
rect 32195 17920 32205 17955
rect 32240 17920 32250 17955
rect 32285 17920 32295 17955
rect 32330 17920 32340 17955
rect 32375 17920 32385 17955
rect 32420 17920 32430 17955
rect 32465 17920 32475 17955
rect 32510 17920 32520 17955
rect 32555 17920 32565 17955
rect 32600 17920 32610 17955
rect 32645 17920 32655 17955
rect 32690 17920 32700 17955
rect 32735 17920 32745 17955
rect 32780 17920 32790 17955
rect 32825 17920 32835 17955
rect 32870 17920 32890 17955
rect 2070 17910 32890 17920
rect 2070 17870 2110 17910
rect 2150 17870 6700 17910
rect 6740 17875 31305 17910
rect 31340 17875 31350 17910
rect 31385 17875 31395 17910
rect 31430 17875 31440 17910
rect 31475 17875 31485 17910
rect 31520 17875 31530 17910
rect 31565 17875 31575 17910
rect 31610 17875 31620 17910
rect 31655 17875 31665 17910
rect 31700 17875 31710 17910
rect 31745 17875 31755 17910
rect 31790 17875 31800 17910
rect 31835 17875 31845 17910
rect 31880 17875 31890 17910
rect 31925 17875 31935 17910
rect 31970 17875 31980 17910
rect 32015 17875 32025 17910
rect 32060 17875 32070 17910
rect 32105 17875 32115 17910
rect 32150 17875 32160 17910
rect 32195 17875 32205 17910
rect 32240 17875 32250 17910
rect 32285 17875 32295 17910
rect 32330 17875 32340 17910
rect 32375 17875 32385 17910
rect 32420 17875 32430 17910
rect 32465 17875 32475 17910
rect 32510 17875 32520 17910
rect 32555 17875 32565 17910
rect 32600 17875 32610 17910
rect 32645 17875 32655 17910
rect 32690 17875 32700 17910
rect 32735 17875 32745 17910
rect 32780 17875 32790 17910
rect 32825 17875 32835 17910
rect 32870 17875 32890 17910
rect 6740 17870 32890 17875
rect 2070 17865 32890 17870
rect 2070 17840 31305 17865
rect 2070 17800 2110 17840
rect 2150 17800 6700 17840
rect 6740 17830 31305 17840
rect 31340 17830 31350 17865
rect 31385 17830 31395 17865
rect 31430 17830 31440 17865
rect 31475 17830 31485 17865
rect 31520 17830 31530 17865
rect 31565 17830 31575 17865
rect 31610 17830 31620 17865
rect 31655 17830 31665 17865
rect 31700 17830 31710 17865
rect 31745 17830 31755 17865
rect 31790 17830 31800 17865
rect 31835 17830 31845 17865
rect 31880 17830 31890 17865
rect 31925 17830 31935 17865
rect 31970 17830 31980 17865
rect 32015 17830 32025 17865
rect 32060 17830 32070 17865
rect 32105 17830 32115 17865
rect 32150 17830 32160 17865
rect 32195 17830 32205 17865
rect 32240 17830 32250 17865
rect 32285 17830 32295 17865
rect 32330 17830 32340 17865
rect 32375 17830 32385 17865
rect 32420 17830 32430 17865
rect 32465 17830 32475 17865
rect 32510 17830 32520 17865
rect 32555 17830 32565 17865
rect 32600 17830 32610 17865
rect 32645 17830 32655 17865
rect 32690 17830 32700 17865
rect 32735 17830 32745 17865
rect 32780 17830 32790 17865
rect 32825 17830 32835 17865
rect 32870 17830 32890 17865
rect 6740 17820 32890 17830
rect 6740 17800 31305 17820
rect 2070 17785 31305 17800
rect 31340 17785 31350 17820
rect 31385 17785 31395 17820
rect 31430 17785 31440 17820
rect 31475 17785 31485 17820
rect 31520 17785 31530 17820
rect 31565 17785 31575 17820
rect 31610 17785 31620 17820
rect 31655 17785 31665 17820
rect 31700 17785 31710 17820
rect 31745 17785 31755 17820
rect 31790 17785 31800 17820
rect 31835 17785 31845 17820
rect 31880 17785 31890 17820
rect 31925 17785 31935 17820
rect 31970 17785 31980 17820
rect 32015 17785 32025 17820
rect 32060 17785 32070 17820
rect 32105 17785 32115 17820
rect 32150 17785 32160 17820
rect 32195 17785 32205 17820
rect 32240 17785 32250 17820
rect 32285 17785 32295 17820
rect 32330 17785 32340 17820
rect 32375 17785 32385 17820
rect 32420 17785 32430 17820
rect 32465 17785 32475 17820
rect 32510 17785 32520 17820
rect 32555 17785 32565 17820
rect 32600 17785 32610 17820
rect 32645 17785 32655 17820
rect 32690 17785 32700 17820
rect 32735 17785 32745 17820
rect 32780 17785 32790 17820
rect 32825 17785 32835 17820
rect 32870 17785 32890 17820
rect 2070 17775 32890 17785
rect 2070 17735 2110 17775
rect 2150 17735 6700 17775
rect 6740 17740 31305 17775
rect 31340 17740 31350 17775
rect 31385 17740 31395 17775
rect 31430 17740 31440 17775
rect 31475 17740 31485 17775
rect 31520 17740 31530 17775
rect 31565 17740 31575 17775
rect 31610 17740 31620 17775
rect 31655 17740 31665 17775
rect 31700 17740 31710 17775
rect 31745 17740 31755 17775
rect 31790 17740 31800 17775
rect 31835 17740 31845 17775
rect 31880 17740 31890 17775
rect 31925 17740 31935 17775
rect 31970 17740 31980 17775
rect 32015 17740 32025 17775
rect 32060 17740 32070 17775
rect 32105 17740 32115 17775
rect 32150 17740 32160 17775
rect 32195 17740 32205 17775
rect 32240 17740 32250 17775
rect 32285 17740 32295 17775
rect 32330 17740 32340 17775
rect 32375 17740 32385 17775
rect 32420 17740 32430 17775
rect 32465 17740 32475 17775
rect 32510 17740 32520 17775
rect 32555 17740 32565 17775
rect 32600 17740 32610 17775
rect 32645 17740 32655 17775
rect 32690 17740 32700 17775
rect 32735 17740 32745 17775
rect 32780 17740 32790 17775
rect 32825 17740 32835 17775
rect 32870 17740 32890 17775
rect 6740 17735 32890 17740
rect 2070 17725 32890 17735
rect 31290 10530 35620 10550
rect 31290 10495 31305 10530
rect 31340 10495 31350 10530
rect 31385 10495 31395 10530
rect 31430 10495 31440 10530
rect 31475 10495 31485 10530
rect 31520 10495 31530 10530
rect 31565 10495 31575 10530
rect 31610 10495 31620 10530
rect 31655 10495 31665 10530
rect 31700 10495 31710 10530
rect 31745 10495 31755 10530
rect 31790 10495 31800 10530
rect 31835 10495 31845 10530
rect 31880 10495 31890 10530
rect 31925 10495 31935 10530
rect 31970 10495 31980 10530
rect 32015 10495 32025 10530
rect 32060 10495 32070 10530
rect 32105 10495 32115 10530
rect 32150 10495 32160 10530
rect 32195 10495 32205 10530
rect 32240 10495 32250 10530
rect 32285 10495 32295 10530
rect 32330 10495 32340 10530
rect 32375 10495 32385 10530
rect 32420 10495 32430 10530
rect 32465 10495 32475 10530
rect 32510 10495 32520 10530
rect 32555 10495 32565 10530
rect 32600 10495 32610 10530
rect 32645 10495 32655 10530
rect 32690 10495 32700 10530
rect 32735 10495 32745 10530
rect 32780 10495 32790 10530
rect 32825 10495 32835 10530
rect 32870 10495 35620 10530
rect 31290 10485 35620 10495
rect 31290 10450 31305 10485
rect 31340 10450 31350 10485
rect 31385 10450 31395 10485
rect 31430 10450 31440 10485
rect 31475 10450 31485 10485
rect 31520 10450 31530 10485
rect 31565 10450 31575 10485
rect 31610 10450 31620 10485
rect 31655 10450 31665 10485
rect 31700 10450 31710 10485
rect 31745 10450 31755 10485
rect 31790 10450 31800 10485
rect 31835 10450 31845 10485
rect 31880 10450 31890 10485
rect 31925 10450 31935 10485
rect 31970 10450 31980 10485
rect 32015 10450 32025 10485
rect 32060 10450 32070 10485
rect 32105 10450 32115 10485
rect 32150 10450 32160 10485
rect 32195 10450 32205 10485
rect 32240 10450 32250 10485
rect 32285 10450 32295 10485
rect 32330 10450 32340 10485
rect 32375 10450 32385 10485
rect 32420 10450 32430 10485
rect 32465 10450 32475 10485
rect 32510 10450 32520 10485
rect 32555 10450 32565 10485
rect 32600 10450 32610 10485
rect 32645 10450 32655 10485
rect 32690 10450 32700 10485
rect 32735 10450 32745 10485
rect 32780 10450 32790 10485
rect 32825 10450 32835 10485
rect 32870 10450 35620 10485
rect 31290 10440 35620 10450
rect 31290 10405 31305 10440
rect 31340 10405 31350 10440
rect 31385 10405 31395 10440
rect 31430 10405 31440 10440
rect 31475 10405 31485 10440
rect 31520 10405 31530 10440
rect 31565 10405 31575 10440
rect 31610 10405 31620 10440
rect 31655 10405 31665 10440
rect 31700 10405 31710 10440
rect 31745 10405 31755 10440
rect 31790 10405 31800 10440
rect 31835 10405 31845 10440
rect 31880 10405 31890 10440
rect 31925 10405 31935 10440
rect 31970 10405 31980 10440
rect 32015 10405 32025 10440
rect 32060 10405 32070 10440
rect 32105 10405 32115 10440
rect 32150 10405 32160 10440
rect 32195 10405 32205 10440
rect 32240 10405 32250 10440
rect 32285 10405 32295 10440
rect 32330 10405 32340 10440
rect 32375 10405 32385 10440
rect 32420 10405 32430 10440
rect 32465 10405 32475 10440
rect 32510 10405 32520 10440
rect 32555 10405 32565 10440
rect 32600 10405 32610 10440
rect 32645 10405 32655 10440
rect 32690 10405 32700 10440
rect 32735 10405 32745 10440
rect 32780 10405 32790 10440
rect 32825 10405 32835 10440
rect 32870 10405 35620 10440
rect 31290 10395 35620 10405
rect 31290 10360 31305 10395
rect 31340 10360 31350 10395
rect 31385 10360 31395 10395
rect 31430 10360 31440 10395
rect 31475 10360 31485 10395
rect 31520 10360 31530 10395
rect 31565 10360 31575 10395
rect 31610 10360 31620 10395
rect 31655 10360 31665 10395
rect 31700 10360 31710 10395
rect 31745 10360 31755 10395
rect 31790 10360 31800 10395
rect 31835 10360 31845 10395
rect 31880 10360 31890 10395
rect 31925 10360 31935 10395
rect 31970 10360 31980 10395
rect 32015 10360 32025 10395
rect 32060 10360 32070 10395
rect 32105 10360 32115 10395
rect 32150 10360 32160 10395
rect 32195 10360 32205 10395
rect 32240 10360 32250 10395
rect 32285 10360 32295 10395
rect 32330 10360 32340 10395
rect 32375 10360 32385 10395
rect 32420 10360 32430 10395
rect 32465 10360 32475 10395
rect 32510 10360 32520 10395
rect 32555 10360 32565 10395
rect 32600 10360 32610 10395
rect 32645 10360 32655 10395
rect 32690 10360 32700 10395
rect 32735 10360 32745 10395
rect 32780 10360 32790 10395
rect 32825 10360 32835 10395
rect 32870 10360 35620 10395
rect 31290 10350 35620 10360
rect 31290 10315 31305 10350
rect 31340 10315 31350 10350
rect 31385 10315 31395 10350
rect 31430 10315 31440 10350
rect 31475 10315 31485 10350
rect 31520 10315 31530 10350
rect 31565 10315 31575 10350
rect 31610 10315 31620 10350
rect 31655 10315 31665 10350
rect 31700 10315 31710 10350
rect 31745 10315 31755 10350
rect 31790 10315 31800 10350
rect 31835 10315 31845 10350
rect 31880 10315 31890 10350
rect 31925 10315 31935 10350
rect 31970 10315 31980 10350
rect 32015 10315 32025 10350
rect 32060 10315 32070 10350
rect 32105 10315 32115 10350
rect 32150 10315 32160 10350
rect 32195 10315 32205 10350
rect 32240 10315 32250 10350
rect 32285 10315 32295 10350
rect 32330 10315 32340 10350
rect 32375 10315 32385 10350
rect 32420 10315 32430 10350
rect 32465 10315 32475 10350
rect 32510 10315 32520 10350
rect 32555 10315 32565 10350
rect 32600 10315 32610 10350
rect 32645 10315 32655 10350
rect 32690 10315 32700 10350
rect 32735 10315 32745 10350
rect 32780 10315 32790 10350
rect 32825 10315 32835 10350
rect 32870 10315 35620 10350
rect 31290 10305 35620 10315
rect 31290 10270 31305 10305
rect 31340 10270 31350 10305
rect 31385 10270 31395 10305
rect 31430 10270 31440 10305
rect 31475 10270 31485 10305
rect 31520 10270 31530 10305
rect 31565 10270 31575 10305
rect 31610 10270 31620 10305
rect 31655 10270 31665 10305
rect 31700 10270 31710 10305
rect 31745 10270 31755 10305
rect 31790 10270 31800 10305
rect 31835 10270 31845 10305
rect 31880 10270 31890 10305
rect 31925 10270 31935 10305
rect 31970 10270 31980 10305
rect 32015 10270 32025 10305
rect 32060 10270 32070 10305
rect 32105 10270 32115 10305
rect 32150 10270 32160 10305
rect 32195 10270 32205 10305
rect 32240 10270 32250 10305
rect 32285 10270 32295 10305
rect 32330 10270 32340 10305
rect 32375 10270 32385 10305
rect 32420 10270 32430 10305
rect 32465 10270 32475 10305
rect 32510 10270 32520 10305
rect 32555 10270 32565 10305
rect 32600 10270 32610 10305
rect 32645 10270 32655 10305
rect 32690 10270 32700 10305
rect 32735 10270 32745 10305
rect 32780 10270 32790 10305
rect 32825 10270 32835 10305
rect 32870 10270 35620 10305
rect 31290 10260 35620 10270
rect 31290 10225 31305 10260
rect 31340 10225 31350 10260
rect 31385 10225 31395 10260
rect 31430 10225 31440 10260
rect 31475 10225 31485 10260
rect 31520 10225 31530 10260
rect 31565 10225 31575 10260
rect 31610 10225 31620 10260
rect 31655 10225 31665 10260
rect 31700 10225 31710 10260
rect 31745 10225 31755 10260
rect 31790 10225 31800 10260
rect 31835 10225 31845 10260
rect 31880 10225 31890 10260
rect 31925 10225 31935 10260
rect 31970 10225 31980 10260
rect 32015 10225 32025 10260
rect 32060 10225 32070 10260
rect 32105 10225 32115 10260
rect 32150 10225 32160 10260
rect 32195 10225 32205 10260
rect 32240 10225 32250 10260
rect 32285 10225 32295 10260
rect 32330 10225 32340 10260
rect 32375 10225 32385 10260
rect 32420 10225 32430 10260
rect 32465 10225 32475 10260
rect 32510 10225 32520 10260
rect 32555 10225 32565 10260
rect 32600 10225 32610 10260
rect 32645 10225 32655 10260
rect 32690 10225 32700 10260
rect 32735 10225 32745 10260
rect 32780 10225 32790 10260
rect 32825 10225 32835 10260
rect 32870 10225 35620 10260
rect 31290 10215 35620 10225
rect 31290 10180 31305 10215
rect 31340 10180 31350 10215
rect 31385 10180 31395 10215
rect 31430 10180 31440 10215
rect 31475 10180 31485 10215
rect 31520 10180 31530 10215
rect 31565 10180 31575 10215
rect 31610 10180 31620 10215
rect 31655 10180 31665 10215
rect 31700 10180 31710 10215
rect 31745 10180 31755 10215
rect 31790 10180 31800 10215
rect 31835 10180 31845 10215
rect 31880 10180 31890 10215
rect 31925 10180 31935 10215
rect 31970 10180 31980 10215
rect 32015 10180 32025 10215
rect 32060 10180 32070 10215
rect 32105 10180 32115 10215
rect 32150 10180 32160 10215
rect 32195 10180 32205 10215
rect 32240 10180 32250 10215
rect 32285 10180 32295 10215
rect 32330 10180 32340 10215
rect 32375 10180 32385 10215
rect 32420 10180 32430 10215
rect 32465 10180 32475 10215
rect 32510 10180 32520 10215
rect 32555 10180 32565 10215
rect 32600 10180 32610 10215
rect 32645 10180 32655 10215
rect 32690 10180 32700 10215
rect 32735 10180 32745 10215
rect 32780 10180 32790 10215
rect 32825 10180 32835 10215
rect 32870 10180 35620 10215
rect 31290 10170 35620 10180
rect 31290 10135 31305 10170
rect 31340 10135 31350 10170
rect 31385 10135 31395 10170
rect 31430 10135 31440 10170
rect 31475 10135 31485 10170
rect 31520 10135 31530 10170
rect 31565 10135 31575 10170
rect 31610 10135 31620 10170
rect 31655 10135 31665 10170
rect 31700 10135 31710 10170
rect 31745 10135 31755 10170
rect 31790 10135 31800 10170
rect 31835 10135 31845 10170
rect 31880 10135 31890 10170
rect 31925 10135 31935 10170
rect 31970 10135 31980 10170
rect 32015 10135 32025 10170
rect 32060 10135 32070 10170
rect 32105 10135 32115 10170
rect 32150 10135 32160 10170
rect 32195 10135 32205 10170
rect 32240 10135 32250 10170
rect 32285 10135 32295 10170
rect 32330 10135 32340 10170
rect 32375 10135 32385 10170
rect 32420 10135 32430 10170
rect 32465 10135 32475 10170
rect 32510 10135 32520 10170
rect 32555 10135 32565 10170
rect 32600 10135 32610 10170
rect 32645 10135 32655 10170
rect 32690 10135 32700 10170
rect 32735 10135 32745 10170
rect 32780 10135 32790 10170
rect 32825 10135 32835 10170
rect 32870 10135 35620 10170
rect 31290 10125 35620 10135
rect 31290 10090 31305 10125
rect 31340 10090 31350 10125
rect 31385 10090 31395 10125
rect 31430 10090 31440 10125
rect 31475 10090 31485 10125
rect 31520 10090 31530 10125
rect 31565 10090 31575 10125
rect 31610 10090 31620 10125
rect 31655 10090 31665 10125
rect 31700 10090 31710 10125
rect 31745 10090 31755 10125
rect 31790 10090 31800 10125
rect 31835 10090 31845 10125
rect 31880 10090 31890 10125
rect 31925 10090 31935 10125
rect 31970 10090 31980 10125
rect 32015 10090 32025 10125
rect 32060 10090 32070 10125
rect 32105 10090 32115 10125
rect 32150 10090 32160 10125
rect 32195 10090 32205 10125
rect 32240 10090 32250 10125
rect 32285 10090 32295 10125
rect 32330 10090 32340 10125
rect 32375 10090 32385 10125
rect 32420 10090 32430 10125
rect 32465 10090 32475 10125
rect 32510 10090 32520 10125
rect 32555 10090 32565 10125
rect 32600 10090 32610 10125
rect 32645 10090 32655 10125
rect 32690 10090 32700 10125
rect 32735 10090 32745 10125
rect 32780 10090 32790 10125
rect 32825 10090 32835 10125
rect 32870 10090 35620 10125
rect 31290 10080 35620 10090
rect 31290 10045 31305 10080
rect 31340 10045 31350 10080
rect 31385 10045 31395 10080
rect 31430 10045 31440 10080
rect 31475 10045 31485 10080
rect 31520 10045 31530 10080
rect 31565 10045 31575 10080
rect 31610 10045 31620 10080
rect 31655 10045 31665 10080
rect 31700 10045 31710 10080
rect 31745 10045 31755 10080
rect 31790 10045 31800 10080
rect 31835 10045 31845 10080
rect 31880 10045 31890 10080
rect 31925 10045 31935 10080
rect 31970 10045 31980 10080
rect 32015 10045 32025 10080
rect 32060 10045 32070 10080
rect 32105 10045 32115 10080
rect 32150 10045 32160 10080
rect 32195 10045 32205 10080
rect 32240 10045 32250 10080
rect 32285 10045 32295 10080
rect 32330 10045 32340 10080
rect 32375 10045 32385 10080
rect 32420 10045 32430 10080
rect 32465 10045 32475 10080
rect 32510 10045 32520 10080
rect 32555 10045 32565 10080
rect 32600 10045 32610 10080
rect 32645 10045 32655 10080
rect 32690 10045 32700 10080
rect 32735 10045 32745 10080
rect 32780 10045 32790 10080
rect 32825 10045 32835 10080
rect 32870 10045 35620 10080
rect 31290 10035 35620 10045
rect 31290 10000 31305 10035
rect 31340 10000 31350 10035
rect 31385 10000 31395 10035
rect 31430 10000 31440 10035
rect 31475 10000 31485 10035
rect 31520 10000 31530 10035
rect 31565 10000 31575 10035
rect 31610 10000 31620 10035
rect 31655 10000 31665 10035
rect 31700 10000 31710 10035
rect 31745 10000 31755 10035
rect 31790 10000 31800 10035
rect 31835 10000 31845 10035
rect 31880 10000 31890 10035
rect 31925 10000 31935 10035
rect 31970 10000 31980 10035
rect 32015 10000 32025 10035
rect 32060 10000 32070 10035
rect 32105 10000 32115 10035
rect 32150 10000 32160 10035
rect 32195 10000 32205 10035
rect 32240 10000 32250 10035
rect 32285 10000 32295 10035
rect 32330 10000 32340 10035
rect 32375 10000 32385 10035
rect 32420 10000 32430 10035
rect 32465 10000 32475 10035
rect 32510 10000 32520 10035
rect 32555 10000 32565 10035
rect 32600 10000 32610 10035
rect 32645 10000 32655 10035
rect 32690 10000 32700 10035
rect 32735 10000 32745 10035
rect 32780 10000 32790 10035
rect 32825 10000 32835 10035
rect 32870 10000 35620 10035
rect 31290 9990 35620 10000
rect 31290 9955 31305 9990
rect 31340 9955 31350 9990
rect 31385 9955 31395 9990
rect 31430 9955 31440 9990
rect 31475 9955 31485 9990
rect 31520 9955 31530 9990
rect 31565 9955 31575 9990
rect 31610 9955 31620 9990
rect 31655 9955 31665 9990
rect 31700 9955 31710 9990
rect 31745 9955 31755 9990
rect 31790 9955 31800 9990
rect 31835 9955 31845 9990
rect 31880 9955 31890 9990
rect 31925 9955 31935 9990
rect 31970 9955 31980 9990
rect 32015 9955 32025 9990
rect 32060 9955 32070 9990
rect 32105 9955 32115 9990
rect 32150 9955 32160 9990
rect 32195 9955 32205 9990
rect 32240 9955 32250 9990
rect 32285 9955 32295 9990
rect 32330 9955 32340 9990
rect 32375 9955 32385 9990
rect 32420 9955 32430 9990
rect 32465 9955 32475 9990
rect 32510 9955 32520 9990
rect 32555 9955 32565 9990
rect 32600 9955 32610 9990
rect 32645 9955 32655 9990
rect 32690 9955 32700 9990
rect 32735 9955 32745 9990
rect 32780 9955 32790 9990
rect 32825 9955 32835 9990
rect 32870 9955 35620 9990
rect 31290 9945 35620 9955
rect 31290 9910 31305 9945
rect 31340 9910 31350 9945
rect 31385 9910 31395 9945
rect 31430 9910 31440 9945
rect 31475 9910 31485 9945
rect 31520 9910 31530 9945
rect 31565 9910 31575 9945
rect 31610 9910 31620 9945
rect 31655 9910 31665 9945
rect 31700 9910 31710 9945
rect 31745 9910 31755 9945
rect 31790 9910 31800 9945
rect 31835 9910 31845 9945
rect 31880 9910 31890 9945
rect 31925 9910 31935 9945
rect 31970 9910 31980 9945
rect 32015 9910 32025 9945
rect 32060 9910 32070 9945
rect 32105 9910 32115 9945
rect 32150 9910 32160 9945
rect 32195 9910 32205 9945
rect 32240 9910 32250 9945
rect 32285 9910 32295 9945
rect 32330 9910 32340 9945
rect 32375 9910 32385 9945
rect 32420 9910 32430 9945
rect 32465 9910 32475 9945
rect 32510 9910 32520 9945
rect 32555 9910 32565 9945
rect 32600 9910 32610 9945
rect 32645 9910 32655 9945
rect 32690 9910 32700 9945
rect 32735 9910 32745 9945
rect 32780 9910 32790 9945
rect 32825 9910 32835 9945
rect 32870 9910 35620 9945
rect 31290 9900 35620 9910
rect 31290 9865 31305 9900
rect 31340 9865 31350 9900
rect 31385 9865 31395 9900
rect 31430 9865 31440 9900
rect 31475 9865 31485 9900
rect 31520 9865 31530 9900
rect 31565 9865 31575 9900
rect 31610 9865 31620 9900
rect 31655 9865 31665 9900
rect 31700 9865 31710 9900
rect 31745 9865 31755 9900
rect 31790 9865 31800 9900
rect 31835 9865 31845 9900
rect 31880 9865 31890 9900
rect 31925 9865 31935 9900
rect 31970 9865 31980 9900
rect 32015 9865 32025 9900
rect 32060 9865 32070 9900
rect 32105 9865 32115 9900
rect 32150 9865 32160 9900
rect 32195 9865 32205 9900
rect 32240 9865 32250 9900
rect 32285 9865 32295 9900
rect 32330 9865 32340 9900
rect 32375 9865 32385 9900
rect 32420 9865 32430 9900
rect 32465 9865 32475 9900
rect 32510 9865 32520 9900
rect 32555 9865 32565 9900
rect 32600 9865 32610 9900
rect 32645 9865 32655 9900
rect 32690 9865 32700 9900
rect 32735 9865 32745 9900
rect 32780 9865 32790 9900
rect 32825 9865 32835 9900
rect 32870 9865 35620 9900
rect 31290 9855 35620 9865
rect 31290 9820 31305 9855
rect 31340 9820 31350 9855
rect 31385 9820 31395 9855
rect 31430 9820 31440 9855
rect 31475 9820 31485 9855
rect 31520 9820 31530 9855
rect 31565 9820 31575 9855
rect 31610 9820 31620 9855
rect 31655 9820 31665 9855
rect 31700 9820 31710 9855
rect 31745 9820 31755 9855
rect 31790 9820 31800 9855
rect 31835 9820 31845 9855
rect 31880 9820 31890 9855
rect 31925 9820 31935 9855
rect 31970 9820 31980 9855
rect 32015 9820 32025 9855
rect 32060 9820 32070 9855
rect 32105 9820 32115 9855
rect 32150 9820 32160 9855
rect 32195 9820 32205 9855
rect 32240 9820 32250 9855
rect 32285 9820 32295 9855
rect 32330 9820 32340 9855
rect 32375 9820 32385 9855
rect 32420 9820 32430 9855
rect 32465 9820 32475 9855
rect 32510 9820 32520 9855
rect 32555 9820 32565 9855
rect 32600 9820 32610 9855
rect 32645 9820 32655 9855
rect 32690 9820 32700 9855
rect 32735 9820 32745 9855
rect 32780 9820 32790 9855
rect 32825 9820 32835 9855
rect 32870 9820 35620 9855
rect 31290 9810 35620 9820
rect 31290 9775 31305 9810
rect 31340 9775 31350 9810
rect 31385 9775 31395 9810
rect 31430 9775 31440 9810
rect 31475 9775 31485 9810
rect 31520 9775 31530 9810
rect 31565 9775 31575 9810
rect 31610 9775 31620 9810
rect 31655 9775 31665 9810
rect 31700 9775 31710 9810
rect 31745 9775 31755 9810
rect 31790 9775 31800 9810
rect 31835 9775 31845 9810
rect 31880 9775 31890 9810
rect 31925 9775 31935 9810
rect 31970 9775 31980 9810
rect 32015 9775 32025 9810
rect 32060 9775 32070 9810
rect 32105 9775 32115 9810
rect 32150 9775 32160 9810
rect 32195 9775 32205 9810
rect 32240 9775 32250 9810
rect 32285 9775 32295 9810
rect 32330 9775 32340 9810
rect 32375 9775 32385 9810
rect 32420 9775 32430 9810
rect 32465 9775 32475 9810
rect 32510 9775 32520 9810
rect 32555 9775 32565 9810
rect 32600 9775 32610 9810
rect 32645 9775 32655 9810
rect 32690 9775 32700 9810
rect 32735 9775 32745 9810
rect 32780 9775 32790 9810
rect 32825 9775 32835 9810
rect 32870 9775 35620 9810
rect 31290 9765 35620 9775
rect 31290 9730 31305 9765
rect 31340 9730 31350 9765
rect 31385 9730 31395 9765
rect 31430 9730 31440 9765
rect 31475 9730 31485 9765
rect 31520 9730 31530 9765
rect 31565 9730 31575 9765
rect 31610 9730 31620 9765
rect 31655 9730 31665 9765
rect 31700 9730 31710 9765
rect 31745 9730 31755 9765
rect 31790 9730 31800 9765
rect 31835 9730 31845 9765
rect 31880 9730 31890 9765
rect 31925 9730 31935 9765
rect 31970 9730 31980 9765
rect 32015 9730 32025 9765
rect 32060 9730 32070 9765
rect 32105 9730 32115 9765
rect 32150 9730 32160 9765
rect 32195 9730 32205 9765
rect 32240 9730 32250 9765
rect 32285 9730 32295 9765
rect 32330 9730 32340 9765
rect 32375 9730 32385 9765
rect 32420 9730 32430 9765
rect 32465 9730 32475 9765
rect 32510 9730 32520 9765
rect 32555 9730 32565 9765
rect 32600 9730 32610 9765
rect 32645 9730 32655 9765
rect 32690 9730 32700 9765
rect 32735 9730 32745 9765
rect 32780 9730 32790 9765
rect 32825 9730 32835 9765
rect 32870 9730 35620 9765
rect 31290 9720 35620 9730
rect 31290 9685 31305 9720
rect 31340 9685 31350 9720
rect 31385 9685 31395 9720
rect 31430 9685 31440 9720
rect 31475 9685 31485 9720
rect 31520 9685 31530 9720
rect 31565 9685 31575 9720
rect 31610 9685 31620 9720
rect 31655 9685 31665 9720
rect 31700 9685 31710 9720
rect 31745 9685 31755 9720
rect 31790 9685 31800 9720
rect 31835 9685 31845 9720
rect 31880 9685 31890 9720
rect 31925 9685 31935 9720
rect 31970 9685 31980 9720
rect 32015 9685 32025 9720
rect 32060 9685 32070 9720
rect 32105 9685 32115 9720
rect 32150 9685 32160 9720
rect 32195 9685 32205 9720
rect 32240 9685 32250 9720
rect 32285 9685 32295 9720
rect 32330 9685 32340 9720
rect 32375 9685 32385 9720
rect 32420 9685 32430 9720
rect 32465 9685 32475 9720
rect 32510 9685 32520 9720
rect 32555 9685 32565 9720
rect 32600 9685 32610 9720
rect 32645 9685 32655 9720
rect 32690 9685 32700 9720
rect 32735 9685 32745 9720
rect 32780 9685 32790 9720
rect 32825 9685 32835 9720
rect 32870 9685 35620 9720
rect 31290 9675 35620 9685
rect -38770 9640 7700 9650
rect -38770 9630 1320 9640
rect -38770 9595 -38755 9630
rect -38720 9595 -38710 9630
rect -38675 9595 -38665 9630
rect -38630 9595 -38620 9630
rect -38585 9595 -38575 9630
rect -38540 9595 -38530 9630
rect -38495 9595 -38485 9630
rect -38450 9595 -38440 9630
rect -38405 9595 -38395 9630
rect -38360 9595 -38350 9630
rect -38315 9595 -38305 9630
rect -38270 9595 -38260 9630
rect -38225 9595 -38215 9630
rect -38180 9595 -38170 9630
rect -38135 9595 -38125 9630
rect -38090 9595 -38080 9630
rect -38045 9595 -38035 9630
rect -38000 9595 -37990 9630
rect -37955 9595 -37945 9630
rect -37910 9595 -37900 9630
rect -37865 9595 -37855 9630
rect -37820 9595 -37810 9630
rect -37775 9595 -37765 9630
rect -37730 9595 -37720 9630
rect -37685 9595 -37675 9630
rect -37640 9595 -37630 9630
rect -37595 9595 -37585 9630
rect -37550 9595 -37540 9630
rect -37505 9595 -37495 9630
rect -37460 9595 -37450 9630
rect -37415 9595 -37405 9630
rect -37370 9595 -37360 9630
rect -37325 9595 -37315 9630
rect -37280 9595 -37270 9630
rect -37235 9595 -37225 9630
rect -37190 9600 1320 9630
rect 1360 9600 2245 9640
rect 2285 9600 3175 9640
rect 3215 9600 6700 9640
rect 6740 9600 7620 9640
rect 7660 9600 7700 9640
rect -37190 9595 7700 9600
rect -38770 9585 7700 9595
rect -38770 9550 -38755 9585
rect -38720 9550 -38710 9585
rect -38675 9550 -38665 9585
rect -38630 9550 -38620 9585
rect -38585 9550 -38575 9585
rect -38540 9550 -38530 9585
rect -38495 9550 -38485 9585
rect -38450 9550 -38440 9585
rect -38405 9550 -38395 9585
rect -38360 9550 -38350 9585
rect -38315 9550 -38305 9585
rect -38270 9550 -38260 9585
rect -38225 9550 -38215 9585
rect -38180 9550 -38170 9585
rect -38135 9550 -38125 9585
rect -38090 9550 -38080 9585
rect -38045 9550 -38035 9585
rect -38000 9550 -37990 9585
rect -37955 9550 -37945 9585
rect -37910 9550 -37900 9585
rect -37865 9550 -37855 9585
rect -37820 9550 -37810 9585
rect -37775 9550 -37765 9585
rect -37730 9550 -37720 9585
rect -37685 9550 -37675 9585
rect -37640 9550 -37630 9585
rect -37595 9550 -37585 9585
rect -37550 9550 -37540 9585
rect -37505 9550 -37495 9585
rect -37460 9550 -37450 9585
rect -37415 9550 -37405 9585
rect -37370 9550 -37360 9585
rect -37325 9550 -37315 9585
rect -37280 9550 -37270 9585
rect -37235 9550 -37225 9585
rect -37190 9575 7700 9585
rect -37190 9550 1320 9575
rect -38770 9540 1320 9550
rect -38770 9505 -38755 9540
rect -38720 9505 -38710 9540
rect -38675 9505 -38665 9540
rect -38630 9505 -38620 9540
rect -38585 9505 -38575 9540
rect -38540 9505 -38530 9540
rect -38495 9505 -38485 9540
rect -38450 9505 -38440 9540
rect -38405 9505 -38395 9540
rect -38360 9505 -38350 9540
rect -38315 9505 -38305 9540
rect -38270 9505 -38260 9540
rect -38225 9505 -38215 9540
rect -38180 9505 -38170 9540
rect -38135 9505 -38125 9540
rect -38090 9505 -38080 9540
rect -38045 9505 -38035 9540
rect -38000 9505 -37990 9540
rect -37955 9505 -37945 9540
rect -37910 9505 -37900 9540
rect -37865 9505 -37855 9540
rect -37820 9505 -37810 9540
rect -37775 9505 -37765 9540
rect -37730 9505 -37720 9540
rect -37685 9505 -37675 9540
rect -37640 9505 -37630 9540
rect -37595 9505 -37585 9540
rect -37550 9505 -37540 9540
rect -37505 9505 -37495 9540
rect -37460 9505 -37450 9540
rect -37415 9505 -37405 9540
rect -37370 9505 -37360 9540
rect -37325 9505 -37315 9540
rect -37280 9505 -37270 9540
rect -37235 9505 -37225 9540
rect -37190 9535 1320 9540
rect 1360 9535 2245 9575
rect 2285 9535 3175 9575
rect 3215 9535 6700 9575
rect 6740 9535 7620 9575
rect 7660 9535 7700 9575
rect -37190 9505 7700 9535
rect -38770 9495 1320 9505
rect -38770 9460 -38755 9495
rect -38720 9460 -38710 9495
rect -38675 9460 -38665 9495
rect -38630 9460 -38620 9495
rect -38585 9460 -38575 9495
rect -38540 9460 -38530 9495
rect -38495 9460 -38485 9495
rect -38450 9460 -38440 9495
rect -38405 9460 -38395 9495
rect -38360 9460 -38350 9495
rect -38315 9460 -38305 9495
rect -38270 9460 -38260 9495
rect -38225 9460 -38215 9495
rect -38180 9460 -38170 9495
rect -38135 9460 -38125 9495
rect -38090 9460 -38080 9495
rect -38045 9460 -38035 9495
rect -38000 9460 -37990 9495
rect -37955 9460 -37945 9495
rect -37910 9460 -37900 9495
rect -37865 9460 -37855 9495
rect -37820 9460 -37810 9495
rect -37775 9460 -37765 9495
rect -37730 9460 -37720 9495
rect -37685 9460 -37675 9495
rect -37640 9460 -37630 9495
rect -37595 9460 -37585 9495
rect -37550 9460 -37540 9495
rect -37505 9460 -37495 9495
rect -37460 9460 -37450 9495
rect -37415 9460 -37405 9495
rect -37370 9460 -37360 9495
rect -37325 9460 -37315 9495
rect -37280 9460 -37270 9495
rect -37235 9460 -37225 9495
rect -37190 9465 1320 9495
rect 1360 9465 2245 9505
rect 2285 9465 3175 9505
rect 3215 9465 6700 9505
rect 6740 9465 7620 9505
rect 7660 9465 7700 9505
rect -37190 9460 7700 9465
rect -38770 9450 7700 9460
rect -38770 9415 -38755 9450
rect -38720 9415 -38710 9450
rect -38675 9415 -38665 9450
rect -38630 9415 -38620 9450
rect -38585 9415 -38575 9450
rect -38540 9415 -38530 9450
rect -38495 9415 -38485 9450
rect -38450 9415 -38440 9450
rect -38405 9415 -38395 9450
rect -38360 9415 -38350 9450
rect -38315 9415 -38305 9450
rect -38270 9415 -38260 9450
rect -38225 9415 -38215 9450
rect -38180 9415 -38170 9450
rect -38135 9415 -38125 9450
rect -38090 9415 -38080 9450
rect -38045 9415 -38035 9450
rect -38000 9415 -37990 9450
rect -37955 9415 -37945 9450
rect -37910 9415 -37900 9450
rect -37865 9415 -37855 9450
rect -37820 9415 -37810 9450
rect -37775 9415 -37765 9450
rect -37730 9415 -37720 9450
rect -37685 9415 -37675 9450
rect -37640 9415 -37630 9450
rect -37595 9415 -37585 9450
rect -37550 9415 -37540 9450
rect -37505 9415 -37495 9450
rect -37460 9415 -37450 9450
rect -37415 9415 -37405 9450
rect -37370 9415 -37360 9450
rect -37325 9415 -37315 9450
rect -37280 9415 -37270 9450
rect -37235 9415 -37225 9450
rect -37190 9435 7700 9450
rect -37190 9415 1320 9435
rect -38770 9405 1320 9415
rect -38770 9370 -38755 9405
rect -38720 9370 -38710 9405
rect -38675 9370 -38665 9405
rect -38630 9370 -38620 9405
rect -38585 9370 -38575 9405
rect -38540 9370 -38530 9405
rect -38495 9370 -38485 9405
rect -38450 9370 -38440 9405
rect -38405 9370 -38395 9405
rect -38360 9370 -38350 9405
rect -38315 9370 -38305 9405
rect -38270 9370 -38260 9405
rect -38225 9370 -38215 9405
rect -38180 9370 -38170 9405
rect -38135 9370 -38125 9405
rect -38090 9370 -38080 9405
rect -38045 9370 -38035 9405
rect -38000 9370 -37990 9405
rect -37955 9370 -37945 9405
rect -37910 9370 -37900 9405
rect -37865 9370 -37855 9405
rect -37820 9370 -37810 9405
rect -37775 9370 -37765 9405
rect -37730 9370 -37720 9405
rect -37685 9370 -37675 9405
rect -37640 9370 -37630 9405
rect -37595 9370 -37585 9405
rect -37550 9370 -37540 9405
rect -37505 9370 -37495 9405
rect -37460 9370 -37450 9405
rect -37415 9370 -37405 9405
rect -37370 9370 -37360 9405
rect -37325 9370 -37315 9405
rect -37280 9370 -37270 9405
rect -37235 9370 -37225 9405
rect -37190 9395 1320 9405
rect 1360 9395 2245 9435
rect 2285 9395 3175 9435
rect 3215 9395 6700 9435
rect 6740 9395 7620 9435
rect 7660 9395 7700 9435
rect -37190 9370 7700 9395
rect -38770 9365 7700 9370
rect -38770 9360 1320 9365
rect -38770 9325 -38755 9360
rect -38720 9325 -38710 9360
rect -38675 9325 -38665 9360
rect -38630 9325 -38620 9360
rect -38585 9325 -38575 9360
rect -38540 9325 -38530 9360
rect -38495 9325 -38485 9360
rect -38450 9325 -38440 9360
rect -38405 9325 -38395 9360
rect -38360 9325 -38350 9360
rect -38315 9325 -38305 9360
rect -38270 9325 -38260 9360
rect -38225 9325 -38215 9360
rect -38180 9325 -38170 9360
rect -38135 9325 -38125 9360
rect -38090 9325 -38080 9360
rect -38045 9325 -38035 9360
rect -38000 9325 -37990 9360
rect -37955 9325 -37945 9360
rect -37910 9325 -37900 9360
rect -37865 9325 -37855 9360
rect -37820 9325 -37810 9360
rect -37775 9325 -37765 9360
rect -37730 9325 -37720 9360
rect -37685 9325 -37675 9360
rect -37640 9325 -37630 9360
rect -37595 9325 -37585 9360
rect -37550 9325 -37540 9360
rect -37505 9325 -37495 9360
rect -37460 9325 -37450 9360
rect -37415 9325 -37405 9360
rect -37370 9325 -37360 9360
rect -37325 9325 -37315 9360
rect -37280 9325 -37270 9360
rect -37235 9325 -37225 9360
rect -37190 9325 1320 9360
rect 1360 9325 2245 9365
rect 2285 9325 3175 9365
rect 3215 9325 6700 9365
rect 6740 9325 7620 9365
rect 7660 9325 7700 9365
rect -38770 9315 7700 9325
rect -38770 9280 -38755 9315
rect -38720 9280 -38710 9315
rect -38675 9280 -38665 9315
rect -38630 9280 -38620 9315
rect -38585 9280 -38575 9315
rect -38540 9280 -38530 9315
rect -38495 9280 -38485 9315
rect -38450 9280 -38440 9315
rect -38405 9280 -38395 9315
rect -38360 9280 -38350 9315
rect -38315 9280 -38305 9315
rect -38270 9280 -38260 9315
rect -38225 9280 -38215 9315
rect -38180 9280 -38170 9315
rect -38135 9280 -38125 9315
rect -38090 9280 -38080 9315
rect -38045 9280 -38035 9315
rect -38000 9280 -37990 9315
rect -37955 9280 -37945 9315
rect -37910 9280 -37900 9315
rect -37865 9280 -37855 9315
rect -37820 9280 -37810 9315
rect -37775 9280 -37765 9315
rect -37730 9280 -37720 9315
rect -37685 9280 -37675 9315
rect -37640 9280 -37630 9315
rect -37595 9280 -37585 9315
rect -37550 9280 -37540 9315
rect -37505 9280 -37495 9315
rect -37460 9280 -37450 9315
rect -37415 9280 -37405 9315
rect -37370 9280 -37360 9315
rect -37325 9280 -37315 9315
rect -37280 9280 -37270 9315
rect -37235 9280 -37225 9315
rect -37190 9300 7700 9315
rect -37190 9280 1320 9300
rect -38770 9270 1320 9280
rect -38770 9235 -38755 9270
rect -38720 9235 -38710 9270
rect -38675 9235 -38665 9270
rect -38630 9235 -38620 9270
rect -38585 9235 -38575 9270
rect -38540 9235 -38530 9270
rect -38495 9235 -38485 9270
rect -38450 9235 -38440 9270
rect -38405 9235 -38395 9270
rect -38360 9235 -38350 9270
rect -38315 9235 -38305 9270
rect -38270 9235 -38260 9270
rect -38225 9235 -38215 9270
rect -38180 9235 -38170 9270
rect -38135 9235 -38125 9270
rect -38090 9235 -38080 9270
rect -38045 9235 -38035 9270
rect -38000 9235 -37990 9270
rect -37955 9235 -37945 9270
rect -37910 9235 -37900 9270
rect -37865 9235 -37855 9270
rect -37820 9235 -37810 9270
rect -37775 9235 -37765 9270
rect -37730 9235 -37720 9270
rect -37685 9235 -37675 9270
rect -37640 9235 -37630 9270
rect -37595 9235 -37585 9270
rect -37550 9235 -37540 9270
rect -37505 9235 -37495 9270
rect -37460 9235 -37450 9270
rect -37415 9235 -37405 9270
rect -37370 9235 -37360 9270
rect -37325 9235 -37315 9270
rect -37280 9235 -37270 9270
rect -37235 9235 -37225 9270
rect -37190 9260 1320 9270
rect 1360 9260 2245 9300
rect 2285 9260 3175 9300
rect 3215 9260 6700 9300
rect 6740 9260 7620 9300
rect 7660 9260 7700 9300
rect -37190 9240 7700 9260
rect -37190 9235 1320 9240
rect -38770 9225 1320 9235
rect -38770 9190 -38755 9225
rect -38720 9190 -38710 9225
rect -38675 9190 -38665 9225
rect -38630 9190 -38620 9225
rect -38585 9190 -38575 9225
rect -38540 9190 -38530 9225
rect -38495 9190 -38485 9225
rect -38450 9190 -38440 9225
rect -38405 9190 -38395 9225
rect -38360 9190 -38350 9225
rect -38315 9190 -38305 9225
rect -38270 9190 -38260 9225
rect -38225 9190 -38215 9225
rect -38180 9190 -38170 9225
rect -38135 9190 -38125 9225
rect -38090 9190 -38080 9225
rect -38045 9190 -38035 9225
rect -38000 9190 -37990 9225
rect -37955 9190 -37945 9225
rect -37910 9190 -37900 9225
rect -37865 9190 -37855 9225
rect -37820 9190 -37810 9225
rect -37775 9190 -37765 9225
rect -37730 9190 -37720 9225
rect -37685 9190 -37675 9225
rect -37640 9190 -37630 9225
rect -37595 9190 -37585 9225
rect -37550 9190 -37540 9225
rect -37505 9190 -37495 9225
rect -37460 9190 -37450 9225
rect -37415 9190 -37405 9225
rect -37370 9190 -37360 9225
rect -37325 9190 -37315 9225
rect -37280 9190 -37270 9225
rect -37235 9190 -37225 9225
rect -37190 9200 1320 9225
rect 1360 9200 2245 9240
rect 2285 9200 3175 9240
rect 3215 9200 6700 9240
rect 6740 9200 7620 9240
rect 7660 9200 7700 9240
rect -37190 9190 7700 9200
rect -38770 9180 7700 9190
rect -38770 9145 -38755 9180
rect -38720 9145 -38710 9180
rect -38675 9145 -38665 9180
rect -38630 9145 -38620 9180
rect -38585 9145 -38575 9180
rect -38540 9145 -38530 9180
rect -38495 9145 -38485 9180
rect -38450 9145 -38440 9180
rect -38405 9145 -38395 9180
rect -38360 9145 -38350 9180
rect -38315 9145 -38305 9180
rect -38270 9145 -38260 9180
rect -38225 9145 -38215 9180
rect -38180 9145 -38170 9180
rect -38135 9145 -38125 9180
rect -38090 9145 -38080 9180
rect -38045 9145 -38035 9180
rect -38000 9145 -37990 9180
rect -37955 9145 -37945 9180
rect -37910 9145 -37900 9180
rect -37865 9145 -37855 9180
rect -37820 9145 -37810 9180
rect -37775 9145 -37765 9180
rect -37730 9145 -37720 9180
rect -37685 9145 -37675 9180
rect -37640 9145 -37630 9180
rect -37595 9145 -37585 9180
rect -37550 9145 -37540 9180
rect -37505 9145 -37495 9180
rect -37460 9145 -37450 9180
rect -37415 9145 -37405 9180
rect -37370 9145 -37360 9180
rect -37325 9145 -37315 9180
rect -37280 9145 -37270 9180
rect -37235 9145 -37225 9180
rect -37190 9175 7700 9180
rect -37190 9145 1320 9175
rect -38770 9135 1320 9145
rect 1360 9135 2245 9175
rect 2285 9135 3175 9175
rect 3215 9135 6700 9175
rect 6740 9135 7620 9175
rect 7660 9135 7700 9175
rect -38770 9100 -38755 9135
rect -38720 9100 -38710 9135
rect -38675 9100 -38665 9135
rect -38630 9100 -38620 9135
rect -38585 9100 -38575 9135
rect -38540 9100 -38530 9135
rect -38495 9100 -38485 9135
rect -38450 9100 -38440 9135
rect -38405 9100 -38395 9135
rect -38360 9100 -38350 9135
rect -38315 9100 -38305 9135
rect -38270 9100 -38260 9135
rect -38225 9100 -38215 9135
rect -38180 9100 -38170 9135
rect -38135 9100 -38125 9135
rect -38090 9100 -38080 9135
rect -38045 9100 -38035 9135
rect -38000 9100 -37990 9135
rect -37955 9100 -37945 9135
rect -37910 9100 -37900 9135
rect -37865 9100 -37855 9135
rect -37820 9100 -37810 9135
rect -37775 9100 -37765 9135
rect -37730 9100 -37720 9135
rect -37685 9100 -37675 9135
rect -37640 9100 -37630 9135
rect -37595 9100 -37585 9135
rect -37550 9100 -37540 9135
rect -37505 9100 -37495 9135
rect -37460 9100 -37450 9135
rect -37415 9100 -37405 9135
rect -37370 9100 -37360 9135
rect -37325 9100 -37315 9135
rect -37280 9100 -37270 9135
rect -37235 9100 -37225 9135
rect -37190 9105 7700 9135
rect -37190 9100 1320 9105
rect -38770 9090 1320 9100
rect -38770 9055 -38755 9090
rect -38720 9055 -38710 9090
rect -38675 9055 -38665 9090
rect -38630 9055 -38620 9090
rect -38585 9055 -38575 9090
rect -38540 9055 -38530 9090
rect -38495 9055 -38485 9090
rect -38450 9055 -38440 9090
rect -38405 9055 -38395 9090
rect -38360 9055 -38350 9090
rect -38315 9055 -38305 9090
rect -38270 9055 -38260 9090
rect -38225 9055 -38215 9090
rect -38180 9055 -38170 9090
rect -38135 9055 -38125 9090
rect -38090 9055 -38080 9090
rect -38045 9055 -38035 9090
rect -38000 9055 -37990 9090
rect -37955 9055 -37945 9090
rect -37910 9055 -37900 9090
rect -37865 9055 -37855 9090
rect -37820 9055 -37810 9090
rect -37775 9055 -37765 9090
rect -37730 9055 -37720 9090
rect -37685 9055 -37675 9090
rect -37640 9055 -37630 9090
rect -37595 9055 -37585 9090
rect -37550 9055 -37540 9090
rect -37505 9055 -37495 9090
rect -37460 9055 -37450 9090
rect -37415 9055 -37405 9090
rect -37370 9055 -37360 9090
rect -37325 9055 -37315 9090
rect -37280 9055 -37270 9090
rect -37235 9055 -37225 9090
rect -37190 9065 1320 9090
rect 1360 9065 2245 9105
rect 2285 9065 3175 9105
rect 3215 9065 6700 9105
rect 6740 9065 7620 9105
rect 7660 9065 7700 9105
rect -37190 9055 7700 9065
rect -38770 9045 7700 9055
rect -38770 9010 -38755 9045
rect -38720 9010 -38710 9045
rect -38675 9010 -38665 9045
rect -38630 9010 -38620 9045
rect -38585 9010 -38575 9045
rect -38540 9010 -38530 9045
rect -38495 9010 -38485 9045
rect -38450 9010 -38440 9045
rect -38405 9010 -38395 9045
rect -38360 9010 -38350 9045
rect -38315 9010 -38305 9045
rect -38270 9010 -38260 9045
rect -38225 9010 -38215 9045
rect -38180 9010 -38170 9045
rect -38135 9010 -38125 9045
rect -38090 9010 -38080 9045
rect -38045 9010 -38035 9045
rect -38000 9010 -37990 9045
rect -37955 9010 -37945 9045
rect -37910 9010 -37900 9045
rect -37865 9010 -37855 9045
rect -37820 9010 -37810 9045
rect -37775 9010 -37765 9045
rect -37730 9010 -37720 9045
rect -37685 9010 -37675 9045
rect -37640 9010 -37630 9045
rect -37595 9010 -37585 9045
rect -37550 9010 -37540 9045
rect -37505 9010 -37495 9045
rect -37460 9010 -37450 9045
rect -37415 9010 -37405 9045
rect -37370 9010 -37360 9045
rect -37325 9010 -37315 9045
rect -37280 9010 -37270 9045
rect -37235 9010 -37225 9045
rect -37190 9035 7700 9045
rect -37190 9010 1320 9035
rect -38770 9000 1320 9010
rect -38770 8965 -38755 9000
rect -38720 8965 -38710 9000
rect -38675 8965 -38665 9000
rect -38630 8965 -38620 9000
rect -38585 8965 -38575 9000
rect -38540 8965 -38530 9000
rect -38495 8965 -38485 9000
rect -38450 8965 -38440 9000
rect -38405 8965 -38395 9000
rect -38360 8965 -38350 9000
rect -38315 8965 -38305 9000
rect -38270 8965 -38260 9000
rect -38225 8965 -38215 9000
rect -38180 8965 -38170 9000
rect -38135 8965 -38125 9000
rect -38090 8965 -38080 9000
rect -38045 8965 -38035 9000
rect -38000 8965 -37990 9000
rect -37955 8965 -37945 9000
rect -37910 8965 -37900 9000
rect -37865 8965 -37855 9000
rect -37820 8965 -37810 9000
rect -37775 8965 -37765 9000
rect -37730 8965 -37720 9000
rect -37685 8965 -37675 9000
rect -37640 8965 -37630 9000
rect -37595 8965 -37585 9000
rect -37550 8965 -37540 9000
rect -37505 8965 -37495 9000
rect -37460 8965 -37450 9000
rect -37415 8965 -37405 9000
rect -37370 8965 -37360 9000
rect -37325 8965 -37315 9000
rect -37280 8965 -37270 9000
rect -37235 8965 -37225 9000
rect -37190 8995 1320 9000
rect 1360 8995 2245 9035
rect 2285 8995 3175 9035
rect 3215 8995 6700 9035
rect 6740 8995 7620 9035
rect 7660 8995 7700 9035
rect -37190 8965 7700 8995
rect -38770 8955 1320 8965
rect -38770 8920 -38755 8955
rect -38720 8920 -38710 8955
rect -38675 8920 -38665 8955
rect -38630 8920 -38620 8955
rect -38585 8920 -38575 8955
rect -38540 8920 -38530 8955
rect -38495 8920 -38485 8955
rect -38450 8920 -38440 8955
rect -38405 8920 -38395 8955
rect -38360 8920 -38350 8955
rect -38315 8920 -38305 8955
rect -38270 8920 -38260 8955
rect -38225 8920 -38215 8955
rect -38180 8920 -38170 8955
rect -38135 8920 -38125 8955
rect -38090 8920 -38080 8955
rect -38045 8920 -38035 8955
rect -38000 8920 -37990 8955
rect -37955 8920 -37945 8955
rect -37910 8920 -37900 8955
rect -37865 8920 -37855 8955
rect -37820 8920 -37810 8955
rect -37775 8920 -37765 8955
rect -37730 8920 -37720 8955
rect -37685 8920 -37675 8955
rect -37640 8920 -37630 8955
rect -37595 8920 -37585 8955
rect -37550 8920 -37540 8955
rect -37505 8920 -37495 8955
rect -37460 8920 -37450 8955
rect -37415 8920 -37405 8955
rect -37370 8920 -37360 8955
rect -37325 8920 -37315 8955
rect -37280 8920 -37270 8955
rect -37235 8920 -37225 8955
rect -37190 8925 1320 8955
rect 1360 8925 2245 8965
rect 2285 8925 3175 8965
rect 3215 8925 6700 8965
rect 6740 8925 7620 8965
rect 7660 8925 7700 8965
rect 31290 9640 31305 9675
rect 31340 9640 31350 9675
rect 31385 9640 31395 9675
rect 31430 9640 31440 9675
rect 31475 9640 31485 9675
rect 31520 9640 31530 9675
rect 31565 9640 31575 9675
rect 31610 9640 31620 9675
rect 31655 9640 31665 9675
rect 31700 9640 31710 9675
rect 31745 9640 31755 9675
rect 31790 9640 31800 9675
rect 31835 9640 31845 9675
rect 31880 9640 31890 9675
rect 31925 9640 31935 9675
rect 31970 9640 31980 9675
rect 32015 9640 32025 9675
rect 32060 9640 32070 9675
rect 32105 9640 32115 9675
rect 32150 9640 32160 9675
rect 32195 9640 32205 9675
rect 32240 9640 32250 9675
rect 32285 9640 32295 9675
rect 32330 9640 32340 9675
rect 32375 9640 32385 9675
rect 32420 9640 32430 9675
rect 32465 9640 32475 9675
rect 32510 9640 32520 9675
rect 32555 9640 32565 9675
rect 32600 9640 32610 9675
rect 32645 9640 32655 9675
rect 32690 9640 32700 9675
rect 32735 9640 32745 9675
rect 32780 9640 32790 9675
rect 32825 9640 32835 9675
rect 32870 9640 35620 9675
rect 31290 9630 35620 9640
rect 31290 9595 31305 9630
rect 31340 9595 31350 9630
rect 31385 9595 31395 9630
rect 31430 9595 31440 9630
rect 31475 9595 31485 9630
rect 31520 9595 31530 9630
rect 31565 9595 31575 9630
rect 31610 9595 31620 9630
rect 31655 9595 31665 9630
rect 31700 9595 31710 9630
rect 31745 9595 31755 9630
rect 31790 9595 31800 9630
rect 31835 9595 31845 9630
rect 31880 9595 31890 9630
rect 31925 9595 31935 9630
rect 31970 9595 31980 9630
rect 32015 9595 32025 9630
rect 32060 9595 32070 9630
rect 32105 9595 32115 9630
rect 32150 9595 32160 9630
rect 32195 9595 32205 9630
rect 32240 9595 32250 9630
rect 32285 9595 32295 9630
rect 32330 9595 32340 9630
rect 32375 9595 32385 9630
rect 32420 9595 32430 9630
rect 32465 9595 32475 9630
rect 32510 9595 32520 9630
rect 32555 9595 32565 9630
rect 32600 9595 32610 9630
rect 32645 9595 32655 9630
rect 32690 9595 32700 9630
rect 32735 9595 32745 9630
rect 32780 9595 32790 9630
rect 32825 9595 32835 9630
rect 32870 9595 35620 9630
rect 31290 9585 35620 9595
rect 31290 9550 31305 9585
rect 31340 9550 31350 9585
rect 31385 9550 31395 9585
rect 31430 9550 31440 9585
rect 31475 9550 31485 9585
rect 31520 9550 31530 9585
rect 31565 9550 31575 9585
rect 31610 9550 31620 9585
rect 31655 9550 31665 9585
rect 31700 9550 31710 9585
rect 31745 9550 31755 9585
rect 31790 9550 31800 9585
rect 31835 9550 31845 9585
rect 31880 9550 31890 9585
rect 31925 9550 31935 9585
rect 31970 9550 31980 9585
rect 32015 9550 32025 9585
rect 32060 9550 32070 9585
rect 32105 9550 32115 9585
rect 32150 9550 32160 9585
rect 32195 9550 32205 9585
rect 32240 9550 32250 9585
rect 32285 9550 32295 9585
rect 32330 9550 32340 9585
rect 32375 9550 32385 9585
rect 32420 9550 32430 9585
rect 32465 9550 32475 9585
rect 32510 9550 32520 9585
rect 32555 9550 32565 9585
rect 32600 9550 32610 9585
rect 32645 9550 32655 9585
rect 32690 9550 32700 9585
rect 32735 9550 32745 9585
rect 32780 9550 32790 9585
rect 32825 9550 32835 9585
rect 32870 9550 35620 9585
rect 31290 9540 35620 9550
rect 31290 9505 31305 9540
rect 31340 9505 31350 9540
rect 31385 9505 31395 9540
rect 31430 9505 31440 9540
rect 31475 9505 31485 9540
rect 31520 9505 31530 9540
rect 31565 9505 31575 9540
rect 31610 9505 31620 9540
rect 31655 9505 31665 9540
rect 31700 9505 31710 9540
rect 31745 9505 31755 9540
rect 31790 9505 31800 9540
rect 31835 9505 31845 9540
rect 31880 9505 31890 9540
rect 31925 9505 31935 9540
rect 31970 9505 31980 9540
rect 32015 9505 32025 9540
rect 32060 9505 32070 9540
rect 32105 9505 32115 9540
rect 32150 9505 32160 9540
rect 32195 9505 32205 9540
rect 32240 9505 32250 9540
rect 32285 9505 32295 9540
rect 32330 9505 32340 9540
rect 32375 9505 32385 9540
rect 32420 9505 32430 9540
rect 32465 9505 32475 9540
rect 32510 9505 32520 9540
rect 32555 9505 32565 9540
rect 32600 9505 32610 9540
rect 32645 9505 32655 9540
rect 32690 9505 32700 9540
rect 32735 9505 32745 9540
rect 32780 9505 32790 9540
rect 32825 9505 32835 9540
rect 32870 9505 35620 9540
rect 31290 9495 35620 9505
rect 31290 9460 31305 9495
rect 31340 9460 31350 9495
rect 31385 9460 31395 9495
rect 31430 9460 31440 9495
rect 31475 9460 31485 9495
rect 31520 9460 31530 9495
rect 31565 9460 31575 9495
rect 31610 9460 31620 9495
rect 31655 9460 31665 9495
rect 31700 9460 31710 9495
rect 31745 9460 31755 9495
rect 31790 9460 31800 9495
rect 31835 9460 31845 9495
rect 31880 9460 31890 9495
rect 31925 9460 31935 9495
rect 31970 9460 31980 9495
rect 32015 9460 32025 9495
rect 32060 9460 32070 9495
rect 32105 9460 32115 9495
rect 32150 9460 32160 9495
rect 32195 9460 32205 9495
rect 32240 9460 32250 9495
rect 32285 9460 32295 9495
rect 32330 9460 32340 9495
rect 32375 9460 32385 9495
rect 32420 9460 32430 9495
rect 32465 9460 32475 9495
rect 32510 9460 32520 9495
rect 32555 9460 32565 9495
rect 32600 9460 32610 9495
rect 32645 9460 32655 9495
rect 32690 9460 32700 9495
rect 32735 9460 32745 9495
rect 32780 9460 32790 9495
rect 32825 9460 32835 9495
rect 32870 9460 35620 9495
rect 31290 9450 35620 9460
rect 31290 9415 31305 9450
rect 31340 9415 31350 9450
rect 31385 9415 31395 9450
rect 31430 9415 31440 9450
rect 31475 9415 31485 9450
rect 31520 9415 31530 9450
rect 31565 9415 31575 9450
rect 31610 9415 31620 9450
rect 31655 9415 31665 9450
rect 31700 9415 31710 9450
rect 31745 9415 31755 9450
rect 31790 9415 31800 9450
rect 31835 9415 31845 9450
rect 31880 9415 31890 9450
rect 31925 9415 31935 9450
rect 31970 9415 31980 9450
rect 32015 9415 32025 9450
rect 32060 9415 32070 9450
rect 32105 9415 32115 9450
rect 32150 9415 32160 9450
rect 32195 9415 32205 9450
rect 32240 9415 32250 9450
rect 32285 9415 32295 9450
rect 32330 9415 32340 9450
rect 32375 9415 32385 9450
rect 32420 9415 32430 9450
rect 32465 9415 32475 9450
rect 32510 9415 32520 9450
rect 32555 9415 32565 9450
rect 32600 9415 32610 9450
rect 32645 9415 32655 9450
rect 32690 9415 32700 9450
rect 32735 9415 32745 9450
rect 32780 9415 32790 9450
rect 32825 9415 32835 9450
rect 32870 9415 35620 9450
rect 31290 9405 35620 9415
rect 31290 9370 31305 9405
rect 31340 9370 31350 9405
rect 31385 9370 31395 9405
rect 31430 9370 31440 9405
rect 31475 9370 31485 9405
rect 31520 9370 31530 9405
rect 31565 9370 31575 9405
rect 31610 9370 31620 9405
rect 31655 9370 31665 9405
rect 31700 9370 31710 9405
rect 31745 9370 31755 9405
rect 31790 9370 31800 9405
rect 31835 9370 31845 9405
rect 31880 9370 31890 9405
rect 31925 9370 31935 9405
rect 31970 9370 31980 9405
rect 32015 9370 32025 9405
rect 32060 9370 32070 9405
rect 32105 9370 32115 9405
rect 32150 9370 32160 9405
rect 32195 9370 32205 9405
rect 32240 9370 32250 9405
rect 32285 9370 32295 9405
rect 32330 9370 32340 9405
rect 32375 9370 32385 9405
rect 32420 9370 32430 9405
rect 32465 9370 32475 9405
rect 32510 9370 32520 9405
rect 32555 9370 32565 9405
rect 32600 9370 32610 9405
rect 32645 9370 32655 9405
rect 32690 9370 32700 9405
rect 32735 9370 32745 9405
rect 32780 9370 32790 9405
rect 32825 9370 32835 9405
rect 32870 9370 35620 9405
rect 31290 9360 35620 9370
rect 31290 9325 31305 9360
rect 31340 9325 31350 9360
rect 31385 9325 31395 9360
rect 31430 9325 31440 9360
rect 31475 9325 31485 9360
rect 31520 9325 31530 9360
rect 31565 9325 31575 9360
rect 31610 9325 31620 9360
rect 31655 9325 31665 9360
rect 31700 9325 31710 9360
rect 31745 9325 31755 9360
rect 31790 9325 31800 9360
rect 31835 9325 31845 9360
rect 31880 9325 31890 9360
rect 31925 9325 31935 9360
rect 31970 9325 31980 9360
rect 32015 9325 32025 9360
rect 32060 9325 32070 9360
rect 32105 9325 32115 9360
rect 32150 9325 32160 9360
rect 32195 9325 32205 9360
rect 32240 9325 32250 9360
rect 32285 9325 32295 9360
rect 32330 9325 32340 9360
rect 32375 9325 32385 9360
rect 32420 9325 32430 9360
rect 32465 9325 32475 9360
rect 32510 9325 32520 9360
rect 32555 9325 32565 9360
rect 32600 9325 32610 9360
rect 32645 9325 32655 9360
rect 32690 9325 32700 9360
rect 32735 9325 32745 9360
rect 32780 9325 32790 9360
rect 32825 9325 32835 9360
rect 32870 9325 35620 9360
rect 31290 9315 35620 9325
rect 31290 9280 31305 9315
rect 31340 9280 31350 9315
rect 31385 9280 31395 9315
rect 31430 9280 31440 9315
rect 31475 9280 31485 9315
rect 31520 9280 31530 9315
rect 31565 9280 31575 9315
rect 31610 9280 31620 9315
rect 31655 9280 31665 9315
rect 31700 9280 31710 9315
rect 31745 9280 31755 9315
rect 31790 9280 31800 9315
rect 31835 9280 31845 9315
rect 31880 9280 31890 9315
rect 31925 9280 31935 9315
rect 31970 9280 31980 9315
rect 32015 9280 32025 9315
rect 32060 9280 32070 9315
rect 32105 9280 32115 9315
rect 32150 9280 32160 9315
rect 32195 9280 32205 9315
rect 32240 9280 32250 9315
rect 32285 9280 32295 9315
rect 32330 9280 32340 9315
rect 32375 9280 32385 9315
rect 32420 9280 32430 9315
rect 32465 9280 32475 9315
rect 32510 9280 32520 9315
rect 32555 9280 32565 9315
rect 32600 9280 32610 9315
rect 32645 9280 32655 9315
rect 32690 9280 32700 9315
rect 32735 9280 32745 9315
rect 32780 9280 32790 9315
rect 32825 9280 32835 9315
rect 32870 9280 35620 9315
rect 31290 9270 35620 9280
rect 31290 9235 31305 9270
rect 31340 9235 31350 9270
rect 31385 9235 31395 9270
rect 31430 9235 31440 9270
rect 31475 9235 31485 9270
rect 31520 9235 31530 9270
rect 31565 9235 31575 9270
rect 31610 9235 31620 9270
rect 31655 9235 31665 9270
rect 31700 9235 31710 9270
rect 31745 9235 31755 9270
rect 31790 9235 31800 9270
rect 31835 9235 31845 9270
rect 31880 9235 31890 9270
rect 31925 9235 31935 9270
rect 31970 9235 31980 9270
rect 32015 9235 32025 9270
rect 32060 9235 32070 9270
rect 32105 9235 32115 9270
rect 32150 9235 32160 9270
rect 32195 9235 32205 9270
rect 32240 9235 32250 9270
rect 32285 9235 32295 9270
rect 32330 9235 32340 9270
rect 32375 9235 32385 9270
rect 32420 9235 32430 9270
rect 32465 9235 32475 9270
rect 32510 9235 32520 9270
rect 32555 9235 32565 9270
rect 32600 9235 32610 9270
rect 32645 9235 32655 9270
rect 32690 9235 32700 9270
rect 32735 9235 32745 9270
rect 32780 9235 32790 9270
rect 32825 9235 32835 9270
rect 32870 9235 35620 9270
rect 31290 9225 35620 9235
rect 31290 9190 31305 9225
rect 31340 9190 31350 9225
rect 31385 9190 31395 9225
rect 31430 9190 31440 9225
rect 31475 9190 31485 9225
rect 31520 9190 31530 9225
rect 31565 9190 31575 9225
rect 31610 9190 31620 9225
rect 31655 9190 31665 9225
rect 31700 9190 31710 9225
rect 31745 9190 31755 9225
rect 31790 9190 31800 9225
rect 31835 9190 31845 9225
rect 31880 9190 31890 9225
rect 31925 9190 31935 9225
rect 31970 9190 31980 9225
rect 32015 9190 32025 9225
rect 32060 9190 32070 9225
rect 32105 9190 32115 9225
rect 32150 9190 32160 9225
rect 32195 9190 32205 9225
rect 32240 9190 32250 9225
rect 32285 9190 32295 9225
rect 32330 9190 32340 9225
rect 32375 9190 32385 9225
rect 32420 9190 32430 9225
rect 32465 9190 32475 9225
rect 32510 9190 32520 9225
rect 32555 9190 32565 9225
rect 32600 9190 32610 9225
rect 32645 9190 32655 9225
rect 32690 9190 32700 9225
rect 32735 9190 32745 9225
rect 32780 9190 32790 9225
rect 32825 9190 32835 9225
rect 32870 9190 35620 9225
rect 31290 9180 35620 9190
rect 31290 9145 31305 9180
rect 31340 9145 31350 9180
rect 31385 9145 31395 9180
rect 31430 9145 31440 9180
rect 31475 9145 31485 9180
rect 31520 9145 31530 9180
rect 31565 9145 31575 9180
rect 31610 9145 31620 9180
rect 31655 9145 31665 9180
rect 31700 9145 31710 9180
rect 31745 9145 31755 9180
rect 31790 9145 31800 9180
rect 31835 9145 31845 9180
rect 31880 9145 31890 9180
rect 31925 9145 31935 9180
rect 31970 9145 31980 9180
rect 32015 9145 32025 9180
rect 32060 9145 32070 9180
rect 32105 9145 32115 9180
rect 32150 9145 32160 9180
rect 32195 9145 32205 9180
rect 32240 9145 32250 9180
rect 32285 9145 32295 9180
rect 32330 9145 32340 9180
rect 32375 9145 32385 9180
rect 32420 9145 32430 9180
rect 32465 9145 32475 9180
rect 32510 9145 32520 9180
rect 32555 9145 32565 9180
rect 32600 9145 32610 9180
rect 32645 9145 32655 9180
rect 32690 9145 32700 9180
rect 32735 9145 32745 9180
rect 32780 9145 32790 9180
rect 32825 9145 32835 9180
rect 32870 9145 35620 9180
rect 31290 9135 35620 9145
rect 31290 9100 31305 9135
rect 31340 9100 31350 9135
rect 31385 9100 31395 9135
rect 31430 9100 31440 9135
rect 31475 9100 31485 9135
rect 31520 9100 31530 9135
rect 31565 9100 31575 9135
rect 31610 9100 31620 9135
rect 31655 9100 31665 9135
rect 31700 9100 31710 9135
rect 31745 9100 31755 9135
rect 31790 9100 31800 9135
rect 31835 9100 31845 9135
rect 31880 9100 31890 9135
rect 31925 9100 31935 9135
rect 31970 9100 31980 9135
rect 32015 9100 32025 9135
rect 32060 9100 32070 9135
rect 32105 9100 32115 9135
rect 32150 9100 32160 9135
rect 32195 9100 32205 9135
rect 32240 9100 32250 9135
rect 32285 9100 32295 9135
rect 32330 9100 32340 9135
rect 32375 9100 32385 9135
rect 32420 9100 32430 9135
rect 32465 9100 32475 9135
rect 32510 9100 32520 9135
rect 32555 9100 32565 9135
rect 32600 9100 32610 9135
rect 32645 9100 32655 9135
rect 32690 9100 32700 9135
rect 32735 9100 32745 9135
rect 32780 9100 32790 9135
rect 32825 9100 32835 9135
rect 32870 9100 35620 9135
rect 31290 9090 35620 9100
rect 31290 9055 31305 9090
rect 31340 9055 31350 9090
rect 31385 9055 31395 9090
rect 31430 9055 31440 9090
rect 31475 9055 31485 9090
rect 31520 9055 31530 9090
rect 31565 9055 31575 9090
rect 31610 9055 31620 9090
rect 31655 9055 31665 9090
rect 31700 9055 31710 9090
rect 31745 9055 31755 9090
rect 31790 9055 31800 9090
rect 31835 9055 31845 9090
rect 31880 9055 31890 9090
rect 31925 9055 31935 9090
rect 31970 9055 31980 9090
rect 32015 9055 32025 9090
rect 32060 9055 32070 9090
rect 32105 9055 32115 9090
rect 32150 9055 32160 9090
rect 32195 9055 32205 9090
rect 32240 9055 32250 9090
rect 32285 9055 32295 9090
rect 32330 9055 32340 9090
rect 32375 9055 32385 9090
rect 32420 9055 32430 9090
rect 32465 9055 32475 9090
rect 32510 9055 32520 9090
rect 32555 9055 32565 9090
rect 32600 9055 32610 9090
rect 32645 9055 32655 9090
rect 32690 9055 32700 9090
rect 32735 9055 32745 9090
rect 32780 9055 32790 9090
rect 32825 9055 32835 9090
rect 32870 9055 35620 9090
rect 31290 9045 35620 9055
rect 31290 9010 31305 9045
rect 31340 9010 31350 9045
rect 31385 9010 31395 9045
rect 31430 9010 31440 9045
rect 31475 9010 31485 9045
rect 31520 9010 31530 9045
rect 31565 9010 31575 9045
rect 31610 9010 31620 9045
rect 31655 9010 31665 9045
rect 31700 9010 31710 9045
rect 31745 9010 31755 9045
rect 31790 9010 31800 9045
rect 31835 9010 31845 9045
rect 31880 9010 31890 9045
rect 31925 9010 31935 9045
rect 31970 9010 31980 9045
rect 32015 9010 32025 9045
rect 32060 9010 32070 9045
rect 32105 9010 32115 9045
rect 32150 9010 32160 9045
rect 32195 9010 32205 9045
rect 32240 9010 32250 9045
rect 32285 9010 32295 9045
rect 32330 9010 32340 9045
rect 32375 9010 32385 9045
rect 32420 9010 32430 9045
rect 32465 9010 32475 9045
rect 32510 9010 32520 9045
rect 32555 9010 32565 9045
rect 32600 9010 32610 9045
rect 32645 9010 32655 9045
rect 32690 9010 32700 9045
rect 32735 9010 32745 9045
rect 32780 9010 32790 9045
rect 32825 9010 32835 9045
rect 32870 9010 35620 9045
rect 31290 9000 35620 9010
rect 31290 8965 31305 9000
rect 31340 8965 31350 9000
rect 31385 8965 31395 9000
rect 31430 8965 31440 9000
rect 31475 8965 31485 9000
rect 31520 8965 31530 9000
rect 31565 8965 31575 9000
rect 31610 8965 31620 9000
rect 31655 8965 31665 9000
rect 31700 8965 31710 9000
rect 31745 8965 31755 9000
rect 31790 8965 31800 9000
rect 31835 8965 31845 9000
rect 31880 8965 31890 9000
rect 31925 8965 31935 9000
rect 31970 8965 31980 9000
rect 32015 8965 32025 9000
rect 32060 8965 32070 9000
rect 32105 8965 32115 9000
rect 32150 8965 32160 9000
rect 32195 8965 32205 9000
rect 32240 8965 32250 9000
rect 32285 8965 32295 9000
rect 32330 8965 32340 9000
rect 32375 8965 32385 9000
rect 32420 8965 32430 9000
rect 32465 8965 32475 9000
rect 32510 8965 32520 9000
rect 32555 8965 32565 9000
rect 32600 8965 32610 9000
rect 32645 8965 32655 9000
rect 32690 8965 32700 9000
rect 32735 8965 32745 9000
rect 32780 8965 32790 9000
rect 32825 8965 32835 9000
rect 32870 8965 35620 9000
rect 31290 8950 35620 8965
rect -37190 8920 7700 8925
rect -38770 8910 7700 8920
rect -38770 8875 -38755 8910
rect -38720 8875 -38710 8910
rect -38675 8875 -38665 8910
rect -38630 8875 -38620 8910
rect -38585 8875 -38575 8910
rect -38540 8875 -38530 8910
rect -38495 8875 -38485 8910
rect -38450 8875 -38440 8910
rect -38405 8875 -38395 8910
rect -38360 8875 -38350 8910
rect -38315 8875 -38305 8910
rect -38270 8875 -38260 8910
rect -38225 8875 -38215 8910
rect -38180 8875 -38170 8910
rect -38135 8875 -38125 8910
rect -38090 8875 -38080 8910
rect -38045 8875 -38035 8910
rect -38000 8875 -37990 8910
rect -37955 8875 -37945 8910
rect -37910 8875 -37900 8910
rect -37865 8875 -37855 8910
rect -37820 8875 -37810 8910
rect -37775 8875 -37765 8910
rect -37730 8875 -37720 8910
rect -37685 8875 -37675 8910
rect -37640 8875 -37630 8910
rect -37595 8875 -37585 8910
rect -37550 8875 -37540 8910
rect -37505 8875 -37495 8910
rect -37460 8875 -37450 8910
rect -37415 8875 -37405 8910
rect -37370 8875 -37360 8910
rect -37325 8875 -37315 8910
rect -37280 8875 -37270 8910
rect -37235 8875 -37225 8910
rect -37190 8900 7700 8910
rect -37190 8875 1320 8900
rect -38770 8865 1320 8875
rect -38770 8830 -38755 8865
rect -38720 8830 -38710 8865
rect -38675 8830 -38665 8865
rect -38630 8830 -38620 8865
rect -38585 8830 -38575 8865
rect -38540 8830 -38530 8865
rect -38495 8830 -38485 8865
rect -38450 8830 -38440 8865
rect -38405 8830 -38395 8865
rect -38360 8830 -38350 8865
rect -38315 8830 -38305 8865
rect -38270 8830 -38260 8865
rect -38225 8830 -38215 8865
rect -38180 8830 -38170 8865
rect -38135 8830 -38125 8865
rect -38090 8830 -38080 8865
rect -38045 8830 -38035 8865
rect -38000 8830 -37990 8865
rect -37955 8830 -37945 8865
rect -37910 8830 -37900 8865
rect -37865 8830 -37855 8865
rect -37820 8830 -37810 8865
rect -37775 8830 -37765 8865
rect -37730 8830 -37720 8865
rect -37685 8830 -37675 8865
rect -37640 8830 -37630 8865
rect -37595 8830 -37585 8865
rect -37550 8830 -37540 8865
rect -37505 8830 -37495 8865
rect -37460 8830 -37450 8865
rect -37415 8830 -37405 8865
rect -37370 8830 -37360 8865
rect -37325 8830 -37315 8865
rect -37280 8830 -37270 8865
rect -37235 8830 -37225 8865
rect -37190 8860 1320 8865
rect 1360 8860 2245 8900
rect 2285 8860 3175 8900
rect 3215 8860 6700 8900
rect 6740 8860 7620 8900
rect 7660 8860 7700 8900
rect -37190 8840 7700 8860
rect -37190 8830 1320 8840
rect -38770 8820 1320 8830
rect -38770 8785 -38755 8820
rect -38720 8785 -38710 8820
rect -38675 8785 -38665 8820
rect -38630 8785 -38620 8820
rect -38585 8785 -38575 8820
rect -38540 8785 -38530 8820
rect -38495 8785 -38485 8820
rect -38450 8785 -38440 8820
rect -38405 8785 -38395 8820
rect -38360 8785 -38350 8820
rect -38315 8785 -38305 8820
rect -38270 8785 -38260 8820
rect -38225 8785 -38215 8820
rect -38180 8785 -38170 8820
rect -38135 8785 -38125 8820
rect -38090 8785 -38080 8820
rect -38045 8785 -38035 8820
rect -38000 8785 -37990 8820
rect -37955 8785 -37945 8820
rect -37910 8785 -37900 8820
rect -37865 8785 -37855 8820
rect -37820 8785 -37810 8820
rect -37775 8785 -37765 8820
rect -37730 8785 -37720 8820
rect -37685 8785 -37675 8820
rect -37640 8785 -37630 8820
rect -37595 8785 -37585 8820
rect -37550 8785 -37540 8820
rect -37505 8785 -37495 8820
rect -37460 8785 -37450 8820
rect -37415 8785 -37405 8820
rect -37370 8785 -37360 8820
rect -37325 8785 -37315 8820
rect -37280 8785 -37270 8820
rect -37235 8785 -37225 8820
rect -37190 8800 1320 8820
rect 1360 8800 2245 8840
rect 2285 8800 3175 8840
rect 3215 8800 6700 8840
rect 6740 8800 7620 8840
rect 7660 8800 7700 8840
rect -37190 8785 7700 8800
rect -38770 8775 7700 8785
rect -38770 8740 -38755 8775
rect -38720 8740 -38710 8775
rect -38675 8740 -38665 8775
rect -38630 8740 -38620 8775
rect -38585 8740 -38575 8775
rect -38540 8740 -38530 8775
rect -38495 8740 -38485 8775
rect -38450 8740 -38440 8775
rect -38405 8740 -38395 8775
rect -38360 8740 -38350 8775
rect -38315 8740 -38305 8775
rect -38270 8740 -38260 8775
rect -38225 8740 -38215 8775
rect -38180 8740 -38170 8775
rect -38135 8740 -38125 8775
rect -38090 8740 -38080 8775
rect -38045 8740 -38035 8775
rect -38000 8740 -37990 8775
rect -37955 8740 -37945 8775
rect -37910 8740 -37900 8775
rect -37865 8740 -37855 8775
rect -37820 8740 -37810 8775
rect -37775 8740 -37765 8775
rect -37730 8740 -37720 8775
rect -37685 8740 -37675 8775
rect -37640 8740 -37630 8775
rect -37595 8740 -37585 8775
rect -37550 8740 -37540 8775
rect -37505 8740 -37495 8775
rect -37460 8740 -37450 8775
rect -37415 8740 -37405 8775
rect -37370 8740 -37360 8775
rect -37325 8740 -37315 8775
rect -37280 8740 -37270 8775
rect -37235 8740 -37225 8775
rect -37190 8740 1320 8775
rect -38770 8735 1320 8740
rect 1360 8735 2245 8775
rect 2285 8735 3175 8775
rect 3215 8735 6700 8775
rect 6740 8735 7620 8775
rect 7660 8735 7700 8775
rect -38770 8730 7700 8735
rect -38770 8695 -38755 8730
rect -38720 8695 -38710 8730
rect -38675 8695 -38665 8730
rect -38630 8695 -38620 8730
rect -38585 8695 -38575 8730
rect -38540 8695 -38530 8730
rect -38495 8695 -38485 8730
rect -38450 8695 -38440 8730
rect -38405 8695 -38395 8730
rect -38360 8695 -38350 8730
rect -38315 8695 -38305 8730
rect -38270 8695 -38260 8730
rect -38225 8695 -38215 8730
rect -38180 8695 -38170 8730
rect -38135 8695 -38125 8730
rect -38090 8695 -38080 8730
rect -38045 8695 -38035 8730
rect -38000 8695 -37990 8730
rect -37955 8695 -37945 8730
rect -37910 8695 -37900 8730
rect -37865 8695 -37855 8730
rect -37820 8695 -37810 8730
rect -37775 8695 -37765 8730
rect -37730 8695 -37720 8730
rect -37685 8695 -37675 8730
rect -37640 8695 -37630 8730
rect -37595 8695 -37585 8730
rect -37550 8695 -37540 8730
rect -37505 8695 -37495 8730
rect -37460 8695 -37450 8730
rect -37415 8695 -37405 8730
rect -37370 8695 -37360 8730
rect -37325 8695 -37315 8730
rect -37280 8695 -37270 8730
rect -37235 8695 -37225 8730
rect -37190 8705 7700 8730
rect -37190 8695 1320 8705
rect -38770 8685 1320 8695
rect -38770 8650 -38755 8685
rect -38720 8650 -38710 8685
rect -38675 8650 -38665 8685
rect -38630 8650 -38620 8685
rect -38585 8650 -38575 8685
rect -38540 8650 -38530 8685
rect -38495 8650 -38485 8685
rect -38450 8650 -38440 8685
rect -38405 8650 -38395 8685
rect -38360 8650 -38350 8685
rect -38315 8650 -38305 8685
rect -38270 8650 -38260 8685
rect -38225 8650 -38215 8685
rect -38180 8650 -38170 8685
rect -38135 8650 -38125 8685
rect -38090 8650 -38080 8685
rect -38045 8650 -38035 8685
rect -38000 8650 -37990 8685
rect -37955 8650 -37945 8685
rect -37910 8650 -37900 8685
rect -37865 8650 -37855 8685
rect -37820 8650 -37810 8685
rect -37775 8650 -37765 8685
rect -37730 8650 -37720 8685
rect -37685 8650 -37675 8685
rect -37640 8650 -37630 8685
rect -37595 8650 -37585 8685
rect -37550 8650 -37540 8685
rect -37505 8650 -37495 8685
rect -37460 8650 -37450 8685
rect -37415 8650 -37405 8685
rect -37370 8650 -37360 8685
rect -37325 8650 -37315 8685
rect -37280 8650 -37270 8685
rect -37235 8650 -37225 8685
rect -37190 8665 1320 8685
rect 1360 8665 2245 8705
rect 2285 8665 3175 8705
rect 3215 8665 6700 8705
rect 6740 8665 7620 8705
rect 7660 8665 7700 8705
rect -37190 8650 7700 8665
rect -38770 8640 7700 8650
rect -38770 8605 -38755 8640
rect -38720 8605 -38710 8640
rect -38675 8605 -38665 8640
rect -38630 8605 -38620 8640
rect -38585 8605 -38575 8640
rect -38540 8605 -38530 8640
rect -38495 8605 -38485 8640
rect -38450 8605 -38440 8640
rect -38405 8605 -38395 8640
rect -38360 8605 -38350 8640
rect -38315 8605 -38305 8640
rect -38270 8605 -38260 8640
rect -38225 8605 -38215 8640
rect -38180 8605 -38170 8640
rect -38135 8605 -38125 8640
rect -38090 8605 -38080 8640
rect -38045 8605 -38035 8640
rect -38000 8605 -37990 8640
rect -37955 8605 -37945 8640
rect -37910 8605 -37900 8640
rect -37865 8605 -37855 8640
rect -37820 8605 -37810 8640
rect -37775 8605 -37765 8640
rect -37730 8605 -37720 8640
rect -37685 8605 -37675 8640
rect -37640 8605 -37630 8640
rect -37595 8605 -37585 8640
rect -37550 8605 -37540 8640
rect -37505 8605 -37495 8640
rect -37460 8605 -37450 8640
rect -37415 8605 -37405 8640
rect -37370 8605 -37360 8640
rect -37325 8605 -37315 8640
rect -37280 8605 -37270 8640
rect -37235 8605 -37225 8640
rect -37190 8635 7700 8640
rect -37190 8605 1320 8635
rect -38770 8595 1320 8605
rect 1360 8595 2245 8635
rect 2285 8595 3175 8635
rect 3215 8595 6700 8635
rect 6740 8595 7620 8635
rect 7660 8595 7700 8635
rect -38770 8560 -38755 8595
rect -38720 8560 -38710 8595
rect -38675 8560 -38665 8595
rect -38630 8560 -38620 8595
rect -38585 8560 -38575 8595
rect -38540 8560 -38530 8595
rect -38495 8560 -38485 8595
rect -38450 8560 -38440 8595
rect -38405 8560 -38395 8595
rect -38360 8560 -38350 8595
rect -38315 8560 -38305 8595
rect -38270 8560 -38260 8595
rect -38225 8560 -38215 8595
rect -38180 8560 -38170 8595
rect -38135 8560 -38125 8595
rect -38090 8560 -38080 8595
rect -38045 8560 -38035 8595
rect -38000 8560 -37990 8595
rect -37955 8560 -37945 8595
rect -37910 8560 -37900 8595
rect -37865 8560 -37855 8595
rect -37820 8560 -37810 8595
rect -37775 8560 -37765 8595
rect -37730 8560 -37720 8595
rect -37685 8560 -37675 8595
rect -37640 8560 -37630 8595
rect -37595 8560 -37585 8595
rect -37550 8560 -37540 8595
rect -37505 8560 -37495 8595
rect -37460 8560 -37450 8595
rect -37415 8560 -37405 8595
rect -37370 8560 -37360 8595
rect -37325 8560 -37315 8595
rect -37280 8560 -37270 8595
rect -37235 8560 -37225 8595
rect -37190 8565 7700 8595
rect -37190 8560 1320 8565
rect -38770 8550 1320 8560
rect -38770 8515 -38755 8550
rect -38720 8515 -38710 8550
rect -38675 8515 -38665 8550
rect -38630 8515 -38620 8550
rect -38585 8515 -38575 8550
rect -38540 8515 -38530 8550
rect -38495 8515 -38485 8550
rect -38450 8515 -38440 8550
rect -38405 8515 -38395 8550
rect -38360 8515 -38350 8550
rect -38315 8515 -38305 8550
rect -38270 8515 -38260 8550
rect -38225 8515 -38215 8550
rect -38180 8515 -38170 8550
rect -38135 8515 -38125 8550
rect -38090 8515 -38080 8550
rect -38045 8515 -38035 8550
rect -38000 8515 -37990 8550
rect -37955 8515 -37945 8550
rect -37910 8515 -37900 8550
rect -37865 8515 -37855 8550
rect -37820 8515 -37810 8550
rect -37775 8515 -37765 8550
rect -37730 8515 -37720 8550
rect -37685 8515 -37675 8550
rect -37640 8515 -37630 8550
rect -37595 8515 -37585 8550
rect -37550 8515 -37540 8550
rect -37505 8515 -37495 8550
rect -37460 8515 -37450 8550
rect -37415 8515 -37405 8550
rect -37370 8515 -37360 8550
rect -37325 8515 -37315 8550
rect -37280 8515 -37270 8550
rect -37235 8515 -37225 8550
rect -37190 8525 1320 8550
rect 1360 8525 2245 8565
rect 2285 8525 3175 8565
rect 3215 8525 6700 8565
rect 6740 8525 7620 8565
rect 7660 8525 7700 8565
rect -37190 8515 7700 8525
rect -38770 8505 7700 8515
rect -38770 8470 -38755 8505
rect -38720 8470 -38710 8505
rect -38675 8470 -38665 8505
rect -38630 8470 -38620 8505
rect -38585 8470 -38575 8505
rect -38540 8470 -38530 8505
rect -38495 8470 -38485 8505
rect -38450 8470 -38440 8505
rect -38405 8470 -38395 8505
rect -38360 8470 -38350 8505
rect -38315 8470 -38305 8505
rect -38270 8470 -38260 8505
rect -38225 8470 -38215 8505
rect -38180 8470 -38170 8505
rect -38135 8470 -38125 8505
rect -38090 8470 -38080 8505
rect -38045 8470 -38035 8505
rect -38000 8470 -37990 8505
rect -37955 8470 -37945 8505
rect -37910 8470 -37900 8505
rect -37865 8470 -37855 8505
rect -37820 8470 -37810 8505
rect -37775 8470 -37765 8505
rect -37730 8470 -37720 8505
rect -37685 8470 -37675 8505
rect -37640 8470 -37630 8505
rect -37595 8470 -37585 8505
rect -37550 8470 -37540 8505
rect -37505 8470 -37495 8505
rect -37460 8470 -37450 8505
rect -37415 8470 -37405 8505
rect -37370 8470 -37360 8505
rect -37325 8470 -37315 8505
rect -37280 8470 -37270 8505
rect -37235 8470 -37225 8505
rect -37190 8500 7700 8505
rect -37190 8470 1320 8500
rect -38770 8460 1320 8470
rect 1360 8460 2245 8500
rect 2285 8460 3175 8500
rect 3215 8460 6700 8500
rect 6740 8460 7620 8500
rect 7660 8460 7700 8500
rect -38770 8425 -38755 8460
rect -38720 8425 -38710 8460
rect -38675 8425 -38665 8460
rect -38630 8425 -38620 8460
rect -38585 8425 -38575 8460
rect -38540 8425 -38530 8460
rect -38495 8425 -38485 8460
rect -38450 8425 -38440 8460
rect -38405 8425 -38395 8460
rect -38360 8425 -38350 8460
rect -38315 8425 -38305 8460
rect -38270 8425 -38260 8460
rect -38225 8425 -38215 8460
rect -38180 8425 -38170 8460
rect -38135 8425 -38125 8460
rect -38090 8425 -38080 8460
rect -38045 8425 -38035 8460
rect -38000 8425 -37990 8460
rect -37955 8425 -37945 8460
rect -37910 8425 -37900 8460
rect -37865 8425 -37855 8460
rect -37820 8425 -37810 8460
rect -37775 8425 -37765 8460
rect -37730 8425 -37720 8460
rect -37685 8425 -37675 8460
rect -37640 8425 -37630 8460
rect -37595 8425 -37585 8460
rect -37550 8425 -37540 8460
rect -37505 8425 -37495 8460
rect -37460 8425 -37450 8460
rect -37415 8425 -37405 8460
rect -37370 8425 -37360 8460
rect -37325 8425 -37315 8460
rect -37280 8425 -37270 8460
rect -37235 8425 -37225 8460
rect -37190 8440 7700 8460
rect -37190 8425 1320 8440
rect -38770 8415 1320 8425
rect -38770 8380 -38755 8415
rect -38720 8380 -38710 8415
rect -38675 8380 -38665 8415
rect -38630 8380 -38620 8415
rect -38585 8380 -38575 8415
rect -38540 8380 -38530 8415
rect -38495 8380 -38485 8415
rect -38450 8380 -38440 8415
rect -38405 8380 -38395 8415
rect -38360 8380 -38350 8415
rect -38315 8380 -38305 8415
rect -38270 8380 -38260 8415
rect -38225 8380 -38215 8415
rect -38180 8380 -38170 8415
rect -38135 8380 -38125 8415
rect -38090 8380 -38080 8415
rect -38045 8380 -38035 8415
rect -38000 8380 -37990 8415
rect -37955 8380 -37945 8415
rect -37910 8380 -37900 8415
rect -37865 8380 -37855 8415
rect -37820 8380 -37810 8415
rect -37775 8380 -37765 8415
rect -37730 8380 -37720 8415
rect -37685 8380 -37675 8415
rect -37640 8380 -37630 8415
rect -37595 8380 -37585 8415
rect -37550 8380 -37540 8415
rect -37505 8380 -37495 8415
rect -37460 8380 -37450 8415
rect -37415 8380 -37405 8415
rect -37370 8380 -37360 8415
rect -37325 8380 -37315 8415
rect -37280 8380 -37270 8415
rect -37235 8380 -37225 8415
rect -37190 8400 1320 8415
rect 1360 8400 2245 8440
rect 2285 8400 3175 8440
rect 3215 8400 6700 8440
rect 6740 8400 7620 8440
rect 7660 8400 7700 8440
rect -37190 8380 7700 8400
rect -38770 8375 7700 8380
rect -38770 8370 1320 8375
rect -38770 8335 -38755 8370
rect -38720 8335 -38710 8370
rect -38675 8335 -38665 8370
rect -38630 8335 -38620 8370
rect -38585 8335 -38575 8370
rect -38540 8335 -38530 8370
rect -38495 8335 -38485 8370
rect -38450 8335 -38440 8370
rect -38405 8335 -38395 8370
rect -38360 8335 -38350 8370
rect -38315 8335 -38305 8370
rect -38270 8335 -38260 8370
rect -38225 8335 -38215 8370
rect -38180 8335 -38170 8370
rect -38135 8335 -38125 8370
rect -38090 8335 -38080 8370
rect -38045 8335 -38035 8370
rect -38000 8335 -37990 8370
rect -37955 8335 -37945 8370
rect -37910 8335 -37900 8370
rect -37865 8335 -37855 8370
rect -37820 8335 -37810 8370
rect -37775 8335 -37765 8370
rect -37730 8335 -37720 8370
rect -37685 8335 -37675 8370
rect -37640 8335 -37630 8370
rect -37595 8335 -37585 8370
rect -37550 8335 -37540 8370
rect -37505 8335 -37495 8370
rect -37460 8335 -37450 8370
rect -37415 8335 -37405 8370
rect -37370 8335 -37360 8370
rect -37325 8335 -37315 8370
rect -37280 8335 -37270 8370
rect -37235 8335 -37225 8370
rect -37190 8335 1320 8370
rect 1360 8335 2245 8375
rect 2285 8335 3175 8375
rect 3215 8335 6700 8375
rect 6740 8335 7620 8375
rect 7660 8335 7700 8375
rect -38770 8325 7700 8335
rect -38770 8290 -38755 8325
rect -38720 8290 -38710 8325
rect -38675 8290 -38665 8325
rect -38630 8290 -38620 8325
rect -38585 8290 -38575 8325
rect -38540 8290 -38530 8325
rect -38495 8290 -38485 8325
rect -38450 8290 -38440 8325
rect -38405 8290 -38395 8325
rect -38360 8290 -38350 8325
rect -38315 8290 -38305 8325
rect -38270 8290 -38260 8325
rect -38225 8290 -38215 8325
rect -38180 8290 -38170 8325
rect -38135 8290 -38125 8325
rect -38090 8290 -38080 8325
rect -38045 8290 -38035 8325
rect -38000 8290 -37990 8325
rect -37955 8290 -37945 8325
rect -37910 8290 -37900 8325
rect -37865 8290 -37855 8325
rect -37820 8290 -37810 8325
rect -37775 8290 -37765 8325
rect -37730 8290 -37720 8325
rect -37685 8290 -37675 8325
rect -37640 8290 -37630 8325
rect -37595 8290 -37585 8325
rect -37550 8290 -37540 8325
rect -37505 8290 -37495 8325
rect -37460 8290 -37450 8325
rect -37415 8290 -37405 8325
rect -37370 8290 -37360 8325
rect -37325 8290 -37315 8325
rect -37280 8290 -37270 8325
rect -37235 8290 -37225 8325
rect -37190 8305 7700 8325
rect -37190 8290 1320 8305
rect -38770 8280 1320 8290
rect -38770 8245 -38755 8280
rect -38720 8245 -38710 8280
rect -38675 8245 -38665 8280
rect -38630 8245 -38620 8280
rect -38585 8245 -38575 8280
rect -38540 8245 -38530 8280
rect -38495 8245 -38485 8280
rect -38450 8245 -38440 8280
rect -38405 8245 -38395 8280
rect -38360 8245 -38350 8280
rect -38315 8245 -38305 8280
rect -38270 8245 -38260 8280
rect -38225 8245 -38215 8280
rect -38180 8245 -38170 8280
rect -38135 8245 -38125 8280
rect -38090 8245 -38080 8280
rect -38045 8245 -38035 8280
rect -38000 8245 -37990 8280
rect -37955 8245 -37945 8280
rect -37910 8245 -37900 8280
rect -37865 8245 -37855 8280
rect -37820 8245 -37810 8280
rect -37775 8245 -37765 8280
rect -37730 8245 -37720 8280
rect -37685 8245 -37675 8280
rect -37640 8245 -37630 8280
rect -37595 8245 -37585 8280
rect -37550 8245 -37540 8280
rect -37505 8245 -37495 8280
rect -37460 8245 -37450 8280
rect -37415 8245 -37405 8280
rect -37370 8245 -37360 8280
rect -37325 8245 -37315 8280
rect -37280 8245 -37270 8280
rect -37235 8245 -37225 8280
rect -37190 8265 1320 8280
rect 1360 8265 2245 8305
rect 2285 8265 3175 8305
rect 3215 8265 6700 8305
rect 6740 8265 7620 8305
rect 7660 8265 7700 8305
rect -37190 8245 7700 8265
rect -38770 8235 7700 8245
rect -38770 8200 -38755 8235
rect -38720 8200 -38710 8235
rect -38675 8200 -38665 8235
rect -38630 8200 -38620 8235
rect -38585 8200 -38575 8235
rect -38540 8200 -38530 8235
rect -38495 8200 -38485 8235
rect -38450 8200 -38440 8235
rect -38405 8200 -38395 8235
rect -38360 8200 -38350 8235
rect -38315 8200 -38305 8235
rect -38270 8200 -38260 8235
rect -38225 8200 -38215 8235
rect -38180 8200 -38170 8235
rect -38135 8200 -38125 8235
rect -38090 8200 -38080 8235
rect -38045 8200 -38035 8235
rect -38000 8200 -37990 8235
rect -37955 8200 -37945 8235
rect -37910 8200 -37900 8235
rect -37865 8200 -37855 8235
rect -37820 8200 -37810 8235
rect -37775 8200 -37765 8235
rect -37730 8200 -37720 8235
rect -37685 8200 -37675 8235
rect -37640 8200 -37630 8235
rect -37595 8200 -37585 8235
rect -37550 8200 -37540 8235
rect -37505 8200 -37495 8235
rect -37460 8200 -37450 8235
rect -37415 8200 -37405 8235
rect -37370 8200 -37360 8235
rect -37325 8200 -37315 8235
rect -37280 8200 -37270 8235
rect -37235 8200 -37225 8235
rect -37190 8200 1320 8235
rect -38770 8195 1320 8200
rect 1360 8195 2245 8235
rect 2285 8195 3175 8235
rect 3215 8195 6700 8235
rect 6740 8195 7620 8235
rect 7660 8195 7700 8235
rect -38770 8190 7700 8195
rect -38770 8155 -38755 8190
rect -38720 8155 -38710 8190
rect -38675 8155 -38665 8190
rect -38630 8155 -38620 8190
rect -38585 8155 -38575 8190
rect -38540 8155 -38530 8190
rect -38495 8155 -38485 8190
rect -38450 8155 -38440 8190
rect -38405 8155 -38395 8190
rect -38360 8155 -38350 8190
rect -38315 8155 -38305 8190
rect -38270 8155 -38260 8190
rect -38225 8155 -38215 8190
rect -38180 8155 -38170 8190
rect -38135 8155 -38125 8190
rect -38090 8155 -38080 8190
rect -38045 8155 -38035 8190
rect -38000 8155 -37990 8190
rect -37955 8155 -37945 8190
rect -37910 8155 -37900 8190
rect -37865 8155 -37855 8190
rect -37820 8155 -37810 8190
rect -37775 8155 -37765 8190
rect -37730 8155 -37720 8190
rect -37685 8155 -37675 8190
rect -37640 8155 -37630 8190
rect -37595 8155 -37585 8190
rect -37550 8155 -37540 8190
rect -37505 8155 -37495 8190
rect -37460 8155 -37450 8190
rect -37415 8155 -37405 8190
rect -37370 8155 -37360 8190
rect -37325 8155 -37315 8190
rect -37280 8155 -37270 8190
rect -37235 8155 -37225 8190
rect -37190 8165 7700 8190
rect -37190 8155 1320 8165
rect -38770 8145 1320 8155
rect -38770 8110 -38755 8145
rect -38720 8110 -38710 8145
rect -38675 8110 -38665 8145
rect -38630 8110 -38620 8145
rect -38585 8110 -38575 8145
rect -38540 8110 -38530 8145
rect -38495 8110 -38485 8145
rect -38450 8110 -38440 8145
rect -38405 8110 -38395 8145
rect -38360 8110 -38350 8145
rect -38315 8110 -38305 8145
rect -38270 8110 -38260 8145
rect -38225 8110 -38215 8145
rect -38180 8110 -38170 8145
rect -38135 8110 -38125 8145
rect -38090 8110 -38080 8145
rect -38045 8110 -38035 8145
rect -38000 8110 -37990 8145
rect -37955 8110 -37945 8145
rect -37910 8110 -37900 8145
rect -37865 8110 -37855 8145
rect -37820 8110 -37810 8145
rect -37775 8110 -37765 8145
rect -37730 8110 -37720 8145
rect -37685 8110 -37675 8145
rect -37640 8110 -37630 8145
rect -37595 8110 -37585 8145
rect -37550 8110 -37540 8145
rect -37505 8110 -37495 8145
rect -37460 8110 -37450 8145
rect -37415 8110 -37405 8145
rect -37370 8110 -37360 8145
rect -37325 8110 -37315 8145
rect -37280 8110 -37270 8145
rect -37235 8110 -37225 8145
rect -37190 8125 1320 8145
rect 1360 8125 2245 8165
rect 2285 8125 3175 8165
rect 3215 8125 6700 8165
rect 6740 8125 7620 8165
rect 7660 8125 7700 8165
rect -37190 8110 7700 8125
rect -38770 8105 7700 8110
rect -120 230 32890 240
rect -120 190 -80 230
rect -40 190 270 230
rect 310 190 620 230
rect 660 190 970 230
rect 1010 190 1320 230
rect 1360 190 1670 230
rect 1710 190 2020 230
rect 2060 190 2370 230
rect 2410 190 2720 230
rect 2760 190 3070 230
rect 3110 190 3420 230
rect 3460 190 3770 230
rect 3810 190 4120 230
rect 4160 190 4470 230
rect 4510 190 4820 230
rect 4860 190 5170 230
rect 5210 190 5520 230
rect 5560 190 5870 230
rect 5910 190 6220 230
rect 6260 190 6570 230
rect 6610 190 6920 230
rect 6960 190 7270 230
rect 7310 190 7620 230
rect 7660 190 7970 230
rect 8010 190 8320 230
rect 8360 190 8670 230
rect 8710 190 9020 230
rect 9060 220 32890 230
rect 9060 190 31305 220
rect -120 185 31305 190
rect 31340 185 31350 220
rect 31385 185 31395 220
rect 31430 185 31440 220
rect 31475 185 31485 220
rect 31520 185 31530 220
rect 31565 185 31575 220
rect 31610 185 31620 220
rect 31655 185 31665 220
rect 31700 185 31710 220
rect 31745 185 31755 220
rect 31790 185 31800 220
rect 31835 185 31845 220
rect 31880 185 31890 220
rect 31925 185 31935 220
rect 31970 185 31980 220
rect 32015 185 32025 220
rect 32060 185 32070 220
rect 32105 185 32115 220
rect 32150 185 32160 220
rect 32195 185 32205 220
rect 32240 185 32250 220
rect 32285 185 32295 220
rect 32330 185 32340 220
rect 32375 185 32385 220
rect 32420 185 32430 220
rect 32465 185 32475 220
rect 32510 185 32520 220
rect 32555 185 32565 220
rect 32600 185 32610 220
rect 32645 185 32655 220
rect 32690 185 32700 220
rect 32735 185 32745 220
rect 32780 185 32790 220
rect 32825 185 32835 220
rect 32870 185 32890 220
rect -120 175 32890 185
rect -120 165 31305 175
rect -120 125 -80 165
rect -40 125 270 165
rect 310 125 620 165
rect 660 125 970 165
rect 1010 125 1320 165
rect 1360 125 1670 165
rect 1710 125 2020 165
rect 2060 125 2370 165
rect 2410 125 2720 165
rect 2760 125 3070 165
rect 3110 125 3420 165
rect 3460 125 3770 165
rect 3810 125 4120 165
rect 4160 125 4470 165
rect 4510 125 4820 165
rect 4860 125 5170 165
rect 5210 125 5520 165
rect 5560 125 5870 165
rect 5910 125 6220 165
rect 6260 125 6570 165
rect 6610 125 6920 165
rect 6960 125 7270 165
rect 7310 125 7620 165
rect 7660 125 7970 165
rect 8010 125 8320 165
rect 8360 125 8670 165
rect 8710 125 9020 165
rect 9060 140 31305 165
rect 31340 140 31350 175
rect 31385 140 31395 175
rect 31430 140 31440 175
rect 31475 140 31485 175
rect 31520 140 31530 175
rect 31565 140 31575 175
rect 31610 140 31620 175
rect 31655 140 31665 175
rect 31700 140 31710 175
rect 31745 140 31755 175
rect 31790 140 31800 175
rect 31835 140 31845 175
rect 31880 140 31890 175
rect 31925 140 31935 175
rect 31970 140 31980 175
rect 32015 140 32025 175
rect 32060 140 32070 175
rect 32105 140 32115 175
rect 32150 140 32160 175
rect 32195 140 32205 175
rect 32240 140 32250 175
rect 32285 140 32295 175
rect 32330 140 32340 175
rect 32375 140 32385 175
rect 32420 140 32430 175
rect 32465 140 32475 175
rect 32510 140 32520 175
rect 32555 140 32565 175
rect 32600 140 32610 175
rect 32645 140 32655 175
rect 32690 140 32700 175
rect 32735 140 32745 175
rect 32780 140 32790 175
rect 32825 140 32835 175
rect 32870 140 32890 175
rect 9060 130 32890 140
rect 9060 125 31305 130
rect -120 95 31305 125
rect 31340 95 31350 130
rect 31385 95 31395 130
rect 31430 95 31440 130
rect 31475 95 31485 130
rect 31520 95 31530 130
rect 31565 95 31575 130
rect 31610 95 31620 130
rect 31655 95 31665 130
rect 31700 95 31710 130
rect 31745 95 31755 130
rect 31790 95 31800 130
rect 31835 95 31845 130
rect 31880 95 31890 130
rect 31925 95 31935 130
rect 31970 95 31980 130
rect 32015 95 32025 130
rect 32060 95 32070 130
rect 32105 95 32115 130
rect 32150 95 32160 130
rect 32195 95 32205 130
rect 32240 95 32250 130
rect 32285 95 32295 130
rect 32330 95 32340 130
rect 32375 95 32385 130
rect 32420 95 32430 130
rect 32465 95 32475 130
rect 32510 95 32520 130
rect 32555 95 32565 130
rect 32600 95 32610 130
rect 32645 95 32655 130
rect 32690 95 32700 130
rect 32735 95 32745 130
rect 32780 95 32790 130
rect 32825 95 32835 130
rect 32870 95 32890 130
rect -120 55 -80 95
rect -40 55 270 95
rect 310 55 620 95
rect 660 55 970 95
rect 1010 55 1320 95
rect 1360 55 1670 95
rect 1710 55 2020 95
rect 2060 55 2370 95
rect 2410 55 2720 95
rect 2760 55 3070 95
rect 3110 55 3420 95
rect 3460 55 3770 95
rect 3810 55 4120 95
rect 4160 55 4470 95
rect 4510 55 4820 95
rect 4860 55 5170 95
rect 5210 55 5520 95
rect 5560 55 5870 95
rect 5910 55 6220 95
rect 6260 55 6570 95
rect 6610 55 6920 95
rect 6960 55 7270 95
rect 7310 55 7620 95
rect 7660 55 7970 95
rect 8010 55 8320 95
rect 8360 55 8670 95
rect 8710 55 9020 95
rect 9060 85 32890 95
rect 9060 55 31305 85
rect -120 50 31305 55
rect 31340 50 31350 85
rect 31385 50 31395 85
rect 31430 50 31440 85
rect 31475 50 31485 85
rect 31520 50 31530 85
rect 31565 50 31575 85
rect 31610 50 31620 85
rect 31655 50 31665 85
rect 31700 50 31710 85
rect 31745 50 31755 85
rect 31790 50 31800 85
rect 31835 50 31845 85
rect 31880 50 31890 85
rect 31925 50 31935 85
rect 31970 50 31980 85
rect 32015 50 32025 85
rect 32060 50 32070 85
rect 32105 50 32115 85
rect 32150 50 32160 85
rect 32195 50 32205 85
rect 32240 50 32250 85
rect 32285 50 32295 85
rect 32330 50 32340 85
rect 32375 50 32385 85
rect 32420 50 32430 85
rect 32465 50 32475 85
rect 32510 50 32520 85
rect 32555 50 32565 85
rect 32600 50 32610 85
rect 32645 50 32655 85
rect 32690 50 32700 85
rect 32735 50 32745 85
rect 32780 50 32790 85
rect 32825 50 32835 85
rect 32870 50 32890 85
rect -120 40 32890 50
rect -120 25 31305 40
rect -120 -15 -80 25
rect -40 -15 270 25
rect 310 -15 620 25
rect 660 -15 970 25
rect 1010 -15 1320 25
rect 1360 -15 1670 25
rect 1710 -15 2020 25
rect 2060 -15 2370 25
rect 2410 -15 2720 25
rect 2760 -15 3070 25
rect 3110 -15 3420 25
rect 3460 -15 3770 25
rect 3810 -15 4120 25
rect 4160 -15 4470 25
rect 4510 -15 4820 25
rect 4860 -15 5170 25
rect 5210 -15 5520 25
rect 5560 -15 5870 25
rect 5910 -15 6220 25
rect 6260 -15 6570 25
rect 6610 -15 6920 25
rect 6960 -15 7270 25
rect 7310 -15 7620 25
rect 7660 -15 7970 25
rect 8010 -15 8320 25
rect 8360 -15 8670 25
rect 8710 -15 9020 25
rect 9060 5 31305 25
rect 31340 5 31350 40
rect 31385 5 31395 40
rect 31430 5 31440 40
rect 31475 5 31485 40
rect 31520 5 31530 40
rect 31565 5 31575 40
rect 31610 5 31620 40
rect 31655 5 31665 40
rect 31700 5 31710 40
rect 31745 5 31755 40
rect 31790 5 31800 40
rect 31835 5 31845 40
rect 31880 5 31890 40
rect 31925 5 31935 40
rect 31970 5 31980 40
rect 32015 5 32025 40
rect 32060 5 32070 40
rect 32105 5 32115 40
rect 32150 5 32160 40
rect 32195 5 32205 40
rect 32240 5 32250 40
rect 32285 5 32295 40
rect 32330 5 32340 40
rect 32375 5 32385 40
rect 32420 5 32430 40
rect 32465 5 32475 40
rect 32510 5 32520 40
rect 32555 5 32565 40
rect 32600 5 32610 40
rect 32645 5 32655 40
rect 32690 5 32700 40
rect 32735 5 32745 40
rect 32780 5 32790 40
rect 32825 5 32835 40
rect 32870 5 32890 40
rect 9060 -5 32890 5
rect 9060 -15 31305 -5
rect -120 -40 31305 -15
rect 31340 -40 31350 -5
rect 31385 -40 31395 -5
rect 31430 -40 31440 -5
rect 31475 -40 31485 -5
rect 31520 -40 31530 -5
rect 31565 -40 31575 -5
rect 31610 -40 31620 -5
rect 31655 -40 31665 -5
rect 31700 -40 31710 -5
rect 31745 -40 31755 -5
rect 31790 -40 31800 -5
rect 31835 -40 31845 -5
rect 31880 -40 31890 -5
rect 31925 -40 31935 -5
rect 31970 -40 31980 -5
rect 32015 -40 32025 -5
rect 32060 -40 32070 -5
rect 32105 -40 32115 -5
rect 32150 -40 32160 -5
rect 32195 -40 32205 -5
rect 32240 -40 32250 -5
rect 32285 -40 32295 -5
rect 32330 -40 32340 -5
rect 32375 -40 32385 -5
rect 32420 -40 32430 -5
rect 32465 -40 32475 -5
rect 32510 -40 32520 -5
rect 32555 -40 32565 -5
rect 32600 -40 32610 -5
rect 32645 -40 32655 -5
rect 32690 -40 32700 -5
rect 32735 -40 32745 -5
rect 32780 -40 32790 -5
rect 32825 -40 32835 -5
rect 32870 -40 32890 -5
rect -120 -45 32890 -40
rect -120 -85 -80 -45
rect -40 -85 270 -45
rect 310 -85 620 -45
rect 660 -85 970 -45
rect 1010 -85 1320 -45
rect 1360 -85 1670 -45
rect 1710 -85 2020 -45
rect 2060 -85 2370 -45
rect 2410 -85 2720 -45
rect 2760 -85 3070 -45
rect 3110 -85 3420 -45
rect 3460 -85 3770 -45
rect 3810 -85 4120 -45
rect 4160 -85 4470 -45
rect 4510 -85 4820 -45
rect 4860 -85 5170 -45
rect 5210 -85 5520 -45
rect 5560 -85 5870 -45
rect 5910 -85 6220 -45
rect 6260 -85 6570 -45
rect 6610 -85 6920 -45
rect 6960 -85 7270 -45
rect 7310 -85 7620 -45
rect 7660 -85 7970 -45
rect 8010 -85 8320 -45
rect 8360 -85 8670 -45
rect 8710 -85 9020 -45
rect 9060 -50 32890 -45
rect 9060 -85 31305 -50
rect 31340 -85 31350 -50
rect 31385 -85 31395 -50
rect 31430 -85 31440 -50
rect 31475 -85 31485 -50
rect 31520 -85 31530 -50
rect 31565 -85 31575 -50
rect 31610 -85 31620 -50
rect 31655 -85 31665 -50
rect 31700 -85 31710 -50
rect 31745 -85 31755 -50
rect 31790 -85 31800 -50
rect 31835 -85 31845 -50
rect 31880 -85 31890 -50
rect 31925 -85 31935 -50
rect 31970 -85 31980 -50
rect 32015 -85 32025 -50
rect 32060 -85 32070 -50
rect 32105 -85 32115 -50
rect 32150 -85 32160 -50
rect 32195 -85 32205 -50
rect 32240 -85 32250 -50
rect 32285 -85 32295 -50
rect 32330 -85 32340 -50
rect 32375 -85 32385 -50
rect 32420 -85 32430 -50
rect 32465 -85 32475 -50
rect 32510 -85 32520 -50
rect 32555 -85 32565 -50
rect 32600 -85 32610 -50
rect 32645 -85 32655 -50
rect 32690 -85 32700 -50
rect 32735 -85 32745 -50
rect 32780 -85 32790 -50
rect 32825 -85 32835 -50
rect 32870 -85 32890 -50
rect -120 -95 32890 -85
rect -120 -110 31305 -95
rect -120 -150 -80 -110
rect -40 -150 270 -110
rect 310 -150 620 -110
rect 660 -150 970 -110
rect 1010 -150 1320 -110
rect 1360 -150 1670 -110
rect 1710 -150 2020 -110
rect 2060 -150 2370 -110
rect 2410 -150 2720 -110
rect 2760 -150 3070 -110
rect 3110 -150 3420 -110
rect 3460 -150 3770 -110
rect 3810 -150 4120 -110
rect 4160 -150 4470 -110
rect 4510 -150 4820 -110
rect 4860 -150 5170 -110
rect 5210 -150 5520 -110
rect 5560 -150 5870 -110
rect 5910 -150 6220 -110
rect 6260 -150 6570 -110
rect 6610 -150 6920 -110
rect 6960 -150 7270 -110
rect 7310 -150 7620 -110
rect 7660 -150 7970 -110
rect 8010 -150 8320 -110
rect 8360 -150 8670 -110
rect 8710 -150 9020 -110
rect 9060 -130 31305 -110
rect 31340 -130 31350 -95
rect 31385 -130 31395 -95
rect 31430 -130 31440 -95
rect 31475 -130 31485 -95
rect 31520 -130 31530 -95
rect 31565 -130 31575 -95
rect 31610 -130 31620 -95
rect 31655 -130 31665 -95
rect 31700 -130 31710 -95
rect 31745 -130 31755 -95
rect 31790 -130 31800 -95
rect 31835 -130 31845 -95
rect 31880 -130 31890 -95
rect 31925 -130 31935 -95
rect 31970 -130 31980 -95
rect 32015 -130 32025 -95
rect 32060 -130 32070 -95
rect 32105 -130 32115 -95
rect 32150 -130 32160 -95
rect 32195 -130 32205 -95
rect 32240 -130 32250 -95
rect 32285 -130 32295 -95
rect 32330 -130 32340 -95
rect 32375 -130 32385 -95
rect 32420 -130 32430 -95
rect 32465 -130 32475 -95
rect 32510 -130 32520 -95
rect 32555 -130 32565 -95
rect 32600 -130 32610 -95
rect 32645 -130 32655 -95
rect 32690 -130 32700 -95
rect 32735 -130 32745 -95
rect 32780 -130 32790 -95
rect 32825 -130 32835 -95
rect 32870 -130 32890 -95
rect 9060 -140 32890 -130
rect 9060 -150 31305 -140
rect -120 -170 31305 -150
rect -120 -210 -80 -170
rect -40 -210 270 -170
rect 310 -210 620 -170
rect 660 -210 970 -170
rect 1010 -210 1320 -170
rect 1360 -210 1670 -170
rect 1710 -210 2020 -170
rect 2060 -210 2370 -170
rect 2410 -210 2720 -170
rect 2760 -210 3070 -170
rect 3110 -210 3420 -170
rect 3460 -210 3770 -170
rect 3810 -210 4120 -170
rect 4160 -210 4470 -170
rect 4510 -210 4820 -170
rect 4860 -210 5170 -170
rect 5210 -210 5520 -170
rect 5560 -210 5870 -170
rect 5910 -210 6220 -170
rect 6260 -210 6570 -170
rect 6610 -210 6920 -170
rect 6960 -210 7270 -170
rect 7310 -210 7620 -170
rect 7660 -210 7970 -170
rect 8010 -210 8320 -170
rect 8360 -210 8670 -170
rect 8710 -210 9020 -170
rect 9060 -175 31305 -170
rect 31340 -175 31350 -140
rect 31385 -175 31395 -140
rect 31430 -175 31440 -140
rect 31475 -175 31485 -140
rect 31520 -175 31530 -140
rect 31565 -175 31575 -140
rect 31610 -175 31620 -140
rect 31655 -175 31665 -140
rect 31700 -175 31710 -140
rect 31745 -175 31755 -140
rect 31790 -175 31800 -140
rect 31835 -175 31845 -140
rect 31880 -175 31890 -140
rect 31925 -175 31935 -140
rect 31970 -175 31980 -140
rect 32015 -175 32025 -140
rect 32060 -175 32070 -140
rect 32105 -175 32115 -140
rect 32150 -175 32160 -140
rect 32195 -175 32205 -140
rect 32240 -175 32250 -140
rect 32285 -175 32295 -140
rect 32330 -175 32340 -140
rect 32375 -175 32385 -140
rect 32420 -175 32430 -140
rect 32465 -175 32475 -140
rect 32510 -175 32520 -140
rect 32555 -175 32565 -140
rect 32600 -175 32610 -140
rect 32645 -175 32655 -140
rect 32690 -175 32700 -140
rect 32735 -175 32745 -140
rect 32780 -175 32790 -140
rect 32825 -175 32835 -140
rect 32870 -175 32890 -140
rect 9060 -185 32890 -175
rect 9060 -210 31305 -185
rect -120 -220 31305 -210
rect 31340 -220 31350 -185
rect 31385 -220 31395 -185
rect 31430 -220 31440 -185
rect 31475 -220 31485 -185
rect 31520 -220 31530 -185
rect 31565 -220 31575 -185
rect 31610 -220 31620 -185
rect 31655 -220 31665 -185
rect 31700 -220 31710 -185
rect 31745 -220 31755 -185
rect 31790 -220 31800 -185
rect 31835 -220 31845 -185
rect 31880 -220 31890 -185
rect 31925 -220 31935 -185
rect 31970 -220 31980 -185
rect 32015 -220 32025 -185
rect 32060 -220 32070 -185
rect 32105 -220 32115 -185
rect 32150 -220 32160 -185
rect 32195 -220 32205 -185
rect 32240 -220 32250 -185
rect 32285 -220 32295 -185
rect 32330 -220 32340 -185
rect 32375 -220 32385 -185
rect 32420 -220 32430 -185
rect 32465 -220 32475 -185
rect 32510 -220 32520 -185
rect 32555 -220 32565 -185
rect 32600 -220 32610 -185
rect 32645 -220 32655 -185
rect 32690 -220 32700 -185
rect 32735 -220 32745 -185
rect 32780 -220 32790 -185
rect 32825 -220 32835 -185
rect 32870 -220 32890 -185
rect -120 -230 32890 -220
rect -120 -235 31305 -230
rect -120 -275 -80 -235
rect -40 -275 270 -235
rect 310 -275 620 -235
rect 660 -275 970 -235
rect 1010 -275 1320 -235
rect 1360 -275 1670 -235
rect 1710 -275 2020 -235
rect 2060 -275 2370 -235
rect 2410 -275 2720 -235
rect 2760 -275 3070 -235
rect 3110 -275 3420 -235
rect 3460 -275 3770 -235
rect 3810 -275 4120 -235
rect 4160 -275 4470 -235
rect 4510 -275 4820 -235
rect 4860 -275 5170 -235
rect 5210 -275 5520 -235
rect 5560 -275 5870 -235
rect 5910 -275 6220 -235
rect 6260 -275 6570 -235
rect 6610 -275 6920 -235
rect 6960 -275 7270 -235
rect 7310 -275 7620 -235
rect 7660 -275 7970 -235
rect 8010 -275 8320 -235
rect 8360 -275 8670 -235
rect 8710 -275 9020 -235
rect 9060 -265 31305 -235
rect 31340 -265 31350 -230
rect 31385 -265 31395 -230
rect 31430 -265 31440 -230
rect 31475 -265 31485 -230
rect 31520 -265 31530 -230
rect 31565 -265 31575 -230
rect 31610 -265 31620 -230
rect 31655 -265 31665 -230
rect 31700 -265 31710 -230
rect 31745 -265 31755 -230
rect 31790 -265 31800 -230
rect 31835 -265 31845 -230
rect 31880 -265 31890 -230
rect 31925 -265 31935 -230
rect 31970 -265 31980 -230
rect 32015 -265 32025 -230
rect 32060 -265 32070 -230
rect 32105 -265 32115 -230
rect 32150 -265 32160 -230
rect 32195 -265 32205 -230
rect 32240 -265 32250 -230
rect 32285 -265 32295 -230
rect 32330 -265 32340 -230
rect 32375 -265 32385 -230
rect 32420 -265 32430 -230
rect 32465 -265 32475 -230
rect 32510 -265 32520 -230
rect 32555 -265 32565 -230
rect 32600 -265 32610 -230
rect 32645 -265 32655 -230
rect 32690 -265 32700 -230
rect 32735 -265 32745 -230
rect 32780 -265 32790 -230
rect 32825 -265 32835 -230
rect 32870 -265 32890 -230
rect 9060 -275 32890 -265
rect -120 -305 31305 -275
rect -120 -345 -80 -305
rect -40 -345 270 -305
rect 310 -345 620 -305
rect 660 -345 970 -305
rect 1010 -345 1320 -305
rect 1360 -345 1670 -305
rect 1710 -345 2020 -305
rect 2060 -345 2370 -305
rect 2410 -345 2720 -305
rect 2760 -345 3070 -305
rect 3110 -345 3420 -305
rect 3460 -345 3770 -305
rect 3810 -345 4120 -305
rect 4160 -345 4470 -305
rect 4510 -345 4820 -305
rect 4860 -345 5170 -305
rect 5210 -345 5520 -305
rect 5560 -345 5870 -305
rect 5910 -345 6220 -305
rect 6260 -345 6570 -305
rect 6610 -345 6920 -305
rect 6960 -345 7270 -305
rect 7310 -345 7620 -305
rect 7660 -345 7970 -305
rect 8010 -345 8320 -305
rect 8360 -345 8670 -305
rect 8710 -345 9020 -305
rect 9060 -310 31305 -305
rect 31340 -310 31350 -275
rect 31385 -310 31395 -275
rect 31430 -310 31440 -275
rect 31475 -310 31485 -275
rect 31520 -310 31530 -275
rect 31565 -310 31575 -275
rect 31610 -310 31620 -275
rect 31655 -310 31665 -275
rect 31700 -310 31710 -275
rect 31745 -310 31755 -275
rect 31790 -310 31800 -275
rect 31835 -310 31845 -275
rect 31880 -310 31890 -275
rect 31925 -310 31935 -275
rect 31970 -310 31980 -275
rect 32015 -310 32025 -275
rect 32060 -310 32070 -275
rect 32105 -310 32115 -275
rect 32150 -310 32160 -275
rect 32195 -310 32205 -275
rect 32240 -310 32250 -275
rect 32285 -310 32295 -275
rect 32330 -310 32340 -275
rect 32375 -310 32385 -275
rect 32420 -310 32430 -275
rect 32465 -310 32475 -275
rect 32510 -310 32520 -275
rect 32555 -310 32565 -275
rect 32600 -310 32610 -275
rect 32645 -310 32655 -275
rect 32690 -310 32700 -275
rect 32735 -310 32745 -275
rect 32780 -310 32790 -275
rect 32825 -310 32835 -275
rect 32870 -310 32890 -275
rect 9060 -320 32890 -310
rect 9060 -345 31305 -320
rect -120 -355 31305 -345
rect 31340 -355 31350 -320
rect 31385 -355 31395 -320
rect 31430 -355 31440 -320
rect 31475 -355 31485 -320
rect 31520 -355 31530 -320
rect 31565 -355 31575 -320
rect 31610 -355 31620 -320
rect 31655 -355 31665 -320
rect 31700 -355 31710 -320
rect 31745 -355 31755 -320
rect 31790 -355 31800 -320
rect 31835 -355 31845 -320
rect 31880 -355 31890 -320
rect 31925 -355 31935 -320
rect 31970 -355 31980 -320
rect 32015 -355 32025 -320
rect 32060 -355 32070 -320
rect 32105 -355 32115 -320
rect 32150 -355 32160 -320
rect 32195 -355 32205 -320
rect 32240 -355 32250 -320
rect 32285 -355 32295 -320
rect 32330 -355 32340 -320
rect 32375 -355 32385 -320
rect 32420 -355 32430 -320
rect 32465 -355 32475 -320
rect 32510 -355 32520 -320
rect 32555 -355 32565 -320
rect 32600 -355 32610 -320
rect 32645 -355 32655 -320
rect 32690 -355 32700 -320
rect 32735 -355 32745 -320
rect 32780 -355 32790 -320
rect 32825 -355 32835 -320
rect 32870 -355 32890 -320
rect -120 -365 32890 -355
rect -120 -375 31305 -365
rect -120 -415 -80 -375
rect -40 -415 270 -375
rect 310 -415 620 -375
rect 660 -415 970 -375
rect 1010 -415 1320 -375
rect 1360 -415 1670 -375
rect 1710 -415 2020 -375
rect 2060 -415 2370 -375
rect 2410 -415 2720 -375
rect 2760 -415 3070 -375
rect 3110 -415 3420 -375
rect 3460 -415 3770 -375
rect 3810 -415 4120 -375
rect 4160 -415 4470 -375
rect 4510 -415 4820 -375
rect 4860 -415 5170 -375
rect 5210 -415 5520 -375
rect 5560 -415 5870 -375
rect 5910 -415 6220 -375
rect 6260 -415 6570 -375
rect 6610 -415 6920 -375
rect 6960 -415 7270 -375
rect 7310 -415 7620 -375
rect 7660 -415 7970 -375
rect 8010 -415 8320 -375
rect 8360 -415 8670 -375
rect 8710 -415 9020 -375
rect 9060 -400 31305 -375
rect 31340 -400 31350 -365
rect 31385 -400 31395 -365
rect 31430 -400 31440 -365
rect 31475 -400 31485 -365
rect 31520 -400 31530 -365
rect 31565 -400 31575 -365
rect 31610 -400 31620 -365
rect 31655 -400 31665 -365
rect 31700 -400 31710 -365
rect 31745 -400 31755 -365
rect 31790 -400 31800 -365
rect 31835 -400 31845 -365
rect 31880 -400 31890 -365
rect 31925 -400 31935 -365
rect 31970 -400 31980 -365
rect 32015 -400 32025 -365
rect 32060 -400 32070 -365
rect 32105 -400 32115 -365
rect 32150 -400 32160 -365
rect 32195 -400 32205 -365
rect 32240 -400 32250 -365
rect 32285 -400 32295 -365
rect 32330 -400 32340 -365
rect 32375 -400 32385 -365
rect 32420 -400 32430 -365
rect 32465 -400 32475 -365
rect 32510 -400 32520 -365
rect 32555 -400 32565 -365
rect 32600 -400 32610 -365
rect 32645 -400 32655 -365
rect 32690 -400 32700 -365
rect 32735 -400 32745 -365
rect 32780 -400 32790 -365
rect 32825 -400 32835 -365
rect 32870 -400 32890 -365
rect 9060 -410 32890 -400
rect 9060 -415 31305 -410
rect -120 -445 31305 -415
rect 31340 -445 31350 -410
rect 31385 -445 31395 -410
rect 31430 -445 31440 -410
rect 31475 -445 31485 -410
rect 31520 -445 31530 -410
rect 31565 -445 31575 -410
rect 31610 -445 31620 -410
rect 31655 -445 31665 -410
rect 31700 -445 31710 -410
rect 31745 -445 31755 -410
rect 31790 -445 31800 -410
rect 31835 -445 31845 -410
rect 31880 -445 31890 -410
rect 31925 -445 31935 -410
rect 31970 -445 31980 -410
rect 32015 -445 32025 -410
rect 32060 -445 32070 -410
rect 32105 -445 32115 -410
rect 32150 -445 32160 -410
rect 32195 -445 32205 -410
rect 32240 -445 32250 -410
rect 32285 -445 32295 -410
rect 32330 -445 32340 -410
rect 32375 -445 32385 -410
rect 32420 -445 32430 -410
rect 32465 -445 32475 -410
rect 32510 -445 32520 -410
rect 32555 -445 32565 -410
rect 32600 -445 32610 -410
rect 32645 -445 32655 -410
rect 32690 -445 32700 -410
rect 32735 -445 32745 -410
rect 32780 -445 32790 -410
rect 32825 -445 32835 -410
rect 32870 -445 32890 -410
rect -120 -485 -80 -445
rect -40 -485 270 -445
rect 310 -485 620 -445
rect 660 -485 970 -445
rect 1010 -485 1320 -445
rect 1360 -485 1670 -445
rect 1710 -485 2020 -445
rect 2060 -485 2370 -445
rect 2410 -485 2720 -445
rect 2760 -485 3070 -445
rect 3110 -485 3420 -445
rect 3460 -485 3770 -445
rect 3810 -485 4120 -445
rect 4160 -485 4470 -445
rect 4510 -485 4820 -445
rect 4860 -485 5170 -445
rect 5210 -485 5520 -445
rect 5560 -485 5870 -445
rect 5910 -485 6220 -445
rect 6260 -485 6570 -445
rect 6610 -485 6920 -445
rect 6960 -485 7270 -445
rect 7310 -485 7620 -445
rect 7660 -485 7970 -445
rect 8010 -485 8320 -445
rect 8360 -485 8670 -445
rect 8710 -485 9020 -445
rect 9060 -455 32890 -445
rect 9060 -485 31305 -455
rect -120 -490 31305 -485
rect 31340 -490 31350 -455
rect 31385 -490 31395 -455
rect 31430 -490 31440 -455
rect 31475 -490 31485 -455
rect 31520 -490 31530 -455
rect 31565 -490 31575 -455
rect 31610 -490 31620 -455
rect 31655 -490 31665 -455
rect 31700 -490 31710 -455
rect 31745 -490 31755 -455
rect 31790 -490 31800 -455
rect 31835 -490 31845 -455
rect 31880 -490 31890 -455
rect 31925 -490 31935 -455
rect 31970 -490 31980 -455
rect 32015 -490 32025 -455
rect 32060 -490 32070 -455
rect 32105 -490 32115 -455
rect 32150 -490 32160 -455
rect 32195 -490 32205 -455
rect 32240 -490 32250 -455
rect 32285 -490 32295 -455
rect 32330 -490 32340 -455
rect 32375 -490 32385 -455
rect 32420 -490 32430 -455
rect 32465 -490 32475 -455
rect 32510 -490 32520 -455
rect 32555 -490 32565 -455
rect 32600 -490 32610 -455
rect 32645 -490 32655 -455
rect 32690 -490 32700 -455
rect 32735 -490 32745 -455
rect 32780 -490 32790 -455
rect 32825 -490 32835 -455
rect 32870 -490 32890 -455
rect -120 -500 32890 -490
rect -120 -510 31305 -500
rect -120 -550 -80 -510
rect -40 -550 270 -510
rect 310 -550 620 -510
rect 660 -550 970 -510
rect 1010 -550 1320 -510
rect 1360 -550 1670 -510
rect 1710 -550 2020 -510
rect 2060 -550 2370 -510
rect 2410 -550 2720 -510
rect 2760 -550 3070 -510
rect 3110 -550 3420 -510
rect 3460 -550 3770 -510
rect 3810 -550 4120 -510
rect 4160 -550 4470 -510
rect 4510 -550 4820 -510
rect 4860 -550 5170 -510
rect 5210 -550 5520 -510
rect 5560 -550 5870 -510
rect 5910 -550 6220 -510
rect 6260 -550 6570 -510
rect 6610 -550 6920 -510
rect 6960 -550 7270 -510
rect 7310 -550 7620 -510
rect 7660 -550 7970 -510
rect 8010 -550 8320 -510
rect 8360 -550 8670 -510
rect 8710 -550 9020 -510
rect 9060 -535 31305 -510
rect 31340 -535 31350 -500
rect 31385 -535 31395 -500
rect 31430 -535 31440 -500
rect 31475 -535 31485 -500
rect 31520 -535 31530 -500
rect 31565 -535 31575 -500
rect 31610 -535 31620 -500
rect 31655 -535 31665 -500
rect 31700 -535 31710 -500
rect 31745 -535 31755 -500
rect 31790 -535 31800 -500
rect 31835 -535 31845 -500
rect 31880 -535 31890 -500
rect 31925 -535 31935 -500
rect 31970 -535 31980 -500
rect 32015 -535 32025 -500
rect 32060 -535 32070 -500
rect 32105 -535 32115 -500
rect 32150 -535 32160 -500
rect 32195 -535 32205 -500
rect 32240 -535 32250 -500
rect 32285 -535 32295 -500
rect 32330 -535 32340 -500
rect 32375 -535 32385 -500
rect 32420 -535 32430 -500
rect 32465 -535 32475 -500
rect 32510 -535 32520 -500
rect 32555 -535 32565 -500
rect 32600 -535 32610 -500
rect 32645 -535 32655 -500
rect 32690 -535 32700 -500
rect 32735 -535 32745 -500
rect 32780 -535 32790 -500
rect 32825 -535 32835 -500
rect 32870 -535 32890 -500
rect 9060 -545 32890 -535
rect 9060 -550 31305 -545
rect -120 -570 31305 -550
rect -120 -610 -80 -570
rect -40 -610 270 -570
rect 310 -610 620 -570
rect 660 -610 970 -570
rect 1010 -610 1320 -570
rect 1360 -610 1670 -570
rect 1710 -610 2020 -570
rect 2060 -610 2370 -570
rect 2410 -610 2720 -570
rect 2760 -610 3070 -570
rect 3110 -610 3420 -570
rect 3460 -610 3770 -570
rect 3810 -610 4120 -570
rect 4160 -610 4470 -570
rect 4510 -610 4820 -570
rect 4860 -610 5170 -570
rect 5210 -610 5520 -570
rect 5560 -610 5870 -570
rect 5910 -610 6220 -570
rect 6260 -610 6570 -570
rect 6610 -610 6920 -570
rect 6960 -610 7270 -570
rect 7310 -610 7620 -570
rect 7660 -610 7970 -570
rect 8010 -610 8320 -570
rect 8360 -610 8670 -570
rect 8710 -610 9020 -570
rect 9060 -580 31305 -570
rect 31340 -580 31350 -545
rect 31385 -580 31395 -545
rect 31430 -580 31440 -545
rect 31475 -580 31485 -545
rect 31520 -580 31530 -545
rect 31565 -580 31575 -545
rect 31610 -580 31620 -545
rect 31655 -580 31665 -545
rect 31700 -580 31710 -545
rect 31745 -580 31755 -545
rect 31790 -580 31800 -545
rect 31835 -580 31845 -545
rect 31880 -580 31890 -545
rect 31925 -580 31935 -545
rect 31970 -580 31980 -545
rect 32015 -580 32025 -545
rect 32060 -580 32070 -545
rect 32105 -580 32115 -545
rect 32150 -580 32160 -545
rect 32195 -580 32205 -545
rect 32240 -580 32250 -545
rect 32285 -580 32295 -545
rect 32330 -580 32340 -545
rect 32375 -580 32385 -545
rect 32420 -580 32430 -545
rect 32465 -580 32475 -545
rect 32510 -580 32520 -545
rect 32555 -580 32565 -545
rect 32600 -580 32610 -545
rect 32645 -580 32655 -545
rect 32690 -580 32700 -545
rect 32735 -580 32745 -545
rect 32780 -580 32790 -545
rect 32825 -580 32835 -545
rect 32870 -580 32890 -545
rect 9060 -590 32890 -580
rect 9060 -610 31305 -590
rect -120 -625 31305 -610
rect 31340 -625 31350 -590
rect 31385 -625 31395 -590
rect 31430 -625 31440 -590
rect 31475 -625 31485 -590
rect 31520 -625 31530 -590
rect 31565 -625 31575 -590
rect 31610 -625 31620 -590
rect 31655 -625 31665 -590
rect 31700 -625 31710 -590
rect 31745 -625 31755 -590
rect 31790 -625 31800 -590
rect 31835 -625 31845 -590
rect 31880 -625 31890 -590
rect 31925 -625 31935 -590
rect 31970 -625 31980 -590
rect 32015 -625 32025 -590
rect 32060 -625 32070 -590
rect 32105 -625 32115 -590
rect 32150 -625 32160 -590
rect 32195 -625 32205 -590
rect 32240 -625 32250 -590
rect 32285 -625 32295 -590
rect 32330 -625 32340 -590
rect 32375 -625 32385 -590
rect 32420 -625 32430 -590
rect 32465 -625 32475 -590
rect 32510 -625 32520 -590
rect 32555 -625 32565 -590
rect 32600 -625 32610 -590
rect 32645 -625 32655 -590
rect 32690 -625 32700 -590
rect 32735 -625 32745 -590
rect 32780 -625 32790 -590
rect 32825 -625 32835 -590
rect 32870 -625 32890 -590
rect -120 -635 32890 -625
rect -120 -675 -80 -635
rect -40 -675 270 -635
rect 310 -675 620 -635
rect 660 -675 970 -635
rect 1010 -675 1320 -635
rect 1360 -675 1670 -635
rect 1710 -675 2020 -635
rect 2060 -675 2370 -635
rect 2410 -675 2720 -635
rect 2760 -675 3070 -635
rect 3110 -675 3420 -635
rect 3460 -675 3770 -635
rect 3810 -675 4120 -635
rect 4160 -675 4470 -635
rect 4510 -675 4820 -635
rect 4860 -675 5170 -635
rect 5210 -675 5520 -635
rect 5560 -675 5870 -635
rect 5910 -675 6220 -635
rect 6260 -675 6570 -635
rect 6610 -675 6920 -635
rect 6960 -675 7270 -635
rect 7310 -675 7620 -635
rect 7660 -675 7970 -635
rect 8010 -675 8320 -635
rect 8360 -675 8670 -635
rect 8710 -675 9020 -635
rect 9060 -670 31305 -635
rect 31340 -670 31350 -635
rect 31385 -670 31395 -635
rect 31430 -670 31440 -635
rect 31475 -670 31485 -635
rect 31520 -670 31530 -635
rect 31565 -670 31575 -635
rect 31610 -670 31620 -635
rect 31655 -670 31665 -635
rect 31700 -670 31710 -635
rect 31745 -670 31755 -635
rect 31790 -670 31800 -635
rect 31835 -670 31845 -635
rect 31880 -670 31890 -635
rect 31925 -670 31935 -635
rect 31970 -670 31980 -635
rect 32015 -670 32025 -635
rect 32060 -670 32070 -635
rect 32105 -670 32115 -635
rect 32150 -670 32160 -635
rect 32195 -670 32205 -635
rect 32240 -670 32250 -635
rect 32285 -670 32295 -635
rect 32330 -670 32340 -635
rect 32375 -670 32385 -635
rect 32420 -670 32430 -635
rect 32465 -670 32475 -635
rect 32510 -670 32520 -635
rect 32555 -670 32565 -635
rect 32600 -670 32610 -635
rect 32645 -670 32655 -635
rect 32690 -670 32700 -635
rect 32735 -670 32745 -635
rect 32780 -670 32790 -635
rect 32825 -670 32835 -635
rect 32870 -670 32890 -635
rect 9060 -675 32890 -670
rect -120 -680 32890 -675
rect -120 -705 31305 -680
rect -120 -745 -80 -705
rect -40 -745 270 -705
rect 310 -745 620 -705
rect 660 -745 970 -705
rect 1010 -745 1320 -705
rect 1360 -745 1670 -705
rect 1710 -745 2020 -705
rect 2060 -745 2370 -705
rect 2410 -745 2720 -705
rect 2760 -745 3070 -705
rect 3110 -745 3420 -705
rect 3460 -745 3770 -705
rect 3810 -745 4120 -705
rect 4160 -745 4470 -705
rect 4510 -745 4820 -705
rect 4860 -745 5170 -705
rect 5210 -745 5520 -705
rect 5560 -745 5870 -705
rect 5910 -745 6220 -705
rect 6260 -745 6570 -705
rect 6610 -745 6920 -705
rect 6960 -745 7270 -705
rect 7310 -745 7620 -705
rect 7660 -745 7970 -705
rect 8010 -745 8320 -705
rect 8360 -745 8670 -705
rect 8710 -745 9020 -705
rect 9060 -715 31305 -705
rect 31340 -715 31350 -680
rect 31385 -715 31395 -680
rect 31430 -715 31440 -680
rect 31475 -715 31485 -680
rect 31520 -715 31530 -680
rect 31565 -715 31575 -680
rect 31610 -715 31620 -680
rect 31655 -715 31665 -680
rect 31700 -715 31710 -680
rect 31745 -715 31755 -680
rect 31790 -715 31800 -680
rect 31835 -715 31845 -680
rect 31880 -715 31890 -680
rect 31925 -715 31935 -680
rect 31970 -715 31980 -680
rect 32015 -715 32025 -680
rect 32060 -715 32070 -680
rect 32105 -715 32115 -680
rect 32150 -715 32160 -680
rect 32195 -715 32205 -680
rect 32240 -715 32250 -680
rect 32285 -715 32295 -680
rect 32330 -715 32340 -680
rect 32375 -715 32385 -680
rect 32420 -715 32430 -680
rect 32465 -715 32475 -680
rect 32510 -715 32520 -680
rect 32555 -715 32565 -680
rect 32600 -715 32610 -680
rect 32645 -715 32655 -680
rect 32690 -715 32700 -680
rect 32735 -715 32745 -680
rect 32780 -715 32790 -680
rect 32825 -715 32835 -680
rect 32870 -715 32890 -680
rect 9060 -725 32890 -715
rect 9060 -745 31305 -725
rect -120 -760 31305 -745
rect 31340 -760 31350 -725
rect 31385 -760 31395 -725
rect 31430 -760 31440 -725
rect 31475 -760 31485 -725
rect 31520 -760 31530 -725
rect 31565 -760 31575 -725
rect 31610 -760 31620 -725
rect 31655 -760 31665 -725
rect 31700 -760 31710 -725
rect 31745 -760 31755 -725
rect 31790 -760 31800 -725
rect 31835 -760 31845 -725
rect 31880 -760 31890 -725
rect 31925 -760 31935 -725
rect 31970 -760 31980 -725
rect 32015 -760 32025 -725
rect 32060 -760 32070 -725
rect 32105 -760 32115 -725
rect 32150 -760 32160 -725
rect 32195 -760 32205 -725
rect 32240 -760 32250 -725
rect 32285 -760 32295 -725
rect 32330 -760 32340 -725
rect 32375 -760 32385 -725
rect 32420 -760 32430 -725
rect 32465 -760 32475 -725
rect 32510 -760 32520 -725
rect 32555 -760 32565 -725
rect 32600 -760 32610 -725
rect 32645 -760 32655 -725
rect 32690 -760 32700 -725
rect 32735 -760 32745 -725
rect 32780 -760 32790 -725
rect 32825 -760 32835 -725
rect 32870 -760 32890 -725
rect -120 -770 32890 -760
rect -120 -775 31305 -770
rect -120 -815 -80 -775
rect -40 -815 270 -775
rect 310 -815 620 -775
rect 660 -815 970 -775
rect 1010 -815 1320 -775
rect 1360 -815 1670 -775
rect 1710 -815 2020 -775
rect 2060 -815 2370 -775
rect 2410 -815 2720 -775
rect 2760 -815 3070 -775
rect 3110 -815 3420 -775
rect 3460 -815 3770 -775
rect 3810 -815 4120 -775
rect 4160 -815 4470 -775
rect 4510 -815 4820 -775
rect 4860 -815 5170 -775
rect 5210 -815 5520 -775
rect 5560 -815 5870 -775
rect 5910 -815 6220 -775
rect 6260 -815 6570 -775
rect 6610 -815 6920 -775
rect 6960 -815 7270 -775
rect 7310 -815 7620 -775
rect 7660 -815 7970 -775
rect 8010 -815 8320 -775
rect 8360 -815 8670 -775
rect 8710 -815 9020 -775
rect 9060 -805 31305 -775
rect 31340 -805 31350 -770
rect 31385 -805 31395 -770
rect 31430 -805 31440 -770
rect 31475 -805 31485 -770
rect 31520 -805 31530 -770
rect 31565 -805 31575 -770
rect 31610 -805 31620 -770
rect 31655 -805 31665 -770
rect 31700 -805 31710 -770
rect 31745 -805 31755 -770
rect 31790 -805 31800 -770
rect 31835 -805 31845 -770
rect 31880 -805 31890 -770
rect 31925 -805 31935 -770
rect 31970 -805 31980 -770
rect 32015 -805 32025 -770
rect 32060 -805 32070 -770
rect 32105 -805 32115 -770
rect 32150 -805 32160 -770
rect 32195 -805 32205 -770
rect 32240 -805 32250 -770
rect 32285 -805 32295 -770
rect 32330 -805 32340 -770
rect 32375 -805 32385 -770
rect 32420 -805 32430 -770
rect 32465 -805 32475 -770
rect 32510 -805 32520 -770
rect 32555 -805 32565 -770
rect 32600 -805 32610 -770
rect 32645 -805 32655 -770
rect 32690 -805 32700 -770
rect 32735 -805 32745 -770
rect 32780 -805 32790 -770
rect 32825 -805 32835 -770
rect 32870 -805 32890 -770
rect 9060 -815 32890 -805
rect -120 -845 31305 -815
rect -120 -885 -80 -845
rect -40 -885 270 -845
rect 310 -885 620 -845
rect 660 -885 970 -845
rect 1010 -885 1320 -845
rect 1360 -885 1670 -845
rect 1710 -885 2020 -845
rect 2060 -885 2370 -845
rect 2410 -885 2720 -845
rect 2760 -885 3070 -845
rect 3110 -885 3420 -845
rect 3460 -885 3770 -845
rect 3810 -885 4120 -845
rect 4160 -885 4470 -845
rect 4510 -885 4820 -845
rect 4860 -885 5170 -845
rect 5210 -885 5520 -845
rect 5560 -885 5870 -845
rect 5910 -885 6220 -845
rect 6260 -885 6570 -845
rect 6610 -885 6920 -845
rect 6960 -885 7270 -845
rect 7310 -885 7620 -845
rect 7660 -885 7970 -845
rect 8010 -885 8320 -845
rect 8360 -885 8670 -845
rect 8710 -885 9020 -845
rect 9060 -850 31305 -845
rect 31340 -850 31350 -815
rect 31385 -850 31395 -815
rect 31430 -850 31440 -815
rect 31475 -850 31485 -815
rect 31520 -850 31530 -815
rect 31565 -850 31575 -815
rect 31610 -850 31620 -815
rect 31655 -850 31665 -815
rect 31700 -850 31710 -815
rect 31745 -850 31755 -815
rect 31790 -850 31800 -815
rect 31835 -850 31845 -815
rect 31880 -850 31890 -815
rect 31925 -850 31935 -815
rect 31970 -850 31980 -815
rect 32015 -850 32025 -815
rect 32060 -850 32070 -815
rect 32105 -850 32115 -815
rect 32150 -850 32160 -815
rect 32195 -850 32205 -815
rect 32240 -850 32250 -815
rect 32285 -850 32295 -815
rect 32330 -850 32340 -815
rect 32375 -850 32385 -815
rect 32420 -850 32430 -815
rect 32465 -850 32475 -815
rect 32510 -850 32520 -815
rect 32555 -850 32565 -815
rect 32600 -850 32610 -815
rect 32645 -850 32655 -815
rect 32690 -850 32700 -815
rect 32735 -850 32745 -815
rect 32780 -850 32790 -815
rect 32825 -850 32835 -815
rect 32870 -850 32890 -815
rect 9060 -860 32890 -850
rect 9060 -885 31305 -860
rect -120 -895 31305 -885
rect 31340 -895 31350 -860
rect 31385 -895 31395 -860
rect 31430 -895 31440 -860
rect 31475 -895 31485 -860
rect 31520 -895 31530 -860
rect 31565 -895 31575 -860
rect 31610 -895 31620 -860
rect 31655 -895 31665 -860
rect 31700 -895 31710 -860
rect 31745 -895 31755 -860
rect 31790 -895 31800 -860
rect 31835 -895 31845 -860
rect 31880 -895 31890 -860
rect 31925 -895 31935 -860
rect 31970 -895 31980 -860
rect 32015 -895 32025 -860
rect 32060 -895 32070 -860
rect 32105 -895 32115 -860
rect 32150 -895 32160 -860
rect 32195 -895 32205 -860
rect 32240 -895 32250 -860
rect 32285 -895 32295 -860
rect 32330 -895 32340 -860
rect 32375 -895 32385 -860
rect 32420 -895 32430 -860
rect 32465 -895 32475 -860
rect 32510 -895 32520 -860
rect 32555 -895 32565 -860
rect 32600 -895 32610 -860
rect 32645 -895 32655 -860
rect 32690 -895 32700 -860
rect 32735 -895 32745 -860
rect 32780 -895 32790 -860
rect 32825 -895 32835 -860
rect 32870 -895 32890 -860
rect -120 -905 32890 -895
rect -120 -910 31305 -905
rect -120 -950 -80 -910
rect -40 -950 270 -910
rect 310 -950 620 -910
rect 660 -950 970 -910
rect 1010 -950 1320 -910
rect 1360 -950 1670 -910
rect 1710 -950 2020 -910
rect 2060 -950 2370 -910
rect 2410 -950 2720 -910
rect 2760 -950 3070 -910
rect 3110 -950 3420 -910
rect 3460 -950 3770 -910
rect 3810 -950 4120 -910
rect 4160 -950 4470 -910
rect 4510 -950 4820 -910
rect 4860 -950 5170 -910
rect 5210 -950 5520 -910
rect 5560 -950 5870 -910
rect 5910 -950 6220 -910
rect 6260 -950 6570 -910
rect 6610 -950 6920 -910
rect 6960 -950 7270 -910
rect 7310 -950 7620 -910
rect 7660 -950 7970 -910
rect 8010 -950 8320 -910
rect 8360 -950 8670 -910
rect 8710 -950 9020 -910
rect 9060 -940 31305 -910
rect 31340 -940 31350 -905
rect 31385 -940 31395 -905
rect 31430 -940 31440 -905
rect 31475 -940 31485 -905
rect 31520 -940 31530 -905
rect 31565 -940 31575 -905
rect 31610 -940 31620 -905
rect 31655 -940 31665 -905
rect 31700 -940 31710 -905
rect 31745 -940 31755 -905
rect 31790 -940 31800 -905
rect 31835 -940 31845 -905
rect 31880 -940 31890 -905
rect 31925 -940 31935 -905
rect 31970 -940 31980 -905
rect 32015 -940 32025 -905
rect 32060 -940 32070 -905
rect 32105 -940 32115 -905
rect 32150 -940 32160 -905
rect 32195 -940 32205 -905
rect 32240 -940 32250 -905
rect 32285 -940 32295 -905
rect 32330 -940 32340 -905
rect 32375 -940 32385 -905
rect 32420 -940 32430 -905
rect 32465 -940 32475 -905
rect 32510 -940 32520 -905
rect 32555 -940 32565 -905
rect 32600 -940 32610 -905
rect 32645 -940 32655 -905
rect 32690 -940 32700 -905
rect 32735 -940 32745 -905
rect 32780 -940 32790 -905
rect 32825 -940 32835 -905
rect 32870 -940 32890 -905
rect 9060 -950 32890 -940
rect -120 -970 31305 -950
rect -120 -1010 -80 -970
rect -40 -1010 270 -970
rect 310 -1010 620 -970
rect 660 -1010 970 -970
rect 1010 -1010 1320 -970
rect 1360 -1010 1670 -970
rect 1710 -1010 2020 -970
rect 2060 -1010 2370 -970
rect 2410 -1010 2720 -970
rect 2760 -1010 3070 -970
rect 3110 -1010 3420 -970
rect 3460 -1010 3770 -970
rect 3810 -1010 4120 -970
rect 4160 -1010 4470 -970
rect 4510 -1010 4820 -970
rect 4860 -1010 5170 -970
rect 5210 -1010 5520 -970
rect 5560 -1010 5870 -970
rect 5910 -1010 6220 -970
rect 6260 -1010 6570 -970
rect 6610 -1010 6920 -970
rect 6960 -1010 7270 -970
rect 7310 -1010 7620 -970
rect 7660 -1010 7970 -970
rect 8010 -1010 8320 -970
rect 8360 -1010 8670 -970
rect 8710 -1010 9020 -970
rect 9060 -985 31305 -970
rect 31340 -985 31350 -950
rect 31385 -985 31395 -950
rect 31430 -985 31440 -950
rect 31475 -985 31485 -950
rect 31520 -985 31530 -950
rect 31565 -985 31575 -950
rect 31610 -985 31620 -950
rect 31655 -985 31665 -950
rect 31700 -985 31710 -950
rect 31745 -985 31755 -950
rect 31790 -985 31800 -950
rect 31835 -985 31845 -950
rect 31880 -985 31890 -950
rect 31925 -985 31935 -950
rect 31970 -985 31980 -950
rect 32015 -985 32025 -950
rect 32060 -985 32070 -950
rect 32105 -985 32115 -950
rect 32150 -985 32160 -950
rect 32195 -985 32205 -950
rect 32240 -985 32250 -950
rect 32285 -985 32295 -950
rect 32330 -985 32340 -950
rect 32375 -985 32385 -950
rect 32420 -985 32430 -950
rect 32465 -985 32475 -950
rect 32510 -985 32520 -950
rect 32555 -985 32565 -950
rect 32600 -985 32610 -950
rect 32645 -985 32655 -950
rect 32690 -985 32700 -950
rect 32735 -985 32745 -950
rect 32780 -985 32790 -950
rect 32825 -985 32835 -950
rect 32870 -985 32890 -950
rect 9060 -995 32890 -985
rect 9060 -1010 31305 -995
rect -120 -1030 31305 -1010
rect 31340 -1030 31350 -995
rect 31385 -1030 31395 -995
rect 31430 -1030 31440 -995
rect 31475 -1030 31485 -995
rect 31520 -1030 31530 -995
rect 31565 -1030 31575 -995
rect 31610 -1030 31620 -995
rect 31655 -1030 31665 -995
rect 31700 -1030 31710 -995
rect 31745 -1030 31755 -995
rect 31790 -1030 31800 -995
rect 31835 -1030 31845 -995
rect 31880 -1030 31890 -995
rect 31925 -1030 31935 -995
rect 31970 -1030 31980 -995
rect 32015 -1030 32025 -995
rect 32060 -1030 32070 -995
rect 32105 -1030 32115 -995
rect 32150 -1030 32160 -995
rect 32195 -1030 32205 -995
rect 32240 -1030 32250 -995
rect 32285 -1030 32295 -995
rect 32330 -1030 32340 -995
rect 32375 -1030 32385 -995
rect 32420 -1030 32430 -995
rect 32465 -1030 32475 -995
rect 32510 -1030 32520 -995
rect 32555 -1030 32565 -995
rect 32600 -1030 32610 -995
rect 32645 -1030 32655 -995
rect 32690 -1030 32700 -995
rect 32735 -1030 32745 -995
rect 32780 -1030 32790 -995
rect 32825 -1030 32835 -995
rect 32870 -1030 32890 -995
rect -120 -1035 32890 -1030
rect -120 -1075 -80 -1035
rect -40 -1075 270 -1035
rect 310 -1075 620 -1035
rect 660 -1075 970 -1035
rect 1010 -1075 1320 -1035
rect 1360 -1075 1670 -1035
rect 1710 -1075 2020 -1035
rect 2060 -1075 2370 -1035
rect 2410 -1075 2720 -1035
rect 2760 -1075 3070 -1035
rect 3110 -1075 3420 -1035
rect 3460 -1075 3770 -1035
rect 3810 -1075 4120 -1035
rect 4160 -1075 4470 -1035
rect 4510 -1075 4820 -1035
rect 4860 -1075 5170 -1035
rect 5210 -1075 5520 -1035
rect 5560 -1075 5870 -1035
rect 5910 -1075 6220 -1035
rect 6260 -1075 6570 -1035
rect 6610 -1075 6920 -1035
rect 6960 -1075 7270 -1035
rect 7310 -1075 7620 -1035
rect 7660 -1075 7970 -1035
rect 8010 -1075 8320 -1035
rect 8360 -1075 8670 -1035
rect 8710 -1075 9020 -1035
rect 9060 -1040 32890 -1035
rect 9060 -1075 31305 -1040
rect 31340 -1075 31350 -1040
rect 31385 -1075 31395 -1040
rect 31430 -1075 31440 -1040
rect 31475 -1075 31485 -1040
rect 31520 -1075 31530 -1040
rect 31565 -1075 31575 -1040
rect 31610 -1075 31620 -1040
rect 31655 -1075 31665 -1040
rect 31700 -1075 31710 -1040
rect 31745 -1075 31755 -1040
rect 31790 -1075 31800 -1040
rect 31835 -1075 31845 -1040
rect 31880 -1075 31890 -1040
rect 31925 -1075 31935 -1040
rect 31970 -1075 31980 -1040
rect 32015 -1075 32025 -1040
rect 32060 -1075 32070 -1040
rect 32105 -1075 32115 -1040
rect 32150 -1075 32160 -1040
rect 32195 -1075 32205 -1040
rect 32240 -1075 32250 -1040
rect 32285 -1075 32295 -1040
rect 32330 -1075 32340 -1040
rect 32375 -1075 32385 -1040
rect 32420 -1075 32430 -1040
rect 32465 -1075 32475 -1040
rect 32510 -1075 32520 -1040
rect 32555 -1075 32565 -1040
rect 32600 -1075 32610 -1040
rect 32645 -1075 32655 -1040
rect 32690 -1075 32700 -1040
rect 32735 -1075 32745 -1040
rect 32780 -1075 32790 -1040
rect 32825 -1075 32835 -1040
rect 32870 -1075 32890 -1040
rect -120 -1085 32890 -1075
rect -120 -1105 31305 -1085
rect -120 -1145 -80 -1105
rect -40 -1145 270 -1105
rect 310 -1145 620 -1105
rect 660 -1145 970 -1105
rect 1010 -1145 1320 -1105
rect 1360 -1145 1670 -1105
rect 1710 -1145 2020 -1105
rect 2060 -1145 2370 -1105
rect 2410 -1145 2720 -1105
rect 2760 -1145 3070 -1105
rect 3110 -1145 3420 -1105
rect 3460 -1145 3770 -1105
rect 3810 -1145 4120 -1105
rect 4160 -1145 4470 -1105
rect 4510 -1145 4820 -1105
rect 4860 -1145 5170 -1105
rect 5210 -1145 5520 -1105
rect 5560 -1145 5870 -1105
rect 5910 -1145 6220 -1105
rect 6260 -1145 6570 -1105
rect 6610 -1145 6920 -1105
rect 6960 -1145 7270 -1105
rect 7310 -1145 7620 -1105
rect 7660 -1145 7970 -1105
rect 8010 -1145 8320 -1105
rect 8360 -1145 8670 -1105
rect 8710 -1145 9020 -1105
rect 9060 -1120 31305 -1105
rect 31340 -1120 31350 -1085
rect 31385 -1120 31395 -1085
rect 31430 -1120 31440 -1085
rect 31475 -1120 31485 -1085
rect 31520 -1120 31530 -1085
rect 31565 -1120 31575 -1085
rect 31610 -1120 31620 -1085
rect 31655 -1120 31665 -1085
rect 31700 -1120 31710 -1085
rect 31745 -1120 31755 -1085
rect 31790 -1120 31800 -1085
rect 31835 -1120 31845 -1085
rect 31880 -1120 31890 -1085
rect 31925 -1120 31935 -1085
rect 31970 -1120 31980 -1085
rect 32015 -1120 32025 -1085
rect 32060 -1120 32070 -1085
rect 32105 -1120 32115 -1085
rect 32150 -1120 32160 -1085
rect 32195 -1120 32205 -1085
rect 32240 -1120 32250 -1085
rect 32285 -1120 32295 -1085
rect 32330 -1120 32340 -1085
rect 32375 -1120 32385 -1085
rect 32420 -1120 32430 -1085
rect 32465 -1120 32475 -1085
rect 32510 -1120 32520 -1085
rect 32555 -1120 32565 -1085
rect 32600 -1120 32610 -1085
rect 32645 -1120 32655 -1085
rect 32690 -1120 32700 -1085
rect 32735 -1120 32745 -1085
rect 32780 -1120 32790 -1085
rect 32825 -1120 32835 -1085
rect 32870 -1120 32890 -1085
rect 9060 -1130 32890 -1120
rect 9060 -1145 31305 -1130
rect -120 -1165 31305 -1145
rect 31340 -1165 31350 -1130
rect 31385 -1165 31395 -1130
rect 31430 -1165 31440 -1130
rect 31475 -1165 31485 -1130
rect 31520 -1165 31530 -1130
rect 31565 -1165 31575 -1130
rect 31610 -1165 31620 -1130
rect 31655 -1165 31665 -1130
rect 31700 -1165 31710 -1130
rect 31745 -1165 31755 -1130
rect 31790 -1165 31800 -1130
rect 31835 -1165 31845 -1130
rect 31880 -1165 31890 -1130
rect 31925 -1165 31935 -1130
rect 31970 -1165 31980 -1130
rect 32015 -1165 32025 -1130
rect 32060 -1165 32070 -1130
rect 32105 -1165 32115 -1130
rect 32150 -1165 32160 -1130
rect 32195 -1165 32205 -1130
rect 32240 -1165 32250 -1130
rect 32285 -1165 32295 -1130
rect 32330 -1165 32340 -1130
rect 32375 -1165 32385 -1130
rect 32420 -1165 32430 -1130
rect 32465 -1165 32475 -1130
rect 32510 -1165 32520 -1130
rect 32555 -1165 32565 -1130
rect 32600 -1165 32610 -1130
rect 32645 -1165 32655 -1130
rect 32690 -1165 32700 -1130
rect 32735 -1165 32745 -1130
rect 32780 -1165 32790 -1130
rect 32825 -1165 32835 -1130
rect 32870 -1165 32890 -1130
rect -120 -1175 32890 -1165
rect -120 -1215 -80 -1175
rect -40 -1215 270 -1175
rect 310 -1215 620 -1175
rect 660 -1215 970 -1175
rect 1010 -1215 1320 -1175
rect 1360 -1215 1670 -1175
rect 1710 -1215 2020 -1175
rect 2060 -1215 2370 -1175
rect 2410 -1215 2720 -1175
rect 2760 -1215 3070 -1175
rect 3110 -1215 3420 -1175
rect 3460 -1215 3770 -1175
rect 3810 -1215 4120 -1175
rect 4160 -1215 4470 -1175
rect 4510 -1215 4820 -1175
rect 4860 -1215 5170 -1175
rect 5210 -1215 5520 -1175
rect 5560 -1215 5870 -1175
rect 5910 -1215 6220 -1175
rect 6260 -1215 6570 -1175
rect 6610 -1215 6920 -1175
rect 6960 -1215 7270 -1175
rect 7310 -1215 7620 -1175
rect 7660 -1215 7970 -1175
rect 8010 -1215 8320 -1175
rect 8360 -1215 8670 -1175
rect 8710 -1215 9020 -1175
rect 9060 -1210 31305 -1175
rect 31340 -1210 31350 -1175
rect 31385 -1210 31395 -1175
rect 31430 -1210 31440 -1175
rect 31475 -1210 31485 -1175
rect 31520 -1210 31530 -1175
rect 31565 -1210 31575 -1175
rect 31610 -1210 31620 -1175
rect 31655 -1210 31665 -1175
rect 31700 -1210 31710 -1175
rect 31745 -1210 31755 -1175
rect 31790 -1210 31800 -1175
rect 31835 -1210 31845 -1175
rect 31880 -1210 31890 -1175
rect 31925 -1210 31935 -1175
rect 31970 -1210 31980 -1175
rect 32015 -1210 32025 -1175
rect 32060 -1210 32070 -1175
rect 32105 -1210 32115 -1175
rect 32150 -1210 32160 -1175
rect 32195 -1210 32205 -1175
rect 32240 -1210 32250 -1175
rect 32285 -1210 32295 -1175
rect 32330 -1210 32340 -1175
rect 32375 -1210 32385 -1175
rect 32420 -1210 32430 -1175
rect 32465 -1210 32475 -1175
rect 32510 -1210 32520 -1175
rect 32555 -1210 32565 -1175
rect 32600 -1210 32610 -1175
rect 32645 -1210 32655 -1175
rect 32690 -1210 32700 -1175
rect 32735 -1210 32745 -1175
rect 32780 -1210 32790 -1175
rect 32825 -1210 32835 -1175
rect 32870 -1210 32890 -1175
rect 9060 -1215 32890 -1210
rect -120 -1220 32890 -1215
rect -120 -1245 31305 -1220
rect -120 -1285 -80 -1245
rect -40 -1285 270 -1245
rect 310 -1285 620 -1245
rect 660 -1285 970 -1245
rect 1010 -1285 1320 -1245
rect 1360 -1285 1670 -1245
rect 1710 -1285 2020 -1245
rect 2060 -1285 2370 -1245
rect 2410 -1285 2720 -1245
rect 2760 -1285 3070 -1245
rect 3110 -1285 3420 -1245
rect 3460 -1285 3770 -1245
rect 3810 -1285 4120 -1245
rect 4160 -1285 4470 -1245
rect 4510 -1285 4820 -1245
rect 4860 -1285 5170 -1245
rect 5210 -1285 5520 -1245
rect 5560 -1285 5870 -1245
rect 5910 -1285 6220 -1245
rect 6260 -1285 6570 -1245
rect 6610 -1285 6920 -1245
rect 6960 -1285 7270 -1245
rect 7310 -1285 7620 -1245
rect 7660 -1285 7970 -1245
rect 8010 -1285 8320 -1245
rect 8360 -1285 8670 -1245
rect 8710 -1285 9020 -1245
rect 9060 -1255 31305 -1245
rect 31340 -1255 31350 -1220
rect 31385 -1255 31395 -1220
rect 31430 -1255 31440 -1220
rect 31475 -1255 31485 -1220
rect 31520 -1255 31530 -1220
rect 31565 -1255 31575 -1220
rect 31610 -1255 31620 -1220
rect 31655 -1255 31665 -1220
rect 31700 -1255 31710 -1220
rect 31745 -1255 31755 -1220
rect 31790 -1255 31800 -1220
rect 31835 -1255 31845 -1220
rect 31880 -1255 31890 -1220
rect 31925 -1255 31935 -1220
rect 31970 -1255 31980 -1220
rect 32015 -1255 32025 -1220
rect 32060 -1255 32070 -1220
rect 32105 -1255 32115 -1220
rect 32150 -1255 32160 -1220
rect 32195 -1255 32205 -1220
rect 32240 -1255 32250 -1220
rect 32285 -1255 32295 -1220
rect 32330 -1255 32340 -1220
rect 32375 -1255 32385 -1220
rect 32420 -1255 32430 -1220
rect 32465 -1255 32475 -1220
rect 32510 -1255 32520 -1220
rect 32555 -1255 32565 -1220
rect 32600 -1255 32610 -1220
rect 32645 -1255 32655 -1220
rect 32690 -1255 32700 -1220
rect 32735 -1255 32745 -1220
rect 32780 -1255 32790 -1220
rect 32825 -1255 32835 -1220
rect 32870 -1255 32890 -1220
rect 9060 -1265 32890 -1255
rect 9060 -1285 31305 -1265
rect -120 -1300 31305 -1285
rect 31340 -1300 31350 -1265
rect 31385 -1300 31395 -1265
rect 31430 -1300 31440 -1265
rect 31475 -1300 31485 -1265
rect 31520 -1300 31530 -1265
rect 31565 -1300 31575 -1265
rect 31610 -1300 31620 -1265
rect 31655 -1300 31665 -1265
rect 31700 -1300 31710 -1265
rect 31745 -1300 31755 -1265
rect 31790 -1300 31800 -1265
rect 31835 -1300 31845 -1265
rect 31880 -1300 31890 -1265
rect 31925 -1300 31935 -1265
rect 31970 -1300 31980 -1265
rect 32015 -1300 32025 -1265
rect 32060 -1300 32070 -1265
rect 32105 -1300 32115 -1265
rect 32150 -1300 32160 -1265
rect 32195 -1300 32205 -1265
rect 32240 -1300 32250 -1265
rect 32285 -1300 32295 -1265
rect 32330 -1300 32340 -1265
rect 32375 -1300 32385 -1265
rect 32420 -1300 32430 -1265
rect 32465 -1300 32475 -1265
rect 32510 -1300 32520 -1265
rect 32555 -1300 32565 -1265
rect 32600 -1300 32610 -1265
rect 32645 -1300 32655 -1265
rect 32690 -1300 32700 -1265
rect 32735 -1300 32745 -1265
rect 32780 -1300 32790 -1265
rect 32825 -1300 32835 -1265
rect 32870 -1300 32890 -1265
rect -120 -1310 32890 -1300
rect -120 -1350 -80 -1310
rect -40 -1350 270 -1310
rect 310 -1350 620 -1310
rect 660 -1350 970 -1310
rect 1010 -1350 1320 -1310
rect 1360 -1350 1670 -1310
rect 1710 -1350 2020 -1310
rect 2060 -1350 2370 -1310
rect 2410 -1350 2720 -1310
rect 2760 -1350 3070 -1310
rect 3110 -1350 3420 -1310
rect 3460 -1350 3770 -1310
rect 3810 -1350 4120 -1310
rect 4160 -1350 4470 -1310
rect 4510 -1350 4820 -1310
rect 4860 -1350 5170 -1310
rect 5210 -1350 5520 -1310
rect 5560 -1350 5870 -1310
rect 5910 -1350 6220 -1310
rect 6260 -1350 6570 -1310
rect 6610 -1350 6920 -1310
rect 6960 -1350 7270 -1310
rect 7310 -1350 7620 -1310
rect 7660 -1350 7970 -1310
rect 8010 -1350 8320 -1310
rect 8360 -1350 8670 -1310
rect 8710 -1350 9020 -1310
rect 9060 -1345 31305 -1310
rect 31340 -1345 31350 -1310
rect 31385 -1345 31395 -1310
rect 31430 -1345 31440 -1310
rect 31475 -1345 31485 -1310
rect 31520 -1345 31530 -1310
rect 31565 -1345 31575 -1310
rect 31610 -1345 31620 -1310
rect 31655 -1345 31665 -1310
rect 31700 -1345 31710 -1310
rect 31745 -1345 31755 -1310
rect 31790 -1345 31800 -1310
rect 31835 -1345 31845 -1310
rect 31880 -1345 31890 -1310
rect 31925 -1345 31935 -1310
rect 31970 -1345 31980 -1310
rect 32015 -1345 32025 -1310
rect 32060 -1345 32070 -1310
rect 32105 -1345 32115 -1310
rect 32150 -1345 32160 -1310
rect 32195 -1345 32205 -1310
rect 32240 -1345 32250 -1310
rect 32285 -1345 32295 -1310
rect 32330 -1345 32340 -1310
rect 32375 -1345 32385 -1310
rect 32420 -1345 32430 -1310
rect 32465 -1345 32475 -1310
rect 32510 -1345 32520 -1310
rect 32555 -1345 32565 -1310
rect 32600 -1345 32610 -1310
rect 32645 -1345 32655 -1310
rect 32690 -1345 32700 -1310
rect 32735 -1345 32745 -1310
rect 32780 -1345 32790 -1310
rect 32825 -1345 32835 -1310
rect 32870 -1345 32890 -1310
rect 9060 -1350 32890 -1345
rect -120 -1360 32890 -1350
use bgr_11  bgr_11_0
timestamp 1756070769
transform -1 0 22290 0 -1 11375
box 15640 -6260 19905 1640
use two_stage_opamp_dummy_magic_29  two_stage_opamp_dummy_magic_29_0
timestamp 1756064335
transform 1 0 -52410 0 1 1630
box 51710 -1500 62090 6110
<< labels >>
flabel metal3 -37570 10155 -37570 10155 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal4 35620 9150 35620 9150 3 FreeSans 800 0 320 0 GNDA
port 2 e
flabel metal2 3605 3135 3605 3135 7 FreeSans 400 0 -160 0 VIN+
port 5 w
flabel metal2 5375 3135 5375 3135 3 FreeSans 400 0 160 0 VIN-
port 6 e
flabel metal2 2185 2395 2185 2395 5 FreeSans 800 0 0 -400 VOUT+
port 3 s
flabel metal2 6795 2395 6795 2395 5 FreeSans 800 0 0 -400 VOUT-
port 4 s
<< end >>
