magic
tech sky130A
magscale 1 2
timestamp 1750177877
<< nwell >>
rect 25930 5820 30470 6490
rect 25450 4780 25870 5150
rect 26360 4490 29970 5560
rect 25270 3570 28030 4230
rect 28310 3570 31070 4230
<< pwell >>
rect 20230 4867 21570 5020
rect 20230 3833 20383 4867
rect 21417 3833 21570 4867
rect 20230 3680 21570 3833
rect 21590 4867 22930 5020
rect 21590 3833 21743 4867
rect 22777 3833 22930 4867
rect 21590 3680 22930 3833
rect 22950 4867 24290 5020
rect 22950 3833 23103 4867
rect 24137 3833 24290 4867
rect 22950 3680 24290 3833
rect 20230 3507 21570 3660
rect 20230 3050 20383 3507
rect 19910 2970 20383 3050
rect 20230 2473 20383 2970
rect 21417 2473 21570 3507
rect 20230 2320 21570 2473
rect 21590 3507 22930 3660
rect 21590 2473 21743 3507
rect 22777 2473 22930 3507
rect 21590 2320 22930 2473
rect 22950 3507 24290 3660
rect 22950 2473 23103 3507
rect 24137 2473 24290 3507
rect 26160 2950 27660 3540
rect 28680 2950 30180 3540
rect 22950 2320 24290 2473
rect 20230 2147 21570 2300
rect 20230 1113 20383 2147
rect 21417 1113 21570 2147
rect 20230 960 21570 1113
rect 21590 2147 22930 2300
rect 21590 1113 21743 2147
rect 22777 1113 22930 2147
rect 21590 960 22930 1113
rect 22950 2147 24290 2300
rect 22950 1113 23103 2147
rect 24137 1113 24290 2147
rect 25680 2000 28140 2890
rect 28200 2000 30660 2890
rect 25880 1900 30540 1910
rect 25880 1410 30530 1900
rect 25880 1400 30540 1410
rect 28609 1360 29212 1362
rect 22950 960 24290 1113
rect 25280 760 27020 1360
rect 27120 760 29220 1360
rect 29280 760 31020 1360
<< nbase >>
rect 20383 3833 21417 4867
rect 21743 3833 22777 4867
rect 23103 3833 24137 4867
rect 20383 2473 21417 3507
rect 21743 2473 22777 3507
rect 23103 2473 24137 3507
rect 20383 1113 21417 2147
rect 21743 1113 22777 2147
rect 23103 1113 24137 2147
<< nmos >>
rect 26350 3150 26390 3250
rect 26470 3150 26510 3250
rect 26590 3150 26630 3250
rect 26710 3150 26750 3250
rect 26830 3150 26870 3250
rect 26950 3150 26990 3250
rect 27070 3150 27110 3250
rect 27190 3150 27230 3250
rect 27310 3150 27350 3250
rect 27430 3150 27470 3250
rect 28870 3150 28910 3250
rect 28990 3150 29030 3250
rect 29110 3150 29150 3250
rect 29230 3150 29270 3250
rect 29350 3150 29390 3250
rect 29470 3150 29510 3250
rect 29590 3150 29630 3250
rect 29710 3150 29750 3250
rect 29830 3150 29870 3250
rect 29950 3150 29990 3250
rect 25870 2200 26870 2700
rect 26950 2200 27950 2700
rect 28390 2200 29390 2700
rect 29470 2200 30470 2700
rect 26130 1510 28130 1710
rect 28210 1510 30210 1710
rect 25470 960 25570 1160
rect 25650 960 25750 1160
rect 25830 960 25930 1160
rect 26010 960 26110 1160
rect 26190 960 26290 1160
rect 26370 960 26470 1160
rect 26550 960 26650 1160
rect 26730 960 26830 1160
rect 27310 960 27410 1160
rect 27490 960 27590 1160
rect 27670 960 27770 1160
rect 27850 960 27950 1160
rect 28030 960 28130 1160
rect 28210 960 28310 1160
rect 28390 960 28490 1160
rect 28570 960 28670 1160
rect 28750 960 28850 1160
rect 28930 960 29030 1160
rect 29470 960 29570 1160
rect 29650 960 29750 1160
rect 29830 960 29930 1160
rect 30010 960 30110 1160
rect 30190 960 30290 1160
rect 30370 960 30470 1160
rect 30550 960 30650 1160
rect 30730 960 30830 1160
<< pmos >>
rect 26230 6050 26330 6250
rect 26410 6050 26510 6250
rect 26590 6050 26690 6250
rect 26770 6050 26870 6250
rect 26950 6050 27050 6250
rect 27130 6050 27230 6250
rect 27310 6050 27410 6250
rect 27490 6050 27590 6250
rect 27670 6050 27770 6250
rect 27850 6050 27950 6250
rect 28030 6050 28130 6250
rect 28210 6050 28310 6250
rect 28390 6050 28490 6250
rect 28570 6050 28670 6250
rect 28750 6050 28850 6250
rect 28930 6050 29030 6250
rect 29110 6050 29210 6250
rect 29290 6050 29390 6250
rect 29470 6050 29570 6250
rect 29650 6050 29750 6250
rect 29830 6050 29930 6250
rect 30010 6050 30110 6250
rect 25590 4900 25620 5100
rect 25700 4900 25730 5100
rect 26590 4730 26690 5330
rect 26770 4730 26870 5330
rect 26950 4730 27050 5330
rect 27130 4730 27230 5330
rect 27310 4730 27410 5330
rect 27490 4730 27590 5330
rect 27670 4730 27770 5330
rect 27850 4730 27950 5330
rect 28030 4730 28130 5330
rect 28210 4730 28310 5330
rect 28390 4730 28490 5330
rect 28570 4730 28670 5330
rect 28750 4730 28850 5330
rect 28930 4730 29030 5330
rect 29110 4730 29210 5330
rect 29290 4730 29390 5330
rect 29470 4730 29570 5330
rect 29650 4730 29750 5330
rect 25490 3800 25530 4000
rect 25610 3800 25650 4000
rect 25730 3800 25770 4000
rect 25850 3800 25890 4000
rect 25970 3800 26010 4000
rect 26090 3800 26130 4000
rect 26210 3800 26250 4000
rect 26330 3800 26370 4000
rect 26450 3800 26490 4000
rect 26570 3800 26610 4000
rect 26690 3800 26730 4000
rect 26810 3800 26850 4000
rect 26930 3800 26970 4000
rect 27050 3800 27090 4000
rect 27170 3800 27210 4000
rect 27290 3800 27330 4000
rect 27410 3800 27450 4000
rect 27530 3800 27570 4000
rect 27650 3800 27690 4000
rect 27770 3800 27810 4000
rect 28530 3800 28570 4000
rect 28650 3800 28690 4000
rect 28770 3800 28810 4000
rect 28890 3800 28930 4000
rect 29010 3800 29050 4000
rect 29130 3800 29170 4000
rect 29250 3800 29290 4000
rect 29370 3800 29410 4000
rect 29490 3800 29530 4000
rect 29610 3800 29650 4000
rect 29730 3800 29770 4000
rect 29850 3800 29890 4000
rect 29970 3800 30010 4000
rect 30090 3800 30130 4000
rect 30210 3800 30250 4000
rect 30330 3800 30370 4000
rect 30450 3800 30490 4000
rect 30570 3800 30610 4000
rect 30690 3800 30730 4000
rect 30810 3800 30850 4000
<< ndiff >>
rect 26270 3220 26350 3250
rect 26270 3180 26290 3220
rect 26330 3180 26350 3220
rect 26270 3150 26350 3180
rect 26390 3220 26470 3250
rect 26390 3180 26410 3220
rect 26450 3180 26470 3220
rect 26390 3150 26470 3180
rect 26510 3220 26590 3250
rect 26510 3180 26530 3220
rect 26570 3180 26590 3220
rect 26510 3150 26590 3180
rect 26630 3220 26710 3250
rect 26630 3180 26650 3220
rect 26690 3180 26710 3220
rect 26630 3150 26710 3180
rect 26750 3220 26830 3250
rect 26750 3180 26770 3220
rect 26810 3180 26830 3220
rect 26750 3150 26830 3180
rect 26870 3220 26950 3250
rect 26870 3180 26890 3220
rect 26930 3180 26950 3220
rect 26870 3150 26950 3180
rect 26990 3220 27070 3250
rect 26990 3180 27010 3220
rect 27050 3180 27070 3220
rect 26990 3150 27070 3180
rect 27110 3220 27190 3250
rect 27110 3180 27130 3220
rect 27170 3180 27190 3220
rect 27110 3150 27190 3180
rect 27230 3220 27310 3250
rect 27230 3180 27250 3220
rect 27290 3180 27310 3220
rect 27230 3150 27310 3180
rect 27350 3220 27430 3250
rect 27350 3180 27370 3220
rect 27410 3180 27430 3220
rect 27350 3150 27430 3180
rect 27470 3220 27550 3250
rect 27470 3180 27490 3220
rect 27530 3180 27550 3220
rect 27470 3150 27550 3180
rect 28790 3220 28870 3250
rect 28790 3180 28810 3220
rect 28850 3180 28870 3220
rect 28790 3150 28870 3180
rect 28910 3220 28990 3250
rect 28910 3180 28930 3220
rect 28970 3180 28990 3220
rect 28910 3150 28990 3180
rect 29030 3220 29110 3250
rect 29030 3180 29050 3220
rect 29090 3180 29110 3220
rect 29030 3150 29110 3180
rect 29150 3220 29230 3250
rect 29150 3180 29170 3220
rect 29210 3180 29230 3220
rect 29150 3150 29230 3180
rect 29270 3220 29350 3250
rect 29270 3180 29290 3220
rect 29330 3180 29350 3220
rect 29270 3150 29350 3180
rect 29390 3220 29470 3250
rect 29390 3180 29410 3220
rect 29450 3180 29470 3220
rect 29390 3150 29470 3180
rect 29510 3220 29590 3250
rect 29510 3180 29530 3220
rect 29570 3180 29590 3220
rect 29510 3150 29590 3180
rect 29630 3220 29710 3250
rect 29630 3180 29650 3220
rect 29690 3180 29710 3220
rect 29630 3150 29710 3180
rect 29750 3220 29830 3250
rect 29750 3180 29770 3220
rect 29810 3180 29830 3220
rect 29750 3150 29830 3180
rect 29870 3220 29950 3250
rect 29870 3180 29890 3220
rect 29930 3180 29950 3220
rect 29870 3150 29950 3180
rect 29990 3220 30070 3250
rect 29990 3180 30010 3220
rect 30050 3180 30070 3220
rect 29990 3150 30070 3180
rect 25790 2670 25870 2700
rect 25790 2630 25810 2670
rect 25850 2630 25870 2670
rect 25790 2570 25870 2630
rect 25790 2530 25810 2570
rect 25850 2530 25870 2570
rect 25790 2470 25870 2530
rect 25790 2430 25810 2470
rect 25850 2430 25870 2470
rect 25790 2370 25870 2430
rect 25790 2330 25810 2370
rect 25850 2330 25870 2370
rect 25790 2270 25870 2330
rect 25790 2230 25810 2270
rect 25850 2230 25870 2270
rect 25790 2200 25870 2230
rect 26870 2670 26950 2700
rect 26870 2630 26890 2670
rect 26930 2630 26950 2670
rect 26870 2570 26950 2630
rect 26870 2530 26890 2570
rect 26930 2530 26950 2570
rect 26870 2470 26950 2530
rect 26870 2430 26890 2470
rect 26930 2430 26950 2470
rect 26870 2370 26950 2430
rect 26870 2330 26890 2370
rect 26930 2330 26950 2370
rect 26870 2270 26950 2330
rect 26870 2230 26890 2270
rect 26930 2230 26950 2270
rect 26870 2200 26950 2230
rect 27950 2670 28030 2700
rect 27950 2630 27970 2670
rect 28010 2630 28030 2670
rect 27950 2570 28030 2630
rect 27950 2530 27970 2570
rect 28010 2530 28030 2570
rect 27950 2470 28030 2530
rect 27950 2430 27970 2470
rect 28010 2430 28030 2470
rect 27950 2370 28030 2430
rect 27950 2330 27970 2370
rect 28010 2330 28030 2370
rect 27950 2270 28030 2330
rect 27950 2230 27970 2270
rect 28010 2230 28030 2270
rect 27950 2200 28030 2230
rect 28310 2670 28390 2700
rect 28310 2630 28330 2670
rect 28370 2630 28390 2670
rect 28310 2570 28390 2630
rect 28310 2530 28330 2570
rect 28370 2530 28390 2570
rect 28310 2470 28390 2530
rect 28310 2430 28330 2470
rect 28370 2430 28390 2470
rect 28310 2370 28390 2430
rect 28310 2330 28330 2370
rect 28370 2330 28390 2370
rect 28310 2270 28390 2330
rect 28310 2230 28330 2270
rect 28370 2230 28390 2270
rect 28310 2200 28390 2230
rect 29390 2670 29470 2700
rect 29390 2630 29410 2670
rect 29450 2630 29470 2670
rect 29390 2570 29470 2630
rect 29390 2530 29410 2570
rect 29450 2530 29470 2570
rect 29390 2470 29470 2530
rect 29390 2430 29410 2470
rect 29450 2430 29470 2470
rect 29390 2370 29470 2430
rect 29390 2330 29410 2370
rect 29450 2330 29470 2370
rect 29390 2270 29470 2330
rect 29390 2230 29410 2270
rect 29450 2230 29470 2270
rect 29390 2200 29470 2230
rect 30470 2670 30550 2700
rect 30470 2630 30490 2670
rect 30530 2630 30550 2670
rect 30470 2570 30550 2630
rect 30470 2530 30490 2570
rect 30530 2530 30550 2570
rect 30470 2470 30550 2530
rect 30470 2430 30490 2470
rect 30530 2430 30550 2470
rect 30470 2370 30550 2430
rect 30470 2330 30490 2370
rect 30530 2330 30550 2370
rect 30470 2270 30550 2330
rect 30470 2230 30490 2270
rect 30530 2230 30550 2270
rect 30470 2200 30550 2230
rect 26050 1680 26130 1710
rect 26050 1640 26070 1680
rect 26110 1640 26130 1680
rect 26050 1580 26130 1640
rect 26050 1540 26070 1580
rect 26110 1540 26130 1580
rect 26050 1510 26130 1540
rect 28130 1680 28210 1710
rect 28130 1640 28150 1680
rect 28190 1640 28210 1680
rect 28130 1580 28210 1640
rect 28130 1540 28150 1580
rect 28190 1540 28210 1580
rect 28130 1510 28210 1540
rect 30210 1680 30290 1710
rect 30210 1640 30230 1680
rect 30270 1640 30290 1680
rect 30210 1580 30290 1640
rect 30210 1540 30230 1580
rect 30270 1540 30290 1580
rect 30210 1510 30290 1540
rect 25390 1130 25470 1160
rect 25390 1090 25410 1130
rect 25450 1090 25470 1130
rect 25390 1030 25470 1090
rect 25390 990 25410 1030
rect 25450 990 25470 1030
rect 25390 960 25470 990
rect 25570 1130 25650 1160
rect 25570 1090 25590 1130
rect 25630 1090 25650 1130
rect 25570 1030 25650 1090
rect 25570 990 25590 1030
rect 25630 990 25650 1030
rect 25570 960 25650 990
rect 25750 1130 25830 1160
rect 25750 1090 25770 1130
rect 25810 1090 25830 1130
rect 25750 1030 25830 1090
rect 25750 990 25770 1030
rect 25810 990 25830 1030
rect 25750 960 25830 990
rect 25930 1130 26010 1160
rect 25930 1090 25950 1130
rect 25990 1090 26010 1130
rect 25930 1030 26010 1090
rect 25930 990 25950 1030
rect 25990 990 26010 1030
rect 25930 960 26010 990
rect 26110 1130 26190 1160
rect 26110 1090 26130 1130
rect 26170 1090 26190 1130
rect 26110 1030 26190 1090
rect 26110 990 26130 1030
rect 26170 990 26190 1030
rect 26110 960 26190 990
rect 26290 1130 26370 1160
rect 26290 1090 26310 1130
rect 26350 1090 26370 1130
rect 26290 1030 26370 1090
rect 26290 990 26310 1030
rect 26350 990 26370 1030
rect 26290 960 26370 990
rect 26470 1130 26550 1160
rect 26470 1090 26490 1130
rect 26530 1090 26550 1130
rect 26470 1030 26550 1090
rect 26470 990 26490 1030
rect 26530 990 26550 1030
rect 26470 960 26550 990
rect 26650 1130 26730 1160
rect 26650 1090 26670 1130
rect 26710 1090 26730 1130
rect 26650 1030 26730 1090
rect 26650 990 26670 1030
rect 26710 990 26730 1030
rect 26650 960 26730 990
rect 26830 1130 26910 1160
rect 26830 1090 26850 1130
rect 26890 1090 26910 1130
rect 26830 1030 26910 1090
rect 26830 990 26850 1030
rect 26890 990 26910 1030
rect 26830 960 26910 990
rect 27230 1130 27310 1160
rect 27230 1090 27250 1130
rect 27290 1090 27310 1130
rect 27230 1030 27310 1090
rect 27230 990 27250 1030
rect 27290 990 27310 1030
rect 27230 960 27310 990
rect 27410 1130 27490 1160
rect 27410 1090 27430 1130
rect 27470 1090 27490 1130
rect 27410 1030 27490 1090
rect 27410 990 27430 1030
rect 27470 990 27490 1030
rect 27410 960 27490 990
rect 27590 1130 27670 1160
rect 27590 1090 27610 1130
rect 27650 1090 27670 1130
rect 27590 1030 27670 1090
rect 27590 990 27610 1030
rect 27650 990 27670 1030
rect 27590 960 27670 990
rect 27770 1130 27850 1160
rect 27770 1090 27790 1130
rect 27830 1090 27850 1130
rect 27770 1030 27850 1090
rect 27770 990 27790 1030
rect 27830 990 27850 1030
rect 27770 960 27850 990
rect 27950 1130 28030 1160
rect 27950 1090 27970 1130
rect 28010 1090 28030 1130
rect 27950 1030 28030 1090
rect 27950 990 27970 1030
rect 28010 990 28030 1030
rect 27950 960 28030 990
rect 28130 1130 28210 1160
rect 28130 1090 28150 1130
rect 28190 1090 28210 1130
rect 28130 1030 28210 1090
rect 28130 990 28150 1030
rect 28190 990 28210 1030
rect 28130 960 28210 990
rect 28310 1130 28390 1160
rect 28310 1090 28330 1130
rect 28370 1090 28390 1130
rect 28310 1030 28390 1090
rect 28310 990 28330 1030
rect 28370 990 28390 1030
rect 28310 960 28390 990
rect 28490 1130 28570 1160
rect 28490 1090 28510 1130
rect 28550 1090 28570 1130
rect 28490 1030 28570 1090
rect 28490 990 28510 1030
rect 28550 990 28570 1030
rect 28490 960 28570 990
rect 28670 1130 28750 1160
rect 28670 1090 28690 1130
rect 28730 1090 28750 1130
rect 28670 1030 28750 1090
rect 28670 990 28690 1030
rect 28730 990 28750 1030
rect 28670 960 28750 990
rect 28850 1130 28930 1160
rect 28850 1090 28870 1130
rect 28910 1090 28930 1130
rect 28850 1030 28930 1090
rect 28850 990 28870 1030
rect 28910 990 28930 1030
rect 28850 960 28930 990
rect 29030 1130 29110 1160
rect 29030 1090 29050 1130
rect 29090 1090 29110 1130
rect 29030 1030 29110 1090
rect 29030 990 29050 1030
rect 29090 990 29110 1030
rect 29030 960 29110 990
rect 29390 1130 29470 1160
rect 29390 1090 29410 1130
rect 29450 1090 29470 1130
rect 29390 1030 29470 1090
rect 29390 990 29410 1030
rect 29450 990 29470 1030
rect 29390 960 29470 990
rect 29570 1130 29650 1160
rect 29570 1090 29590 1130
rect 29630 1090 29650 1130
rect 29570 1030 29650 1090
rect 29570 990 29590 1030
rect 29630 990 29650 1030
rect 29570 960 29650 990
rect 29750 1130 29830 1160
rect 29750 1090 29770 1130
rect 29810 1090 29830 1130
rect 29750 1030 29830 1090
rect 29750 990 29770 1030
rect 29810 990 29830 1030
rect 29750 960 29830 990
rect 29930 1130 30010 1160
rect 29930 1090 29950 1130
rect 29990 1090 30010 1130
rect 29930 1030 30010 1090
rect 29930 990 29950 1030
rect 29990 990 30010 1030
rect 29930 960 30010 990
rect 30110 1130 30190 1160
rect 30110 1090 30130 1130
rect 30170 1090 30190 1130
rect 30110 1030 30190 1090
rect 30110 990 30130 1030
rect 30170 990 30190 1030
rect 30110 960 30190 990
rect 30290 1130 30370 1160
rect 30290 1090 30310 1130
rect 30350 1090 30370 1130
rect 30290 1030 30370 1090
rect 30290 990 30310 1030
rect 30350 990 30370 1030
rect 30290 960 30370 990
rect 30470 1130 30550 1160
rect 30470 1090 30490 1130
rect 30530 1090 30550 1130
rect 30470 1030 30550 1090
rect 30470 990 30490 1030
rect 30530 990 30550 1030
rect 30470 960 30550 990
rect 30650 1130 30730 1160
rect 30650 1090 30670 1130
rect 30710 1090 30730 1130
rect 30650 1030 30730 1090
rect 30650 990 30670 1030
rect 30710 990 30730 1030
rect 30650 960 30730 990
rect 30830 1130 30910 1160
rect 30830 1090 30850 1130
rect 30890 1090 30910 1130
rect 30830 1030 30910 1090
rect 30830 990 30850 1030
rect 30890 990 30910 1030
rect 30830 960 30910 990
<< pdiff >>
rect 26150 6220 26230 6250
rect 26150 6180 26170 6220
rect 26210 6180 26230 6220
rect 26150 6120 26230 6180
rect 26150 6080 26170 6120
rect 26210 6080 26230 6120
rect 26150 6050 26230 6080
rect 26330 6220 26410 6250
rect 26330 6180 26350 6220
rect 26390 6180 26410 6220
rect 26330 6120 26410 6180
rect 26330 6080 26350 6120
rect 26390 6080 26410 6120
rect 26330 6050 26410 6080
rect 26510 6220 26590 6250
rect 26510 6180 26530 6220
rect 26570 6180 26590 6220
rect 26510 6120 26590 6180
rect 26510 6080 26530 6120
rect 26570 6080 26590 6120
rect 26510 6050 26590 6080
rect 26690 6220 26770 6250
rect 26690 6180 26710 6220
rect 26750 6180 26770 6220
rect 26690 6120 26770 6180
rect 26690 6080 26710 6120
rect 26750 6080 26770 6120
rect 26690 6050 26770 6080
rect 26870 6220 26950 6250
rect 26870 6180 26890 6220
rect 26930 6180 26950 6220
rect 26870 6120 26950 6180
rect 26870 6080 26890 6120
rect 26930 6080 26950 6120
rect 26870 6050 26950 6080
rect 27050 6220 27130 6250
rect 27050 6180 27070 6220
rect 27110 6180 27130 6220
rect 27050 6120 27130 6180
rect 27050 6080 27070 6120
rect 27110 6080 27130 6120
rect 27050 6050 27130 6080
rect 27230 6220 27310 6250
rect 27230 6180 27250 6220
rect 27290 6180 27310 6220
rect 27230 6120 27310 6180
rect 27230 6080 27250 6120
rect 27290 6080 27310 6120
rect 27230 6050 27310 6080
rect 27410 6220 27490 6250
rect 27410 6180 27430 6220
rect 27470 6180 27490 6220
rect 27410 6120 27490 6180
rect 27410 6080 27430 6120
rect 27470 6080 27490 6120
rect 27410 6050 27490 6080
rect 27590 6220 27670 6250
rect 27590 6180 27610 6220
rect 27650 6180 27670 6220
rect 27590 6120 27670 6180
rect 27590 6080 27610 6120
rect 27650 6080 27670 6120
rect 27590 6050 27670 6080
rect 27770 6220 27850 6250
rect 27770 6180 27790 6220
rect 27830 6180 27850 6220
rect 27770 6120 27850 6180
rect 27770 6080 27790 6120
rect 27830 6080 27850 6120
rect 27770 6050 27850 6080
rect 27950 6220 28030 6250
rect 27950 6180 27970 6220
rect 28010 6180 28030 6220
rect 27950 6120 28030 6180
rect 27950 6080 27970 6120
rect 28010 6080 28030 6120
rect 27950 6050 28030 6080
rect 28130 6220 28210 6250
rect 28130 6180 28150 6220
rect 28190 6180 28210 6220
rect 28130 6120 28210 6180
rect 28130 6080 28150 6120
rect 28190 6080 28210 6120
rect 28130 6050 28210 6080
rect 28310 6220 28390 6250
rect 28310 6180 28330 6220
rect 28370 6180 28390 6220
rect 28310 6120 28390 6180
rect 28310 6080 28330 6120
rect 28370 6080 28390 6120
rect 28310 6050 28390 6080
rect 28490 6220 28570 6250
rect 28490 6180 28510 6220
rect 28550 6180 28570 6220
rect 28490 6120 28570 6180
rect 28490 6080 28510 6120
rect 28550 6080 28570 6120
rect 28490 6050 28570 6080
rect 28670 6220 28750 6250
rect 28670 6180 28690 6220
rect 28730 6180 28750 6220
rect 28670 6120 28750 6180
rect 28670 6080 28690 6120
rect 28730 6080 28750 6120
rect 28670 6050 28750 6080
rect 28850 6220 28930 6250
rect 28850 6180 28870 6220
rect 28910 6180 28930 6220
rect 28850 6120 28930 6180
rect 28850 6080 28870 6120
rect 28910 6080 28930 6120
rect 28850 6050 28930 6080
rect 29030 6220 29110 6250
rect 29030 6180 29050 6220
rect 29090 6180 29110 6220
rect 29030 6120 29110 6180
rect 29030 6080 29050 6120
rect 29090 6080 29110 6120
rect 29030 6050 29110 6080
rect 29210 6220 29290 6250
rect 29210 6180 29230 6220
rect 29270 6180 29290 6220
rect 29210 6120 29290 6180
rect 29210 6080 29230 6120
rect 29270 6080 29290 6120
rect 29210 6050 29290 6080
rect 29390 6220 29470 6250
rect 29390 6180 29410 6220
rect 29450 6180 29470 6220
rect 29390 6120 29470 6180
rect 29390 6080 29410 6120
rect 29450 6080 29470 6120
rect 29390 6050 29470 6080
rect 29570 6220 29650 6250
rect 29570 6180 29590 6220
rect 29630 6180 29650 6220
rect 29570 6120 29650 6180
rect 29570 6080 29590 6120
rect 29630 6080 29650 6120
rect 29570 6050 29650 6080
rect 29750 6220 29830 6250
rect 29750 6180 29770 6220
rect 29810 6180 29830 6220
rect 29750 6120 29830 6180
rect 29750 6080 29770 6120
rect 29810 6080 29830 6120
rect 29750 6050 29830 6080
rect 29930 6220 30010 6250
rect 29930 6180 29950 6220
rect 29990 6180 30010 6220
rect 29930 6120 30010 6180
rect 29930 6080 29950 6120
rect 29990 6080 30010 6120
rect 29930 6050 30010 6080
rect 30110 6220 30190 6250
rect 30110 6180 30130 6220
rect 30170 6180 30190 6220
rect 30110 6120 30190 6180
rect 30110 6080 30130 6120
rect 30170 6080 30190 6120
rect 30110 6050 30190 6080
rect 25510 5070 25590 5100
rect 25510 5030 25530 5070
rect 25570 5030 25590 5070
rect 20560 4638 21240 4690
rect 20560 4604 20614 4638
rect 20648 4604 20704 4638
rect 20738 4604 20794 4638
rect 20828 4604 20884 4638
rect 20918 4604 20974 4638
rect 21008 4604 21064 4638
rect 21098 4604 21154 4638
rect 21188 4604 21240 4638
rect 20560 4548 21240 4604
rect 20560 4514 20614 4548
rect 20648 4514 20704 4548
rect 20738 4514 20794 4548
rect 20828 4514 20884 4548
rect 20918 4514 20974 4548
rect 21008 4514 21064 4548
rect 21098 4514 21154 4548
rect 21188 4514 21240 4548
rect 20560 4458 21240 4514
rect 20560 4424 20614 4458
rect 20648 4424 20704 4458
rect 20738 4424 20794 4458
rect 20828 4424 20884 4458
rect 20918 4424 20974 4458
rect 21008 4424 21064 4458
rect 21098 4424 21154 4458
rect 21188 4424 21240 4458
rect 20560 4368 21240 4424
rect 20560 4334 20614 4368
rect 20648 4334 20704 4368
rect 20738 4334 20794 4368
rect 20828 4334 20884 4368
rect 20918 4334 20974 4368
rect 21008 4334 21064 4368
rect 21098 4334 21154 4368
rect 21188 4334 21240 4368
rect 20560 4278 21240 4334
rect 20560 4244 20614 4278
rect 20648 4244 20704 4278
rect 20738 4244 20794 4278
rect 20828 4244 20884 4278
rect 20918 4244 20974 4278
rect 21008 4244 21064 4278
rect 21098 4244 21154 4278
rect 21188 4244 21240 4278
rect 20560 4188 21240 4244
rect 20560 4154 20614 4188
rect 20648 4154 20704 4188
rect 20738 4154 20794 4188
rect 20828 4154 20884 4188
rect 20918 4154 20974 4188
rect 21008 4154 21064 4188
rect 21098 4154 21154 4188
rect 21188 4154 21240 4188
rect 20560 4098 21240 4154
rect 20560 4064 20614 4098
rect 20648 4064 20704 4098
rect 20738 4064 20794 4098
rect 20828 4064 20884 4098
rect 20918 4064 20974 4098
rect 21008 4064 21064 4098
rect 21098 4064 21154 4098
rect 21188 4064 21240 4098
rect 20560 4010 21240 4064
rect 21920 4638 22600 4690
rect 21920 4604 21974 4638
rect 22008 4604 22064 4638
rect 22098 4604 22154 4638
rect 22188 4604 22244 4638
rect 22278 4604 22334 4638
rect 22368 4604 22424 4638
rect 22458 4604 22514 4638
rect 22548 4604 22600 4638
rect 21920 4548 22600 4604
rect 21920 4514 21974 4548
rect 22008 4514 22064 4548
rect 22098 4514 22154 4548
rect 22188 4514 22244 4548
rect 22278 4514 22334 4548
rect 22368 4514 22424 4548
rect 22458 4514 22514 4548
rect 22548 4514 22600 4548
rect 21920 4458 22600 4514
rect 21920 4424 21974 4458
rect 22008 4424 22064 4458
rect 22098 4424 22154 4458
rect 22188 4424 22244 4458
rect 22278 4424 22334 4458
rect 22368 4424 22424 4458
rect 22458 4424 22514 4458
rect 22548 4424 22600 4458
rect 21920 4368 22600 4424
rect 21920 4334 21974 4368
rect 22008 4334 22064 4368
rect 22098 4334 22154 4368
rect 22188 4334 22244 4368
rect 22278 4334 22334 4368
rect 22368 4334 22424 4368
rect 22458 4334 22514 4368
rect 22548 4334 22600 4368
rect 21920 4278 22600 4334
rect 21920 4244 21974 4278
rect 22008 4244 22064 4278
rect 22098 4244 22154 4278
rect 22188 4244 22244 4278
rect 22278 4244 22334 4278
rect 22368 4244 22424 4278
rect 22458 4244 22514 4278
rect 22548 4244 22600 4278
rect 21920 4188 22600 4244
rect 21920 4154 21974 4188
rect 22008 4154 22064 4188
rect 22098 4154 22154 4188
rect 22188 4154 22244 4188
rect 22278 4154 22334 4188
rect 22368 4154 22424 4188
rect 22458 4154 22514 4188
rect 22548 4154 22600 4188
rect 21920 4098 22600 4154
rect 21920 4064 21974 4098
rect 22008 4064 22064 4098
rect 22098 4064 22154 4098
rect 22188 4064 22244 4098
rect 22278 4064 22334 4098
rect 22368 4064 22424 4098
rect 22458 4064 22514 4098
rect 22548 4064 22600 4098
rect 21920 4010 22600 4064
rect 25510 4970 25590 5030
rect 25510 4930 25530 4970
rect 25570 4930 25590 4970
rect 25510 4900 25590 4930
rect 25620 5070 25700 5100
rect 25620 5030 25640 5070
rect 25680 5030 25700 5070
rect 25620 4970 25700 5030
rect 25620 4930 25640 4970
rect 25680 4930 25700 4970
rect 25620 4900 25700 4930
rect 25730 5070 25810 5100
rect 25730 5030 25750 5070
rect 25790 5030 25810 5070
rect 25730 4970 25810 5030
rect 25730 4930 25750 4970
rect 25790 4930 25810 4970
rect 25730 4900 25810 4930
rect 23280 4638 23960 4690
rect 23280 4604 23334 4638
rect 23368 4604 23424 4638
rect 23458 4604 23514 4638
rect 23548 4604 23604 4638
rect 23638 4604 23694 4638
rect 23728 4604 23784 4638
rect 23818 4604 23874 4638
rect 23908 4604 23960 4638
rect 23280 4548 23960 4604
rect 23280 4514 23334 4548
rect 23368 4514 23424 4548
rect 23458 4514 23514 4548
rect 23548 4514 23604 4548
rect 23638 4514 23694 4548
rect 23728 4514 23784 4548
rect 23818 4514 23874 4548
rect 23908 4514 23960 4548
rect 23280 4458 23960 4514
rect 23280 4424 23334 4458
rect 23368 4424 23424 4458
rect 23458 4424 23514 4458
rect 23548 4424 23604 4458
rect 23638 4424 23694 4458
rect 23728 4424 23784 4458
rect 23818 4424 23874 4458
rect 23908 4424 23960 4458
rect 23280 4368 23960 4424
rect 23280 4334 23334 4368
rect 23368 4334 23424 4368
rect 23458 4334 23514 4368
rect 23548 4334 23604 4368
rect 23638 4334 23694 4368
rect 23728 4334 23784 4368
rect 23818 4334 23874 4368
rect 23908 4334 23960 4368
rect 23280 4278 23960 4334
rect 23280 4244 23334 4278
rect 23368 4244 23424 4278
rect 23458 4244 23514 4278
rect 23548 4244 23604 4278
rect 23638 4244 23694 4278
rect 23728 4244 23784 4278
rect 23818 4244 23874 4278
rect 23908 4244 23960 4278
rect 23280 4188 23960 4244
rect 23280 4154 23334 4188
rect 23368 4154 23424 4188
rect 23458 4154 23514 4188
rect 23548 4154 23604 4188
rect 23638 4154 23694 4188
rect 23728 4154 23784 4188
rect 23818 4154 23874 4188
rect 23908 4154 23960 4188
rect 23280 4098 23960 4154
rect 23280 4064 23334 4098
rect 23368 4064 23424 4098
rect 23458 4064 23514 4098
rect 23548 4064 23604 4098
rect 23638 4064 23694 4098
rect 23728 4064 23784 4098
rect 23818 4064 23874 4098
rect 23908 4064 23960 4098
rect 23280 4010 23960 4064
rect 26500 5300 26590 5330
rect 26500 5260 26530 5300
rect 26570 5260 26590 5300
rect 26500 5200 26590 5260
rect 26500 5160 26530 5200
rect 26570 5160 26590 5200
rect 26500 5100 26590 5160
rect 26500 5060 26530 5100
rect 26570 5060 26590 5100
rect 26500 5000 26590 5060
rect 26500 4960 26530 5000
rect 26570 4960 26590 5000
rect 26500 4900 26590 4960
rect 26500 4860 26530 4900
rect 26570 4860 26590 4900
rect 26500 4800 26590 4860
rect 26500 4760 26530 4800
rect 26570 4760 26590 4800
rect 26500 4730 26590 4760
rect 26690 5300 26770 5330
rect 26690 5260 26710 5300
rect 26750 5260 26770 5300
rect 26690 5200 26770 5260
rect 26690 5160 26710 5200
rect 26750 5160 26770 5200
rect 26690 5100 26770 5160
rect 26690 5060 26710 5100
rect 26750 5060 26770 5100
rect 26690 5000 26770 5060
rect 26690 4960 26710 5000
rect 26750 4960 26770 5000
rect 26690 4900 26770 4960
rect 26690 4860 26710 4900
rect 26750 4860 26770 4900
rect 26690 4800 26770 4860
rect 26690 4760 26710 4800
rect 26750 4760 26770 4800
rect 26690 4730 26770 4760
rect 26870 5300 26950 5330
rect 26870 5260 26890 5300
rect 26930 5260 26950 5300
rect 26870 5200 26950 5260
rect 26870 5160 26890 5200
rect 26930 5160 26950 5200
rect 26870 5100 26950 5160
rect 26870 5060 26890 5100
rect 26930 5060 26950 5100
rect 26870 5000 26950 5060
rect 26870 4960 26890 5000
rect 26930 4960 26950 5000
rect 26870 4900 26950 4960
rect 26870 4860 26890 4900
rect 26930 4860 26950 4900
rect 26870 4800 26950 4860
rect 26870 4760 26890 4800
rect 26930 4760 26950 4800
rect 26870 4730 26950 4760
rect 27050 5300 27130 5330
rect 27050 5260 27070 5300
rect 27110 5260 27130 5300
rect 27050 5200 27130 5260
rect 27050 5160 27070 5200
rect 27110 5160 27130 5200
rect 27050 5100 27130 5160
rect 27050 5060 27070 5100
rect 27110 5060 27130 5100
rect 27050 5000 27130 5060
rect 27050 4960 27070 5000
rect 27110 4960 27130 5000
rect 27050 4900 27130 4960
rect 27050 4860 27070 4900
rect 27110 4860 27130 4900
rect 27050 4800 27130 4860
rect 27050 4760 27070 4800
rect 27110 4760 27130 4800
rect 27050 4730 27130 4760
rect 27230 5300 27310 5330
rect 27230 5260 27250 5300
rect 27290 5260 27310 5300
rect 27230 5200 27310 5260
rect 27230 5160 27250 5200
rect 27290 5160 27310 5200
rect 27230 5100 27310 5160
rect 27230 5060 27250 5100
rect 27290 5060 27310 5100
rect 27230 5000 27310 5060
rect 27230 4960 27250 5000
rect 27290 4960 27310 5000
rect 27230 4900 27310 4960
rect 27230 4860 27250 4900
rect 27290 4860 27310 4900
rect 27230 4800 27310 4860
rect 27230 4760 27250 4800
rect 27290 4760 27310 4800
rect 27230 4730 27310 4760
rect 27410 5300 27490 5330
rect 27410 5260 27430 5300
rect 27470 5260 27490 5300
rect 27410 5200 27490 5260
rect 27410 5160 27430 5200
rect 27470 5160 27490 5200
rect 27410 5100 27490 5160
rect 27410 5060 27430 5100
rect 27470 5060 27490 5100
rect 27410 5000 27490 5060
rect 27410 4960 27430 5000
rect 27470 4960 27490 5000
rect 27410 4900 27490 4960
rect 27410 4860 27430 4900
rect 27470 4860 27490 4900
rect 27410 4800 27490 4860
rect 27410 4760 27430 4800
rect 27470 4760 27490 4800
rect 27410 4730 27490 4760
rect 27590 5300 27670 5330
rect 27590 5260 27610 5300
rect 27650 5260 27670 5300
rect 27590 5200 27670 5260
rect 27590 5160 27610 5200
rect 27650 5160 27670 5200
rect 27590 5100 27670 5160
rect 27590 5060 27610 5100
rect 27650 5060 27670 5100
rect 27590 5000 27670 5060
rect 27590 4960 27610 5000
rect 27650 4960 27670 5000
rect 27590 4900 27670 4960
rect 27590 4860 27610 4900
rect 27650 4860 27670 4900
rect 27590 4800 27670 4860
rect 27590 4760 27610 4800
rect 27650 4760 27670 4800
rect 27590 4730 27670 4760
rect 27770 5300 27850 5330
rect 27770 5260 27790 5300
rect 27830 5260 27850 5300
rect 27770 5200 27850 5260
rect 27770 5160 27790 5200
rect 27830 5160 27850 5200
rect 27770 5100 27850 5160
rect 27770 5060 27790 5100
rect 27830 5060 27850 5100
rect 27770 5000 27850 5060
rect 27770 4960 27790 5000
rect 27830 4960 27850 5000
rect 27770 4900 27850 4960
rect 27770 4860 27790 4900
rect 27830 4860 27850 4900
rect 27770 4800 27850 4860
rect 27770 4760 27790 4800
rect 27830 4760 27850 4800
rect 27770 4730 27850 4760
rect 27950 5300 28030 5330
rect 27950 5260 27970 5300
rect 28010 5260 28030 5300
rect 27950 5200 28030 5260
rect 27950 5160 27970 5200
rect 28010 5160 28030 5200
rect 27950 5100 28030 5160
rect 27950 5060 27970 5100
rect 28010 5060 28030 5100
rect 27950 5000 28030 5060
rect 27950 4960 27970 5000
rect 28010 4960 28030 5000
rect 27950 4900 28030 4960
rect 27950 4860 27970 4900
rect 28010 4860 28030 4900
rect 27950 4800 28030 4860
rect 27950 4760 27970 4800
rect 28010 4760 28030 4800
rect 27950 4730 28030 4760
rect 28130 5300 28210 5330
rect 28130 5260 28150 5300
rect 28190 5260 28210 5300
rect 28130 5200 28210 5260
rect 28130 5160 28150 5200
rect 28190 5160 28210 5200
rect 28130 5100 28210 5160
rect 28130 5060 28150 5100
rect 28190 5060 28210 5100
rect 28130 5000 28210 5060
rect 28130 4960 28150 5000
rect 28190 4960 28210 5000
rect 28130 4900 28210 4960
rect 28130 4860 28150 4900
rect 28190 4860 28210 4900
rect 28130 4800 28210 4860
rect 28130 4760 28150 4800
rect 28190 4760 28210 4800
rect 28130 4730 28210 4760
rect 28310 5300 28390 5330
rect 28310 5260 28330 5300
rect 28370 5260 28390 5300
rect 28310 5200 28390 5260
rect 28310 5160 28330 5200
rect 28370 5160 28390 5200
rect 28310 5100 28390 5160
rect 28310 5060 28330 5100
rect 28370 5060 28390 5100
rect 28310 5000 28390 5060
rect 28310 4960 28330 5000
rect 28370 4960 28390 5000
rect 28310 4900 28390 4960
rect 28310 4860 28330 4900
rect 28370 4860 28390 4900
rect 28310 4800 28390 4860
rect 28310 4760 28330 4800
rect 28370 4760 28390 4800
rect 28310 4730 28390 4760
rect 28490 5300 28570 5330
rect 28490 5260 28510 5300
rect 28550 5260 28570 5300
rect 28490 5200 28570 5260
rect 28490 5160 28510 5200
rect 28550 5160 28570 5200
rect 28490 5100 28570 5160
rect 28490 5060 28510 5100
rect 28550 5060 28570 5100
rect 28490 5000 28570 5060
rect 28490 4960 28510 5000
rect 28550 4960 28570 5000
rect 28490 4900 28570 4960
rect 28490 4860 28510 4900
rect 28550 4860 28570 4900
rect 28490 4800 28570 4860
rect 28490 4760 28510 4800
rect 28550 4760 28570 4800
rect 28490 4730 28570 4760
rect 28670 5300 28750 5330
rect 28670 5260 28690 5300
rect 28730 5260 28750 5300
rect 28670 5200 28750 5260
rect 28670 5160 28690 5200
rect 28730 5160 28750 5200
rect 28670 5100 28750 5160
rect 28670 5060 28690 5100
rect 28730 5060 28750 5100
rect 28670 5000 28750 5060
rect 28670 4960 28690 5000
rect 28730 4960 28750 5000
rect 28670 4900 28750 4960
rect 28670 4860 28690 4900
rect 28730 4860 28750 4900
rect 28670 4800 28750 4860
rect 28670 4760 28690 4800
rect 28730 4760 28750 4800
rect 28670 4730 28750 4760
rect 28850 5300 28930 5330
rect 28850 5260 28870 5300
rect 28910 5260 28930 5300
rect 28850 5200 28930 5260
rect 28850 5160 28870 5200
rect 28910 5160 28930 5200
rect 28850 5100 28930 5160
rect 28850 5060 28870 5100
rect 28910 5060 28930 5100
rect 28850 5000 28930 5060
rect 28850 4960 28870 5000
rect 28910 4960 28930 5000
rect 28850 4900 28930 4960
rect 28850 4860 28870 4900
rect 28910 4860 28930 4900
rect 28850 4800 28930 4860
rect 28850 4760 28870 4800
rect 28910 4760 28930 4800
rect 28850 4730 28930 4760
rect 29030 5300 29110 5330
rect 29030 5260 29050 5300
rect 29090 5260 29110 5300
rect 29030 5200 29110 5260
rect 29030 5160 29050 5200
rect 29090 5160 29110 5200
rect 29030 5100 29110 5160
rect 29030 5060 29050 5100
rect 29090 5060 29110 5100
rect 29030 5000 29110 5060
rect 29030 4960 29050 5000
rect 29090 4960 29110 5000
rect 29030 4900 29110 4960
rect 29030 4860 29050 4900
rect 29090 4860 29110 4900
rect 29030 4800 29110 4860
rect 29030 4760 29050 4800
rect 29090 4760 29110 4800
rect 29030 4730 29110 4760
rect 29210 5300 29290 5330
rect 29210 5260 29230 5300
rect 29270 5260 29290 5300
rect 29210 5200 29290 5260
rect 29210 5160 29230 5200
rect 29270 5160 29290 5200
rect 29210 5100 29290 5160
rect 29210 5060 29230 5100
rect 29270 5060 29290 5100
rect 29210 5000 29290 5060
rect 29210 4960 29230 5000
rect 29270 4960 29290 5000
rect 29210 4900 29290 4960
rect 29210 4860 29230 4900
rect 29270 4860 29290 4900
rect 29210 4800 29290 4860
rect 29210 4760 29230 4800
rect 29270 4760 29290 4800
rect 29210 4730 29290 4760
rect 29390 5300 29470 5330
rect 29390 5260 29410 5300
rect 29450 5260 29470 5300
rect 29390 5200 29470 5260
rect 29390 5160 29410 5200
rect 29450 5160 29470 5200
rect 29390 5100 29470 5160
rect 29390 5060 29410 5100
rect 29450 5060 29470 5100
rect 29390 5000 29470 5060
rect 29390 4960 29410 5000
rect 29450 4960 29470 5000
rect 29390 4900 29470 4960
rect 29390 4860 29410 4900
rect 29450 4860 29470 4900
rect 29390 4800 29470 4860
rect 29390 4760 29410 4800
rect 29450 4760 29470 4800
rect 29390 4730 29470 4760
rect 29570 5300 29650 5330
rect 29570 5260 29590 5300
rect 29630 5260 29650 5300
rect 29570 5200 29650 5260
rect 29570 5160 29590 5200
rect 29630 5160 29650 5200
rect 29570 5100 29650 5160
rect 29570 5060 29590 5100
rect 29630 5060 29650 5100
rect 29570 5000 29650 5060
rect 29570 4960 29590 5000
rect 29630 4960 29650 5000
rect 29570 4900 29650 4960
rect 29570 4860 29590 4900
rect 29630 4860 29650 4900
rect 29570 4800 29650 4860
rect 29570 4760 29590 4800
rect 29630 4760 29650 4800
rect 29570 4730 29650 4760
rect 29750 5300 29830 5330
rect 29750 5260 29770 5300
rect 29810 5260 29830 5300
rect 29750 5200 29830 5260
rect 29750 5160 29770 5200
rect 29810 5160 29830 5200
rect 29750 5100 29830 5160
rect 29750 5060 29770 5100
rect 29810 5060 29830 5100
rect 29750 5000 29830 5060
rect 29750 4960 29770 5000
rect 29810 4960 29830 5000
rect 29750 4900 29830 4960
rect 29750 4860 29770 4900
rect 29810 4860 29830 4900
rect 29750 4800 29830 4860
rect 29750 4760 29770 4800
rect 29810 4760 29830 4800
rect 29750 4730 29830 4760
rect 25410 3970 25490 4000
rect 25410 3930 25430 3970
rect 25470 3930 25490 3970
rect 25410 3870 25490 3930
rect 25410 3830 25430 3870
rect 25470 3830 25490 3870
rect 25410 3800 25490 3830
rect 25530 3970 25610 4000
rect 25530 3930 25550 3970
rect 25590 3930 25610 3970
rect 25530 3870 25610 3930
rect 25530 3830 25550 3870
rect 25590 3830 25610 3870
rect 25530 3800 25610 3830
rect 25650 3970 25730 4000
rect 25650 3930 25670 3970
rect 25710 3930 25730 3970
rect 25650 3870 25730 3930
rect 25650 3830 25670 3870
rect 25710 3830 25730 3870
rect 25650 3800 25730 3830
rect 25770 3970 25850 4000
rect 25770 3930 25790 3970
rect 25830 3930 25850 3970
rect 25770 3870 25850 3930
rect 25770 3830 25790 3870
rect 25830 3830 25850 3870
rect 25770 3800 25850 3830
rect 25890 3970 25970 4000
rect 25890 3930 25910 3970
rect 25950 3930 25970 3970
rect 25890 3870 25970 3930
rect 25890 3830 25910 3870
rect 25950 3830 25970 3870
rect 25890 3800 25970 3830
rect 26010 3970 26090 4000
rect 26010 3930 26030 3970
rect 26070 3930 26090 3970
rect 26010 3870 26090 3930
rect 26010 3830 26030 3870
rect 26070 3830 26090 3870
rect 26010 3800 26090 3830
rect 26130 3970 26210 4000
rect 26130 3930 26150 3970
rect 26190 3930 26210 3970
rect 26130 3870 26210 3930
rect 26130 3830 26150 3870
rect 26190 3830 26210 3870
rect 26130 3800 26210 3830
rect 26250 3970 26330 4000
rect 26250 3930 26270 3970
rect 26310 3930 26330 3970
rect 26250 3870 26330 3930
rect 26250 3830 26270 3870
rect 26310 3830 26330 3870
rect 26250 3800 26330 3830
rect 26370 3970 26450 4000
rect 26370 3930 26390 3970
rect 26430 3930 26450 3970
rect 26370 3870 26450 3930
rect 26370 3830 26390 3870
rect 26430 3830 26450 3870
rect 26370 3800 26450 3830
rect 26490 3970 26570 4000
rect 26490 3930 26510 3970
rect 26550 3930 26570 3970
rect 26490 3870 26570 3930
rect 26490 3830 26510 3870
rect 26550 3830 26570 3870
rect 26490 3800 26570 3830
rect 26610 3970 26690 4000
rect 26610 3930 26630 3970
rect 26670 3930 26690 3970
rect 26610 3870 26690 3930
rect 26610 3830 26630 3870
rect 26670 3830 26690 3870
rect 26610 3800 26690 3830
rect 26730 3970 26810 4000
rect 26730 3930 26750 3970
rect 26790 3930 26810 3970
rect 26730 3870 26810 3930
rect 26730 3830 26750 3870
rect 26790 3830 26810 3870
rect 26730 3800 26810 3830
rect 26850 3970 26930 4000
rect 26850 3930 26870 3970
rect 26910 3930 26930 3970
rect 26850 3870 26930 3930
rect 26850 3830 26870 3870
rect 26910 3830 26930 3870
rect 26850 3800 26930 3830
rect 26970 3970 27050 4000
rect 26970 3930 26990 3970
rect 27030 3930 27050 3970
rect 26970 3870 27050 3930
rect 26970 3830 26990 3870
rect 27030 3830 27050 3870
rect 26970 3800 27050 3830
rect 27090 3970 27170 4000
rect 27090 3930 27110 3970
rect 27150 3930 27170 3970
rect 27090 3870 27170 3930
rect 27090 3830 27110 3870
rect 27150 3830 27170 3870
rect 27090 3800 27170 3830
rect 27210 3970 27290 4000
rect 27210 3930 27230 3970
rect 27270 3930 27290 3970
rect 27210 3870 27290 3930
rect 27210 3830 27230 3870
rect 27270 3830 27290 3870
rect 27210 3800 27290 3830
rect 27330 3970 27410 4000
rect 27330 3930 27350 3970
rect 27390 3930 27410 3970
rect 27330 3870 27410 3930
rect 27330 3830 27350 3870
rect 27390 3830 27410 3870
rect 27330 3800 27410 3830
rect 27450 3970 27530 4000
rect 27450 3930 27470 3970
rect 27510 3930 27530 3970
rect 27450 3870 27530 3930
rect 27450 3830 27470 3870
rect 27510 3830 27530 3870
rect 27450 3800 27530 3830
rect 27570 3970 27650 4000
rect 27570 3930 27590 3970
rect 27630 3930 27650 3970
rect 27570 3870 27650 3930
rect 27570 3830 27590 3870
rect 27630 3830 27650 3870
rect 27570 3800 27650 3830
rect 27690 3970 27770 4000
rect 27690 3930 27710 3970
rect 27750 3930 27770 3970
rect 27690 3870 27770 3930
rect 27690 3830 27710 3870
rect 27750 3830 27770 3870
rect 27690 3800 27770 3830
rect 27810 3970 27890 4000
rect 27810 3930 27830 3970
rect 27870 3930 27890 3970
rect 27810 3870 27890 3930
rect 27810 3830 27830 3870
rect 27870 3830 27890 3870
rect 27810 3800 27890 3830
rect 20560 3278 21240 3330
rect 20560 3244 20614 3278
rect 20648 3244 20704 3278
rect 20738 3244 20794 3278
rect 20828 3244 20884 3278
rect 20918 3244 20974 3278
rect 21008 3244 21064 3278
rect 21098 3244 21154 3278
rect 21188 3244 21240 3278
rect 20560 3188 21240 3244
rect 20560 3154 20614 3188
rect 20648 3154 20704 3188
rect 20738 3154 20794 3188
rect 20828 3154 20884 3188
rect 20918 3154 20974 3188
rect 21008 3154 21064 3188
rect 21098 3154 21154 3188
rect 21188 3154 21240 3188
rect 20560 3098 21240 3154
rect 20560 3064 20614 3098
rect 20648 3064 20704 3098
rect 20738 3064 20794 3098
rect 20828 3064 20884 3098
rect 20918 3064 20974 3098
rect 21008 3064 21064 3098
rect 21098 3064 21154 3098
rect 21188 3064 21240 3098
rect 20560 3008 21240 3064
rect 20560 2974 20614 3008
rect 20648 2974 20704 3008
rect 20738 2974 20794 3008
rect 20828 2974 20884 3008
rect 20918 2974 20974 3008
rect 21008 2974 21064 3008
rect 21098 2974 21154 3008
rect 21188 2974 21240 3008
rect 20560 2918 21240 2974
rect 20560 2884 20614 2918
rect 20648 2884 20704 2918
rect 20738 2884 20794 2918
rect 20828 2884 20884 2918
rect 20918 2884 20974 2918
rect 21008 2884 21064 2918
rect 21098 2884 21154 2918
rect 21188 2884 21240 2918
rect 20560 2828 21240 2884
rect 20560 2794 20614 2828
rect 20648 2794 20704 2828
rect 20738 2794 20794 2828
rect 20828 2794 20884 2828
rect 20918 2794 20974 2828
rect 21008 2794 21064 2828
rect 21098 2794 21154 2828
rect 21188 2794 21240 2828
rect 20560 2738 21240 2794
rect 20560 2704 20614 2738
rect 20648 2704 20704 2738
rect 20738 2704 20794 2738
rect 20828 2704 20884 2738
rect 20918 2704 20974 2738
rect 21008 2704 21064 2738
rect 21098 2704 21154 2738
rect 21188 2704 21240 2738
rect 20560 2650 21240 2704
rect 21920 3278 22600 3330
rect 21920 3244 21974 3278
rect 22008 3244 22064 3278
rect 22098 3244 22154 3278
rect 22188 3244 22244 3278
rect 22278 3244 22334 3278
rect 22368 3244 22424 3278
rect 22458 3244 22514 3278
rect 22548 3244 22600 3278
rect 21920 3188 22600 3244
rect 21920 3154 21974 3188
rect 22008 3154 22064 3188
rect 22098 3154 22154 3188
rect 22188 3154 22244 3188
rect 22278 3154 22334 3188
rect 22368 3154 22424 3188
rect 22458 3154 22514 3188
rect 22548 3154 22600 3188
rect 21920 3098 22600 3154
rect 21920 3064 21974 3098
rect 22008 3064 22064 3098
rect 22098 3064 22154 3098
rect 22188 3064 22244 3098
rect 22278 3064 22334 3098
rect 22368 3064 22424 3098
rect 22458 3064 22514 3098
rect 22548 3064 22600 3098
rect 21920 3008 22600 3064
rect 21920 2974 21974 3008
rect 22008 2974 22064 3008
rect 22098 2974 22154 3008
rect 22188 2974 22244 3008
rect 22278 2974 22334 3008
rect 22368 2974 22424 3008
rect 22458 2974 22514 3008
rect 22548 2974 22600 3008
rect 21920 2918 22600 2974
rect 21920 2884 21974 2918
rect 22008 2884 22064 2918
rect 22098 2884 22154 2918
rect 22188 2884 22244 2918
rect 22278 2884 22334 2918
rect 22368 2884 22424 2918
rect 22458 2884 22514 2918
rect 22548 2884 22600 2918
rect 21920 2828 22600 2884
rect 21920 2794 21974 2828
rect 22008 2794 22064 2828
rect 22098 2794 22154 2828
rect 22188 2794 22244 2828
rect 22278 2794 22334 2828
rect 22368 2794 22424 2828
rect 22458 2794 22514 2828
rect 22548 2794 22600 2828
rect 21920 2738 22600 2794
rect 21920 2704 21974 2738
rect 22008 2704 22064 2738
rect 22098 2704 22154 2738
rect 22188 2704 22244 2738
rect 22278 2704 22334 2738
rect 22368 2704 22424 2738
rect 22458 2704 22514 2738
rect 22548 2704 22600 2738
rect 21920 2650 22600 2704
rect 28450 3970 28530 4000
rect 28450 3930 28470 3970
rect 28510 3930 28530 3970
rect 28450 3870 28530 3930
rect 28450 3830 28470 3870
rect 28510 3830 28530 3870
rect 28450 3800 28530 3830
rect 28570 3970 28650 4000
rect 28570 3930 28590 3970
rect 28630 3930 28650 3970
rect 28570 3870 28650 3930
rect 28570 3830 28590 3870
rect 28630 3830 28650 3870
rect 28570 3800 28650 3830
rect 28690 3970 28770 4000
rect 28690 3930 28710 3970
rect 28750 3930 28770 3970
rect 28690 3870 28770 3930
rect 28690 3830 28710 3870
rect 28750 3830 28770 3870
rect 28690 3800 28770 3830
rect 28810 3970 28890 4000
rect 28810 3930 28830 3970
rect 28870 3930 28890 3970
rect 28810 3870 28890 3930
rect 28810 3830 28830 3870
rect 28870 3830 28890 3870
rect 28810 3800 28890 3830
rect 28930 3970 29010 4000
rect 28930 3930 28950 3970
rect 28990 3930 29010 3970
rect 28930 3870 29010 3930
rect 28930 3830 28950 3870
rect 28990 3830 29010 3870
rect 28930 3800 29010 3830
rect 29050 3970 29130 4000
rect 29050 3930 29070 3970
rect 29110 3930 29130 3970
rect 29050 3870 29130 3930
rect 29050 3830 29070 3870
rect 29110 3830 29130 3870
rect 29050 3800 29130 3830
rect 29170 3970 29250 4000
rect 29170 3930 29190 3970
rect 29230 3930 29250 3970
rect 29170 3870 29250 3930
rect 29170 3830 29190 3870
rect 29230 3830 29250 3870
rect 29170 3800 29250 3830
rect 29290 3970 29370 4000
rect 29290 3930 29310 3970
rect 29350 3930 29370 3970
rect 29290 3870 29370 3930
rect 29290 3830 29310 3870
rect 29350 3830 29370 3870
rect 29290 3800 29370 3830
rect 29410 3970 29490 4000
rect 29410 3930 29430 3970
rect 29470 3930 29490 3970
rect 29410 3870 29490 3930
rect 29410 3830 29430 3870
rect 29470 3830 29490 3870
rect 29410 3800 29490 3830
rect 29530 3970 29610 4000
rect 29530 3930 29550 3970
rect 29590 3930 29610 3970
rect 29530 3870 29610 3930
rect 29530 3830 29550 3870
rect 29590 3830 29610 3870
rect 29530 3800 29610 3830
rect 29650 3970 29730 4000
rect 29650 3930 29670 3970
rect 29710 3930 29730 3970
rect 29650 3870 29730 3930
rect 29650 3830 29670 3870
rect 29710 3830 29730 3870
rect 29650 3800 29730 3830
rect 29770 3970 29850 4000
rect 29770 3930 29790 3970
rect 29830 3930 29850 3970
rect 29770 3870 29850 3930
rect 29770 3830 29790 3870
rect 29830 3830 29850 3870
rect 29770 3800 29850 3830
rect 29890 3970 29970 4000
rect 29890 3930 29910 3970
rect 29950 3930 29970 3970
rect 29890 3870 29970 3930
rect 29890 3830 29910 3870
rect 29950 3830 29970 3870
rect 29890 3800 29970 3830
rect 30010 3970 30090 4000
rect 30010 3930 30030 3970
rect 30070 3930 30090 3970
rect 30010 3870 30090 3930
rect 30010 3830 30030 3870
rect 30070 3830 30090 3870
rect 30010 3800 30090 3830
rect 30130 3970 30210 4000
rect 30130 3930 30150 3970
rect 30190 3930 30210 3970
rect 30130 3870 30210 3930
rect 30130 3830 30150 3870
rect 30190 3830 30210 3870
rect 30130 3800 30210 3830
rect 30250 3970 30330 4000
rect 30250 3930 30270 3970
rect 30310 3930 30330 3970
rect 30250 3870 30330 3930
rect 30250 3830 30270 3870
rect 30310 3830 30330 3870
rect 30250 3800 30330 3830
rect 30370 3970 30450 4000
rect 30370 3930 30390 3970
rect 30430 3930 30450 3970
rect 30370 3870 30450 3930
rect 30370 3830 30390 3870
rect 30430 3830 30450 3870
rect 30370 3800 30450 3830
rect 30490 3970 30570 4000
rect 30490 3930 30510 3970
rect 30550 3930 30570 3970
rect 30490 3870 30570 3930
rect 30490 3830 30510 3870
rect 30550 3830 30570 3870
rect 30490 3800 30570 3830
rect 30610 3970 30690 4000
rect 30610 3930 30630 3970
rect 30670 3930 30690 3970
rect 30610 3870 30690 3930
rect 30610 3830 30630 3870
rect 30670 3830 30690 3870
rect 30610 3800 30690 3830
rect 30730 3970 30810 4000
rect 30730 3930 30750 3970
rect 30790 3930 30810 3970
rect 30730 3870 30810 3930
rect 30730 3830 30750 3870
rect 30790 3830 30810 3870
rect 30730 3800 30810 3830
rect 30850 3970 30930 4000
rect 30850 3930 30870 3970
rect 30910 3930 30930 3970
rect 30850 3870 30930 3930
rect 30850 3830 30870 3870
rect 30910 3830 30930 3870
rect 30850 3800 30930 3830
rect 23280 3278 23960 3330
rect 23280 3244 23334 3278
rect 23368 3244 23424 3278
rect 23458 3244 23514 3278
rect 23548 3244 23604 3278
rect 23638 3244 23694 3278
rect 23728 3244 23784 3278
rect 23818 3244 23874 3278
rect 23908 3244 23960 3278
rect 23280 3188 23960 3244
rect 23280 3154 23334 3188
rect 23368 3154 23424 3188
rect 23458 3154 23514 3188
rect 23548 3154 23604 3188
rect 23638 3154 23694 3188
rect 23728 3154 23784 3188
rect 23818 3154 23874 3188
rect 23908 3154 23960 3188
rect 23280 3098 23960 3154
rect 23280 3064 23334 3098
rect 23368 3064 23424 3098
rect 23458 3064 23514 3098
rect 23548 3064 23604 3098
rect 23638 3064 23694 3098
rect 23728 3064 23784 3098
rect 23818 3064 23874 3098
rect 23908 3064 23960 3098
rect 23280 3008 23960 3064
rect 23280 2974 23334 3008
rect 23368 2974 23424 3008
rect 23458 2974 23514 3008
rect 23548 2974 23604 3008
rect 23638 2974 23694 3008
rect 23728 2974 23784 3008
rect 23818 2974 23874 3008
rect 23908 2974 23960 3008
rect 23280 2918 23960 2974
rect 23280 2884 23334 2918
rect 23368 2884 23424 2918
rect 23458 2884 23514 2918
rect 23548 2884 23604 2918
rect 23638 2884 23694 2918
rect 23728 2884 23784 2918
rect 23818 2884 23874 2918
rect 23908 2884 23960 2918
rect 23280 2828 23960 2884
rect 23280 2794 23334 2828
rect 23368 2794 23424 2828
rect 23458 2794 23514 2828
rect 23548 2794 23604 2828
rect 23638 2794 23694 2828
rect 23728 2794 23784 2828
rect 23818 2794 23874 2828
rect 23908 2794 23960 2828
rect 23280 2738 23960 2794
rect 23280 2704 23334 2738
rect 23368 2704 23424 2738
rect 23458 2704 23514 2738
rect 23548 2704 23604 2738
rect 23638 2704 23694 2738
rect 23728 2704 23784 2738
rect 23818 2704 23874 2738
rect 23908 2704 23960 2738
rect 23280 2650 23960 2704
rect 20560 1918 21240 1970
rect 20560 1884 20614 1918
rect 20648 1884 20704 1918
rect 20738 1884 20794 1918
rect 20828 1884 20884 1918
rect 20918 1884 20974 1918
rect 21008 1884 21064 1918
rect 21098 1884 21154 1918
rect 21188 1884 21240 1918
rect 20560 1828 21240 1884
rect 20560 1794 20614 1828
rect 20648 1794 20704 1828
rect 20738 1794 20794 1828
rect 20828 1794 20884 1828
rect 20918 1794 20974 1828
rect 21008 1794 21064 1828
rect 21098 1794 21154 1828
rect 21188 1794 21240 1828
rect 20560 1738 21240 1794
rect 20560 1704 20614 1738
rect 20648 1704 20704 1738
rect 20738 1704 20794 1738
rect 20828 1704 20884 1738
rect 20918 1704 20974 1738
rect 21008 1704 21064 1738
rect 21098 1704 21154 1738
rect 21188 1704 21240 1738
rect 20560 1648 21240 1704
rect 20560 1614 20614 1648
rect 20648 1614 20704 1648
rect 20738 1614 20794 1648
rect 20828 1614 20884 1648
rect 20918 1614 20974 1648
rect 21008 1614 21064 1648
rect 21098 1614 21154 1648
rect 21188 1614 21240 1648
rect 20560 1558 21240 1614
rect 20560 1524 20614 1558
rect 20648 1524 20704 1558
rect 20738 1524 20794 1558
rect 20828 1524 20884 1558
rect 20918 1524 20974 1558
rect 21008 1524 21064 1558
rect 21098 1524 21154 1558
rect 21188 1524 21240 1558
rect 20560 1468 21240 1524
rect 20560 1434 20614 1468
rect 20648 1434 20704 1468
rect 20738 1434 20794 1468
rect 20828 1434 20884 1468
rect 20918 1434 20974 1468
rect 21008 1434 21064 1468
rect 21098 1434 21154 1468
rect 21188 1434 21240 1468
rect 20560 1378 21240 1434
rect 20560 1344 20614 1378
rect 20648 1344 20704 1378
rect 20738 1344 20794 1378
rect 20828 1344 20884 1378
rect 20918 1344 20974 1378
rect 21008 1344 21064 1378
rect 21098 1344 21154 1378
rect 21188 1344 21240 1378
rect 20560 1290 21240 1344
rect 21920 1918 22600 1970
rect 21920 1884 21974 1918
rect 22008 1884 22064 1918
rect 22098 1884 22154 1918
rect 22188 1884 22244 1918
rect 22278 1884 22334 1918
rect 22368 1884 22424 1918
rect 22458 1884 22514 1918
rect 22548 1884 22600 1918
rect 21920 1828 22600 1884
rect 21920 1794 21974 1828
rect 22008 1794 22064 1828
rect 22098 1794 22154 1828
rect 22188 1794 22244 1828
rect 22278 1794 22334 1828
rect 22368 1794 22424 1828
rect 22458 1794 22514 1828
rect 22548 1794 22600 1828
rect 21920 1738 22600 1794
rect 21920 1704 21974 1738
rect 22008 1704 22064 1738
rect 22098 1704 22154 1738
rect 22188 1704 22244 1738
rect 22278 1704 22334 1738
rect 22368 1704 22424 1738
rect 22458 1704 22514 1738
rect 22548 1704 22600 1738
rect 21920 1648 22600 1704
rect 21920 1614 21974 1648
rect 22008 1614 22064 1648
rect 22098 1614 22154 1648
rect 22188 1614 22244 1648
rect 22278 1614 22334 1648
rect 22368 1614 22424 1648
rect 22458 1614 22514 1648
rect 22548 1614 22600 1648
rect 21920 1558 22600 1614
rect 21920 1524 21974 1558
rect 22008 1524 22064 1558
rect 22098 1524 22154 1558
rect 22188 1524 22244 1558
rect 22278 1524 22334 1558
rect 22368 1524 22424 1558
rect 22458 1524 22514 1558
rect 22548 1524 22600 1558
rect 21920 1468 22600 1524
rect 21920 1434 21974 1468
rect 22008 1434 22064 1468
rect 22098 1434 22154 1468
rect 22188 1434 22244 1468
rect 22278 1434 22334 1468
rect 22368 1434 22424 1468
rect 22458 1434 22514 1468
rect 22548 1434 22600 1468
rect 21920 1378 22600 1434
rect 21920 1344 21974 1378
rect 22008 1344 22064 1378
rect 22098 1344 22154 1378
rect 22188 1344 22244 1378
rect 22278 1344 22334 1378
rect 22368 1344 22424 1378
rect 22458 1344 22514 1378
rect 22548 1344 22600 1378
rect 21920 1290 22600 1344
rect 23280 1918 23960 1970
rect 23280 1884 23334 1918
rect 23368 1884 23424 1918
rect 23458 1884 23514 1918
rect 23548 1884 23604 1918
rect 23638 1884 23694 1918
rect 23728 1884 23784 1918
rect 23818 1884 23874 1918
rect 23908 1884 23960 1918
rect 23280 1828 23960 1884
rect 23280 1794 23334 1828
rect 23368 1794 23424 1828
rect 23458 1794 23514 1828
rect 23548 1794 23604 1828
rect 23638 1794 23694 1828
rect 23728 1794 23784 1828
rect 23818 1794 23874 1828
rect 23908 1794 23960 1828
rect 23280 1738 23960 1794
rect 23280 1704 23334 1738
rect 23368 1704 23424 1738
rect 23458 1704 23514 1738
rect 23548 1704 23604 1738
rect 23638 1704 23694 1738
rect 23728 1704 23784 1738
rect 23818 1704 23874 1738
rect 23908 1704 23960 1738
rect 23280 1648 23960 1704
rect 23280 1614 23334 1648
rect 23368 1614 23424 1648
rect 23458 1614 23514 1648
rect 23548 1614 23604 1648
rect 23638 1614 23694 1648
rect 23728 1614 23784 1648
rect 23818 1614 23874 1648
rect 23908 1614 23960 1648
rect 23280 1558 23960 1614
rect 23280 1524 23334 1558
rect 23368 1524 23424 1558
rect 23458 1524 23514 1558
rect 23548 1524 23604 1558
rect 23638 1524 23694 1558
rect 23728 1524 23784 1558
rect 23818 1524 23874 1558
rect 23908 1524 23960 1558
rect 23280 1468 23960 1524
rect 23280 1434 23334 1468
rect 23368 1434 23424 1468
rect 23458 1434 23514 1468
rect 23548 1434 23604 1468
rect 23638 1434 23694 1468
rect 23728 1434 23784 1468
rect 23818 1434 23874 1468
rect 23908 1434 23960 1468
rect 23280 1378 23960 1434
rect 23280 1344 23334 1378
rect 23368 1344 23424 1378
rect 23458 1344 23514 1378
rect 23548 1344 23604 1378
rect 23638 1344 23694 1378
rect 23728 1344 23784 1378
rect 23818 1344 23874 1378
rect 23908 1344 23960 1378
rect 23280 1290 23960 1344
<< ndiffc >>
rect 26290 3180 26330 3220
rect 26410 3180 26450 3220
rect 26530 3180 26570 3220
rect 26650 3180 26690 3220
rect 26770 3180 26810 3220
rect 26890 3180 26930 3220
rect 27010 3180 27050 3220
rect 27130 3180 27170 3220
rect 27250 3180 27290 3220
rect 27370 3180 27410 3220
rect 27490 3180 27530 3220
rect 28810 3180 28850 3220
rect 28930 3180 28970 3220
rect 29050 3180 29090 3220
rect 29170 3180 29210 3220
rect 29290 3180 29330 3220
rect 29410 3180 29450 3220
rect 29530 3180 29570 3220
rect 29650 3180 29690 3220
rect 29770 3180 29810 3220
rect 29890 3180 29930 3220
rect 30010 3180 30050 3220
rect 25810 2630 25850 2670
rect 25810 2530 25850 2570
rect 25810 2430 25850 2470
rect 25810 2330 25850 2370
rect 25810 2230 25850 2270
rect 26890 2630 26930 2670
rect 26890 2530 26930 2570
rect 26890 2430 26930 2470
rect 26890 2330 26930 2370
rect 26890 2230 26930 2270
rect 27970 2630 28010 2670
rect 27970 2530 28010 2570
rect 27970 2430 28010 2470
rect 27970 2330 28010 2370
rect 27970 2230 28010 2270
rect 28330 2630 28370 2670
rect 28330 2530 28370 2570
rect 28330 2430 28370 2470
rect 28330 2330 28370 2370
rect 28330 2230 28370 2270
rect 29410 2630 29450 2670
rect 29410 2530 29450 2570
rect 29410 2430 29450 2470
rect 29410 2330 29450 2370
rect 29410 2230 29450 2270
rect 30490 2630 30530 2670
rect 30490 2530 30530 2570
rect 30490 2430 30530 2470
rect 30490 2330 30530 2370
rect 30490 2230 30530 2270
rect 26070 1640 26110 1680
rect 26070 1540 26110 1580
rect 28150 1640 28190 1680
rect 28150 1540 28190 1580
rect 30230 1640 30270 1680
rect 30230 1540 30270 1580
rect 25410 1090 25450 1130
rect 25410 990 25450 1030
rect 25590 1090 25630 1130
rect 25590 990 25630 1030
rect 25770 1090 25810 1130
rect 25770 990 25810 1030
rect 25950 1090 25990 1130
rect 25950 990 25990 1030
rect 26130 1090 26170 1130
rect 26130 990 26170 1030
rect 26310 1090 26350 1130
rect 26310 990 26350 1030
rect 26490 1090 26530 1130
rect 26490 990 26530 1030
rect 26670 1090 26710 1130
rect 26670 990 26710 1030
rect 26850 1090 26890 1130
rect 26850 990 26890 1030
rect 27250 1090 27290 1130
rect 27250 990 27290 1030
rect 27430 1090 27470 1130
rect 27430 990 27470 1030
rect 27610 1090 27650 1130
rect 27610 990 27650 1030
rect 27790 1090 27830 1130
rect 27790 990 27830 1030
rect 27970 1090 28010 1130
rect 27970 990 28010 1030
rect 28150 1090 28190 1130
rect 28150 990 28190 1030
rect 28330 1090 28370 1130
rect 28330 990 28370 1030
rect 28510 1090 28550 1130
rect 28510 990 28550 1030
rect 28690 1090 28730 1130
rect 28690 990 28730 1030
rect 28870 1090 28910 1130
rect 28870 990 28910 1030
rect 29050 1090 29090 1130
rect 29050 990 29090 1030
rect 29410 1090 29450 1130
rect 29410 990 29450 1030
rect 29590 1090 29630 1130
rect 29590 990 29630 1030
rect 29770 1090 29810 1130
rect 29770 990 29810 1030
rect 29950 1090 29990 1130
rect 29950 990 29990 1030
rect 30130 1090 30170 1130
rect 30130 990 30170 1030
rect 30310 1090 30350 1130
rect 30310 990 30350 1030
rect 30490 1090 30530 1130
rect 30490 990 30530 1030
rect 30670 1090 30710 1130
rect 30670 990 30710 1030
rect 30850 1090 30890 1130
rect 30850 990 30890 1030
<< pdiffc >>
rect 26170 6180 26210 6220
rect 26170 6080 26210 6120
rect 26350 6180 26390 6220
rect 26350 6080 26390 6120
rect 26530 6180 26570 6220
rect 26530 6080 26570 6120
rect 26710 6180 26750 6220
rect 26710 6080 26750 6120
rect 26890 6180 26930 6220
rect 26890 6080 26930 6120
rect 27070 6180 27110 6220
rect 27070 6080 27110 6120
rect 27250 6180 27290 6220
rect 27250 6080 27290 6120
rect 27430 6180 27470 6220
rect 27430 6080 27470 6120
rect 27610 6180 27650 6220
rect 27610 6080 27650 6120
rect 27790 6180 27830 6220
rect 27790 6080 27830 6120
rect 27970 6180 28010 6220
rect 27970 6080 28010 6120
rect 28150 6180 28190 6220
rect 28150 6080 28190 6120
rect 28330 6180 28370 6220
rect 28330 6080 28370 6120
rect 28510 6180 28550 6220
rect 28510 6080 28550 6120
rect 28690 6180 28730 6220
rect 28690 6080 28730 6120
rect 28870 6180 28910 6220
rect 28870 6080 28910 6120
rect 29050 6180 29090 6220
rect 29050 6080 29090 6120
rect 29230 6180 29270 6220
rect 29230 6080 29270 6120
rect 29410 6180 29450 6220
rect 29410 6080 29450 6120
rect 29590 6180 29630 6220
rect 29590 6080 29630 6120
rect 29770 6180 29810 6220
rect 29770 6080 29810 6120
rect 29950 6180 29990 6220
rect 29950 6080 29990 6120
rect 30130 6180 30170 6220
rect 30130 6080 30170 6120
rect 25530 5030 25570 5070
rect 20614 4604 20648 4638
rect 20704 4604 20738 4638
rect 20794 4604 20828 4638
rect 20884 4604 20918 4638
rect 20974 4604 21008 4638
rect 21064 4604 21098 4638
rect 21154 4604 21188 4638
rect 20614 4514 20648 4548
rect 20704 4514 20738 4548
rect 20794 4514 20828 4548
rect 20884 4514 20918 4548
rect 20974 4514 21008 4548
rect 21064 4514 21098 4548
rect 21154 4514 21188 4548
rect 20614 4424 20648 4458
rect 20704 4424 20738 4458
rect 20794 4424 20828 4458
rect 20884 4424 20918 4458
rect 20974 4424 21008 4458
rect 21064 4424 21098 4458
rect 21154 4424 21188 4458
rect 20614 4334 20648 4368
rect 20704 4334 20738 4368
rect 20794 4334 20828 4368
rect 20884 4334 20918 4368
rect 20974 4334 21008 4368
rect 21064 4334 21098 4368
rect 21154 4334 21188 4368
rect 20614 4244 20648 4278
rect 20704 4244 20738 4278
rect 20794 4244 20828 4278
rect 20884 4244 20918 4278
rect 20974 4244 21008 4278
rect 21064 4244 21098 4278
rect 21154 4244 21188 4278
rect 20614 4154 20648 4188
rect 20704 4154 20738 4188
rect 20794 4154 20828 4188
rect 20884 4154 20918 4188
rect 20974 4154 21008 4188
rect 21064 4154 21098 4188
rect 21154 4154 21188 4188
rect 20614 4064 20648 4098
rect 20704 4064 20738 4098
rect 20794 4064 20828 4098
rect 20884 4064 20918 4098
rect 20974 4064 21008 4098
rect 21064 4064 21098 4098
rect 21154 4064 21188 4098
rect 21974 4604 22008 4638
rect 22064 4604 22098 4638
rect 22154 4604 22188 4638
rect 22244 4604 22278 4638
rect 22334 4604 22368 4638
rect 22424 4604 22458 4638
rect 22514 4604 22548 4638
rect 21974 4514 22008 4548
rect 22064 4514 22098 4548
rect 22154 4514 22188 4548
rect 22244 4514 22278 4548
rect 22334 4514 22368 4548
rect 22424 4514 22458 4548
rect 22514 4514 22548 4548
rect 21974 4424 22008 4458
rect 22064 4424 22098 4458
rect 22154 4424 22188 4458
rect 22244 4424 22278 4458
rect 22334 4424 22368 4458
rect 22424 4424 22458 4458
rect 22514 4424 22548 4458
rect 21974 4334 22008 4368
rect 22064 4334 22098 4368
rect 22154 4334 22188 4368
rect 22244 4334 22278 4368
rect 22334 4334 22368 4368
rect 22424 4334 22458 4368
rect 22514 4334 22548 4368
rect 21974 4244 22008 4278
rect 22064 4244 22098 4278
rect 22154 4244 22188 4278
rect 22244 4244 22278 4278
rect 22334 4244 22368 4278
rect 22424 4244 22458 4278
rect 22514 4244 22548 4278
rect 21974 4154 22008 4188
rect 22064 4154 22098 4188
rect 22154 4154 22188 4188
rect 22244 4154 22278 4188
rect 22334 4154 22368 4188
rect 22424 4154 22458 4188
rect 22514 4154 22548 4188
rect 21974 4064 22008 4098
rect 22064 4064 22098 4098
rect 22154 4064 22188 4098
rect 22244 4064 22278 4098
rect 22334 4064 22368 4098
rect 22424 4064 22458 4098
rect 22514 4064 22548 4098
rect 25530 4930 25570 4970
rect 25640 5030 25680 5070
rect 25640 4930 25680 4970
rect 25750 5030 25790 5070
rect 25750 4930 25790 4970
rect 23334 4604 23368 4638
rect 23424 4604 23458 4638
rect 23514 4604 23548 4638
rect 23604 4604 23638 4638
rect 23694 4604 23728 4638
rect 23784 4604 23818 4638
rect 23874 4604 23908 4638
rect 23334 4514 23368 4548
rect 23424 4514 23458 4548
rect 23514 4514 23548 4548
rect 23604 4514 23638 4548
rect 23694 4514 23728 4548
rect 23784 4514 23818 4548
rect 23874 4514 23908 4548
rect 23334 4424 23368 4458
rect 23424 4424 23458 4458
rect 23514 4424 23548 4458
rect 23604 4424 23638 4458
rect 23694 4424 23728 4458
rect 23784 4424 23818 4458
rect 23874 4424 23908 4458
rect 23334 4334 23368 4368
rect 23424 4334 23458 4368
rect 23514 4334 23548 4368
rect 23604 4334 23638 4368
rect 23694 4334 23728 4368
rect 23784 4334 23818 4368
rect 23874 4334 23908 4368
rect 23334 4244 23368 4278
rect 23424 4244 23458 4278
rect 23514 4244 23548 4278
rect 23604 4244 23638 4278
rect 23694 4244 23728 4278
rect 23784 4244 23818 4278
rect 23874 4244 23908 4278
rect 23334 4154 23368 4188
rect 23424 4154 23458 4188
rect 23514 4154 23548 4188
rect 23604 4154 23638 4188
rect 23694 4154 23728 4188
rect 23784 4154 23818 4188
rect 23874 4154 23908 4188
rect 23334 4064 23368 4098
rect 23424 4064 23458 4098
rect 23514 4064 23548 4098
rect 23604 4064 23638 4098
rect 23694 4064 23728 4098
rect 23784 4064 23818 4098
rect 23874 4064 23908 4098
rect 26530 5260 26570 5300
rect 26530 5160 26570 5200
rect 26530 5060 26570 5100
rect 26530 4960 26570 5000
rect 26530 4860 26570 4900
rect 26530 4760 26570 4800
rect 26710 5260 26750 5300
rect 26710 5160 26750 5200
rect 26710 5060 26750 5100
rect 26710 4960 26750 5000
rect 26710 4860 26750 4900
rect 26710 4760 26750 4800
rect 26890 5260 26930 5300
rect 26890 5160 26930 5200
rect 26890 5060 26930 5100
rect 26890 4960 26930 5000
rect 26890 4860 26930 4900
rect 26890 4760 26930 4800
rect 27070 5260 27110 5300
rect 27070 5160 27110 5200
rect 27070 5060 27110 5100
rect 27070 4960 27110 5000
rect 27070 4860 27110 4900
rect 27070 4760 27110 4800
rect 27250 5260 27290 5300
rect 27250 5160 27290 5200
rect 27250 5060 27290 5100
rect 27250 4960 27290 5000
rect 27250 4860 27290 4900
rect 27250 4760 27290 4800
rect 27430 5260 27470 5300
rect 27430 5160 27470 5200
rect 27430 5060 27470 5100
rect 27430 4960 27470 5000
rect 27430 4860 27470 4900
rect 27430 4760 27470 4800
rect 27610 5260 27650 5300
rect 27610 5160 27650 5200
rect 27610 5060 27650 5100
rect 27610 4960 27650 5000
rect 27610 4860 27650 4900
rect 27610 4760 27650 4800
rect 27790 5260 27830 5300
rect 27790 5160 27830 5200
rect 27790 5060 27830 5100
rect 27790 4960 27830 5000
rect 27790 4860 27830 4900
rect 27790 4760 27830 4800
rect 27970 5260 28010 5300
rect 27970 5160 28010 5200
rect 27970 5060 28010 5100
rect 27970 4960 28010 5000
rect 27970 4860 28010 4900
rect 27970 4760 28010 4800
rect 28150 5260 28190 5300
rect 28150 5160 28190 5200
rect 28150 5060 28190 5100
rect 28150 4960 28190 5000
rect 28150 4860 28190 4900
rect 28150 4760 28190 4800
rect 28330 5260 28370 5300
rect 28330 5160 28370 5200
rect 28330 5060 28370 5100
rect 28330 4960 28370 5000
rect 28330 4860 28370 4900
rect 28330 4760 28370 4800
rect 28510 5260 28550 5300
rect 28510 5160 28550 5200
rect 28510 5060 28550 5100
rect 28510 4960 28550 5000
rect 28510 4860 28550 4900
rect 28510 4760 28550 4800
rect 28690 5260 28730 5300
rect 28690 5160 28730 5200
rect 28690 5060 28730 5100
rect 28690 4960 28730 5000
rect 28690 4860 28730 4900
rect 28690 4760 28730 4800
rect 28870 5260 28910 5300
rect 28870 5160 28910 5200
rect 28870 5060 28910 5100
rect 28870 4960 28910 5000
rect 28870 4860 28910 4900
rect 28870 4760 28910 4800
rect 29050 5260 29090 5300
rect 29050 5160 29090 5200
rect 29050 5060 29090 5100
rect 29050 4960 29090 5000
rect 29050 4860 29090 4900
rect 29050 4760 29090 4800
rect 29230 5260 29270 5300
rect 29230 5160 29270 5200
rect 29230 5060 29270 5100
rect 29230 4960 29270 5000
rect 29230 4860 29270 4900
rect 29230 4760 29270 4800
rect 29410 5260 29450 5300
rect 29410 5160 29450 5200
rect 29410 5060 29450 5100
rect 29410 4960 29450 5000
rect 29410 4860 29450 4900
rect 29410 4760 29450 4800
rect 29590 5260 29630 5300
rect 29590 5160 29630 5200
rect 29590 5060 29630 5100
rect 29590 4960 29630 5000
rect 29590 4860 29630 4900
rect 29590 4760 29630 4800
rect 29770 5260 29810 5300
rect 29770 5160 29810 5200
rect 29770 5060 29810 5100
rect 29770 4960 29810 5000
rect 29770 4860 29810 4900
rect 29770 4760 29810 4800
rect 25430 3930 25470 3970
rect 25430 3830 25470 3870
rect 25550 3930 25590 3970
rect 25550 3830 25590 3870
rect 25670 3930 25710 3970
rect 25670 3830 25710 3870
rect 25790 3930 25830 3970
rect 25790 3830 25830 3870
rect 25910 3930 25950 3970
rect 25910 3830 25950 3870
rect 26030 3930 26070 3970
rect 26030 3830 26070 3870
rect 26150 3930 26190 3970
rect 26150 3830 26190 3870
rect 26270 3930 26310 3970
rect 26270 3830 26310 3870
rect 26390 3930 26430 3970
rect 26390 3830 26430 3870
rect 26510 3930 26550 3970
rect 26510 3830 26550 3870
rect 26630 3930 26670 3970
rect 26630 3830 26670 3870
rect 26750 3930 26790 3970
rect 26750 3830 26790 3870
rect 26870 3930 26910 3970
rect 26870 3830 26910 3870
rect 26990 3930 27030 3970
rect 26990 3830 27030 3870
rect 27110 3930 27150 3970
rect 27110 3830 27150 3870
rect 27230 3930 27270 3970
rect 27230 3830 27270 3870
rect 27350 3930 27390 3970
rect 27350 3830 27390 3870
rect 27470 3930 27510 3970
rect 27470 3830 27510 3870
rect 27590 3930 27630 3970
rect 27590 3830 27630 3870
rect 27710 3930 27750 3970
rect 27710 3830 27750 3870
rect 27830 3930 27870 3970
rect 27830 3830 27870 3870
rect 20614 3244 20648 3278
rect 20704 3244 20738 3278
rect 20794 3244 20828 3278
rect 20884 3244 20918 3278
rect 20974 3244 21008 3278
rect 21064 3244 21098 3278
rect 21154 3244 21188 3278
rect 20614 3154 20648 3188
rect 20704 3154 20738 3188
rect 20794 3154 20828 3188
rect 20884 3154 20918 3188
rect 20974 3154 21008 3188
rect 21064 3154 21098 3188
rect 21154 3154 21188 3188
rect 20614 3064 20648 3098
rect 20704 3064 20738 3098
rect 20794 3064 20828 3098
rect 20884 3064 20918 3098
rect 20974 3064 21008 3098
rect 21064 3064 21098 3098
rect 21154 3064 21188 3098
rect 20614 2974 20648 3008
rect 20704 2974 20738 3008
rect 20794 2974 20828 3008
rect 20884 2974 20918 3008
rect 20974 2974 21008 3008
rect 21064 2974 21098 3008
rect 21154 2974 21188 3008
rect 20614 2884 20648 2918
rect 20704 2884 20738 2918
rect 20794 2884 20828 2918
rect 20884 2884 20918 2918
rect 20974 2884 21008 2918
rect 21064 2884 21098 2918
rect 21154 2884 21188 2918
rect 20614 2794 20648 2828
rect 20704 2794 20738 2828
rect 20794 2794 20828 2828
rect 20884 2794 20918 2828
rect 20974 2794 21008 2828
rect 21064 2794 21098 2828
rect 21154 2794 21188 2828
rect 20614 2704 20648 2738
rect 20704 2704 20738 2738
rect 20794 2704 20828 2738
rect 20884 2704 20918 2738
rect 20974 2704 21008 2738
rect 21064 2704 21098 2738
rect 21154 2704 21188 2738
rect 21974 3244 22008 3278
rect 22064 3244 22098 3278
rect 22154 3244 22188 3278
rect 22244 3244 22278 3278
rect 22334 3244 22368 3278
rect 22424 3244 22458 3278
rect 22514 3244 22548 3278
rect 21974 3154 22008 3188
rect 22064 3154 22098 3188
rect 22154 3154 22188 3188
rect 22244 3154 22278 3188
rect 22334 3154 22368 3188
rect 22424 3154 22458 3188
rect 22514 3154 22548 3188
rect 21974 3064 22008 3098
rect 22064 3064 22098 3098
rect 22154 3064 22188 3098
rect 22244 3064 22278 3098
rect 22334 3064 22368 3098
rect 22424 3064 22458 3098
rect 22514 3064 22548 3098
rect 21974 2974 22008 3008
rect 22064 2974 22098 3008
rect 22154 2974 22188 3008
rect 22244 2974 22278 3008
rect 22334 2974 22368 3008
rect 22424 2974 22458 3008
rect 22514 2974 22548 3008
rect 21974 2884 22008 2918
rect 22064 2884 22098 2918
rect 22154 2884 22188 2918
rect 22244 2884 22278 2918
rect 22334 2884 22368 2918
rect 22424 2884 22458 2918
rect 22514 2884 22548 2918
rect 21974 2794 22008 2828
rect 22064 2794 22098 2828
rect 22154 2794 22188 2828
rect 22244 2794 22278 2828
rect 22334 2794 22368 2828
rect 22424 2794 22458 2828
rect 22514 2794 22548 2828
rect 21974 2704 22008 2738
rect 22064 2704 22098 2738
rect 22154 2704 22188 2738
rect 22244 2704 22278 2738
rect 22334 2704 22368 2738
rect 22424 2704 22458 2738
rect 22514 2704 22548 2738
rect 28470 3930 28510 3970
rect 28470 3830 28510 3870
rect 28590 3930 28630 3970
rect 28590 3830 28630 3870
rect 28710 3930 28750 3970
rect 28710 3830 28750 3870
rect 28830 3930 28870 3970
rect 28830 3830 28870 3870
rect 28950 3930 28990 3970
rect 28950 3830 28990 3870
rect 29070 3930 29110 3970
rect 29070 3830 29110 3870
rect 29190 3930 29230 3970
rect 29190 3830 29230 3870
rect 29310 3930 29350 3970
rect 29310 3830 29350 3870
rect 29430 3930 29470 3970
rect 29430 3830 29470 3870
rect 29550 3930 29590 3970
rect 29550 3830 29590 3870
rect 29670 3930 29710 3970
rect 29670 3830 29710 3870
rect 29790 3930 29830 3970
rect 29790 3830 29830 3870
rect 29910 3930 29950 3970
rect 29910 3830 29950 3870
rect 30030 3930 30070 3970
rect 30030 3830 30070 3870
rect 30150 3930 30190 3970
rect 30150 3830 30190 3870
rect 30270 3930 30310 3970
rect 30270 3830 30310 3870
rect 30390 3930 30430 3970
rect 30390 3830 30430 3870
rect 30510 3930 30550 3970
rect 30510 3830 30550 3870
rect 30630 3930 30670 3970
rect 30630 3830 30670 3870
rect 30750 3930 30790 3970
rect 30750 3830 30790 3870
rect 30870 3930 30910 3970
rect 30870 3830 30910 3870
rect 23334 3244 23368 3278
rect 23424 3244 23458 3278
rect 23514 3244 23548 3278
rect 23604 3244 23638 3278
rect 23694 3244 23728 3278
rect 23784 3244 23818 3278
rect 23874 3244 23908 3278
rect 23334 3154 23368 3188
rect 23424 3154 23458 3188
rect 23514 3154 23548 3188
rect 23604 3154 23638 3188
rect 23694 3154 23728 3188
rect 23784 3154 23818 3188
rect 23874 3154 23908 3188
rect 23334 3064 23368 3098
rect 23424 3064 23458 3098
rect 23514 3064 23548 3098
rect 23604 3064 23638 3098
rect 23694 3064 23728 3098
rect 23784 3064 23818 3098
rect 23874 3064 23908 3098
rect 23334 2974 23368 3008
rect 23424 2974 23458 3008
rect 23514 2974 23548 3008
rect 23604 2974 23638 3008
rect 23694 2974 23728 3008
rect 23784 2974 23818 3008
rect 23874 2974 23908 3008
rect 23334 2884 23368 2918
rect 23424 2884 23458 2918
rect 23514 2884 23548 2918
rect 23604 2884 23638 2918
rect 23694 2884 23728 2918
rect 23784 2884 23818 2918
rect 23874 2884 23908 2918
rect 23334 2794 23368 2828
rect 23424 2794 23458 2828
rect 23514 2794 23548 2828
rect 23604 2794 23638 2828
rect 23694 2794 23728 2828
rect 23784 2794 23818 2828
rect 23874 2794 23908 2828
rect 23334 2704 23368 2738
rect 23424 2704 23458 2738
rect 23514 2704 23548 2738
rect 23604 2704 23638 2738
rect 23694 2704 23728 2738
rect 23784 2704 23818 2738
rect 23874 2704 23908 2738
rect 20614 1884 20648 1918
rect 20704 1884 20738 1918
rect 20794 1884 20828 1918
rect 20884 1884 20918 1918
rect 20974 1884 21008 1918
rect 21064 1884 21098 1918
rect 21154 1884 21188 1918
rect 20614 1794 20648 1828
rect 20704 1794 20738 1828
rect 20794 1794 20828 1828
rect 20884 1794 20918 1828
rect 20974 1794 21008 1828
rect 21064 1794 21098 1828
rect 21154 1794 21188 1828
rect 20614 1704 20648 1738
rect 20704 1704 20738 1738
rect 20794 1704 20828 1738
rect 20884 1704 20918 1738
rect 20974 1704 21008 1738
rect 21064 1704 21098 1738
rect 21154 1704 21188 1738
rect 20614 1614 20648 1648
rect 20704 1614 20738 1648
rect 20794 1614 20828 1648
rect 20884 1614 20918 1648
rect 20974 1614 21008 1648
rect 21064 1614 21098 1648
rect 21154 1614 21188 1648
rect 20614 1524 20648 1558
rect 20704 1524 20738 1558
rect 20794 1524 20828 1558
rect 20884 1524 20918 1558
rect 20974 1524 21008 1558
rect 21064 1524 21098 1558
rect 21154 1524 21188 1558
rect 20614 1434 20648 1468
rect 20704 1434 20738 1468
rect 20794 1434 20828 1468
rect 20884 1434 20918 1468
rect 20974 1434 21008 1468
rect 21064 1434 21098 1468
rect 21154 1434 21188 1468
rect 20614 1344 20648 1378
rect 20704 1344 20738 1378
rect 20794 1344 20828 1378
rect 20884 1344 20918 1378
rect 20974 1344 21008 1378
rect 21064 1344 21098 1378
rect 21154 1344 21188 1378
rect 21974 1884 22008 1918
rect 22064 1884 22098 1918
rect 22154 1884 22188 1918
rect 22244 1884 22278 1918
rect 22334 1884 22368 1918
rect 22424 1884 22458 1918
rect 22514 1884 22548 1918
rect 21974 1794 22008 1828
rect 22064 1794 22098 1828
rect 22154 1794 22188 1828
rect 22244 1794 22278 1828
rect 22334 1794 22368 1828
rect 22424 1794 22458 1828
rect 22514 1794 22548 1828
rect 21974 1704 22008 1738
rect 22064 1704 22098 1738
rect 22154 1704 22188 1738
rect 22244 1704 22278 1738
rect 22334 1704 22368 1738
rect 22424 1704 22458 1738
rect 22514 1704 22548 1738
rect 21974 1614 22008 1648
rect 22064 1614 22098 1648
rect 22154 1614 22188 1648
rect 22244 1614 22278 1648
rect 22334 1614 22368 1648
rect 22424 1614 22458 1648
rect 22514 1614 22548 1648
rect 21974 1524 22008 1558
rect 22064 1524 22098 1558
rect 22154 1524 22188 1558
rect 22244 1524 22278 1558
rect 22334 1524 22368 1558
rect 22424 1524 22458 1558
rect 22514 1524 22548 1558
rect 21974 1434 22008 1468
rect 22064 1434 22098 1468
rect 22154 1434 22188 1468
rect 22244 1434 22278 1468
rect 22334 1434 22368 1468
rect 22424 1434 22458 1468
rect 22514 1434 22548 1468
rect 21974 1344 22008 1378
rect 22064 1344 22098 1378
rect 22154 1344 22188 1378
rect 22244 1344 22278 1378
rect 22334 1344 22368 1378
rect 22424 1344 22458 1378
rect 22514 1344 22548 1378
rect 23334 1884 23368 1918
rect 23424 1884 23458 1918
rect 23514 1884 23548 1918
rect 23604 1884 23638 1918
rect 23694 1884 23728 1918
rect 23784 1884 23818 1918
rect 23874 1884 23908 1918
rect 23334 1794 23368 1828
rect 23424 1794 23458 1828
rect 23514 1794 23548 1828
rect 23604 1794 23638 1828
rect 23694 1794 23728 1828
rect 23784 1794 23818 1828
rect 23874 1794 23908 1828
rect 23334 1704 23368 1738
rect 23424 1704 23458 1738
rect 23514 1704 23548 1738
rect 23604 1704 23638 1738
rect 23694 1704 23728 1738
rect 23784 1704 23818 1738
rect 23874 1704 23908 1738
rect 23334 1614 23368 1648
rect 23424 1614 23458 1648
rect 23514 1614 23548 1648
rect 23604 1614 23638 1648
rect 23694 1614 23728 1648
rect 23784 1614 23818 1648
rect 23874 1614 23908 1648
rect 23334 1524 23368 1558
rect 23424 1524 23458 1558
rect 23514 1524 23548 1558
rect 23604 1524 23638 1558
rect 23694 1524 23728 1558
rect 23784 1524 23818 1558
rect 23874 1524 23908 1558
rect 23334 1434 23368 1468
rect 23424 1434 23458 1468
rect 23514 1434 23548 1468
rect 23604 1434 23638 1468
rect 23694 1434 23728 1468
rect 23784 1434 23818 1468
rect 23874 1434 23908 1468
rect 23334 1344 23368 1378
rect 23424 1344 23458 1378
rect 23514 1344 23548 1378
rect 23604 1344 23638 1378
rect 23694 1344 23728 1378
rect 23784 1344 23818 1378
rect 23874 1344 23908 1378
<< psubdiff >>
rect 21810 5820 22250 5840
rect 21810 5760 21840 5820
rect 21900 5760 22000 5820
rect 22060 5760 22160 5820
rect 22220 5760 22250 5820
rect 21810 5740 22250 5760
rect 20256 4959 21544 4994
rect 20256 4936 20386 4959
rect 20256 4902 20290 4936
rect 20324 4925 20386 4936
rect 20420 4925 20476 4959
rect 20510 4925 20566 4959
rect 20600 4925 20656 4959
rect 20690 4925 20746 4959
rect 20780 4925 20836 4959
rect 20870 4925 20926 4959
rect 20960 4925 21016 4959
rect 21050 4925 21106 4959
rect 21140 4925 21196 4959
rect 21230 4925 21286 4959
rect 21320 4925 21376 4959
rect 21410 4936 21544 4959
rect 21410 4925 21477 4936
rect 20324 4902 21477 4925
rect 21511 4902 21544 4936
rect 20256 4893 21544 4902
rect 20256 4846 20357 4893
rect 20256 4812 20290 4846
rect 20324 4812 20357 4846
rect 21443 4846 21544 4893
rect 20256 4756 20357 4812
rect 20256 4722 20290 4756
rect 20324 4722 20357 4756
rect 20256 4666 20357 4722
rect 20256 4632 20290 4666
rect 20324 4632 20357 4666
rect 20256 4576 20357 4632
rect 20256 4542 20290 4576
rect 20324 4542 20357 4576
rect 20256 4486 20357 4542
rect 20256 4452 20290 4486
rect 20324 4452 20357 4486
rect 20256 4396 20357 4452
rect 20256 4362 20290 4396
rect 20324 4362 20357 4396
rect 20256 4306 20357 4362
rect 20256 4272 20290 4306
rect 20324 4272 20357 4306
rect 20256 4216 20357 4272
rect 20256 4182 20290 4216
rect 20324 4182 20357 4216
rect 20256 4126 20357 4182
rect 20256 4092 20290 4126
rect 20324 4092 20357 4126
rect 20256 4036 20357 4092
rect 20256 4002 20290 4036
rect 20324 4002 20357 4036
rect 20256 3946 20357 4002
rect 20256 3912 20290 3946
rect 20324 3912 20357 3946
rect 20256 3856 20357 3912
rect 21443 4812 21477 4846
rect 21511 4812 21544 4846
rect 21443 4756 21544 4812
rect 21443 4722 21477 4756
rect 21511 4722 21544 4756
rect 21443 4666 21544 4722
rect 21443 4632 21477 4666
rect 21511 4632 21544 4666
rect 21443 4576 21544 4632
rect 21443 4542 21477 4576
rect 21511 4542 21544 4576
rect 21443 4486 21544 4542
rect 21443 4452 21477 4486
rect 21511 4452 21544 4486
rect 21443 4396 21544 4452
rect 21443 4362 21477 4396
rect 21511 4362 21544 4396
rect 21443 4306 21544 4362
rect 21443 4272 21477 4306
rect 21511 4272 21544 4306
rect 21443 4216 21544 4272
rect 21443 4182 21477 4216
rect 21511 4182 21544 4216
rect 21443 4126 21544 4182
rect 21443 4092 21477 4126
rect 21511 4092 21544 4126
rect 21443 4036 21544 4092
rect 21443 4002 21477 4036
rect 21511 4002 21544 4036
rect 21443 3946 21544 4002
rect 21443 3912 21477 3946
rect 21511 3912 21544 3946
rect 20256 3822 20290 3856
rect 20324 3822 20357 3856
rect 20256 3807 20357 3822
rect 21443 3856 21544 3912
rect 21443 3822 21477 3856
rect 21511 3822 21544 3856
rect 21443 3807 21544 3822
rect 20256 3772 21544 3807
rect 20256 3738 20386 3772
rect 20420 3738 20476 3772
rect 20510 3738 20566 3772
rect 20600 3738 20656 3772
rect 20690 3738 20746 3772
rect 20780 3738 20836 3772
rect 20870 3738 20926 3772
rect 20960 3738 21016 3772
rect 21050 3738 21106 3772
rect 21140 3738 21196 3772
rect 21230 3738 21286 3772
rect 21320 3738 21376 3772
rect 21410 3738 21544 3772
rect 20256 3706 21544 3738
rect 21616 4959 22904 4994
rect 21616 4936 21746 4959
rect 21616 4902 21650 4936
rect 21684 4925 21746 4936
rect 21780 4925 21836 4959
rect 21870 4925 21926 4959
rect 21960 4925 22016 4959
rect 22050 4925 22106 4959
rect 22140 4925 22196 4959
rect 22230 4925 22286 4959
rect 22320 4925 22376 4959
rect 22410 4925 22466 4959
rect 22500 4925 22556 4959
rect 22590 4925 22646 4959
rect 22680 4925 22736 4959
rect 22770 4936 22904 4959
rect 22770 4925 22837 4936
rect 21684 4902 22837 4925
rect 22871 4902 22904 4936
rect 21616 4893 22904 4902
rect 21616 4846 21717 4893
rect 21616 4812 21650 4846
rect 21684 4812 21717 4846
rect 22803 4846 22904 4893
rect 21616 4756 21717 4812
rect 21616 4722 21650 4756
rect 21684 4722 21717 4756
rect 21616 4666 21717 4722
rect 21616 4632 21650 4666
rect 21684 4632 21717 4666
rect 21616 4576 21717 4632
rect 21616 4542 21650 4576
rect 21684 4542 21717 4576
rect 21616 4486 21717 4542
rect 21616 4452 21650 4486
rect 21684 4452 21717 4486
rect 21616 4396 21717 4452
rect 21616 4362 21650 4396
rect 21684 4362 21717 4396
rect 21616 4306 21717 4362
rect 21616 4272 21650 4306
rect 21684 4272 21717 4306
rect 21616 4216 21717 4272
rect 21616 4182 21650 4216
rect 21684 4182 21717 4216
rect 21616 4126 21717 4182
rect 21616 4092 21650 4126
rect 21684 4092 21717 4126
rect 21616 4036 21717 4092
rect 21616 4002 21650 4036
rect 21684 4002 21717 4036
rect 21616 3946 21717 4002
rect 21616 3912 21650 3946
rect 21684 3912 21717 3946
rect 21616 3856 21717 3912
rect 22803 4812 22837 4846
rect 22871 4812 22904 4846
rect 22803 4756 22904 4812
rect 22803 4722 22837 4756
rect 22871 4722 22904 4756
rect 22803 4666 22904 4722
rect 22803 4632 22837 4666
rect 22871 4632 22904 4666
rect 22803 4576 22904 4632
rect 22803 4542 22837 4576
rect 22871 4542 22904 4576
rect 22803 4486 22904 4542
rect 22803 4452 22837 4486
rect 22871 4452 22904 4486
rect 22803 4396 22904 4452
rect 22803 4362 22837 4396
rect 22871 4362 22904 4396
rect 22803 4306 22904 4362
rect 22803 4272 22837 4306
rect 22871 4272 22904 4306
rect 22803 4216 22904 4272
rect 22803 4182 22837 4216
rect 22871 4182 22904 4216
rect 22803 4126 22904 4182
rect 22803 4092 22837 4126
rect 22871 4092 22904 4126
rect 22803 4036 22904 4092
rect 22803 4002 22837 4036
rect 22871 4002 22904 4036
rect 22803 3946 22904 4002
rect 22803 3912 22837 3946
rect 22871 3912 22904 3946
rect 21616 3822 21650 3856
rect 21684 3822 21717 3856
rect 21616 3807 21717 3822
rect 22803 3856 22904 3912
rect 22803 3822 22837 3856
rect 22871 3822 22904 3856
rect 22803 3807 22904 3822
rect 21616 3772 22904 3807
rect 21616 3738 21746 3772
rect 21780 3738 21836 3772
rect 21870 3738 21926 3772
rect 21960 3738 22016 3772
rect 22050 3738 22106 3772
rect 22140 3738 22196 3772
rect 22230 3738 22286 3772
rect 22320 3738 22376 3772
rect 22410 3738 22466 3772
rect 22500 3738 22556 3772
rect 22590 3738 22646 3772
rect 22680 3738 22736 3772
rect 22770 3738 22904 3772
rect 21616 3706 22904 3738
rect 22976 4959 24264 4994
rect 22976 4936 23106 4959
rect 22976 4902 23010 4936
rect 23044 4925 23106 4936
rect 23140 4925 23196 4959
rect 23230 4925 23286 4959
rect 23320 4925 23376 4959
rect 23410 4925 23466 4959
rect 23500 4925 23556 4959
rect 23590 4925 23646 4959
rect 23680 4925 23736 4959
rect 23770 4925 23826 4959
rect 23860 4925 23916 4959
rect 23950 4925 24006 4959
rect 24040 4925 24096 4959
rect 24130 4936 24264 4959
rect 24130 4925 24197 4936
rect 23044 4902 24197 4925
rect 24231 4902 24264 4936
rect 22976 4893 24264 4902
rect 22976 4846 23077 4893
rect 22976 4812 23010 4846
rect 23044 4812 23077 4846
rect 24163 4846 24264 4893
rect 22976 4756 23077 4812
rect 22976 4722 23010 4756
rect 23044 4722 23077 4756
rect 22976 4666 23077 4722
rect 22976 4632 23010 4666
rect 23044 4632 23077 4666
rect 22976 4576 23077 4632
rect 22976 4542 23010 4576
rect 23044 4542 23077 4576
rect 22976 4486 23077 4542
rect 22976 4452 23010 4486
rect 23044 4452 23077 4486
rect 22976 4396 23077 4452
rect 22976 4362 23010 4396
rect 23044 4362 23077 4396
rect 22976 4306 23077 4362
rect 22976 4272 23010 4306
rect 23044 4272 23077 4306
rect 22976 4216 23077 4272
rect 22976 4182 23010 4216
rect 23044 4182 23077 4216
rect 22976 4126 23077 4182
rect 22976 4092 23010 4126
rect 23044 4092 23077 4126
rect 22976 4036 23077 4092
rect 22976 4002 23010 4036
rect 23044 4002 23077 4036
rect 22976 3946 23077 4002
rect 22976 3912 23010 3946
rect 23044 3912 23077 3946
rect 22976 3856 23077 3912
rect 24163 4812 24197 4846
rect 24231 4812 24264 4846
rect 24163 4756 24264 4812
rect 24163 4722 24197 4756
rect 24231 4722 24264 4756
rect 24163 4666 24264 4722
rect 24163 4632 24197 4666
rect 24231 4632 24264 4666
rect 24163 4576 24264 4632
rect 24163 4542 24197 4576
rect 24231 4542 24264 4576
rect 24163 4486 24264 4542
rect 24163 4452 24197 4486
rect 24231 4452 24264 4486
rect 24163 4396 24264 4452
rect 24163 4362 24197 4396
rect 24231 4362 24264 4396
rect 24163 4306 24264 4362
rect 24163 4272 24197 4306
rect 24231 4272 24264 4306
rect 24163 4216 24264 4272
rect 24163 4182 24197 4216
rect 24231 4182 24264 4216
rect 24163 4126 24264 4182
rect 24163 4092 24197 4126
rect 24231 4092 24264 4126
rect 24163 4036 24264 4092
rect 24163 4002 24197 4036
rect 24231 4002 24264 4036
rect 24163 3946 24264 4002
rect 24163 3912 24197 3946
rect 24231 3912 24264 3946
rect 22976 3822 23010 3856
rect 23044 3822 23077 3856
rect 22976 3807 23077 3822
rect 24163 3856 24264 3912
rect 24163 3822 24197 3856
rect 24231 3822 24264 3856
rect 24163 3807 24264 3822
rect 22976 3772 24264 3807
rect 22976 3738 23106 3772
rect 23140 3738 23196 3772
rect 23230 3738 23286 3772
rect 23320 3738 23376 3772
rect 23410 3738 23466 3772
rect 23500 3738 23556 3772
rect 23590 3738 23646 3772
rect 23680 3738 23736 3772
rect 23770 3738 23826 3772
rect 23860 3738 23916 3772
rect 23950 3738 24006 3772
rect 24040 3738 24096 3772
rect 24130 3738 24264 3772
rect 22976 3706 24264 3738
rect 20256 3599 21544 3634
rect 20256 3576 20386 3599
rect 20256 3542 20290 3576
rect 20324 3565 20386 3576
rect 20420 3565 20476 3599
rect 20510 3565 20566 3599
rect 20600 3565 20656 3599
rect 20690 3565 20746 3599
rect 20780 3565 20836 3599
rect 20870 3565 20926 3599
rect 20960 3565 21016 3599
rect 21050 3565 21106 3599
rect 21140 3565 21196 3599
rect 21230 3565 21286 3599
rect 21320 3565 21376 3599
rect 21410 3576 21544 3599
rect 21410 3565 21477 3576
rect 20324 3542 21477 3565
rect 21511 3542 21544 3576
rect 20256 3533 21544 3542
rect 20256 3486 20357 3533
rect 20256 3452 20290 3486
rect 20324 3452 20357 3486
rect 21443 3486 21544 3533
rect 20256 3396 20357 3452
rect 20256 3362 20290 3396
rect 20324 3362 20357 3396
rect 20256 3306 20357 3362
rect 20256 3272 20290 3306
rect 20324 3272 20357 3306
rect 20256 3216 20357 3272
rect 20256 3182 20290 3216
rect 20324 3182 20357 3216
rect 20256 3126 20357 3182
rect 20256 3092 20290 3126
rect 20324 3092 20357 3126
rect 19900 3030 20200 3060
rect 19900 2990 19930 3030
rect 19970 2990 20030 3030
rect 20070 2990 20130 3030
rect 20170 2990 20200 3030
rect 19900 2960 20200 2990
rect 20256 3036 20357 3092
rect 20256 3002 20290 3036
rect 20324 3002 20357 3036
rect 20256 2946 20357 3002
rect 20256 2912 20290 2946
rect 20324 2912 20357 2946
rect 20256 2856 20357 2912
rect 20256 2822 20290 2856
rect 20324 2822 20357 2856
rect 20256 2766 20357 2822
rect 20256 2732 20290 2766
rect 20324 2732 20357 2766
rect 20256 2676 20357 2732
rect 20256 2642 20290 2676
rect 20324 2642 20357 2676
rect 20256 2586 20357 2642
rect 20256 2552 20290 2586
rect 20324 2552 20357 2586
rect 20256 2496 20357 2552
rect 21443 3452 21477 3486
rect 21511 3452 21544 3486
rect 21443 3396 21544 3452
rect 21443 3362 21477 3396
rect 21511 3362 21544 3396
rect 21443 3306 21544 3362
rect 21443 3272 21477 3306
rect 21511 3272 21544 3306
rect 21443 3216 21544 3272
rect 21443 3182 21477 3216
rect 21511 3182 21544 3216
rect 21443 3126 21544 3182
rect 21443 3092 21477 3126
rect 21511 3092 21544 3126
rect 21443 3036 21544 3092
rect 21443 3002 21477 3036
rect 21511 3002 21544 3036
rect 21443 2946 21544 3002
rect 21443 2912 21477 2946
rect 21511 2912 21544 2946
rect 21443 2856 21544 2912
rect 21443 2822 21477 2856
rect 21511 2822 21544 2856
rect 21443 2766 21544 2822
rect 21443 2732 21477 2766
rect 21511 2732 21544 2766
rect 21443 2676 21544 2732
rect 21443 2642 21477 2676
rect 21511 2642 21544 2676
rect 21443 2586 21544 2642
rect 21443 2552 21477 2586
rect 21511 2552 21544 2586
rect 20256 2462 20290 2496
rect 20324 2462 20357 2496
rect 20256 2447 20357 2462
rect 21443 2496 21544 2552
rect 21443 2462 21477 2496
rect 21511 2462 21544 2496
rect 21443 2447 21544 2462
rect 20256 2412 21544 2447
rect 20256 2378 20386 2412
rect 20420 2378 20476 2412
rect 20510 2378 20566 2412
rect 20600 2378 20656 2412
rect 20690 2378 20746 2412
rect 20780 2378 20836 2412
rect 20870 2378 20926 2412
rect 20960 2378 21016 2412
rect 21050 2378 21106 2412
rect 21140 2378 21196 2412
rect 21230 2378 21286 2412
rect 21320 2378 21376 2412
rect 21410 2378 21544 2412
rect 20256 2346 21544 2378
rect 21616 3599 22904 3634
rect 21616 3576 21746 3599
rect 21616 3542 21650 3576
rect 21684 3565 21746 3576
rect 21780 3565 21836 3599
rect 21870 3565 21926 3599
rect 21960 3565 22016 3599
rect 22050 3565 22106 3599
rect 22140 3565 22196 3599
rect 22230 3565 22286 3599
rect 22320 3565 22376 3599
rect 22410 3565 22466 3599
rect 22500 3565 22556 3599
rect 22590 3565 22646 3599
rect 22680 3565 22736 3599
rect 22770 3576 22904 3599
rect 22770 3565 22837 3576
rect 21684 3542 22837 3565
rect 22871 3542 22904 3576
rect 21616 3533 22904 3542
rect 21616 3486 21717 3533
rect 21616 3452 21650 3486
rect 21684 3452 21717 3486
rect 22803 3486 22904 3533
rect 21616 3396 21717 3452
rect 21616 3362 21650 3396
rect 21684 3362 21717 3396
rect 21616 3306 21717 3362
rect 21616 3272 21650 3306
rect 21684 3272 21717 3306
rect 21616 3216 21717 3272
rect 21616 3182 21650 3216
rect 21684 3182 21717 3216
rect 21616 3126 21717 3182
rect 21616 3092 21650 3126
rect 21684 3092 21717 3126
rect 21616 3036 21717 3092
rect 21616 3002 21650 3036
rect 21684 3002 21717 3036
rect 21616 2946 21717 3002
rect 21616 2912 21650 2946
rect 21684 2912 21717 2946
rect 21616 2856 21717 2912
rect 21616 2822 21650 2856
rect 21684 2822 21717 2856
rect 21616 2766 21717 2822
rect 21616 2732 21650 2766
rect 21684 2732 21717 2766
rect 21616 2676 21717 2732
rect 21616 2642 21650 2676
rect 21684 2642 21717 2676
rect 21616 2586 21717 2642
rect 21616 2552 21650 2586
rect 21684 2552 21717 2586
rect 21616 2496 21717 2552
rect 22803 3452 22837 3486
rect 22871 3452 22904 3486
rect 22803 3396 22904 3452
rect 22803 3362 22837 3396
rect 22871 3362 22904 3396
rect 22803 3306 22904 3362
rect 22803 3272 22837 3306
rect 22871 3272 22904 3306
rect 22803 3216 22904 3272
rect 22803 3182 22837 3216
rect 22871 3182 22904 3216
rect 22803 3126 22904 3182
rect 22803 3092 22837 3126
rect 22871 3092 22904 3126
rect 22803 3036 22904 3092
rect 22803 3002 22837 3036
rect 22871 3002 22904 3036
rect 22803 2946 22904 3002
rect 22803 2912 22837 2946
rect 22871 2912 22904 2946
rect 22803 2856 22904 2912
rect 22803 2822 22837 2856
rect 22871 2822 22904 2856
rect 22803 2766 22904 2822
rect 22803 2732 22837 2766
rect 22871 2732 22904 2766
rect 22803 2676 22904 2732
rect 22803 2642 22837 2676
rect 22871 2642 22904 2676
rect 22803 2586 22904 2642
rect 22803 2552 22837 2586
rect 22871 2552 22904 2586
rect 21616 2462 21650 2496
rect 21684 2462 21717 2496
rect 21616 2447 21717 2462
rect 22803 2496 22904 2552
rect 22803 2462 22837 2496
rect 22871 2462 22904 2496
rect 22803 2447 22904 2462
rect 21616 2412 22904 2447
rect 21616 2378 21746 2412
rect 21780 2378 21836 2412
rect 21870 2378 21926 2412
rect 21960 2378 22016 2412
rect 22050 2378 22106 2412
rect 22140 2378 22196 2412
rect 22230 2378 22286 2412
rect 22320 2378 22376 2412
rect 22410 2378 22466 2412
rect 22500 2378 22556 2412
rect 22590 2378 22646 2412
rect 22680 2378 22736 2412
rect 22770 2378 22904 2412
rect 21616 2346 22904 2378
rect 22976 3599 24264 3634
rect 22976 3576 23106 3599
rect 22976 3542 23010 3576
rect 23044 3565 23106 3576
rect 23140 3565 23196 3599
rect 23230 3565 23286 3599
rect 23320 3565 23376 3599
rect 23410 3565 23466 3599
rect 23500 3565 23556 3599
rect 23590 3565 23646 3599
rect 23680 3565 23736 3599
rect 23770 3565 23826 3599
rect 23860 3565 23916 3599
rect 23950 3565 24006 3599
rect 24040 3565 24096 3599
rect 24130 3576 24264 3599
rect 24130 3565 24197 3576
rect 23044 3542 24197 3565
rect 24231 3542 24264 3576
rect 22976 3533 24264 3542
rect 22976 3486 23077 3533
rect 22976 3452 23010 3486
rect 23044 3452 23077 3486
rect 24163 3486 24264 3533
rect 22976 3396 23077 3452
rect 22976 3362 23010 3396
rect 23044 3362 23077 3396
rect 22976 3306 23077 3362
rect 22976 3272 23010 3306
rect 23044 3272 23077 3306
rect 22976 3216 23077 3272
rect 22976 3182 23010 3216
rect 23044 3182 23077 3216
rect 22976 3126 23077 3182
rect 22976 3092 23010 3126
rect 23044 3092 23077 3126
rect 22976 3036 23077 3092
rect 22976 3002 23010 3036
rect 23044 3002 23077 3036
rect 22976 2946 23077 3002
rect 22976 2912 23010 2946
rect 23044 2912 23077 2946
rect 22976 2856 23077 2912
rect 22976 2822 23010 2856
rect 23044 2822 23077 2856
rect 22976 2766 23077 2822
rect 22976 2732 23010 2766
rect 23044 2732 23077 2766
rect 22976 2676 23077 2732
rect 22976 2642 23010 2676
rect 23044 2642 23077 2676
rect 22976 2586 23077 2642
rect 22976 2552 23010 2586
rect 23044 2552 23077 2586
rect 22976 2496 23077 2552
rect 24163 3452 24197 3486
rect 24231 3452 24264 3486
rect 24163 3396 24264 3452
rect 24163 3362 24197 3396
rect 24231 3362 24264 3396
rect 24163 3306 24264 3362
rect 24163 3272 24197 3306
rect 24231 3272 24264 3306
rect 24163 3216 24264 3272
rect 24163 3182 24197 3216
rect 24231 3182 24264 3216
rect 24163 3126 24264 3182
rect 24163 3092 24197 3126
rect 24231 3092 24264 3126
rect 24163 3036 24264 3092
rect 24163 3002 24197 3036
rect 24231 3002 24264 3036
rect 24163 2946 24264 3002
rect 26170 3490 26830 3530
rect 26990 3490 27650 3530
rect 26170 3280 26210 3490
rect 27610 3280 27650 3490
rect 26170 3000 26210 3120
rect 27610 3000 27650 3120
rect 26170 2960 26830 3000
rect 26990 2960 27650 3000
rect 28690 3490 29350 3530
rect 29510 3490 30170 3530
rect 28690 3280 28730 3490
rect 30130 3280 30170 3490
rect 28690 3000 28730 3120
rect 30130 3000 30170 3120
rect 28690 2960 30170 3000
rect 24163 2912 24197 2946
rect 24231 2912 24264 2946
rect 24163 2856 24264 2912
rect 24163 2822 24197 2856
rect 24231 2822 24264 2856
rect 24163 2766 24264 2822
rect 24163 2732 24197 2766
rect 24231 2732 24264 2766
rect 24163 2676 24264 2732
rect 24163 2642 24197 2676
rect 24231 2642 24264 2676
rect 24163 2586 24264 2642
rect 24163 2552 24197 2586
rect 24231 2552 24264 2586
rect 22976 2462 23010 2496
rect 23044 2462 23077 2496
rect 22976 2447 23077 2462
rect 24163 2496 24264 2552
rect 24163 2462 24197 2496
rect 24231 2462 24264 2496
rect 24163 2447 24264 2462
rect 22976 2412 24264 2447
rect 22976 2378 23106 2412
rect 23140 2378 23196 2412
rect 23230 2378 23286 2412
rect 23320 2378 23376 2412
rect 23410 2378 23466 2412
rect 23500 2378 23556 2412
rect 23590 2378 23646 2412
rect 23680 2378 23736 2412
rect 23770 2378 23826 2412
rect 23860 2378 23916 2412
rect 23950 2378 24006 2412
rect 24040 2378 24096 2412
rect 24130 2378 24264 2412
rect 22976 2346 24264 2378
rect 25690 2840 26830 2880
rect 26990 2840 28130 2880
rect 25690 2530 25730 2840
rect 20256 2239 21544 2274
rect 20256 2216 20386 2239
rect 20256 2182 20290 2216
rect 20324 2205 20386 2216
rect 20420 2205 20476 2239
rect 20510 2205 20566 2239
rect 20600 2205 20656 2239
rect 20690 2205 20746 2239
rect 20780 2205 20836 2239
rect 20870 2205 20926 2239
rect 20960 2205 21016 2239
rect 21050 2205 21106 2239
rect 21140 2205 21196 2239
rect 21230 2205 21286 2239
rect 21320 2205 21376 2239
rect 21410 2216 21544 2239
rect 21410 2205 21477 2216
rect 20324 2182 21477 2205
rect 21511 2182 21544 2216
rect 20256 2173 21544 2182
rect 20256 2126 20357 2173
rect 20256 2092 20290 2126
rect 20324 2092 20357 2126
rect 21443 2126 21544 2173
rect 20256 2036 20357 2092
rect 20256 2002 20290 2036
rect 20324 2002 20357 2036
rect 20256 1946 20357 2002
rect 20256 1912 20290 1946
rect 20324 1912 20357 1946
rect 20256 1856 20357 1912
rect 20256 1822 20290 1856
rect 20324 1822 20357 1856
rect 20256 1766 20357 1822
rect 20256 1732 20290 1766
rect 20324 1732 20357 1766
rect 20256 1676 20357 1732
rect 20256 1642 20290 1676
rect 20324 1642 20357 1676
rect 20256 1586 20357 1642
rect 20256 1552 20290 1586
rect 20324 1552 20357 1586
rect 20256 1496 20357 1552
rect 20256 1462 20290 1496
rect 20324 1462 20357 1496
rect 20256 1406 20357 1462
rect 20256 1372 20290 1406
rect 20324 1372 20357 1406
rect 20256 1316 20357 1372
rect 20256 1282 20290 1316
rect 20324 1282 20357 1316
rect 20256 1226 20357 1282
rect 20256 1192 20290 1226
rect 20324 1192 20357 1226
rect 20256 1136 20357 1192
rect 21443 2092 21477 2126
rect 21511 2092 21544 2126
rect 21443 2036 21544 2092
rect 21443 2002 21477 2036
rect 21511 2002 21544 2036
rect 21443 1946 21544 2002
rect 21443 1912 21477 1946
rect 21511 1912 21544 1946
rect 21443 1856 21544 1912
rect 21443 1822 21477 1856
rect 21511 1822 21544 1856
rect 21443 1766 21544 1822
rect 21443 1732 21477 1766
rect 21511 1732 21544 1766
rect 21443 1676 21544 1732
rect 21443 1642 21477 1676
rect 21511 1642 21544 1676
rect 21443 1586 21544 1642
rect 21443 1552 21477 1586
rect 21511 1552 21544 1586
rect 21443 1496 21544 1552
rect 21443 1462 21477 1496
rect 21511 1462 21544 1496
rect 21443 1406 21544 1462
rect 21443 1372 21477 1406
rect 21511 1372 21544 1406
rect 21443 1316 21544 1372
rect 21443 1282 21477 1316
rect 21511 1282 21544 1316
rect 21443 1226 21544 1282
rect 21443 1192 21477 1226
rect 21511 1192 21544 1226
rect 20256 1102 20290 1136
rect 20324 1102 20357 1136
rect 20256 1087 20357 1102
rect 21443 1136 21544 1192
rect 21443 1102 21477 1136
rect 21511 1102 21544 1136
rect 21443 1087 21544 1102
rect 20256 1052 21544 1087
rect 20256 1018 20386 1052
rect 20420 1018 20476 1052
rect 20510 1018 20566 1052
rect 20600 1018 20656 1052
rect 20690 1018 20746 1052
rect 20780 1018 20836 1052
rect 20870 1018 20926 1052
rect 20960 1018 21016 1052
rect 21050 1018 21106 1052
rect 21140 1018 21196 1052
rect 21230 1018 21286 1052
rect 21320 1018 21376 1052
rect 21410 1018 21544 1052
rect 20256 986 21544 1018
rect 21616 2239 22904 2274
rect 21616 2216 21746 2239
rect 21616 2182 21650 2216
rect 21684 2205 21746 2216
rect 21780 2205 21836 2239
rect 21870 2205 21926 2239
rect 21960 2205 22016 2239
rect 22050 2205 22106 2239
rect 22140 2205 22196 2239
rect 22230 2205 22286 2239
rect 22320 2205 22376 2239
rect 22410 2205 22466 2239
rect 22500 2205 22556 2239
rect 22590 2205 22646 2239
rect 22680 2205 22736 2239
rect 22770 2216 22904 2239
rect 22770 2205 22837 2216
rect 21684 2182 22837 2205
rect 22871 2182 22904 2216
rect 21616 2173 22904 2182
rect 21616 2126 21717 2173
rect 21616 2092 21650 2126
rect 21684 2092 21717 2126
rect 22803 2126 22904 2173
rect 21616 2036 21717 2092
rect 21616 2002 21650 2036
rect 21684 2002 21717 2036
rect 21616 1946 21717 2002
rect 21616 1912 21650 1946
rect 21684 1912 21717 1946
rect 21616 1856 21717 1912
rect 21616 1822 21650 1856
rect 21684 1822 21717 1856
rect 21616 1766 21717 1822
rect 21616 1732 21650 1766
rect 21684 1732 21717 1766
rect 21616 1676 21717 1732
rect 21616 1642 21650 1676
rect 21684 1642 21717 1676
rect 21616 1586 21717 1642
rect 21616 1552 21650 1586
rect 21684 1552 21717 1586
rect 21616 1496 21717 1552
rect 21616 1462 21650 1496
rect 21684 1462 21717 1496
rect 21616 1406 21717 1462
rect 21616 1372 21650 1406
rect 21684 1372 21717 1406
rect 21616 1316 21717 1372
rect 21616 1282 21650 1316
rect 21684 1282 21717 1316
rect 21616 1226 21717 1282
rect 21616 1192 21650 1226
rect 21684 1192 21717 1226
rect 21616 1136 21717 1192
rect 22803 2092 22837 2126
rect 22871 2092 22904 2126
rect 22803 2036 22904 2092
rect 22803 2002 22837 2036
rect 22871 2002 22904 2036
rect 22803 1946 22904 2002
rect 22803 1912 22837 1946
rect 22871 1912 22904 1946
rect 22803 1856 22904 1912
rect 22803 1822 22837 1856
rect 22871 1822 22904 1856
rect 22803 1766 22904 1822
rect 22803 1732 22837 1766
rect 22871 1732 22904 1766
rect 22803 1676 22904 1732
rect 22803 1642 22837 1676
rect 22871 1642 22904 1676
rect 22803 1586 22904 1642
rect 22803 1552 22837 1586
rect 22871 1552 22904 1586
rect 22803 1496 22904 1552
rect 22803 1462 22837 1496
rect 22871 1462 22904 1496
rect 22803 1406 22904 1462
rect 22803 1372 22837 1406
rect 22871 1372 22904 1406
rect 22803 1316 22904 1372
rect 22803 1282 22837 1316
rect 22871 1282 22904 1316
rect 22803 1226 22904 1282
rect 22803 1192 22837 1226
rect 22871 1192 22904 1226
rect 21616 1102 21650 1136
rect 21684 1102 21717 1136
rect 21616 1087 21717 1102
rect 22803 1136 22904 1192
rect 22803 1102 22837 1136
rect 22871 1102 22904 1136
rect 22803 1087 22904 1102
rect 21616 1052 22904 1087
rect 21616 1018 21746 1052
rect 21780 1018 21836 1052
rect 21870 1018 21926 1052
rect 21960 1018 22016 1052
rect 22050 1018 22106 1052
rect 22140 1018 22196 1052
rect 22230 1018 22286 1052
rect 22320 1018 22376 1052
rect 22410 1018 22466 1052
rect 22500 1018 22556 1052
rect 22590 1018 22646 1052
rect 22680 1018 22736 1052
rect 22770 1018 22904 1052
rect 21616 986 22904 1018
rect 22976 2239 24264 2274
rect 22976 2216 23106 2239
rect 22976 2182 23010 2216
rect 23044 2205 23106 2216
rect 23140 2205 23196 2239
rect 23230 2205 23286 2239
rect 23320 2205 23376 2239
rect 23410 2205 23466 2239
rect 23500 2205 23556 2239
rect 23590 2205 23646 2239
rect 23680 2205 23736 2239
rect 23770 2205 23826 2239
rect 23860 2205 23916 2239
rect 23950 2205 24006 2239
rect 24040 2205 24096 2239
rect 24130 2216 24264 2239
rect 24130 2205 24197 2216
rect 23044 2182 24197 2205
rect 24231 2182 24264 2216
rect 22976 2173 24264 2182
rect 22976 2126 23077 2173
rect 22976 2092 23010 2126
rect 23044 2092 23077 2126
rect 24163 2126 24264 2173
rect 22976 2036 23077 2092
rect 22976 2002 23010 2036
rect 23044 2002 23077 2036
rect 22976 1946 23077 2002
rect 22976 1912 23010 1946
rect 23044 1912 23077 1946
rect 22976 1856 23077 1912
rect 22976 1822 23010 1856
rect 23044 1822 23077 1856
rect 22976 1766 23077 1822
rect 22976 1732 23010 1766
rect 23044 1732 23077 1766
rect 22976 1676 23077 1732
rect 22976 1642 23010 1676
rect 23044 1642 23077 1676
rect 22976 1586 23077 1642
rect 22976 1552 23010 1586
rect 23044 1552 23077 1586
rect 22976 1496 23077 1552
rect 22976 1462 23010 1496
rect 23044 1462 23077 1496
rect 22976 1406 23077 1462
rect 22976 1372 23010 1406
rect 23044 1372 23077 1406
rect 22976 1316 23077 1372
rect 22976 1282 23010 1316
rect 23044 1282 23077 1316
rect 22976 1226 23077 1282
rect 22976 1192 23010 1226
rect 23044 1192 23077 1226
rect 22976 1136 23077 1192
rect 24163 2092 24197 2126
rect 24231 2092 24264 2126
rect 24163 2036 24264 2092
rect 24163 2002 24197 2036
rect 24231 2002 24264 2036
rect 25690 2050 25730 2370
rect 28090 2530 28130 2840
rect 28090 2050 28130 2370
rect 25690 2010 26830 2050
rect 26990 2010 28130 2050
rect 28210 2840 29350 2880
rect 29510 2840 30650 2880
rect 28210 2530 28250 2840
rect 28210 2050 28250 2370
rect 30610 2530 30650 2840
rect 30610 2050 30650 2370
rect 28210 2010 29350 2050
rect 29510 2010 30650 2050
rect 24163 1946 24264 2002
rect 24163 1912 24197 1946
rect 24231 1912 24264 1946
rect 24163 1856 24264 1912
rect 24163 1822 24197 1856
rect 24231 1822 24264 1856
rect 24163 1766 24264 1822
rect 24163 1732 24197 1766
rect 24231 1732 24264 1766
rect 24163 1676 24264 1732
rect 24163 1642 24197 1676
rect 24231 1642 24264 1676
rect 24163 1586 24264 1642
rect 24163 1552 24197 1586
rect 24231 1552 24264 1586
rect 24163 1496 24264 1552
rect 24163 1462 24197 1496
rect 24231 1462 24264 1496
rect 24163 1406 24264 1462
rect 25890 1860 28090 1900
rect 28250 1860 30530 1900
rect 25890 1690 25930 1860
rect 25890 1450 25930 1530
rect 30290 1680 30370 1710
rect 30290 1640 30310 1680
rect 30350 1640 30370 1680
rect 30290 1580 30370 1640
rect 30290 1540 30310 1580
rect 30350 1540 30370 1580
rect 30290 1510 30370 1540
rect 30490 1690 30530 1860
rect 30490 1450 30530 1530
rect 25890 1410 28090 1450
rect 28250 1410 30530 1450
rect 24163 1372 24197 1406
rect 24231 1372 24264 1406
rect 24163 1316 24264 1372
rect 24163 1282 24197 1316
rect 24231 1282 24264 1316
rect 24163 1226 24264 1282
rect 24163 1192 24197 1226
rect 24231 1192 24264 1226
rect 22976 1102 23010 1136
rect 23044 1102 23077 1136
rect 22976 1087 23077 1102
rect 24163 1136 24264 1192
rect 24163 1102 24197 1136
rect 24231 1102 24264 1136
rect 24163 1087 24264 1102
rect 22976 1052 24264 1087
rect 22976 1018 23106 1052
rect 23140 1018 23196 1052
rect 23230 1018 23286 1052
rect 23320 1018 23376 1052
rect 23410 1018 23466 1052
rect 23500 1018 23556 1052
rect 23590 1018 23646 1052
rect 23680 1018 23736 1052
rect 23770 1018 23826 1052
rect 23860 1018 23916 1052
rect 23950 1018 24006 1052
rect 24040 1018 24096 1052
rect 24130 1018 24264 1052
rect 22976 986 24264 1018
rect 25290 1310 26070 1350
rect 26230 1310 27010 1350
rect 25290 1140 25330 1310
rect 25290 810 25330 980
rect 26970 1140 27010 1310
rect 26970 810 27010 980
rect 25290 770 26070 810
rect 26230 770 27010 810
rect 27130 1310 28090 1350
rect 28250 1310 29210 1350
rect 27130 1140 27170 1310
rect 27130 810 27170 980
rect 29170 1140 29210 1310
rect 29170 810 29210 980
rect 27130 770 28090 810
rect 28250 770 29210 810
rect 29290 1310 30070 1350
rect 30230 1310 31010 1350
rect 29290 1140 29330 1310
rect 29290 810 29330 980
rect 30970 1140 31010 1310
rect 30970 810 31010 980
rect 29290 770 30070 810
rect 30230 770 31010 810
<< nsubdiff >>
rect 25970 6400 30370 6440
rect 25970 5900 26010 6400
rect 26070 6220 26150 6250
rect 26070 6180 26090 6220
rect 26130 6180 26150 6220
rect 26070 6120 26150 6180
rect 26070 6080 26090 6120
rect 26130 6080 26150 6120
rect 26070 6050 26150 6080
rect 30190 6220 30270 6250
rect 30190 6180 30210 6220
rect 30250 6180 30270 6220
rect 30190 6120 30270 6180
rect 30190 6080 30210 6120
rect 30250 6080 30270 6120
rect 30190 6050 30270 6080
rect 30330 5900 30370 6400
rect 25970 5860 30370 5900
rect 26400 5480 29930 5520
rect 20419 4812 21381 4831
rect 20419 4778 20550 4812
rect 20584 4778 20640 4812
rect 20674 4778 20730 4812
rect 20764 4778 20820 4812
rect 20854 4778 20910 4812
rect 20944 4778 21000 4812
rect 21034 4778 21090 4812
rect 21124 4778 21180 4812
rect 21214 4778 21270 4812
rect 21304 4778 21381 4812
rect 20419 4759 21381 4778
rect 20419 4755 20491 4759
rect 20419 4721 20438 4755
rect 20472 4721 20491 4755
rect 20419 4665 20491 4721
rect 21309 4736 21381 4759
rect 21309 4702 21328 4736
rect 21362 4702 21381 4736
rect 20419 4631 20438 4665
rect 20472 4631 20491 4665
rect 20419 4575 20491 4631
rect 20419 4541 20438 4575
rect 20472 4541 20491 4575
rect 20419 4485 20491 4541
rect 20419 4451 20438 4485
rect 20472 4451 20491 4485
rect 20419 4395 20491 4451
rect 20419 4361 20438 4395
rect 20472 4361 20491 4395
rect 20419 4305 20491 4361
rect 20419 4271 20438 4305
rect 20472 4271 20491 4305
rect 20419 4215 20491 4271
rect 20419 4181 20438 4215
rect 20472 4181 20491 4215
rect 20419 4125 20491 4181
rect 20419 4091 20438 4125
rect 20472 4091 20491 4125
rect 20419 4035 20491 4091
rect 20419 4001 20438 4035
rect 20472 4001 20491 4035
rect 21309 4646 21381 4702
rect 21309 4612 21328 4646
rect 21362 4612 21381 4646
rect 21309 4556 21381 4612
rect 21309 4522 21328 4556
rect 21362 4522 21381 4556
rect 21309 4466 21381 4522
rect 21309 4432 21328 4466
rect 21362 4432 21381 4466
rect 21309 4376 21381 4432
rect 21309 4342 21328 4376
rect 21362 4342 21381 4376
rect 21309 4286 21381 4342
rect 21309 4252 21328 4286
rect 21362 4252 21381 4286
rect 21309 4196 21381 4252
rect 21309 4162 21328 4196
rect 21362 4162 21381 4196
rect 21309 4106 21381 4162
rect 21309 4072 21328 4106
rect 21362 4072 21381 4106
rect 21309 4016 21381 4072
rect 20419 3941 20491 4001
rect 21309 3982 21328 4016
rect 21362 3982 21381 4016
rect 21309 3941 21381 3982
rect 20419 3922 21381 3941
rect 20419 3888 20516 3922
rect 20550 3888 20606 3922
rect 20640 3888 20696 3922
rect 20730 3888 20786 3922
rect 20820 3888 20876 3922
rect 20910 3888 20966 3922
rect 21000 3888 21056 3922
rect 21090 3888 21146 3922
rect 21180 3888 21236 3922
rect 21270 3888 21381 3922
rect 20419 3869 21381 3888
rect 21779 4812 22741 4831
rect 21779 4778 21910 4812
rect 21944 4778 22000 4812
rect 22034 4778 22090 4812
rect 22124 4778 22180 4812
rect 22214 4778 22270 4812
rect 22304 4778 22360 4812
rect 22394 4778 22450 4812
rect 22484 4778 22540 4812
rect 22574 4778 22630 4812
rect 22664 4778 22741 4812
rect 21779 4759 22741 4778
rect 21779 4755 21851 4759
rect 21779 4721 21798 4755
rect 21832 4721 21851 4755
rect 21779 4665 21851 4721
rect 22669 4736 22741 4759
rect 22669 4702 22688 4736
rect 22722 4702 22741 4736
rect 21779 4631 21798 4665
rect 21832 4631 21851 4665
rect 21779 4575 21851 4631
rect 21779 4541 21798 4575
rect 21832 4541 21851 4575
rect 21779 4485 21851 4541
rect 21779 4451 21798 4485
rect 21832 4451 21851 4485
rect 21779 4395 21851 4451
rect 21779 4361 21798 4395
rect 21832 4361 21851 4395
rect 21779 4305 21851 4361
rect 21779 4271 21798 4305
rect 21832 4271 21851 4305
rect 21779 4215 21851 4271
rect 21779 4181 21798 4215
rect 21832 4181 21851 4215
rect 21779 4125 21851 4181
rect 21779 4091 21798 4125
rect 21832 4091 21851 4125
rect 21779 4035 21851 4091
rect 21779 4001 21798 4035
rect 21832 4001 21851 4035
rect 22669 4646 22741 4702
rect 22669 4612 22688 4646
rect 22722 4612 22741 4646
rect 22669 4556 22741 4612
rect 22669 4522 22688 4556
rect 22722 4522 22741 4556
rect 22669 4466 22741 4522
rect 22669 4432 22688 4466
rect 22722 4432 22741 4466
rect 22669 4376 22741 4432
rect 22669 4342 22688 4376
rect 22722 4342 22741 4376
rect 22669 4286 22741 4342
rect 22669 4252 22688 4286
rect 22722 4252 22741 4286
rect 22669 4196 22741 4252
rect 22669 4162 22688 4196
rect 22722 4162 22741 4196
rect 22669 4106 22741 4162
rect 22669 4072 22688 4106
rect 22722 4072 22741 4106
rect 22669 4016 22741 4072
rect 21779 3941 21851 4001
rect 22669 3982 22688 4016
rect 22722 3982 22741 4016
rect 22669 3941 22741 3982
rect 21779 3922 22741 3941
rect 21779 3888 21876 3922
rect 21910 3888 21966 3922
rect 22000 3888 22056 3922
rect 22090 3888 22146 3922
rect 22180 3888 22236 3922
rect 22270 3888 22326 3922
rect 22360 3888 22416 3922
rect 22450 3888 22506 3922
rect 22540 3888 22596 3922
rect 22630 3888 22741 3922
rect 21779 3869 22741 3888
rect 23139 4812 24101 4831
rect 23139 4778 23270 4812
rect 23304 4778 23360 4812
rect 23394 4778 23450 4812
rect 23484 4778 23540 4812
rect 23574 4778 23630 4812
rect 23664 4778 23720 4812
rect 23754 4778 23810 4812
rect 23844 4778 23900 4812
rect 23934 4778 23990 4812
rect 24024 4778 24101 4812
rect 23139 4759 24101 4778
rect 23139 4755 23211 4759
rect 23139 4721 23158 4755
rect 23192 4721 23211 4755
rect 23139 4665 23211 4721
rect 24029 4736 24101 4759
rect 24029 4702 24048 4736
rect 24082 4702 24101 4736
rect 23139 4631 23158 4665
rect 23192 4631 23211 4665
rect 23139 4575 23211 4631
rect 23139 4541 23158 4575
rect 23192 4541 23211 4575
rect 23139 4485 23211 4541
rect 23139 4451 23158 4485
rect 23192 4451 23211 4485
rect 23139 4395 23211 4451
rect 23139 4361 23158 4395
rect 23192 4361 23211 4395
rect 23139 4305 23211 4361
rect 23139 4271 23158 4305
rect 23192 4271 23211 4305
rect 23139 4215 23211 4271
rect 23139 4181 23158 4215
rect 23192 4181 23211 4215
rect 23139 4125 23211 4181
rect 23139 4091 23158 4125
rect 23192 4091 23211 4125
rect 23139 4035 23211 4091
rect 23139 4001 23158 4035
rect 23192 4001 23211 4035
rect 24029 4646 24101 4702
rect 24029 4612 24048 4646
rect 24082 4612 24101 4646
rect 24029 4556 24101 4612
rect 24029 4522 24048 4556
rect 24082 4522 24101 4556
rect 24029 4466 24101 4522
rect 24029 4432 24048 4466
rect 24082 4432 24101 4466
rect 24029 4376 24101 4432
rect 24029 4342 24048 4376
rect 24082 4342 24101 4376
rect 24029 4286 24101 4342
rect 24029 4252 24048 4286
rect 24082 4252 24101 4286
rect 24029 4196 24101 4252
rect 24029 4162 24048 4196
rect 24082 4162 24101 4196
rect 24029 4106 24101 4162
rect 24029 4072 24048 4106
rect 24082 4072 24101 4106
rect 24029 4016 24101 4072
rect 23139 3941 23211 4001
rect 24029 3982 24048 4016
rect 24082 3982 24101 4016
rect 24029 3941 24101 3982
rect 23139 3922 24101 3941
rect 23139 3888 23236 3922
rect 23270 3888 23326 3922
rect 23360 3888 23416 3922
rect 23450 3888 23506 3922
rect 23540 3888 23596 3922
rect 23630 3888 23686 3922
rect 23720 3888 23776 3922
rect 23810 3888 23866 3922
rect 23900 3888 23956 3922
rect 23990 3888 24101 3922
rect 23139 3869 24101 3888
rect 26400 4570 26440 5480
rect 29890 4570 29930 5480
rect 26400 4530 29930 4570
rect 25310 4150 26570 4190
rect 26730 4150 27990 4190
rect 25310 3980 25350 4150
rect 25310 3650 25350 3820
rect 27950 3980 27990 4150
rect 27950 3650 27990 3820
rect 20419 3452 21381 3471
rect 20419 3418 20550 3452
rect 20584 3418 20640 3452
rect 20674 3418 20730 3452
rect 20764 3418 20820 3452
rect 20854 3418 20910 3452
rect 20944 3418 21000 3452
rect 21034 3418 21090 3452
rect 21124 3418 21180 3452
rect 21214 3418 21270 3452
rect 21304 3418 21381 3452
rect 20419 3399 21381 3418
rect 20419 3395 20491 3399
rect 20419 3361 20438 3395
rect 20472 3361 20491 3395
rect 20419 3305 20491 3361
rect 21309 3376 21381 3399
rect 21309 3342 21328 3376
rect 21362 3342 21381 3376
rect 20419 3271 20438 3305
rect 20472 3271 20491 3305
rect 20419 3215 20491 3271
rect 20419 3181 20438 3215
rect 20472 3181 20491 3215
rect 20419 3125 20491 3181
rect 20419 3091 20438 3125
rect 20472 3091 20491 3125
rect 20419 3035 20491 3091
rect 20419 3001 20438 3035
rect 20472 3001 20491 3035
rect 20419 2945 20491 3001
rect 20419 2911 20438 2945
rect 20472 2911 20491 2945
rect 20419 2855 20491 2911
rect 20419 2821 20438 2855
rect 20472 2821 20491 2855
rect 20419 2765 20491 2821
rect 20419 2731 20438 2765
rect 20472 2731 20491 2765
rect 20419 2675 20491 2731
rect 20419 2641 20438 2675
rect 20472 2641 20491 2675
rect 21309 3286 21381 3342
rect 21309 3252 21328 3286
rect 21362 3252 21381 3286
rect 21309 3196 21381 3252
rect 21309 3162 21328 3196
rect 21362 3162 21381 3196
rect 21309 3106 21381 3162
rect 21309 3072 21328 3106
rect 21362 3072 21381 3106
rect 21309 3016 21381 3072
rect 21309 2982 21328 3016
rect 21362 2982 21381 3016
rect 21309 2926 21381 2982
rect 21309 2892 21328 2926
rect 21362 2892 21381 2926
rect 21309 2836 21381 2892
rect 21309 2802 21328 2836
rect 21362 2802 21381 2836
rect 21309 2746 21381 2802
rect 21309 2712 21328 2746
rect 21362 2712 21381 2746
rect 21309 2656 21381 2712
rect 20419 2581 20491 2641
rect 21309 2622 21328 2656
rect 21362 2622 21381 2656
rect 21309 2581 21381 2622
rect 20419 2562 21381 2581
rect 20419 2528 20516 2562
rect 20550 2528 20606 2562
rect 20640 2528 20696 2562
rect 20730 2528 20786 2562
rect 20820 2528 20876 2562
rect 20910 2528 20966 2562
rect 21000 2528 21056 2562
rect 21090 2528 21146 2562
rect 21180 2528 21236 2562
rect 21270 2528 21381 2562
rect 20419 2509 21381 2528
rect 21779 3452 22741 3471
rect 21779 3418 21910 3452
rect 21944 3418 22000 3452
rect 22034 3418 22090 3452
rect 22124 3418 22180 3452
rect 22214 3418 22270 3452
rect 22304 3418 22360 3452
rect 22394 3418 22450 3452
rect 22484 3418 22540 3452
rect 22574 3418 22630 3452
rect 22664 3418 22741 3452
rect 21779 3399 22741 3418
rect 21779 3395 21851 3399
rect 21779 3361 21798 3395
rect 21832 3361 21851 3395
rect 21779 3305 21851 3361
rect 22669 3376 22741 3399
rect 22669 3342 22688 3376
rect 22722 3342 22741 3376
rect 21779 3271 21798 3305
rect 21832 3271 21851 3305
rect 21779 3215 21851 3271
rect 21779 3181 21798 3215
rect 21832 3181 21851 3215
rect 21779 3125 21851 3181
rect 21779 3091 21798 3125
rect 21832 3091 21851 3125
rect 21779 3035 21851 3091
rect 21779 3001 21798 3035
rect 21832 3001 21851 3035
rect 21779 2945 21851 3001
rect 21779 2911 21798 2945
rect 21832 2911 21851 2945
rect 21779 2855 21851 2911
rect 21779 2821 21798 2855
rect 21832 2821 21851 2855
rect 21779 2765 21851 2821
rect 21779 2731 21798 2765
rect 21832 2731 21851 2765
rect 21779 2675 21851 2731
rect 21779 2641 21798 2675
rect 21832 2641 21851 2675
rect 22669 3286 22741 3342
rect 22669 3252 22688 3286
rect 22722 3252 22741 3286
rect 22669 3196 22741 3252
rect 22669 3162 22688 3196
rect 22722 3162 22741 3196
rect 22669 3106 22741 3162
rect 22669 3072 22688 3106
rect 22722 3072 22741 3106
rect 22669 3016 22741 3072
rect 22669 2982 22688 3016
rect 22722 2982 22741 3016
rect 22669 2926 22741 2982
rect 22669 2892 22688 2926
rect 22722 2892 22741 2926
rect 22669 2836 22741 2892
rect 22669 2802 22688 2836
rect 22722 2802 22741 2836
rect 22669 2746 22741 2802
rect 22669 2712 22688 2746
rect 22722 2712 22741 2746
rect 22669 2656 22741 2712
rect 21779 2581 21851 2641
rect 22669 2622 22688 2656
rect 22722 2622 22741 2656
rect 22669 2581 22741 2622
rect 21779 2562 22741 2581
rect 21779 2528 21876 2562
rect 21910 2528 21966 2562
rect 22000 2528 22056 2562
rect 22090 2528 22146 2562
rect 22180 2528 22236 2562
rect 22270 2528 22326 2562
rect 22360 2528 22416 2562
rect 22450 2528 22506 2562
rect 22540 2528 22596 2562
rect 22630 2528 22741 2562
rect 21779 2509 22741 2528
rect 25310 3610 26570 3650
rect 26730 3610 27990 3650
rect 28350 4150 29610 4190
rect 29770 4150 31030 4190
rect 28350 3980 28390 4150
rect 28350 3650 28390 3820
rect 30990 3980 31030 4150
rect 30990 3650 31030 3820
rect 28350 3610 29610 3650
rect 29770 3610 31030 3650
rect 23139 3452 24101 3471
rect 23139 3418 23270 3452
rect 23304 3418 23360 3452
rect 23394 3418 23450 3452
rect 23484 3418 23540 3452
rect 23574 3418 23630 3452
rect 23664 3418 23720 3452
rect 23754 3418 23810 3452
rect 23844 3418 23900 3452
rect 23934 3418 23990 3452
rect 24024 3418 24101 3452
rect 23139 3399 24101 3418
rect 23139 3395 23211 3399
rect 23139 3361 23158 3395
rect 23192 3361 23211 3395
rect 23139 3305 23211 3361
rect 24029 3376 24101 3399
rect 24029 3342 24048 3376
rect 24082 3342 24101 3376
rect 23139 3271 23158 3305
rect 23192 3271 23211 3305
rect 23139 3215 23211 3271
rect 23139 3181 23158 3215
rect 23192 3181 23211 3215
rect 23139 3125 23211 3181
rect 23139 3091 23158 3125
rect 23192 3091 23211 3125
rect 23139 3035 23211 3091
rect 23139 3001 23158 3035
rect 23192 3001 23211 3035
rect 23139 2945 23211 3001
rect 23139 2911 23158 2945
rect 23192 2911 23211 2945
rect 23139 2855 23211 2911
rect 23139 2821 23158 2855
rect 23192 2821 23211 2855
rect 23139 2765 23211 2821
rect 23139 2731 23158 2765
rect 23192 2731 23211 2765
rect 23139 2675 23211 2731
rect 23139 2641 23158 2675
rect 23192 2641 23211 2675
rect 24029 3286 24101 3342
rect 24029 3252 24048 3286
rect 24082 3252 24101 3286
rect 24029 3196 24101 3252
rect 24029 3162 24048 3196
rect 24082 3162 24101 3196
rect 24029 3106 24101 3162
rect 24029 3072 24048 3106
rect 24082 3072 24101 3106
rect 24029 3016 24101 3072
rect 24029 2982 24048 3016
rect 24082 2982 24101 3016
rect 24029 2926 24101 2982
rect 24029 2892 24048 2926
rect 24082 2892 24101 2926
rect 24029 2836 24101 2892
rect 24029 2802 24048 2836
rect 24082 2802 24101 2836
rect 24029 2746 24101 2802
rect 24029 2712 24048 2746
rect 24082 2712 24101 2746
rect 24029 2656 24101 2712
rect 23139 2581 23211 2641
rect 24029 2622 24048 2656
rect 24082 2622 24101 2656
rect 24029 2581 24101 2622
rect 23139 2562 24101 2581
rect 23139 2528 23236 2562
rect 23270 2528 23326 2562
rect 23360 2528 23416 2562
rect 23450 2528 23506 2562
rect 23540 2528 23596 2562
rect 23630 2528 23686 2562
rect 23720 2528 23776 2562
rect 23810 2528 23866 2562
rect 23900 2528 23956 2562
rect 23990 2528 24101 2562
rect 23139 2509 24101 2528
rect 20419 2092 21381 2111
rect 20419 2058 20550 2092
rect 20584 2058 20640 2092
rect 20674 2058 20730 2092
rect 20764 2058 20820 2092
rect 20854 2058 20910 2092
rect 20944 2058 21000 2092
rect 21034 2058 21090 2092
rect 21124 2058 21180 2092
rect 21214 2058 21270 2092
rect 21304 2058 21381 2092
rect 20419 2039 21381 2058
rect 20419 2035 20491 2039
rect 20419 2001 20438 2035
rect 20472 2001 20491 2035
rect 20419 1945 20491 2001
rect 21309 2016 21381 2039
rect 21309 1982 21328 2016
rect 21362 1982 21381 2016
rect 20419 1911 20438 1945
rect 20472 1911 20491 1945
rect 20419 1855 20491 1911
rect 20419 1821 20438 1855
rect 20472 1821 20491 1855
rect 20419 1765 20491 1821
rect 20419 1731 20438 1765
rect 20472 1731 20491 1765
rect 20419 1675 20491 1731
rect 20419 1641 20438 1675
rect 20472 1641 20491 1675
rect 20419 1585 20491 1641
rect 20419 1551 20438 1585
rect 20472 1551 20491 1585
rect 20419 1495 20491 1551
rect 20419 1461 20438 1495
rect 20472 1461 20491 1495
rect 20419 1405 20491 1461
rect 20419 1371 20438 1405
rect 20472 1371 20491 1405
rect 20419 1315 20491 1371
rect 20419 1281 20438 1315
rect 20472 1281 20491 1315
rect 21309 1926 21381 1982
rect 21309 1892 21328 1926
rect 21362 1892 21381 1926
rect 21309 1836 21381 1892
rect 21309 1802 21328 1836
rect 21362 1802 21381 1836
rect 21309 1746 21381 1802
rect 21309 1712 21328 1746
rect 21362 1712 21381 1746
rect 21309 1656 21381 1712
rect 21309 1622 21328 1656
rect 21362 1622 21381 1656
rect 21309 1566 21381 1622
rect 21309 1532 21328 1566
rect 21362 1532 21381 1566
rect 21309 1476 21381 1532
rect 21309 1442 21328 1476
rect 21362 1442 21381 1476
rect 21309 1386 21381 1442
rect 21309 1352 21328 1386
rect 21362 1352 21381 1386
rect 21309 1296 21381 1352
rect 20419 1221 20491 1281
rect 21309 1262 21328 1296
rect 21362 1262 21381 1296
rect 21309 1221 21381 1262
rect 20419 1202 21381 1221
rect 20419 1168 20516 1202
rect 20550 1168 20606 1202
rect 20640 1168 20696 1202
rect 20730 1168 20786 1202
rect 20820 1168 20876 1202
rect 20910 1168 20966 1202
rect 21000 1168 21056 1202
rect 21090 1168 21146 1202
rect 21180 1168 21236 1202
rect 21270 1168 21381 1202
rect 20419 1149 21381 1168
rect 21779 2092 22741 2111
rect 21779 2058 21910 2092
rect 21944 2058 22000 2092
rect 22034 2058 22090 2092
rect 22124 2058 22180 2092
rect 22214 2058 22270 2092
rect 22304 2058 22360 2092
rect 22394 2058 22450 2092
rect 22484 2058 22540 2092
rect 22574 2058 22630 2092
rect 22664 2058 22741 2092
rect 21779 2039 22741 2058
rect 21779 2035 21851 2039
rect 21779 2001 21798 2035
rect 21832 2001 21851 2035
rect 21779 1945 21851 2001
rect 22669 2016 22741 2039
rect 22669 1982 22688 2016
rect 22722 1982 22741 2016
rect 21779 1911 21798 1945
rect 21832 1911 21851 1945
rect 21779 1855 21851 1911
rect 21779 1821 21798 1855
rect 21832 1821 21851 1855
rect 21779 1765 21851 1821
rect 21779 1731 21798 1765
rect 21832 1731 21851 1765
rect 21779 1675 21851 1731
rect 21779 1641 21798 1675
rect 21832 1641 21851 1675
rect 21779 1585 21851 1641
rect 21779 1551 21798 1585
rect 21832 1551 21851 1585
rect 21779 1495 21851 1551
rect 21779 1461 21798 1495
rect 21832 1461 21851 1495
rect 21779 1405 21851 1461
rect 21779 1371 21798 1405
rect 21832 1371 21851 1405
rect 21779 1315 21851 1371
rect 21779 1281 21798 1315
rect 21832 1281 21851 1315
rect 22669 1926 22741 1982
rect 22669 1892 22688 1926
rect 22722 1892 22741 1926
rect 22669 1836 22741 1892
rect 22669 1802 22688 1836
rect 22722 1802 22741 1836
rect 22669 1746 22741 1802
rect 22669 1712 22688 1746
rect 22722 1712 22741 1746
rect 22669 1656 22741 1712
rect 22669 1622 22688 1656
rect 22722 1622 22741 1656
rect 22669 1566 22741 1622
rect 22669 1532 22688 1566
rect 22722 1532 22741 1566
rect 22669 1476 22741 1532
rect 22669 1442 22688 1476
rect 22722 1442 22741 1476
rect 22669 1386 22741 1442
rect 22669 1352 22688 1386
rect 22722 1352 22741 1386
rect 22669 1296 22741 1352
rect 21779 1221 21851 1281
rect 22669 1262 22688 1296
rect 22722 1262 22741 1296
rect 22669 1221 22741 1262
rect 21779 1202 22741 1221
rect 21779 1168 21876 1202
rect 21910 1168 21966 1202
rect 22000 1168 22056 1202
rect 22090 1168 22146 1202
rect 22180 1168 22236 1202
rect 22270 1168 22326 1202
rect 22360 1168 22416 1202
rect 22450 1168 22506 1202
rect 22540 1168 22596 1202
rect 22630 1168 22741 1202
rect 21779 1149 22741 1168
rect 23139 2092 24101 2111
rect 23139 2058 23270 2092
rect 23304 2058 23360 2092
rect 23394 2058 23450 2092
rect 23484 2058 23540 2092
rect 23574 2058 23630 2092
rect 23664 2058 23720 2092
rect 23754 2058 23810 2092
rect 23844 2058 23900 2092
rect 23934 2058 23990 2092
rect 24024 2058 24101 2092
rect 23139 2039 24101 2058
rect 23139 2035 23211 2039
rect 23139 2001 23158 2035
rect 23192 2001 23211 2035
rect 23139 1945 23211 2001
rect 24029 2016 24101 2039
rect 24029 1982 24048 2016
rect 24082 1982 24101 2016
rect 23139 1911 23158 1945
rect 23192 1911 23211 1945
rect 23139 1855 23211 1911
rect 23139 1821 23158 1855
rect 23192 1821 23211 1855
rect 23139 1765 23211 1821
rect 23139 1731 23158 1765
rect 23192 1731 23211 1765
rect 23139 1675 23211 1731
rect 23139 1641 23158 1675
rect 23192 1641 23211 1675
rect 23139 1585 23211 1641
rect 23139 1551 23158 1585
rect 23192 1551 23211 1585
rect 23139 1495 23211 1551
rect 23139 1461 23158 1495
rect 23192 1461 23211 1495
rect 23139 1405 23211 1461
rect 23139 1371 23158 1405
rect 23192 1371 23211 1405
rect 23139 1315 23211 1371
rect 23139 1281 23158 1315
rect 23192 1281 23211 1315
rect 24029 1926 24101 1982
rect 24029 1892 24048 1926
rect 24082 1892 24101 1926
rect 24029 1836 24101 1892
rect 24029 1802 24048 1836
rect 24082 1802 24101 1836
rect 24029 1746 24101 1802
rect 24029 1712 24048 1746
rect 24082 1712 24101 1746
rect 24029 1656 24101 1712
rect 24029 1622 24048 1656
rect 24082 1622 24101 1656
rect 24029 1566 24101 1622
rect 24029 1532 24048 1566
rect 24082 1532 24101 1566
rect 24029 1476 24101 1532
rect 24029 1442 24048 1476
rect 24082 1442 24101 1476
rect 24029 1386 24101 1442
rect 24029 1352 24048 1386
rect 24082 1352 24101 1386
rect 24029 1296 24101 1352
rect 23139 1221 23211 1281
rect 24029 1262 24048 1296
rect 24082 1262 24101 1296
rect 24029 1221 24101 1262
rect 23139 1202 24101 1221
rect 23139 1168 23236 1202
rect 23270 1168 23326 1202
rect 23360 1168 23416 1202
rect 23450 1168 23506 1202
rect 23540 1168 23596 1202
rect 23630 1168 23686 1202
rect 23720 1168 23776 1202
rect 23810 1168 23866 1202
rect 23900 1168 23956 1202
rect 23990 1168 24101 1202
rect 23139 1149 24101 1168
<< psubdiffcont >>
rect 21840 5760 21900 5820
rect 22000 5760 22060 5820
rect 22160 5760 22220 5820
rect 20290 4902 20324 4936
rect 20386 4925 20420 4959
rect 20476 4925 20510 4959
rect 20566 4925 20600 4959
rect 20656 4925 20690 4959
rect 20746 4925 20780 4959
rect 20836 4925 20870 4959
rect 20926 4925 20960 4959
rect 21016 4925 21050 4959
rect 21106 4925 21140 4959
rect 21196 4925 21230 4959
rect 21286 4925 21320 4959
rect 21376 4925 21410 4959
rect 21477 4902 21511 4936
rect 20290 4812 20324 4846
rect 20290 4722 20324 4756
rect 20290 4632 20324 4666
rect 20290 4542 20324 4576
rect 20290 4452 20324 4486
rect 20290 4362 20324 4396
rect 20290 4272 20324 4306
rect 20290 4182 20324 4216
rect 20290 4092 20324 4126
rect 20290 4002 20324 4036
rect 20290 3912 20324 3946
rect 21477 4812 21511 4846
rect 21477 4722 21511 4756
rect 21477 4632 21511 4666
rect 21477 4542 21511 4576
rect 21477 4452 21511 4486
rect 21477 4362 21511 4396
rect 21477 4272 21511 4306
rect 21477 4182 21511 4216
rect 21477 4092 21511 4126
rect 21477 4002 21511 4036
rect 21477 3912 21511 3946
rect 20290 3822 20324 3856
rect 21477 3822 21511 3856
rect 20386 3738 20420 3772
rect 20476 3738 20510 3772
rect 20566 3738 20600 3772
rect 20656 3738 20690 3772
rect 20746 3738 20780 3772
rect 20836 3738 20870 3772
rect 20926 3738 20960 3772
rect 21016 3738 21050 3772
rect 21106 3738 21140 3772
rect 21196 3738 21230 3772
rect 21286 3738 21320 3772
rect 21376 3738 21410 3772
rect 21650 4902 21684 4936
rect 21746 4925 21780 4959
rect 21836 4925 21870 4959
rect 21926 4925 21960 4959
rect 22016 4925 22050 4959
rect 22106 4925 22140 4959
rect 22196 4925 22230 4959
rect 22286 4925 22320 4959
rect 22376 4925 22410 4959
rect 22466 4925 22500 4959
rect 22556 4925 22590 4959
rect 22646 4925 22680 4959
rect 22736 4925 22770 4959
rect 22837 4902 22871 4936
rect 21650 4812 21684 4846
rect 21650 4722 21684 4756
rect 21650 4632 21684 4666
rect 21650 4542 21684 4576
rect 21650 4452 21684 4486
rect 21650 4362 21684 4396
rect 21650 4272 21684 4306
rect 21650 4182 21684 4216
rect 21650 4092 21684 4126
rect 21650 4002 21684 4036
rect 21650 3912 21684 3946
rect 22837 4812 22871 4846
rect 22837 4722 22871 4756
rect 22837 4632 22871 4666
rect 22837 4542 22871 4576
rect 22837 4452 22871 4486
rect 22837 4362 22871 4396
rect 22837 4272 22871 4306
rect 22837 4182 22871 4216
rect 22837 4092 22871 4126
rect 22837 4002 22871 4036
rect 22837 3912 22871 3946
rect 21650 3822 21684 3856
rect 22837 3822 22871 3856
rect 21746 3738 21780 3772
rect 21836 3738 21870 3772
rect 21926 3738 21960 3772
rect 22016 3738 22050 3772
rect 22106 3738 22140 3772
rect 22196 3738 22230 3772
rect 22286 3738 22320 3772
rect 22376 3738 22410 3772
rect 22466 3738 22500 3772
rect 22556 3738 22590 3772
rect 22646 3738 22680 3772
rect 22736 3738 22770 3772
rect 23010 4902 23044 4936
rect 23106 4925 23140 4959
rect 23196 4925 23230 4959
rect 23286 4925 23320 4959
rect 23376 4925 23410 4959
rect 23466 4925 23500 4959
rect 23556 4925 23590 4959
rect 23646 4925 23680 4959
rect 23736 4925 23770 4959
rect 23826 4925 23860 4959
rect 23916 4925 23950 4959
rect 24006 4925 24040 4959
rect 24096 4925 24130 4959
rect 24197 4902 24231 4936
rect 23010 4812 23044 4846
rect 23010 4722 23044 4756
rect 23010 4632 23044 4666
rect 23010 4542 23044 4576
rect 23010 4452 23044 4486
rect 23010 4362 23044 4396
rect 23010 4272 23044 4306
rect 23010 4182 23044 4216
rect 23010 4092 23044 4126
rect 23010 4002 23044 4036
rect 23010 3912 23044 3946
rect 24197 4812 24231 4846
rect 24197 4722 24231 4756
rect 24197 4632 24231 4666
rect 24197 4542 24231 4576
rect 24197 4452 24231 4486
rect 24197 4362 24231 4396
rect 24197 4272 24231 4306
rect 24197 4182 24231 4216
rect 24197 4092 24231 4126
rect 24197 4002 24231 4036
rect 24197 3912 24231 3946
rect 23010 3822 23044 3856
rect 24197 3822 24231 3856
rect 23106 3738 23140 3772
rect 23196 3738 23230 3772
rect 23286 3738 23320 3772
rect 23376 3738 23410 3772
rect 23466 3738 23500 3772
rect 23556 3738 23590 3772
rect 23646 3738 23680 3772
rect 23736 3738 23770 3772
rect 23826 3738 23860 3772
rect 23916 3738 23950 3772
rect 24006 3738 24040 3772
rect 24096 3738 24130 3772
rect 20290 3542 20324 3576
rect 20386 3565 20420 3599
rect 20476 3565 20510 3599
rect 20566 3565 20600 3599
rect 20656 3565 20690 3599
rect 20746 3565 20780 3599
rect 20836 3565 20870 3599
rect 20926 3565 20960 3599
rect 21016 3565 21050 3599
rect 21106 3565 21140 3599
rect 21196 3565 21230 3599
rect 21286 3565 21320 3599
rect 21376 3565 21410 3599
rect 21477 3542 21511 3576
rect 20290 3452 20324 3486
rect 20290 3362 20324 3396
rect 20290 3272 20324 3306
rect 20290 3182 20324 3216
rect 20290 3092 20324 3126
rect 19930 2990 19970 3030
rect 20030 2990 20070 3030
rect 20130 2990 20170 3030
rect 20290 3002 20324 3036
rect 20290 2912 20324 2946
rect 20290 2822 20324 2856
rect 20290 2732 20324 2766
rect 20290 2642 20324 2676
rect 20290 2552 20324 2586
rect 21477 3452 21511 3486
rect 21477 3362 21511 3396
rect 21477 3272 21511 3306
rect 21477 3182 21511 3216
rect 21477 3092 21511 3126
rect 21477 3002 21511 3036
rect 21477 2912 21511 2946
rect 21477 2822 21511 2856
rect 21477 2732 21511 2766
rect 21477 2642 21511 2676
rect 21477 2552 21511 2586
rect 20290 2462 20324 2496
rect 21477 2462 21511 2496
rect 20386 2378 20420 2412
rect 20476 2378 20510 2412
rect 20566 2378 20600 2412
rect 20656 2378 20690 2412
rect 20746 2378 20780 2412
rect 20836 2378 20870 2412
rect 20926 2378 20960 2412
rect 21016 2378 21050 2412
rect 21106 2378 21140 2412
rect 21196 2378 21230 2412
rect 21286 2378 21320 2412
rect 21376 2378 21410 2412
rect 21650 3542 21684 3576
rect 21746 3565 21780 3599
rect 21836 3565 21870 3599
rect 21926 3565 21960 3599
rect 22016 3565 22050 3599
rect 22106 3565 22140 3599
rect 22196 3565 22230 3599
rect 22286 3565 22320 3599
rect 22376 3565 22410 3599
rect 22466 3565 22500 3599
rect 22556 3565 22590 3599
rect 22646 3565 22680 3599
rect 22736 3565 22770 3599
rect 22837 3542 22871 3576
rect 21650 3452 21684 3486
rect 21650 3362 21684 3396
rect 21650 3272 21684 3306
rect 21650 3182 21684 3216
rect 21650 3092 21684 3126
rect 21650 3002 21684 3036
rect 21650 2912 21684 2946
rect 21650 2822 21684 2856
rect 21650 2732 21684 2766
rect 21650 2642 21684 2676
rect 21650 2552 21684 2586
rect 22837 3452 22871 3486
rect 22837 3362 22871 3396
rect 22837 3272 22871 3306
rect 22837 3182 22871 3216
rect 22837 3092 22871 3126
rect 22837 3002 22871 3036
rect 22837 2912 22871 2946
rect 22837 2822 22871 2856
rect 22837 2732 22871 2766
rect 22837 2642 22871 2676
rect 22837 2552 22871 2586
rect 21650 2462 21684 2496
rect 22837 2462 22871 2496
rect 21746 2378 21780 2412
rect 21836 2378 21870 2412
rect 21926 2378 21960 2412
rect 22016 2378 22050 2412
rect 22106 2378 22140 2412
rect 22196 2378 22230 2412
rect 22286 2378 22320 2412
rect 22376 2378 22410 2412
rect 22466 2378 22500 2412
rect 22556 2378 22590 2412
rect 22646 2378 22680 2412
rect 22736 2378 22770 2412
rect 23010 3542 23044 3576
rect 23106 3565 23140 3599
rect 23196 3565 23230 3599
rect 23286 3565 23320 3599
rect 23376 3565 23410 3599
rect 23466 3565 23500 3599
rect 23556 3565 23590 3599
rect 23646 3565 23680 3599
rect 23736 3565 23770 3599
rect 23826 3565 23860 3599
rect 23916 3565 23950 3599
rect 24006 3565 24040 3599
rect 24096 3565 24130 3599
rect 24197 3542 24231 3576
rect 23010 3452 23044 3486
rect 23010 3362 23044 3396
rect 23010 3272 23044 3306
rect 23010 3182 23044 3216
rect 23010 3092 23044 3126
rect 23010 3002 23044 3036
rect 23010 2912 23044 2946
rect 23010 2822 23044 2856
rect 23010 2732 23044 2766
rect 23010 2642 23044 2676
rect 23010 2552 23044 2586
rect 24197 3452 24231 3486
rect 24197 3362 24231 3396
rect 24197 3272 24231 3306
rect 24197 3182 24231 3216
rect 24197 3092 24231 3126
rect 24197 3002 24231 3036
rect 26830 3490 26990 3530
rect 26170 3120 26210 3280
rect 27610 3120 27650 3280
rect 26830 2960 26990 3000
rect 29350 3490 29510 3530
rect 28690 3120 28730 3280
rect 30130 3120 30170 3280
rect 24197 2912 24231 2946
rect 24197 2822 24231 2856
rect 24197 2732 24231 2766
rect 24197 2642 24231 2676
rect 24197 2552 24231 2586
rect 23010 2462 23044 2496
rect 24197 2462 24231 2496
rect 23106 2378 23140 2412
rect 23196 2378 23230 2412
rect 23286 2378 23320 2412
rect 23376 2378 23410 2412
rect 23466 2378 23500 2412
rect 23556 2378 23590 2412
rect 23646 2378 23680 2412
rect 23736 2378 23770 2412
rect 23826 2378 23860 2412
rect 23916 2378 23950 2412
rect 24006 2378 24040 2412
rect 24096 2378 24130 2412
rect 26830 2840 26990 2880
rect 25690 2370 25730 2530
rect 20290 2182 20324 2216
rect 20386 2205 20420 2239
rect 20476 2205 20510 2239
rect 20566 2205 20600 2239
rect 20656 2205 20690 2239
rect 20746 2205 20780 2239
rect 20836 2205 20870 2239
rect 20926 2205 20960 2239
rect 21016 2205 21050 2239
rect 21106 2205 21140 2239
rect 21196 2205 21230 2239
rect 21286 2205 21320 2239
rect 21376 2205 21410 2239
rect 21477 2182 21511 2216
rect 20290 2092 20324 2126
rect 20290 2002 20324 2036
rect 20290 1912 20324 1946
rect 20290 1822 20324 1856
rect 20290 1732 20324 1766
rect 20290 1642 20324 1676
rect 20290 1552 20324 1586
rect 20290 1462 20324 1496
rect 20290 1372 20324 1406
rect 20290 1282 20324 1316
rect 20290 1192 20324 1226
rect 21477 2092 21511 2126
rect 21477 2002 21511 2036
rect 21477 1912 21511 1946
rect 21477 1822 21511 1856
rect 21477 1732 21511 1766
rect 21477 1642 21511 1676
rect 21477 1552 21511 1586
rect 21477 1462 21511 1496
rect 21477 1372 21511 1406
rect 21477 1282 21511 1316
rect 21477 1192 21511 1226
rect 20290 1102 20324 1136
rect 21477 1102 21511 1136
rect 20386 1018 20420 1052
rect 20476 1018 20510 1052
rect 20566 1018 20600 1052
rect 20656 1018 20690 1052
rect 20746 1018 20780 1052
rect 20836 1018 20870 1052
rect 20926 1018 20960 1052
rect 21016 1018 21050 1052
rect 21106 1018 21140 1052
rect 21196 1018 21230 1052
rect 21286 1018 21320 1052
rect 21376 1018 21410 1052
rect 21650 2182 21684 2216
rect 21746 2205 21780 2239
rect 21836 2205 21870 2239
rect 21926 2205 21960 2239
rect 22016 2205 22050 2239
rect 22106 2205 22140 2239
rect 22196 2205 22230 2239
rect 22286 2205 22320 2239
rect 22376 2205 22410 2239
rect 22466 2205 22500 2239
rect 22556 2205 22590 2239
rect 22646 2205 22680 2239
rect 22736 2205 22770 2239
rect 22837 2182 22871 2216
rect 21650 2092 21684 2126
rect 21650 2002 21684 2036
rect 21650 1912 21684 1946
rect 21650 1822 21684 1856
rect 21650 1732 21684 1766
rect 21650 1642 21684 1676
rect 21650 1552 21684 1586
rect 21650 1462 21684 1496
rect 21650 1372 21684 1406
rect 21650 1282 21684 1316
rect 21650 1192 21684 1226
rect 22837 2092 22871 2126
rect 22837 2002 22871 2036
rect 22837 1912 22871 1946
rect 22837 1822 22871 1856
rect 22837 1732 22871 1766
rect 22837 1642 22871 1676
rect 22837 1552 22871 1586
rect 22837 1462 22871 1496
rect 22837 1372 22871 1406
rect 22837 1282 22871 1316
rect 22837 1192 22871 1226
rect 21650 1102 21684 1136
rect 22837 1102 22871 1136
rect 21746 1018 21780 1052
rect 21836 1018 21870 1052
rect 21926 1018 21960 1052
rect 22016 1018 22050 1052
rect 22106 1018 22140 1052
rect 22196 1018 22230 1052
rect 22286 1018 22320 1052
rect 22376 1018 22410 1052
rect 22466 1018 22500 1052
rect 22556 1018 22590 1052
rect 22646 1018 22680 1052
rect 22736 1018 22770 1052
rect 23010 2182 23044 2216
rect 23106 2205 23140 2239
rect 23196 2205 23230 2239
rect 23286 2205 23320 2239
rect 23376 2205 23410 2239
rect 23466 2205 23500 2239
rect 23556 2205 23590 2239
rect 23646 2205 23680 2239
rect 23736 2205 23770 2239
rect 23826 2205 23860 2239
rect 23916 2205 23950 2239
rect 24006 2205 24040 2239
rect 24096 2205 24130 2239
rect 24197 2182 24231 2216
rect 23010 2092 23044 2126
rect 23010 2002 23044 2036
rect 23010 1912 23044 1946
rect 23010 1822 23044 1856
rect 23010 1732 23044 1766
rect 23010 1642 23044 1676
rect 23010 1552 23044 1586
rect 23010 1462 23044 1496
rect 23010 1372 23044 1406
rect 23010 1282 23044 1316
rect 23010 1192 23044 1226
rect 24197 2092 24231 2126
rect 24197 2002 24231 2036
rect 28090 2370 28130 2530
rect 26830 2010 26990 2050
rect 29350 2840 29510 2880
rect 28210 2370 28250 2530
rect 30610 2370 30650 2530
rect 29350 2010 29510 2050
rect 24197 1912 24231 1946
rect 24197 1822 24231 1856
rect 24197 1732 24231 1766
rect 24197 1642 24231 1676
rect 24197 1552 24231 1586
rect 24197 1462 24231 1496
rect 28090 1860 28250 1900
rect 25890 1530 25930 1690
rect 30310 1640 30350 1680
rect 30310 1540 30350 1580
rect 30490 1530 30530 1690
rect 28090 1410 28250 1450
rect 24197 1372 24231 1406
rect 24197 1282 24231 1316
rect 24197 1192 24231 1226
rect 23010 1102 23044 1136
rect 24197 1102 24231 1136
rect 23106 1018 23140 1052
rect 23196 1018 23230 1052
rect 23286 1018 23320 1052
rect 23376 1018 23410 1052
rect 23466 1018 23500 1052
rect 23556 1018 23590 1052
rect 23646 1018 23680 1052
rect 23736 1018 23770 1052
rect 23826 1018 23860 1052
rect 23916 1018 23950 1052
rect 24006 1018 24040 1052
rect 24096 1018 24130 1052
rect 26070 1310 26230 1350
rect 25290 980 25330 1140
rect 26970 980 27010 1140
rect 26070 770 26230 810
rect 28090 1310 28250 1350
rect 27130 980 27170 1140
rect 29170 980 29210 1140
rect 28090 770 28250 810
rect 30070 1310 30230 1350
rect 29290 980 29330 1140
rect 30970 980 31010 1140
rect 30070 770 30230 810
<< nsubdiffcont >>
rect 26090 6180 26130 6220
rect 26090 6080 26130 6120
rect 30210 6180 30250 6220
rect 30210 6080 30250 6120
rect 20550 4778 20584 4812
rect 20640 4778 20674 4812
rect 20730 4778 20764 4812
rect 20820 4778 20854 4812
rect 20910 4778 20944 4812
rect 21000 4778 21034 4812
rect 21090 4778 21124 4812
rect 21180 4778 21214 4812
rect 21270 4778 21304 4812
rect 20438 4721 20472 4755
rect 21328 4702 21362 4736
rect 20438 4631 20472 4665
rect 20438 4541 20472 4575
rect 20438 4451 20472 4485
rect 20438 4361 20472 4395
rect 20438 4271 20472 4305
rect 20438 4181 20472 4215
rect 20438 4091 20472 4125
rect 20438 4001 20472 4035
rect 21328 4612 21362 4646
rect 21328 4522 21362 4556
rect 21328 4432 21362 4466
rect 21328 4342 21362 4376
rect 21328 4252 21362 4286
rect 21328 4162 21362 4196
rect 21328 4072 21362 4106
rect 21328 3982 21362 4016
rect 20516 3888 20550 3922
rect 20606 3888 20640 3922
rect 20696 3888 20730 3922
rect 20786 3888 20820 3922
rect 20876 3888 20910 3922
rect 20966 3888 21000 3922
rect 21056 3888 21090 3922
rect 21146 3888 21180 3922
rect 21236 3888 21270 3922
rect 21910 4778 21944 4812
rect 22000 4778 22034 4812
rect 22090 4778 22124 4812
rect 22180 4778 22214 4812
rect 22270 4778 22304 4812
rect 22360 4778 22394 4812
rect 22450 4778 22484 4812
rect 22540 4778 22574 4812
rect 22630 4778 22664 4812
rect 21798 4721 21832 4755
rect 22688 4702 22722 4736
rect 21798 4631 21832 4665
rect 21798 4541 21832 4575
rect 21798 4451 21832 4485
rect 21798 4361 21832 4395
rect 21798 4271 21832 4305
rect 21798 4181 21832 4215
rect 21798 4091 21832 4125
rect 21798 4001 21832 4035
rect 22688 4612 22722 4646
rect 22688 4522 22722 4556
rect 22688 4432 22722 4466
rect 22688 4342 22722 4376
rect 22688 4252 22722 4286
rect 22688 4162 22722 4196
rect 22688 4072 22722 4106
rect 22688 3982 22722 4016
rect 21876 3888 21910 3922
rect 21966 3888 22000 3922
rect 22056 3888 22090 3922
rect 22146 3888 22180 3922
rect 22236 3888 22270 3922
rect 22326 3888 22360 3922
rect 22416 3888 22450 3922
rect 22506 3888 22540 3922
rect 22596 3888 22630 3922
rect 23270 4778 23304 4812
rect 23360 4778 23394 4812
rect 23450 4778 23484 4812
rect 23540 4778 23574 4812
rect 23630 4778 23664 4812
rect 23720 4778 23754 4812
rect 23810 4778 23844 4812
rect 23900 4778 23934 4812
rect 23990 4778 24024 4812
rect 23158 4721 23192 4755
rect 24048 4702 24082 4736
rect 23158 4631 23192 4665
rect 23158 4541 23192 4575
rect 23158 4451 23192 4485
rect 23158 4361 23192 4395
rect 23158 4271 23192 4305
rect 23158 4181 23192 4215
rect 23158 4091 23192 4125
rect 23158 4001 23192 4035
rect 24048 4612 24082 4646
rect 24048 4522 24082 4556
rect 24048 4432 24082 4466
rect 24048 4342 24082 4376
rect 24048 4252 24082 4286
rect 24048 4162 24082 4196
rect 24048 4072 24082 4106
rect 24048 3982 24082 4016
rect 23236 3888 23270 3922
rect 23326 3888 23360 3922
rect 23416 3888 23450 3922
rect 23506 3888 23540 3922
rect 23596 3888 23630 3922
rect 23686 3888 23720 3922
rect 23776 3888 23810 3922
rect 23866 3888 23900 3922
rect 23956 3888 23990 3922
rect 26570 4150 26730 4190
rect 25310 3820 25350 3980
rect 27950 3820 27990 3980
rect 20550 3418 20584 3452
rect 20640 3418 20674 3452
rect 20730 3418 20764 3452
rect 20820 3418 20854 3452
rect 20910 3418 20944 3452
rect 21000 3418 21034 3452
rect 21090 3418 21124 3452
rect 21180 3418 21214 3452
rect 21270 3418 21304 3452
rect 20438 3361 20472 3395
rect 21328 3342 21362 3376
rect 20438 3271 20472 3305
rect 20438 3181 20472 3215
rect 20438 3091 20472 3125
rect 20438 3001 20472 3035
rect 20438 2911 20472 2945
rect 20438 2821 20472 2855
rect 20438 2731 20472 2765
rect 20438 2641 20472 2675
rect 21328 3252 21362 3286
rect 21328 3162 21362 3196
rect 21328 3072 21362 3106
rect 21328 2982 21362 3016
rect 21328 2892 21362 2926
rect 21328 2802 21362 2836
rect 21328 2712 21362 2746
rect 21328 2622 21362 2656
rect 20516 2528 20550 2562
rect 20606 2528 20640 2562
rect 20696 2528 20730 2562
rect 20786 2528 20820 2562
rect 20876 2528 20910 2562
rect 20966 2528 21000 2562
rect 21056 2528 21090 2562
rect 21146 2528 21180 2562
rect 21236 2528 21270 2562
rect 21910 3418 21944 3452
rect 22000 3418 22034 3452
rect 22090 3418 22124 3452
rect 22180 3418 22214 3452
rect 22270 3418 22304 3452
rect 22360 3418 22394 3452
rect 22450 3418 22484 3452
rect 22540 3418 22574 3452
rect 22630 3418 22664 3452
rect 21798 3361 21832 3395
rect 22688 3342 22722 3376
rect 21798 3271 21832 3305
rect 21798 3181 21832 3215
rect 21798 3091 21832 3125
rect 21798 3001 21832 3035
rect 21798 2911 21832 2945
rect 21798 2821 21832 2855
rect 21798 2731 21832 2765
rect 21798 2641 21832 2675
rect 22688 3252 22722 3286
rect 22688 3162 22722 3196
rect 22688 3072 22722 3106
rect 22688 2982 22722 3016
rect 22688 2892 22722 2926
rect 22688 2802 22722 2836
rect 22688 2712 22722 2746
rect 22688 2622 22722 2656
rect 21876 2528 21910 2562
rect 21966 2528 22000 2562
rect 22056 2528 22090 2562
rect 22146 2528 22180 2562
rect 22236 2528 22270 2562
rect 22326 2528 22360 2562
rect 22416 2528 22450 2562
rect 22506 2528 22540 2562
rect 22596 2528 22630 2562
rect 26570 3610 26730 3650
rect 29610 4150 29770 4190
rect 28350 3820 28390 3980
rect 30990 3820 31030 3980
rect 29610 3610 29770 3650
rect 23270 3418 23304 3452
rect 23360 3418 23394 3452
rect 23450 3418 23484 3452
rect 23540 3418 23574 3452
rect 23630 3418 23664 3452
rect 23720 3418 23754 3452
rect 23810 3418 23844 3452
rect 23900 3418 23934 3452
rect 23990 3418 24024 3452
rect 23158 3361 23192 3395
rect 24048 3342 24082 3376
rect 23158 3271 23192 3305
rect 23158 3181 23192 3215
rect 23158 3091 23192 3125
rect 23158 3001 23192 3035
rect 23158 2911 23192 2945
rect 23158 2821 23192 2855
rect 23158 2731 23192 2765
rect 23158 2641 23192 2675
rect 24048 3252 24082 3286
rect 24048 3162 24082 3196
rect 24048 3072 24082 3106
rect 24048 2982 24082 3016
rect 24048 2892 24082 2926
rect 24048 2802 24082 2836
rect 24048 2712 24082 2746
rect 24048 2622 24082 2656
rect 23236 2528 23270 2562
rect 23326 2528 23360 2562
rect 23416 2528 23450 2562
rect 23506 2528 23540 2562
rect 23596 2528 23630 2562
rect 23686 2528 23720 2562
rect 23776 2528 23810 2562
rect 23866 2528 23900 2562
rect 23956 2528 23990 2562
rect 20550 2058 20584 2092
rect 20640 2058 20674 2092
rect 20730 2058 20764 2092
rect 20820 2058 20854 2092
rect 20910 2058 20944 2092
rect 21000 2058 21034 2092
rect 21090 2058 21124 2092
rect 21180 2058 21214 2092
rect 21270 2058 21304 2092
rect 20438 2001 20472 2035
rect 21328 1982 21362 2016
rect 20438 1911 20472 1945
rect 20438 1821 20472 1855
rect 20438 1731 20472 1765
rect 20438 1641 20472 1675
rect 20438 1551 20472 1585
rect 20438 1461 20472 1495
rect 20438 1371 20472 1405
rect 20438 1281 20472 1315
rect 21328 1892 21362 1926
rect 21328 1802 21362 1836
rect 21328 1712 21362 1746
rect 21328 1622 21362 1656
rect 21328 1532 21362 1566
rect 21328 1442 21362 1476
rect 21328 1352 21362 1386
rect 21328 1262 21362 1296
rect 20516 1168 20550 1202
rect 20606 1168 20640 1202
rect 20696 1168 20730 1202
rect 20786 1168 20820 1202
rect 20876 1168 20910 1202
rect 20966 1168 21000 1202
rect 21056 1168 21090 1202
rect 21146 1168 21180 1202
rect 21236 1168 21270 1202
rect 21910 2058 21944 2092
rect 22000 2058 22034 2092
rect 22090 2058 22124 2092
rect 22180 2058 22214 2092
rect 22270 2058 22304 2092
rect 22360 2058 22394 2092
rect 22450 2058 22484 2092
rect 22540 2058 22574 2092
rect 22630 2058 22664 2092
rect 21798 2001 21832 2035
rect 22688 1982 22722 2016
rect 21798 1911 21832 1945
rect 21798 1821 21832 1855
rect 21798 1731 21832 1765
rect 21798 1641 21832 1675
rect 21798 1551 21832 1585
rect 21798 1461 21832 1495
rect 21798 1371 21832 1405
rect 21798 1281 21832 1315
rect 22688 1892 22722 1926
rect 22688 1802 22722 1836
rect 22688 1712 22722 1746
rect 22688 1622 22722 1656
rect 22688 1532 22722 1566
rect 22688 1442 22722 1476
rect 22688 1352 22722 1386
rect 22688 1262 22722 1296
rect 21876 1168 21910 1202
rect 21966 1168 22000 1202
rect 22056 1168 22090 1202
rect 22146 1168 22180 1202
rect 22236 1168 22270 1202
rect 22326 1168 22360 1202
rect 22416 1168 22450 1202
rect 22506 1168 22540 1202
rect 22596 1168 22630 1202
rect 23270 2058 23304 2092
rect 23360 2058 23394 2092
rect 23450 2058 23484 2092
rect 23540 2058 23574 2092
rect 23630 2058 23664 2092
rect 23720 2058 23754 2092
rect 23810 2058 23844 2092
rect 23900 2058 23934 2092
rect 23990 2058 24024 2092
rect 23158 2001 23192 2035
rect 24048 1982 24082 2016
rect 23158 1911 23192 1945
rect 23158 1821 23192 1855
rect 23158 1731 23192 1765
rect 23158 1641 23192 1675
rect 23158 1551 23192 1585
rect 23158 1461 23192 1495
rect 23158 1371 23192 1405
rect 23158 1281 23192 1315
rect 24048 1892 24082 1926
rect 24048 1802 24082 1836
rect 24048 1712 24082 1746
rect 24048 1622 24082 1656
rect 24048 1532 24082 1566
rect 24048 1442 24082 1476
rect 24048 1352 24082 1386
rect 24048 1262 24082 1296
rect 23236 1168 23270 1202
rect 23326 1168 23360 1202
rect 23416 1168 23450 1202
rect 23506 1168 23540 1202
rect 23596 1168 23630 1202
rect 23686 1168 23720 1202
rect 23776 1168 23810 1202
rect 23866 1168 23900 1202
rect 23956 1168 23990 1202
<< poly >>
rect 29830 6340 29900 6360
rect 29830 6300 29850 6340
rect 29890 6300 29900 6340
rect 29830 6280 29900 6300
rect 26230 6250 26330 6280
rect 26410 6250 26510 6280
rect 26590 6250 26690 6280
rect 26770 6250 26870 6280
rect 26950 6250 27050 6280
rect 27130 6250 27230 6280
rect 27310 6250 27410 6280
rect 27490 6250 27590 6280
rect 27670 6250 27770 6280
rect 27850 6250 27950 6280
rect 28030 6250 28130 6280
rect 28210 6250 28310 6280
rect 28390 6250 28490 6280
rect 28570 6250 28670 6280
rect 28750 6250 28850 6280
rect 28930 6250 29030 6280
rect 29110 6250 29210 6280
rect 29290 6250 29390 6280
rect 29470 6250 29570 6280
rect 29650 6250 29750 6280
rect 29830 6250 29930 6280
rect 30010 6250 30110 6280
rect 26230 6020 26330 6050
rect 26150 6000 26330 6020
rect 26410 6030 26510 6050
rect 26590 6030 26690 6050
rect 26770 6030 26870 6050
rect 26950 6030 27050 6050
rect 27130 6030 27230 6050
rect 27310 6030 27410 6050
rect 27490 6030 27590 6050
rect 27670 6030 27770 6050
rect 27850 6030 27950 6050
rect 28030 6030 28130 6050
rect 28210 6030 28310 6050
rect 28390 6030 28490 6050
rect 28570 6030 28670 6050
rect 28750 6030 28850 6050
rect 28930 6030 29030 6050
rect 29110 6030 29210 6050
rect 29290 6030 29390 6050
rect 29470 6030 29570 6050
rect 29650 6030 29750 6050
rect 29830 6030 29930 6050
rect 26410 6020 29930 6030
rect 30010 6020 30110 6050
rect 26410 6000 29950 6020
rect 26150 5960 26170 6000
rect 26210 5990 26330 6000
rect 26210 5960 26230 5990
rect 26150 5940 26230 5960
rect 29890 5960 29900 6000
rect 29940 5960 29950 6000
rect 30010 6000 30190 6020
rect 30010 5990 30130 6000
rect 29890 5940 29950 5960
rect 30110 5960 30130 5990
rect 30170 5960 30190 6000
rect 30110 5940 30190 5960
rect 25590 5100 25620 5130
rect 25700 5100 25730 5130
rect 25590 4880 25620 4900
rect 25700 4880 25730 4900
rect 25590 4850 25730 4880
rect 25620 4810 25640 4850
rect 25680 4810 25700 4850
rect 25620 4790 25700 4810
rect 26510 5420 26590 5440
rect 26510 5380 26530 5420
rect 26570 5390 26590 5420
rect 29750 5420 29830 5440
rect 29750 5390 29770 5420
rect 26570 5380 26690 5390
rect 26510 5360 26690 5380
rect 29650 5380 29770 5390
rect 29810 5380 29830 5420
rect 29650 5360 29830 5380
rect 26590 5330 26690 5360
rect 26770 5330 26870 5360
rect 26950 5330 27050 5360
rect 27130 5330 27230 5360
rect 27310 5330 27410 5360
rect 27490 5330 27590 5360
rect 27670 5330 27770 5360
rect 27850 5330 27950 5360
rect 28030 5330 28130 5360
rect 28210 5330 28310 5360
rect 28390 5330 28490 5360
rect 28570 5330 28670 5360
rect 28750 5330 28850 5360
rect 28930 5330 29030 5360
rect 29110 5330 29210 5360
rect 29290 5330 29390 5360
rect 29470 5330 29570 5360
rect 29650 5330 29750 5360
rect 26590 4700 26690 4730
rect 26770 4710 26870 4730
rect 26950 4710 27050 4730
rect 27130 4710 27230 4730
rect 27310 4710 27410 4730
rect 27490 4710 27590 4730
rect 27670 4710 27770 4730
rect 27850 4710 27950 4730
rect 28030 4710 28130 4730
rect 28210 4710 28310 4730
rect 28390 4710 28490 4730
rect 28570 4710 28670 4730
rect 28750 4710 28850 4730
rect 28930 4710 29030 4730
rect 29110 4710 29210 4730
rect 29290 4710 29390 4730
rect 29470 4710 29570 4730
rect 26770 4680 29570 4710
rect 29650 4700 29750 4730
rect 27650 4640 27670 4680
rect 27710 4640 27730 4680
rect 27650 4620 27730 4640
rect 29390 4640 29410 4680
rect 29450 4640 29470 4680
rect 29390 4620 29470 4640
rect 25490 4000 25530 4030
rect 25610 4000 25650 4030
rect 25730 4000 25770 4030
rect 25850 4000 25890 4030
rect 25970 4000 26010 4030
rect 26090 4000 26130 4030
rect 26210 4000 26250 4030
rect 26330 4000 26370 4030
rect 26450 4000 26490 4030
rect 26570 4000 26610 4030
rect 26690 4000 26730 4030
rect 26810 4000 26850 4030
rect 26930 4000 26970 4030
rect 27050 4000 27090 4030
rect 27170 4000 27210 4030
rect 27290 4000 27330 4030
rect 27410 4000 27450 4030
rect 27530 4000 27570 4030
rect 27650 4000 27690 4030
rect 27770 4000 27810 4030
rect 25490 3780 25530 3800
rect 25420 3750 25530 3780
rect 25610 3770 25650 3800
rect 25730 3780 25770 3800
rect 25850 3780 25890 3800
rect 25970 3780 26010 3800
rect 26090 3780 26130 3800
rect 25590 3750 25670 3770
rect 25730 3750 26130 3780
rect 26210 3780 26250 3800
rect 26330 3780 26370 3800
rect 26210 3750 26370 3780
rect 26450 3780 26490 3800
rect 26570 3780 26610 3800
rect 26690 3780 26730 3800
rect 26810 3780 26850 3800
rect 26450 3750 26850 3780
rect 26930 3780 26970 3800
rect 27050 3780 27090 3800
rect 26930 3750 27090 3780
rect 27170 3780 27210 3800
rect 27290 3780 27330 3800
rect 27410 3780 27450 3800
rect 27530 3780 27570 3800
rect 27170 3750 27570 3780
rect 27650 3770 27690 3800
rect 27770 3780 27810 3800
rect 27640 3750 27700 3770
rect 27770 3750 27880 3780
rect 25420 3710 25430 3750
rect 25470 3710 25480 3750
rect 25420 3690 25480 3710
rect 25590 3710 25610 3750
rect 25650 3710 25670 3750
rect 25590 3690 25670 3710
rect 25770 3710 25790 3750
rect 25830 3710 25850 3750
rect 25770 3690 25850 3710
rect 26250 3710 26270 3750
rect 26310 3710 26330 3750
rect 26250 3690 26330 3710
rect 26490 3710 26510 3750
rect 26550 3710 26570 3750
rect 26490 3690 26570 3710
rect 26970 3710 26990 3750
rect 27030 3710 27050 3750
rect 26970 3690 27050 3710
rect 27210 3710 27230 3750
rect 27270 3710 27290 3750
rect 27210 3690 27290 3710
rect 27640 3710 27650 3750
rect 27690 3710 27700 3750
rect 27640 3690 27700 3710
rect 27820 3710 27830 3750
rect 27870 3710 27880 3750
rect 27820 3690 27880 3710
rect 28530 4000 28570 4030
rect 28650 4000 28690 4030
rect 28770 4000 28810 4030
rect 28890 4000 28930 4030
rect 29010 4000 29050 4030
rect 29130 4000 29170 4030
rect 29250 4000 29290 4030
rect 29370 4000 29410 4030
rect 29490 4000 29530 4030
rect 29610 4000 29650 4030
rect 29730 4000 29770 4030
rect 29850 4000 29890 4030
rect 29970 4000 30010 4030
rect 30090 4000 30130 4030
rect 30210 4000 30250 4030
rect 30330 4000 30370 4030
rect 30450 4000 30490 4030
rect 30570 4000 30610 4030
rect 30690 4000 30730 4030
rect 30810 4000 30850 4030
rect 28530 3750 28570 3800
rect 28650 3770 28690 3800
rect 28770 3780 28810 3800
rect 28890 3780 28930 3800
rect 29010 3780 29050 3800
rect 29130 3780 29170 3800
rect 28640 3750 28700 3770
rect 28770 3750 29170 3780
rect 29250 3780 29290 3800
rect 29370 3780 29410 3800
rect 29250 3750 29410 3780
rect 29490 3780 29530 3800
rect 29610 3780 29650 3800
rect 29730 3780 29770 3800
rect 29850 3780 29890 3800
rect 29490 3750 29890 3780
rect 29970 3780 30010 3800
rect 30090 3780 30130 3800
rect 29970 3750 30130 3780
rect 30210 3780 30250 3800
rect 30330 3780 30370 3800
rect 30450 3780 30490 3800
rect 30570 3780 30610 3800
rect 30210 3750 30610 3780
rect 30690 3770 30730 3800
rect 30810 3780 30850 3800
rect 30670 3750 30750 3770
rect 30810 3750 30920 3780
rect 28640 3710 28650 3750
rect 28690 3710 28700 3750
rect 28640 3690 28700 3710
rect 29050 3710 29070 3750
rect 29110 3710 29130 3750
rect 29050 3690 29130 3710
rect 29290 3710 29310 3750
rect 29350 3710 29370 3750
rect 29290 3690 29370 3710
rect 29770 3710 29790 3750
rect 29830 3710 29850 3750
rect 29770 3690 29850 3710
rect 30010 3710 30030 3750
rect 30070 3710 30090 3750
rect 30010 3690 30090 3710
rect 30490 3710 30510 3750
rect 30550 3710 30570 3750
rect 30490 3690 30570 3710
rect 30670 3710 30690 3750
rect 30730 3710 30750 3750
rect 30670 3690 30750 3710
rect 30860 3710 30870 3750
rect 30910 3710 30920 3750
rect 30860 3690 30920 3710
rect 26390 3430 26470 3450
rect 26390 3390 26410 3430
rect 26450 3390 26470 3430
rect 26390 3360 26470 3390
rect 26390 3330 27470 3360
rect 26350 3250 26390 3280
rect 26470 3250 26510 3330
rect 26590 3250 26630 3330
rect 26710 3250 26750 3280
rect 26830 3250 26870 3280
rect 26950 3250 26990 3330
rect 27070 3250 27110 3330
rect 27190 3250 27230 3280
rect 27310 3250 27350 3280
rect 27430 3250 27470 3330
rect 26350 3120 26390 3150
rect 26470 3120 26510 3150
rect 26590 3120 26630 3150
rect 26270 3100 26390 3120
rect 26270 3060 26290 3100
rect 26330 3070 26390 3100
rect 26710 3070 26750 3150
rect 26830 3070 26870 3150
rect 26950 3120 26990 3150
rect 27070 3120 27110 3150
rect 27190 3070 27230 3150
rect 27310 3070 27350 3150
rect 27430 3120 27470 3150
rect 26330 3060 27350 3070
rect 26270 3040 27350 3060
rect 29870 3430 29950 3450
rect 29870 3390 29890 3430
rect 29930 3390 29950 3430
rect 29870 3360 29950 3390
rect 28870 3330 29950 3360
rect 28870 3250 28910 3330
rect 28990 3250 29030 3280
rect 29110 3250 29150 3280
rect 29230 3250 29270 3330
rect 29350 3250 29390 3330
rect 29470 3250 29510 3280
rect 29590 3250 29630 3280
rect 29710 3250 29750 3330
rect 29830 3250 29870 3330
rect 29950 3250 29990 3280
rect 28870 3120 28910 3150
rect 28990 3070 29030 3150
rect 29110 3070 29150 3150
rect 29230 3120 29270 3150
rect 29350 3120 29390 3150
rect 29470 3070 29510 3150
rect 29590 3070 29630 3150
rect 29710 3120 29750 3150
rect 29830 3120 29870 3150
rect 29950 3120 29990 3150
rect 29950 3100 30070 3120
rect 29950 3070 30010 3100
rect 28990 3060 30010 3070
rect 30050 3060 30070 3100
rect 28990 3040 30070 3060
rect 25970 2780 26050 2800
rect 25970 2740 25990 2780
rect 26030 2740 26050 2780
rect 25970 2730 26050 2740
rect 26210 2780 26290 2800
rect 26210 2740 26230 2780
rect 26270 2740 26290 2780
rect 26210 2730 26290 2740
rect 26450 2780 26530 2800
rect 26450 2740 26470 2780
rect 26510 2740 26530 2780
rect 26450 2730 26530 2740
rect 26690 2780 26770 2800
rect 26690 2740 26710 2780
rect 26750 2740 26770 2780
rect 26690 2730 26770 2740
rect 27170 2780 27250 2800
rect 27170 2740 27190 2780
rect 27230 2740 27250 2780
rect 27170 2730 27250 2740
rect 27410 2780 27490 2800
rect 27410 2740 27430 2780
rect 27470 2740 27490 2780
rect 27410 2730 27490 2740
rect 27650 2780 27730 2800
rect 27650 2740 27670 2780
rect 27710 2740 27730 2780
rect 27650 2730 27730 2740
rect 25870 2700 26870 2730
rect 26950 2700 27950 2730
rect 25870 2170 26870 2200
rect 26950 2170 27950 2200
rect 28610 2780 28690 2800
rect 28610 2740 28630 2780
rect 28670 2740 28690 2780
rect 28610 2730 28690 2740
rect 28850 2780 28930 2800
rect 28850 2740 28870 2780
rect 28910 2740 28930 2780
rect 28850 2730 28930 2740
rect 29090 2780 29170 2800
rect 29090 2740 29110 2780
rect 29150 2740 29170 2780
rect 29090 2730 29170 2740
rect 29570 2780 29650 2800
rect 29570 2740 29590 2780
rect 29630 2740 29650 2780
rect 29570 2730 29650 2740
rect 29810 2780 29890 2800
rect 29810 2740 29830 2780
rect 29870 2740 29890 2780
rect 29810 2730 29890 2740
rect 30050 2780 30130 2800
rect 30050 2740 30070 2780
rect 30110 2740 30130 2780
rect 30050 2730 30130 2740
rect 30290 2780 30370 2800
rect 30290 2740 30310 2780
rect 30350 2740 30370 2780
rect 30290 2730 30370 2740
rect 28390 2700 29390 2730
rect 29470 2700 30470 2730
rect 28390 2170 29390 2200
rect 29470 2170 30470 2200
rect 26210 1800 26290 1820
rect 26210 1760 26230 1800
rect 26270 1760 26290 1800
rect 26210 1740 26290 1760
rect 26370 1800 26450 1820
rect 26370 1760 26390 1800
rect 26430 1760 26450 1800
rect 26370 1740 26450 1760
rect 26530 1800 26610 1820
rect 26530 1760 26550 1800
rect 26590 1760 26610 1800
rect 26530 1740 26610 1760
rect 26690 1800 26770 1820
rect 26690 1760 26710 1800
rect 26750 1760 26770 1800
rect 26690 1740 26770 1760
rect 26850 1800 26930 1820
rect 26850 1760 26870 1800
rect 26910 1760 26930 1800
rect 26850 1740 26930 1760
rect 27010 1800 27090 1820
rect 27010 1760 27030 1800
rect 27070 1760 27090 1800
rect 27010 1740 27090 1760
rect 27170 1800 27250 1820
rect 27170 1760 27190 1800
rect 27230 1760 27250 1800
rect 27170 1740 27250 1760
rect 27330 1800 27410 1820
rect 27330 1760 27350 1800
rect 27390 1760 27410 1800
rect 27330 1740 27410 1760
rect 27490 1800 27570 1820
rect 27490 1760 27510 1800
rect 27550 1760 27570 1800
rect 27490 1740 27570 1760
rect 27650 1800 27730 1820
rect 27650 1760 27670 1800
rect 27710 1760 27730 1800
rect 27650 1740 27730 1760
rect 27810 1800 27890 1820
rect 27810 1760 27830 1800
rect 27870 1760 27890 1800
rect 27810 1740 27890 1760
rect 27970 1800 28050 1820
rect 27970 1760 27990 1800
rect 28030 1760 28050 1800
rect 27970 1740 28050 1760
rect 28290 1800 28370 1820
rect 28290 1760 28310 1800
rect 28350 1760 28370 1800
rect 28290 1740 28370 1760
rect 28450 1800 28530 1820
rect 28450 1760 28470 1800
rect 28510 1760 28530 1800
rect 28450 1740 28530 1760
rect 28610 1800 28690 1820
rect 28610 1760 28630 1800
rect 28670 1760 28690 1800
rect 28610 1740 28690 1760
rect 28770 1800 28850 1820
rect 28770 1760 28790 1800
rect 28830 1760 28850 1800
rect 28770 1740 28850 1760
rect 28930 1800 29010 1820
rect 28930 1760 28950 1800
rect 28990 1760 29010 1800
rect 28930 1740 29010 1760
rect 29090 1800 29170 1820
rect 29090 1760 29110 1800
rect 29150 1760 29170 1800
rect 29090 1740 29170 1760
rect 29250 1800 29330 1820
rect 29250 1760 29270 1800
rect 29310 1760 29330 1800
rect 29250 1740 29330 1760
rect 29410 1800 29490 1820
rect 29410 1760 29430 1800
rect 29470 1760 29490 1800
rect 29410 1740 29490 1760
rect 29570 1800 29650 1820
rect 29570 1760 29590 1800
rect 29630 1760 29650 1800
rect 29570 1740 29650 1760
rect 29730 1800 29810 1820
rect 29730 1760 29750 1800
rect 29790 1760 29810 1800
rect 29730 1740 29810 1760
rect 29890 1800 29970 1820
rect 29890 1760 29910 1800
rect 29950 1760 29970 1800
rect 29890 1740 29970 1760
rect 30050 1800 30130 1820
rect 30050 1760 30070 1800
rect 30110 1760 30130 1800
rect 30050 1740 30130 1760
rect 26130 1710 28130 1740
rect 28210 1710 30210 1740
rect 26130 1480 28130 1510
rect 28210 1480 30210 1510
rect 25470 1160 25570 1190
rect 25650 1180 26650 1210
rect 25650 1160 25750 1180
rect 25830 1160 25930 1180
rect 26010 1160 26110 1180
rect 26190 1160 26290 1180
rect 26370 1160 26470 1180
rect 26550 1160 26650 1180
rect 26730 1160 26830 1190
rect 25470 930 25570 960
rect 25650 930 25750 960
rect 25830 930 25930 960
rect 26010 930 26110 960
rect 26190 930 26290 960
rect 26370 930 26470 960
rect 26550 930 26650 960
rect 26730 930 26830 960
rect 27310 1160 27410 1190
rect 27490 1180 28850 1210
rect 27490 1160 27590 1180
rect 27670 1160 27770 1180
rect 27850 1160 27950 1180
rect 28030 1160 28130 1180
rect 28210 1160 28310 1180
rect 28390 1160 28490 1180
rect 28570 1160 28670 1180
rect 28750 1160 28850 1180
rect 28930 1160 29030 1190
rect 27310 930 27410 960
rect 27490 930 27590 960
rect 27670 930 27770 960
rect 27850 930 27950 960
rect 28030 930 28130 960
rect 28210 930 28310 960
rect 28390 930 28490 960
rect 28570 930 28670 960
rect 28750 930 28850 960
rect 28930 930 29030 960
rect 29470 1160 29570 1190
rect 29650 1180 30650 1210
rect 29650 1160 29750 1180
rect 29830 1160 29930 1180
rect 30010 1160 30110 1180
rect 30190 1160 30290 1180
rect 30370 1160 30470 1180
rect 30550 1160 30650 1180
rect 30730 1160 30830 1190
rect 29470 930 29570 960
rect 29650 930 29750 960
rect 29830 930 29930 960
rect 30010 930 30110 960
rect 30190 930 30290 960
rect 30370 930 30470 960
rect 30550 930 30650 960
rect 30730 930 30830 960
<< polycont >>
rect 29850 6300 29890 6340
rect 26170 5960 26210 6000
rect 29900 5960 29940 6000
rect 30130 5960 30170 6000
rect 25640 4810 25680 4850
rect 26530 5380 26570 5420
rect 29770 5380 29810 5420
rect 27670 4640 27710 4680
rect 29410 4640 29450 4680
rect 25430 3710 25470 3750
rect 25610 3710 25650 3750
rect 25790 3710 25830 3750
rect 26270 3710 26310 3750
rect 26510 3710 26550 3750
rect 26990 3710 27030 3750
rect 27230 3710 27270 3750
rect 27650 3710 27690 3750
rect 27830 3710 27870 3750
rect 28650 3710 28690 3750
rect 29070 3710 29110 3750
rect 29310 3710 29350 3750
rect 29790 3710 29830 3750
rect 30030 3710 30070 3750
rect 30510 3710 30550 3750
rect 30690 3710 30730 3750
rect 30870 3710 30910 3750
rect 26410 3390 26450 3430
rect 26290 3060 26330 3100
rect 29890 3390 29930 3430
rect 30010 3060 30050 3100
rect 25990 2740 26030 2780
rect 26230 2740 26270 2780
rect 26470 2740 26510 2780
rect 26710 2740 26750 2780
rect 27190 2740 27230 2780
rect 27430 2740 27470 2780
rect 27670 2740 27710 2780
rect 28630 2740 28670 2780
rect 28870 2740 28910 2780
rect 29110 2740 29150 2780
rect 29590 2740 29630 2780
rect 29830 2740 29870 2780
rect 30070 2740 30110 2780
rect 30310 2740 30350 2780
rect 26230 1760 26270 1800
rect 26390 1760 26430 1800
rect 26550 1760 26590 1800
rect 26710 1760 26750 1800
rect 26870 1760 26910 1800
rect 27030 1760 27070 1800
rect 27190 1760 27230 1800
rect 27350 1760 27390 1800
rect 27510 1760 27550 1800
rect 27670 1760 27710 1800
rect 27830 1760 27870 1800
rect 27990 1760 28030 1800
rect 28310 1760 28350 1800
rect 28470 1760 28510 1800
rect 28630 1760 28670 1800
rect 28790 1760 28830 1800
rect 28950 1760 28990 1800
rect 29110 1760 29150 1800
rect 29270 1760 29310 1800
rect 29430 1760 29470 1800
rect 29590 1760 29630 1800
rect 29750 1760 29790 1800
rect 29910 1760 29950 1800
rect 30070 1760 30110 1800
<< xpolycontact >>
rect 20182 6340 20622 6410
rect 21850 6340 22290 6410
rect 22612 6330 23052 6400
rect 24220 6330 24660 6400
rect 20182 6220 20622 6290
rect 21850 6220 22290 6290
rect 22612 6210 23052 6280
rect 24220 6210 24660 6280
rect 20182 6060 20622 6130
rect 21790 6060 22230 6130
rect 22612 6090 23052 6160
rect 24220 6090 24660 6160
rect 20182 5940 20622 6010
rect 21790 5940 22230 6010
rect 22612 5970 23052 6040
rect 24220 5970 24660 6040
rect 22612 5850 23052 5920
rect 24220 5850 24660 5920
rect 22612 5730 23052 5800
rect 24220 5730 24660 5800
rect 20192 5620 20630 5690
rect 21008 5620 21448 5690
rect 22612 5610 23052 5680
rect 23480 5610 23920 5680
rect 20192 5500 20630 5570
rect 21008 5500 21448 5570
<< ppolyres >>
rect 20630 5620 21008 5690
rect 20630 5500 21008 5570
<< xpolyres >>
rect 20622 6340 21850 6410
rect 23052 6330 24220 6400
rect 20622 6220 21850 6290
rect 23052 6210 24220 6280
rect 20622 6060 21790 6130
rect 23052 6090 24220 6160
rect 20622 5940 21790 6010
rect 23052 5970 24220 6040
rect 23052 5850 24220 5920
rect 23052 5730 24220 5800
rect 23052 5610 23480 5680
<< locali >>
rect 28890 6930 28950 6990
rect 21890 6830 21950 6890
rect 23290 6830 23350 6890
rect 30290 6830 30350 6890
rect 25390 6720 25450 6780
rect 26790 6610 26850 6670
rect 20092 6400 20182 6410
rect 20092 6350 20112 6400
rect 20162 6350 20182 6400
rect 20092 6340 20182 6350
rect 25970 6400 30370 6440
rect 22220 6290 22290 6340
rect 22522 6390 22612 6400
rect 22522 6340 22542 6390
rect 22592 6340 22612 6390
rect 22522 6330 22612 6340
rect 24660 6330 24740 6400
rect 20092 6280 20182 6290
rect 20092 6230 20112 6280
rect 20162 6230 20182 6280
rect 20092 6220 20182 6230
rect 22522 6270 22612 6280
rect 22522 6220 22542 6270
rect 22592 6220 22612 6270
rect 22522 6210 22612 6220
rect 24590 6160 24660 6210
rect 20092 6120 20182 6130
rect 20092 6070 20112 6120
rect 20162 6070 20182 6120
rect 20092 6060 20182 6070
rect 22160 6010 22230 6060
rect 20092 6000 20182 6010
rect 20092 5950 20112 6000
rect 20162 5950 20182 6000
rect 20092 5940 20182 5950
rect 22532 6090 22612 6160
rect 21820 5820 22240 5830
rect 21820 5760 21840 5820
rect 21900 5760 22000 5820
rect 22060 5760 22160 5820
rect 22220 5760 22240 5820
rect 21820 5750 22240 5760
rect 22532 5800 22572 6090
rect 24700 6040 24740 6330
rect 24660 5970 24740 6040
rect 22612 5920 22682 5970
rect 24660 5910 24750 5920
rect 24660 5860 24680 5910
rect 24730 5860 24750 5910
rect 25970 5900 26010 6400
rect 26320 6340 26400 6360
rect 26320 6300 26340 6340
rect 26380 6300 26400 6340
rect 26320 6280 26400 6300
rect 26690 6340 26770 6360
rect 26690 6300 26710 6340
rect 26750 6300 26770 6340
rect 26690 6280 26770 6300
rect 27050 6340 27130 6360
rect 27050 6300 27070 6340
rect 27110 6300 27130 6340
rect 27050 6280 27130 6300
rect 27410 6340 27490 6360
rect 27410 6300 27430 6340
rect 27470 6300 27490 6340
rect 27410 6280 27490 6300
rect 27770 6340 27850 6360
rect 27770 6300 27790 6340
rect 27830 6300 27850 6340
rect 27770 6280 27850 6300
rect 28130 6340 28210 6360
rect 28130 6300 28150 6340
rect 28190 6300 28210 6340
rect 28130 6280 28210 6300
rect 28490 6340 28570 6360
rect 28490 6300 28510 6340
rect 28550 6300 28570 6340
rect 28490 6280 28570 6300
rect 28850 6340 28930 6360
rect 28850 6300 28870 6340
rect 28910 6300 28930 6340
rect 28850 6280 28930 6300
rect 29210 6340 29290 6360
rect 29210 6300 29230 6340
rect 29270 6300 29290 6340
rect 29210 6280 29290 6300
rect 29570 6340 29650 6360
rect 29570 6300 29590 6340
rect 29630 6300 29650 6340
rect 29570 6280 29650 6300
rect 29830 6340 29900 6360
rect 29830 6300 29850 6340
rect 29890 6300 29900 6340
rect 29830 6280 29900 6300
rect 29940 6340 30010 6360
rect 29940 6300 29950 6340
rect 29990 6300 30010 6340
rect 29940 6280 30010 6300
rect 26350 6240 26390 6280
rect 26710 6240 26750 6280
rect 27070 6240 27110 6280
rect 27430 6240 27470 6280
rect 27790 6240 27830 6280
rect 28150 6240 28190 6280
rect 28510 6240 28550 6280
rect 28870 6240 28910 6280
rect 29230 6240 29270 6280
rect 29590 6240 29630 6280
rect 29950 6240 29990 6280
rect 26080 6220 26220 6240
rect 26080 6180 26090 6220
rect 26130 6180 26170 6220
rect 26210 6180 26220 6220
rect 26080 6120 26220 6180
rect 26080 6080 26090 6120
rect 26130 6080 26170 6120
rect 26210 6080 26220 6120
rect 26080 6060 26220 6080
rect 26340 6220 26400 6240
rect 26340 6180 26350 6220
rect 26390 6180 26400 6220
rect 26340 6120 26400 6180
rect 26340 6080 26350 6120
rect 26390 6080 26400 6120
rect 26340 6060 26400 6080
rect 26520 6220 26580 6240
rect 26520 6180 26530 6220
rect 26570 6180 26580 6220
rect 26520 6120 26580 6180
rect 26520 6080 26530 6120
rect 26570 6080 26580 6120
rect 26520 6060 26580 6080
rect 26700 6220 26760 6240
rect 26700 6180 26710 6220
rect 26750 6180 26760 6220
rect 26700 6120 26760 6180
rect 26700 6080 26710 6120
rect 26750 6080 26760 6120
rect 26700 6060 26760 6080
rect 26880 6220 26940 6240
rect 26880 6180 26890 6220
rect 26930 6180 26940 6220
rect 26880 6120 26940 6180
rect 26880 6080 26890 6120
rect 26930 6080 26940 6120
rect 26880 6060 26940 6080
rect 27060 6220 27120 6240
rect 27060 6180 27070 6220
rect 27110 6180 27120 6220
rect 27060 6120 27120 6180
rect 27060 6080 27070 6120
rect 27110 6080 27120 6120
rect 27060 6060 27120 6080
rect 27240 6220 27300 6240
rect 27240 6180 27250 6220
rect 27290 6180 27300 6220
rect 27240 6120 27300 6180
rect 27240 6080 27250 6120
rect 27290 6080 27300 6120
rect 27240 6060 27300 6080
rect 27420 6220 27480 6240
rect 27420 6180 27430 6220
rect 27470 6180 27480 6220
rect 27420 6120 27480 6180
rect 27420 6080 27430 6120
rect 27470 6080 27480 6120
rect 27420 6060 27480 6080
rect 27600 6220 27660 6240
rect 27600 6180 27610 6220
rect 27650 6180 27660 6220
rect 27600 6120 27660 6180
rect 27600 6080 27610 6120
rect 27650 6080 27660 6120
rect 27600 6060 27660 6080
rect 27780 6220 27840 6240
rect 27780 6180 27790 6220
rect 27830 6180 27840 6220
rect 27780 6120 27840 6180
rect 27780 6080 27790 6120
rect 27830 6080 27840 6120
rect 27780 6060 27840 6080
rect 27960 6220 28020 6240
rect 27960 6180 27970 6220
rect 28010 6180 28020 6220
rect 27960 6120 28020 6180
rect 27960 6080 27970 6120
rect 28010 6080 28020 6120
rect 27960 6060 28020 6080
rect 28140 6220 28200 6240
rect 28140 6180 28150 6220
rect 28190 6180 28200 6220
rect 28140 6120 28200 6180
rect 28140 6080 28150 6120
rect 28190 6080 28200 6120
rect 28140 6060 28200 6080
rect 28320 6220 28380 6240
rect 28320 6180 28330 6220
rect 28370 6180 28380 6220
rect 28320 6120 28380 6180
rect 28320 6080 28330 6120
rect 28370 6080 28380 6120
rect 28320 6060 28380 6080
rect 28500 6220 28560 6240
rect 28500 6180 28510 6220
rect 28550 6180 28560 6220
rect 28500 6120 28560 6180
rect 28500 6080 28510 6120
rect 28550 6080 28560 6120
rect 28500 6060 28560 6080
rect 28680 6220 28740 6240
rect 28680 6180 28690 6220
rect 28730 6180 28740 6220
rect 28680 6120 28740 6180
rect 28680 6080 28690 6120
rect 28730 6080 28740 6120
rect 28680 6060 28740 6080
rect 28860 6220 28920 6240
rect 28860 6180 28870 6220
rect 28910 6180 28920 6220
rect 28860 6120 28920 6180
rect 28860 6080 28870 6120
rect 28910 6080 28920 6120
rect 28860 6060 28920 6080
rect 29040 6220 29100 6240
rect 29040 6180 29050 6220
rect 29090 6180 29100 6220
rect 29040 6120 29100 6180
rect 29040 6080 29050 6120
rect 29090 6080 29100 6120
rect 29040 6060 29100 6080
rect 29220 6220 29280 6240
rect 29220 6180 29230 6220
rect 29270 6180 29280 6220
rect 29220 6120 29280 6180
rect 29220 6080 29230 6120
rect 29270 6080 29280 6120
rect 29220 6060 29280 6080
rect 29400 6220 29460 6240
rect 29400 6180 29410 6220
rect 29450 6180 29460 6220
rect 29400 6120 29460 6180
rect 29400 6080 29410 6120
rect 29450 6080 29460 6120
rect 29400 6060 29460 6080
rect 29580 6220 29640 6240
rect 29580 6180 29590 6220
rect 29630 6180 29640 6220
rect 29580 6120 29640 6180
rect 29580 6080 29590 6120
rect 29630 6080 29640 6120
rect 29580 6060 29640 6080
rect 29760 6220 29820 6240
rect 29760 6180 29770 6220
rect 29810 6180 29820 6220
rect 29760 6120 29820 6180
rect 29760 6080 29770 6120
rect 29810 6080 29820 6120
rect 29760 6060 29820 6080
rect 29940 6220 30000 6240
rect 29940 6180 29950 6220
rect 29990 6180 30000 6220
rect 29940 6120 30000 6180
rect 29940 6080 29950 6120
rect 29990 6080 30000 6120
rect 29940 6060 30000 6080
rect 30120 6220 30260 6240
rect 30120 6180 30130 6220
rect 30170 6180 30210 6220
rect 30250 6180 30260 6220
rect 30120 6120 30260 6180
rect 30120 6080 30130 6120
rect 30170 6080 30210 6120
rect 30250 6080 30260 6120
rect 30120 6060 30260 6080
rect 26170 6020 26210 6060
rect 26530 6020 26570 6060
rect 26890 6020 26930 6060
rect 27250 6020 27290 6060
rect 27610 6020 27650 6060
rect 27970 6020 28010 6060
rect 28330 6020 28370 6060
rect 28690 6020 28730 6060
rect 29050 6020 29090 6060
rect 29410 6020 29450 6060
rect 29770 6020 29810 6060
rect 30130 6020 30170 6060
rect 26150 6000 26230 6020
rect 26150 5960 26170 6000
rect 26210 5960 26230 6000
rect 26150 5940 26230 5960
rect 26510 6000 26590 6020
rect 26510 5960 26530 6000
rect 26570 5960 26590 6000
rect 26510 5940 26590 5960
rect 26870 6000 26950 6020
rect 26870 5960 26890 6000
rect 26930 5960 26950 6000
rect 26870 5940 26950 5960
rect 27230 6000 27310 6020
rect 27230 5960 27250 6000
rect 27290 5960 27310 6000
rect 27230 5940 27310 5960
rect 27590 6000 27670 6020
rect 27590 5960 27610 6000
rect 27650 5960 27670 6000
rect 27590 5940 27670 5960
rect 27950 6000 28030 6020
rect 27950 5960 27970 6000
rect 28010 5960 28030 6000
rect 27950 5940 28030 5960
rect 28310 6000 28390 6020
rect 28310 5960 28330 6000
rect 28370 5960 28390 6000
rect 28310 5940 28390 5960
rect 28670 6000 28750 6020
rect 28670 5960 28690 6000
rect 28730 5960 28750 6000
rect 28670 5940 28750 5960
rect 29030 6000 29110 6020
rect 29030 5960 29050 6000
rect 29090 5960 29110 6000
rect 29030 5940 29110 5960
rect 29390 6000 29470 6020
rect 29390 5960 29410 6000
rect 29450 5960 29470 6000
rect 29390 5940 29470 5960
rect 29750 6000 29830 6020
rect 29750 5960 29770 6000
rect 29810 5960 29830 6000
rect 29750 5940 29830 5960
rect 29890 6000 29950 6020
rect 29890 5960 29900 6000
rect 29940 5960 29950 6000
rect 29890 5940 29950 5960
rect 30110 6000 30190 6020
rect 30110 5960 30130 6000
rect 30170 5960 30190 6000
rect 30110 5940 30190 5960
rect 30330 5900 30370 6400
rect 25970 5860 30370 5900
rect 24660 5850 24750 5860
rect 22532 5730 22612 5800
rect 24660 5790 24750 5810
rect 24660 5740 24680 5790
rect 24730 5740 24750 5790
rect 24660 5720 24750 5740
rect 20102 5680 20192 5690
rect 20102 5630 20122 5680
rect 20172 5630 20192 5680
rect 20102 5620 20192 5630
rect 21448 5680 21538 5690
rect 21448 5630 21468 5680
rect 21518 5630 21538 5680
rect 21448 5620 21538 5630
rect 22522 5670 22612 5680
rect 22522 5620 22542 5670
rect 22592 5620 22612 5670
rect 22522 5610 22612 5620
rect 23920 5670 24010 5680
rect 23920 5620 23940 5670
rect 23990 5620 24010 5670
rect 23920 5610 24010 5620
rect 20102 5560 20192 5570
rect 20102 5510 20122 5560
rect 20172 5510 20192 5560
rect 20102 5500 20192 5510
rect 21448 5560 21538 5570
rect 21448 5510 21468 5560
rect 21518 5510 21538 5560
rect 21448 5500 21538 5510
rect 26400 5480 29930 5520
rect 25520 5070 25580 5090
rect 25520 5030 25530 5070
rect 25570 5030 25580 5070
rect 21300 4994 21550 5000
rect 22660 4994 22910 5000
rect 24020 4994 24270 5000
rect 20256 4959 21550 4994
rect 20256 4936 20386 4959
rect 20256 4902 20290 4936
rect 20324 4925 20386 4936
rect 20420 4925 20476 4959
rect 20510 4925 20566 4959
rect 20600 4925 20656 4959
rect 20690 4925 20746 4959
rect 20780 4925 20836 4959
rect 20870 4925 20926 4959
rect 20960 4925 21016 4959
rect 21050 4925 21106 4959
rect 21140 4925 21196 4959
rect 21230 4925 21286 4959
rect 21320 4925 21376 4959
rect 21410 4936 21550 4959
rect 21410 4925 21477 4936
rect 20324 4902 21477 4925
rect 21511 4902 21550 4936
rect 20256 4895 21550 4902
rect 20256 4846 20355 4895
rect 20256 4812 20290 4846
rect 20324 4812 20355 4846
rect 21300 4846 21550 4895
rect 21300 4831 21477 4846
rect 20256 4756 20355 4812
rect 20256 4722 20290 4756
rect 20324 4722 20355 4756
rect 20256 4666 20355 4722
rect 20256 4632 20290 4666
rect 20324 4632 20355 4666
rect 20256 4576 20355 4632
rect 20256 4542 20290 4576
rect 20324 4542 20355 4576
rect 20256 4486 20355 4542
rect 20256 4452 20290 4486
rect 20324 4452 20355 4486
rect 20256 4396 20355 4452
rect 20256 4362 20290 4396
rect 20324 4362 20355 4396
rect 20256 4306 20355 4362
rect 20256 4272 20290 4306
rect 20324 4272 20355 4306
rect 20256 4216 20355 4272
rect 20256 4182 20290 4216
rect 20324 4182 20355 4216
rect 20256 4126 20355 4182
rect 20256 4092 20290 4126
rect 20324 4092 20355 4126
rect 20256 4036 20355 4092
rect 20256 4002 20290 4036
rect 20324 4002 20355 4036
rect 20256 3946 20355 4002
rect 20256 3912 20290 3946
rect 20324 3912 20355 3946
rect 20256 3856 20355 3912
rect 20419 4812 21477 4831
rect 21511 4812 21550 4846
rect 20419 4778 20550 4812
rect 20584 4778 20640 4812
rect 20674 4778 20730 4812
rect 20764 4778 20820 4812
rect 20854 4778 20910 4812
rect 20944 4778 21000 4812
rect 21034 4778 21090 4812
rect 21124 4778 21180 4812
rect 21214 4778 21270 4812
rect 21304 4778 21550 4812
rect 20419 4759 21550 4778
rect 20419 4755 20491 4759
rect 20419 4721 20438 4755
rect 20472 4721 20491 4755
rect 20419 4665 20491 4721
rect 21300 4756 21550 4759
rect 21300 4736 21477 4756
rect 21300 4702 21328 4736
rect 21362 4722 21477 4736
rect 21511 4722 21550 4756
rect 21362 4702 21550 4722
rect 20419 4631 20438 4665
rect 20472 4631 20491 4665
rect 20419 4575 20491 4631
rect 20419 4541 20438 4575
rect 20472 4541 20491 4575
rect 20419 4485 20491 4541
rect 20419 4451 20438 4485
rect 20472 4451 20491 4485
rect 20419 4395 20491 4451
rect 20419 4361 20438 4395
rect 20472 4361 20491 4395
rect 20419 4305 20491 4361
rect 20419 4271 20438 4305
rect 20472 4271 20491 4305
rect 20419 4215 20491 4271
rect 20419 4181 20438 4215
rect 20472 4181 20491 4215
rect 20419 4125 20491 4181
rect 20419 4091 20438 4125
rect 20472 4091 20491 4125
rect 20419 4035 20491 4091
rect 20419 4001 20438 4035
rect 20472 4001 20491 4035
rect 20553 4638 21247 4697
rect 20553 4604 20614 4638
rect 20648 4610 20704 4638
rect 20738 4610 20794 4638
rect 20828 4610 20884 4638
rect 20660 4604 20704 4610
rect 20760 4604 20794 4610
rect 20860 4604 20884 4610
rect 20918 4610 20974 4638
rect 20918 4604 20926 4610
rect 20553 4576 20626 4604
rect 20660 4576 20726 4604
rect 20760 4576 20826 4604
rect 20860 4576 20926 4604
rect 20960 4604 20974 4610
rect 21008 4610 21064 4638
rect 21008 4604 21026 4610
rect 20960 4576 21026 4604
rect 21060 4604 21064 4610
rect 21098 4610 21154 4638
rect 21098 4604 21126 4610
rect 21188 4604 21247 4638
rect 21060 4576 21126 4604
rect 21160 4576 21247 4604
rect 20553 4548 21247 4576
rect 20553 4514 20614 4548
rect 20648 4514 20704 4548
rect 20738 4514 20794 4548
rect 20828 4514 20884 4548
rect 20918 4514 20974 4548
rect 21008 4514 21064 4548
rect 21098 4514 21154 4548
rect 21188 4514 21247 4548
rect 20553 4510 21247 4514
rect 20553 4476 20626 4510
rect 20660 4476 20726 4510
rect 20760 4476 20826 4510
rect 20860 4476 20926 4510
rect 20960 4476 21026 4510
rect 21060 4476 21126 4510
rect 21160 4476 21247 4510
rect 20553 4458 21247 4476
rect 20553 4424 20614 4458
rect 20648 4424 20704 4458
rect 20738 4424 20794 4458
rect 20828 4424 20884 4458
rect 20918 4424 20974 4458
rect 21008 4424 21064 4458
rect 21098 4424 21154 4458
rect 21188 4424 21247 4458
rect 20553 4410 21247 4424
rect 20553 4376 20626 4410
rect 20660 4376 20726 4410
rect 20760 4376 20826 4410
rect 20860 4376 20926 4410
rect 20960 4376 21026 4410
rect 21060 4376 21126 4410
rect 21160 4376 21247 4410
rect 20553 4368 21247 4376
rect 20553 4334 20614 4368
rect 20648 4334 20704 4368
rect 20738 4334 20794 4368
rect 20828 4334 20884 4368
rect 20918 4334 20974 4368
rect 21008 4334 21064 4368
rect 21098 4334 21154 4368
rect 21188 4334 21247 4368
rect 20553 4310 21247 4334
rect 20553 4278 20626 4310
rect 20660 4278 20726 4310
rect 20760 4278 20826 4310
rect 20860 4278 20926 4310
rect 20553 4244 20614 4278
rect 20660 4276 20704 4278
rect 20760 4276 20794 4278
rect 20860 4276 20884 4278
rect 20648 4244 20704 4276
rect 20738 4244 20794 4276
rect 20828 4244 20884 4276
rect 20918 4276 20926 4278
rect 20960 4278 21026 4310
rect 20960 4276 20974 4278
rect 20918 4244 20974 4276
rect 21008 4276 21026 4278
rect 21060 4278 21126 4310
rect 21160 4278 21247 4310
rect 21060 4276 21064 4278
rect 21008 4244 21064 4276
rect 21098 4276 21126 4278
rect 21098 4244 21154 4276
rect 21188 4244 21247 4278
rect 20553 4210 21247 4244
rect 20553 4188 20626 4210
rect 20660 4188 20726 4210
rect 20760 4188 20826 4210
rect 20860 4188 20926 4210
rect 20553 4154 20614 4188
rect 20660 4176 20704 4188
rect 20760 4176 20794 4188
rect 20860 4176 20884 4188
rect 20648 4154 20704 4176
rect 20738 4154 20794 4176
rect 20828 4154 20884 4176
rect 20918 4176 20926 4188
rect 20960 4188 21026 4210
rect 20960 4176 20974 4188
rect 20918 4154 20974 4176
rect 21008 4176 21026 4188
rect 21060 4188 21126 4210
rect 21160 4188 21247 4210
rect 21060 4176 21064 4188
rect 21008 4154 21064 4176
rect 21098 4176 21126 4188
rect 21098 4154 21154 4176
rect 21188 4154 21247 4188
rect 20553 4110 21247 4154
rect 20553 4098 20626 4110
rect 20660 4098 20726 4110
rect 20760 4098 20826 4110
rect 20860 4098 20926 4110
rect 20553 4064 20614 4098
rect 20660 4076 20704 4098
rect 20760 4076 20794 4098
rect 20860 4076 20884 4098
rect 20648 4064 20704 4076
rect 20738 4064 20794 4076
rect 20828 4064 20884 4076
rect 20918 4076 20926 4098
rect 20960 4098 21026 4110
rect 20960 4076 20974 4098
rect 20918 4064 20974 4076
rect 21008 4076 21026 4098
rect 21060 4098 21126 4110
rect 21160 4098 21247 4110
rect 21060 4076 21064 4098
rect 21008 4064 21064 4076
rect 21098 4076 21126 4098
rect 21098 4064 21154 4076
rect 21188 4064 21247 4098
rect 20553 4003 21247 4064
rect 21300 4666 21550 4702
rect 21300 4646 21477 4666
rect 21300 4612 21328 4646
rect 21362 4632 21477 4646
rect 21511 4632 21550 4666
rect 21362 4612 21550 4632
rect 21300 4576 21550 4612
rect 21300 4556 21477 4576
rect 21300 4522 21328 4556
rect 21362 4542 21477 4556
rect 21511 4542 21550 4576
rect 21362 4522 21550 4542
rect 21300 4486 21550 4522
rect 21300 4466 21477 4486
rect 21300 4432 21328 4466
rect 21362 4452 21477 4466
rect 21511 4452 21550 4486
rect 21362 4432 21550 4452
rect 21300 4396 21550 4432
rect 21300 4376 21477 4396
rect 21300 4342 21328 4376
rect 21362 4362 21477 4376
rect 21511 4362 21550 4396
rect 21362 4342 21550 4362
rect 21300 4306 21550 4342
rect 21300 4286 21477 4306
rect 21300 4252 21328 4286
rect 21362 4272 21477 4286
rect 21511 4272 21550 4306
rect 21362 4252 21550 4272
rect 21300 4216 21550 4252
rect 21300 4196 21477 4216
rect 21300 4162 21328 4196
rect 21362 4182 21477 4196
rect 21511 4182 21550 4216
rect 21362 4162 21550 4182
rect 21300 4126 21550 4162
rect 21300 4106 21477 4126
rect 21300 4072 21328 4106
rect 21362 4092 21477 4106
rect 21511 4092 21550 4126
rect 21362 4072 21550 4092
rect 21300 4036 21550 4072
rect 21300 4016 21477 4036
rect 20419 3941 20491 4001
rect 21300 3982 21328 4016
rect 21362 4002 21477 4016
rect 21511 4002 21550 4036
rect 21362 3982 21550 4002
rect 21300 3946 21550 3982
rect 21300 3941 21477 3946
rect 20419 3922 21477 3941
rect 20419 3888 20516 3922
rect 20550 3888 20606 3922
rect 20640 3888 20696 3922
rect 20730 3888 20786 3922
rect 20820 3888 20876 3922
rect 20910 3888 20966 3922
rect 21000 3888 21056 3922
rect 21090 3888 21146 3922
rect 21180 3888 21236 3922
rect 21270 3912 21477 3922
rect 21511 3912 21550 3946
rect 21270 3888 21550 3912
rect 20419 3869 21550 3888
rect 20256 3822 20290 3856
rect 20324 3822 20355 3856
rect 20256 3805 20355 3822
rect 21300 3856 21550 3869
rect 21300 3822 21477 3856
rect 21511 3822 21550 3856
rect 21300 3805 21550 3822
rect 20256 3772 21550 3805
rect 20256 3738 20386 3772
rect 20420 3738 20476 3772
rect 20510 3738 20566 3772
rect 20600 3738 20656 3772
rect 20690 3738 20746 3772
rect 20780 3738 20836 3772
rect 20870 3738 20926 3772
rect 20960 3738 21016 3772
rect 21050 3738 21106 3772
rect 21140 3738 21196 3772
rect 21230 3738 21286 3772
rect 21320 3738 21376 3772
rect 21410 3738 21550 3772
rect 20256 3710 21550 3738
rect 21616 4959 22910 4994
rect 21616 4936 21746 4959
rect 21616 4902 21650 4936
rect 21684 4925 21746 4936
rect 21780 4925 21836 4959
rect 21870 4925 21926 4959
rect 21960 4925 22016 4959
rect 22050 4925 22106 4959
rect 22140 4925 22196 4959
rect 22230 4925 22286 4959
rect 22320 4925 22376 4959
rect 22410 4925 22466 4959
rect 22500 4925 22556 4959
rect 22590 4925 22646 4959
rect 22680 4925 22736 4959
rect 22770 4936 22910 4959
rect 22770 4925 22837 4936
rect 21684 4902 22837 4925
rect 22871 4902 22910 4936
rect 21616 4895 22910 4902
rect 21616 4846 21715 4895
rect 21616 4812 21650 4846
rect 21684 4812 21715 4846
rect 22660 4846 22910 4895
rect 22660 4831 22837 4846
rect 21616 4756 21715 4812
rect 21616 4722 21650 4756
rect 21684 4722 21715 4756
rect 21616 4666 21715 4722
rect 21616 4632 21650 4666
rect 21684 4632 21715 4666
rect 21616 4576 21715 4632
rect 21616 4542 21650 4576
rect 21684 4542 21715 4576
rect 21616 4486 21715 4542
rect 21616 4452 21650 4486
rect 21684 4452 21715 4486
rect 21616 4396 21715 4452
rect 21616 4362 21650 4396
rect 21684 4362 21715 4396
rect 21616 4306 21715 4362
rect 21616 4272 21650 4306
rect 21684 4272 21715 4306
rect 21616 4216 21715 4272
rect 21616 4182 21650 4216
rect 21684 4182 21715 4216
rect 21616 4126 21715 4182
rect 21616 4092 21650 4126
rect 21684 4092 21715 4126
rect 21616 4036 21715 4092
rect 21616 4002 21650 4036
rect 21684 4002 21715 4036
rect 21616 3946 21715 4002
rect 21616 3912 21650 3946
rect 21684 3912 21715 3946
rect 21616 3856 21715 3912
rect 21779 4812 22837 4831
rect 22871 4812 22910 4846
rect 21779 4778 21910 4812
rect 21944 4778 22000 4812
rect 22034 4778 22090 4812
rect 22124 4778 22180 4812
rect 22214 4778 22270 4812
rect 22304 4778 22360 4812
rect 22394 4778 22450 4812
rect 22484 4778 22540 4812
rect 22574 4778 22630 4812
rect 22664 4778 22910 4812
rect 21779 4759 22910 4778
rect 21779 4755 21851 4759
rect 21779 4721 21798 4755
rect 21832 4721 21851 4755
rect 21779 4665 21851 4721
rect 22660 4756 22910 4759
rect 22660 4736 22837 4756
rect 22660 4702 22688 4736
rect 22722 4722 22837 4736
rect 22871 4722 22910 4756
rect 22722 4702 22910 4722
rect 21779 4631 21798 4665
rect 21832 4631 21851 4665
rect 21779 4575 21851 4631
rect 21779 4541 21798 4575
rect 21832 4541 21851 4575
rect 21779 4485 21851 4541
rect 21779 4451 21798 4485
rect 21832 4451 21851 4485
rect 21779 4395 21851 4451
rect 21779 4361 21798 4395
rect 21832 4361 21851 4395
rect 21779 4305 21851 4361
rect 21779 4271 21798 4305
rect 21832 4271 21851 4305
rect 21779 4215 21851 4271
rect 21779 4181 21798 4215
rect 21832 4181 21851 4215
rect 21779 4125 21851 4181
rect 21779 4091 21798 4125
rect 21832 4091 21851 4125
rect 21779 4035 21851 4091
rect 21779 4001 21798 4035
rect 21832 4001 21851 4035
rect 21913 4638 22607 4697
rect 21913 4604 21974 4638
rect 22008 4610 22064 4638
rect 22098 4610 22154 4638
rect 22188 4610 22244 4638
rect 22020 4604 22064 4610
rect 22120 4604 22154 4610
rect 22220 4604 22244 4610
rect 22278 4610 22334 4638
rect 22278 4604 22286 4610
rect 21913 4576 21986 4604
rect 22020 4576 22086 4604
rect 22120 4576 22186 4604
rect 22220 4576 22286 4604
rect 22320 4604 22334 4610
rect 22368 4610 22424 4638
rect 22368 4604 22386 4610
rect 22320 4576 22386 4604
rect 22420 4604 22424 4610
rect 22458 4610 22514 4638
rect 22458 4604 22486 4610
rect 22548 4604 22607 4638
rect 22420 4576 22486 4604
rect 22520 4576 22607 4604
rect 21913 4548 22607 4576
rect 21913 4514 21974 4548
rect 22008 4514 22064 4548
rect 22098 4514 22154 4548
rect 22188 4514 22244 4548
rect 22278 4514 22334 4548
rect 22368 4514 22424 4548
rect 22458 4514 22514 4548
rect 22548 4514 22607 4548
rect 21913 4510 22607 4514
rect 21913 4476 21986 4510
rect 22020 4476 22086 4510
rect 22120 4476 22186 4510
rect 22220 4476 22286 4510
rect 22320 4476 22386 4510
rect 22420 4476 22486 4510
rect 22520 4476 22607 4510
rect 21913 4458 22607 4476
rect 21913 4424 21974 4458
rect 22008 4424 22064 4458
rect 22098 4424 22154 4458
rect 22188 4424 22244 4458
rect 22278 4424 22334 4458
rect 22368 4424 22424 4458
rect 22458 4424 22514 4458
rect 22548 4424 22607 4458
rect 21913 4410 22607 4424
rect 21913 4376 21986 4410
rect 22020 4376 22086 4410
rect 22120 4376 22186 4410
rect 22220 4376 22286 4410
rect 22320 4376 22386 4410
rect 22420 4376 22486 4410
rect 22520 4376 22607 4410
rect 21913 4368 22607 4376
rect 21913 4334 21974 4368
rect 22008 4334 22064 4368
rect 22098 4334 22154 4368
rect 22188 4334 22244 4368
rect 22278 4334 22334 4368
rect 22368 4334 22424 4368
rect 22458 4334 22514 4368
rect 22548 4334 22607 4368
rect 21913 4310 22607 4334
rect 21913 4278 21986 4310
rect 22020 4278 22086 4310
rect 22120 4278 22186 4310
rect 22220 4278 22286 4310
rect 21913 4244 21974 4278
rect 22020 4276 22064 4278
rect 22120 4276 22154 4278
rect 22220 4276 22244 4278
rect 22008 4244 22064 4276
rect 22098 4244 22154 4276
rect 22188 4244 22244 4276
rect 22278 4276 22286 4278
rect 22320 4278 22386 4310
rect 22320 4276 22334 4278
rect 22278 4244 22334 4276
rect 22368 4276 22386 4278
rect 22420 4278 22486 4310
rect 22520 4278 22607 4310
rect 22420 4276 22424 4278
rect 22368 4244 22424 4276
rect 22458 4276 22486 4278
rect 22458 4244 22514 4276
rect 22548 4244 22607 4278
rect 21913 4210 22607 4244
rect 21913 4188 21986 4210
rect 22020 4188 22086 4210
rect 22120 4188 22186 4210
rect 22220 4188 22286 4210
rect 21913 4154 21974 4188
rect 22020 4176 22064 4188
rect 22120 4176 22154 4188
rect 22220 4176 22244 4188
rect 22008 4154 22064 4176
rect 22098 4154 22154 4176
rect 22188 4154 22244 4176
rect 22278 4176 22286 4188
rect 22320 4188 22386 4210
rect 22320 4176 22334 4188
rect 22278 4154 22334 4176
rect 22368 4176 22386 4188
rect 22420 4188 22486 4210
rect 22520 4188 22607 4210
rect 22420 4176 22424 4188
rect 22368 4154 22424 4176
rect 22458 4176 22486 4188
rect 22458 4154 22514 4176
rect 22548 4154 22607 4188
rect 21913 4110 22607 4154
rect 21913 4098 21986 4110
rect 22020 4098 22086 4110
rect 22120 4098 22186 4110
rect 22220 4098 22286 4110
rect 21913 4064 21974 4098
rect 22020 4076 22064 4098
rect 22120 4076 22154 4098
rect 22220 4076 22244 4098
rect 22008 4064 22064 4076
rect 22098 4064 22154 4076
rect 22188 4064 22244 4076
rect 22278 4076 22286 4098
rect 22320 4098 22386 4110
rect 22320 4076 22334 4098
rect 22278 4064 22334 4076
rect 22368 4076 22386 4098
rect 22420 4098 22486 4110
rect 22520 4098 22607 4110
rect 22420 4076 22424 4098
rect 22368 4064 22424 4076
rect 22458 4076 22486 4098
rect 22458 4064 22514 4076
rect 22548 4064 22607 4098
rect 21913 4003 22607 4064
rect 22660 4666 22910 4702
rect 22660 4646 22837 4666
rect 22660 4612 22688 4646
rect 22722 4632 22837 4646
rect 22871 4632 22910 4666
rect 22722 4612 22910 4632
rect 22660 4576 22910 4612
rect 22660 4556 22837 4576
rect 22660 4522 22688 4556
rect 22722 4542 22837 4556
rect 22871 4542 22910 4576
rect 22722 4522 22910 4542
rect 22660 4486 22910 4522
rect 22660 4466 22837 4486
rect 22660 4432 22688 4466
rect 22722 4452 22837 4466
rect 22871 4452 22910 4486
rect 22722 4432 22910 4452
rect 22660 4396 22910 4432
rect 22660 4376 22837 4396
rect 22660 4342 22688 4376
rect 22722 4362 22837 4376
rect 22871 4362 22910 4396
rect 22722 4342 22910 4362
rect 22660 4306 22910 4342
rect 22660 4286 22837 4306
rect 22660 4252 22688 4286
rect 22722 4272 22837 4286
rect 22871 4272 22910 4306
rect 22722 4252 22910 4272
rect 22660 4216 22910 4252
rect 22660 4196 22837 4216
rect 22660 4162 22688 4196
rect 22722 4182 22837 4196
rect 22871 4182 22910 4216
rect 22722 4162 22910 4182
rect 22660 4126 22910 4162
rect 22660 4106 22837 4126
rect 22660 4072 22688 4106
rect 22722 4092 22837 4106
rect 22871 4092 22910 4126
rect 22722 4072 22910 4092
rect 22660 4036 22910 4072
rect 22660 4016 22837 4036
rect 21779 3941 21851 4001
rect 22660 3982 22688 4016
rect 22722 4002 22837 4016
rect 22871 4002 22910 4036
rect 22722 3982 22910 4002
rect 22660 3946 22910 3982
rect 22660 3941 22837 3946
rect 21779 3922 22837 3941
rect 21779 3888 21876 3922
rect 21910 3888 21966 3922
rect 22000 3888 22056 3922
rect 22090 3888 22146 3922
rect 22180 3888 22236 3922
rect 22270 3888 22326 3922
rect 22360 3888 22416 3922
rect 22450 3888 22506 3922
rect 22540 3888 22596 3922
rect 22630 3912 22837 3922
rect 22871 3912 22910 3946
rect 22630 3888 22910 3912
rect 21779 3869 22910 3888
rect 21616 3822 21650 3856
rect 21684 3822 21715 3856
rect 21616 3805 21715 3822
rect 22660 3856 22910 3869
rect 22660 3822 22837 3856
rect 22871 3822 22910 3856
rect 22660 3805 22910 3822
rect 21616 3772 22910 3805
rect 21616 3738 21746 3772
rect 21780 3738 21836 3772
rect 21870 3738 21926 3772
rect 21960 3738 22016 3772
rect 22050 3738 22106 3772
rect 22140 3738 22196 3772
rect 22230 3738 22286 3772
rect 22320 3738 22376 3772
rect 22410 3738 22466 3772
rect 22500 3738 22556 3772
rect 22590 3738 22646 3772
rect 22680 3738 22736 3772
rect 22770 3738 22910 3772
rect 21616 3710 22910 3738
rect 22976 4959 24270 4994
rect 22976 4936 23106 4959
rect 22976 4902 23010 4936
rect 23044 4925 23106 4936
rect 23140 4925 23196 4959
rect 23230 4925 23286 4959
rect 23320 4925 23376 4959
rect 23410 4925 23466 4959
rect 23500 4925 23556 4959
rect 23590 4925 23646 4959
rect 23680 4925 23736 4959
rect 23770 4925 23826 4959
rect 23860 4925 23916 4959
rect 23950 4925 24006 4959
rect 24040 4925 24096 4959
rect 24130 4936 24270 4959
rect 24130 4925 24197 4936
rect 23044 4902 24197 4925
rect 24231 4902 24270 4936
rect 25520 4970 25580 5030
rect 25520 4930 25530 4970
rect 25570 4930 25580 4970
rect 25520 4910 25580 4930
rect 25630 5070 25690 5090
rect 25630 5030 25640 5070
rect 25680 5030 25690 5070
rect 25630 4970 25690 5030
rect 25630 4930 25640 4970
rect 25680 4930 25690 4970
rect 25630 4910 25690 4930
rect 25740 5070 25800 5090
rect 25740 5030 25750 5070
rect 25790 5030 25800 5070
rect 25740 4970 25800 5030
rect 25740 4930 25750 4970
rect 25790 4930 25800 4970
rect 25740 4910 25800 4930
rect 22976 4895 24270 4902
rect 22976 4846 23075 4895
rect 22976 4812 23010 4846
rect 23044 4812 23075 4846
rect 24020 4846 24270 4895
rect 25530 4870 25570 4910
rect 25750 4870 25790 4910
rect 24020 4831 24197 4846
rect 22976 4756 23075 4812
rect 22976 4722 23010 4756
rect 23044 4722 23075 4756
rect 22976 4666 23075 4722
rect 22976 4632 23010 4666
rect 23044 4632 23075 4666
rect 22976 4576 23075 4632
rect 22976 4542 23010 4576
rect 23044 4542 23075 4576
rect 22976 4486 23075 4542
rect 22976 4452 23010 4486
rect 23044 4452 23075 4486
rect 22976 4396 23075 4452
rect 22976 4362 23010 4396
rect 23044 4362 23075 4396
rect 22976 4306 23075 4362
rect 22976 4272 23010 4306
rect 23044 4272 23075 4306
rect 22976 4216 23075 4272
rect 22976 4182 23010 4216
rect 23044 4182 23075 4216
rect 22976 4126 23075 4182
rect 22976 4092 23010 4126
rect 23044 4092 23075 4126
rect 22976 4036 23075 4092
rect 22976 4002 23010 4036
rect 23044 4002 23075 4036
rect 22976 3946 23075 4002
rect 22976 3912 23010 3946
rect 23044 3912 23075 3946
rect 22976 3856 23075 3912
rect 23139 4812 24197 4831
rect 24231 4812 24270 4846
rect 23139 4778 23270 4812
rect 23304 4778 23360 4812
rect 23394 4778 23450 4812
rect 23484 4778 23540 4812
rect 23574 4778 23630 4812
rect 23664 4778 23720 4812
rect 23754 4778 23810 4812
rect 23844 4778 23900 4812
rect 23934 4778 23990 4812
rect 24024 4778 24270 4812
rect 25490 4850 25570 4870
rect 25490 4810 25510 4850
rect 25550 4810 25570 4850
rect 25490 4790 25570 4810
rect 25620 4850 25700 4870
rect 25620 4810 25640 4850
rect 25680 4810 25700 4850
rect 25620 4790 25700 4810
rect 25750 4850 25830 4870
rect 25750 4810 25770 4850
rect 25810 4810 25830 4850
rect 25750 4790 25830 4810
rect 23139 4759 24270 4778
rect 23139 4755 23211 4759
rect 23139 4721 23158 4755
rect 23192 4721 23211 4755
rect 23139 4665 23211 4721
rect 24020 4756 24270 4759
rect 24020 4736 24197 4756
rect 24020 4702 24048 4736
rect 24082 4722 24197 4736
rect 24231 4722 24270 4756
rect 24082 4702 24270 4722
rect 23139 4631 23158 4665
rect 23192 4631 23211 4665
rect 23139 4575 23211 4631
rect 23139 4541 23158 4575
rect 23192 4541 23211 4575
rect 23139 4485 23211 4541
rect 23139 4451 23158 4485
rect 23192 4451 23211 4485
rect 23139 4395 23211 4451
rect 23139 4361 23158 4395
rect 23192 4361 23211 4395
rect 23139 4305 23211 4361
rect 23139 4271 23158 4305
rect 23192 4271 23211 4305
rect 23139 4215 23211 4271
rect 23139 4181 23158 4215
rect 23192 4181 23211 4215
rect 23139 4125 23211 4181
rect 23139 4091 23158 4125
rect 23192 4091 23211 4125
rect 23139 4035 23211 4091
rect 23139 4001 23158 4035
rect 23192 4001 23211 4035
rect 23273 4638 23967 4697
rect 23273 4604 23334 4638
rect 23368 4610 23424 4638
rect 23458 4610 23514 4638
rect 23548 4610 23604 4638
rect 23380 4604 23424 4610
rect 23480 4604 23514 4610
rect 23580 4604 23604 4610
rect 23638 4610 23694 4638
rect 23638 4604 23646 4610
rect 23273 4576 23346 4604
rect 23380 4576 23446 4604
rect 23480 4576 23546 4604
rect 23580 4576 23646 4604
rect 23680 4604 23694 4610
rect 23728 4610 23784 4638
rect 23728 4604 23746 4610
rect 23680 4576 23746 4604
rect 23780 4604 23784 4610
rect 23818 4610 23874 4638
rect 23818 4604 23846 4610
rect 23908 4604 23967 4638
rect 23780 4576 23846 4604
rect 23880 4576 23967 4604
rect 23273 4548 23967 4576
rect 23273 4514 23334 4548
rect 23368 4514 23424 4548
rect 23458 4514 23514 4548
rect 23548 4514 23604 4548
rect 23638 4514 23694 4548
rect 23728 4514 23784 4548
rect 23818 4514 23874 4548
rect 23908 4514 23967 4548
rect 23273 4510 23967 4514
rect 23273 4476 23346 4510
rect 23380 4476 23446 4510
rect 23480 4476 23546 4510
rect 23580 4476 23646 4510
rect 23680 4476 23746 4510
rect 23780 4476 23846 4510
rect 23880 4476 23967 4510
rect 23273 4458 23967 4476
rect 23273 4424 23334 4458
rect 23368 4424 23424 4458
rect 23458 4424 23514 4458
rect 23548 4424 23604 4458
rect 23638 4424 23694 4458
rect 23728 4424 23784 4458
rect 23818 4424 23874 4458
rect 23908 4424 23967 4458
rect 23273 4410 23967 4424
rect 23273 4376 23346 4410
rect 23380 4376 23446 4410
rect 23480 4376 23546 4410
rect 23580 4376 23646 4410
rect 23680 4376 23746 4410
rect 23780 4376 23846 4410
rect 23880 4376 23967 4410
rect 23273 4368 23967 4376
rect 23273 4334 23334 4368
rect 23368 4334 23424 4368
rect 23458 4334 23514 4368
rect 23548 4334 23604 4368
rect 23638 4334 23694 4368
rect 23728 4334 23784 4368
rect 23818 4334 23874 4368
rect 23908 4334 23967 4368
rect 23273 4310 23967 4334
rect 23273 4278 23346 4310
rect 23380 4278 23446 4310
rect 23480 4278 23546 4310
rect 23580 4278 23646 4310
rect 23273 4244 23334 4278
rect 23380 4276 23424 4278
rect 23480 4276 23514 4278
rect 23580 4276 23604 4278
rect 23368 4244 23424 4276
rect 23458 4244 23514 4276
rect 23548 4244 23604 4276
rect 23638 4276 23646 4278
rect 23680 4278 23746 4310
rect 23680 4276 23694 4278
rect 23638 4244 23694 4276
rect 23728 4276 23746 4278
rect 23780 4278 23846 4310
rect 23880 4278 23967 4310
rect 23780 4276 23784 4278
rect 23728 4244 23784 4276
rect 23818 4276 23846 4278
rect 23818 4244 23874 4276
rect 23908 4244 23967 4278
rect 23273 4210 23967 4244
rect 23273 4188 23346 4210
rect 23380 4188 23446 4210
rect 23480 4188 23546 4210
rect 23580 4188 23646 4210
rect 23273 4154 23334 4188
rect 23380 4176 23424 4188
rect 23480 4176 23514 4188
rect 23580 4176 23604 4188
rect 23368 4154 23424 4176
rect 23458 4154 23514 4176
rect 23548 4154 23604 4176
rect 23638 4176 23646 4188
rect 23680 4188 23746 4210
rect 23680 4176 23694 4188
rect 23638 4154 23694 4176
rect 23728 4176 23746 4188
rect 23780 4188 23846 4210
rect 23880 4188 23967 4210
rect 23780 4176 23784 4188
rect 23728 4154 23784 4176
rect 23818 4176 23846 4188
rect 23818 4154 23874 4176
rect 23908 4154 23967 4188
rect 23273 4110 23967 4154
rect 23273 4098 23346 4110
rect 23380 4098 23446 4110
rect 23480 4098 23546 4110
rect 23580 4098 23646 4110
rect 23273 4064 23334 4098
rect 23380 4076 23424 4098
rect 23480 4076 23514 4098
rect 23580 4076 23604 4098
rect 23368 4064 23424 4076
rect 23458 4064 23514 4076
rect 23548 4064 23604 4076
rect 23638 4076 23646 4098
rect 23680 4098 23746 4110
rect 23680 4076 23694 4098
rect 23638 4064 23694 4076
rect 23728 4076 23746 4098
rect 23780 4098 23846 4110
rect 23880 4098 23967 4110
rect 23780 4076 23784 4098
rect 23728 4064 23784 4076
rect 23818 4076 23846 4098
rect 23818 4064 23874 4076
rect 23908 4064 23967 4098
rect 23273 4003 23967 4064
rect 24020 4666 24270 4702
rect 24020 4646 24197 4666
rect 24020 4612 24048 4646
rect 24082 4632 24197 4646
rect 24231 4632 24270 4666
rect 24082 4612 24270 4632
rect 24020 4576 24270 4612
rect 24020 4556 24197 4576
rect 24020 4522 24048 4556
rect 24082 4542 24197 4556
rect 24231 4542 24270 4576
rect 24082 4522 24270 4542
rect 26400 4570 26440 5480
rect 26530 5440 26570 5480
rect 29770 5440 29810 5480
rect 26510 5420 26590 5440
rect 26510 5380 26530 5420
rect 26570 5380 26590 5420
rect 26510 5360 26590 5380
rect 26870 5420 26950 5440
rect 26870 5380 26890 5420
rect 26930 5380 26950 5420
rect 26870 5360 26950 5380
rect 27230 5420 27310 5440
rect 27230 5380 27250 5420
rect 27290 5380 27310 5420
rect 27230 5360 27310 5380
rect 27590 5420 27670 5440
rect 27590 5380 27610 5420
rect 27650 5380 27670 5420
rect 27590 5360 27670 5380
rect 27950 5420 28030 5440
rect 27950 5380 27970 5420
rect 28010 5380 28030 5420
rect 27950 5360 28030 5380
rect 28310 5420 28390 5440
rect 28310 5380 28330 5420
rect 28370 5380 28390 5420
rect 28310 5360 28390 5380
rect 28670 5420 28750 5440
rect 28670 5380 28690 5420
rect 28730 5380 28750 5420
rect 28670 5360 28750 5380
rect 29030 5420 29110 5440
rect 29030 5380 29050 5420
rect 29090 5380 29110 5420
rect 29030 5360 29110 5380
rect 29390 5420 29470 5440
rect 29390 5380 29410 5420
rect 29450 5380 29470 5420
rect 29390 5360 29470 5380
rect 29750 5420 29830 5440
rect 29750 5380 29770 5420
rect 29810 5380 29830 5420
rect 29750 5360 29830 5380
rect 26530 5320 26570 5360
rect 26890 5320 26930 5360
rect 27250 5320 27290 5360
rect 27610 5320 27650 5360
rect 27970 5320 28010 5360
rect 28330 5320 28370 5360
rect 28690 5320 28730 5360
rect 29050 5320 29090 5360
rect 29410 5320 29450 5360
rect 29770 5320 29810 5360
rect 26510 5300 26580 5320
rect 26510 5260 26530 5300
rect 26570 5260 26580 5300
rect 26510 5200 26580 5260
rect 26510 5160 26530 5200
rect 26570 5160 26580 5200
rect 26510 5100 26580 5160
rect 26510 5060 26530 5100
rect 26570 5060 26580 5100
rect 26510 5000 26580 5060
rect 26510 4960 26530 5000
rect 26570 4960 26580 5000
rect 26510 4900 26580 4960
rect 26510 4860 26530 4900
rect 26570 4860 26580 4900
rect 26510 4800 26580 4860
rect 26510 4760 26530 4800
rect 26570 4760 26580 4800
rect 26510 4740 26580 4760
rect 26700 5300 26760 5320
rect 26700 5260 26710 5300
rect 26750 5260 26760 5300
rect 26700 5200 26760 5260
rect 26700 5160 26710 5200
rect 26750 5160 26760 5200
rect 26700 5100 26760 5160
rect 26700 5060 26710 5100
rect 26750 5060 26760 5100
rect 26700 5000 26760 5060
rect 26700 4960 26710 5000
rect 26750 4960 26760 5000
rect 26700 4900 26760 4960
rect 26700 4860 26710 4900
rect 26750 4860 26760 4900
rect 26700 4800 26760 4860
rect 26700 4760 26710 4800
rect 26750 4760 26760 4800
rect 26700 4740 26760 4760
rect 26880 5300 26940 5320
rect 26880 5260 26890 5300
rect 26930 5260 26940 5300
rect 26880 5200 26940 5260
rect 26880 5160 26890 5200
rect 26930 5160 26940 5200
rect 26880 5100 26940 5160
rect 26880 5060 26890 5100
rect 26930 5060 26940 5100
rect 26880 5000 26940 5060
rect 26880 4960 26890 5000
rect 26930 4960 26940 5000
rect 26880 4900 26940 4960
rect 26880 4860 26890 4900
rect 26930 4860 26940 4900
rect 26880 4800 26940 4860
rect 26880 4760 26890 4800
rect 26930 4760 26940 4800
rect 26880 4740 26940 4760
rect 27060 5300 27120 5320
rect 27060 5260 27070 5300
rect 27110 5260 27120 5300
rect 27060 5200 27120 5260
rect 27060 5160 27070 5200
rect 27110 5160 27120 5200
rect 27060 5100 27120 5160
rect 27060 5060 27070 5100
rect 27110 5060 27120 5100
rect 27060 5000 27120 5060
rect 27060 4960 27070 5000
rect 27110 4960 27120 5000
rect 27060 4900 27120 4960
rect 27060 4860 27070 4900
rect 27110 4860 27120 4900
rect 27060 4800 27120 4860
rect 27060 4760 27070 4800
rect 27110 4760 27120 4800
rect 27060 4740 27120 4760
rect 27240 5300 27300 5320
rect 27240 5260 27250 5300
rect 27290 5260 27300 5300
rect 27240 5200 27300 5260
rect 27240 5160 27250 5200
rect 27290 5160 27300 5200
rect 27240 5100 27300 5160
rect 27240 5060 27250 5100
rect 27290 5060 27300 5100
rect 27240 5000 27300 5060
rect 27240 4960 27250 5000
rect 27290 4960 27300 5000
rect 27240 4900 27300 4960
rect 27240 4860 27250 4900
rect 27290 4860 27300 4900
rect 27240 4800 27300 4860
rect 27240 4760 27250 4800
rect 27290 4760 27300 4800
rect 27240 4740 27300 4760
rect 27420 5300 27480 5320
rect 27420 5260 27430 5300
rect 27470 5260 27480 5300
rect 27420 5200 27480 5260
rect 27420 5160 27430 5200
rect 27470 5160 27480 5200
rect 27420 5100 27480 5160
rect 27420 5060 27430 5100
rect 27470 5060 27480 5100
rect 27420 5000 27480 5060
rect 27420 4960 27430 5000
rect 27470 4960 27480 5000
rect 27420 4900 27480 4960
rect 27420 4860 27430 4900
rect 27470 4860 27480 4900
rect 27420 4800 27480 4860
rect 27420 4760 27430 4800
rect 27470 4760 27480 4800
rect 27420 4740 27480 4760
rect 27600 5300 27660 5320
rect 27600 5260 27610 5300
rect 27650 5260 27660 5300
rect 27600 5200 27660 5260
rect 27600 5160 27610 5200
rect 27650 5160 27660 5200
rect 27600 5100 27660 5160
rect 27600 5060 27610 5100
rect 27650 5060 27660 5100
rect 27600 5000 27660 5060
rect 27600 4960 27610 5000
rect 27650 4960 27660 5000
rect 27600 4900 27660 4960
rect 27600 4860 27610 4900
rect 27650 4860 27660 4900
rect 27600 4800 27660 4860
rect 27600 4760 27610 4800
rect 27650 4760 27660 4800
rect 27600 4740 27660 4760
rect 27780 5300 27840 5320
rect 27780 5260 27790 5300
rect 27830 5260 27840 5300
rect 27780 5200 27840 5260
rect 27780 5160 27790 5200
rect 27830 5160 27840 5200
rect 27780 5100 27840 5160
rect 27780 5060 27790 5100
rect 27830 5060 27840 5100
rect 27780 5000 27840 5060
rect 27780 4960 27790 5000
rect 27830 4960 27840 5000
rect 27780 4900 27840 4960
rect 27780 4860 27790 4900
rect 27830 4860 27840 4900
rect 27780 4800 27840 4860
rect 27780 4760 27790 4800
rect 27830 4760 27840 4800
rect 27780 4740 27840 4760
rect 27960 5300 28020 5320
rect 27960 5260 27970 5300
rect 28010 5260 28020 5300
rect 27960 5200 28020 5260
rect 27960 5160 27970 5200
rect 28010 5160 28020 5200
rect 27960 5100 28020 5160
rect 27960 5060 27970 5100
rect 28010 5060 28020 5100
rect 27960 5000 28020 5060
rect 27960 4960 27970 5000
rect 28010 4960 28020 5000
rect 27960 4900 28020 4960
rect 27960 4860 27970 4900
rect 28010 4860 28020 4900
rect 27960 4800 28020 4860
rect 27960 4760 27970 4800
rect 28010 4760 28020 4800
rect 27960 4740 28020 4760
rect 28140 5300 28200 5320
rect 28140 5260 28150 5300
rect 28190 5260 28200 5300
rect 28140 5200 28200 5260
rect 28140 5160 28150 5200
rect 28190 5160 28200 5200
rect 28140 5100 28200 5160
rect 28140 5060 28150 5100
rect 28190 5060 28200 5100
rect 28140 5000 28200 5060
rect 28140 4960 28150 5000
rect 28190 4960 28200 5000
rect 28140 4900 28200 4960
rect 28140 4860 28150 4900
rect 28190 4860 28200 4900
rect 28140 4800 28200 4860
rect 28140 4760 28150 4800
rect 28190 4760 28200 4800
rect 28140 4740 28200 4760
rect 28320 5300 28380 5320
rect 28320 5260 28330 5300
rect 28370 5260 28380 5300
rect 28320 5200 28380 5260
rect 28320 5160 28330 5200
rect 28370 5160 28380 5200
rect 28320 5100 28380 5160
rect 28320 5060 28330 5100
rect 28370 5060 28380 5100
rect 28320 5000 28380 5060
rect 28320 4960 28330 5000
rect 28370 4960 28380 5000
rect 28320 4900 28380 4960
rect 28320 4860 28330 4900
rect 28370 4860 28380 4900
rect 28320 4800 28380 4860
rect 28320 4760 28330 4800
rect 28370 4760 28380 4800
rect 28320 4740 28380 4760
rect 28500 5300 28560 5320
rect 28500 5260 28510 5300
rect 28550 5260 28560 5300
rect 28500 5200 28560 5260
rect 28500 5160 28510 5200
rect 28550 5160 28560 5200
rect 28500 5100 28560 5160
rect 28500 5060 28510 5100
rect 28550 5060 28560 5100
rect 28500 5000 28560 5060
rect 28500 4960 28510 5000
rect 28550 4960 28560 5000
rect 28500 4900 28560 4960
rect 28500 4860 28510 4900
rect 28550 4860 28560 4900
rect 28500 4800 28560 4860
rect 28500 4760 28510 4800
rect 28550 4760 28560 4800
rect 28500 4740 28560 4760
rect 28680 5300 28740 5320
rect 28680 5260 28690 5300
rect 28730 5260 28740 5300
rect 28680 5200 28740 5260
rect 28680 5160 28690 5200
rect 28730 5160 28740 5200
rect 28680 5100 28740 5160
rect 28680 5060 28690 5100
rect 28730 5060 28740 5100
rect 28680 5000 28740 5060
rect 28680 4960 28690 5000
rect 28730 4960 28740 5000
rect 28680 4900 28740 4960
rect 28680 4860 28690 4900
rect 28730 4860 28740 4900
rect 28680 4800 28740 4860
rect 28680 4760 28690 4800
rect 28730 4760 28740 4800
rect 28680 4740 28740 4760
rect 28860 5300 28920 5320
rect 28860 5260 28870 5300
rect 28910 5260 28920 5300
rect 28860 5200 28920 5260
rect 28860 5160 28870 5200
rect 28910 5160 28920 5200
rect 28860 5100 28920 5160
rect 28860 5060 28870 5100
rect 28910 5060 28920 5100
rect 28860 5000 28920 5060
rect 28860 4960 28870 5000
rect 28910 4960 28920 5000
rect 28860 4900 28920 4960
rect 28860 4860 28870 4900
rect 28910 4860 28920 4900
rect 28860 4800 28920 4860
rect 28860 4760 28870 4800
rect 28910 4760 28920 4800
rect 28860 4740 28920 4760
rect 29040 5300 29100 5320
rect 29040 5260 29050 5300
rect 29090 5260 29100 5300
rect 29040 5200 29100 5260
rect 29040 5160 29050 5200
rect 29090 5160 29100 5200
rect 29040 5100 29100 5160
rect 29040 5060 29050 5100
rect 29090 5060 29100 5100
rect 29040 5000 29100 5060
rect 29040 4960 29050 5000
rect 29090 4960 29100 5000
rect 29040 4900 29100 4960
rect 29040 4860 29050 4900
rect 29090 4860 29100 4900
rect 29040 4800 29100 4860
rect 29040 4760 29050 4800
rect 29090 4760 29100 4800
rect 29040 4740 29100 4760
rect 29220 5300 29280 5320
rect 29220 5260 29230 5300
rect 29270 5260 29280 5300
rect 29220 5200 29280 5260
rect 29220 5160 29230 5200
rect 29270 5160 29280 5200
rect 29220 5100 29280 5160
rect 29220 5060 29230 5100
rect 29270 5060 29280 5100
rect 29220 5000 29280 5060
rect 29220 4960 29230 5000
rect 29270 4960 29280 5000
rect 29220 4900 29280 4960
rect 29220 4860 29230 4900
rect 29270 4860 29280 4900
rect 29220 4800 29280 4860
rect 29220 4760 29230 4800
rect 29270 4760 29280 4800
rect 29220 4740 29280 4760
rect 29400 5300 29460 5320
rect 29400 5260 29410 5300
rect 29450 5260 29460 5300
rect 29400 5200 29460 5260
rect 29400 5160 29410 5200
rect 29450 5160 29460 5200
rect 29400 5100 29460 5160
rect 29400 5060 29410 5100
rect 29450 5060 29460 5100
rect 29400 5000 29460 5060
rect 29400 4960 29410 5000
rect 29450 4960 29460 5000
rect 29400 4900 29460 4960
rect 29400 4860 29410 4900
rect 29450 4860 29460 4900
rect 29400 4800 29460 4860
rect 29400 4760 29410 4800
rect 29450 4760 29460 4800
rect 29400 4740 29460 4760
rect 29580 5300 29640 5320
rect 29580 5260 29590 5300
rect 29630 5260 29640 5300
rect 29580 5200 29640 5260
rect 29580 5160 29590 5200
rect 29630 5160 29640 5200
rect 29580 5100 29640 5160
rect 29580 5060 29590 5100
rect 29630 5060 29640 5100
rect 29580 5000 29640 5060
rect 29580 4960 29590 5000
rect 29630 4960 29640 5000
rect 29580 4900 29640 4960
rect 29580 4860 29590 4900
rect 29630 4860 29640 4900
rect 29580 4800 29640 4860
rect 29580 4760 29590 4800
rect 29630 4760 29640 4800
rect 29580 4740 29640 4760
rect 29760 5300 29820 5320
rect 29760 5260 29770 5300
rect 29810 5260 29820 5300
rect 29760 5200 29820 5260
rect 29760 5160 29770 5200
rect 29810 5160 29820 5200
rect 29760 5100 29820 5160
rect 29760 5060 29770 5100
rect 29810 5060 29820 5100
rect 29760 5000 29820 5060
rect 29760 4960 29770 5000
rect 29810 4960 29820 5000
rect 29760 4900 29820 4960
rect 29760 4860 29770 4900
rect 29810 4860 29820 4900
rect 29760 4800 29820 4860
rect 29760 4760 29770 4800
rect 29810 4760 29820 4800
rect 29760 4740 29820 4760
rect 26710 4700 26750 4740
rect 27070 4700 27110 4740
rect 27430 4700 27470 4740
rect 27790 4700 27830 4740
rect 28150 4700 28190 4740
rect 28510 4700 28550 4740
rect 28870 4700 28910 4740
rect 29230 4700 29270 4740
rect 29590 4700 29630 4740
rect 26690 4680 26770 4700
rect 26690 4640 26710 4680
rect 26750 4640 26770 4680
rect 26690 4620 26770 4640
rect 27050 4680 27130 4700
rect 27050 4640 27070 4680
rect 27110 4640 27130 4680
rect 27050 4620 27130 4640
rect 27410 4680 27490 4700
rect 27410 4640 27430 4680
rect 27470 4640 27490 4680
rect 27410 4620 27490 4640
rect 27650 4680 27730 4700
rect 27650 4640 27670 4680
rect 27710 4640 27730 4680
rect 27650 4620 27730 4640
rect 27770 4680 27850 4700
rect 27770 4640 27790 4680
rect 27830 4640 27850 4680
rect 27770 4620 27850 4640
rect 28130 4680 28210 4700
rect 28130 4640 28150 4680
rect 28190 4640 28210 4680
rect 28130 4620 28210 4640
rect 28490 4680 28570 4700
rect 28490 4640 28510 4680
rect 28550 4640 28570 4680
rect 28490 4620 28570 4640
rect 28850 4680 28930 4700
rect 28850 4640 28870 4680
rect 28910 4640 28930 4680
rect 28850 4620 28930 4640
rect 29210 4680 29290 4700
rect 29210 4640 29230 4680
rect 29270 4640 29290 4680
rect 29210 4620 29290 4640
rect 29390 4680 29470 4700
rect 29390 4640 29410 4680
rect 29450 4640 29470 4680
rect 29390 4620 29470 4640
rect 29570 4680 29650 4700
rect 29570 4640 29590 4680
rect 29630 4640 29650 4680
rect 29570 4620 29650 4640
rect 29890 4570 29930 5480
rect 26400 4530 29930 4570
rect 24020 4486 24270 4522
rect 24020 4466 24197 4486
rect 24020 4432 24048 4466
rect 24082 4452 24197 4466
rect 24231 4452 24270 4486
rect 24082 4432 24270 4452
rect 24020 4396 24270 4432
rect 24020 4376 24197 4396
rect 24020 4342 24048 4376
rect 24082 4362 24197 4376
rect 24231 4362 24270 4396
rect 24082 4342 24270 4362
rect 24020 4306 24270 4342
rect 24020 4286 24197 4306
rect 24020 4252 24048 4286
rect 24082 4272 24197 4286
rect 24231 4272 24270 4306
rect 24082 4252 24270 4272
rect 24020 4216 24270 4252
rect 24020 4196 24197 4216
rect 24020 4162 24048 4196
rect 24082 4182 24197 4196
rect 24231 4182 24270 4216
rect 28690 4210 28770 4230
rect 28690 4190 28710 4210
rect 24082 4162 24270 4182
rect 24020 4126 24270 4162
rect 24020 4106 24197 4126
rect 24020 4072 24048 4106
rect 24082 4092 24197 4106
rect 24231 4092 24270 4126
rect 24082 4072 24270 4092
rect 24020 4036 24270 4072
rect 24020 4016 24197 4036
rect 23139 3941 23211 4001
rect 24020 3982 24048 4016
rect 24082 4002 24197 4016
rect 24231 4002 24270 4036
rect 24082 3982 24270 4002
rect 24020 3946 24270 3982
rect 24020 3941 24197 3946
rect 23139 3922 24197 3941
rect 23139 3888 23236 3922
rect 23270 3888 23326 3922
rect 23360 3888 23416 3922
rect 23450 3888 23506 3922
rect 23540 3888 23596 3922
rect 23630 3888 23686 3922
rect 23720 3888 23776 3922
rect 23810 3888 23866 3922
rect 23900 3888 23956 3922
rect 23990 3912 24197 3922
rect 24231 3912 24270 3946
rect 23990 3888 24270 3912
rect 23139 3869 24270 3888
rect 22976 3822 23010 3856
rect 23044 3822 23075 3856
rect 22976 3805 23075 3822
rect 24020 3856 24270 3869
rect 24020 3822 24197 3856
rect 24231 3822 24270 3856
rect 24020 3805 24270 3822
rect 22976 3772 24270 3805
rect 22976 3738 23106 3772
rect 23140 3738 23196 3772
rect 23230 3738 23286 3772
rect 23320 3738 23376 3772
rect 23410 3738 23466 3772
rect 23500 3738 23556 3772
rect 23590 3738 23646 3772
rect 23680 3738 23736 3772
rect 23770 3738 23826 3772
rect 23860 3738 23916 3772
rect 23950 3738 24006 3772
rect 24040 3738 24096 3772
rect 24130 3738 24270 3772
rect 22976 3710 24270 3738
rect 20250 3630 24270 3710
rect 20256 3599 21550 3630
rect 20256 3576 20386 3599
rect 20256 3542 20290 3576
rect 20324 3565 20386 3576
rect 20420 3565 20476 3599
rect 20510 3565 20566 3599
rect 20600 3565 20656 3599
rect 20690 3565 20746 3599
rect 20780 3565 20836 3599
rect 20870 3565 20926 3599
rect 20960 3565 21016 3599
rect 21050 3565 21106 3599
rect 21140 3565 21196 3599
rect 21230 3565 21286 3599
rect 21320 3565 21376 3599
rect 21410 3576 21550 3599
rect 21410 3565 21477 3576
rect 20324 3542 21477 3565
rect 21511 3542 21550 3576
rect 20256 3535 21550 3542
rect 20256 3486 20355 3535
rect 20256 3452 20290 3486
rect 20324 3452 20355 3486
rect 21300 3486 21550 3535
rect 21300 3471 21477 3486
rect 20256 3396 20355 3452
rect 20256 3362 20290 3396
rect 20324 3362 20355 3396
rect 20256 3306 20355 3362
rect 20256 3272 20290 3306
rect 20324 3272 20355 3306
rect 20256 3216 20355 3272
rect 20256 3182 20290 3216
rect 20324 3182 20355 3216
rect 20256 3126 20355 3182
rect 20256 3092 20290 3126
rect 20324 3092 20355 3126
rect 20256 3050 20355 3092
rect 19910 3036 20355 3050
rect 19910 3030 20290 3036
rect 19910 2990 19930 3030
rect 19970 2990 20030 3030
rect 20070 2990 20130 3030
rect 20170 3002 20290 3030
rect 20324 3002 20355 3036
rect 20170 2990 20355 3002
rect 19910 2970 20355 2990
rect 20256 2946 20355 2970
rect 20256 2912 20290 2946
rect 20324 2912 20355 2946
rect 20256 2856 20355 2912
rect 20256 2822 20290 2856
rect 20324 2822 20355 2856
rect 20256 2766 20355 2822
rect 20256 2732 20290 2766
rect 20324 2732 20355 2766
rect 20256 2676 20355 2732
rect 20256 2642 20290 2676
rect 20324 2642 20355 2676
rect 20256 2586 20355 2642
rect 20256 2552 20290 2586
rect 20324 2552 20355 2586
rect 20256 2496 20355 2552
rect 20419 3452 21477 3471
rect 21511 3452 21550 3486
rect 20419 3418 20550 3452
rect 20584 3418 20640 3452
rect 20674 3418 20730 3452
rect 20764 3418 20820 3452
rect 20854 3418 20910 3452
rect 20944 3418 21000 3452
rect 21034 3418 21090 3452
rect 21124 3418 21180 3452
rect 21214 3418 21270 3452
rect 21304 3418 21550 3452
rect 20419 3399 21550 3418
rect 20419 3395 20491 3399
rect 20419 3361 20438 3395
rect 20472 3361 20491 3395
rect 20419 3305 20491 3361
rect 21300 3396 21550 3399
rect 21300 3376 21477 3396
rect 21300 3342 21328 3376
rect 21362 3362 21477 3376
rect 21511 3362 21550 3396
rect 21362 3342 21550 3362
rect 20419 3271 20438 3305
rect 20472 3271 20491 3305
rect 20419 3215 20491 3271
rect 20419 3181 20438 3215
rect 20472 3181 20491 3215
rect 20419 3125 20491 3181
rect 20419 3091 20438 3125
rect 20472 3091 20491 3125
rect 20419 3035 20491 3091
rect 20419 3001 20438 3035
rect 20472 3001 20491 3035
rect 20419 2945 20491 3001
rect 20419 2911 20438 2945
rect 20472 2911 20491 2945
rect 20419 2855 20491 2911
rect 20419 2821 20438 2855
rect 20472 2821 20491 2855
rect 20419 2765 20491 2821
rect 20419 2731 20438 2765
rect 20472 2731 20491 2765
rect 20419 2675 20491 2731
rect 20419 2641 20438 2675
rect 20472 2641 20491 2675
rect 20553 3278 21247 3337
rect 20553 3244 20614 3278
rect 20648 3250 20704 3278
rect 20738 3250 20794 3278
rect 20828 3250 20884 3278
rect 20660 3244 20704 3250
rect 20760 3244 20794 3250
rect 20860 3244 20884 3250
rect 20918 3250 20974 3278
rect 20918 3244 20926 3250
rect 20553 3216 20626 3244
rect 20660 3216 20726 3244
rect 20760 3216 20826 3244
rect 20860 3216 20926 3244
rect 20960 3244 20974 3250
rect 21008 3250 21064 3278
rect 21008 3244 21026 3250
rect 20960 3216 21026 3244
rect 21060 3244 21064 3250
rect 21098 3250 21154 3278
rect 21098 3244 21126 3250
rect 21188 3244 21247 3278
rect 21060 3216 21126 3244
rect 21160 3216 21247 3244
rect 20553 3188 21247 3216
rect 20553 3154 20614 3188
rect 20648 3154 20704 3188
rect 20738 3154 20794 3188
rect 20828 3154 20884 3188
rect 20918 3154 20974 3188
rect 21008 3154 21064 3188
rect 21098 3154 21154 3188
rect 21188 3154 21247 3188
rect 20553 3150 21247 3154
rect 20553 3116 20626 3150
rect 20660 3116 20726 3150
rect 20760 3116 20826 3150
rect 20860 3116 20926 3150
rect 20960 3116 21026 3150
rect 21060 3116 21126 3150
rect 21160 3116 21247 3150
rect 20553 3098 21247 3116
rect 20553 3064 20614 3098
rect 20648 3064 20704 3098
rect 20738 3064 20794 3098
rect 20828 3064 20884 3098
rect 20918 3064 20974 3098
rect 21008 3064 21064 3098
rect 21098 3064 21154 3098
rect 21188 3064 21247 3098
rect 20553 3050 21247 3064
rect 20553 3016 20626 3050
rect 20660 3016 20726 3050
rect 20760 3016 20826 3050
rect 20860 3016 20926 3050
rect 20960 3016 21026 3050
rect 21060 3016 21126 3050
rect 21160 3016 21247 3050
rect 20553 3008 21247 3016
rect 20553 2974 20614 3008
rect 20648 2974 20704 3008
rect 20738 2974 20794 3008
rect 20828 2974 20884 3008
rect 20918 2974 20974 3008
rect 21008 2974 21064 3008
rect 21098 2974 21154 3008
rect 21188 2974 21247 3008
rect 20553 2950 21247 2974
rect 20553 2918 20626 2950
rect 20660 2918 20726 2950
rect 20760 2918 20826 2950
rect 20860 2918 20926 2950
rect 20553 2884 20614 2918
rect 20660 2916 20704 2918
rect 20760 2916 20794 2918
rect 20860 2916 20884 2918
rect 20648 2884 20704 2916
rect 20738 2884 20794 2916
rect 20828 2884 20884 2916
rect 20918 2916 20926 2918
rect 20960 2918 21026 2950
rect 20960 2916 20974 2918
rect 20918 2884 20974 2916
rect 21008 2916 21026 2918
rect 21060 2918 21126 2950
rect 21160 2918 21247 2950
rect 21060 2916 21064 2918
rect 21008 2884 21064 2916
rect 21098 2916 21126 2918
rect 21098 2884 21154 2916
rect 21188 2884 21247 2918
rect 20553 2850 21247 2884
rect 20553 2828 20626 2850
rect 20660 2828 20726 2850
rect 20760 2828 20826 2850
rect 20860 2828 20926 2850
rect 20553 2794 20614 2828
rect 20660 2816 20704 2828
rect 20760 2816 20794 2828
rect 20860 2816 20884 2828
rect 20648 2794 20704 2816
rect 20738 2794 20794 2816
rect 20828 2794 20884 2816
rect 20918 2816 20926 2828
rect 20960 2828 21026 2850
rect 20960 2816 20974 2828
rect 20918 2794 20974 2816
rect 21008 2816 21026 2828
rect 21060 2828 21126 2850
rect 21160 2828 21247 2850
rect 21060 2816 21064 2828
rect 21008 2794 21064 2816
rect 21098 2816 21126 2828
rect 21098 2794 21154 2816
rect 21188 2794 21247 2828
rect 20553 2750 21247 2794
rect 20553 2738 20626 2750
rect 20660 2738 20726 2750
rect 20760 2738 20826 2750
rect 20860 2738 20926 2750
rect 20553 2704 20614 2738
rect 20660 2716 20704 2738
rect 20760 2716 20794 2738
rect 20860 2716 20884 2738
rect 20648 2704 20704 2716
rect 20738 2704 20794 2716
rect 20828 2704 20884 2716
rect 20918 2716 20926 2738
rect 20960 2738 21026 2750
rect 20960 2716 20974 2738
rect 20918 2704 20974 2716
rect 21008 2716 21026 2738
rect 21060 2738 21126 2750
rect 21160 2738 21247 2750
rect 21060 2716 21064 2738
rect 21008 2704 21064 2716
rect 21098 2716 21126 2738
rect 21098 2704 21154 2716
rect 21188 2704 21247 2738
rect 20553 2643 21247 2704
rect 21300 3306 21550 3342
rect 21300 3286 21477 3306
rect 21300 3252 21328 3286
rect 21362 3272 21477 3286
rect 21511 3272 21550 3306
rect 21362 3252 21550 3272
rect 21300 3216 21550 3252
rect 21300 3196 21477 3216
rect 21300 3162 21328 3196
rect 21362 3182 21477 3196
rect 21511 3182 21550 3216
rect 21362 3162 21550 3182
rect 21300 3126 21550 3162
rect 21300 3106 21477 3126
rect 21300 3072 21328 3106
rect 21362 3092 21477 3106
rect 21511 3092 21550 3126
rect 21362 3072 21550 3092
rect 21300 3036 21550 3072
rect 21300 3016 21477 3036
rect 21300 2982 21328 3016
rect 21362 3002 21477 3016
rect 21511 3002 21550 3036
rect 21362 2982 21550 3002
rect 21300 2946 21550 2982
rect 21300 2926 21477 2946
rect 21300 2892 21328 2926
rect 21362 2912 21477 2926
rect 21511 2912 21550 2946
rect 21362 2892 21550 2912
rect 21300 2856 21550 2892
rect 21300 2836 21477 2856
rect 21300 2802 21328 2836
rect 21362 2822 21477 2836
rect 21511 2822 21550 2856
rect 21362 2802 21550 2822
rect 21300 2766 21550 2802
rect 21300 2746 21477 2766
rect 21300 2712 21328 2746
rect 21362 2732 21477 2746
rect 21511 2732 21550 2766
rect 21362 2712 21550 2732
rect 21300 2676 21550 2712
rect 21300 2656 21477 2676
rect 20419 2581 20491 2641
rect 21300 2622 21328 2656
rect 21362 2642 21477 2656
rect 21511 2642 21550 2676
rect 21362 2622 21550 2642
rect 21300 2586 21550 2622
rect 21300 2581 21477 2586
rect 20419 2562 21477 2581
rect 20419 2528 20516 2562
rect 20550 2528 20606 2562
rect 20640 2528 20696 2562
rect 20730 2528 20786 2562
rect 20820 2528 20876 2562
rect 20910 2528 20966 2562
rect 21000 2528 21056 2562
rect 21090 2528 21146 2562
rect 21180 2528 21236 2562
rect 21270 2552 21477 2562
rect 21511 2552 21550 2586
rect 21270 2528 21550 2552
rect 20419 2509 21550 2528
rect 20256 2462 20290 2496
rect 20324 2462 20355 2496
rect 20256 2445 20355 2462
rect 21300 2496 21550 2509
rect 21300 2462 21477 2496
rect 21511 2462 21550 2496
rect 21300 2445 21550 2462
rect 20256 2412 21550 2445
rect 20256 2378 20386 2412
rect 20420 2378 20476 2412
rect 20510 2378 20566 2412
rect 20600 2378 20656 2412
rect 20690 2378 20746 2412
rect 20780 2378 20836 2412
rect 20870 2378 20926 2412
rect 20960 2378 21016 2412
rect 21050 2378 21106 2412
rect 21140 2378 21196 2412
rect 21230 2378 21286 2412
rect 21320 2378 21376 2412
rect 21410 2378 21550 2412
rect 20256 2350 21550 2378
rect 21616 3599 22910 3630
rect 21616 3576 21746 3599
rect 21616 3542 21650 3576
rect 21684 3565 21746 3576
rect 21780 3565 21836 3599
rect 21870 3565 21926 3599
rect 21960 3565 22016 3599
rect 22050 3565 22106 3599
rect 22140 3565 22196 3599
rect 22230 3565 22286 3599
rect 22320 3565 22376 3599
rect 22410 3565 22466 3599
rect 22500 3565 22556 3599
rect 22590 3565 22646 3599
rect 22680 3565 22736 3599
rect 22770 3576 22910 3599
rect 22770 3565 22837 3576
rect 21684 3542 22837 3565
rect 22871 3542 22910 3576
rect 21616 3535 22910 3542
rect 21616 3486 21715 3535
rect 21616 3452 21650 3486
rect 21684 3452 21715 3486
rect 22660 3486 22910 3535
rect 22660 3471 22837 3486
rect 21616 3396 21715 3452
rect 21616 3362 21650 3396
rect 21684 3362 21715 3396
rect 21616 3306 21715 3362
rect 21616 3272 21650 3306
rect 21684 3272 21715 3306
rect 21616 3216 21715 3272
rect 21616 3182 21650 3216
rect 21684 3182 21715 3216
rect 21616 3126 21715 3182
rect 21616 3092 21650 3126
rect 21684 3092 21715 3126
rect 21616 3036 21715 3092
rect 21616 3002 21650 3036
rect 21684 3002 21715 3036
rect 21616 2946 21715 3002
rect 21616 2912 21650 2946
rect 21684 2912 21715 2946
rect 21616 2856 21715 2912
rect 21616 2822 21650 2856
rect 21684 2822 21715 2856
rect 21616 2766 21715 2822
rect 21616 2732 21650 2766
rect 21684 2732 21715 2766
rect 21616 2676 21715 2732
rect 21616 2642 21650 2676
rect 21684 2642 21715 2676
rect 21616 2586 21715 2642
rect 21616 2552 21650 2586
rect 21684 2552 21715 2586
rect 21616 2496 21715 2552
rect 21779 3452 22837 3471
rect 22871 3452 22910 3486
rect 21779 3418 21910 3452
rect 21944 3418 22000 3452
rect 22034 3418 22090 3452
rect 22124 3418 22180 3452
rect 22214 3418 22270 3452
rect 22304 3418 22360 3452
rect 22394 3418 22450 3452
rect 22484 3418 22540 3452
rect 22574 3418 22630 3452
rect 22664 3418 22910 3452
rect 21779 3399 22910 3418
rect 21779 3395 21851 3399
rect 21779 3361 21798 3395
rect 21832 3361 21851 3395
rect 21779 3305 21851 3361
rect 22660 3396 22910 3399
rect 22660 3376 22837 3396
rect 22660 3342 22688 3376
rect 22722 3362 22837 3376
rect 22871 3362 22910 3396
rect 22722 3342 22910 3362
rect 21779 3271 21798 3305
rect 21832 3271 21851 3305
rect 21779 3215 21851 3271
rect 21779 3181 21798 3215
rect 21832 3181 21851 3215
rect 21779 3125 21851 3181
rect 21779 3091 21798 3125
rect 21832 3091 21851 3125
rect 21779 3035 21851 3091
rect 21779 3001 21798 3035
rect 21832 3001 21851 3035
rect 21779 2945 21851 3001
rect 21779 2911 21798 2945
rect 21832 2911 21851 2945
rect 21779 2855 21851 2911
rect 21779 2821 21798 2855
rect 21832 2821 21851 2855
rect 21779 2765 21851 2821
rect 21779 2731 21798 2765
rect 21832 2731 21851 2765
rect 21779 2675 21851 2731
rect 21779 2641 21798 2675
rect 21832 2641 21851 2675
rect 21913 3278 22607 3337
rect 21913 3244 21974 3278
rect 22008 3250 22064 3278
rect 22098 3250 22154 3278
rect 22188 3250 22244 3278
rect 22020 3244 22064 3250
rect 22120 3244 22154 3250
rect 22220 3244 22244 3250
rect 22278 3250 22334 3278
rect 22278 3244 22286 3250
rect 21913 3216 21986 3244
rect 22020 3216 22086 3244
rect 22120 3216 22186 3244
rect 22220 3216 22286 3244
rect 22320 3244 22334 3250
rect 22368 3250 22424 3278
rect 22368 3244 22386 3250
rect 22320 3216 22386 3244
rect 22420 3244 22424 3250
rect 22458 3250 22514 3278
rect 22458 3244 22486 3250
rect 22548 3244 22607 3278
rect 22420 3216 22486 3244
rect 22520 3216 22607 3244
rect 21913 3188 22607 3216
rect 21913 3154 21974 3188
rect 22008 3154 22064 3188
rect 22098 3154 22154 3188
rect 22188 3154 22244 3188
rect 22278 3154 22334 3188
rect 22368 3154 22424 3188
rect 22458 3154 22514 3188
rect 22548 3154 22607 3188
rect 21913 3150 22607 3154
rect 21913 3116 21986 3150
rect 22020 3116 22086 3150
rect 22120 3116 22186 3150
rect 22220 3116 22286 3150
rect 22320 3116 22386 3150
rect 22420 3116 22486 3150
rect 22520 3116 22607 3150
rect 21913 3098 22607 3116
rect 21913 3064 21974 3098
rect 22008 3064 22064 3098
rect 22098 3064 22154 3098
rect 22188 3064 22244 3098
rect 22278 3064 22334 3098
rect 22368 3064 22424 3098
rect 22458 3064 22514 3098
rect 22548 3064 22607 3098
rect 21913 3050 22607 3064
rect 21913 3016 21986 3050
rect 22020 3016 22086 3050
rect 22120 3016 22186 3050
rect 22220 3016 22286 3050
rect 22320 3016 22386 3050
rect 22420 3016 22486 3050
rect 22520 3016 22607 3050
rect 21913 3008 22607 3016
rect 21913 2974 21974 3008
rect 22008 2974 22064 3008
rect 22098 2974 22154 3008
rect 22188 2974 22244 3008
rect 22278 2974 22334 3008
rect 22368 2974 22424 3008
rect 22458 2974 22514 3008
rect 22548 2974 22607 3008
rect 21913 2950 22607 2974
rect 21913 2918 21986 2950
rect 22020 2918 22086 2950
rect 22120 2918 22186 2950
rect 22220 2918 22286 2950
rect 21913 2884 21974 2918
rect 22020 2916 22064 2918
rect 22120 2916 22154 2918
rect 22220 2916 22244 2918
rect 22008 2884 22064 2916
rect 22098 2884 22154 2916
rect 22188 2884 22244 2916
rect 22278 2916 22286 2918
rect 22320 2918 22386 2950
rect 22320 2916 22334 2918
rect 22278 2884 22334 2916
rect 22368 2916 22386 2918
rect 22420 2918 22486 2950
rect 22520 2918 22607 2950
rect 22420 2916 22424 2918
rect 22368 2884 22424 2916
rect 22458 2916 22486 2918
rect 22458 2884 22514 2916
rect 22548 2884 22607 2918
rect 21913 2850 22607 2884
rect 21913 2828 21986 2850
rect 22020 2828 22086 2850
rect 22120 2828 22186 2850
rect 22220 2828 22286 2850
rect 21913 2794 21974 2828
rect 22020 2816 22064 2828
rect 22120 2816 22154 2828
rect 22220 2816 22244 2828
rect 22008 2794 22064 2816
rect 22098 2794 22154 2816
rect 22188 2794 22244 2816
rect 22278 2816 22286 2828
rect 22320 2828 22386 2850
rect 22320 2816 22334 2828
rect 22278 2794 22334 2816
rect 22368 2816 22386 2828
rect 22420 2828 22486 2850
rect 22520 2828 22607 2850
rect 22420 2816 22424 2828
rect 22368 2794 22424 2816
rect 22458 2816 22486 2828
rect 22458 2794 22514 2816
rect 22548 2794 22607 2828
rect 21913 2750 22607 2794
rect 21913 2738 21986 2750
rect 22020 2738 22086 2750
rect 22120 2738 22186 2750
rect 22220 2738 22286 2750
rect 21913 2704 21974 2738
rect 22020 2716 22064 2738
rect 22120 2716 22154 2738
rect 22220 2716 22244 2738
rect 22008 2704 22064 2716
rect 22098 2704 22154 2716
rect 22188 2704 22244 2716
rect 22278 2716 22286 2738
rect 22320 2738 22386 2750
rect 22320 2716 22334 2738
rect 22278 2704 22334 2716
rect 22368 2716 22386 2738
rect 22420 2738 22486 2750
rect 22520 2738 22607 2750
rect 22420 2716 22424 2738
rect 22368 2704 22424 2716
rect 22458 2716 22486 2738
rect 22458 2704 22514 2716
rect 22548 2704 22607 2738
rect 21913 2643 22607 2704
rect 22660 3306 22910 3342
rect 22660 3286 22837 3306
rect 22660 3252 22688 3286
rect 22722 3272 22837 3286
rect 22871 3272 22910 3306
rect 22722 3252 22910 3272
rect 22660 3216 22910 3252
rect 22660 3196 22837 3216
rect 22660 3162 22688 3196
rect 22722 3182 22837 3196
rect 22871 3182 22910 3216
rect 22722 3162 22910 3182
rect 22660 3126 22910 3162
rect 22660 3106 22837 3126
rect 22660 3072 22688 3106
rect 22722 3092 22837 3106
rect 22871 3092 22910 3126
rect 22722 3072 22910 3092
rect 22660 3036 22910 3072
rect 22660 3016 22837 3036
rect 22660 2982 22688 3016
rect 22722 3002 22837 3016
rect 22871 3002 22910 3036
rect 22722 2982 22910 3002
rect 22660 2946 22910 2982
rect 22660 2926 22837 2946
rect 22660 2892 22688 2926
rect 22722 2912 22837 2926
rect 22871 2912 22910 2946
rect 22722 2892 22910 2912
rect 22660 2856 22910 2892
rect 22660 2836 22837 2856
rect 22660 2802 22688 2836
rect 22722 2822 22837 2836
rect 22871 2822 22910 2856
rect 22722 2802 22910 2822
rect 22660 2766 22910 2802
rect 22660 2746 22837 2766
rect 22660 2712 22688 2746
rect 22722 2732 22837 2746
rect 22871 2732 22910 2766
rect 22722 2712 22910 2732
rect 22660 2676 22910 2712
rect 22660 2656 22837 2676
rect 21779 2581 21851 2641
rect 22660 2622 22688 2656
rect 22722 2642 22837 2656
rect 22871 2642 22910 2676
rect 22722 2622 22910 2642
rect 22660 2586 22910 2622
rect 22660 2581 22837 2586
rect 21779 2562 22837 2581
rect 21779 2528 21876 2562
rect 21910 2528 21966 2562
rect 22000 2528 22056 2562
rect 22090 2528 22146 2562
rect 22180 2528 22236 2562
rect 22270 2528 22326 2562
rect 22360 2528 22416 2562
rect 22450 2528 22506 2562
rect 22540 2528 22596 2562
rect 22630 2552 22837 2562
rect 22871 2552 22910 2586
rect 22630 2528 22910 2552
rect 21779 2509 22910 2528
rect 21616 2462 21650 2496
rect 21684 2462 21715 2496
rect 21616 2445 21715 2462
rect 22660 2496 22910 2509
rect 22660 2462 22837 2496
rect 22871 2462 22910 2496
rect 22660 2445 22910 2462
rect 21616 2412 22910 2445
rect 21616 2378 21746 2412
rect 21780 2378 21836 2412
rect 21870 2378 21926 2412
rect 21960 2378 22016 2412
rect 22050 2378 22106 2412
rect 22140 2378 22196 2412
rect 22230 2378 22286 2412
rect 22320 2378 22376 2412
rect 22410 2378 22466 2412
rect 22500 2378 22556 2412
rect 22590 2378 22646 2412
rect 22680 2378 22736 2412
rect 22770 2378 22910 2412
rect 21616 2350 22910 2378
rect 22976 3599 24270 3630
rect 25310 4150 26570 4190
rect 26730 4150 27990 4190
rect 25310 3980 25350 4150
rect 25420 4090 25480 4110
rect 25420 4050 25430 4090
rect 25470 4050 25480 4090
rect 25420 4030 25480 4050
rect 25530 4090 25610 4110
rect 25530 4050 25550 4090
rect 25590 4050 25610 4090
rect 25530 4030 25610 4050
rect 25660 4090 25720 4110
rect 25660 4050 25670 4090
rect 25710 4050 25720 4090
rect 25660 4030 25720 4050
rect 25900 4090 25960 4110
rect 25900 4050 25910 4090
rect 25950 4050 25960 4090
rect 25900 4030 25960 4050
rect 26140 4090 26200 4110
rect 26140 4050 26150 4090
rect 26190 4050 26200 4090
rect 26140 4030 26200 4050
rect 26250 4090 26330 4110
rect 26250 4050 26270 4090
rect 26310 4050 26330 4090
rect 26250 4030 26330 4050
rect 26380 4090 26440 4110
rect 26380 4050 26390 4090
rect 26430 4050 26440 4090
rect 26380 4030 26440 4050
rect 26620 4090 26680 4110
rect 26620 4050 26630 4090
rect 26670 4050 26680 4090
rect 26620 4030 26680 4050
rect 26860 4090 26920 4110
rect 26860 4050 26870 4090
rect 26910 4050 26920 4090
rect 26860 4030 26920 4050
rect 26970 4090 27050 4110
rect 26970 4050 26990 4090
rect 27030 4050 27050 4090
rect 26970 4030 27050 4050
rect 27100 4090 27160 4110
rect 27100 4050 27110 4090
rect 27150 4050 27160 4090
rect 27100 4030 27160 4050
rect 27340 4090 27400 4110
rect 27340 4050 27350 4090
rect 27390 4050 27400 4090
rect 27340 4030 27400 4050
rect 27580 4090 27640 4110
rect 27580 4050 27590 4090
rect 27630 4050 27640 4090
rect 27580 4030 27640 4050
rect 27690 4090 27770 4110
rect 27690 4050 27710 4090
rect 27750 4050 27770 4090
rect 27690 4030 27770 4050
rect 25430 3990 25470 4030
rect 25550 3990 25590 4030
rect 25670 3990 25710 4030
rect 25910 3990 25950 4030
rect 26150 3990 26190 4030
rect 26270 3990 26310 4030
rect 26390 3990 26430 4030
rect 26630 3990 26670 4030
rect 26870 3990 26910 4030
rect 26990 3990 27030 4030
rect 27110 3990 27150 4030
rect 27350 3990 27390 4030
rect 27590 3990 27630 4030
rect 27710 3990 27750 4030
rect 25310 3650 25350 3820
rect 25420 3970 25480 3990
rect 25420 3930 25430 3970
rect 25470 3930 25480 3970
rect 25420 3870 25480 3930
rect 25420 3830 25430 3870
rect 25470 3830 25480 3870
rect 25420 3750 25480 3830
rect 25540 3970 25600 3990
rect 25540 3930 25550 3970
rect 25590 3930 25600 3970
rect 25540 3870 25600 3930
rect 25540 3830 25550 3870
rect 25590 3830 25600 3870
rect 25540 3810 25600 3830
rect 25660 3970 25720 3990
rect 25660 3930 25670 3970
rect 25710 3930 25720 3970
rect 25660 3870 25720 3930
rect 25660 3830 25670 3870
rect 25710 3830 25720 3870
rect 25660 3810 25720 3830
rect 25780 3970 25840 3990
rect 25780 3930 25790 3970
rect 25830 3930 25840 3970
rect 25780 3870 25840 3930
rect 25780 3830 25790 3870
rect 25830 3830 25840 3870
rect 25780 3810 25840 3830
rect 25900 3970 25960 3990
rect 25900 3930 25910 3970
rect 25950 3930 25960 3970
rect 25900 3870 25960 3930
rect 25900 3830 25910 3870
rect 25950 3830 25960 3870
rect 25900 3810 25960 3830
rect 26020 3970 26080 3990
rect 26020 3930 26030 3970
rect 26070 3930 26080 3970
rect 26020 3870 26080 3930
rect 26020 3830 26030 3870
rect 26070 3830 26080 3870
rect 26020 3810 26080 3830
rect 26140 3970 26200 3990
rect 26140 3930 26150 3970
rect 26190 3930 26200 3970
rect 26140 3870 26200 3930
rect 26140 3830 26150 3870
rect 26190 3830 26200 3870
rect 26140 3810 26200 3830
rect 26260 3970 26320 3990
rect 26260 3930 26270 3970
rect 26310 3930 26320 3970
rect 26260 3870 26320 3930
rect 26260 3830 26270 3870
rect 26310 3830 26320 3870
rect 26260 3810 26320 3830
rect 26380 3970 26440 3990
rect 26380 3930 26390 3970
rect 26430 3930 26440 3970
rect 26380 3870 26440 3930
rect 26380 3830 26390 3870
rect 26430 3830 26440 3870
rect 26380 3810 26440 3830
rect 26500 3970 26560 3990
rect 26500 3930 26510 3970
rect 26550 3930 26560 3970
rect 26500 3870 26560 3930
rect 26500 3830 26510 3870
rect 26550 3830 26560 3870
rect 26500 3810 26560 3830
rect 26620 3970 26680 3990
rect 26620 3930 26630 3970
rect 26670 3930 26680 3970
rect 26620 3870 26680 3930
rect 26620 3830 26630 3870
rect 26670 3830 26680 3870
rect 26620 3810 26680 3830
rect 26740 3970 26800 3990
rect 26740 3930 26750 3970
rect 26790 3930 26800 3970
rect 26740 3870 26800 3930
rect 26740 3830 26750 3870
rect 26790 3830 26800 3870
rect 26740 3810 26800 3830
rect 26860 3970 26920 3990
rect 26860 3930 26870 3970
rect 26910 3930 26920 3970
rect 26860 3870 26920 3930
rect 26860 3830 26870 3870
rect 26910 3830 26920 3870
rect 26860 3810 26920 3830
rect 26980 3970 27040 3990
rect 26980 3930 26990 3970
rect 27030 3930 27040 3970
rect 26980 3870 27040 3930
rect 26980 3830 26990 3870
rect 27030 3830 27040 3870
rect 26980 3810 27040 3830
rect 27100 3970 27160 3990
rect 27100 3930 27110 3970
rect 27150 3930 27160 3970
rect 27100 3870 27160 3930
rect 27100 3830 27110 3870
rect 27150 3830 27160 3870
rect 27100 3810 27160 3830
rect 27220 3970 27280 3990
rect 27220 3930 27230 3970
rect 27270 3930 27280 3970
rect 27220 3870 27280 3930
rect 27220 3830 27230 3870
rect 27270 3830 27280 3870
rect 27220 3810 27280 3830
rect 27340 3970 27400 3990
rect 27340 3930 27350 3970
rect 27390 3930 27400 3970
rect 27340 3870 27400 3930
rect 27340 3830 27350 3870
rect 27390 3830 27400 3870
rect 27340 3810 27400 3830
rect 27460 3970 27520 3990
rect 27460 3930 27470 3970
rect 27510 3930 27520 3970
rect 27460 3870 27520 3930
rect 27460 3830 27470 3870
rect 27510 3830 27520 3870
rect 27460 3810 27520 3830
rect 27580 3970 27640 3990
rect 27580 3930 27590 3970
rect 27630 3930 27640 3970
rect 27580 3870 27640 3930
rect 27580 3830 27590 3870
rect 27630 3830 27640 3870
rect 27580 3810 27640 3830
rect 27700 3970 27760 3990
rect 27700 3930 27710 3970
rect 27750 3930 27760 3970
rect 27700 3870 27760 3930
rect 27700 3830 27710 3870
rect 27750 3830 27760 3870
rect 27700 3810 27760 3830
rect 27820 3970 27880 3990
rect 27820 3930 27830 3970
rect 27870 3930 27880 3970
rect 27820 3870 27880 3930
rect 27820 3830 27830 3870
rect 27870 3830 27880 3870
rect 25790 3770 25830 3810
rect 26030 3770 26070 3810
rect 26510 3770 26550 3810
rect 26750 3770 26790 3810
rect 27230 3770 27270 3810
rect 27470 3770 27510 3810
rect 25420 3710 25430 3750
rect 25470 3710 25480 3750
rect 25420 3690 25480 3710
rect 25590 3750 25670 3770
rect 25590 3710 25610 3750
rect 25650 3710 25670 3750
rect 25590 3690 25670 3710
rect 25770 3750 25850 3770
rect 25770 3710 25790 3750
rect 25830 3710 25850 3750
rect 25770 3690 25850 3710
rect 26010 3750 26090 3770
rect 26010 3710 26030 3750
rect 26070 3710 26090 3750
rect 26010 3690 26090 3710
rect 26250 3750 26330 3770
rect 26250 3710 26270 3750
rect 26310 3710 26330 3750
rect 26250 3690 26330 3710
rect 26490 3750 26570 3770
rect 26490 3710 26510 3750
rect 26550 3710 26570 3750
rect 26490 3690 26570 3710
rect 26730 3750 26810 3770
rect 26730 3710 26750 3750
rect 26790 3710 26810 3750
rect 26730 3690 26810 3710
rect 26970 3750 27050 3770
rect 26970 3710 26990 3750
rect 27030 3710 27050 3750
rect 26970 3690 27050 3710
rect 27210 3750 27290 3770
rect 27210 3710 27230 3750
rect 27270 3710 27290 3750
rect 27210 3690 27290 3710
rect 27450 3750 27530 3770
rect 27450 3710 27470 3750
rect 27510 3710 27530 3750
rect 27450 3690 27530 3710
rect 27640 3750 27700 3770
rect 27640 3710 27650 3750
rect 27690 3710 27700 3750
rect 27640 3690 27700 3710
rect 27820 3750 27880 3830
rect 27820 3710 27830 3750
rect 27870 3710 27880 3750
rect 27820 3690 27880 3710
rect 27950 3980 27990 4150
rect 25430 3650 25470 3690
rect 27830 3650 27870 3690
rect 27950 3650 27990 3820
rect 25310 3610 26570 3650
rect 26730 3610 27990 3650
rect 28350 4170 28710 4190
rect 28750 4190 28770 4210
rect 28930 4210 29010 4230
rect 28930 4190 28950 4210
rect 28750 4170 28950 4190
rect 28990 4190 29010 4210
rect 29170 4210 29250 4230
rect 29170 4190 29190 4210
rect 28990 4170 29190 4190
rect 29230 4190 29250 4210
rect 29410 4210 29490 4230
rect 29410 4190 29430 4210
rect 29230 4170 29430 4190
rect 29470 4190 29490 4210
rect 29650 4210 29730 4230
rect 29650 4190 29670 4210
rect 29710 4190 29730 4210
rect 29890 4210 29970 4230
rect 29890 4190 29910 4210
rect 29470 4170 29610 4190
rect 29770 4170 29910 4190
rect 29950 4190 29970 4210
rect 30130 4210 30210 4230
rect 30130 4190 30150 4210
rect 29950 4170 30150 4190
rect 30190 4190 30210 4210
rect 30370 4210 30450 4230
rect 30370 4190 30390 4210
rect 30190 4170 30390 4190
rect 30430 4190 30450 4210
rect 30610 4210 30690 4230
rect 30610 4190 30630 4210
rect 30430 4170 30630 4190
rect 30670 4190 30690 4210
rect 30850 4210 30930 4230
rect 30850 4190 30870 4210
rect 30670 4170 30870 4190
rect 30910 4190 30930 4210
rect 30910 4170 31030 4190
rect 28350 4150 29610 4170
rect 29770 4150 31030 4170
rect 28350 3980 28390 4150
rect 28570 4090 28650 4110
rect 28570 4050 28590 4090
rect 28630 4050 28650 4090
rect 28570 4030 28650 4050
rect 28700 4090 28760 4110
rect 28700 4050 28710 4090
rect 28750 4050 28760 4090
rect 28700 4030 28760 4050
rect 28940 4090 29000 4110
rect 28940 4050 28950 4090
rect 28990 4050 29000 4090
rect 28940 4030 29000 4050
rect 29180 4090 29240 4110
rect 29180 4050 29190 4090
rect 29230 4050 29240 4090
rect 29180 4030 29240 4050
rect 29290 4090 29370 4110
rect 29290 4050 29310 4090
rect 29350 4050 29370 4090
rect 29290 4030 29370 4050
rect 29420 4090 29480 4110
rect 29420 4050 29430 4090
rect 29470 4050 29480 4090
rect 29420 4030 29480 4050
rect 29660 4090 29720 4110
rect 29660 4050 29670 4090
rect 29710 4050 29720 4090
rect 29660 4030 29720 4050
rect 29900 4090 29960 4110
rect 29900 4050 29910 4090
rect 29950 4050 29960 4090
rect 29900 4030 29960 4050
rect 30010 4090 30090 4110
rect 30010 4050 30030 4090
rect 30070 4050 30090 4090
rect 30010 4030 30090 4050
rect 30140 4090 30200 4110
rect 30140 4050 30150 4090
rect 30190 4050 30200 4090
rect 30140 4030 30200 4050
rect 30380 4090 30440 4110
rect 30380 4050 30390 4090
rect 30430 4050 30440 4090
rect 30380 4030 30440 4050
rect 30620 4090 30680 4110
rect 30620 4050 30630 4090
rect 30670 4050 30680 4090
rect 30620 4030 30680 4050
rect 30730 4090 30810 4110
rect 30730 4050 30750 4090
rect 30790 4050 30810 4090
rect 30730 4030 30810 4050
rect 30860 4090 30920 4110
rect 30860 4050 30870 4090
rect 30910 4050 30920 4090
rect 30860 4030 30920 4050
rect 28590 3990 28630 4030
rect 28710 3990 28750 4030
rect 28950 3990 28990 4030
rect 29190 3990 29230 4030
rect 29310 3990 29350 4030
rect 29430 3990 29470 4030
rect 29670 3990 29710 4030
rect 29910 3990 29950 4030
rect 30030 3990 30070 4030
rect 30150 3990 30190 4030
rect 30390 3990 30430 4030
rect 30630 3990 30670 4030
rect 30750 3990 30790 4030
rect 30870 3990 30910 4030
rect 28350 3650 28390 3820
rect 28460 3970 28520 3990
rect 28460 3930 28470 3970
rect 28510 3930 28520 3970
rect 28460 3870 28520 3930
rect 28460 3830 28470 3870
rect 28510 3830 28520 3870
rect 28460 3810 28520 3830
rect 28580 3970 28640 3990
rect 28580 3930 28590 3970
rect 28630 3930 28640 3970
rect 28580 3870 28640 3930
rect 28580 3830 28590 3870
rect 28630 3830 28640 3870
rect 28580 3810 28640 3830
rect 28700 3970 28760 3990
rect 28700 3930 28710 3970
rect 28750 3930 28760 3970
rect 28700 3870 28760 3930
rect 28700 3830 28710 3870
rect 28750 3830 28760 3870
rect 28700 3810 28760 3830
rect 28820 3970 28880 3990
rect 28820 3930 28830 3970
rect 28870 3930 28880 3970
rect 28820 3870 28880 3930
rect 28820 3830 28830 3870
rect 28870 3830 28880 3870
rect 28820 3810 28880 3830
rect 28940 3970 29000 3990
rect 28940 3930 28950 3970
rect 28990 3930 29000 3970
rect 28940 3870 29000 3930
rect 28940 3830 28950 3870
rect 28990 3830 29000 3870
rect 28940 3810 29000 3830
rect 29060 3970 29120 3990
rect 29060 3930 29070 3970
rect 29110 3930 29120 3970
rect 29060 3870 29120 3930
rect 29060 3830 29070 3870
rect 29110 3830 29120 3870
rect 29060 3810 29120 3830
rect 29180 3970 29240 3990
rect 29180 3930 29190 3970
rect 29230 3930 29240 3970
rect 29180 3870 29240 3930
rect 29180 3830 29190 3870
rect 29230 3830 29240 3870
rect 29180 3810 29240 3830
rect 29300 3970 29360 3990
rect 29300 3930 29310 3970
rect 29350 3930 29360 3970
rect 29300 3870 29360 3930
rect 29300 3830 29310 3870
rect 29350 3830 29360 3870
rect 29300 3810 29360 3830
rect 29420 3970 29480 3990
rect 29420 3930 29430 3970
rect 29470 3930 29480 3970
rect 29420 3870 29480 3930
rect 29420 3830 29430 3870
rect 29470 3830 29480 3870
rect 29420 3810 29480 3830
rect 29540 3970 29600 3990
rect 29540 3930 29550 3970
rect 29590 3930 29600 3970
rect 29540 3870 29600 3930
rect 29540 3830 29550 3870
rect 29590 3830 29600 3870
rect 29540 3810 29600 3830
rect 29660 3970 29720 3990
rect 29660 3930 29670 3970
rect 29710 3930 29720 3970
rect 29660 3870 29720 3930
rect 29660 3830 29670 3870
rect 29710 3830 29720 3870
rect 29660 3810 29720 3830
rect 29780 3970 29840 3990
rect 29780 3930 29790 3970
rect 29830 3930 29840 3970
rect 29780 3870 29840 3930
rect 29780 3830 29790 3870
rect 29830 3830 29840 3870
rect 29780 3810 29840 3830
rect 29900 3970 29960 3990
rect 29900 3930 29910 3970
rect 29950 3930 29960 3970
rect 29900 3870 29960 3930
rect 29900 3830 29910 3870
rect 29950 3830 29960 3870
rect 29900 3810 29960 3830
rect 30020 3970 30080 3990
rect 30020 3930 30030 3970
rect 30070 3930 30080 3970
rect 30020 3870 30080 3930
rect 30020 3830 30030 3870
rect 30070 3830 30080 3870
rect 30020 3810 30080 3830
rect 30140 3970 30200 3990
rect 30140 3930 30150 3970
rect 30190 3930 30200 3970
rect 30140 3870 30200 3930
rect 30140 3830 30150 3870
rect 30190 3830 30200 3870
rect 30140 3810 30200 3830
rect 30260 3970 30320 3990
rect 30260 3930 30270 3970
rect 30310 3930 30320 3970
rect 30260 3870 30320 3930
rect 30260 3830 30270 3870
rect 30310 3830 30320 3870
rect 30260 3810 30320 3830
rect 30380 3970 30440 3990
rect 30380 3930 30390 3970
rect 30430 3930 30440 3970
rect 30380 3870 30440 3930
rect 30380 3830 30390 3870
rect 30430 3830 30440 3870
rect 30380 3810 30440 3830
rect 30500 3970 30560 3990
rect 30500 3930 30510 3970
rect 30550 3930 30560 3970
rect 30500 3870 30560 3930
rect 30500 3830 30510 3870
rect 30550 3830 30560 3870
rect 30500 3810 30560 3830
rect 30620 3970 30680 3990
rect 30620 3930 30630 3970
rect 30670 3930 30680 3970
rect 30620 3870 30680 3930
rect 30620 3830 30630 3870
rect 30670 3830 30680 3870
rect 30620 3810 30680 3830
rect 30740 3970 30800 3990
rect 30740 3930 30750 3970
rect 30790 3930 30800 3970
rect 30740 3870 30800 3930
rect 30740 3830 30750 3870
rect 30790 3830 30800 3870
rect 30740 3810 30800 3830
rect 30860 3970 30920 3990
rect 30860 3930 30870 3970
rect 30910 3930 30920 3970
rect 30860 3870 30920 3930
rect 30860 3830 30870 3870
rect 30910 3830 30920 3870
rect 28830 3770 28870 3810
rect 29070 3770 29110 3810
rect 29550 3770 29590 3810
rect 29790 3770 29830 3810
rect 30270 3770 30310 3810
rect 30510 3770 30550 3810
rect 28640 3750 28700 3770
rect 28640 3710 28650 3750
rect 28690 3710 28700 3750
rect 28640 3690 28700 3710
rect 28810 3750 28890 3770
rect 28810 3710 28830 3750
rect 28870 3710 28890 3750
rect 28810 3690 28890 3710
rect 29050 3750 29130 3770
rect 29050 3710 29070 3750
rect 29110 3710 29130 3750
rect 29050 3690 29130 3710
rect 29290 3750 29370 3770
rect 29290 3710 29310 3750
rect 29350 3710 29370 3750
rect 29290 3690 29370 3710
rect 29530 3750 29610 3770
rect 29530 3710 29550 3750
rect 29590 3710 29610 3750
rect 29530 3690 29610 3710
rect 29770 3750 29850 3770
rect 29770 3710 29790 3750
rect 29830 3710 29850 3750
rect 29770 3690 29850 3710
rect 30010 3750 30090 3770
rect 30010 3710 30030 3750
rect 30070 3710 30090 3750
rect 30010 3690 30090 3710
rect 30250 3750 30330 3770
rect 30250 3710 30270 3750
rect 30310 3710 30330 3750
rect 30250 3690 30330 3710
rect 30490 3750 30570 3770
rect 30490 3710 30510 3750
rect 30550 3710 30570 3750
rect 30490 3690 30570 3710
rect 30670 3750 30750 3770
rect 30670 3710 30690 3750
rect 30730 3710 30750 3750
rect 30670 3690 30750 3710
rect 30860 3750 30920 3830
rect 30860 3710 30870 3750
rect 30910 3710 30920 3750
rect 30860 3690 30920 3710
rect 30990 3980 31030 4150
rect 30870 3650 30910 3690
rect 30990 3650 31030 3820
rect 28350 3610 29610 3650
rect 29770 3610 31030 3650
rect 22976 3576 23106 3599
rect 22976 3542 23010 3576
rect 23044 3565 23106 3576
rect 23140 3565 23196 3599
rect 23230 3565 23286 3599
rect 23320 3565 23376 3599
rect 23410 3565 23466 3599
rect 23500 3565 23556 3599
rect 23590 3565 23646 3599
rect 23680 3565 23736 3599
rect 23770 3565 23826 3599
rect 23860 3565 23916 3599
rect 23950 3565 24006 3599
rect 24040 3565 24096 3599
rect 24130 3576 24270 3599
rect 24130 3565 24197 3576
rect 23044 3542 24197 3565
rect 24231 3542 24270 3576
rect 22976 3535 24270 3542
rect 22976 3486 23075 3535
rect 22976 3452 23010 3486
rect 23044 3452 23075 3486
rect 24020 3486 24270 3535
rect 24020 3471 24197 3486
rect 22976 3396 23075 3452
rect 22976 3362 23010 3396
rect 23044 3362 23075 3396
rect 22976 3306 23075 3362
rect 22976 3272 23010 3306
rect 23044 3272 23075 3306
rect 22976 3216 23075 3272
rect 22976 3182 23010 3216
rect 23044 3182 23075 3216
rect 22976 3126 23075 3182
rect 22976 3092 23010 3126
rect 23044 3092 23075 3126
rect 22976 3036 23075 3092
rect 22976 3002 23010 3036
rect 23044 3002 23075 3036
rect 22976 2946 23075 3002
rect 22976 2912 23010 2946
rect 23044 2912 23075 2946
rect 22976 2856 23075 2912
rect 22976 2822 23010 2856
rect 23044 2822 23075 2856
rect 22976 2766 23075 2822
rect 22976 2732 23010 2766
rect 23044 2732 23075 2766
rect 22976 2676 23075 2732
rect 22976 2642 23010 2676
rect 23044 2642 23075 2676
rect 22976 2586 23075 2642
rect 22976 2552 23010 2586
rect 23044 2552 23075 2586
rect 22976 2496 23075 2552
rect 23139 3452 24197 3471
rect 24231 3452 24270 3486
rect 23139 3418 23270 3452
rect 23304 3418 23360 3452
rect 23394 3418 23450 3452
rect 23484 3418 23540 3452
rect 23574 3418 23630 3452
rect 23664 3418 23720 3452
rect 23754 3418 23810 3452
rect 23844 3418 23900 3452
rect 23934 3418 23990 3452
rect 24024 3418 24270 3452
rect 23139 3399 24270 3418
rect 23139 3395 23211 3399
rect 23139 3361 23158 3395
rect 23192 3361 23211 3395
rect 23139 3305 23211 3361
rect 24020 3396 24270 3399
rect 24020 3376 24197 3396
rect 24020 3342 24048 3376
rect 24082 3362 24197 3376
rect 24231 3362 24270 3396
rect 24082 3342 24270 3362
rect 23139 3271 23158 3305
rect 23192 3271 23211 3305
rect 23139 3215 23211 3271
rect 23139 3181 23158 3215
rect 23192 3181 23211 3215
rect 23139 3125 23211 3181
rect 23139 3091 23158 3125
rect 23192 3091 23211 3125
rect 23139 3035 23211 3091
rect 23139 3001 23158 3035
rect 23192 3001 23211 3035
rect 23139 2945 23211 3001
rect 23139 2911 23158 2945
rect 23192 2911 23211 2945
rect 23139 2855 23211 2911
rect 23139 2821 23158 2855
rect 23192 2821 23211 2855
rect 23139 2765 23211 2821
rect 23139 2731 23158 2765
rect 23192 2731 23211 2765
rect 23139 2675 23211 2731
rect 23139 2641 23158 2675
rect 23192 2641 23211 2675
rect 23273 3278 23967 3337
rect 23273 3244 23334 3278
rect 23368 3250 23424 3278
rect 23458 3250 23514 3278
rect 23548 3250 23604 3278
rect 23380 3244 23424 3250
rect 23480 3244 23514 3250
rect 23580 3244 23604 3250
rect 23638 3250 23694 3278
rect 23638 3244 23646 3250
rect 23273 3216 23346 3244
rect 23380 3216 23446 3244
rect 23480 3216 23546 3244
rect 23580 3216 23646 3244
rect 23680 3244 23694 3250
rect 23728 3250 23784 3278
rect 23728 3244 23746 3250
rect 23680 3216 23746 3244
rect 23780 3244 23784 3250
rect 23818 3250 23874 3278
rect 23818 3244 23846 3250
rect 23908 3244 23967 3278
rect 23780 3216 23846 3244
rect 23880 3216 23967 3244
rect 23273 3188 23967 3216
rect 23273 3154 23334 3188
rect 23368 3154 23424 3188
rect 23458 3154 23514 3188
rect 23548 3154 23604 3188
rect 23638 3154 23694 3188
rect 23728 3154 23784 3188
rect 23818 3154 23874 3188
rect 23908 3154 23967 3188
rect 23273 3150 23967 3154
rect 23273 3116 23346 3150
rect 23380 3116 23446 3150
rect 23480 3116 23546 3150
rect 23580 3116 23646 3150
rect 23680 3116 23746 3150
rect 23780 3116 23846 3150
rect 23880 3116 23967 3150
rect 23273 3098 23967 3116
rect 23273 3064 23334 3098
rect 23368 3064 23424 3098
rect 23458 3064 23514 3098
rect 23548 3064 23604 3098
rect 23638 3064 23694 3098
rect 23728 3064 23784 3098
rect 23818 3064 23874 3098
rect 23908 3064 23967 3098
rect 23273 3050 23967 3064
rect 23273 3016 23346 3050
rect 23380 3016 23446 3050
rect 23480 3016 23546 3050
rect 23580 3016 23646 3050
rect 23680 3016 23746 3050
rect 23780 3016 23846 3050
rect 23880 3016 23967 3050
rect 23273 3008 23967 3016
rect 23273 2974 23334 3008
rect 23368 2974 23424 3008
rect 23458 2974 23514 3008
rect 23548 2974 23604 3008
rect 23638 2974 23694 3008
rect 23728 2974 23784 3008
rect 23818 2974 23874 3008
rect 23908 2974 23967 3008
rect 23273 2950 23967 2974
rect 23273 2918 23346 2950
rect 23380 2918 23446 2950
rect 23480 2918 23546 2950
rect 23580 2918 23646 2950
rect 23273 2884 23334 2918
rect 23380 2916 23424 2918
rect 23480 2916 23514 2918
rect 23580 2916 23604 2918
rect 23368 2884 23424 2916
rect 23458 2884 23514 2916
rect 23548 2884 23604 2916
rect 23638 2916 23646 2918
rect 23680 2918 23746 2950
rect 23680 2916 23694 2918
rect 23638 2884 23694 2916
rect 23728 2916 23746 2918
rect 23780 2918 23846 2950
rect 23880 2918 23967 2950
rect 23780 2916 23784 2918
rect 23728 2884 23784 2916
rect 23818 2916 23846 2918
rect 23818 2884 23874 2916
rect 23908 2884 23967 2918
rect 23273 2850 23967 2884
rect 23273 2828 23346 2850
rect 23380 2828 23446 2850
rect 23480 2828 23546 2850
rect 23580 2828 23646 2850
rect 23273 2794 23334 2828
rect 23380 2816 23424 2828
rect 23480 2816 23514 2828
rect 23580 2816 23604 2828
rect 23368 2794 23424 2816
rect 23458 2794 23514 2816
rect 23548 2794 23604 2816
rect 23638 2816 23646 2828
rect 23680 2828 23746 2850
rect 23680 2816 23694 2828
rect 23638 2794 23694 2816
rect 23728 2816 23746 2828
rect 23780 2828 23846 2850
rect 23880 2828 23967 2850
rect 23780 2816 23784 2828
rect 23728 2794 23784 2816
rect 23818 2816 23846 2828
rect 23818 2794 23874 2816
rect 23908 2794 23967 2828
rect 23273 2750 23967 2794
rect 23273 2738 23346 2750
rect 23380 2738 23446 2750
rect 23480 2738 23546 2750
rect 23580 2738 23646 2750
rect 23273 2704 23334 2738
rect 23380 2716 23424 2738
rect 23480 2716 23514 2738
rect 23580 2716 23604 2738
rect 23368 2704 23424 2716
rect 23458 2704 23514 2716
rect 23548 2704 23604 2716
rect 23638 2716 23646 2738
rect 23680 2738 23746 2750
rect 23680 2716 23694 2738
rect 23638 2704 23694 2716
rect 23728 2716 23746 2738
rect 23780 2738 23846 2750
rect 23880 2738 23967 2750
rect 23780 2716 23784 2738
rect 23728 2704 23784 2716
rect 23818 2716 23846 2738
rect 23818 2704 23874 2716
rect 23908 2704 23967 2738
rect 23273 2643 23967 2704
rect 24020 3306 24270 3342
rect 24020 3286 24197 3306
rect 24020 3252 24048 3286
rect 24082 3272 24197 3286
rect 24231 3272 24270 3306
rect 24082 3252 24270 3272
rect 24020 3216 24270 3252
rect 24020 3196 24197 3216
rect 24020 3162 24048 3196
rect 24082 3182 24197 3196
rect 24231 3182 24270 3216
rect 24082 3162 24270 3182
rect 24020 3126 24270 3162
rect 24020 3106 24197 3126
rect 24020 3072 24048 3106
rect 24082 3092 24197 3106
rect 24231 3092 24270 3126
rect 24082 3072 24270 3092
rect 24020 3036 24270 3072
rect 24020 3016 24197 3036
rect 24020 2982 24048 3016
rect 24082 3002 24197 3016
rect 24231 3002 24270 3036
rect 24082 2982 24270 3002
rect 24020 2946 24270 2982
rect 26170 3490 26830 3530
rect 26990 3490 27650 3530
rect 26170 3280 26210 3490
rect 26390 3430 26470 3450
rect 26390 3390 26410 3430
rect 26450 3390 26470 3430
rect 26390 3370 26470 3390
rect 26270 3340 26350 3360
rect 26270 3300 26290 3340
rect 26330 3300 26350 3340
rect 26270 3280 26350 3300
rect 26520 3340 26580 3360
rect 26520 3300 26530 3340
rect 26570 3300 26580 3340
rect 26520 3280 26580 3300
rect 26750 3340 26830 3360
rect 26750 3300 26770 3340
rect 26810 3300 26830 3340
rect 26750 3280 26830 3300
rect 27000 3340 27060 3360
rect 27000 3300 27010 3340
rect 27050 3300 27060 3340
rect 27000 3280 27060 3300
rect 27230 3340 27310 3360
rect 27230 3300 27250 3340
rect 27290 3300 27310 3340
rect 27230 3280 27310 3300
rect 27480 3340 27540 3360
rect 27480 3300 27490 3340
rect 27530 3300 27540 3340
rect 27480 3280 27540 3300
rect 27610 3280 27650 3490
rect 26290 3240 26330 3280
rect 26530 3240 26570 3280
rect 26770 3240 26810 3280
rect 27010 3240 27050 3280
rect 27250 3240 27290 3280
rect 27490 3240 27530 3280
rect 26280 3220 26340 3240
rect 26280 3180 26290 3220
rect 26330 3180 26340 3220
rect 26280 3160 26340 3180
rect 26400 3220 26460 3240
rect 26400 3180 26410 3220
rect 26450 3180 26460 3220
rect 26400 3160 26460 3180
rect 26520 3220 26580 3240
rect 26520 3180 26530 3220
rect 26570 3180 26580 3220
rect 26520 3160 26580 3180
rect 26640 3220 26700 3240
rect 26640 3180 26650 3220
rect 26690 3180 26700 3220
rect 26640 3160 26700 3180
rect 26760 3220 26820 3240
rect 26760 3180 26770 3220
rect 26810 3180 26820 3220
rect 26760 3160 26820 3180
rect 26880 3220 26940 3240
rect 26880 3180 26890 3220
rect 26930 3180 26940 3220
rect 26880 3160 26940 3180
rect 27000 3220 27060 3240
rect 27000 3180 27010 3220
rect 27050 3180 27060 3220
rect 27000 3160 27060 3180
rect 27120 3220 27180 3240
rect 27120 3180 27130 3220
rect 27170 3180 27180 3220
rect 27120 3160 27180 3180
rect 27240 3220 27300 3240
rect 27240 3180 27250 3220
rect 27290 3180 27300 3220
rect 27240 3160 27300 3180
rect 27360 3220 27420 3240
rect 27360 3180 27370 3220
rect 27410 3180 27420 3220
rect 27360 3160 27420 3180
rect 27480 3220 27540 3240
rect 27480 3180 27490 3220
rect 27530 3180 27540 3220
rect 27480 3160 27540 3180
rect 26410 3120 26450 3160
rect 26650 3120 26690 3160
rect 26890 3120 26930 3160
rect 27130 3120 27170 3160
rect 27370 3120 27410 3160
rect 26170 3000 26210 3120
rect 26270 3100 26350 3120
rect 26270 3060 26290 3100
rect 26330 3060 26350 3100
rect 26270 3040 26350 3060
rect 26400 3100 26460 3120
rect 26400 3060 26410 3100
rect 26450 3060 26460 3100
rect 26400 3040 26460 3060
rect 26640 3100 26700 3120
rect 26640 3060 26650 3100
rect 26690 3060 26700 3100
rect 26640 3040 26700 3060
rect 26880 3100 26940 3120
rect 26880 3060 26890 3100
rect 26930 3060 26940 3100
rect 26880 3040 26940 3060
rect 27120 3100 27180 3120
rect 27120 3060 27130 3100
rect 27170 3060 27180 3100
rect 27120 3040 27180 3060
rect 27360 3100 27420 3120
rect 27360 3060 27370 3100
rect 27410 3060 27420 3100
rect 27360 3040 27420 3060
rect 27610 3000 27650 3120
rect 26170 2960 26830 3000
rect 26990 2980 27650 3000
rect 26990 2960 27370 2980
rect 24020 2926 24197 2946
rect 24020 2892 24048 2926
rect 24082 2912 24197 2926
rect 24231 2912 24270 2946
rect 26390 2920 26470 2960
rect 26630 2920 26710 2960
rect 26870 2920 26950 2960
rect 27110 2920 27190 2960
rect 27350 2940 27370 2960
rect 27410 2960 27650 2980
rect 28690 3490 29350 3530
rect 29510 3490 30170 3530
rect 28690 3280 28730 3490
rect 29870 3430 29950 3450
rect 29870 3390 29890 3430
rect 29930 3390 29950 3430
rect 29870 3370 29950 3390
rect 28800 3340 28860 3360
rect 28800 3300 28810 3340
rect 28850 3300 28860 3340
rect 28800 3280 28860 3300
rect 29030 3340 29110 3360
rect 29030 3300 29050 3340
rect 29090 3300 29110 3340
rect 29030 3280 29110 3300
rect 29280 3340 29340 3360
rect 29280 3300 29290 3340
rect 29330 3300 29340 3340
rect 29280 3280 29340 3300
rect 29510 3340 29590 3360
rect 29510 3300 29530 3340
rect 29570 3300 29590 3340
rect 29510 3280 29590 3300
rect 29760 3340 29820 3360
rect 29760 3300 29770 3340
rect 29810 3300 29820 3340
rect 29760 3280 29820 3300
rect 29990 3340 30070 3360
rect 29990 3300 30010 3340
rect 30050 3300 30070 3340
rect 29990 3280 30070 3300
rect 30130 3280 30170 3490
rect 28810 3240 28850 3280
rect 29050 3240 29090 3280
rect 29290 3240 29330 3280
rect 29530 3240 29570 3280
rect 29770 3240 29810 3280
rect 30010 3240 30050 3280
rect 28800 3220 28860 3240
rect 28800 3180 28810 3220
rect 28850 3180 28860 3220
rect 28800 3160 28860 3180
rect 28920 3220 28980 3240
rect 28920 3180 28930 3220
rect 28970 3180 28980 3220
rect 28920 3160 28980 3180
rect 29040 3220 29100 3240
rect 29040 3180 29050 3220
rect 29090 3180 29100 3220
rect 29040 3160 29100 3180
rect 29160 3220 29220 3240
rect 29160 3180 29170 3220
rect 29210 3180 29220 3220
rect 29160 3160 29220 3180
rect 29280 3220 29340 3240
rect 29280 3180 29290 3220
rect 29330 3180 29340 3220
rect 29280 3160 29340 3180
rect 29400 3220 29460 3240
rect 29400 3180 29410 3220
rect 29450 3180 29460 3220
rect 29400 3160 29460 3180
rect 29520 3220 29580 3240
rect 29520 3180 29530 3220
rect 29570 3180 29580 3220
rect 29520 3160 29580 3180
rect 29640 3220 29700 3240
rect 29640 3180 29650 3220
rect 29690 3180 29700 3220
rect 29640 3160 29700 3180
rect 29760 3220 29820 3240
rect 29760 3180 29770 3220
rect 29810 3180 29820 3220
rect 29760 3160 29820 3180
rect 29880 3220 29940 3240
rect 29880 3180 29890 3220
rect 29930 3180 29940 3220
rect 29880 3160 29940 3180
rect 30000 3220 30060 3240
rect 30000 3180 30010 3220
rect 30050 3180 30060 3220
rect 30000 3160 30060 3180
rect 28930 3120 28970 3160
rect 29170 3120 29210 3160
rect 29410 3120 29450 3160
rect 29650 3120 29690 3160
rect 29890 3120 29930 3160
rect 28690 3000 28730 3120
rect 28920 3100 28980 3120
rect 28920 3060 28930 3100
rect 28970 3060 28980 3100
rect 28920 3040 28980 3060
rect 29160 3100 29220 3120
rect 29160 3060 29170 3100
rect 29210 3060 29220 3100
rect 29160 3040 29220 3060
rect 29400 3100 29460 3120
rect 29400 3060 29410 3100
rect 29450 3060 29460 3100
rect 29400 3040 29460 3060
rect 29640 3100 29700 3120
rect 29640 3060 29650 3100
rect 29690 3060 29700 3100
rect 29640 3040 29700 3060
rect 29880 3100 29940 3120
rect 29880 3060 29890 3100
rect 29930 3060 29940 3100
rect 29880 3040 29940 3060
rect 29990 3100 30070 3120
rect 29990 3060 30010 3100
rect 30050 3060 30070 3100
rect 29990 3040 30070 3060
rect 30130 3000 30170 3120
rect 28690 2960 30170 3000
rect 27410 2940 27430 2960
rect 27350 2920 27430 2940
rect 29870 2920 29950 2960
rect 24082 2892 24270 2912
rect 24020 2856 24270 2892
rect 24020 2836 24197 2856
rect 24020 2802 24048 2836
rect 24082 2822 24197 2836
rect 24231 2822 24270 2856
rect 24082 2802 24270 2822
rect 24020 2766 24270 2802
rect 24020 2746 24197 2766
rect 24020 2712 24048 2746
rect 24082 2732 24197 2746
rect 24231 2732 24270 2766
rect 24082 2712 24270 2732
rect 24020 2676 24270 2712
rect 24020 2656 24197 2676
rect 23139 2581 23211 2641
rect 24020 2622 24048 2656
rect 24082 2642 24197 2656
rect 24231 2642 24270 2676
rect 24082 2622 24270 2642
rect 24020 2586 24270 2622
rect 24020 2581 24197 2586
rect 23139 2562 24197 2581
rect 23139 2528 23236 2562
rect 23270 2528 23326 2562
rect 23360 2528 23416 2562
rect 23450 2528 23506 2562
rect 23540 2528 23596 2562
rect 23630 2528 23686 2562
rect 23720 2528 23776 2562
rect 23810 2528 23866 2562
rect 23900 2528 23956 2562
rect 23990 2552 24197 2562
rect 24231 2552 24270 2586
rect 23990 2528 24270 2552
rect 23139 2509 24270 2528
rect 22976 2462 23010 2496
rect 23044 2462 23075 2496
rect 22976 2445 23075 2462
rect 24020 2496 24270 2509
rect 24020 2462 24197 2496
rect 24231 2462 24270 2496
rect 24020 2445 24270 2462
rect 22976 2412 24270 2445
rect 22976 2378 23106 2412
rect 23140 2378 23196 2412
rect 23230 2378 23286 2412
rect 23320 2378 23376 2412
rect 23410 2378 23466 2412
rect 23500 2378 23556 2412
rect 23590 2378 23646 2412
rect 23680 2378 23736 2412
rect 23770 2378 23826 2412
rect 23860 2378 23916 2412
rect 23950 2378 24006 2412
rect 24040 2378 24096 2412
rect 24130 2378 24270 2412
rect 22976 2350 24270 2378
rect 20250 2270 24270 2350
rect 20256 2239 21550 2270
rect 20256 2216 20386 2239
rect 20256 2182 20290 2216
rect 20324 2205 20386 2216
rect 20420 2205 20476 2239
rect 20510 2205 20566 2239
rect 20600 2205 20656 2239
rect 20690 2205 20746 2239
rect 20780 2205 20836 2239
rect 20870 2205 20926 2239
rect 20960 2205 21016 2239
rect 21050 2205 21106 2239
rect 21140 2205 21196 2239
rect 21230 2205 21286 2239
rect 21320 2205 21376 2239
rect 21410 2216 21550 2239
rect 21410 2205 21477 2216
rect 20324 2182 21477 2205
rect 21511 2182 21550 2216
rect 20256 2175 21550 2182
rect 20256 2126 20355 2175
rect 20256 2092 20290 2126
rect 20324 2092 20355 2126
rect 21300 2126 21550 2175
rect 21300 2111 21477 2126
rect 20256 2036 20355 2092
rect 20256 2002 20290 2036
rect 20324 2002 20355 2036
rect 20256 1946 20355 2002
rect 20256 1912 20290 1946
rect 20324 1912 20355 1946
rect 20256 1856 20355 1912
rect 20256 1822 20290 1856
rect 20324 1822 20355 1856
rect 20256 1766 20355 1822
rect 20256 1732 20290 1766
rect 20324 1732 20355 1766
rect 20256 1676 20355 1732
rect 20256 1642 20290 1676
rect 20324 1642 20355 1676
rect 20256 1586 20355 1642
rect 20256 1552 20290 1586
rect 20324 1552 20355 1586
rect 20256 1496 20355 1552
rect 20256 1462 20290 1496
rect 20324 1462 20355 1496
rect 20256 1406 20355 1462
rect 20256 1372 20290 1406
rect 20324 1372 20355 1406
rect 20256 1316 20355 1372
rect 20256 1282 20290 1316
rect 20324 1282 20355 1316
rect 20256 1226 20355 1282
rect 20256 1192 20290 1226
rect 20324 1192 20355 1226
rect 20256 1136 20355 1192
rect 20419 2092 21477 2111
rect 21511 2092 21550 2126
rect 20419 2058 20550 2092
rect 20584 2058 20640 2092
rect 20674 2058 20730 2092
rect 20764 2058 20820 2092
rect 20854 2058 20910 2092
rect 20944 2058 21000 2092
rect 21034 2058 21090 2092
rect 21124 2058 21180 2092
rect 21214 2058 21270 2092
rect 21304 2058 21550 2092
rect 20419 2039 21550 2058
rect 20419 2035 20491 2039
rect 20419 2001 20438 2035
rect 20472 2001 20491 2035
rect 20419 1945 20491 2001
rect 21300 2036 21550 2039
rect 21300 2016 21477 2036
rect 21300 1982 21328 2016
rect 21362 2002 21477 2016
rect 21511 2002 21550 2036
rect 21362 1982 21550 2002
rect 20419 1911 20438 1945
rect 20472 1911 20491 1945
rect 20419 1855 20491 1911
rect 20419 1821 20438 1855
rect 20472 1821 20491 1855
rect 20419 1765 20491 1821
rect 20419 1731 20438 1765
rect 20472 1731 20491 1765
rect 20419 1675 20491 1731
rect 20419 1641 20438 1675
rect 20472 1641 20491 1675
rect 20419 1585 20491 1641
rect 20419 1551 20438 1585
rect 20472 1551 20491 1585
rect 20419 1495 20491 1551
rect 20419 1461 20438 1495
rect 20472 1461 20491 1495
rect 20419 1405 20491 1461
rect 20419 1371 20438 1405
rect 20472 1371 20491 1405
rect 20419 1315 20491 1371
rect 20419 1281 20438 1315
rect 20472 1281 20491 1315
rect 20553 1918 21247 1977
rect 20553 1884 20614 1918
rect 20648 1890 20704 1918
rect 20738 1890 20794 1918
rect 20828 1890 20884 1918
rect 20660 1884 20704 1890
rect 20760 1884 20794 1890
rect 20860 1884 20884 1890
rect 20918 1890 20974 1918
rect 20918 1884 20926 1890
rect 20553 1856 20626 1884
rect 20660 1856 20726 1884
rect 20760 1856 20826 1884
rect 20860 1856 20926 1884
rect 20960 1884 20974 1890
rect 21008 1890 21064 1918
rect 21008 1884 21026 1890
rect 20960 1856 21026 1884
rect 21060 1884 21064 1890
rect 21098 1890 21154 1918
rect 21098 1884 21126 1890
rect 21188 1884 21247 1918
rect 21060 1856 21126 1884
rect 21160 1856 21247 1884
rect 20553 1828 21247 1856
rect 20553 1794 20614 1828
rect 20648 1794 20704 1828
rect 20738 1794 20794 1828
rect 20828 1794 20884 1828
rect 20918 1794 20974 1828
rect 21008 1794 21064 1828
rect 21098 1794 21154 1828
rect 21188 1794 21247 1828
rect 20553 1790 21247 1794
rect 20553 1756 20626 1790
rect 20660 1756 20726 1790
rect 20760 1756 20826 1790
rect 20860 1756 20926 1790
rect 20960 1756 21026 1790
rect 21060 1756 21126 1790
rect 21160 1756 21247 1790
rect 20553 1738 21247 1756
rect 20553 1704 20614 1738
rect 20648 1704 20704 1738
rect 20738 1704 20794 1738
rect 20828 1704 20884 1738
rect 20918 1704 20974 1738
rect 21008 1704 21064 1738
rect 21098 1704 21154 1738
rect 21188 1704 21247 1738
rect 20553 1690 21247 1704
rect 20553 1656 20626 1690
rect 20660 1656 20726 1690
rect 20760 1656 20826 1690
rect 20860 1656 20926 1690
rect 20960 1656 21026 1690
rect 21060 1656 21126 1690
rect 21160 1656 21247 1690
rect 20553 1648 21247 1656
rect 20553 1614 20614 1648
rect 20648 1614 20704 1648
rect 20738 1614 20794 1648
rect 20828 1614 20884 1648
rect 20918 1614 20974 1648
rect 21008 1614 21064 1648
rect 21098 1614 21154 1648
rect 21188 1614 21247 1648
rect 20553 1590 21247 1614
rect 20553 1558 20626 1590
rect 20660 1558 20726 1590
rect 20760 1558 20826 1590
rect 20860 1558 20926 1590
rect 20553 1524 20614 1558
rect 20660 1556 20704 1558
rect 20760 1556 20794 1558
rect 20860 1556 20884 1558
rect 20648 1524 20704 1556
rect 20738 1524 20794 1556
rect 20828 1524 20884 1556
rect 20918 1556 20926 1558
rect 20960 1558 21026 1590
rect 20960 1556 20974 1558
rect 20918 1524 20974 1556
rect 21008 1556 21026 1558
rect 21060 1558 21126 1590
rect 21160 1558 21247 1590
rect 21060 1556 21064 1558
rect 21008 1524 21064 1556
rect 21098 1556 21126 1558
rect 21098 1524 21154 1556
rect 21188 1524 21247 1558
rect 20553 1490 21247 1524
rect 20553 1468 20626 1490
rect 20660 1468 20726 1490
rect 20760 1468 20826 1490
rect 20860 1468 20926 1490
rect 20553 1434 20614 1468
rect 20660 1456 20704 1468
rect 20760 1456 20794 1468
rect 20860 1456 20884 1468
rect 20648 1434 20704 1456
rect 20738 1434 20794 1456
rect 20828 1434 20884 1456
rect 20918 1456 20926 1468
rect 20960 1468 21026 1490
rect 20960 1456 20974 1468
rect 20918 1434 20974 1456
rect 21008 1456 21026 1468
rect 21060 1468 21126 1490
rect 21160 1468 21247 1490
rect 21060 1456 21064 1468
rect 21008 1434 21064 1456
rect 21098 1456 21126 1468
rect 21098 1434 21154 1456
rect 21188 1434 21247 1468
rect 20553 1390 21247 1434
rect 20553 1378 20626 1390
rect 20660 1378 20726 1390
rect 20760 1378 20826 1390
rect 20860 1378 20926 1390
rect 20553 1344 20614 1378
rect 20660 1356 20704 1378
rect 20760 1356 20794 1378
rect 20860 1356 20884 1378
rect 20648 1344 20704 1356
rect 20738 1344 20794 1356
rect 20828 1344 20884 1356
rect 20918 1356 20926 1378
rect 20960 1378 21026 1390
rect 20960 1356 20974 1378
rect 20918 1344 20974 1356
rect 21008 1356 21026 1378
rect 21060 1378 21126 1390
rect 21160 1378 21247 1390
rect 21060 1356 21064 1378
rect 21008 1344 21064 1356
rect 21098 1356 21126 1378
rect 21098 1344 21154 1356
rect 21188 1344 21247 1378
rect 20553 1283 21247 1344
rect 21300 1946 21550 1982
rect 21300 1926 21477 1946
rect 21300 1892 21328 1926
rect 21362 1912 21477 1926
rect 21511 1912 21550 1946
rect 21362 1892 21550 1912
rect 21300 1856 21550 1892
rect 21300 1836 21477 1856
rect 21300 1802 21328 1836
rect 21362 1822 21477 1836
rect 21511 1822 21550 1856
rect 21362 1802 21550 1822
rect 21300 1766 21550 1802
rect 21300 1746 21477 1766
rect 21300 1712 21328 1746
rect 21362 1732 21477 1746
rect 21511 1732 21550 1766
rect 21362 1712 21550 1732
rect 21300 1676 21550 1712
rect 21300 1656 21477 1676
rect 21300 1622 21328 1656
rect 21362 1642 21477 1656
rect 21511 1642 21550 1676
rect 21362 1622 21550 1642
rect 21300 1586 21550 1622
rect 21300 1566 21477 1586
rect 21300 1532 21328 1566
rect 21362 1552 21477 1566
rect 21511 1552 21550 1586
rect 21362 1532 21550 1552
rect 21300 1496 21550 1532
rect 21300 1476 21477 1496
rect 21300 1442 21328 1476
rect 21362 1462 21477 1476
rect 21511 1462 21550 1496
rect 21362 1442 21550 1462
rect 21300 1406 21550 1442
rect 21300 1386 21477 1406
rect 21300 1352 21328 1386
rect 21362 1372 21477 1386
rect 21511 1372 21550 1406
rect 21362 1352 21550 1372
rect 21300 1316 21550 1352
rect 21300 1296 21477 1316
rect 20419 1221 20491 1281
rect 21300 1262 21328 1296
rect 21362 1282 21477 1296
rect 21511 1282 21550 1316
rect 21362 1262 21550 1282
rect 21300 1226 21550 1262
rect 21300 1221 21477 1226
rect 20419 1202 21477 1221
rect 20419 1168 20516 1202
rect 20550 1168 20606 1202
rect 20640 1168 20696 1202
rect 20730 1168 20786 1202
rect 20820 1168 20876 1202
rect 20910 1168 20966 1202
rect 21000 1168 21056 1202
rect 21090 1168 21146 1202
rect 21180 1168 21236 1202
rect 21270 1192 21477 1202
rect 21511 1192 21550 1226
rect 21270 1168 21550 1192
rect 20419 1149 21550 1168
rect 20256 1102 20290 1136
rect 20324 1102 20355 1136
rect 20256 1085 20355 1102
rect 21300 1136 21550 1149
rect 21300 1102 21477 1136
rect 21511 1102 21550 1136
rect 21300 1085 21550 1102
rect 20256 1052 21550 1085
rect 20256 1018 20386 1052
rect 20420 1018 20476 1052
rect 20510 1018 20566 1052
rect 20600 1018 20656 1052
rect 20690 1018 20746 1052
rect 20780 1018 20836 1052
rect 20870 1018 20926 1052
rect 20960 1018 21016 1052
rect 21050 1018 21106 1052
rect 21140 1018 21196 1052
rect 21230 1018 21286 1052
rect 21320 1018 21376 1052
rect 21410 1018 21550 1052
rect 20256 986 21550 1018
rect 21616 2239 22910 2270
rect 21616 2216 21746 2239
rect 21616 2182 21650 2216
rect 21684 2205 21746 2216
rect 21780 2205 21836 2239
rect 21870 2205 21926 2239
rect 21960 2205 22016 2239
rect 22050 2205 22106 2239
rect 22140 2205 22196 2239
rect 22230 2205 22286 2239
rect 22320 2205 22376 2239
rect 22410 2205 22466 2239
rect 22500 2205 22556 2239
rect 22590 2205 22646 2239
rect 22680 2205 22736 2239
rect 22770 2216 22910 2239
rect 22770 2205 22837 2216
rect 21684 2182 22837 2205
rect 22871 2182 22910 2216
rect 21616 2175 22910 2182
rect 21616 2126 21715 2175
rect 21616 2092 21650 2126
rect 21684 2092 21715 2126
rect 22660 2126 22910 2175
rect 22660 2111 22837 2126
rect 21616 2036 21715 2092
rect 21616 2002 21650 2036
rect 21684 2002 21715 2036
rect 21616 1946 21715 2002
rect 21616 1912 21650 1946
rect 21684 1912 21715 1946
rect 21616 1856 21715 1912
rect 21616 1822 21650 1856
rect 21684 1822 21715 1856
rect 21616 1766 21715 1822
rect 21616 1732 21650 1766
rect 21684 1732 21715 1766
rect 21616 1676 21715 1732
rect 21616 1642 21650 1676
rect 21684 1642 21715 1676
rect 21616 1586 21715 1642
rect 21616 1552 21650 1586
rect 21684 1552 21715 1586
rect 21616 1496 21715 1552
rect 21616 1462 21650 1496
rect 21684 1462 21715 1496
rect 21616 1406 21715 1462
rect 21616 1372 21650 1406
rect 21684 1372 21715 1406
rect 21616 1316 21715 1372
rect 21616 1282 21650 1316
rect 21684 1282 21715 1316
rect 21616 1226 21715 1282
rect 21616 1192 21650 1226
rect 21684 1192 21715 1226
rect 21616 1136 21715 1192
rect 21779 2092 22837 2111
rect 22871 2092 22910 2126
rect 21779 2058 21910 2092
rect 21944 2058 22000 2092
rect 22034 2058 22090 2092
rect 22124 2058 22180 2092
rect 22214 2058 22270 2092
rect 22304 2058 22360 2092
rect 22394 2058 22450 2092
rect 22484 2058 22540 2092
rect 22574 2058 22630 2092
rect 22664 2058 22910 2092
rect 21779 2039 22910 2058
rect 21779 2035 21851 2039
rect 21779 2001 21798 2035
rect 21832 2001 21851 2035
rect 21779 1945 21851 2001
rect 22660 2036 22910 2039
rect 22660 2016 22837 2036
rect 22660 1982 22688 2016
rect 22722 2002 22837 2016
rect 22871 2002 22910 2036
rect 22722 1982 22910 2002
rect 21779 1911 21798 1945
rect 21832 1911 21851 1945
rect 21779 1855 21851 1911
rect 21779 1821 21798 1855
rect 21832 1821 21851 1855
rect 21779 1765 21851 1821
rect 21779 1731 21798 1765
rect 21832 1731 21851 1765
rect 21779 1675 21851 1731
rect 21779 1641 21798 1675
rect 21832 1641 21851 1675
rect 21779 1585 21851 1641
rect 21779 1551 21798 1585
rect 21832 1551 21851 1585
rect 21779 1495 21851 1551
rect 21779 1461 21798 1495
rect 21832 1461 21851 1495
rect 21779 1405 21851 1461
rect 21779 1371 21798 1405
rect 21832 1371 21851 1405
rect 21779 1315 21851 1371
rect 21779 1281 21798 1315
rect 21832 1281 21851 1315
rect 21913 1918 22607 1977
rect 21913 1884 21974 1918
rect 22008 1890 22064 1918
rect 22098 1890 22154 1918
rect 22188 1890 22244 1918
rect 22020 1884 22064 1890
rect 22120 1884 22154 1890
rect 22220 1884 22244 1890
rect 22278 1890 22334 1918
rect 22278 1884 22286 1890
rect 21913 1856 21986 1884
rect 22020 1856 22086 1884
rect 22120 1856 22186 1884
rect 22220 1856 22286 1884
rect 22320 1884 22334 1890
rect 22368 1890 22424 1918
rect 22368 1884 22386 1890
rect 22320 1856 22386 1884
rect 22420 1884 22424 1890
rect 22458 1890 22514 1918
rect 22458 1884 22486 1890
rect 22548 1884 22607 1918
rect 22420 1856 22486 1884
rect 22520 1856 22607 1884
rect 21913 1828 22607 1856
rect 21913 1794 21974 1828
rect 22008 1794 22064 1828
rect 22098 1794 22154 1828
rect 22188 1794 22244 1828
rect 22278 1794 22334 1828
rect 22368 1794 22424 1828
rect 22458 1794 22514 1828
rect 22548 1794 22607 1828
rect 21913 1790 22607 1794
rect 21913 1756 21986 1790
rect 22020 1756 22086 1790
rect 22120 1756 22186 1790
rect 22220 1756 22286 1790
rect 22320 1756 22386 1790
rect 22420 1756 22486 1790
rect 22520 1756 22607 1790
rect 21913 1738 22607 1756
rect 21913 1704 21974 1738
rect 22008 1704 22064 1738
rect 22098 1704 22154 1738
rect 22188 1704 22244 1738
rect 22278 1704 22334 1738
rect 22368 1704 22424 1738
rect 22458 1704 22514 1738
rect 22548 1704 22607 1738
rect 21913 1690 22607 1704
rect 21913 1656 21986 1690
rect 22020 1656 22086 1690
rect 22120 1656 22186 1690
rect 22220 1656 22286 1690
rect 22320 1656 22386 1690
rect 22420 1656 22486 1690
rect 22520 1656 22607 1690
rect 21913 1648 22607 1656
rect 21913 1614 21974 1648
rect 22008 1614 22064 1648
rect 22098 1614 22154 1648
rect 22188 1614 22244 1648
rect 22278 1614 22334 1648
rect 22368 1614 22424 1648
rect 22458 1614 22514 1648
rect 22548 1614 22607 1648
rect 21913 1590 22607 1614
rect 21913 1558 21986 1590
rect 22020 1558 22086 1590
rect 22120 1558 22186 1590
rect 22220 1558 22286 1590
rect 21913 1524 21974 1558
rect 22020 1556 22064 1558
rect 22120 1556 22154 1558
rect 22220 1556 22244 1558
rect 22008 1524 22064 1556
rect 22098 1524 22154 1556
rect 22188 1524 22244 1556
rect 22278 1556 22286 1558
rect 22320 1558 22386 1590
rect 22320 1556 22334 1558
rect 22278 1524 22334 1556
rect 22368 1556 22386 1558
rect 22420 1558 22486 1590
rect 22520 1558 22607 1590
rect 22420 1556 22424 1558
rect 22368 1524 22424 1556
rect 22458 1556 22486 1558
rect 22458 1524 22514 1556
rect 22548 1524 22607 1558
rect 21913 1490 22607 1524
rect 21913 1468 21986 1490
rect 22020 1468 22086 1490
rect 22120 1468 22186 1490
rect 22220 1468 22286 1490
rect 21913 1434 21974 1468
rect 22020 1456 22064 1468
rect 22120 1456 22154 1468
rect 22220 1456 22244 1468
rect 22008 1434 22064 1456
rect 22098 1434 22154 1456
rect 22188 1434 22244 1456
rect 22278 1456 22286 1468
rect 22320 1468 22386 1490
rect 22320 1456 22334 1468
rect 22278 1434 22334 1456
rect 22368 1456 22386 1468
rect 22420 1468 22486 1490
rect 22520 1468 22607 1490
rect 22420 1456 22424 1468
rect 22368 1434 22424 1456
rect 22458 1456 22486 1468
rect 22458 1434 22514 1456
rect 22548 1434 22607 1468
rect 21913 1390 22607 1434
rect 21913 1378 21986 1390
rect 22020 1378 22086 1390
rect 22120 1378 22186 1390
rect 22220 1378 22286 1390
rect 21913 1344 21974 1378
rect 22020 1356 22064 1378
rect 22120 1356 22154 1378
rect 22220 1356 22244 1378
rect 22008 1344 22064 1356
rect 22098 1344 22154 1356
rect 22188 1344 22244 1356
rect 22278 1356 22286 1378
rect 22320 1378 22386 1390
rect 22320 1356 22334 1378
rect 22278 1344 22334 1356
rect 22368 1356 22386 1378
rect 22420 1378 22486 1390
rect 22520 1378 22607 1390
rect 22420 1356 22424 1378
rect 22368 1344 22424 1356
rect 22458 1356 22486 1378
rect 22458 1344 22514 1356
rect 22548 1344 22607 1378
rect 21913 1283 22607 1344
rect 22660 1946 22910 1982
rect 22660 1926 22837 1946
rect 22660 1892 22688 1926
rect 22722 1912 22837 1926
rect 22871 1912 22910 1946
rect 22722 1892 22910 1912
rect 22660 1856 22910 1892
rect 22660 1836 22837 1856
rect 22660 1802 22688 1836
rect 22722 1822 22837 1836
rect 22871 1822 22910 1856
rect 22722 1802 22910 1822
rect 22660 1766 22910 1802
rect 22660 1746 22837 1766
rect 22660 1712 22688 1746
rect 22722 1732 22837 1746
rect 22871 1732 22910 1766
rect 22722 1712 22910 1732
rect 22660 1676 22910 1712
rect 22660 1656 22837 1676
rect 22660 1622 22688 1656
rect 22722 1642 22837 1656
rect 22871 1642 22910 1676
rect 22722 1622 22910 1642
rect 22660 1586 22910 1622
rect 22660 1566 22837 1586
rect 22660 1532 22688 1566
rect 22722 1552 22837 1566
rect 22871 1552 22910 1586
rect 22722 1532 22910 1552
rect 22660 1496 22910 1532
rect 22660 1476 22837 1496
rect 22660 1442 22688 1476
rect 22722 1462 22837 1476
rect 22871 1462 22910 1496
rect 22722 1442 22910 1462
rect 22660 1406 22910 1442
rect 22660 1386 22837 1406
rect 22660 1352 22688 1386
rect 22722 1372 22837 1386
rect 22871 1372 22910 1406
rect 22722 1352 22910 1372
rect 22660 1316 22910 1352
rect 22660 1296 22837 1316
rect 21779 1221 21851 1281
rect 22660 1262 22688 1296
rect 22722 1282 22837 1296
rect 22871 1282 22910 1316
rect 22722 1262 22910 1282
rect 22660 1226 22910 1262
rect 22660 1221 22837 1226
rect 21779 1202 22837 1221
rect 21779 1168 21876 1202
rect 21910 1168 21966 1202
rect 22000 1168 22056 1202
rect 22090 1168 22146 1202
rect 22180 1168 22236 1202
rect 22270 1168 22326 1202
rect 22360 1168 22416 1202
rect 22450 1168 22506 1202
rect 22540 1168 22596 1202
rect 22630 1192 22837 1202
rect 22871 1192 22910 1226
rect 22630 1168 22910 1192
rect 21779 1149 22910 1168
rect 21616 1102 21650 1136
rect 21684 1102 21715 1136
rect 21616 1085 21715 1102
rect 22660 1136 22910 1149
rect 22660 1102 22837 1136
rect 22871 1102 22910 1136
rect 22660 1085 22910 1102
rect 21616 1052 22910 1085
rect 21616 1018 21746 1052
rect 21780 1018 21836 1052
rect 21870 1018 21926 1052
rect 21960 1018 22016 1052
rect 22050 1018 22106 1052
rect 22140 1018 22196 1052
rect 22230 1018 22286 1052
rect 22320 1018 22376 1052
rect 22410 1018 22466 1052
rect 22500 1018 22556 1052
rect 22590 1018 22646 1052
rect 22680 1018 22736 1052
rect 22770 1018 22910 1052
rect 21616 986 22910 1018
rect 22976 2239 24270 2270
rect 22976 2216 23106 2239
rect 22976 2182 23010 2216
rect 23044 2205 23106 2216
rect 23140 2205 23196 2239
rect 23230 2205 23286 2239
rect 23320 2205 23376 2239
rect 23410 2205 23466 2239
rect 23500 2205 23556 2239
rect 23590 2205 23646 2239
rect 23680 2205 23736 2239
rect 23770 2205 23826 2239
rect 23860 2205 23916 2239
rect 23950 2205 24006 2239
rect 24040 2205 24096 2239
rect 24130 2216 24270 2239
rect 24130 2205 24197 2216
rect 23044 2182 24197 2205
rect 24231 2182 24270 2216
rect 22976 2175 24270 2182
rect 22976 2126 23075 2175
rect 22976 2092 23010 2126
rect 23044 2092 23075 2126
rect 24020 2126 24270 2175
rect 24020 2111 24197 2126
rect 22976 2036 23075 2092
rect 22976 2002 23010 2036
rect 23044 2002 23075 2036
rect 22976 1946 23075 2002
rect 22976 1912 23010 1946
rect 23044 1912 23075 1946
rect 22976 1856 23075 1912
rect 22976 1822 23010 1856
rect 23044 1822 23075 1856
rect 22976 1766 23075 1822
rect 22976 1732 23010 1766
rect 23044 1732 23075 1766
rect 22976 1676 23075 1732
rect 22976 1642 23010 1676
rect 23044 1642 23075 1676
rect 22976 1586 23075 1642
rect 22976 1552 23010 1586
rect 23044 1552 23075 1586
rect 22976 1496 23075 1552
rect 22976 1462 23010 1496
rect 23044 1462 23075 1496
rect 22976 1406 23075 1462
rect 22976 1372 23010 1406
rect 23044 1372 23075 1406
rect 22976 1316 23075 1372
rect 22976 1282 23010 1316
rect 23044 1282 23075 1316
rect 22976 1226 23075 1282
rect 22976 1192 23010 1226
rect 23044 1192 23075 1226
rect 22976 1136 23075 1192
rect 23139 2092 24197 2111
rect 24231 2092 24270 2126
rect 23139 2058 23270 2092
rect 23304 2058 23360 2092
rect 23394 2058 23450 2092
rect 23484 2058 23540 2092
rect 23574 2058 23630 2092
rect 23664 2058 23720 2092
rect 23754 2058 23810 2092
rect 23844 2058 23900 2092
rect 23934 2058 23990 2092
rect 24024 2058 24270 2092
rect 23139 2039 24270 2058
rect 23139 2035 23211 2039
rect 23139 2001 23158 2035
rect 23192 2001 23211 2035
rect 23139 1945 23211 2001
rect 24020 2036 24270 2039
rect 24020 2016 24197 2036
rect 24020 1982 24048 2016
rect 24082 2002 24197 2016
rect 24231 2002 24270 2036
rect 25690 2840 26830 2880
rect 26990 2840 28130 2880
rect 25690 2530 25730 2840
rect 25970 2780 26050 2800
rect 25790 2750 25870 2770
rect 25790 2710 25810 2750
rect 25850 2710 25870 2750
rect 25970 2740 25990 2780
rect 26030 2740 26050 2780
rect 25970 2720 26050 2740
rect 26210 2780 26290 2800
rect 26210 2740 26230 2780
rect 26270 2740 26290 2780
rect 26210 2720 26290 2740
rect 26450 2780 26530 2800
rect 26450 2740 26470 2780
rect 26510 2740 26530 2780
rect 26450 2720 26530 2740
rect 26690 2780 26770 2800
rect 26690 2740 26710 2780
rect 26750 2740 26770 2780
rect 26690 2720 26770 2740
rect 27170 2780 27250 2800
rect 27170 2740 27190 2780
rect 27230 2740 27250 2780
rect 27170 2720 27250 2740
rect 27410 2780 27490 2800
rect 27410 2740 27430 2780
rect 27470 2740 27490 2780
rect 27410 2720 27490 2740
rect 27650 2780 27730 2800
rect 27650 2740 27670 2780
rect 27710 2740 27730 2780
rect 27650 2720 27730 2740
rect 27950 2750 28030 2770
rect 25790 2690 25870 2710
rect 27950 2710 27970 2750
rect 28010 2710 28030 2750
rect 27950 2690 28030 2710
rect 25690 2050 25730 2370
rect 25800 2670 25860 2690
rect 25800 2630 25810 2670
rect 25850 2630 25860 2670
rect 25800 2570 25860 2630
rect 25800 2530 25810 2570
rect 25850 2530 25860 2570
rect 25800 2470 25860 2530
rect 25800 2430 25810 2470
rect 25850 2430 25860 2470
rect 25800 2370 25860 2430
rect 25800 2330 25810 2370
rect 25850 2330 25860 2370
rect 25800 2270 25860 2330
rect 25800 2230 25810 2270
rect 25850 2230 25860 2270
rect 25800 2210 25860 2230
rect 26880 2670 26940 2690
rect 26880 2630 26890 2670
rect 26930 2630 26940 2670
rect 26880 2570 26940 2630
rect 26880 2530 26890 2570
rect 26930 2530 26940 2570
rect 26880 2470 26940 2530
rect 26880 2430 26890 2470
rect 26930 2430 26940 2470
rect 26880 2370 26940 2430
rect 26880 2330 26890 2370
rect 26930 2330 26940 2370
rect 26880 2270 26940 2330
rect 26880 2230 26890 2270
rect 26930 2230 26940 2270
rect 26880 2210 26940 2230
rect 27960 2670 28020 2690
rect 27960 2630 27970 2670
rect 28010 2630 28020 2670
rect 27960 2570 28020 2630
rect 27960 2530 27970 2570
rect 28010 2530 28020 2570
rect 27960 2470 28020 2530
rect 27960 2430 27970 2470
rect 28010 2430 28020 2470
rect 27960 2370 28020 2430
rect 27960 2330 27970 2370
rect 28010 2330 28020 2370
rect 27960 2270 28020 2330
rect 27960 2230 27970 2270
rect 28010 2230 28020 2270
rect 27960 2210 28020 2230
rect 28090 2530 28130 2840
rect 26890 2170 26930 2210
rect 26870 2150 26950 2170
rect 26870 2110 26890 2150
rect 26930 2110 26950 2150
rect 26870 2090 26950 2110
rect 28090 2050 28130 2370
rect 25690 2010 26830 2050
rect 26990 2010 28130 2050
rect 28210 2840 29350 2880
rect 29510 2840 30650 2880
rect 28210 2530 28250 2840
rect 28610 2780 28690 2800
rect 28310 2750 28390 2770
rect 28310 2710 28330 2750
rect 28370 2710 28390 2750
rect 28610 2740 28630 2780
rect 28670 2740 28690 2780
rect 28610 2720 28690 2740
rect 28850 2780 28930 2800
rect 28850 2740 28870 2780
rect 28910 2740 28930 2780
rect 28850 2720 28930 2740
rect 29090 2780 29170 2800
rect 29090 2740 29110 2780
rect 29150 2740 29170 2780
rect 29090 2720 29170 2740
rect 29570 2780 29650 2800
rect 29570 2740 29590 2780
rect 29630 2740 29650 2780
rect 29570 2720 29650 2740
rect 29810 2780 29890 2800
rect 29810 2740 29830 2780
rect 29870 2740 29890 2780
rect 29810 2720 29890 2740
rect 30050 2780 30130 2800
rect 30050 2740 30070 2780
rect 30110 2740 30130 2780
rect 30050 2720 30130 2740
rect 30290 2780 30370 2800
rect 30290 2740 30310 2780
rect 30350 2740 30370 2780
rect 30290 2720 30370 2740
rect 30470 2750 30550 2770
rect 28310 2690 28390 2710
rect 30470 2710 30490 2750
rect 30530 2710 30550 2750
rect 30470 2690 30550 2710
rect 28210 2050 28250 2370
rect 28320 2670 28380 2690
rect 28320 2630 28330 2670
rect 28370 2630 28380 2670
rect 28320 2570 28380 2630
rect 28320 2530 28330 2570
rect 28370 2530 28380 2570
rect 28320 2470 28380 2530
rect 28320 2430 28330 2470
rect 28370 2430 28380 2470
rect 28320 2370 28380 2430
rect 28320 2330 28330 2370
rect 28370 2330 28380 2370
rect 28320 2270 28380 2330
rect 28320 2230 28330 2270
rect 28370 2230 28380 2270
rect 28320 2210 28380 2230
rect 29400 2670 29460 2690
rect 29400 2630 29410 2670
rect 29450 2630 29460 2670
rect 29400 2570 29460 2630
rect 29400 2530 29410 2570
rect 29450 2530 29460 2570
rect 29400 2470 29460 2530
rect 29400 2430 29410 2470
rect 29450 2430 29460 2470
rect 29400 2370 29460 2430
rect 29400 2330 29410 2370
rect 29450 2330 29460 2370
rect 29400 2270 29460 2330
rect 29400 2230 29410 2270
rect 29450 2230 29460 2270
rect 29400 2210 29460 2230
rect 30480 2670 30540 2690
rect 30480 2630 30490 2670
rect 30530 2630 30540 2670
rect 30480 2570 30540 2630
rect 30480 2530 30490 2570
rect 30530 2530 30540 2570
rect 30480 2470 30540 2530
rect 30480 2430 30490 2470
rect 30530 2430 30540 2470
rect 30480 2370 30540 2430
rect 30480 2330 30490 2370
rect 30530 2330 30540 2370
rect 30480 2270 30540 2330
rect 30480 2230 30490 2270
rect 30530 2230 30540 2270
rect 30480 2210 30540 2230
rect 30610 2530 30650 2840
rect 29410 2170 29450 2210
rect 29390 2150 29470 2170
rect 29390 2110 29410 2150
rect 29450 2110 29470 2150
rect 29390 2090 29470 2110
rect 30610 2050 30650 2370
rect 28210 2010 29350 2050
rect 29510 2010 30650 2050
rect 24082 1982 24270 2002
rect 23139 1911 23158 1945
rect 23192 1911 23211 1945
rect 23139 1855 23211 1911
rect 23139 1821 23158 1855
rect 23192 1821 23211 1855
rect 23139 1765 23211 1821
rect 23139 1731 23158 1765
rect 23192 1731 23211 1765
rect 23139 1675 23211 1731
rect 23139 1641 23158 1675
rect 23192 1641 23211 1675
rect 23139 1585 23211 1641
rect 23139 1551 23158 1585
rect 23192 1551 23211 1585
rect 23139 1495 23211 1551
rect 23139 1461 23158 1495
rect 23192 1461 23211 1495
rect 23139 1405 23211 1461
rect 23139 1371 23158 1405
rect 23192 1371 23211 1405
rect 23139 1315 23211 1371
rect 23139 1281 23158 1315
rect 23192 1281 23211 1315
rect 23273 1918 23967 1977
rect 23273 1884 23334 1918
rect 23368 1890 23424 1918
rect 23458 1890 23514 1918
rect 23548 1890 23604 1918
rect 23380 1884 23424 1890
rect 23480 1884 23514 1890
rect 23580 1884 23604 1890
rect 23638 1890 23694 1918
rect 23638 1884 23646 1890
rect 23273 1856 23346 1884
rect 23380 1856 23446 1884
rect 23480 1856 23546 1884
rect 23580 1856 23646 1884
rect 23680 1884 23694 1890
rect 23728 1890 23784 1918
rect 23728 1884 23746 1890
rect 23680 1856 23746 1884
rect 23780 1884 23784 1890
rect 23818 1890 23874 1918
rect 23818 1884 23846 1890
rect 23908 1884 23967 1918
rect 23780 1856 23846 1884
rect 23880 1856 23967 1884
rect 23273 1828 23967 1856
rect 23273 1794 23334 1828
rect 23368 1794 23424 1828
rect 23458 1794 23514 1828
rect 23548 1794 23604 1828
rect 23638 1794 23694 1828
rect 23728 1794 23784 1828
rect 23818 1794 23874 1828
rect 23908 1794 23967 1828
rect 23273 1790 23967 1794
rect 23273 1756 23346 1790
rect 23380 1756 23446 1790
rect 23480 1756 23546 1790
rect 23580 1756 23646 1790
rect 23680 1756 23746 1790
rect 23780 1756 23846 1790
rect 23880 1756 23967 1790
rect 23273 1738 23967 1756
rect 23273 1704 23334 1738
rect 23368 1704 23424 1738
rect 23458 1704 23514 1738
rect 23548 1704 23604 1738
rect 23638 1704 23694 1738
rect 23728 1704 23784 1738
rect 23818 1704 23874 1738
rect 23908 1704 23967 1738
rect 23273 1690 23967 1704
rect 23273 1656 23346 1690
rect 23380 1656 23446 1690
rect 23480 1656 23546 1690
rect 23580 1656 23646 1690
rect 23680 1656 23746 1690
rect 23780 1656 23846 1690
rect 23880 1656 23967 1690
rect 23273 1648 23967 1656
rect 23273 1614 23334 1648
rect 23368 1614 23424 1648
rect 23458 1614 23514 1648
rect 23548 1614 23604 1648
rect 23638 1614 23694 1648
rect 23728 1614 23784 1648
rect 23818 1614 23874 1648
rect 23908 1614 23967 1648
rect 23273 1590 23967 1614
rect 23273 1558 23346 1590
rect 23380 1558 23446 1590
rect 23480 1558 23546 1590
rect 23580 1558 23646 1590
rect 23273 1524 23334 1558
rect 23380 1556 23424 1558
rect 23480 1556 23514 1558
rect 23580 1556 23604 1558
rect 23368 1524 23424 1556
rect 23458 1524 23514 1556
rect 23548 1524 23604 1556
rect 23638 1556 23646 1558
rect 23680 1558 23746 1590
rect 23680 1556 23694 1558
rect 23638 1524 23694 1556
rect 23728 1556 23746 1558
rect 23780 1558 23846 1590
rect 23880 1558 23967 1590
rect 23780 1556 23784 1558
rect 23728 1524 23784 1556
rect 23818 1556 23846 1558
rect 23818 1524 23874 1556
rect 23908 1524 23967 1558
rect 23273 1490 23967 1524
rect 23273 1468 23346 1490
rect 23380 1468 23446 1490
rect 23480 1468 23546 1490
rect 23580 1468 23646 1490
rect 23273 1434 23334 1468
rect 23380 1456 23424 1468
rect 23480 1456 23514 1468
rect 23580 1456 23604 1468
rect 23368 1434 23424 1456
rect 23458 1434 23514 1456
rect 23548 1434 23604 1456
rect 23638 1456 23646 1468
rect 23680 1468 23746 1490
rect 23680 1456 23694 1468
rect 23638 1434 23694 1456
rect 23728 1456 23746 1468
rect 23780 1468 23846 1490
rect 23880 1468 23967 1490
rect 23780 1456 23784 1468
rect 23728 1434 23784 1456
rect 23818 1456 23846 1468
rect 23818 1434 23874 1456
rect 23908 1434 23967 1468
rect 23273 1390 23967 1434
rect 23273 1378 23346 1390
rect 23380 1378 23446 1390
rect 23480 1378 23546 1390
rect 23580 1378 23646 1390
rect 23273 1344 23334 1378
rect 23380 1356 23424 1378
rect 23480 1356 23514 1378
rect 23580 1356 23604 1378
rect 23368 1344 23424 1356
rect 23458 1344 23514 1356
rect 23548 1344 23604 1356
rect 23638 1356 23646 1378
rect 23680 1378 23746 1390
rect 23680 1356 23694 1378
rect 23638 1344 23694 1356
rect 23728 1356 23746 1378
rect 23780 1378 23846 1390
rect 23880 1378 23967 1390
rect 23780 1356 23784 1378
rect 23728 1344 23784 1356
rect 23818 1356 23846 1378
rect 23818 1344 23874 1356
rect 23908 1344 23967 1378
rect 23273 1283 23967 1344
rect 24020 1946 24270 1982
rect 24020 1926 24197 1946
rect 24020 1892 24048 1926
rect 24082 1912 24197 1926
rect 24231 1912 24270 1946
rect 24082 1892 24270 1912
rect 24020 1856 24270 1892
rect 24020 1836 24197 1856
rect 24020 1802 24048 1836
rect 24082 1822 24197 1836
rect 24231 1822 24270 1856
rect 24082 1802 24270 1822
rect 24020 1766 24270 1802
rect 24020 1746 24197 1766
rect 24020 1712 24048 1746
rect 24082 1732 24197 1746
rect 24231 1732 24270 1766
rect 24082 1712 24270 1732
rect 24020 1676 24270 1712
rect 24020 1656 24197 1676
rect 24020 1622 24048 1656
rect 24082 1642 24197 1656
rect 24231 1642 24270 1676
rect 24082 1622 24270 1642
rect 25890 1860 28090 1900
rect 28250 1860 30530 1900
rect 25890 1690 25930 1860
rect 26050 1800 26130 1820
rect 26050 1760 26070 1800
rect 26110 1760 26130 1800
rect 26050 1740 26130 1760
rect 26210 1800 26290 1820
rect 26210 1760 26230 1800
rect 26270 1760 26290 1800
rect 26210 1740 26290 1760
rect 26370 1800 26450 1820
rect 26370 1760 26390 1800
rect 26430 1760 26450 1800
rect 26370 1740 26450 1760
rect 26530 1800 26610 1820
rect 26530 1760 26550 1800
rect 26590 1760 26610 1800
rect 26530 1740 26610 1760
rect 26690 1800 26770 1820
rect 26690 1760 26710 1800
rect 26750 1760 26770 1800
rect 26690 1740 26770 1760
rect 26850 1800 26930 1820
rect 26850 1760 26870 1800
rect 26910 1760 26930 1800
rect 26850 1740 26930 1760
rect 27010 1800 27090 1820
rect 27010 1760 27030 1800
rect 27070 1760 27090 1800
rect 27010 1740 27090 1760
rect 27170 1800 27250 1820
rect 27170 1760 27190 1800
rect 27230 1760 27250 1800
rect 27170 1740 27250 1760
rect 27330 1800 27410 1820
rect 27330 1760 27350 1800
rect 27390 1760 27410 1800
rect 27330 1740 27410 1760
rect 27490 1800 27570 1820
rect 27490 1760 27510 1800
rect 27550 1760 27570 1800
rect 27490 1740 27570 1760
rect 27650 1800 27730 1820
rect 27650 1760 27670 1800
rect 27710 1760 27730 1800
rect 27650 1740 27730 1760
rect 27810 1800 27890 1820
rect 27810 1760 27830 1800
rect 27870 1760 27890 1800
rect 27810 1740 27890 1760
rect 27970 1800 28050 1820
rect 27970 1760 27990 1800
rect 28030 1760 28050 1800
rect 27970 1740 28050 1760
rect 28130 1800 28210 1820
rect 28130 1760 28150 1800
rect 28190 1760 28210 1800
rect 28130 1740 28210 1760
rect 28290 1800 28370 1820
rect 28290 1760 28310 1800
rect 28350 1760 28370 1800
rect 28290 1740 28370 1760
rect 28450 1800 28530 1820
rect 28450 1760 28470 1800
rect 28510 1760 28530 1800
rect 28450 1740 28530 1760
rect 28610 1800 28690 1820
rect 28610 1760 28630 1800
rect 28670 1760 28690 1800
rect 28610 1740 28690 1760
rect 28770 1800 28850 1820
rect 28770 1760 28790 1800
rect 28830 1760 28850 1800
rect 28770 1740 28850 1760
rect 28930 1800 29010 1820
rect 28930 1760 28950 1800
rect 28990 1760 29010 1800
rect 28930 1740 29010 1760
rect 29090 1800 29170 1820
rect 29090 1760 29110 1800
rect 29150 1760 29170 1800
rect 29090 1740 29170 1760
rect 29250 1800 29330 1820
rect 29250 1760 29270 1800
rect 29310 1760 29330 1800
rect 29250 1740 29330 1760
rect 29410 1800 29490 1820
rect 29410 1760 29430 1800
rect 29470 1760 29490 1800
rect 29410 1740 29490 1760
rect 29570 1800 29650 1820
rect 29570 1760 29590 1800
rect 29630 1760 29650 1800
rect 29570 1740 29650 1760
rect 29730 1800 29810 1820
rect 29730 1760 29750 1800
rect 29790 1760 29810 1800
rect 29730 1740 29810 1760
rect 29890 1800 29970 1820
rect 29890 1760 29910 1800
rect 29950 1760 29970 1800
rect 29890 1740 29970 1760
rect 30050 1800 30130 1820
rect 30050 1760 30070 1800
rect 30110 1760 30130 1800
rect 30050 1740 30130 1760
rect 26070 1700 26110 1740
rect 28150 1700 28190 1740
rect 24020 1586 24270 1622
rect 24020 1566 24197 1586
rect 24020 1532 24048 1566
rect 24082 1552 24197 1566
rect 24231 1552 24270 1586
rect 25160 1580 25220 1640
rect 24082 1532 24270 1552
rect 24020 1496 24270 1532
rect 24020 1476 24197 1496
rect 24020 1442 24048 1476
rect 24082 1462 24197 1476
rect 24231 1462 24270 1496
rect 24082 1442 24270 1462
rect 24020 1406 24270 1442
rect 26060 1680 26120 1700
rect 26060 1650 26070 1680
rect 25970 1640 26070 1650
rect 26110 1640 26120 1680
rect 25970 1630 26120 1640
rect 25970 1590 25990 1630
rect 26030 1590 26120 1630
rect 25970 1580 26120 1590
rect 25970 1570 26070 1580
rect 25890 1450 25930 1530
rect 26060 1540 26070 1570
rect 26110 1540 26120 1580
rect 26060 1520 26120 1540
rect 28140 1680 28200 1700
rect 28140 1640 28150 1680
rect 28190 1640 28200 1680
rect 28140 1580 28200 1640
rect 28140 1540 28150 1580
rect 28190 1540 28200 1580
rect 28140 1520 28200 1540
rect 30220 1680 30360 1700
rect 30220 1640 30230 1680
rect 30270 1640 30310 1680
rect 30350 1650 30360 1680
rect 30490 1690 30530 1860
rect 30350 1640 30450 1650
rect 30220 1630 30450 1640
rect 30220 1590 30390 1630
rect 30430 1590 30450 1630
rect 30220 1580 30450 1590
rect 30220 1540 30230 1580
rect 30270 1540 30310 1580
rect 30350 1570 30450 1580
rect 30350 1540 30360 1570
rect 30220 1520 30360 1540
rect 30490 1450 30530 1530
rect 25890 1410 28090 1450
rect 28250 1410 30530 1450
rect 24020 1386 24197 1406
rect 24020 1352 24048 1386
rect 24082 1372 24197 1386
rect 24231 1372 24270 1406
rect 24082 1352 24270 1372
rect 24020 1316 24270 1352
rect 24020 1296 24197 1316
rect 23139 1221 23211 1281
rect 24020 1262 24048 1296
rect 24082 1282 24197 1296
rect 24231 1282 24270 1316
rect 24082 1262 24270 1282
rect 24020 1226 24270 1262
rect 24020 1221 24197 1226
rect 23139 1202 24197 1221
rect 23139 1168 23236 1202
rect 23270 1168 23326 1202
rect 23360 1168 23416 1202
rect 23450 1168 23506 1202
rect 23540 1168 23596 1202
rect 23630 1168 23686 1202
rect 23720 1168 23776 1202
rect 23810 1168 23866 1202
rect 23900 1168 23956 1202
rect 23990 1192 24197 1202
rect 24231 1192 24270 1226
rect 23990 1168 24270 1192
rect 23139 1149 24270 1168
rect 22976 1102 23010 1136
rect 23044 1102 23075 1136
rect 22976 1085 23075 1102
rect 24020 1136 24270 1149
rect 24020 1102 24197 1136
rect 24231 1102 24270 1136
rect 24020 1085 24270 1102
rect 22976 1052 24270 1085
rect 22976 1018 23106 1052
rect 23140 1018 23196 1052
rect 23230 1018 23286 1052
rect 23320 1018 23376 1052
rect 23410 1018 23466 1052
rect 23500 1018 23556 1052
rect 23590 1018 23646 1052
rect 23680 1018 23736 1052
rect 23770 1018 23826 1052
rect 23860 1018 23916 1052
rect 23950 1018 24006 1052
rect 24040 1018 24096 1052
rect 24130 1018 24270 1052
rect 22976 990 24270 1018
rect 25290 1310 26070 1350
rect 26230 1310 27010 1350
rect 25290 1140 25330 1310
rect 25750 1250 25830 1270
rect 25750 1210 25770 1250
rect 25810 1210 25830 1250
rect 25750 1190 25830 1210
rect 26110 1250 26190 1270
rect 26110 1210 26130 1250
rect 26170 1210 26190 1250
rect 26110 1190 26190 1210
rect 26470 1250 26550 1270
rect 26470 1210 26490 1250
rect 26530 1210 26550 1250
rect 26470 1190 26550 1210
rect 25770 1150 25810 1190
rect 26130 1150 26170 1190
rect 26490 1150 26530 1190
rect 22976 986 24264 990
rect 21300 980 21550 986
rect 22660 980 22910 986
rect 25290 810 25330 980
rect 25400 1130 25460 1150
rect 25400 1090 25410 1130
rect 25450 1090 25460 1130
rect 25400 1030 25460 1090
rect 25400 990 25410 1030
rect 25450 990 25460 1030
rect 25400 970 25460 990
rect 25580 1130 25640 1150
rect 25580 1090 25590 1130
rect 25630 1090 25640 1130
rect 25580 1030 25640 1090
rect 25580 990 25590 1030
rect 25630 990 25640 1030
rect 25580 970 25640 990
rect 25760 1130 25820 1150
rect 25760 1090 25770 1130
rect 25810 1090 25820 1130
rect 25760 1030 25820 1090
rect 25760 990 25770 1030
rect 25810 990 25820 1030
rect 25760 970 25820 990
rect 25940 1130 26000 1150
rect 25940 1090 25950 1130
rect 25990 1090 26000 1130
rect 25940 1030 26000 1090
rect 25940 990 25950 1030
rect 25990 990 26000 1030
rect 25940 970 26000 990
rect 26120 1130 26180 1150
rect 26120 1090 26130 1130
rect 26170 1090 26180 1130
rect 26120 1030 26180 1090
rect 26120 990 26130 1030
rect 26170 990 26180 1030
rect 26120 970 26180 990
rect 26300 1130 26360 1150
rect 26300 1090 26310 1130
rect 26350 1090 26360 1130
rect 26300 1030 26360 1090
rect 26300 990 26310 1030
rect 26350 990 26360 1030
rect 26300 970 26360 990
rect 26480 1130 26540 1150
rect 26480 1090 26490 1130
rect 26530 1090 26540 1130
rect 26480 1030 26540 1090
rect 26480 990 26490 1030
rect 26530 990 26540 1030
rect 26480 970 26540 990
rect 26660 1130 26720 1150
rect 26660 1090 26670 1130
rect 26710 1090 26720 1130
rect 26660 1030 26720 1090
rect 26660 990 26670 1030
rect 26710 990 26720 1030
rect 26660 970 26720 990
rect 26840 1130 26900 1150
rect 26840 1090 26850 1130
rect 26890 1090 26900 1130
rect 26840 1030 26900 1090
rect 26840 990 26850 1030
rect 26890 990 26900 1030
rect 26840 970 26900 990
rect 26970 1140 27010 1310
rect 25590 930 25630 970
rect 25950 930 25990 970
rect 26310 930 26350 970
rect 26670 930 26710 970
rect 25570 910 25650 930
rect 25570 870 25590 910
rect 25630 870 25650 910
rect 25570 850 25650 870
rect 25930 910 26010 930
rect 25930 870 25950 910
rect 25990 870 26010 910
rect 25930 850 26010 870
rect 26290 910 26370 930
rect 26290 870 26310 910
rect 26350 870 26370 910
rect 26290 850 26370 870
rect 26650 910 26730 930
rect 26650 870 26670 910
rect 26710 870 26730 910
rect 26650 850 26730 870
rect 26970 810 27010 980
rect 25290 770 26070 810
rect 26230 770 27010 810
rect 27130 1310 28090 1350
rect 28250 1310 29210 1350
rect 27130 1140 27170 1310
rect 27590 1250 27670 1270
rect 27590 1210 27610 1250
rect 27650 1210 27670 1250
rect 27590 1190 27670 1210
rect 27950 1250 28030 1270
rect 27950 1210 27970 1250
rect 28010 1210 28030 1250
rect 27950 1190 28030 1210
rect 28310 1250 28390 1270
rect 28310 1210 28330 1250
rect 28370 1210 28390 1250
rect 28310 1190 28390 1210
rect 28670 1250 28750 1270
rect 28670 1210 28690 1250
rect 28730 1210 28750 1250
rect 28670 1190 28750 1210
rect 27610 1150 27650 1190
rect 27970 1150 28010 1190
rect 28330 1150 28370 1190
rect 28690 1150 28730 1190
rect 27130 810 27170 980
rect 27240 1130 27300 1150
rect 27240 1090 27250 1130
rect 27290 1090 27300 1130
rect 27240 1030 27300 1090
rect 27240 990 27250 1030
rect 27290 990 27300 1030
rect 27240 970 27300 990
rect 27420 1130 27480 1150
rect 27420 1090 27430 1130
rect 27470 1090 27480 1130
rect 27420 1030 27480 1090
rect 27420 990 27430 1030
rect 27470 990 27480 1030
rect 27420 970 27480 990
rect 27600 1130 27660 1150
rect 27600 1090 27610 1130
rect 27650 1090 27660 1130
rect 27600 1030 27660 1090
rect 27600 990 27610 1030
rect 27650 990 27660 1030
rect 27600 970 27660 990
rect 27780 1130 27840 1150
rect 27780 1090 27790 1130
rect 27830 1090 27840 1130
rect 27780 1030 27840 1090
rect 27780 990 27790 1030
rect 27830 990 27840 1030
rect 27780 970 27840 990
rect 27960 1130 28020 1150
rect 27960 1090 27970 1130
rect 28010 1090 28020 1130
rect 27960 1030 28020 1090
rect 27960 990 27970 1030
rect 28010 990 28020 1030
rect 27960 970 28020 990
rect 28140 1130 28200 1150
rect 28140 1090 28150 1130
rect 28190 1090 28200 1130
rect 28140 1030 28200 1090
rect 28140 990 28150 1030
rect 28190 990 28200 1030
rect 28140 970 28200 990
rect 28320 1130 28380 1150
rect 28320 1090 28330 1130
rect 28370 1090 28380 1130
rect 28320 1030 28380 1090
rect 28320 990 28330 1030
rect 28370 990 28380 1030
rect 28320 970 28380 990
rect 28500 1130 28560 1150
rect 28500 1090 28510 1130
rect 28550 1090 28560 1130
rect 28500 1030 28560 1090
rect 28500 990 28510 1030
rect 28550 990 28560 1030
rect 28500 970 28560 990
rect 28680 1130 28740 1150
rect 28680 1090 28690 1130
rect 28730 1090 28740 1130
rect 28680 1030 28740 1090
rect 28680 990 28690 1030
rect 28730 990 28740 1030
rect 28680 970 28740 990
rect 28860 1130 28920 1150
rect 28860 1090 28870 1130
rect 28910 1090 28920 1130
rect 28860 1030 28920 1090
rect 28860 990 28870 1030
rect 28910 990 28920 1030
rect 28860 970 28920 990
rect 29040 1130 29100 1150
rect 29040 1090 29050 1130
rect 29090 1090 29100 1130
rect 29040 1030 29100 1090
rect 29040 990 29050 1030
rect 29090 990 29100 1030
rect 29040 970 29100 990
rect 29170 1140 29210 1310
rect 27430 930 27470 970
rect 27790 930 27830 970
rect 28150 930 28190 970
rect 28510 930 28550 970
rect 28870 930 28910 970
rect 27410 910 27490 930
rect 27410 870 27430 910
rect 27470 870 27490 910
rect 27410 850 27490 870
rect 28130 910 28210 930
rect 28130 870 28150 910
rect 28190 870 28210 910
rect 28130 850 28210 870
rect 28490 910 28570 930
rect 28490 870 28510 910
rect 28550 870 28570 910
rect 28490 850 28570 870
rect 28850 910 28930 930
rect 28850 870 28870 910
rect 28910 870 28930 910
rect 28850 850 28930 870
rect 29170 810 29210 980
rect 27130 770 28090 810
rect 28250 770 29210 810
rect 29290 1310 30070 1350
rect 30230 1310 31010 1350
rect 29290 1140 29330 1310
rect 29750 1250 29830 1270
rect 29750 1210 29770 1250
rect 29810 1210 29830 1250
rect 29750 1190 29830 1210
rect 30110 1250 30190 1270
rect 30110 1210 30130 1250
rect 30170 1210 30190 1250
rect 30110 1190 30190 1210
rect 30470 1250 30550 1270
rect 30470 1210 30490 1250
rect 30530 1210 30550 1250
rect 30470 1190 30550 1210
rect 29770 1150 29810 1190
rect 30130 1150 30170 1190
rect 30490 1150 30530 1190
rect 29290 810 29330 980
rect 29400 1130 29460 1150
rect 29400 1090 29410 1130
rect 29450 1090 29460 1130
rect 29400 1030 29460 1090
rect 29400 990 29410 1030
rect 29450 990 29460 1030
rect 29400 970 29460 990
rect 29580 1130 29640 1150
rect 29580 1090 29590 1130
rect 29630 1090 29640 1130
rect 29580 1030 29640 1090
rect 29580 990 29590 1030
rect 29630 990 29640 1030
rect 29580 970 29640 990
rect 29760 1130 29820 1150
rect 29760 1090 29770 1130
rect 29810 1090 29820 1130
rect 29760 1030 29820 1090
rect 29760 990 29770 1030
rect 29810 990 29820 1030
rect 29760 970 29820 990
rect 29940 1130 30000 1150
rect 29940 1090 29950 1130
rect 29990 1090 30000 1130
rect 29940 1030 30000 1090
rect 29940 990 29950 1030
rect 29990 990 30000 1030
rect 29940 970 30000 990
rect 30120 1130 30180 1150
rect 30120 1090 30130 1130
rect 30170 1090 30180 1130
rect 30120 1030 30180 1090
rect 30120 990 30130 1030
rect 30170 990 30180 1030
rect 30120 970 30180 990
rect 30300 1130 30360 1150
rect 30300 1090 30310 1130
rect 30350 1090 30360 1130
rect 30300 1030 30360 1090
rect 30300 990 30310 1030
rect 30350 990 30360 1030
rect 30300 970 30360 990
rect 30480 1130 30540 1150
rect 30480 1090 30490 1130
rect 30530 1090 30540 1130
rect 30480 1030 30540 1090
rect 30480 990 30490 1030
rect 30530 990 30540 1030
rect 30480 970 30540 990
rect 30660 1130 30720 1150
rect 30660 1090 30670 1130
rect 30710 1090 30720 1130
rect 30660 1030 30720 1090
rect 30660 990 30670 1030
rect 30710 990 30720 1030
rect 30660 970 30720 990
rect 30840 1130 30900 1150
rect 30840 1090 30850 1130
rect 30890 1090 30900 1130
rect 30840 1030 30900 1090
rect 30840 990 30850 1030
rect 30890 990 30900 1030
rect 30840 970 30900 990
rect 30970 1140 31010 1310
rect 29590 930 29630 970
rect 29950 930 29990 970
rect 30310 930 30350 970
rect 30670 930 30710 970
rect 29570 910 29650 930
rect 29570 870 29590 910
rect 29630 870 29650 910
rect 29570 850 29650 870
rect 29930 910 30010 930
rect 29930 870 29950 910
rect 29990 870 30010 910
rect 29930 850 30010 870
rect 30290 910 30370 930
rect 30290 870 30310 910
rect 30350 870 30370 910
rect 30290 850 30370 870
rect 30650 910 30730 930
rect 30650 870 30670 910
rect 30710 870 30730 910
rect 30650 850 30730 870
rect 30970 810 31010 980
rect 29290 770 30070 810
rect 30230 770 31010 810
rect 25940 750 26000 770
rect 26660 750 26720 770
rect 29940 750 30000 770
rect 30660 750 30720 770
rect 25070 660 25130 720
<< viali >>
rect 20112 6350 20162 6400
rect 22542 6340 22592 6390
rect 20112 6230 20162 6280
rect 22542 6220 22592 6270
rect 20112 6070 20162 6120
rect 20112 5950 20162 6000
rect 21840 5760 21900 5820
rect 22000 5760 22060 5820
rect 22160 5760 22220 5820
rect 24680 5860 24730 5910
rect 26340 6300 26380 6340
rect 26710 6300 26750 6340
rect 27070 6300 27110 6340
rect 27430 6300 27470 6340
rect 27790 6300 27830 6340
rect 28150 6300 28190 6340
rect 28510 6300 28550 6340
rect 28870 6300 28910 6340
rect 29230 6300 29270 6340
rect 29590 6300 29630 6340
rect 29850 6300 29890 6340
rect 29950 6300 29990 6340
rect 26170 5960 26210 6000
rect 26530 5960 26570 6000
rect 26890 5960 26930 6000
rect 27250 5960 27290 6000
rect 27610 5960 27650 6000
rect 27970 5960 28010 6000
rect 28330 5960 28370 6000
rect 28690 5960 28730 6000
rect 29050 5960 29090 6000
rect 29410 5960 29450 6000
rect 29770 5960 29810 6000
rect 29900 5960 29940 6000
rect 30130 5960 30170 6000
rect 24680 5740 24730 5790
rect 20122 5630 20172 5680
rect 21468 5630 21518 5680
rect 22542 5620 22592 5670
rect 23940 5620 23990 5670
rect 20122 5510 20172 5560
rect 21468 5510 21518 5560
rect 20626 4604 20648 4610
rect 20648 4604 20660 4610
rect 20726 4604 20738 4610
rect 20738 4604 20760 4610
rect 20826 4604 20828 4610
rect 20828 4604 20860 4610
rect 20626 4576 20660 4604
rect 20726 4576 20760 4604
rect 20826 4576 20860 4604
rect 20926 4576 20960 4610
rect 21026 4576 21060 4610
rect 21126 4604 21154 4610
rect 21154 4604 21160 4610
rect 21126 4576 21160 4604
rect 20626 4476 20660 4510
rect 20726 4476 20760 4510
rect 20826 4476 20860 4510
rect 20926 4476 20960 4510
rect 21026 4476 21060 4510
rect 21126 4476 21160 4510
rect 20626 4376 20660 4410
rect 20726 4376 20760 4410
rect 20826 4376 20860 4410
rect 20926 4376 20960 4410
rect 21026 4376 21060 4410
rect 21126 4376 21160 4410
rect 20626 4278 20660 4310
rect 20726 4278 20760 4310
rect 20826 4278 20860 4310
rect 20626 4276 20648 4278
rect 20648 4276 20660 4278
rect 20726 4276 20738 4278
rect 20738 4276 20760 4278
rect 20826 4276 20828 4278
rect 20828 4276 20860 4278
rect 20926 4276 20960 4310
rect 21026 4276 21060 4310
rect 21126 4278 21160 4310
rect 21126 4276 21154 4278
rect 21154 4276 21160 4278
rect 20626 4188 20660 4210
rect 20726 4188 20760 4210
rect 20826 4188 20860 4210
rect 20626 4176 20648 4188
rect 20648 4176 20660 4188
rect 20726 4176 20738 4188
rect 20738 4176 20760 4188
rect 20826 4176 20828 4188
rect 20828 4176 20860 4188
rect 20926 4176 20960 4210
rect 21026 4176 21060 4210
rect 21126 4188 21160 4210
rect 21126 4176 21154 4188
rect 21154 4176 21160 4188
rect 20626 4098 20660 4110
rect 20726 4098 20760 4110
rect 20826 4098 20860 4110
rect 20626 4076 20648 4098
rect 20648 4076 20660 4098
rect 20726 4076 20738 4098
rect 20738 4076 20760 4098
rect 20826 4076 20828 4098
rect 20828 4076 20860 4098
rect 20926 4076 20960 4110
rect 21026 4076 21060 4110
rect 21126 4098 21160 4110
rect 21126 4076 21154 4098
rect 21154 4076 21160 4098
rect 21986 4604 22008 4610
rect 22008 4604 22020 4610
rect 22086 4604 22098 4610
rect 22098 4604 22120 4610
rect 22186 4604 22188 4610
rect 22188 4604 22220 4610
rect 21986 4576 22020 4604
rect 22086 4576 22120 4604
rect 22186 4576 22220 4604
rect 22286 4576 22320 4610
rect 22386 4576 22420 4610
rect 22486 4604 22514 4610
rect 22514 4604 22520 4610
rect 22486 4576 22520 4604
rect 21986 4476 22020 4510
rect 22086 4476 22120 4510
rect 22186 4476 22220 4510
rect 22286 4476 22320 4510
rect 22386 4476 22420 4510
rect 22486 4476 22520 4510
rect 21986 4376 22020 4410
rect 22086 4376 22120 4410
rect 22186 4376 22220 4410
rect 22286 4376 22320 4410
rect 22386 4376 22420 4410
rect 22486 4376 22520 4410
rect 21986 4278 22020 4310
rect 22086 4278 22120 4310
rect 22186 4278 22220 4310
rect 21986 4276 22008 4278
rect 22008 4276 22020 4278
rect 22086 4276 22098 4278
rect 22098 4276 22120 4278
rect 22186 4276 22188 4278
rect 22188 4276 22220 4278
rect 22286 4276 22320 4310
rect 22386 4276 22420 4310
rect 22486 4278 22520 4310
rect 22486 4276 22514 4278
rect 22514 4276 22520 4278
rect 21986 4188 22020 4210
rect 22086 4188 22120 4210
rect 22186 4188 22220 4210
rect 21986 4176 22008 4188
rect 22008 4176 22020 4188
rect 22086 4176 22098 4188
rect 22098 4176 22120 4188
rect 22186 4176 22188 4188
rect 22188 4176 22220 4188
rect 22286 4176 22320 4210
rect 22386 4176 22420 4210
rect 22486 4188 22520 4210
rect 22486 4176 22514 4188
rect 22514 4176 22520 4188
rect 21986 4098 22020 4110
rect 22086 4098 22120 4110
rect 22186 4098 22220 4110
rect 21986 4076 22008 4098
rect 22008 4076 22020 4098
rect 22086 4076 22098 4098
rect 22098 4076 22120 4098
rect 22186 4076 22188 4098
rect 22188 4076 22220 4098
rect 22286 4076 22320 4110
rect 22386 4076 22420 4110
rect 22486 4098 22520 4110
rect 22486 4076 22514 4098
rect 22514 4076 22520 4098
rect 25510 4810 25550 4850
rect 25640 4810 25680 4850
rect 25770 4810 25810 4850
rect 23346 4604 23368 4610
rect 23368 4604 23380 4610
rect 23446 4604 23458 4610
rect 23458 4604 23480 4610
rect 23546 4604 23548 4610
rect 23548 4604 23580 4610
rect 23346 4576 23380 4604
rect 23446 4576 23480 4604
rect 23546 4576 23580 4604
rect 23646 4576 23680 4610
rect 23746 4576 23780 4610
rect 23846 4604 23874 4610
rect 23874 4604 23880 4610
rect 23846 4576 23880 4604
rect 23346 4476 23380 4510
rect 23446 4476 23480 4510
rect 23546 4476 23580 4510
rect 23646 4476 23680 4510
rect 23746 4476 23780 4510
rect 23846 4476 23880 4510
rect 23346 4376 23380 4410
rect 23446 4376 23480 4410
rect 23546 4376 23580 4410
rect 23646 4376 23680 4410
rect 23746 4376 23780 4410
rect 23846 4376 23880 4410
rect 23346 4278 23380 4310
rect 23446 4278 23480 4310
rect 23546 4278 23580 4310
rect 23346 4276 23368 4278
rect 23368 4276 23380 4278
rect 23446 4276 23458 4278
rect 23458 4276 23480 4278
rect 23546 4276 23548 4278
rect 23548 4276 23580 4278
rect 23646 4276 23680 4310
rect 23746 4276 23780 4310
rect 23846 4278 23880 4310
rect 23846 4276 23874 4278
rect 23874 4276 23880 4278
rect 23346 4188 23380 4210
rect 23446 4188 23480 4210
rect 23546 4188 23580 4210
rect 23346 4176 23368 4188
rect 23368 4176 23380 4188
rect 23446 4176 23458 4188
rect 23458 4176 23480 4188
rect 23546 4176 23548 4188
rect 23548 4176 23580 4188
rect 23646 4176 23680 4210
rect 23746 4176 23780 4210
rect 23846 4188 23880 4210
rect 23846 4176 23874 4188
rect 23874 4176 23880 4188
rect 23346 4098 23380 4110
rect 23446 4098 23480 4110
rect 23546 4098 23580 4110
rect 23346 4076 23368 4098
rect 23368 4076 23380 4098
rect 23446 4076 23458 4098
rect 23458 4076 23480 4098
rect 23546 4076 23548 4098
rect 23548 4076 23580 4098
rect 23646 4076 23680 4110
rect 23746 4076 23780 4110
rect 23846 4098 23880 4110
rect 23846 4076 23874 4098
rect 23874 4076 23880 4098
rect 26890 5380 26930 5420
rect 27250 5380 27290 5420
rect 27610 5380 27650 5420
rect 27970 5380 28010 5420
rect 28330 5380 28370 5420
rect 28690 5380 28730 5420
rect 29050 5380 29090 5420
rect 29410 5380 29450 5420
rect 26710 4640 26750 4680
rect 27070 4640 27110 4680
rect 27430 4640 27470 4680
rect 27670 4640 27710 4680
rect 27790 4640 27830 4680
rect 28150 4640 28190 4680
rect 28510 4640 28550 4680
rect 28870 4640 28910 4680
rect 29230 4640 29270 4680
rect 29410 4640 29450 4680
rect 29590 4640 29630 4680
rect 19930 2990 19970 3030
rect 20626 3244 20648 3250
rect 20648 3244 20660 3250
rect 20726 3244 20738 3250
rect 20738 3244 20760 3250
rect 20826 3244 20828 3250
rect 20828 3244 20860 3250
rect 20626 3216 20660 3244
rect 20726 3216 20760 3244
rect 20826 3216 20860 3244
rect 20926 3216 20960 3250
rect 21026 3216 21060 3250
rect 21126 3244 21154 3250
rect 21154 3244 21160 3250
rect 21126 3216 21160 3244
rect 20626 3116 20660 3150
rect 20726 3116 20760 3150
rect 20826 3116 20860 3150
rect 20926 3116 20960 3150
rect 21026 3116 21060 3150
rect 21126 3116 21160 3150
rect 20626 3016 20660 3050
rect 20726 3016 20760 3050
rect 20826 3016 20860 3050
rect 20926 3016 20960 3050
rect 21026 3016 21060 3050
rect 21126 3016 21160 3050
rect 20626 2918 20660 2950
rect 20726 2918 20760 2950
rect 20826 2918 20860 2950
rect 20626 2916 20648 2918
rect 20648 2916 20660 2918
rect 20726 2916 20738 2918
rect 20738 2916 20760 2918
rect 20826 2916 20828 2918
rect 20828 2916 20860 2918
rect 20926 2916 20960 2950
rect 21026 2916 21060 2950
rect 21126 2918 21160 2950
rect 21126 2916 21154 2918
rect 21154 2916 21160 2918
rect 20626 2828 20660 2850
rect 20726 2828 20760 2850
rect 20826 2828 20860 2850
rect 20626 2816 20648 2828
rect 20648 2816 20660 2828
rect 20726 2816 20738 2828
rect 20738 2816 20760 2828
rect 20826 2816 20828 2828
rect 20828 2816 20860 2828
rect 20926 2816 20960 2850
rect 21026 2816 21060 2850
rect 21126 2828 21160 2850
rect 21126 2816 21154 2828
rect 21154 2816 21160 2828
rect 20626 2738 20660 2750
rect 20726 2738 20760 2750
rect 20826 2738 20860 2750
rect 20626 2716 20648 2738
rect 20648 2716 20660 2738
rect 20726 2716 20738 2738
rect 20738 2716 20760 2738
rect 20826 2716 20828 2738
rect 20828 2716 20860 2738
rect 20926 2716 20960 2750
rect 21026 2716 21060 2750
rect 21126 2738 21160 2750
rect 21126 2716 21154 2738
rect 21154 2716 21160 2738
rect 21986 3244 22008 3250
rect 22008 3244 22020 3250
rect 22086 3244 22098 3250
rect 22098 3244 22120 3250
rect 22186 3244 22188 3250
rect 22188 3244 22220 3250
rect 21986 3216 22020 3244
rect 22086 3216 22120 3244
rect 22186 3216 22220 3244
rect 22286 3216 22320 3250
rect 22386 3216 22420 3250
rect 22486 3244 22514 3250
rect 22514 3244 22520 3250
rect 22486 3216 22520 3244
rect 21986 3116 22020 3150
rect 22086 3116 22120 3150
rect 22186 3116 22220 3150
rect 22286 3116 22320 3150
rect 22386 3116 22420 3150
rect 22486 3116 22520 3150
rect 21986 3016 22020 3050
rect 22086 3016 22120 3050
rect 22186 3016 22220 3050
rect 22286 3016 22320 3050
rect 22386 3016 22420 3050
rect 22486 3016 22520 3050
rect 21986 2918 22020 2950
rect 22086 2918 22120 2950
rect 22186 2918 22220 2950
rect 21986 2916 22008 2918
rect 22008 2916 22020 2918
rect 22086 2916 22098 2918
rect 22098 2916 22120 2918
rect 22186 2916 22188 2918
rect 22188 2916 22220 2918
rect 22286 2916 22320 2950
rect 22386 2916 22420 2950
rect 22486 2918 22520 2950
rect 22486 2916 22514 2918
rect 22514 2916 22520 2918
rect 21986 2828 22020 2850
rect 22086 2828 22120 2850
rect 22186 2828 22220 2850
rect 21986 2816 22008 2828
rect 22008 2816 22020 2828
rect 22086 2816 22098 2828
rect 22098 2816 22120 2828
rect 22186 2816 22188 2828
rect 22188 2816 22220 2828
rect 22286 2816 22320 2850
rect 22386 2816 22420 2850
rect 22486 2828 22520 2850
rect 22486 2816 22514 2828
rect 22514 2816 22520 2828
rect 21986 2738 22020 2750
rect 22086 2738 22120 2750
rect 22186 2738 22220 2750
rect 21986 2716 22008 2738
rect 22008 2716 22020 2738
rect 22086 2716 22098 2738
rect 22098 2716 22120 2738
rect 22186 2716 22188 2738
rect 22188 2716 22220 2738
rect 22286 2716 22320 2750
rect 22386 2716 22420 2750
rect 22486 2738 22520 2750
rect 22486 2716 22514 2738
rect 22514 2716 22520 2738
rect 25430 4050 25470 4090
rect 25550 4050 25590 4090
rect 25670 4050 25710 4090
rect 25910 4050 25950 4090
rect 26150 4050 26190 4090
rect 26270 4050 26310 4090
rect 26390 4050 26430 4090
rect 26630 4050 26670 4090
rect 26870 4050 26910 4090
rect 26990 4050 27030 4090
rect 27110 4050 27150 4090
rect 27350 4050 27390 4090
rect 27590 4050 27630 4090
rect 27710 4050 27750 4090
rect 25610 3710 25650 3750
rect 25790 3710 25830 3750
rect 26030 3710 26070 3750
rect 26270 3710 26310 3750
rect 26510 3710 26550 3750
rect 26750 3710 26790 3750
rect 26990 3710 27030 3750
rect 27230 3710 27270 3750
rect 27470 3710 27510 3750
rect 27650 3710 27690 3750
rect 28710 4170 28750 4210
rect 28950 4170 28990 4210
rect 29190 4170 29230 4210
rect 29430 4170 29470 4210
rect 29670 4190 29710 4210
rect 29670 4170 29710 4190
rect 29910 4170 29950 4210
rect 30150 4170 30190 4210
rect 30390 4170 30430 4210
rect 30630 4170 30670 4210
rect 30870 4170 30910 4210
rect 28590 4050 28630 4090
rect 28710 4050 28750 4090
rect 28950 4050 28990 4090
rect 29190 4050 29230 4090
rect 29310 4050 29350 4090
rect 29430 4050 29470 4090
rect 29670 4050 29710 4090
rect 29910 4050 29950 4090
rect 30030 4050 30070 4090
rect 30150 4050 30190 4090
rect 30390 4050 30430 4090
rect 30630 4050 30670 4090
rect 30750 4050 30790 4090
rect 30870 4050 30910 4090
rect 28650 3710 28690 3750
rect 28830 3710 28870 3750
rect 29070 3710 29110 3750
rect 29310 3710 29350 3750
rect 29550 3710 29590 3750
rect 29790 3710 29830 3750
rect 30030 3710 30070 3750
rect 30270 3710 30310 3750
rect 30510 3710 30550 3750
rect 30690 3710 30730 3750
rect 23346 3244 23368 3250
rect 23368 3244 23380 3250
rect 23446 3244 23458 3250
rect 23458 3244 23480 3250
rect 23546 3244 23548 3250
rect 23548 3244 23580 3250
rect 23346 3216 23380 3244
rect 23446 3216 23480 3244
rect 23546 3216 23580 3244
rect 23646 3216 23680 3250
rect 23746 3216 23780 3250
rect 23846 3244 23874 3250
rect 23874 3244 23880 3250
rect 23846 3216 23880 3244
rect 23346 3116 23380 3150
rect 23446 3116 23480 3150
rect 23546 3116 23580 3150
rect 23646 3116 23680 3150
rect 23746 3116 23780 3150
rect 23846 3116 23880 3150
rect 23346 3016 23380 3050
rect 23446 3016 23480 3050
rect 23546 3016 23580 3050
rect 23646 3016 23680 3050
rect 23746 3016 23780 3050
rect 23846 3016 23880 3050
rect 23346 2918 23380 2950
rect 23446 2918 23480 2950
rect 23546 2918 23580 2950
rect 23346 2916 23368 2918
rect 23368 2916 23380 2918
rect 23446 2916 23458 2918
rect 23458 2916 23480 2918
rect 23546 2916 23548 2918
rect 23548 2916 23580 2918
rect 23646 2916 23680 2950
rect 23746 2916 23780 2950
rect 23846 2918 23880 2950
rect 23846 2916 23874 2918
rect 23874 2916 23880 2918
rect 23346 2828 23380 2850
rect 23446 2828 23480 2850
rect 23546 2828 23580 2850
rect 23346 2816 23368 2828
rect 23368 2816 23380 2828
rect 23446 2816 23458 2828
rect 23458 2816 23480 2828
rect 23546 2816 23548 2828
rect 23548 2816 23580 2828
rect 23646 2816 23680 2850
rect 23746 2816 23780 2850
rect 23846 2828 23880 2850
rect 23846 2816 23874 2828
rect 23874 2816 23880 2828
rect 23346 2738 23380 2750
rect 23446 2738 23480 2750
rect 23546 2738 23580 2750
rect 23346 2716 23368 2738
rect 23368 2716 23380 2738
rect 23446 2716 23458 2738
rect 23458 2716 23480 2738
rect 23546 2716 23548 2738
rect 23548 2716 23580 2738
rect 23646 2716 23680 2750
rect 23746 2716 23780 2750
rect 23846 2738 23880 2750
rect 23846 2716 23874 2738
rect 23874 2716 23880 2738
rect 26410 3390 26450 3430
rect 26290 3300 26330 3340
rect 26530 3300 26570 3340
rect 26770 3300 26810 3340
rect 27010 3300 27050 3340
rect 27250 3300 27290 3340
rect 27490 3300 27530 3340
rect 26290 3060 26330 3100
rect 26410 3060 26450 3100
rect 26650 3060 26690 3100
rect 26890 3060 26930 3100
rect 27130 3060 27170 3100
rect 27370 3060 27410 3100
rect 27370 2940 27410 2980
rect 29890 3390 29930 3430
rect 28810 3300 28850 3340
rect 29050 3300 29090 3340
rect 29290 3300 29330 3340
rect 29530 3300 29570 3340
rect 29770 3300 29810 3340
rect 30010 3300 30050 3340
rect 28930 3060 28970 3100
rect 29170 3060 29210 3100
rect 29410 3060 29450 3100
rect 29650 3060 29690 3100
rect 29890 3060 29930 3100
rect 30010 3060 30050 3100
rect 20626 1884 20648 1890
rect 20648 1884 20660 1890
rect 20726 1884 20738 1890
rect 20738 1884 20760 1890
rect 20826 1884 20828 1890
rect 20828 1884 20860 1890
rect 20626 1856 20660 1884
rect 20726 1856 20760 1884
rect 20826 1856 20860 1884
rect 20926 1856 20960 1890
rect 21026 1856 21060 1890
rect 21126 1884 21154 1890
rect 21154 1884 21160 1890
rect 21126 1856 21160 1884
rect 20626 1756 20660 1790
rect 20726 1756 20760 1790
rect 20826 1756 20860 1790
rect 20926 1756 20960 1790
rect 21026 1756 21060 1790
rect 21126 1756 21160 1790
rect 20626 1656 20660 1690
rect 20726 1656 20760 1690
rect 20826 1656 20860 1690
rect 20926 1656 20960 1690
rect 21026 1656 21060 1690
rect 21126 1656 21160 1690
rect 20626 1558 20660 1590
rect 20726 1558 20760 1590
rect 20826 1558 20860 1590
rect 20626 1556 20648 1558
rect 20648 1556 20660 1558
rect 20726 1556 20738 1558
rect 20738 1556 20760 1558
rect 20826 1556 20828 1558
rect 20828 1556 20860 1558
rect 20926 1556 20960 1590
rect 21026 1556 21060 1590
rect 21126 1558 21160 1590
rect 21126 1556 21154 1558
rect 21154 1556 21160 1558
rect 20626 1468 20660 1490
rect 20726 1468 20760 1490
rect 20826 1468 20860 1490
rect 20626 1456 20648 1468
rect 20648 1456 20660 1468
rect 20726 1456 20738 1468
rect 20738 1456 20760 1468
rect 20826 1456 20828 1468
rect 20828 1456 20860 1468
rect 20926 1456 20960 1490
rect 21026 1456 21060 1490
rect 21126 1468 21160 1490
rect 21126 1456 21154 1468
rect 21154 1456 21160 1468
rect 20626 1378 20660 1390
rect 20726 1378 20760 1390
rect 20826 1378 20860 1390
rect 20626 1356 20648 1378
rect 20648 1356 20660 1378
rect 20726 1356 20738 1378
rect 20738 1356 20760 1378
rect 20826 1356 20828 1378
rect 20828 1356 20860 1378
rect 20926 1356 20960 1390
rect 21026 1356 21060 1390
rect 21126 1378 21160 1390
rect 21126 1356 21154 1378
rect 21154 1356 21160 1378
rect 21986 1884 22008 1890
rect 22008 1884 22020 1890
rect 22086 1884 22098 1890
rect 22098 1884 22120 1890
rect 22186 1884 22188 1890
rect 22188 1884 22220 1890
rect 21986 1856 22020 1884
rect 22086 1856 22120 1884
rect 22186 1856 22220 1884
rect 22286 1856 22320 1890
rect 22386 1856 22420 1890
rect 22486 1884 22514 1890
rect 22514 1884 22520 1890
rect 22486 1856 22520 1884
rect 21986 1756 22020 1790
rect 22086 1756 22120 1790
rect 22186 1756 22220 1790
rect 22286 1756 22320 1790
rect 22386 1756 22420 1790
rect 22486 1756 22520 1790
rect 21986 1656 22020 1690
rect 22086 1656 22120 1690
rect 22186 1656 22220 1690
rect 22286 1656 22320 1690
rect 22386 1656 22420 1690
rect 22486 1656 22520 1690
rect 21986 1558 22020 1590
rect 22086 1558 22120 1590
rect 22186 1558 22220 1590
rect 21986 1556 22008 1558
rect 22008 1556 22020 1558
rect 22086 1556 22098 1558
rect 22098 1556 22120 1558
rect 22186 1556 22188 1558
rect 22188 1556 22220 1558
rect 22286 1556 22320 1590
rect 22386 1556 22420 1590
rect 22486 1558 22520 1590
rect 22486 1556 22514 1558
rect 22514 1556 22520 1558
rect 21986 1468 22020 1490
rect 22086 1468 22120 1490
rect 22186 1468 22220 1490
rect 21986 1456 22008 1468
rect 22008 1456 22020 1468
rect 22086 1456 22098 1468
rect 22098 1456 22120 1468
rect 22186 1456 22188 1468
rect 22188 1456 22220 1468
rect 22286 1456 22320 1490
rect 22386 1456 22420 1490
rect 22486 1468 22520 1490
rect 22486 1456 22514 1468
rect 22514 1456 22520 1468
rect 21986 1378 22020 1390
rect 22086 1378 22120 1390
rect 22186 1378 22220 1390
rect 21986 1356 22008 1378
rect 22008 1356 22020 1378
rect 22086 1356 22098 1378
rect 22098 1356 22120 1378
rect 22186 1356 22188 1378
rect 22188 1356 22220 1378
rect 22286 1356 22320 1390
rect 22386 1356 22420 1390
rect 22486 1378 22520 1390
rect 22486 1356 22514 1378
rect 22514 1356 22520 1378
rect 25810 2710 25850 2750
rect 25990 2740 26030 2780
rect 26230 2740 26270 2780
rect 26470 2740 26510 2780
rect 26710 2740 26750 2780
rect 27190 2740 27230 2780
rect 27430 2740 27470 2780
rect 27670 2740 27710 2780
rect 27970 2710 28010 2750
rect 26890 2110 26930 2150
rect 28330 2710 28370 2750
rect 28630 2740 28670 2780
rect 28870 2740 28910 2780
rect 29110 2740 29150 2780
rect 29590 2740 29630 2780
rect 29830 2740 29870 2780
rect 30070 2740 30110 2780
rect 30310 2740 30350 2780
rect 30490 2710 30530 2750
rect 29410 2110 29450 2150
rect 23346 1884 23368 1890
rect 23368 1884 23380 1890
rect 23446 1884 23458 1890
rect 23458 1884 23480 1890
rect 23546 1884 23548 1890
rect 23548 1884 23580 1890
rect 23346 1856 23380 1884
rect 23446 1856 23480 1884
rect 23546 1856 23580 1884
rect 23646 1856 23680 1890
rect 23746 1856 23780 1890
rect 23846 1884 23874 1890
rect 23874 1884 23880 1890
rect 23846 1856 23880 1884
rect 23346 1756 23380 1790
rect 23446 1756 23480 1790
rect 23546 1756 23580 1790
rect 23646 1756 23680 1790
rect 23746 1756 23780 1790
rect 23846 1756 23880 1790
rect 23346 1656 23380 1690
rect 23446 1656 23480 1690
rect 23546 1656 23580 1690
rect 23646 1656 23680 1690
rect 23746 1656 23780 1690
rect 23846 1656 23880 1690
rect 23346 1558 23380 1590
rect 23446 1558 23480 1590
rect 23546 1558 23580 1590
rect 23346 1556 23368 1558
rect 23368 1556 23380 1558
rect 23446 1556 23458 1558
rect 23458 1556 23480 1558
rect 23546 1556 23548 1558
rect 23548 1556 23580 1558
rect 23646 1556 23680 1590
rect 23746 1556 23780 1590
rect 23846 1558 23880 1590
rect 23846 1556 23874 1558
rect 23874 1556 23880 1558
rect 23346 1468 23380 1490
rect 23446 1468 23480 1490
rect 23546 1468 23580 1490
rect 23346 1456 23368 1468
rect 23368 1456 23380 1468
rect 23446 1456 23458 1468
rect 23458 1456 23480 1468
rect 23546 1456 23548 1468
rect 23548 1456 23580 1468
rect 23646 1456 23680 1490
rect 23746 1456 23780 1490
rect 23846 1468 23880 1490
rect 23846 1456 23874 1468
rect 23874 1456 23880 1468
rect 23346 1378 23380 1390
rect 23446 1378 23480 1390
rect 23546 1378 23580 1390
rect 23346 1356 23368 1378
rect 23368 1356 23380 1378
rect 23446 1356 23458 1378
rect 23458 1356 23480 1378
rect 23546 1356 23548 1378
rect 23548 1356 23580 1378
rect 23646 1356 23680 1390
rect 23746 1356 23780 1390
rect 23846 1378 23880 1390
rect 23846 1356 23874 1378
rect 23874 1356 23880 1378
rect 26070 1760 26110 1800
rect 26230 1760 26270 1800
rect 26390 1760 26430 1800
rect 26550 1760 26590 1800
rect 26710 1760 26750 1800
rect 26870 1760 26910 1800
rect 27030 1760 27070 1800
rect 27190 1760 27230 1800
rect 27350 1760 27390 1800
rect 27510 1760 27550 1800
rect 27670 1760 27710 1800
rect 27830 1760 27870 1800
rect 27990 1760 28030 1800
rect 28150 1760 28190 1800
rect 28310 1760 28350 1800
rect 28470 1760 28510 1800
rect 28630 1760 28670 1800
rect 28790 1760 28830 1800
rect 28950 1760 28990 1800
rect 29110 1760 29150 1800
rect 29270 1760 29310 1800
rect 29430 1760 29470 1800
rect 29590 1760 29630 1800
rect 29750 1760 29790 1800
rect 29910 1760 29950 1800
rect 30070 1760 30110 1800
rect 25990 1590 26030 1630
rect 30390 1590 30430 1630
rect 25770 1210 25810 1250
rect 26130 1210 26170 1250
rect 26490 1210 26530 1250
rect 25590 870 25630 910
rect 25950 870 25990 910
rect 26310 870 26350 910
rect 26670 870 26710 910
rect 27610 1210 27650 1250
rect 27970 1210 28010 1250
rect 28330 1210 28370 1250
rect 28690 1210 28730 1250
rect 27430 870 27470 910
rect 28150 870 28190 910
rect 28510 870 28550 910
rect 28870 870 28910 910
rect 29770 1210 29810 1250
rect 30130 1210 30170 1250
rect 30490 1210 30530 1250
rect 29590 870 29630 910
rect 29950 870 29990 910
rect 30310 870 30350 910
rect 30670 870 30710 910
<< metal1 >>
rect 22522 7050 22602 7060
rect 22522 6990 22532 7050
rect 22592 6990 22602 7050
rect 22522 6980 22602 6990
rect 28880 6990 28960 7000
rect 19970 6890 20050 6900
rect 19970 6830 19980 6890
rect 20040 6830 20050 6890
rect 19970 6820 20050 6830
rect 21880 6890 21960 6900
rect 21880 6830 21890 6890
rect 21950 6830 21960 6890
rect 21880 6820 21960 6830
rect 19880 6780 19960 6790
rect 19880 6720 19890 6780
rect 19950 6720 19960 6780
rect 19880 6710 19960 6720
rect 19900 5700 19940 6710
rect 19880 5690 19960 5700
rect 19880 5630 19890 5690
rect 19950 5630 19960 5690
rect 19880 5620 19960 5630
rect 19990 5580 20030 6820
rect 22410 6680 22490 6690
rect 22410 6620 22420 6680
rect 22480 6620 22490 6680
rect 22410 6610 22490 6620
rect 22320 6570 22400 6580
rect 22320 6510 22330 6570
rect 22390 6510 22400 6570
rect 22320 6500 22400 6510
rect 20092 6340 20102 6410
rect 20172 6340 20182 6410
rect 20092 6220 20102 6290
rect 20172 6220 20182 6290
rect 22340 6210 22380 6500
rect 22320 6200 22400 6210
rect 22320 6140 22330 6200
rect 22390 6140 22400 6200
rect 22320 6130 22400 6140
rect 20092 6060 20102 6130
rect 20172 6060 20182 6130
rect 20092 5940 20102 6010
rect 20172 5940 20182 6010
rect 21810 5820 22250 5840
rect 21810 5760 21840 5820
rect 21900 5760 22000 5820
rect 22060 5760 22160 5820
rect 22220 5760 22250 5820
rect 21810 5740 22250 5760
rect 22430 5690 22470 6610
rect 22542 6400 22582 6980
rect 28880 6930 28890 6990
rect 28950 6930 28960 6990
rect 28880 6920 28960 6930
rect 23270 6890 23370 6910
rect 23270 6830 23290 6890
rect 23350 6830 23370 6890
rect 24840 6900 24920 6910
rect 24840 6840 24850 6900
rect 24910 6840 24920 6900
rect 24840 6830 24920 6840
rect 30270 6890 30370 6910
rect 30270 6830 30290 6890
rect 30350 6830 30370 6890
rect 23270 6810 23370 6830
rect 22522 6330 22532 6400
rect 22602 6330 22612 6400
rect 22542 6280 22582 6330
rect 22522 6210 22532 6280
rect 22602 6210 22612 6280
rect 24660 5850 24670 5920
rect 24740 5850 24750 5920
rect 24660 5800 24750 5810
rect 24660 5730 24670 5800
rect 24740 5730 24750 5800
rect 24660 5720 24750 5730
rect 20102 5620 20112 5690
rect 20182 5620 20192 5690
rect 21448 5620 21458 5690
rect 21528 5620 21538 5690
rect 22410 5680 22490 5690
rect 24680 5680 24720 5720
rect 22410 5620 22420 5680
rect 22480 5620 22490 5680
rect 22410 5610 22490 5620
rect 22522 5610 22532 5680
rect 22602 5610 22612 5680
rect 23920 5610 23930 5680
rect 24000 5610 24010 5680
rect 24660 5670 24740 5680
rect 24660 5610 24670 5670
rect 24730 5610 24740 5670
rect 19970 5570 20050 5580
rect 19970 5510 19980 5570
rect 20040 5510 20050 5570
rect 19970 5500 20050 5510
rect 20102 5500 20112 5570
rect 20182 5500 20192 5570
rect 21448 5500 21458 5570
rect 21528 5500 21538 5570
rect 22542 5100 22582 5610
rect 24660 5600 24740 5610
rect 22522 5090 22602 5100
rect 22522 5030 22532 5090
rect 22592 5030 22602 5090
rect 22522 5020 22602 5030
rect 24300 5090 24380 5100
rect 24300 5030 24310 5090
rect 24370 5030 24380 5090
rect 24300 5020 24380 5030
rect 20550 4610 23970 4700
rect 20550 4576 20626 4610
rect 20660 4576 20726 4610
rect 20760 4576 20826 4610
rect 20860 4576 20926 4610
rect 20960 4576 21026 4610
rect 21060 4576 21126 4610
rect 21160 4576 21986 4610
rect 22020 4576 22086 4610
rect 22120 4576 22186 4610
rect 22220 4576 22286 4610
rect 22320 4576 22386 4610
rect 22420 4576 22486 4610
rect 22520 4576 23346 4610
rect 23380 4576 23446 4610
rect 23480 4576 23546 4610
rect 23580 4576 23646 4610
rect 23680 4576 23746 4610
rect 23780 4576 23846 4610
rect 23880 4576 23970 4610
rect 20550 4510 23970 4576
rect 20550 4476 20626 4510
rect 20660 4476 20726 4510
rect 20760 4476 20826 4510
rect 20860 4476 20926 4510
rect 20960 4476 21026 4510
rect 21060 4476 21126 4510
rect 21160 4476 21986 4510
rect 22020 4476 22086 4510
rect 22120 4476 22186 4510
rect 22220 4476 22286 4510
rect 22320 4476 22386 4510
rect 22420 4476 22486 4510
rect 22520 4476 23346 4510
rect 23380 4476 23446 4510
rect 23480 4476 23546 4510
rect 23580 4476 23646 4510
rect 23680 4476 23746 4510
rect 23780 4476 23846 4510
rect 23880 4476 23970 4510
rect 20550 4410 23970 4476
rect 20550 4376 20626 4410
rect 20660 4376 20726 4410
rect 20760 4376 20826 4410
rect 20860 4376 20926 4410
rect 20960 4376 21026 4410
rect 21060 4376 21126 4410
rect 21160 4376 21986 4410
rect 22020 4376 22086 4410
rect 22120 4376 22186 4410
rect 22220 4376 22286 4410
rect 22320 4376 22386 4410
rect 22420 4376 22486 4410
rect 22520 4376 23346 4410
rect 23380 4376 23446 4410
rect 23480 4376 23546 4410
rect 23580 4376 23646 4410
rect 23680 4376 23746 4410
rect 23780 4376 23846 4410
rect 23880 4376 23970 4410
rect 20550 4310 23970 4376
rect 20550 4276 20626 4310
rect 20660 4276 20726 4310
rect 20760 4276 20826 4310
rect 20860 4276 20926 4310
rect 20960 4276 21026 4310
rect 21060 4276 21126 4310
rect 21160 4276 21986 4310
rect 22020 4276 22086 4310
rect 22120 4276 22186 4310
rect 22220 4276 22286 4310
rect 22320 4276 22386 4310
rect 22420 4276 22486 4310
rect 22520 4276 23346 4310
rect 23380 4276 23446 4310
rect 23480 4276 23546 4310
rect 23580 4276 23646 4310
rect 23680 4276 23746 4310
rect 23780 4276 23846 4310
rect 23880 4276 23970 4310
rect 20550 4210 23970 4276
rect 20550 4176 20626 4210
rect 20660 4176 20726 4210
rect 20760 4176 20826 4210
rect 20860 4176 20926 4210
rect 20960 4176 21026 4210
rect 21060 4176 21126 4210
rect 21160 4176 21986 4210
rect 22020 4176 22086 4210
rect 22120 4176 22186 4210
rect 22220 4176 22286 4210
rect 22320 4176 22386 4210
rect 22420 4176 22486 4210
rect 22520 4176 23346 4210
rect 23380 4176 23446 4210
rect 23480 4176 23546 4210
rect 23580 4176 23646 4210
rect 23680 4176 23746 4210
rect 23780 4176 23846 4210
rect 23880 4176 23970 4210
rect 20550 4110 23970 4176
rect 20550 4076 20626 4110
rect 20660 4076 20726 4110
rect 20760 4076 20826 4110
rect 20860 4076 20926 4110
rect 20960 4076 21026 4110
rect 21060 4076 21126 4110
rect 21160 4076 21986 4110
rect 22020 4076 22086 4110
rect 22120 4076 22186 4110
rect 22220 4076 22286 4110
rect 22320 4076 22386 4110
rect 22420 4076 22486 4110
rect 22520 4076 23346 4110
rect 23380 4076 23446 4110
rect 23480 4076 23546 4110
rect 23580 4076 23646 4110
rect 23680 4076 23746 4110
rect 23780 4076 23846 4110
rect 23880 4076 23970 4110
rect 20550 4000 23970 4076
rect 20550 3250 21250 4000
rect 20550 3216 20626 3250
rect 20660 3216 20726 3250
rect 20760 3216 20826 3250
rect 20860 3216 20926 3250
rect 20960 3216 21026 3250
rect 21060 3216 21126 3250
rect 21160 3216 21250 3250
rect 20550 3150 21250 3216
rect 20550 3116 20626 3150
rect 20660 3116 20726 3150
rect 20760 3116 20826 3150
rect 20860 3116 20926 3150
rect 20960 3116 21026 3150
rect 21060 3116 21126 3150
rect 21160 3116 21250 3150
rect 20550 3050 21250 3116
rect 19780 3040 19860 3050
rect 19780 2980 19790 3040
rect 19850 3030 19860 3040
rect 19910 3040 19990 3050
rect 19910 3030 19920 3040
rect 19850 2990 19920 3030
rect 19850 2980 19860 2990
rect 19780 2970 19860 2980
rect 19910 2980 19920 2990
rect 19980 2980 19990 3040
rect 19910 2970 19990 2980
rect 20550 3016 20626 3050
rect 20660 3016 20726 3050
rect 20760 3016 20826 3050
rect 20860 3016 20926 3050
rect 20960 3016 21026 3050
rect 21060 3016 21126 3050
rect 21160 3016 21250 3050
rect 20550 2950 21250 3016
rect 20550 2916 20626 2950
rect 20660 2916 20726 2950
rect 20760 2916 20826 2950
rect 20860 2916 20926 2950
rect 20960 2916 21026 2950
rect 21060 2916 21126 2950
rect 21160 2916 21250 2950
rect 20550 2850 21250 2916
rect 20550 2816 20626 2850
rect 20660 2816 20726 2850
rect 20760 2816 20826 2850
rect 20860 2816 20926 2850
rect 20960 2816 21026 2850
rect 21060 2816 21126 2850
rect 21160 2816 21250 2850
rect 20550 2750 21250 2816
rect 20550 2716 20626 2750
rect 20660 2716 20726 2750
rect 20760 2716 20826 2750
rect 20860 2716 20926 2750
rect 20960 2716 21026 2750
rect 21060 2716 21126 2750
rect 21160 2716 21250 2750
rect 20550 1980 21250 2716
rect 21904 3250 22604 3340
rect 21904 3216 21986 3250
rect 22020 3216 22086 3250
rect 22120 3216 22186 3250
rect 22220 3216 22286 3250
rect 22320 3216 22386 3250
rect 22420 3216 22486 3250
rect 22520 3216 22604 3250
rect 21904 3150 22604 3216
rect 21904 3116 21986 3150
rect 22020 3116 22086 3150
rect 22120 3116 22186 3150
rect 22220 3116 22286 3150
rect 22320 3116 22386 3150
rect 22420 3116 22486 3150
rect 22520 3116 22604 3150
rect 21904 3050 22604 3116
rect 21904 3016 21986 3050
rect 22020 3016 22086 3050
rect 22120 3016 22186 3050
rect 22220 3016 22286 3050
rect 22320 3016 22386 3050
rect 22420 3016 22486 3050
rect 22520 3020 22604 3050
rect 22520 3016 22540 3020
rect 21904 2960 22540 3016
rect 22594 2960 22604 3020
rect 21904 2950 22604 2960
rect 21904 2916 21986 2950
rect 22020 2916 22086 2950
rect 22120 2916 22186 2950
rect 22220 2916 22286 2950
rect 22320 2916 22386 2950
rect 22420 2916 22486 2950
rect 22520 2916 22604 2950
rect 21904 2850 22604 2916
rect 21904 2816 21986 2850
rect 22020 2816 22086 2850
rect 22120 2816 22186 2850
rect 22220 2816 22286 2850
rect 22320 2816 22386 2850
rect 22420 2816 22486 2850
rect 22520 2816 22604 2850
rect 21904 2750 22604 2816
rect 21904 2716 21986 2750
rect 22020 2716 22086 2750
rect 22120 2716 22186 2750
rect 22220 2716 22286 2750
rect 22320 2716 22386 2750
rect 22420 2716 22486 2750
rect 22520 2716 22604 2750
rect 21904 2640 22604 2716
rect 23270 3250 23970 4000
rect 23270 3216 23346 3250
rect 23380 3216 23446 3250
rect 23480 3216 23546 3250
rect 23580 3216 23646 3250
rect 23680 3216 23746 3250
rect 23780 3216 23846 3250
rect 23880 3216 23970 3250
rect 23270 3150 23970 3216
rect 23270 3116 23346 3150
rect 23380 3116 23446 3150
rect 23480 3116 23546 3150
rect 23580 3116 23646 3150
rect 23680 3116 23746 3150
rect 23780 3116 23846 3150
rect 23880 3116 23970 3150
rect 23270 3050 23970 3116
rect 23270 3016 23346 3050
rect 23380 3016 23446 3050
rect 23480 3016 23546 3050
rect 23580 3016 23646 3050
rect 23680 3016 23746 3050
rect 23780 3016 23846 3050
rect 23880 3016 23970 3050
rect 23270 2950 23970 3016
rect 23270 2916 23346 2950
rect 23380 2916 23446 2950
rect 23480 2916 23546 2950
rect 23580 2916 23646 2950
rect 23680 2916 23746 2950
rect 23780 2916 23846 2950
rect 23880 2916 23970 2950
rect 23270 2850 23970 2916
rect 23270 2816 23346 2850
rect 23380 2816 23446 2850
rect 23480 2816 23546 2850
rect 23580 2816 23646 2850
rect 23680 2816 23746 2850
rect 23780 2816 23846 2850
rect 23880 2816 23970 2850
rect 23270 2750 23970 2816
rect 23270 2716 23346 2750
rect 23380 2716 23446 2750
rect 23480 2716 23546 2750
rect 23580 2716 23646 2750
rect 23680 2716 23746 2750
rect 23780 2716 23846 2750
rect 23880 2716 23970 2750
rect 22660 1980 22910 2290
rect 23270 1980 23970 2716
rect 24320 1980 24360 5020
rect 24680 4700 24720 5600
rect 24750 5560 24830 5570
rect 24750 5500 24760 5560
rect 24820 5500 24830 5560
rect 24750 5490 24830 5500
rect 24660 4690 24740 4700
rect 24660 4630 24670 4690
rect 24730 4630 24740 4690
rect 24660 4620 24740 4630
rect 24390 4580 24470 4590
rect 24390 4520 24400 4580
rect 24460 4520 24470 4580
rect 24390 4510 24470 4520
rect 24410 3030 24450 4510
rect 24770 4110 24810 5490
rect 24750 4100 24830 4110
rect 24750 4040 24760 4100
rect 24820 4040 24830 4100
rect 24750 4030 24830 4040
rect 24860 3650 24900 6830
rect 30270 6810 30370 6830
rect 30620 6890 30700 6900
rect 30620 6830 30630 6890
rect 30690 6830 30700 6890
rect 30620 6820 30700 6830
rect 25380 6780 25460 6790
rect 25380 6720 25390 6780
rect 25450 6720 25460 6780
rect 25380 6710 25460 6720
rect 25240 6680 25320 6690
rect 25240 6620 25250 6680
rect 25310 6620 25320 6680
rect 25240 6610 25320 6620
rect 26770 6670 26870 6690
rect 26770 6610 26790 6670
rect 26850 6610 26870 6670
rect 25060 6350 25140 6360
rect 25060 6290 25070 6350
rect 25130 6290 25140 6350
rect 25060 6280 25140 6290
rect 24930 5910 25010 5920
rect 24930 5850 24940 5910
rect 25000 5850 25010 5910
rect 24930 5840 25010 5850
rect 24950 4590 24990 5840
rect 24930 4580 25010 4590
rect 24930 4520 24940 4580
rect 25000 4520 25010 4580
rect 24930 4510 25010 4520
rect 24840 3640 24920 3650
rect 24840 3580 24850 3640
rect 24910 3580 24920 3640
rect 24840 3570 24920 3580
rect 24390 3020 24470 3030
rect 24390 2960 24400 3020
rect 24460 2960 24470 3020
rect 24390 2950 24470 2960
rect 20550 1890 24360 1980
rect 20550 1856 20626 1890
rect 20660 1856 20726 1890
rect 20760 1856 20826 1890
rect 20860 1856 20926 1890
rect 20960 1856 21026 1890
rect 21060 1856 21126 1890
rect 21160 1856 21986 1890
rect 22020 1856 22086 1890
rect 22120 1856 22186 1890
rect 22220 1856 22286 1890
rect 22320 1856 22386 1890
rect 22420 1856 22486 1890
rect 22520 1856 23346 1890
rect 23380 1856 23446 1890
rect 23480 1856 23546 1890
rect 23580 1856 23646 1890
rect 23680 1856 23746 1890
rect 23780 1856 23846 1890
rect 23880 1856 24360 1890
rect 20550 1790 24360 1856
rect 20550 1756 20626 1790
rect 20660 1756 20726 1790
rect 20760 1756 20826 1790
rect 20860 1756 20926 1790
rect 20960 1756 21026 1790
rect 21060 1756 21126 1790
rect 21160 1756 21986 1790
rect 22020 1756 22086 1790
rect 22120 1756 22186 1790
rect 22220 1756 22286 1790
rect 22320 1756 22386 1790
rect 22420 1756 22486 1790
rect 22520 1756 23346 1790
rect 23380 1756 23446 1790
rect 23480 1756 23546 1790
rect 23580 1756 23646 1790
rect 23680 1756 23746 1790
rect 23780 1756 23846 1790
rect 23880 1756 24360 1790
rect 20550 1690 24360 1756
rect 20550 1656 20626 1690
rect 20660 1656 20726 1690
rect 20760 1656 20826 1690
rect 20860 1656 20926 1690
rect 20960 1656 21026 1690
rect 21060 1656 21126 1690
rect 21160 1656 21986 1690
rect 22020 1656 22086 1690
rect 22120 1656 22186 1690
rect 22220 1656 22286 1690
rect 22320 1656 22386 1690
rect 22420 1656 22486 1690
rect 22520 1656 23346 1690
rect 23380 1656 23446 1690
rect 23480 1656 23546 1690
rect 23580 1656 23646 1690
rect 23680 1656 23746 1690
rect 23780 1656 23846 1690
rect 23880 1656 24360 1690
rect 20550 1590 24360 1656
rect 20550 1556 20626 1590
rect 20660 1556 20726 1590
rect 20760 1556 20826 1590
rect 20860 1556 20926 1590
rect 20960 1556 21026 1590
rect 21060 1556 21126 1590
rect 21160 1556 21986 1590
rect 22020 1556 22086 1590
rect 22120 1556 22186 1590
rect 22220 1556 22286 1590
rect 22320 1556 22386 1590
rect 22420 1556 22486 1590
rect 22520 1556 23346 1590
rect 23380 1556 23446 1590
rect 23480 1556 23546 1590
rect 23580 1556 23646 1590
rect 23680 1556 23746 1590
rect 23780 1556 23846 1590
rect 23880 1556 24360 1590
rect 20550 1490 24360 1556
rect 20550 1456 20626 1490
rect 20660 1456 20726 1490
rect 20760 1456 20826 1490
rect 20860 1456 20926 1490
rect 20960 1456 21026 1490
rect 21060 1456 21126 1490
rect 21160 1456 21986 1490
rect 22020 1456 22086 1490
rect 22120 1456 22186 1490
rect 22220 1456 22286 1490
rect 22320 1456 22386 1490
rect 22420 1456 22486 1490
rect 22520 1456 23346 1490
rect 23380 1456 23446 1490
rect 23480 1456 23546 1490
rect 23580 1456 23646 1490
rect 23680 1456 23746 1490
rect 23780 1456 23846 1490
rect 23880 1456 24360 1490
rect 20550 1390 24360 1456
rect 20550 1356 20626 1390
rect 20660 1356 20726 1390
rect 20760 1356 20826 1390
rect 20860 1356 20926 1390
rect 20960 1356 21026 1390
rect 21060 1356 21126 1390
rect 21160 1356 21986 1390
rect 22020 1356 22086 1390
rect 22120 1356 22186 1390
rect 22220 1356 22286 1390
rect 22320 1356 22386 1390
rect 22420 1356 22486 1390
rect 22520 1356 23346 1390
rect 23380 1356 23446 1390
rect 23480 1356 23546 1390
rect 23580 1356 23646 1390
rect 23680 1356 23746 1390
rect 23780 1356 23846 1390
rect 23880 1356 24360 1390
rect 20550 1280 24360 1356
rect 25080 730 25120 6280
rect 25150 4490 25230 4500
rect 25150 4430 25160 4490
rect 25220 4430 25230 4490
rect 25150 4420 25230 4430
rect 25170 1650 25210 4420
rect 25260 4340 25300 6610
rect 26770 6590 26870 6610
rect 25680 6570 25760 6580
rect 25680 6510 25690 6570
rect 25750 6510 25760 6570
rect 25680 6500 25760 6510
rect 25700 5810 25740 6500
rect 25990 6480 26070 6490
rect 25990 6420 26000 6480
rect 26060 6420 26070 6480
rect 25990 6410 26070 6420
rect 25680 5800 25760 5810
rect 25680 5740 25690 5800
rect 25750 5740 25760 5800
rect 25680 5730 25760 5740
rect 25490 4860 25570 4870
rect 25490 4800 25500 4860
rect 25560 4800 25570 4860
rect 25490 4790 25570 4800
rect 25620 4850 25700 4870
rect 25620 4810 25640 4850
rect 25680 4810 25700 4850
rect 25620 4790 25700 4810
rect 25750 4860 25830 4870
rect 25750 4800 25760 4860
rect 25820 4800 25830 4860
rect 25750 4790 25830 4800
rect 25510 4590 25550 4790
rect 25490 4580 25570 4590
rect 25490 4520 25500 4580
rect 25560 4520 25570 4580
rect 25490 4510 25570 4520
rect 25640 4500 25680 4790
rect 25620 4490 25700 4500
rect 25620 4430 25630 4490
rect 25690 4430 25700 4490
rect 25620 4420 25700 4430
rect 26010 4410 26050 6410
rect 27070 6360 27110 6370
rect 27790 6360 27830 6370
rect 28150 6360 28190 6370
rect 28870 6360 28910 6370
rect 29590 6360 29630 6370
rect 29850 6360 29890 6370
rect 29950 6360 29990 6370
rect 26320 6350 26400 6360
rect 26320 6290 26330 6350
rect 26390 6290 26400 6350
rect 26320 6280 26400 6290
rect 26690 6350 26770 6360
rect 26690 6290 26700 6350
rect 26760 6290 26770 6350
rect 26690 6280 26770 6290
rect 27050 6340 27130 6360
rect 27050 6300 27070 6340
rect 27110 6300 27130 6340
rect 27050 6280 27130 6300
rect 27410 6350 27490 6360
rect 27410 6290 27420 6350
rect 27480 6290 27490 6350
rect 27410 6280 27490 6290
rect 27770 6340 27850 6360
rect 27770 6300 27790 6340
rect 27830 6300 27850 6340
rect 27770 6280 27850 6300
rect 28130 6340 28210 6360
rect 28130 6300 28150 6340
rect 28190 6300 28210 6340
rect 28130 6280 28210 6300
rect 28490 6350 28570 6360
rect 28490 6290 28500 6350
rect 28560 6290 28570 6350
rect 28490 6280 28570 6290
rect 28850 6340 28930 6360
rect 28850 6300 28870 6340
rect 28910 6300 28930 6340
rect 28850 6280 28930 6300
rect 29210 6350 29290 6360
rect 29210 6290 29220 6350
rect 29280 6290 29290 6350
rect 29210 6280 29290 6290
rect 29570 6340 29650 6360
rect 29570 6300 29590 6340
rect 29630 6300 29650 6340
rect 29570 6280 29650 6300
rect 29830 6340 29900 6360
rect 29830 6300 29850 6340
rect 29890 6300 29900 6340
rect 29830 6280 29900 6300
rect 29940 6340 30010 6360
rect 29940 6300 29950 6340
rect 29990 6300 30010 6340
rect 29940 6280 30010 6300
rect 26150 6010 26230 6020
rect 26150 5950 26160 6010
rect 26220 5950 26230 6010
rect 26150 5940 26230 5950
rect 26510 6010 26590 6020
rect 26510 5950 26520 6010
rect 26580 5950 26590 6010
rect 26510 5940 26590 5950
rect 26870 6010 26950 6020
rect 26870 5950 26880 6010
rect 26940 5950 26950 6010
rect 26870 5940 26950 5950
rect 27230 6010 27310 6020
rect 27230 5950 27240 6010
rect 27300 5950 27310 6010
rect 27230 5940 27310 5950
rect 27590 6010 27670 6020
rect 27590 5950 27600 6010
rect 27660 5950 27670 6010
rect 27590 5940 27670 5950
rect 27950 6010 28030 6020
rect 27950 5950 27960 6010
rect 28020 5950 28030 6010
rect 27950 5940 28030 5950
rect 28310 6010 28390 6020
rect 28310 5950 28320 6010
rect 28380 5950 28390 6010
rect 28310 5940 28390 5950
rect 28670 6010 28750 6020
rect 28670 5950 28680 6010
rect 28740 5950 28750 6010
rect 28670 5940 28750 5950
rect 29030 6010 29110 6020
rect 29030 5950 29040 6010
rect 29100 5950 29110 6010
rect 29030 5940 29110 5950
rect 29390 6010 29470 6020
rect 29390 5950 29400 6010
rect 29460 5950 29470 6010
rect 29390 5940 29470 5950
rect 29750 6010 29830 6020
rect 29750 5950 29760 6010
rect 29820 5950 29830 6010
rect 29750 5940 29830 5950
rect 29890 6000 29950 6020
rect 29890 5960 29900 6000
rect 29940 5960 29950 6000
rect 29890 5940 29950 5960
rect 30110 6010 30190 6020
rect 30110 5950 30120 6010
rect 30180 5950 30190 6010
rect 30110 5940 30190 5950
rect 29900 5900 29940 5940
rect 29880 5890 29960 5900
rect 29880 5830 29890 5890
rect 29950 5830 29960 5890
rect 29880 5820 29960 5830
rect 30010 5890 30090 5900
rect 30010 5830 30020 5890
rect 30080 5830 30090 5890
rect 30010 5820 30090 5830
rect 26870 5430 26950 5440
rect 26870 5370 26880 5430
rect 26940 5370 26950 5430
rect 26870 5360 26950 5370
rect 27230 5430 27310 5440
rect 27230 5370 27240 5430
rect 27300 5370 27310 5430
rect 27230 5360 27310 5370
rect 27590 5430 27670 5440
rect 27590 5370 27600 5430
rect 27660 5370 27670 5430
rect 27590 5360 27670 5370
rect 27950 5430 28030 5440
rect 27950 5370 27960 5430
rect 28020 5370 28030 5430
rect 27950 5360 28030 5370
rect 28310 5430 28390 5440
rect 28310 5370 28320 5430
rect 28380 5370 28390 5430
rect 28310 5360 28390 5370
rect 28670 5430 28750 5440
rect 28670 5370 28680 5430
rect 28740 5370 28750 5430
rect 28670 5360 28750 5370
rect 29030 5430 29110 5440
rect 29030 5370 29040 5430
rect 29100 5370 29110 5430
rect 29030 5360 29110 5370
rect 29390 5430 29470 5440
rect 29390 5370 29400 5430
rect 29460 5370 29470 5430
rect 29390 5360 29470 5370
rect 26690 4680 26770 4700
rect 26690 4640 26710 4680
rect 26750 4640 26770 4680
rect 26690 4620 26770 4640
rect 27050 4680 27130 4700
rect 27050 4640 27070 4680
rect 27110 4640 27130 4680
rect 27050 4620 27130 4640
rect 27410 4680 27490 4700
rect 27410 4640 27430 4680
rect 27470 4640 27490 4680
rect 27410 4620 27490 4640
rect 27650 4680 27730 4700
rect 27650 4640 27670 4680
rect 27710 4640 27730 4680
rect 27650 4620 27730 4640
rect 27770 4690 27850 4700
rect 27770 4630 27780 4690
rect 27840 4630 27850 4690
rect 27770 4620 27850 4630
rect 28130 4680 28210 4700
rect 28130 4640 28150 4680
rect 28190 4640 28210 4680
rect 28130 4620 28210 4640
rect 28490 4690 28570 4700
rect 28490 4630 28500 4690
rect 28560 4630 28570 4690
rect 28490 4620 28570 4630
rect 28850 4680 28930 4700
rect 28850 4640 28870 4680
rect 28910 4640 28930 4680
rect 28850 4620 28930 4640
rect 29210 4680 29290 4700
rect 29210 4640 29230 4680
rect 29270 4640 29290 4680
rect 29210 4620 29290 4640
rect 29390 4680 29470 4700
rect 29390 4640 29410 4680
rect 29450 4640 29470 4680
rect 29390 4620 29470 4640
rect 29570 4680 29650 4700
rect 29570 4640 29590 4680
rect 29630 4640 29650 4680
rect 29570 4620 29650 4640
rect 26710 4410 26750 4620
rect 27070 4500 27110 4620
rect 27430 4590 27470 4620
rect 27410 4580 27490 4590
rect 27410 4520 27420 4580
rect 27480 4520 27490 4580
rect 27410 4510 27490 4520
rect 27050 4490 27130 4500
rect 27050 4430 27060 4490
rect 27120 4430 27130 4490
rect 27050 4420 27130 4430
rect 25990 4400 26070 4410
rect 25990 4340 26000 4400
rect 26060 4340 26070 4400
rect 25240 4330 25320 4340
rect 25990 4330 26070 4340
rect 26690 4400 26770 4410
rect 26690 4340 26700 4400
rect 26760 4340 26770 4400
rect 26690 4330 26770 4340
rect 25240 4270 25250 4330
rect 25310 4270 25320 4330
rect 25240 4260 25320 4270
rect 25410 4220 25490 4230
rect 25410 4160 25420 4220
rect 25480 4160 25490 4220
rect 25410 4150 25490 4160
rect 25650 4220 25730 4230
rect 25650 4160 25660 4220
rect 25720 4160 25730 4220
rect 25650 4150 25730 4160
rect 25890 4220 25970 4230
rect 25890 4160 25900 4220
rect 25960 4160 25970 4220
rect 25890 4150 25970 4160
rect 26130 4220 26210 4230
rect 26130 4160 26140 4220
rect 26200 4160 26210 4220
rect 26130 4150 26210 4160
rect 26370 4220 26450 4230
rect 26370 4160 26380 4220
rect 26440 4160 26450 4220
rect 26370 4150 26450 4160
rect 26610 4220 26690 4230
rect 26610 4160 26620 4220
rect 26680 4160 26690 4220
rect 26610 4150 26690 4160
rect 26850 4220 26930 4230
rect 26850 4160 26860 4220
rect 26920 4160 26930 4220
rect 26850 4150 26930 4160
rect 27090 4220 27170 4230
rect 27090 4160 27100 4220
rect 27160 4160 27170 4220
rect 27090 4150 27170 4160
rect 27330 4220 27410 4230
rect 27330 4160 27340 4220
rect 27400 4160 27410 4220
rect 27330 4150 27410 4160
rect 27570 4220 27650 4230
rect 27570 4160 27580 4220
rect 27640 4160 27650 4220
rect 27570 4150 27650 4160
rect 25430 4110 25470 4150
rect 25670 4110 25710 4150
rect 25910 4110 25950 4150
rect 26150 4110 26190 4150
rect 26390 4110 26430 4150
rect 26630 4110 26670 4150
rect 26870 4110 26910 4150
rect 27110 4110 27150 4150
rect 27350 4110 27390 4150
rect 27590 4110 27630 4150
rect 27690 4110 27730 4620
rect 28150 4410 28190 4620
rect 28870 4590 28910 4620
rect 28850 4580 28930 4590
rect 28850 4520 28860 4580
rect 28920 4520 28930 4580
rect 28850 4510 28930 4520
rect 29230 4500 29270 4620
rect 29410 4500 29450 4620
rect 29210 4490 29290 4500
rect 29210 4430 29220 4490
rect 29280 4430 29290 4490
rect 29210 4420 29290 4430
rect 29390 4490 29470 4500
rect 29390 4430 29400 4490
rect 29460 4430 29470 4490
rect 29390 4420 29470 4430
rect 29590 4410 29630 4620
rect 28130 4400 28210 4410
rect 28130 4340 28140 4400
rect 28200 4340 28210 4400
rect 28130 4330 28210 4340
rect 29570 4400 29650 4410
rect 29570 4340 29580 4400
rect 29640 4340 29650 4400
rect 29570 4330 29650 4340
rect 30030 4320 30070 5820
rect 30640 4500 30680 6820
rect 31240 6670 31320 6680
rect 31240 6610 31250 6670
rect 31310 6610 31320 6670
rect 31240 6600 31320 6610
rect 31150 5800 31230 5810
rect 31150 5740 31160 5800
rect 31220 5740 31230 5800
rect 31150 5730 31230 5740
rect 30620 4490 30700 4500
rect 30620 4430 30630 4490
rect 30690 4430 30700 4490
rect 30620 4420 30700 4430
rect 31060 4400 31140 4410
rect 31060 4340 31070 4400
rect 31130 4340 31140 4400
rect 31060 4330 31140 4340
rect 28570 4310 28650 4320
rect 28570 4250 28580 4310
rect 28640 4250 28650 4310
rect 28570 4240 28650 4250
rect 30010 4310 30090 4320
rect 30010 4250 30020 4310
rect 30080 4250 30090 4310
rect 30010 4240 30090 4250
rect 28590 4110 28630 4240
rect 28690 4220 28770 4230
rect 28690 4160 28700 4220
rect 28760 4160 28770 4220
rect 28690 4150 28770 4160
rect 28930 4220 29010 4230
rect 28930 4160 28940 4220
rect 29000 4160 29010 4220
rect 28930 4150 29010 4160
rect 29170 4220 29250 4230
rect 29170 4160 29180 4220
rect 29240 4160 29250 4220
rect 29170 4150 29250 4160
rect 29410 4220 29490 4230
rect 29410 4160 29420 4220
rect 29480 4160 29490 4220
rect 29410 4150 29490 4160
rect 29650 4220 29730 4230
rect 29650 4160 29660 4220
rect 29720 4160 29730 4220
rect 29650 4150 29730 4160
rect 29890 4220 29970 4230
rect 29890 4160 29900 4220
rect 29960 4160 29970 4220
rect 29890 4150 29970 4160
rect 30130 4220 30210 4230
rect 30130 4160 30140 4220
rect 30200 4160 30210 4220
rect 30130 4150 30210 4160
rect 30370 4220 30450 4230
rect 30370 4160 30380 4220
rect 30440 4160 30450 4220
rect 30370 4150 30450 4160
rect 30610 4220 30690 4230
rect 30610 4160 30620 4220
rect 30680 4160 30690 4220
rect 30610 4150 30690 4160
rect 30850 4220 30930 4230
rect 30850 4160 30860 4220
rect 30920 4160 30930 4220
rect 30850 4150 30930 4160
rect 28710 4110 28750 4150
rect 28950 4110 28990 4150
rect 29190 4110 29230 4150
rect 29430 4110 29470 4150
rect 29670 4110 29710 4150
rect 29910 4110 29950 4150
rect 30150 4110 30190 4150
rect 30390 4110 30430 4150
rect 30630 4110 30670 4150
rect 30870 4110 30910 4150
rect 25420 4090 25480 4110
rect 25420 4050 25430 4090
rect 25470 4050 25480 4090
rect 25420 4030 25480 4050
rect 25530 4100 25610 4110
rect 25530 4040 25540 4100
rect 25600 4040 25610 4100
rect 25530 4030 25610 4040
rect 25660 4090 25720 4110
rect 25660 4050 25670 4090
rect 25710 4050 25720 4090
rect 25660 4030 25720 4050
rect 25900 4090 25960 4110
rect 25900 4050 25910 4090
rect 25950 4050 25960 4090
rect 25900 4030 25960 4050
rect 26140 4090 26200 4110
rect 26140 4050 26150 4090
rect 26190 4050 26200 4090
rect 26140 4030 26200 4050
rect 26250 4100 26330 4110
rect 26250 4040 26260 4100
rect 26320 4040 26330 4100
rect 26250 4030 26330 4040
rect 26380 4090 26440 4110
rect 26380 4050 26390 4090
rect 26430 4050 26440 4090
rect 26380 4030 26440 4050
rect 26620 4090 26680 4110
rect 26620 4050 26630 4090
rect 26670 4050 26680 4090
rect 26620 4030 26680 4050
rect 26860 4090 26920 4110
rect 26860 4050 26870 4090
rect 26910 4050 26920 4090
rect 26860 4030 26920 4050
rect 26970 4100 27050 4110
rect 26970 4040 26980 4100
rect 27040 4040 27050 4100
rect 26970 4030 27050 4040
rect 27100 4090 27160 4110
rect 27100 4050 27110 4090
rect 27150 4050 27160 4090
rect 27100 4030 27160 4050
rect 27340 4090 27400 4110
rect 27340 4050 27350 4090
rect 27390 4050 27400 4090
rect 27340 4030 27400 4050
rect 27580 4090 27640 4110
rect 27580 4050 27590 4090
rect 27630 4050 27640 4090
rect 27580 4030 27640 4050
rect 27690 4100 27770 4110
rect 27690 4040 27700 4100
rect 27760 4040 27770 4100
rect 27690 4030 27770 4040
rect 27950 4100 28030 4110
rect 27950 4040 27960 4100
rect 28020 4040 28030 4100
rect 27950 4030 28030 4040
rect 28310 4100 28390 4110
rect 28310 4040 28320 4100
rect 28380 4040 28390 4100
rect 28310 4030 28390 4040
rect 28570 4100 28650 4110
rect 28570 4040 28580 4100
rect 28640 4040 28650 4100
rect 28570 4030 28650 4040
rect 28700 4090 28760 4110
rect 28700 4050 28710 4090
rect 28750 4050 28760 4090
rect 28700 4030 28760 4050
rect 28940 4090 29000 4110
rect 28940 4050 28950 4090
rect 28990 4050 29000 4090
rect 28940 4030 29000 4050
rect 29180 4090 29240 4110
rect 29180 4050 29190 4090
rect 29230 4050 29240 4090
rect 29180 4030 29240 4050
rect 29290 4100 29370 4110
rect 29290 4040 29300 4100
rect 29360 4040 29370 4100
rect 29290 4030 29370 4040
rect 29420 4090 29480 4110
rect 29420 4050 29430 4090
rect 29470 4050 29480 4090
rect 29420 4030 29480 4050
rect 29660 4090 29720 4110
rect 29660 4050 29670 4090
rect 29710 4050 29720 4090
rect 29660 4030 29720 4050
rect 29900 4090 29960 4110
rect 29900 4050 29910 4090
rect 29950 4050 29960 4090
rect 29900 4030 29960 4050
rect 30010 4100 30090 4110
rect 30010 4040 30020 4100
rect 30080 4040 30090 4100
rect 30010 4030 30090 4040
rect 30140 4090 30200 4110
rect 30140 4050 30150 4090
rect 30190 4050 30200 4090
rect 30140 4030 30200 4050
rect 30380 4090 30440 4110
rect 30380 4050 30390 4090
rect 30430 4050 30440 4090
rect 30380 4030 30440 4050
rect 30620 4090 30680 4110
rect 30620 4050 30630 4090
rect 30670 4050 30680 4090
rect 30620 4030 30680 4050
rect 30730 4100 30810 4110
rect 30730 4040 30740 4100
rect 30800 4040 30810 4100
rect 30730 4030 30810 4040
rect 30860 4090 30920 4110
rect 30860 4050 30870 4090
rect 30910 4050 30920 4090
rect 30860 4030 30920 4050
rect 25590 3750 25670 3770
rect 25590 3710 25610 3750
rect 25650 3710 25670 3750
rect 25590 3690 25670 3710
rect 25770 3760 25850 3770
rect 25770 3700 25780 3760
rect 25840 3700 25850 3760
rect 25770 3690 25850 3700
rect 26010 3750 26090 3770
rect 26010 3710 26030 3750
rect 26070 3710 26090 3750
rect 26010 3690 26090 3710
rect 26250 3750 26330 3770
rect 26250 3710 26270 3750
rect 26310 3710 26330 3750
rect 26250 3690 26330 3710
rect 26490 3760 26570 3770
rect 26490 3700 26500 3760
rect 26560 3700 26570 3760
rect 26490 3690 26570 3700
rect 26730 3750 26810 3770
rect 26730 3710 26750 3750
rect 26790 3710 26810 3750
rect 26730 3690 26810 3710
rect 26970 3750 27050 3770
rect 26970 3710 26990 3750
rect 27030 3710 27050 3750
rect 26970 3690 27050 3710
rect 27210 3760 27290 3770
rect 27210 3700 27220 3760
rect 27280 3700 27290 3760
rect 27210 3690 27290 3700
rect 27450 3750 27530 3770
rect 27450 3710 27470 3750
rect 27510 3710 27530 3750
rect 27450 3690 27530 3710
rect 27640 3750 27700 3770
rect 27640 3710 27650 3750
rect 27690 3710 27700 3750
rect 27640 3690 27700 3710
rect 25610 3650 25650 3690
rect 26030 3650 26070 3690
rect 26270 3650 26310 3690
rect 26750 3650 26790 3690
rect 26990 3650 27030 3690
rect 25590 3640 25670 3650
rect 25590 3580 25600 3640
rect 25660 3580 25670 3640
rect 25590 3570 25670 3580
rect 26010 3640 26090 3650
rect 26010 3580 26020 3640
rect 26080 3580 26090 3640
rect 26010 3570 26090 3580
rect 26250 3640 26330 3650
rect 26250 3580 26260 3640
rect 26320 3580 26330 3640
rect 26250 3570 26330 3580
rect 26730 3640 26810 3650
rect 26730 3580 26740 3640
rect 26800 3580 26810 3640
rect 26730 3570 26810 3580
rect 26970 3640 27050 3650
rect 26970 3580 26980 3640
rect 27040 3580 27050 3640
rect 26970 3570 27050 3580
rect 26990 3480 27030 3570
rect 26510 3470 26590 3480
rect 26390 3440 26470 3450
rect 26390 3380 26400 3440
rect 26460 3380 26470 3440
rect 26510 3410 26520 3470
rect 26580 3410 26590 3470
rect 26510 3400 26590 3410
rect 26990 3470 27070 3480
rect 26990 3410 27000 3470
rect 27060 3410 27070 3470
rect 26990 3400 27070 3410
rect 26390 3370 26470 3380
rect 26530 3360 26570 3400
rect 27010 3360 27050 3400
rect 27250 3360 27290 3690
rect 27470 3650 27510 3690
rect 27650 3650 27690 3690
rect 27450 3640 27530 3650
rect 27450 3580 27460 3640
rect 27520 3580 27530 3640
rect 27450 3570 27530 3580
rect 27630 3640 27710 3650
rect 27630 3580 27640 3640
rect 27700 3580 27710 3640
rect 27630 3570 27710 3580
rect 27470 3470 27550 3480
rect 27470 3410 27480 3470
rect 27540 3410 27550 3470
rect 27470 3400 27550 3410
rect 27490 3360 27530 3400
rect 26270 3350 26350 3360
rect 26270 3290 26280 3350
rect 26340 3290 26350 3350
rect 26270 3280 26350 3290
rect 26520 3340 26580 3360
rect 26520 3300 26530 3340
rect 26570 3300 26580 3340
rect 26520 3280 26580 3300
rect 26750 3350 26830 3360
rect 26750 3290 26760 3350
rect 26820 3290 26830 3350
rect 26750 3280 26830 3290
rect 27000 3340 27060 3360
rect 27000 3300 27010 3340
rect 27050 3300 27060 3340
rect 27000 3280 27060 3300
rect 27230 3350 27310 3360
rect 27230 3290 27240 3350
rect 27300 3290 27310 3350
rect 27230 3280 27310 3290
rect 27480 3340 27540 3360
rect 27480 3300 27490 3340
rect 27530 3300 27540 3340
rect 27480 3280 27540 3300
rect 26270 3110 26350 3120
rect 26270 3050 26280 3110
rect 26340 3050 26350 3110
rect 26270 3040 26350 3050
rect 26400 3100 26460 3120
rect 26400 3060 26410 3100
rect 26450 3060 26460 3100
rect 26400 3040 26460 3060
rect 26640 3100 26700 3120
rect 26640 3060 26650 3100
rect 26690 3060 26700 3100
rect 26640 3040 26700 3060
rect 26880 3100 26940 3120
rect 26880 3060 26890 3100
rect 26930 3060 26940 3100
rect 26880 3040 26940 3060
rect 27120 3100 27180 3120
rect 27120 3060 27130 3100
rect 27170 3060 27180 3100
rect 27120 3040 27180 3060
rect 27360 3100 27420 3120
rect 27360 3060 27370 3100
rect 27410 3060 27420 3100
rect 27360 3040 27420 3060
rect 26410 3000 26450 3040
rect 26650 3000 26690 3040
rect 26890 3000 26930 3040
rect 27130 3000 27170 3040
rect 27370 3000 27410 3040
rect 25790 2990 25870 3000
rect 25790 2930 25800 2990
rect 25860 2930 25870 2990
rect 25790 2920 25870 2930
rect 26390 2990 26470 3000
rect 26390 2930 26400 2990
rect 26460 2930 26470 2990
rect 26390 2920 26470 2930
rect 26630 2990 26710 3000
rect 26630 2930 26640 2990
rect 26700 2930 26710 2990
rect 26630 2920 26710 2930
rect 26870 2990 26950 3000
rect 26870 2930 26880 2990
rect 26940 2930 26950 2990
rect 26870 2920 26950 2930
rect 27110 2990 27190 3000
rect 27110 2930 27120 2990
rect 27180 2930 27190 2990
rect 27110 2920 27190 2930
rect 27350 2990 27430 3000
rect 27350 2930 27360 2990
rect 27420 2930 27430 2990
rect 27350 2920 27430 2930
rect 25810 2770 25850 2920
rect 25970 2790 26050 2800
rect 25790 2750 25870 2770
rect 25790 2710 25810 2750
rect 25850 2710 25870 2750
rect 25970 2730 25980 2790
rect 26040 2730 26050 2790
rect 25970 2720 26050 2730
rect 26210 2790 26290 2800
rect 26210 2730 26220 2790
rect 26280 2730 26290 2790
rect 26210 2720 26290 2730
rect 26450 2790 26530 2800
rect 26450 2730 26460 2790
rect 26520 2730 26530 2790
rect 26450 2720 26530 2730
rect 26690 2790 26770 2800
rect 26690 2730 26700 2790
rect 26760 2730 26770 2790
rect 26690 2720 26770 2730
rect 27170 2790 27250 2800
rect 27170 2730 27180 2790
rect 27240 2730 27250 2790
rect 27170 2720 27250 2730
rect 27410 2790 27490 2800
rect 27410 2730 27420 2790
rect 27480 2730 27490 2790
rect 27410 2720 27490 2730
rect 27650 2790 27730 2800
rect 27650 2730 27660 2790
rect 27720 2730 27730 2790
rect 27970 2770 28010 4030
rect 28330 2770 28370 4030
rect 28640 3750 28700 3770
rect 28640 3710 28650 3750
rect 28690 3710 28700 3750
rect 28640 3690 28700 3710
rect 28810 3750 28890 3770
rect 28810 3710 28830 3750
rect 28870 3710 28890 3750
rect 28810 3690 28890 3710
rect 29050 3760 29130 3770
rect 29050 3700 29060 3760
rect 29120 3700 29130 3760
rect 29050 3690 29130 3700
rect 29290 3750 29370 3770
rect 29290 3710 29310 3750
rect 29350 3710 29370 3750
rect 29290 3690 29370 3710
rect 29530 3750 29610 3770
rect 29530 3710 29550 3750
rect 29590 3710 29610 3750
rect 29530 3690 29610 3710
rect 29770 3760 29850 3770
rect 29770 3700 29780 3760
rect 29840 3700 29850 3760
rect 29770 3690 29850 3700
rect 30010 3750 30090 3770
rect 30010 3710 30030 3750
rect 30070 3710 30090 3750
rect 30010 3690 30090 3710
rect 30250 3750 30330 3770
rect 30250 3710 30270 3750
rect 30310 3710 30330 3750
rect 30250 3690 30330 3710
rect 30490 3760 30570 3770
rect 30490 3700 30500 3760
rect 30560 3700 30570 3760
rect 30490 3690 30570 3700
rect 30670 3750 30750 3770
rect 30670 3710 30690 3750
rect 30730 3710 30750 3750
rect 30670 3690 30750 3710
rect 28650 3650 28690 3690
rect 28830 3650 28870 3690
rect 28630 3640 28710 3650
rect 28630 3580 28640 3640
rect 28700 3580 28710 3640
rect 28630 3570 28710 3580
rect 28810 3640 28890 3650
rect 28810 3580 28820 3640
rect 28880 3580 28890 3640
rect 28810 3570 28890 3580
rect 28790 3470 28870 3480
rect 28790 3410 28800 3470
rect 28860 3410 28870 3470
rect 28790 3400 28870 3410
rect 28810 3360 28850 3400
rect 29050 3360 29090 3690
rect 29310 3650 29350 3690
rect 29550 3650 29590 3690
rect 30030 3650 30070 3690
rect 30270 3650 30310 3690
rect 30690 3650 30730 3690
rect 29290 3640 29370 3650
rect 29290 3580 29300 3640
rect 29360 3580 29370 3640
rect 29290 3570 29370 3580
rect 29530 3640 29610 3650
rect 29530 3580 29540 3640
rect 29600 3580 29610 3640
rect 29530 3570 29610 3580
rect 30010 3640 30090 3650
rect 30010 3580 30020 3640
rect 30080 3580 30090 3640
rect 30010 3570 30090 3580
rect 30250 3640 30330 3650
rect 30250 3580 30260 3640
rect 30320 3580 30330 3640
rect 30250 3570 30330 3580
rect 30670 3640 30750 3650
rect 30670 3580 30680 3640
rect 30740 3580 30750 3640
rect 30670 3570 30750 3580
rect 29310 3480 29350 3570
rect 29270 3470 29350 3480
rect 29270 3410 29280 3470
rect 29340 3410 29350 3470
rect 29270 3400 29350 3410
rect 29750 3470 29830 3480
rect 29750 3410 29760 3470
rect 29820 3410 29830 3470
rect 31080 3450 31120 4330
rect 29750 3400 29830 3410
rect 29870 3440 29950 3450
rect 29290 3360 29330 3400
rect 29770 3360 29810 3400
rect 29870 3380 29880 3440
rect 29940 3380 29950 3440
rect 29870 3370 29950 3380
rect 31060 3440 31140 3450
rect 31060 3380 31070 3440
rect 31130 3380 31140 3440
rect 31060 3370 31140 3380
rect 28800 3340 28860 3360
rect 28800 3300 28810 3340
rect 28850 3300 28860 3340
rect 28800 3280 28860 3300
rect 29030 3350 29110 3360
rect 29030 3290 29040 3350
rect 29100 3290 29110 3350
rect 29030 3280 29110 3290
rect 29280 3340 29340 3360
rect 29280 3300 29290 3340
rect 29330 3300 29340 3340
rect 29280 3280 29340 3300
rect 29510 3350 29590 3360
rect 29510 3290 29520 3350
rect 29580 3290 29590 3350
rect 29510 3280 29590 3290
rect 29760 3340 29820 3360
rect 29760 3300 29770 3340
rect 29810 3300 29820 3340
rect 29760 3280 29820 3300
rect 29990 3350 30070 3360
rect 29990 3290 30000 3350
rect 30060 3290 30070 3350
rect 29990 3280 30070 3290
rect 31170 3120 31210 5730
rect 31260 3650 31300 6600
rect 31240 3640 31320 3650
rect 31240 3580 31250 3640
rect 31310 3580 31320 3640
rect 31240 3570 31320 3580
rect 28920 3100 28980 3120
rect 28920 3060 28930 3100
rect 28970 3060 28980 3100
rect 28920 3040 28980 3060
rect 29160 3100 29220 3120
rect 29160 3060 29170 3100
rect 29210 3060 29220 3100
rect 29160 3040 29220 3060
rect 29400 3100 29460 3120
rect 29400 3060 29410 3100
rect 29450 3060 29460 3100
rect 29400 3040 29460 3060
rect 29640 3100 29700 3120
rect 29640 3060 29650 3100
rect 29690 3060 29700 3100
rect 29640 3040 29700 3060
rect 29880 3100 29940 3120
rect 29880 3060 29890 3100
rect 29930 3060 29940 3100
rect 29880 3040 29940 3060
rect 29990 3110 30070 3120
rect 29990 3050 30000 3110
rect 30060 3050 30070 3110
rect 29990 3040 30070 3050
rect 31150 3110 31230 3120
rect 31150 3050 31160 3110
rect 31220 3050 31230 3110
rect 31150 3040 31230 3050
rect 28930 3000 28970 3040
rect 29170 3000 29210 3040
rect 29410 3000 29450 3040
rect 29650 3000 29690 3040
rect 29890 3000 29930 3040
rect 28910 2990 28990 3000
rect 28910 2930 28920 2990
rect 28980 2930 28990 2990
rect 28910 2920 28990 2930
rect 29150 2990 29230 3000
rect 29150 2930 29160 2990
rect 29220 2930 29230 2990
rect 29150 2920 29230 2930
rect 29390 2990 29470 3000
rect 29390 2930 29400 2990
rect 29460 2930 29470 2990
rect 29390 2920 29470 2930
rect 29630 2990 29710 3000
rect 29630 2930 29640 2990
rect 29700 2930 29710 2990
rect 29630 2920 29710 2930
rect 29870 2990 29950 3000
rect 29870 2930 29880 2990
rect 29940 2930 29950 2990
rect 29870 2920 29950 2930
rect 30470 2990 30550 3000
rect 30470 2930 30480 2990
rect 30540 2930 30550 2990
rect 30470 2920 30550 2930
rect 28610 2790 28690 2800
rect 27650 2720 27730 2730
rect 27950 2750 28030 2770
rect 25790 2690 25870 2710
rect 27950 2710 27970 2750
rect 28010 2710 28030 2750
rect 27950 2690 28030 2710
rect 28310 2750 28390 2770
rect 28310 2710 28330 2750
rect 28370 2710 28390 2750
rect 28610 2730 28620 2790
rect 28680 2730 28690 2790
rect 28610 2720 28690 2730
rect 28850 2790 28930 2800
rect 28850 2730 28860 2790
rect 28920 2730 28930 2790
rect 28850 2720 28930 2730
rect 29090 2790 29170 2800
rect 29090 2730 29100 2790
rect 29160 2730 29170 2790
rect 29090 2720 29170 2730
rect 29570 2790 29650 2800
rect 29570 2730 29580 2790
rect 29640 2730 29650 2790
rect 29570 2720 29650 2730
rect 29810 2790 29890 2800
rect 29810 2730 29820 2790
rect 29880 2730 29890 2790
rect 29810 2720 29890 2730
rect 30050 2790 30130 2800
rect 30050 2730 30060 2790
rect 30120 2730 30130 2790
rect 30050 2720 30130 2730
rect 30290 2790 30370 2800
rect 30290 2730 30300 2790
rect 30360 2730 30370 2790
rect 30490 2770 30530 2920
rect 30290 2720 30370 2730
rect 30470 2750 30550 2770
rect 28310 2690 28390 2710
rect 30470 2710 30490 2750
rect 30530 2710 30550 2750
rect 30470 2690 30550 2710
rect 26870 2160 26950 2170
rect 26870 2100 26880 2160
rect 26940 2100 26950 2160
rect 26870 2090 26950 2100
rect 29390 2160 29470 2170
rect 29390 2100 29400 2160
rect 29460 2100 29470 2160
rect 29390 2090 29470 2100
rect 26050 1810 26130 1820
rect 26050 1750 26060 1810
rect 26120 1750 26130 1810
rect 26050 1740 26130 1750
rect 26210 1810 26290 1820
rect 26210 1750 26220 1810
rect 26280 1750 26290 1810
rect 26210 1740 26290 1750
rect 26370 1810 26450 1820
rect 26370 1750 26380 1810
rect 26440 1750 26450 1810
rect 26370 1740 26450 1750
rect 26530 1810 26610 1820
rect 26530 1750 26540 1810
rect 26600 1750 26610 1810
rect 26530 1740 26610 1750
rect 26690 1810 26770 1820
rect 26690 1750 26700 1810
rect 26760 1750 26770 1810
rect 26690 1740 26770 1750
rect 26850 1810 26930 1820
rect 26850 1750 26860 1810
rect 26920 1750 26930 1810
rect 26850 1740 26930 1750
rect 27010 1810 27090 1820
rect 27010 1750 27020 1810
rect 27080 1750 27090 1810
rect 27010 1740 27090 1750
rect 27170 1810 27250 1820
rect 27170 1750 27180 1810
rect 27240 1750 27250 1810
rect 27170 1740 27250 1750
rect 27330 1810 27410 1820
rect 27330 1750 27340 1810
rect 27400 1750 27410 1810
rect 27330 1740 27410 1750
rect 27490 1810 27570 1820
rect 27490 1750 27500 1810
rect 27560 1750 27570 1810
rect 27490 1740 27570 1750
rect 27650 1810 27730 1820
rect 27650 1750 27660 1810
rect 27720 1750 27730 1810
rect 27650 1740 27730 1750
rect 27810 1810 27890 1820
rect 27810 1750 27820 1810
rect 27880 1750 27890 1810
rect 27810 1740 27890 1750
rect 27970 1810 28050 1820
rect 27970 1750 27980 1810
rect 28040 1750 28050 1810
rect 27970 1740 28050 1750
rect 28130 1810 28210 1820
rect 28130 1750 28140 1810
rect 28200 1750 28210 1810
rect 28130 1740 28210 1750
rect 28290 1810 28370 1820
rect 28290 1750 28300 1810
rect 28360 1750 28370 1810
rect 28290 1740 28370 1750
rect 28450 1810 28530 1820
rect 28450 1750 28460 1810
rect 28520 1750 28530 1810
rect 28450 1740 28530 1750
rect 28610 1810 28690 1820
rect 28610 1750 28620 1810
rect 28680 1750 28690 1810
rect 28610 1740 28690 1750
rect 28770 1810 28850 1820
rect 28770 1750 28780 1810
rect 28840 1750 28850 1810
rect 28770 1740 28850 1750
rect 28930 1810 29010 1820
rect 28930 1750 28940 1810
rect 29000 1750 29010 1810
rect 28930 1740 29010 1750
rect 29090 1810 29170 1820
rect 29090 1750 29100 1810
rect 29160 1750 29170 1810
rect 29090 1740 29170 1750
rect 29250 1810 29330 1820
rect 29250 1750 29260 1810
rect 29320 1750 29330 1810
rect 29250 1740 29330 1750
rect 29410 1810 29490 1820
rect 29410 1750 29420 1810
rect 29480 1750 29490 1810
rect 29410 1740 29490 1750
rect 29570 1810 29650 1820
rect 29570 1750 29580 1810
rect 29640 1750 29650 1810
rect 29570 1740 29650 1750
rect 29730 1810 29810 1820
rect 29730 1750 29740 1810
rect 29800 1750 29810 1810
rect 29730 1740 29810 1750
rect 29890 1810 29970 1820
rect 29890 1750 29900 1810
rect 29960 1750 29970 1810
rect 29890 1740 29970 1750
rect 30050 1810 30130 1820
rect 30050 1750 30060 1810
rect 30120 1750 30130 1810
rect 30050 1740 30130 1750
rect 25150 1640 25230 1650
rect 25150 1580 25160 1640
rect 25220 1580 25230 1640
rect 25150 1570 25230 1580
rect 25970 1640 26050 1650
rect 25970 1580 25980 1640
rect 26040 1580 26050 1640
rect 25970 1570 26050 1580
rect 30370 1640 30450 1650
rect 30370 1580 30380 1640
rect 30440 1580 30450 1640
rect 30370 1570 30450 1580
rect 25750 1260 25830 1270
rect 25750 1200 25760 1260
rect 25820 1200 25830 1260
rect 25750 1190 25830 1200
rect 26110 1260 26190 1270
rect 26110 1200 26120 1260
rect 26180 1200 26190 1260
rect 26110 1190 26190 1200
rect 26470 1260 26550 1270
rect 26470 1200 26480 1260
rect 26540 1200 26550 1260
rect 26470 1190 26550 1200
rect 27590 1260 27670 1270
rect 27590 1200 27600 1260
rect 27660 1200 27670 1260
rect 27590 1190 27670 1200
rect 27950 1260 28030 1270
rect 27950 1200 27960 1260
rect 28020 1200 28030 1260
rect 27950 1190 28030 1200
rect 28310 1260 28390 1270
rect 28310 1200 28320 1260
rect 28380 1200 28390 1260
rect 28310 1190 28390 1200
rect 28670 1260 28750 1270
rect 28670 1200 28680 1260
rect 28740 1200 28750 1260
rect 28670 1190 28750 1200
rect 29750 1260 29830 1270
rect 29750 1200 29760 1260
rect 29820 1200 29830 1260
rect 29750 1190 29830 1200
rect 30110 1260 30190 1270
rect 30110 1200 30120 1260
rect 30180 1200 30190 1260
rect 30110 1190 30190 1200
rect 30470 1260 30550 1270
rect 30470 1200 30480 1260
rect 30540 1200 30550 1260
rect 30470 1190 30550 1200
rect 25570 920 25650 930
rect 25570 860 25580 920
rect 25640 860 25650 920
rect 25570 850 25650 860
rect 25930 910 26010 930
rect 25930 870 25950 910
rect 25990 870 26010 910
rect 25930 850 26010 870
rect 26290 920 26370 930
rect 26290 860 26300 920
rect 26360 860 26370 920
rect 26290 850 26370 860
rect 26650 910 26730 930
rect 26650 870 26670 910
rect 26710 870 26730 910
rect 26650 850 26730 870
rect 27410 910 27490 930
rect 27410 870 27430 910
rect 27470 870 27490 910
rect 27410 850 27490 870
rect 28130 920 28210 930
rect 28130 860 28140 920
rect 28200 860 28210 920
rect 28130 850 28210 860
rect 28490 920 28570 930
rect 28490 860 28500 920
rect 28560 860 28570 920
rect 28490 850 28570 860
rect 28850 920 28930 930
rect 28850 860 28860 920
rect 28920 860 28930 920
rect 28850 850 28930 860
rect 29570 920 29650 930
rect 29570 860 29580 920
rect 29640 860 29650 920
rect 29570 850 29650 860
rect 29930 910 30010 930
rect 29930 870 29950 910
rect 29990 870 30010 910
rect 29930 850 30010 870
rect 30290 920 30370 930
rect 30290 860 30300 920
rect 30360 860 30370 920
rect 30290 850 30370 860
rect 30650 910 30730 930
rect 30650 870 30670 910
rect 30710 870 30730 910
rect 30650 850 30730 870
rect 25950 820 25990 850
rect 26670 820 26710 850
rect 25930 810 26010 820
rect 25930 750 25940 810
rect 26000 750 26010 810
rect 25930 740 26010 750
rect 26650 810 26730 820
rect 26650 750 26660 810
rect 26720 750 26730 810
rect 26650 740 26730 750
rect 27430 730 27470 850
rect 29950 820 29990 850
rect 30670 820 30710 850
rect 29930 810 30010 820
rect 29930 750 29940 810
rect 30000 750 30010 810
rect 29930 740 30010 750
rect 30650 810 30730 820
rect 30650 750 30660 810
rect 30720 750 30730 810
rect 30650 740 30730 750
rect 25060 720 25140 730
rect 25060 660 25070 720
rect 25130 660 25140 720
rect 25060 650 25140 660
rect 27410 720 27490 730
rect 27410 660 27420 720
rect 27480 660 27490 720
rect 27410 650 27490 660
rect 26550 -110 26590 640
rect 27630 -110 27670 640
rect 27990 -110 28030 640
rect 29430 -110 29470 640
<< via1 >>
rect 22532 6990 22592 7050
rect 19980 6830 20040 6890
rect 21890 6830 21950 6890
rect 19890 6720 19950 6780
rect 19890 5630 19950 5690
rect 22420 6620 22480 6680
rect 22330 6510 22390 6570
rect 20102 6400 20172 6410
rect 20102 6350 20112 6400
rect 20112 6350 20162 6400
rect 20162 6350 20172 6400
rect 20102 6340 20172 6350
rect 20102 6280 20172 6290
rect 20102 6230 20112 6280
rect 20112 6230 20162 6280
rect 20162 6230 20172 6280
rect 20102 6220 20172 6230
rect 22330 6140 22390 6200
rect 20102 6120 20172 6130
rect 20102 6070 20112 6120
rect 20112 6070 20162 6120
rect 20162 6070 20172 6120
rect 20102 6060 20172 6070
rect 20102 6000 20172 6010
rect 20102 5950 20112 6000
rect 20112 5950 20162 6000
rect 20162 5950 20172 6000
rect 20102 5940 20172 5950
rect 21840 5760 21900 5820
rect 22000 5760 22060 5820
rect 22160 5760 22220 5820
rect 28890 6930 28950 6990
rect 23290 6830 23350 6890
rect 24850 6840 24910 6900
rect 30290 6830 30350 6890
rect 22532 6390 22602 6400
rect 22532 6340 22542 6390
rect 22542 6340 22592 6390
rect 22592 6340 22602 6390
rect 22532 6330 22602 6340
rect 22532 6270 22602 6280
rect 22532 6220 22542 6270
rect 22542 6220 22592 6270
rect 22592 6220 22602 6270
rect 22532 6210 22602 6220
rect 24670 5910 24740 5920
rect 24670 5860 24680 5910
rect 24680 5860 24730 5910
rect 24730 5860 24740 5910
rect 24670 5850 24740 5860
rect 24670 5790 24740 5800
rect 24670 5740 24680 5790
rect 24680 5740 24730 5790
rect 24730 5740 24740 5790
rect 24670 5730 24740 5740
rect 20112 5680 20182 5690
rect 20112 5630 20122 5680
rect 20122 5630 20172 5680
rect 20172 5630 20182 5680
rect 20112 5620 20182 5630
rect 21458 5680 21528 5690
rect 21458 5630 21468 5680
rect 21468 5630 21518 5680
rect 21518 5630 21528 5680
rect 21458 5620 21528 5630
rect 22420 5620 22480 5680
rect 22532 5670 22602 5680
rect 22532 5620 22542 5670
rect 22542 5620 22592 5670
rect 22592 5620 22602 5670
rect 22532 5610 22602 5620
rect 23930 5670 24000 5680
rect 23930 5620 23940 5670
rect 23940 5620 23990 5670
rect 23990 5620 24000 5670
rect 23930 5610 24000 5620
rect 24670 5610 24730 5670
rect 19980 5510 20040 5570
rect 20112 5560 20182 5570
rect 20112 5510 20122 5560
rect 20122 5510 20172 5560
rect 20172 5510 20182 5560
rect 20112 5500 20182 5510
rect 21458 5560 21528 5570
rect 21458 5510 21468 5560
rect 21468 5510 21518 5560
rect 21518 5510 21528 5560
rect 21458 5500 21528 5510
rect 22532 5030 22592 5090
rect 24310 5030 24370 5090
rect 19790 2980 19850 3040
rect 19920 3030 19980 3040
rect 19920 2990 19930 3030
rect 19930 2990 19970 3030
rect 19970 2990 19980 3030
rect 19920 2980 19980 2990
rect 22540 2960 22594 3020
rect 24760 5500 24820 5560
rect 24670 4630 24730 4690
rect 24400 4520 24460 4580
rect 24760 4040 24820 4100
rect 30630 6830 30690 6890
rect 25390 6720 25450 6780
rect 25250 6620 25310 6680
rect 26790 6610 26850 6670
rect 25070 6290 25130 6350
rect 24940 5850 25000 5910
rect 24940 4520 25000 4580
rect 24850 3580 24910 3640
rect 24400 2960 24460 3020
rect 25160 4430 25220 4490
rect 25690 6510 25750 6570
rect 26000 6420 26060 6480
rect 25690 5740 25750 5800
rect 25500 4850 25560 4860
rect 25500 4810 25510 4850
rect 25510 4810 25550 4850
rect 25550 4810 25560 4850
rect 25500 4800 25560 4810
rect 25760 4850 25820 4860
rect 25760 4810 25770 4850
rect 25770 4810 25810 4850
rect 25810 4810 25820 4850
rect 25760 4800 25820 4810
rect 25500 4520 25560 4580
rect 25630 4430 25690 4490
rect 26330 6340 26390 6350
rect 26330 6300 26340 6340
rect 26340 6300 26380 6340
rect 26380 6300 26390 6340
rect 26330 6290 26390 6300
rect 26700 6340 26760 6350
rect 26700 6300 26710 6340
rect 26710 6300 26750 6340
rect 26750 6300 26760 6340
rect 26700 6290 26760 6300
rect 27420 6340 27480 6350
rect 27420 6300 27430 6340
rect 27430 6300 27470 6340
rect 27470 6300 27480 6340
rect 27420 6290 27480 6300
rect 28500 6340 28560 6350
rect 28500 6300 28510 6340
rect 28510 6300 28550 6340
rect 28550 6300 28560 6340
rect 28500 6290 28560 6300
rect 29220 6340 29280 6350
rect 29220 6300 29230 6340
rect 29230 6300 29270 6340
rect 29270 6300 29280 6340
rect 29220 6290 29280 6300
rect 26160 6000 26220 6010
rect 26160 5960 26170 6000
rect 26170 5960 26210 6000
rect 26210 5960 26220 6000
rect 26160 5950 26220 5960
rect 26520 6000 26580 6010
rect 26520 5960 26530 6000
rect 26530 5960 26570 6000
rect 26570 5960 26580 6000
rect 26520 5950 26580 5960
rect 26880 6000 26940 6010
rect 26880 5960 26890 6000
rect 26890 5960 26930 6000
rect 26930 5960 26940 6000
rect 26880 5950 26940 5960
rect 27240 6000 27300 6010
rect 27240 5960 27250 6000
rect 27250 5960 27290 6000
rect 27290 5960 27300 6000
rect 27240 5950 27300 5960
rect 27600 6000 27660 6010
rect 27600 5960 27610 6000
rect 27610 5960 27650 6000
rect 27650 5960 27660 6000
rect 27600 5950 27660 5960
rect 27960 6000 28020 6010
rect 27960 5960 27970 6000
rect 27970 5960 28010 6000
rect 28010 5960 28020 6000
rect 27960 5950 28020 5960
rect 28320 6000 28380 6010
rect 28320 5960 28330 6000
rect 28330 5960 28370 6000
rect 28370 5960 28380 6000
rect 28320 5950 28380 5960
rect 28680 6000 28740 6010
rect 28680 5960 28690 6000
rect 28690 5960 28730 6000
rect 28730 5960 28740 6000
rect 28680 5950 28740 5960
rect 29040 6000 29100 6010
rect 29040 5960 29050 6000
rect 29050 5960 29090 6000
rect 29090 5960 29100 6000
rect 29040 5950 29100 5960
rect 29400 6000 29460 6010
rect 29400 5960 29410 6000
rect 29410 5960 29450 6000
rect 29450 5960 29460 6000
rect 29400 5950 29460 5960
rect 29760 6000 29820 6010
rect 29760 5960 29770 6000
rect 29770 5960 29810 6000
rect 29810 5960 29820 6000
rect 29760 5950 29820 5960
rect 30120 6000 30180 6010
rect 30120 5960 30130 6000
rect 30130 5960 30170 6000
rect 30170 5960 30180 6000
rect 30120 5950 30180 5960
rect 29890 5830 29950 5890
rect 30020 5830 30080 5890
rect 26880 5420 26940 5430
rect 26880 5380 26890 5420
rect 26890 5380 26930 5420
rect 26930 5380 26940 5420
rect 26880 5370 26940 5380
rect 27240 5420 27300 5430
rect 27240 5380 27250 5420
rect 27250 5380 27290 5420
rect 27290 5380 27300 5420
rect 27240 5370 27300 5380
rect 27600 5420 27660 5430
rect 27600 5380 27610 5420
rect 27610 5380 27650 5420
rect 27650 5380 27660 5420
rect 27600 5370 27660 5380
rect 27960 5420 28020 5430
rect 27960 5380 27970 5420
rect 27970 5380 28010 5420
rect 28010 5380 28020 5420
rect 27960 5370 28020 5380
rect 28320 5420 28380 5430
rect 28320 5380 28330 5420
rect 28330 5380 28370 5420
rect 28370 5380 28380 5420
rect 28320 5370 28380 5380
rect 28680 5420 28740 5430
rect 28680 5380 28690 5420
rect 28690 5380 28730 5420
rect 28730 5380 28740 5420
rect 28680 5370 28740 5380
rect 29040 5420 29100 5430
rect 29040 5380 29050 5420
rect 29050 5380 29090 5420
rect 29090 5380 29100 5420
rect 29040 5370 29100 5380
rect 29400 5420 29460 5430
rect 29400 5380 29410 5420
rect 29410 5380 29450 5420
rect 29450 5380 29460 5420
rect 29400 5370 29460 5380
rect 27780 4680 27840 4690
rect 27780 4640 27790 4680
rect 27790 4640 27830 4680
rect 27830 4640 27840 4680
rect 27780 4630 27840 4640
rect 28500 4680 28560 4690
rect 28500 4640 28510 4680
rect 28510 4640 28550 4680
rect 28550 4640 28560 4680
rect 28500 4630 28560 4640
rect 27420 4520 27480 4580
rect 27060 4430 27120 4490
rect 26000 4340 26060 4400
rect 26700 4340 26760 4400
rect 25250 4270 25310 4330
rect 25420 4160 25480 4220
rect 25660 4160 25720 4220
rect 25900 4160 25960 4220
rect 26140 4160 26200 4220
rect 26380 4160 26440 4220
rect 26620 4160 26680 4220
rect 26860 4160 26920 4220
rect 27100 4160 27160 4220
rect 27340 4160 27400 4220
rect 27580 4160 27640 4220
rect 28860 4520 28920 4580
rect 29220 4430 29280 4490
rect 29400 4430 29460 4490
rect 28140 4340 28200 4400
rect 29580 4340 29640 4400
rect 31250 6610 31310 6670
rect 31160 5740 31220 5800
rect 30630 4430 30690 4490
rect 31070 4340 31130 4400
rect 28580 4250 28640 4310
rect 30020 4250 30080 4310
rect 28700 4210 28760 4220
rect 28700 4170 28710 4210
rect 28710 4170 28750 4210
rect 28750 4170 28760 4210
rect 28700 4160 28760 4170
rect 28940 4210 29000 4220
rect 28940 4170 28950 4210
rect 28950 4170 28990 4210
rect 28990 4170 29000 4210
rect 28940 4160 29000 4170
rect 29180 4210 29240 4220
rect 29180 4170 29190 4210
rect 29190 4170 29230 4210
rect 29230 4170 29240 4210
rect 29180 4160 29240 4170
rect 29420 4210 29480 4220
rect 29420 4170 29430 4210
rect 29430 4170 29470 4210
rect 29470 4170 29480 4210
rect 29420 4160 29480 4170
rect 29660 4210 29720 4220
rect 29660 4170 29670 4210
rect 29670 4170 29710 4210
rect 29710 4170 29720 4210
rect 29660 4160 29720 4170
rect 29900 4210 29960 4220
rect 29900 4170 29910 4210
rect 29910 4170 29950 4210
rect 29950 4170 29960 4210
rect 29900 4160 29960 4170
rect 30140 4210 30200 4220
rect 30140 4170 30150 4210
rect 30150 4170 30190 4210
rect 30190 4170 30200 4210
rect 30140 4160 30200 4170
rect 30380 4210 30440 4220
rect 30380 4170 30390 4210
rect 30390 4170 30430 4210
rect 30430 4170 30440 4210
rect 30380 4160 30440 4170
rect 30620 4210 30680 4220
rect 30620 4170 30630 4210
rect 30630 4170 30670 4210
rect 30670 4170 30680 4210
rect 30620 4160 30680 4170
rect 30860 4210 30920 4220
rect 30860 4170 30870 4210
rect 30870 4170 30910 4210
rect 30910 4170 30920 4210
rect 30860 4160 30920 4170
rect 25540 4090 25600 4100
rect 25540 4050 25550 4090
rect 25550 4050 25590 4090
rect 25590 4050 25600 4090
rect 25540 4040 25600 4050
rect 26260 4090 26320 4100
rect 26260 4050 26270 4090
rect 26270 4050 26310 4090
rect 26310 4050 26320 4090
rect 26260 4040 26320 4050
rect 26980 4090 27040 4100
rect 26980 4050 26990 4090
rect 26990 4050 27030 4090
rect 27030 4050 27040 4090
rect 26980 4040 27040 4050
rect 27700 4090 27760 4100
rect 27700 4050 27710 4090
rect 27710 4050 27750 4090
rect 27750 4050 27760 4090
rect 27700 4040 27760 4050
rect 27960 4040 28020 4100
rect 28320 4040 28380 4100
rect 28580 4090 28640 4100
rect 28580 4050 28590 4090
rect 28590 4050 28630 4090
rect 28630 4050 28640 4090
rect 28580 4040 28640 4050
rect 29300 4090 29360 4100
rect 29300 4050 29310 4090
rect 29310 4050 29350 4090
rect 29350 4050 29360 4090
rect 29300 4040 29360 4050
rect 30020 4090 30080 4100
rect 30020 4050 30030 4090
rect 30030 4050 30070 4090
rect 30070 4050 30080 4090
rect 30020 4040 30080 4050
rect 30740 4090 30800 4100
rect 30740 4050 30750 4090
rect 30750 4050 30790 4090
rect 30790 4050 30800 4090
rect 30740 4040 30800 4050
rect 25780 3750 25840 3760
rect 25780 3710 25790 3750
rect 25790 3710 25830 3750
rect 25830 3710 25840 3750
rect 25780 3700 25840 3710
rect 26500 3750 26560 3760
rect 26500 3710 26510 3750
rect 26510 3710 26550 3750
rect 26550 3710 26560 3750
rect 26500 3700 26560 3710
rect 27220 3750 27280 3760
rect 27220 3710 27230 3750
rect 27230 3710 27270 3750
rect 27270 3710 27280 3750
rect 27220 3700 27280 3710
rect 25600 3580 25660 3640
rect 26020 3580 26080 3640
rect 26260 3580 26320 3640
rect 26740 3580 26800 3640
rect 26980 3580 27040 3640
rect 26400 3430 26460 3440
rect 26400 3390 26410 3430
rect 26410 3390 26450 3430
rect 26450 3390 26460 3430
rect 26400 3380 26460 3390
rect 26520 3410 26580 3470
rect 27000 3410 27060 3470
rect 27460 3580 27520 3640
rect 27640 3580 27700 3640
rect 27480 3410 27540 3470
rect 26280 3340 26340 3350
rect 26280 3300 26290 3340
rect 26290 3300 26330 3340
rect 26330 3300 26340 3340
rect 26280 3290 26340 3300
rect 26760 3340 26820 3350
rect 26760 3300 26770 3340
rect 26770 3300 26810 3340
rect 26810 3300 26820 3340
rect 26760 3290 26820 3300
rect 27240 3340 27300 3350
rect 27240 3300 27250 3340
rect 27250 3300 27290 3340
rect 27290 3300 27300 3340
rect 27240 3290 27300 3300
rect 26280 3100 26340 3110
rect 26280 3060 26290 3100
rect 26290 3060 26330 3100
rect 26330 3060 26340 3100
rect 26280 3050 26340 3060
rect 25800 2930 25860 2990
rect 26400 2930 26460 2990
rect 26640 2930 26700 2990
rect 26880 2930 26940 2990
rect 27120 2930 27180 2990
rect 27360 2980 27420 2990
rect 27360 2940 27370 2980
rect 27370 2940 27410 2980
rect 27410 2940 27420 2980
rect 27360 2930 27420 2940
rect 25980 2780 26040 2790
rect 25980 2740 25990 2780
rect 25990 2740 26030 2780
rect 26030 2740 26040 2780
rect 25980 2730 26040 2740
rect 26220 2780 26280 2790
rect 26220 2740 26230 2780
rect 26230 2740 26270 2780
rect 26270 2740 26280 2780
rect 26220 2730 26280 2740
rect 26460 2780 26520 2790
rect 26460 2740 26470 2780
rect 26470 2740 26510 2780
rect 26510 2740 26520 2780
rect 26460 2730 26520 2740
rect 26700 2780 26760 2790
rect 26700 2740 26710 2780
rect 26710 2740 26750 2780
rect 26750 2740 26760 2780
rect 26700 2730 26760 2740
rect 27180 2780 27240 2790
rect 27180 2740 27190 2780
rect 27190 2740 27230 2780
rect 27230 2740 27240 2780
rect 27180 2730 27240 2740
rect 27420 2780 27480 2790
rect 27420 2740 27430 2780
rect 27430 2740 27470 2780
rect 27470 2740 27480 2780
rect 27420 2730 27480 2740
rect 27660 2780 27720 2790
rect 27660 2740 27670 2780
rect 27670 2740 27710 2780
rect 27710 2740 27720 2780
rect 27660 2730 27720 2740
rect 29060 3750 29120 3760
rect 29060 3710 29070 3750
rect 29070 3710 29110 3750
rect 29110 3710 29120 3750
rect 29060 3700 29120 3710
rect 29780 3750 29840 3760
rect 29780 3710 29790 3750
rect 29790 3710 29830 3750
rect 29830 3710 29840 3750
rect 29780 3700 29840 3710
rect 30500 3750 30560 3760
rect 30500 3710 30510 3750
rect 30510 3710 30550 3750
rect 30550 3710 30560 3750
rect 30500 3700 30560 3710
rect 28640 3580 28700 3640
rect 28820 3580 28880 3640
rect 28800 3410 28860 3470
rect 29300 3580 29360 3640
rect 29540 3580 29600 3640
rect 30020 3580 30080 3640
rect 30260 3580 30320 3640
rect 30680 3580 30740 3640
rect 29280 3410 29340 3470
rect 29760 3410 29820 3470
rect 29880 3430 29940 3440
rect 29880 3390 29890 3430
rect 29890 3390 29930 3430
rect 29930 3390 29940 3430
rect 29880 3380 29940 3390
rect 31070 3380 31130 3440
rect 29040 3340 29100 3350
rect 29040 3300 29050 3340
rect 29050 3300 29090 3340
rect 29090 3300 29100 3340
rect 29040 3290 29100 3300
rect 29520 3340 29580 3350
rect 29520 3300 29530 3340
rect 29530 3300 29570 3340
rect 29570 3300 29580 3340
rect 29520 3290 29580 3300
rect 30000 3340 30060 3350
rect 30000 3300 30010 3340
rect 30010 3300 30050 3340
rect 30050 3300 30060 3340
rect 30000 3290 30060 3300
rect 31250 3580 31310 3640
rect 30000 3100 30060 3110
rect 30000 3060 30010 3100
rect 30010 3060 30050 3100
rect 30050 3060 30060 3100
rect 30000 3050 30060 3060
rect 31160 3050 31220 3110
rect 28920 2930 28980 2990
rect 29160 2930 29220 2990
rect 29400 2930 29460 2990
rect 29640 2930 29700 2990
rect 29880 2930 29940 2990
rect 30480 2930 30540 2990
rect 28620 2780 28680 2790
rect 28620 2740 28630 2780
rect 28630 2740 28670 2780
rect 28670 2740 28680 2780
rect 28620 2730 28680 2740
rect 28860 2780 28920 2790
rect 28860 2740 28870 2780
rect 28870 2740 28910 2780
rect 28910 2740 28920 2780
rect 28860 2730 28920 2740
rect 29100 2780 29160 2790
rect 29100 2740 29110 2780
rect 29110 2740 29150 2780
rect 29150 2740 29160 2780
rect 29100 2730 29160 2740
rect 29580 2780 29640 2790
rect 29580 2740 29590 2780
rect 29590 2740 29630 2780
rect 29630 2740 29640 2780
rect 29580 2730 29640 2740
rect 29820 2780 29880 2790
rect 29820 2740 29830 2780
rect 29830 2740 29870 2780
rect 29870 2740 29880 2780
rect 29820 2730 29880 2740
rect 30060 2780 30120 2790
rect 30060 2740 30070 2780
rect 30070 2740 30110 2780
rect 30110 2740 30120 2780
rect 30060 2730 30120 2740
rect 30300 2780 30360 2790
rect 30300 2740 30310 2780
rect 30310 2740 30350 2780
rect 30350 2740 30360 2780
rect 30300 2730 30360 2740
rect 26880 2150 26940 2160
rect 26880 2110 26890 2150
rect 26890 2110 26930 2150
rect 26930 2110 26940 2150
rect 26880 2100 26940 2110
rect 29400 2150 29460 2160
rect 29400 2110 29410 2150
rect 29410 2110 29450 2150
rect 29450 2110 29460 2150
rect 29400 2100 29460 2110
rect 26060 1800 26120 1810
rect 26060 1760 26070 1800
rect 26070 1760 26110 1800
rect 26110 1760 26120 1800
rect 26060 1750 26120 1760
rect 26220 1800 26280 1810
rect 26220 1760 26230 1800
rect 26230 1760 26270 1800
rect 26270 1760 26280 1800
rect 26220 1750 26280 1760
rect 26380 1800 26440 1810
rect 26380 1760 26390 1800
rect 26390 1760 26430 1800
rect 26430 1760 26440 1800
rect 26380 1750 26440 1760
rect 26540 1800 26600 1810
rect 26540 1760 26550 1800
rect 26550 1760 26590 1800
rect 26590 1760 26600 1800
rect 26540 1750 26600 1760
rect 26700 1800 26760 1810
rect 26700 1760 26710 1800
rect 26710 1760 26750 1800
rect 26750 1760 26760 1800
rect 26700 1750 26760 1760
rect 26860 1800 26920 1810
rect 26860 1760 26870 1800
rect 26870 1760 26910 1800
rect 26910 1760 26920 1800
rect 26860 1750 26920 1760
rect 27020 1800 27080 1810
rect 27020 1760 27030 1800
rect 27030 1760 27070 1800
rect 27070 1760 27080 1800
rect 27020 1750 27080 1760
rect 27180 1800 27240 1810
rect 27180 1760 27190 1800
rect 27190 1760 27230 1800
rect 27230 1760 27240 1800
rect 27180 1750 27240 1760
rect 27340 1800 27400 1810
rect 27340 1760 27350 1800
rect 27350 1760 27390 1800
rect 27390 1760 27400 1800
rect 27340 1750 27400 1760
rect 27500 1800 27560 1810
rect 27500 1760 27510 1800
rect 27510 1760 27550 1800
rect 27550 1760 27560 1800
rect 27500 1750 27560 1760
rect 27660 1800 27720 1810
rect 27660 1760 27670 1800
rect 27670 1760 27710 1800
rect 27710 1760 27720 1800
rect 27660 1750 27720 1760
rect 27820 1800 27880 1810
rect 27820 1760 27830 1800
rect 27830 1760 27870 1800
rect 27870 1760 27880 1800
rect 27820 1750 27880 1760
rect 27980 1800 28040 1810
rect 27980 1760 27990 1800
rect 27990 1760 28030 1800
rect 28030 1760 28040 1800
rect 27980 1750 28040 1760
rect 28140 1800 28200 1810
rect 28140 1760 28150 1800
rect 28150 1760 28190 1800
rect 28190 1760 28200 1800
rect 28140 1750 28200 1760
rect 28300 1800 28360 1810
rect 28300 1760 28310 1800
rect 28310 1760 28350 1800
rect 28350 1760 28360 1800
rect 28300 1750 28360 1760
rect 28460 1800 28520 1810
rect 28460 1760 28470 1800
rect 28470 1760 28510 1800
rect 28510 1760 28520 1800
rect 28460 1750 28520 1760
rect 28620 1800 28680 1810
rect 28620 1760 28630 1800
rect 28630 1760 28670 1800
rect 28670 1760 28680 1800
rect 28620 1750 28680 1760
rect 28780 1800 28840 1810
rect 28780 1760 28790 1800
rect 28790 1760 28830 1800
rect 28830 1760 28840 1800
rect 28780 1750 28840 1760
rect 28940 1800 29000 1810
rect 28940 1760 28950 1800
rect 28950 1760 28990 1800
rect 28990 1760 29000 1800
rect 28940 1750 29000 1760
rect 29100 1800 29160 1810
rect 29100 1760 29110 1800
rect 29110 1760 29150 1800
rect 29150 1760 29160 1800
rect 29100 1750 29160 1760
rect 29260 1800 29320 1810
rect 29260 1760 29270 1800
rect 29270 1760 29310 1800
rect 29310 1760 29320 1800
rect 29260 1750 29320 1760
rect 29420 1800 29480 1810
rect 29420 1760 29430 1800
rect 29430 1760 29470 1800
rect 29470 1760 29480 1800
rect 29420 1750 29480 1760
rect 29580 1800 29640 1810
rect 29580 1760 29590 1800
rect 29590 1760 29630 1800
rect 29630 1760 29640 1800
rect 29580 1750 29640 1760
rect 29740 1800 29800 1810
rect 29740 1760 29750 1800
rect 29750 1760 29790 1800
rect 29790 1760 29800 1800
rect 29740 1750 29800 1760
rect 29900 1800 29960 1810
rect 29900 1760 29910 1800
rect 29910 1760 29950 1800
rect 29950 1760 29960 1800
rect 29900 1750 29960 1760
rect 30060 1800 30120 1810
rect 30060 1760 30070 1800
rect 30070 1760 30110 1800
rect 30110 1760 30120 1800
rect 30060 1750 30120 1760
rect 25160 1580 25220 1640
rect 25980 1630 26040 1640
rect 25980 1590 25990 1630
rect 25990 1590 26030 1630
rect 26030 1590 26040 1630
rect 25980 1580 26040 1590
rect 30380 1630 30440 1640
rect 30380 1590 30390 1630
rect 30390 1590 30430 1630
rect 30430 1590 30440 1630
rect 30380 1580 30440 1590
rect 25760 1250 25820 1260
rect 25760 1210 25770 1250
rect 25770 1210 25810 1250
rect 25810 1210 25820 1250
rect 25760 1200 25820 1210
rect 26120 1250 26180 1260
rect 26120 1210 26130 1250
rect 26130 1210 26170 1250
rect 26170 1210 26180 1250
rect 26120 1200 26180 1210
rect 26480 1250 26540 1260
rect 26480 1210 26490 1250
rect 26490 1210 26530 1250
rect 26530 1210 26540 1250
rect 26480 1200 26540 1210
rect 27600 1250 27660 1260
rect 27600 1210 27610 1250
rect 27610 1210 27650 1250
rect 27650 1210 27660 1250
rect 27600 1200 27660 1210
rect 27960 1250 28020 1260
rect 27960 1210 27970 1250
rect 27970 1210 28010 1250
rect 28010 1210 28020 1250
rect 27960 1200 28020 1210
rect 28320 1250 28380 1260
rect 28320 1210 28330 1250
rect 28330 1210 28370 1250
rect 28370 1210 28380 1250
rect 28320 1200 28380 1210
rect 28680 1250 28740 1260
rect 28680 1210 28690 1250
rect 28690 1210 28730 1250
rect 28730 1210 28740 1250
rect 28680 1200 28740 1210
rect 29760 1250 29820 1260
rect 29760 1210 29770 1250
rect 29770 1210 29810 1250
rect 29810 1210 29820 1250
rect 29760 1200 29820 1210
rect 30120 1250 30180 1260
rect 30120 1210 30130 1250
rect 30130 1210 30170 1250
rect 30170 1210 30180 1250
rect 30120 1200 30180 1210
rect 30480 1250 30540 1260
rect 30480 1210 30490 1250
rect 30490 1210 30530 1250
rect 30530 1210 30540 1250
rect 30480 1200 30540 1210
rect 25580 910 25640 920
rect 25580 870 25590 910
rect 25590 870 25630 910
rect 25630 870 25640 910
rect 25580 860 25640 870
rect 26300 910 26360 920
rect 26300 870 26310 910
rect 26310 870 26350 910
rect 26350 870 26360 910
rect 26300 860 26360 870
rect 28140 910 28200 920
rect 28140 870 28150 910
rect 28150 870 28190 910
rect 28190 870 28200 910
rect 28140 860 28200 870
rect 28500 910 28560 920
rect 28500 870 28510 910
rect 28510 870 28550 910
rect 28550 870 28560 910
rect 28500 860 28560 870
rect 28860 910 28920 920
rect 28860 870 28870 910
rect 28870 870 28910 910
rect 28910 870 28920 910
rect 28860 860 28920 870
rect 29580 910 29640 920
rect 29580 870 29590 910
rect 29590 870 29630 910
rect 29630 870 29640 910
rect 29580 860 29640 870
rect 30300 910 30360 920
rect 30300 870 30310 910
rect 30310 870 30350 910
rect 30350 870 30360 910
rect 30300 860 30360 870
rect 25940 750 26000 810
rect 26660 750 26720 810
rect 29940 750 30000 810
rect 30660 750 30720 810
rect 25070 660 25130 720
rect 27420 660 27480 720
<< metal2 >>
rect 19610 9980 19690 9990
rect 19610 9920 19620 9980
rect 19680 9920 19690 9980
rect 19610 9910 19690 9920
rect 31500 9980 31580 9990
rect 31500 9920 31510 9980
rect 31570 9920 31580 9980
rect 31500 9910 31580 9920
rect 19780 7050 19860 7060
rect 19780 6990 19790 7050
rect 19850 7040 19860 7050
rect 22522 7050 22602 7060
rect 22522 7040 22532 7050
rect 19850 7000 22532 7040
rect 19850 6990 19860 7000
rect 19780 6980 19860 6990
rect 22522 6990 22532 7000
rect 22592 6990 22602 7050
rect 22522 6980 22602 6990
rect 28880 6990 28960 7000
rect 28880 6930 28890 6990
rect 28950 6980 28960 6990
rect 31500 6990 31580 7000
rect 31500 6980 31510 6990
rect 28950 6940 31510 6980
rect 28950 6930 28960 6940
rect 28880 6920 28960 6930
rect 31500 6930 31510 6940
rect 31570 6930 31580 6990
rect 31500 6920 31580 6930
rect 19970 6890 20050 6900
rect 19970 6830 19980 6890
rect 20040 6880 20050 6890
rect 21880 6890 21960 6900
rect 21880 6880 21890 6890
rect 20040 6840 21890 6880
rect 20040 6830 20050 6840
rect 19970 6820 20050 6830
rect 21880 6830 21890 6840
rect 21950 6830 21960 6890
rect 21880 6820 21960 6830
rect 23270 6890 23370 6910
rect 24840 6900 24920 6910
rect 24840 6890 24850 6900
rect 23270 6830 23290 6890
rect 23350 6850 24850 6890
rect 23350 6830 23370 6850
rect 24840 6840 24850 6850
rect 24910 6840 24920 6900
rect 24840 6830 24920 6840
rect 30270 6890 30370 6910
rect 30270 6830 30290 6890
rect 30350 6880 30370 6890
rect 30620 6890 30700 6900
rect 30620 6880 30630 6890
rect 30350 6840 30630 6880
rect 30350 6830 30370 6840
rect 23270 6810 23370 6830
rect 30270 6810 30370 6830
rect 30620 6830 30630 6840
rect 30690 6830 30700 6890
rect 30620 6820 30700 6830
rect 19880 6780 19960 6790
rect 19880 6720 19890 6780
rect 19950 6770 19960 6780
rect 25380 6780 25460 6790
rect 25380 6770 25390 6780
rect 19950 6730 25390 6770
rect 19950 6720 19960 6730
rect 19880 6710 19960 6720
rect 25380 6720 25390 6730
rect 25450 6720 25460 6780
rect 25380 6710 25460 6720
rect 22410 6680 22490 6690
rect 22410 6620 22420 6680
rect 22480 6670 22490 6680
rect 25240 6680 25320 6690
rect 25240 6670 25250 6680
rect 22480 6630 25250 6670
rect 22480 6620 22490 6630
rect 22410 6610 22490 6620
rect 25240 6620 25250 6630
rect 25310 6620 25320 6680
rect 25240 6610 25320 6620
rect 26770 6670 26870 6690
rect 26770 6610 26790 6670
rect 26850 6660 26870 6670
rect 31240 6670 31320 6680
rect 31240 6660 31250 6670
rect 26850 6620 31250 6660
rect 26850 6610 26870 6620
rect 26770 6590 26870 6610
rect 31240 6610 31250 6620
rect 31310 6610 31320 6670
rect 31240 6600 31320 6610
rect 22320 6570 22400 6580
rect 22320 6510 22330 6570
rect 22390 6560 22400 6570
rect 25680 6570 25760 6580
rect 25680 6560 25690 6570
rect 22390 6520 25690 6560
rect 22390 6510 22400 6520
rect 22320 6500 22400 6510
rect 25680 6510 25690 6520
rect 25750 6510 25760 6570
rect 25680 6500 25760 6510
rect 25990 6480 26070 6490
rect 25990 6470 26000 6480
rect 20092 6430 26000 6470
rect 20092 6410 20182 6430
rect 25990 6420 26000 6430
rect 26060 6420 26070 6480
rect 25990 6410 26070 6420
rect 20092 6340 20102 6410
rect 20172 6340 20182 6410
rect 22522 6330 22532 6400
rect 22602 6330 22612 6400
rect 25060 6350 25140 6360
rect 25060 6290 25070 6350
rect 25130 6340 25140 6350
rect 26320 6350 26400 6360
rect 26320 6340 26330 6350
rect 25130 6300 26330 6340
rect 25130 6290 25140 6300
rect 19780 6280 19860 6290
rect 19780 6220 19790 6280
rect 19850 6270 19860 6280
rect 20092 6270 20102 6290
rect 19850 6230 20102 6270
rect 19850 6220 19860 6230
rect 20092 6220 20102 6230
rect 20172 6220 20182 6290
rect 25060 6280 25140 6290
rect 26320 6290 26330 6300
rect 26390 6290 26400 6350
rect 26320 6280 26400 6290
rect 26690 6350 26770 6360
rect 26690 6290 26700 6350
rect 26760 6340 26770 6350
rect 27410 6350 27490 6360
rect 27410 6340 27420 6350
rect 26760 6300 27420 6340
rect 26760 6290 26770 6300
rect 26690 6280 26770 6290
rect 27410 6290 27420 6300
rect 27480 6340 27490 6350
rect 28490 6350 28570 6360
rect 28490 6340 28500 6350
rect 27480 6300 28500 6340
rect 27480 6290 27490 6300
rect 27410 6280 27490 6290
rect 28490 6290 28500 6300
rect 28560 6340 28570 6350
rect 29210 6350 29290 6360
rect 29210 6340 29220 6350
rect 28560 6300 29220 6340
rect 28560 6290 28570 6300
rect 28490 6280 28570 6290
rect 29210 6290 29220 6300
rect 29280 6340 29290 6350
rect 29280 6300 30470 6340
rect 29280 6290 29290 6300
rect 29210 6280 29290 6290
rect 19780 6210 19860 6220
rect 22522 6210 22532 6280
rect 22602 6210 22612 6280
rect 22320 6200 22400 6210
rect 22320 6190 22330 6200
rect 20092 6150 22330 6190
rect 20092 6130 20182 6150
rect 22320 6140 22330 6150
rect 22390 6140 22400 6200
rect 22320 6130 22400 6140
rect 20092 6060 20102 6130
rect 20172 6060 20182 6130
rect 31090 6110 32600 6150
rect 31090 6020 32600 6060
rect 26150 6010 26230 6020
rect 19780 6000 19860 6010
rect 19780 5940 19790 6000
rect 19850 5990 19860 6000
rect 20092 5990 20102 6010
rect 19850 5950 20102 5990
rect 19850 5940 19860 5950
rect 20092 5940 20102 5950
rect 20172 5940 20182 6010
rect 26150 5950 26160 6010
rect 26220 6000 26230 6010
rect 26510 6010 26590 6020
rect 26510 6000 26520 6010
rect 26220 5960 26520 6000
rect 26220 5950 26230 5960
rect 26150 5940 26230 5950
rect 26510 5950 26520 5960
rect 26580 6000 26590 6010
rect 26870 6010 26950 6020
rect 26870 6000 26880 6010
rect 26580 5960 26880 6000
rect 26580 5950 26590 5960
rect 26510 5940 26590 5950
rect 26870 5950 26880 5960
rect 26940 6000 26950 6010
rect 27230 6010 27310 6020
rect 27230 6000 27240 6010
rect 26940 5960 27240 6000
rect 26940 5950 26950 5960
rect 26870 5940 26950 5950
rect 27230 5950 27240 5960
rect 27300 6000 27310 6010
rect 27590 6010 27670 6020
rect 27590 6000 27600 6010
rect 27300 5960 27600 6000
rect 27300 5950 27310 5960
rect 27230 5940 27310 5950
rect 27590 5950 27600 5960
rect 27660 6000 27670 6010
rect 27950 6010 28030 6020
rect 27950 6000 27960 6010
rect 27660 5960 27960 6000
rect 27660 5950 27670 5960
rect 27590 5940 27670 5950
rect 27950 5950 27960 5960
rect 28020 6000 28030 6010
rect 28310 6010 28390 6020
rect 28310 6000 28320 6010
rect 28020 5960 28320 6000
rect 28020 5950 28030 5960
rect 27950 5940 28030 5950
rect 28310 5950 28320 5960
rect 28380 6000 28390 6010
rect 28670 6010 28750 6020
rect 28670 6000 28680 6010
rect 28380 5960 28680 6000
rect 28380 5950 28390 5960
rect 28310 5940 28390 5950
rect 28670 5950 28680 5960
rect 28740 6000 28750 6010
rect 29030 6010 29110 6020
rect 29030 6000 29040 6010
rect 28740 5960 29040 6000
rect 28740 5950 28750 5960
rect 28670 5940 28750 5950
rect 29030 5950 29040 5960
rect 29100 6000 29110 6010
rect 29390 6010 29470 6020
rect 29390 6000 29400 6010
rect 29100 5960 29400 6000
rect 29100 5950 29110 5960
rect 29030 5940 29110 5950
rect 29390 5950 29400 5960
rect 29460 6000 29470 6010
rect 29750 6010 29830 6020
rect 29750 6000 29760 6010
rect 29460 5960 29760 6000
rect 29460 5950 29470 5960
rect 29390 5940 29470 5950
rect 29750 5950 29760 5960
rect 29820 6000 29830 6010
rect 30110 6010 30190 6020
rect 30110 6000 30120 6010
rect 29820 5960 30120 6000
rect 29820 5950 29830 5960
rect 29750 5940 29830 5950
rect 30110 5950 30120 5960
rect 30180 6000 30190 6010
rect 30180 5960 30470 6000
rect 30180 5950 30190 5960
rect 30110 5940 30190 5950
rect 19780 5930 19860 5940
rect 24660 5850 24670 5920
rect 24740 5900 24750 5920
rect 24930 5910 25010 5920
rect 31090 5910 32600 5950
rect 24930 5900 24940 5910
rect 24740 5860 24940 5900
rect 24740 5850 24750 5860
rect 24930 5850 24940 5860
rect 25000 5850 25010 5910
rect 24930 5840 25010 5850
rect 29880 5890 29960 5900
rect 19780 5820 19860 5830
rect 19780 5760 19790 5820
rect 19850 5810 19860 5820
rect 21810 5820 22250 5840
rect 29880 5830 29890 5890
rect 29950 5880 29960 5890
rect 30010 5890 30090 5900
rect 30010 5880 30020 5890
rect 29950 5840 30020 5880
rect 29950 5830 29960 5840
rect 29880 5820 29960 5830
rect 30010 5830 30020 5840
rect 30080 5830 30090 5890
rect 30010 5820 30090 5830
rect 21810 5810 21840 5820
rect 19850 5770 21840 5810
rect 19850 5760 19860 5770
rect 19780 5750 19860 5760
rect 21810 5760 21840 5770
rect 21900 5760 22000 5820
rect 22060 5760 22160 5820
rect 22220 5760 22250 5820
rect 21810 5740 22250 5760
rect 24660 5800 24750 5810
rect 24660 5730 24670 5800
rect 24740 5730 24750 5800
rect 25680 5800 25760 5810
rect 25680 5740 25690 5800
rect 25750 5790 25760 5800
rect 31150 5800 31230 5810
rect 31150 5790 31160 5800
rect 25750 5750 31160 5790
rect 25750 5740 25760 5750
rect 25680 5730 25760 5740
rect 31150 5740 31160 5750
rect 31220 5740 31230 5800
rect 31150 5730 31230 5740
rect 24660 5720 24750 5730
rect 19880 5690 19960 5700
rect 19880 5630 19890 5690
rect 19950 5680 19960 5690
rect 20102 5680 20112 5690
rect 19950 5640 20112 5680
rect 19950 5630 19960 5640
rect 19880 5620 19960 5630
rect 20102 5620 20112 5640
rect 20182 5620 20192 5690
rect 21448 5620 21458 5690
rect 21528 5670 21538 5690
rect 22410 5680 22490 5690
rect 22410 5670 22420 5680
rect 21528 5630 22420 5670
rect 21528 5620 21538 5630
rect 22410 5620 22420 5630
rect 22480 5620 22490 5680
rect 22410 5610 22490 5620
rect 22522 5610 22532 5680
rect 22602 5610 22612 5680
rect 23920 5610 23930 5680
rect 24000 5660 24010 5680
rect 24660 5670 24740 5680
rect 24660 5660 24670 5670
rect 24000 5620 24670 5660
rect 24000 5610 24010 5620
rect 24660 5610 24670 5620
rect 24730 5610 24740 5670
rect 31500 5620 31580 5630
rect 31500 5610 31510 5620
rect 24660 5600 24740 5610
rect 19970 5570 20050 5580
rect 31310 5570 31510 5610
rect 19970 5510 19980 5570
rect 20040 5550 20050 5570
rect 20102 5550 20112 5570
rect 20040 5510 20112 5550
rect 19970 5500 20050 5510
rect 20102 5500 20112 5510
rect 20182 5500 20192 5570
rect 21448 5500 21458 5570
rect 21528 5550 21538 5570
rect 24750 5560 24830 5570
rect 24750 5550 24760 5560
rect 21528 5510 24760 5550
rect 21528 5500 21538 5510
rect 24750 5500 24760 5510
rect 24820 5500 24830 5560
rect 31500 5560 31510 5570
rect 31570 5560 31580 5620
rect 31500 5550 31580 5560
rect 24750 5490 24830 5500
rect 26870 5430 26950 5440
rect 26870 5370 26880 5430
rect 26940 5420 26950 5430
rect 27230 5430 27310 5440
rect 27230 5420 27240 5430
rect 26940 5380 27240 5420
rect 26940 5370 26950 5380
rect 26870 5360 26950 5370
rect 27230 5370 27240 5380
rect 27300 5420 27310 5430
rect 27590 5430 27670 5440
rect 27590 5420 27600 5430
rect 27300 5380 27600 5420
rect 27300 5370 27310 5380
rect 27230 5360 27310 5370
rect 27590 5370 27600 5380
rect 27660 5420 27670 5430
rect 27950 5430 28030 5440
rect 27950 5420 27960 5430
rect 27660 5380 27960 5420
rect 27660 5370 27670 5380
rect 27590 5360 27670 5370
rect 27950 5370 27960 5380
rect 28020 5420 28030 5430
rect 28310 5430 28390 5440
rect 28310 5420 28320 5430
rect 28020 5380 28320 5420
rect 28020 5370 28030 5380
rect 27950 5360 28030 5370
rect 28310 5370 28320 5380
rect 28380 5420 28390 5430
rect 28670 5430 28750 5440
rect 28670 5420 28680 5430
rect 28380 5380 28680 5420
rect 28380 5370 28390 5380
rect 28310 5360 28390 5370
rect 28670 5370 28680 5380
rect 28740 5420 28750 5430
rect 29030 5430 29110 5440
rect 29030 5420 29040 5430
rect 28740 5380 29040 5420
rect 28740 5370 28750 5380
rect 28670 5360 28750 5370
rect 29030 5370 29040 5380
rect 29100 5420 29110 5430
rect 29390 5430 29470 5440
rect 29390 5420 29400 5430
rect 29100 5380 29400 5420
rect 29100 5370 29110 5380
rect 29030 5360 29110 5370
rect 29390 5370 29400 5380
rect 29460 5370 29470 5430
rect 29390 5360 29470 5370
rect 22522 5090 22602 5100
rect 22522 5030 22532 5090
rect 22592 5080 22602 5090
rect 24300 5090 24380 5100
rect 24300 5080 24310 5090
rect 22592 5040 24310 5080
rect 22592 5030 22602 5040
rect 22522 5020 22602 5030
rect 24300 5030 24310 5040
rect 24370 5030 24380 5090
rect 24300 5020 24380 5030
rect 25490 4860 25570 4870
rect 25490 4800 25500 4860
rect 25560 4850 25570 4860
rect 25750 4860 25830 4870
rect 25750 4850 25760 4860
rect 25560 4810 25760 4850
rect 25560 4800 25570 4810
rect 25490 4790 25570 4800
rect 25750 4800 25760 4810
rect 25820 4800 25830 4860
rect 25750 4790 25830 4800
rect 24660 4690 24740 4700
rect 24660 4630 24670 4690
rect 24730 4680 24740 4690
rect 27770 4690 27850 4700
rect 27770 4680 27780 4690
rect 24730 4640 27780 4680
rect 24730 4630 24740 4640
rect 24660 4620 24740 4630
rect 27770 4630 27780 4640
rect 27840 4680 27850 4690
rect 28490 4690 28570 4700
rect 28490 4680 28500 4690
rect 27840 4640 28500 4680
rect 27840 4630 27850 4640
rect 27770 4620 27850 4630
rect 28490 4630 28500 4640
rect 28560 4630 28570 4690
rect 28490 4620 28570 4630
rect 24390 4580 24470 4590
rect 24390 4520 24400 4580
rect 24460 4570 24470 4580
rect 24930 4580 25010 4590
rect 24930 4570 24940 4580
rect 24460 4530 24530 4570
rect 24570 4530 24940 4570
rect 24460 4520 24470 4530
rect 24390 4510 24470 4520
rect 24930 4520 24940 4530
rect 25000 4570 25010 4580
rect 25490 4580 25570 4590
rect 25490 4570 25500 4580
rect 25000 4530 25500 4570
rect 25000 4520 25010 4530
rect 24930 4510 25010 4520
rect 25490 4520 25500 4530
rect 25560 4570 25570 4580
rect 27410 4580 27490 4590
rect 27410 4570 27420 4580
rect 25560 4530 27420 4570
rect 25560 4520 25570 4530
rect 25490 4510 25570 4520
rect 27410 4520 27420 4530
rect 27480 4570 27490 4580
rect 28850 4580 28930 4590
rect 28850 4570 28860 4580
rect 27480 4530 28860 4570
rect 27480 4520 27490 4530
rect 27410 4510 27490 4520
rect 28850 4520 28860 4530
rect 28920 4520 28930 4580
rect 28850 4510 28930 4520
rect 25150 4490 25230 4500
rect 25150 4430 25160 4490
rect 25220 4480 25230 4490
rect 25620 4490 25700 4500
rect 25620 4480 25630 4490
rect 25220 4440 25630 4480
rect 25220 4430 25230 4440
rect 25150 4420 25230 4430
rect 25620 4430 25630 4440
rect 25690 4480 25700 4490
rect 27050 4490 27130 4500
rect 27050 4480 27060 4490
rect 25690 4440 27060 4480
rect 25690 4430 25700 4440
rect 25620 4420 25700 4430
rect 27050 4430 27060 4440
rect 27120 4480 27130 4490
rect 29210 4490 29290 4500
rect 29210 4480 29220 4490
rect 27120 4440 29220 4480
rect 27120 4430 27130 4440
rect 27050 4420 27130 4430
rect 29210 4430 29220 4440
rect 29280 4430 29290 4490
rect 29210 4420 29290 4430
rect 29390 4490 29470 4500
rect 29390 4430 29400 4490
rect 29460 4480 29470 4490
rect 30620 4490 30700 4500
rect 30620 4480 30630 4490
rect 29460 4440 30630 4480
rect 29460 4430 29470 4440
rect 29390 4420 29470 4430
rect 30620 4430 30630 4440
rect 30690 4430 30700 4490
rect 30620 4420 30700 4430
rect 25990 4400 26070 4410
rect 25990 4340 26000 4400
rect 26060 4390 26070 4400
rect 26690 4400 26770 4410
rect 26690 4390 26700 4400
rect 26060 4350 26700 4390
rect 26060 4340 26070 4350
rect 25240 4330 25320 4340
rect 25990 4330 26070 4340
rect 26690 4340 26700 4350
rect 26760 4390 26770 4400
rect 28130 4400 28210 4410
rect 28130 4390 28140 4400
rect 26760 4350 28140 4390
rect 26760 4340 26770 4350
rect 26690 4330 26770 4340
rect 28130 4340 28140 4350
rect 28200 4390 28210 4400
rect 29570 4400 29650 4410
rect 29570 4390 29580 4400
rect 28200 4350 29580 4390
rect 28200 4340 28210 4350
rect 28130 4330 28210 4340
rect 29570 4340 29580 4350
rect 29640 4390 29650 4400
rect 31060 4400 31140 4410
rect 31060 4390 31070 4400
rect 29640 4350 31070 4390
rect 29640 4340 29650 4350
rect 29570 4330 29650 4340
rect 31060 4340 31070 4350
rect 31130 4340 31140 4400
rect 31060 4330 31140 4340
rect 25240 4270 25250 4330
rect 25310 4300 25320 4330
rect 28570 4310 28650 4320
rect 28570 4300 28580 4310
rect 25310 4270 28580 4300
rect 25240 4260 28580 4270
rect 28570 4250 28580 4260
rect 28640 4300 28650 4310
rect 30010 4310 30090 4320
rect 30010 4300 30020 4310
rect 28640 4260 30020 4300
rect 28640 4250 28650 4260
rect 28570 4240 28650 4250
rect 30010 4250 30020 4260
rect 30080 4250 30090 4310
rect 30010 4240 30090 4250
rect 25410 4220 25490 4230
rect 25410 4160 25420 4220
rect 25480 4210 25490 4220
rect 25650 4220 25730 4230
rect 25650 4210 25660 4220
rect 25480 4170 25660 4210
rect 25480 4160 25490 4170
rect 25410 4150 25490 4160
rect 25650 4160 25660 4170
rect 25720 4210 25730 4220
rect 25890 4220 25970 4230
rect 25890 4210 25900 4220
rect 25720 4170 25900 4210
rect 25720 4160 25730 4170
rect 25650 4150 25730 4160
rect 25890 4160 25900 4170
rect 25960 4210 25970 4220
rect 26130 4220 26210 4230
rect 26130 4210 26140 4220
rect 25960 4170 26140 4210
rect 25960 4160 25970 4170
rect 25890 4150 25970 4160
rect 26130 4160 26140 4170
rect 26200 4210 26210 4220
rect 26370 4220 26450 4230
rect 26370 4210 26380 4220
rect 26200 4170 26380 4210
rect 26200 4160 26210 4170
rect 26130 4150 26210 4160
rect 26370 4160 26380 4170
rect 26440 4210 26450 4220
rect 26610 4220 26690 4230
rect 26610 4210 26620 4220
rect 26440 4170 26620 4210
rect 26440 4160 26450 4170
rect 26370 4150 26450 4160
rect 26610 4160 26620 4170
rect 26680 4210 26690 4220
rect 26850 4220 26930 4230
rect 26850 4210 26860 4220
rect 26680 4170 26860 4210
rect 26680 4160 26690 4170
rect 26610 4150 26690 4160
rect 26850 4160 26860 4170
rect 26920 4210 26930 4220
rect 27090 4220 27170 4230
rect 27090 4210 27100 4220
rect 26920 4170 27100 4210
rect 26920 4160 26930 4170
rect 26850 4150 26930 4160
rect 27090 4160 27100 4170
rect 27160 4210 27170 4220
rect 27330 4220 27410 4230
rect 27330 4210 27340 4220
rect 27160 4170 27340 4210
rect 27160 4160 27170 4170
rect 27090 4150 27170 4160
rect 27330 4160 27340 4170
rect 27400 4210 27410 4220
rect 27570 4220 27650 4230
rect 27570 4210 27580 4220
rect 27400 4170 27580 4210
rect 27400 4160 27410 4170
rect 27330 4150 27410 4160
rect 27570 4160 27580 4170
rect 27640 4210 27650 4220
rect 28690 4220 28770 4230
rect 28690 4210 28700 4220
rect 27640 4170 28700 4210
rect 27640 4160 27650 4170
rect 27570 4150 27650 4160
rect 28690 4160 28700 4170
rect 28760 4210 28770 4220
rect 28930 4220 29010 4230
rect 28930 4210 28940 4220
rect 28760 4170 28940 4210
rect 28760 4160 28770 4170
rect 28690 4150 28770 4160
rect 28930 4160 28940 4170
rect 29000 4210 29010 4220
rect 29170 4220 29250 4230
rect 29170 4210 29180 4220
rect 29000 4170 29180 4210
rect 29000 4160 29010 4170
rect 28930 4150 29010 4160
rect 29170 4160 29180 4170
rect 29240 4210 29250 4220
rect 29410 4220 29490 4230
rect 29410 4210 29420 4220
rect 29240 4170 29420 4210
rect 29240 4160 29250 4170
rect 29170 4150 29250 4160
rect 29410 4160 29420 4170
rect 29480 4210 29490 4220
rect 29650 4220 29730 4230
rect 29650 4210 29660 4220
rect 29480 4170 29660 4210
rect 29480 4160 29490 4170
rect 29410 4150 29490 4160
rect 29650 4160 29660 4170
rect 29720 4210 29730 4220
rect 29890 4220 29970 4230
rect 29890 4210 29900 4220
rect 29720 4170 29900 4210
rect 29720 4160 29730 4170
rect 29650 4150 29730 4160
rect 29890 4160 29900 4170
rect 29960 4210 29970 4220
rect 30130 4220 30210 4230
rect 30130 4210 30140 4220
rect 29960 4170 30140 4210
rect 29960 4160 29970 4170
rect 29890 4150 29970 4160
rect 30130 4160 30140 4170
rect 30200 4210 30210 4220
rect 30370 4220 30450 4230
rect 30370 4210 30380 4220
rect 30200 4170 30380 4210
rect 30200 4160 30210 4170
rect 30130 4150 30210 4160
rect 30370 4160 30380 4170
rect 30440 4210 30450 4220
rect 30610 4220 30690 4230
rect 30610 4210 30620 4220
rect 30440 4170 30620 4210
rect 30440 4160 30450 4170
rect 30370 4150 30450 4160
rect 30610 4160 30620 4170
rect 30680 4210 30690 4220
rect 30850 4220 30930 4230
rect 30850 4210 30860 4220
rect 30680 4170 30860 4210
rect 30680 4160 30690 4170
rect 30610 4150 30690 4160
rect 30850 4160 30860 4170
rect 30920 4210 30930 4220
rect 31500 4220 31580 4230
rect 31500 4210 31510 4220
rect 30920 4170 31510 4210
rect 30920 4160 30930 4170
rect 30850 4150 30930 4160
rect 31500 4160 31510 4170
rect 31570 4160 31580 4220
rect 31500 4150 31580 4160
rect 24750 4100 24830 4110
rect 24750 4040 24760 4100
rect 24820 4090 24830 4100
rect 25530 4100 25610 4110
rect 25530 4090 25540 4100
rect 24820 4050 25540 4090
rect 24820 4040 24830 4050
rect 24750 4030 24830 4040
rect 25530 4040 25540 4050
rect 25600 4090 25610 4100
rect 26250 4100 26330 4110
rect 26250 4090 26260 4100
rect 25600 4050 26260 4090
rect 25600 4040 25610 4050
rect 25530 4030 25610 4040
rect 26250 4040 26260 4050
rect 26320 4090 26330 4100
rect 26970 4100 27050 4110
rect 26970 4090 26980 4100
rect 26320 4050 26980 4090
rect 26320 4040 26330 4050
rect 26250 4030 26330 4040
rect 26970 4040 26980 4050
rect 27040 4090 27050 4100
rect 27690 4100 27770 4110
rect 27690 4090 27700 4100
rect 27040 4050 27700 4090
rect 27040 4040 27050 4050
rect 26970 4030 27050 4040
rect 27690 4040 27700 4050
rect 27760 4090 27770 4100
rect 27950 4100 28030 4110
rect 27950 4090 27960 4100
rect 27760 4050 27960 4090
rect 27760 4040 27770 4050
rect 27690 4030 27770 4040
rect 27950 4040 27960 4050
rect 28020 4040 28030 4100
rect 27950 4030 28030 4040
rect 28310 4100 28390 4110
rect 28310 4040 28320 4100
rect 28380 4090 28390 4100
rect 28570 4100 28650 4110
rect 28570 4090 28580 4100
rect 28380 4050 28580 4090
rect 28380 4040 28390 4050
rect 28310 4030 28390 4040
rect 28570 4040 28580 4050
rect 28640 4090 28650 4100
rect 29290 4100 29370 4110
rect 29290 4090 29300 4100
rect 28640 4050 29300 4090
rect 28640 4040 28650 4050
rect 28570 4030 28650 4040
rect 29290 4040 29300 4050
rect 29360 4090 29370 4100
rect 30010 4100 30090 4110
rect 30010 4090 30020 4100
rect 29360 4050 30020 4090
rect 29360 4040 29370 4050
rect 29290 4030 29370 4040
rect 30010 4040 30020 4050
rect 30080 4090 30090 4100
rect 30730 4100 30810 4110
rect 30730 4090 30740 4100
rect 30080 4050 30740 4090
rect 30080 4040 30090 4050
rect 30010 4030 30090 4040
rect 30730 4040 30740 4050
rect 30800 4040 30810 4100
rect 30850 4050 30930 4090
rect 30730 4030 30810 4040
rect 25770 3760 25850 3770
rect 25770 3700 25780 3760
rect 25840 3750 25850 3760
rect 26010 3750 26090 3770
rect 26490 3760 26570 3770
rect 26490 3750 26500 3760
rect 25840 3710 26500 3750
rect 25840 3700 25850 3710
rect 25770 3690 25850 3700
rect 26010 3690 26090 3710
rect 26490 3700 26500 3710
rect 26560 3750 26570 3760
rect 26730 3750 26810 3770
rect 27210 3760 27290 3770
rect 27210 3750 27220 3760
rect 26560 3710 27220 3750
rect 26560 3700 26570 3710
rect 26490 3690 26570 3700
rect 26730 3690 26810 3710
rect 27210 3700 27220 3710
rect 27280 3700 27290 3760
rect 27210 3690 27290 3700
rect 27450 3690 27530 3770
rect 28810 3690 28890 3770
rect 29050 3760 29130 3770
rect 29050 3700 29060 3760
rect 29120 3750 29130 3760
rect 29530 3750 29610 3770
rect 29770 3760 29850 3770
rect 29770 3750 29780 3760
rect 29120 3710 29780 3750
rect 29120 3700 29130 3710
rect 29050 3690 29130 3700
rect 29530 3690 29610 3710
rect 29770 3700 29780 3710
rect 29840 3750 29850 3760
rect 30250 3750 30330 3770
rect 30490 3760 30570 3770
rect 30490 3750 30500 3760
rect 29840 3710 30500 3750
rect 29840 3700 29850 3710
rect 29770 3690 29850 3700
rect 30250 3690 30330 3710
rect 30490 3700 30500 3710
rect 30560 3750 30570 3760
rect 30560 3710 30750 3750
rect 30560 3700 30570 3710
rect 30490 3690 30570 3700
rect 24840 3640 24920 3650
rect 24840 3580 24850 3640
rect 24910 3630 24920 3640
rect 25590 3640 25670 3650
rect 25590 3630 25600 3640
rect 24910 3590 25600 3630
rect 24910 3580 24920 3590
rect 24840 3570 24920 3580
rect 25590 3580 25600 3590
rect 25660 3630 25670 3640
rect 26010 3640 26090 3650
rect 26010 3630 26020 3640
rect 25660 3590 26020 3630
rect 25660 3580 25670 3590
rect 25590 3570 25670 3580
rect 26010 3580 26020 3590
rect 26080 3630 26090 3640
rect 26250 3640 26330 3650
rect 26250 3630 26260 3640
rect 26080 3590 26260 3630
rect 26080 3580 26090 3590
rect 26010 3570 26090 3580
rect 26250 3580 26260 3590
rect 26320 3630 26330 3640
rect 26730 3640 26810 3650
rect 26730 3630 26740 3640
rect 26320 3590 26740 3630
rect 26320 3580 26330 3590
rect 26250 3570 26330 3580
rect 26730 3580 26740 3590
rect 26800 3630 26810 3640
rect 26970 3640 27050 3650
rect 26970 3630 26980 3640
rect 26800 3590 26980 3630
rect 26800 3580 26810 3590
rect 26730 3570 26810 3580
rect 26970 3580 26980 3590
rect 27040 3630 27050 3640
rect 27450 3640 27530 3650
rect 27450 3630 27460 3640
rect 27040 3590 27460 3630
rect 27040 3580 27050 3590
rect 26970 3570 27050 3580
rect 27450 3580 27460 3590
rect 27520 3630 27530 3640
rect 27630 3640 27710 3650
rect 27630 3630 27640 3640
rect 27520 3590 27640 3630
rect 27520 3580 27530 3590
rect 27450 3570 27530 3580
rect 27630 3580 27640 3590
rect 27700 3580 27710 3640
rect 27630 3570 27710 3580
rect 28630 3640 28710 3650
rect 28630 3580 28640 3640
rect 28700 3630 28710 3640
rect 28810 3640 28890 3650
rect 28810 3630 28820 3640
rect 28700 3590 28820 3630
rect 28700 3580 28710 3590
rect 28630 3570 28710 3580
rect 28810 3580 28820 3590
rect 28880 3630 28890 3640
rect 29290 3640 29370 3650
rect 29290 3630 29300 3640
rect 28880 3590 29300 3630
rect 28880 3580 28890 3590
rect 28810 3570 28890 3580
rect 29290 3580 29300 3590
rect 29360 3630 29370 3640
rect 29530 3640 29610 3650
rect 29530 3630 29540 3640
rect 29360 3590 29540 3630
rect 29360 3580 29370 3590
rect 29290 3570 29370 3580
rect 29530 3580 29540 3590
rect 29600 3630 29610 3640
rect 30010 3640 30090 3650
rect 30010 3630 30020 3640
rect 29600 3590 30020 3630
rect 29600 3580 29610 3590
rect 29530 3570 29610 3580
rect 30010 3580 30020 3590
rect 30080 3630 30090 3640
rect 30250 3640 30330 3650
rect 30250 3630 30260 3640
rect 30080 3590 30260 3630
rect 30080 3580 30090 3590
rect 30010 3570 30090 3580
rect 30250 3580 30260 3590
rect 30320 3630 30330 3640
rect 30670 3640 30750 3650
rect 30670 3630 30680 3640
rect 30320 3590 30680 3630
rect 30320 3580 30330 3590
rect 30250 3570 30330 3580
rect 30670 3580 30680 3590
rect 30740 3630 30750 3640
rect 31240 3640 31320 3650
rect 31240 3630 31250 3640
rect 30740 3590 31250 3630
rect 30740 3580 30750 3590
rect 30670 3570 30750 3580
rect 31240 3580 31250 3590
rect 31310 3580 31320 3640
rect 31240 3570 31320 3580
rect 26510 3470 26590 3480
rect 26390 3440 26470 3450
rect 26390 3430 26400 3440
rect 26040 3390 26400 3430
rect 26390 3380 26400 3390
rect 26460 3380 26470 3440
rect 26510 3410 26520 3470
rect 26580 3460 26590 3470
rect 26990 3470 27070 3480
rect 26990 3460 27000 3470
rect 26580 3420 27000 3460
rect 26580 3410 26590 3420
rect 26510 3400 26590 3410
rect 26990 3410 27000 3420
rect 27060 3460 27070 3470
rect 27470 3470 27550 3480
rect 27470 3460 27480 3470
rect 27060 3420 27480 3460
rect 27060 3410 27070 3420
rect 26990 3400 27070 3410
rect 27470 3410 27480 3420
rect 27540 3410 27550 3470
rect 27470 3400 27550 3410
rect 28790 3470 28870 3480
rect 28790 3410 28800 3470
rect 28860 3460 28870 3470
rect 29270 3470 29350 3480
rect 29270 3460 29280 3470
rect 28860 3420 29280 3460
rect 28860 3410 28870 3420
rect 28790 3400 28870 3410
rect 29270 3410 29280 3420
rect 29340 3460 29350 3470
rect 29750 3470 29830 3480
rect 29750 3460 29760 3470
rect 29340 3420 29760 3460
rect 29340 3410 29350 3420
rect 29270 3400 29350 3410
rect 29750 3410 29760 3420
rect 29820 3410 29830 3470
rect 29750 3400 29830 3410
rect 29870 3440 29950 3450
rect 26390 3370 26470 3380
rect 29870 3380 29880 3440
rect 29940 3430 29950 3440
rect 31060 3440 31140 3450
rect 31060 3430 31070 3440
rect 29940 3390 31070 3430
rect 29940 3380 29950 3390
rect 29870 3370 29950 3380
rect 31060 3380 31070 3390
rect 31130 3380 31140 3440
rect 31300 3390 32600 3430
rect 31060 3370 31140 3380
rect 26270 3350 26350 3360
rect 26270 3290 26280 3350
rect 26340 3340 26350 3350
rect 26750 3350 26830 3360
rect 26750 3340 26760 3350
rect 26340 3300 26760 3340
rect 26340 3290 26350 3300
rect 26270 3280 26350 3290
rect 26750 3290 26760 3300
rect 26820 3340 26830 3350
rect 27230 3350 27310 3360
rect 27230 3340 27240 3350
rect 26820 3300 27240 3340
rect 26820 3290 26830 3300
rect 26750 3280 26830 3290
rect 27230 3290 27240 3300
rect 27300 3290 27310 3350
rect 27230 3280 27310 3290
rect 29030 3350 29110 3360
rect 29030 3290 29040 3350
rect 29100 3340 29110 3350
rect 29510 3350 29590 3360
rect 29510 3340 29520 3350
rect 29100 3300 29520 3340
rect 29100 3290 29110 3300
rect 29030 3280 29110 3290
rect 29510 3290 29520 3300
rect 29580 3340 29590 3350
rect 29990 3350 30070 3360
rect 29990 3340 30000 3350
rect 29580 3300 30000 3340
rect 29580 3290 29590 3300
rect 29510 3280 29590 3290
rect 29990 3290 30000 3300
rect 30060 3290 30070 3350
rect 29990 3280 30070 3290
rect 26270 3110 26350 3120
rect 26270 3100 26280 3110
rect 26030 3060 26280 3100
rect 26270 3050 26280 3060
rect 26340 3050 26350 3110
rect 19780 3040 19860 3050
rect 19780 2980 19790 3040
rect 19850 2980 19860 3040
rect 19780 2970 19860 2980
rect 19910 3040 19990 3050
rect 26270 3040 26350 3050
rect 29990 3110 30070 3120
rect 29990 3050 30000 3110
rect 30060 3100 30070 3110
rect 31150 3110 31230 3120
rect 31150 3100 31160 3110
rect 30060 3060 31160 3100
rect 30060 3050 30070 3060
rect 29990 3040 30070 3050
rect 31150 3050 31160 3060
rect 31220 3050 31230 3110
rect 31150 3040 31230 3050
rect 19910 2980 19920 3040
rect 19980 2980 19990 3040
rect 19910 2970 19990 2980
rect 22524 3020 22604 3030
rect 22524 2960 22540 3020
rect 22594 3010 22604 3020
rect 24390 3020 24470 3030
rect 24390 3010 24400 3020
rect 22594 2970 24400 3010
rect 22594 2960 22604 2970
rect 22524 2950 22604 2960
rect 24390 2960 24400 2970
rect 24460 2960 24470 3020
rect 24390 2950 24470 2960
rect 25790 2990 25870 3000
rect 25790 2930 25800 2990
rect 25860 2980 25870 2990
rect 26390 2990 26470 3000
rect 26390 2980 26400 2990
rect 25860 2940 26400 2980
rect 25860 2930 25870 2940
rect 25790 2920 25870 2930
rect 26390 2930 26400 2940
rect 26460 2980 26470 2990
rect 26630 2990 26710 3000
rect 26630 2980 26640 2990
rect 26460 2940 26640 2980
rect 26460 2930 26470 2940
rect 26390 2920 26470 2930
rect 26630 2930 26640 2940
rect 26700 2980 26710 2990
rect 26870 2990 26950 3000
rect 26870 2980 26880 2990
rect 26700 2940 26880 2980
rect 26700 2930 26710 2940
rect 26630 2920 26710 2930
rect 26870 2930 26880 2940
rect 26940 2980 26950 2990
rect 27110 2990 27190 3000
rect 27110 2980 27120 2990
rect 26940 2940 27120 2980
rect 26940 2930 26950 2940
rect 26870 2920 26950 2930
rect 27110 2930 27120 2940
rect 27180 2980 27190 2990
rect 27350 2990 27430 3000
rect 27350 2980 27360 2990
rect 27180 2940 27360 2980
rect 27180 2930 27190 2940
rect 27110 2920 27190 2930
rect 27350 2930 27360 2940
rect 27420 2930 27430 2990
rect 27350 2920 27430 2930
rect 28910 2990 28990 3000
rect 28910 2930 28920 2990
rect 28980 2980 28990 2990
rect 29150 2990 29230 3000
rect 29150 2980 29160 2990
rect 28980 2940 29160 2980
rect 28980 2930 28990 2940
rect 28910 2920 28990 2930
rect 29150 2930 29160 2940
rect 29220 2980 29230 2990
rect 29390 2990 29470 3000
rect 29390 2980 29400 2990
rect 29220 2940 29400 2980
rect 29220 2930 29230 2940
rect 29150 2920 29230 2930
rect 29390 2930 29400 2940
rect 29460 2980 29470 2990
rect 29630 2990 29710 3000
rect 29630 2980 29640 2990
rect 29460 2940 29640 2980
rect 29460 2930 29470 2940
rect 29390 2920 29470 2930
rect 29630 2930 29640 2940
rect 29700 2980 29710 2990
rect 29870 2990 29950 3000
rect 29870 2980 29880 2990
rect 29700 2940 29880 2980
rect 29700 2930 29710 2940
rect 29630 2920 29710 2930
rect 29870 2930 29880 2940
rect 29940 2980 29950 2990
rect 30470 2990 30550 3000
rect 30470 2980 30480 2990
rect 29940 2940 30480 2980
rect 29940 2930 29950 2940
rect 29870 2920 29950 2930
rect 30470 2930 30480 2940
rect 30540 2930 30550 2990
rect 30470 2920 30550 2930
rect 25970 2790 26050 2800
rect 25970 2730 25980 2790
rect 26040 2780 26050 2790
rect 26210 2790 26290 2800
rect 26210 2780 26220 2790
rect 26040 2740 26220 2780
rect 26040 2730 26050 2740
rect 25970 2720 26050 2730
rect 26210 2730 26220 2740
rect 26280 2780 26290 2790
rect 26450 2790 26530 2800
rect 26450 2780 26460 2790
rect 26280 2740 26460 2780
rect 26280 2730 26290 2740
rect 26210 2720 26290 2730
rect 26450 2730 26460 2740
rect 26520 2780 26530 2790
rect 26690 2790 26770 2800
rect 26690 2780 26700 2790
rect 26520 2740 26700 2780
rect 26520 2730 26530 2740
rect 26450 2720 26530 2730
rect 26690 2730 26700 2740
rect 26760 2780 26770 2790
rect 27170 2790 27250 2800
rect 27170 2780 27180 2790
rect 26760 2740 27180 2780
rect 26760 2730 26770 2740
rect 26690 2720 26770 2730
rect 27170 2730 27180 2740
rect 27240 2780 27250 2790
rect 27410 2790 27490 2800
rect 27410 2780 27420 2790
rect 27240 2740 27420 2780
rect 27240 2730 27250 2740
rect 27170 2720 27250 2730
rect 27410 2730 27420 2740
rect 27480 2780 27490 2790
rect 27650 2790 27730 2800
rect 27650 2780 27660 2790
rect 27480 2740 27660 2780
rect 27480 2730 27490 2740
rect 27410 2720 27490 2730
rect 27650 2730 27660 2740
rect 27720 2780 27730 2790
rect 28610 2790 28690 2800
rect 28610 2780 28620 2790
rect 27720 2740 28620 2780
rect 27720 2730 27730 2740
rect 27650 2720 27730 2730
rect 28610 2730 28620 2740
rect 28680 2780 28690 2790
rect 28850 2790 28930 2800
rect 28850 2780 28860 2790
rect 28680 2740 28860 2780
rect 28680 2730 28690 2740
rect 28610 2720 28690 2730
rect 28850 2730 28860 2740
rect 28920 2780 28930 2790
rect 29090 2790 29170 2800
rect 29090 2780 29100 2790
rect 28920 2740 29100 2780
rect 28920 2730 28930 2740
rect 28850 2720 28930 2730
rect 29090 2730 29100 2740
rect 29160 2780 29170 2790
rect 29570 2790 29650 2800
rect 29570 2780 29580 2790
rect 29160 2740 29580 2780
rect 29160 2730 29170 2740
rect 29090 2720 29170 2730
rect 29570 2730 29580 2740
rect 29640 2780 29650 2790
rect 29810 2790 29890 2800
rect 29810 2780 29820 2790
rect 29640 2740 29820 2780
rect 29640 2730 29650 2740
rect 29570 2720 29650 2730
rect 29810 2730 29820 2740
rect 29880 2780 29890 2790
rect 30050 2790 30130 2800
rect 30050 2780 30060 2790
rect 29880 2740 30060 2780
rect 29880 2730 29890 2740
rect 29810 2720 29890 2730
rect 30050 2730 30060 2740
rect 30120 2780 30130 2790
rect 30290 2790 30370 2800
rect 30290 2780 30300 2790
rect 30120 2740 30300 2780
rect 30120 2730 30130 2740
rect 30050 2720 30130 2730
rect 30290 2730 30300 2740
rect 30360 2780 30370 2790
rect 31500 2790 31580 2800
rect 31500 2780 31510 2790
rect 30360 2740 31510 2780
rect 30360 2730 30370 2740
rect 30290 2720 30370 2730
rect 31500 2730 31510 2740
rect 31570 2730 31580 2790
rect 31500 2720 31580 2730
rect 26870 2160 26950 2170
rect 26870 2100 26880 2160
rect 26940 2150 26950 2160
rect 29390 2160 29470 2170
rect 29390 2150 29400 2160
rect 26940 2110 29400 2150
rect 26940 2100 26950 2110
rect 26870 2090 26950 2100
rect 29390 2100 29400 2110
rect 29460 2150 29470 2160
rect 31330 2160 31410 2170
rect 31330 2150 31340 2160
rect 29460 2110 31340 2150
rect 29460 2100 29470 2110
rect 29390 2090 29470 2100
rect 31330 2100 31340 2110
rect 31400 2100 31410 2160
rect 31330 2090 31410 2100
rect 26050 1810 26130 1820
rect 26050 1750 26060 1810
rect 26120 1800 26130 1810
rect 26210 1810 26290 1820
rect 26210 1800 26220 1810
rect 26120 1760 26220 1800
rect 26120 1750 26130 1760
rect 26050 1740 26130 1750
rect 26210 1750 26220 1760
rect 26280 1800 26290 1810
rect 26370 1810 26450 1820
rect 26370 1800 26380 1810
rect 26280 1760 26380 1800
rect 26280 1750 26290 1760
rect 26210 1740 26290 1750
rect 26370 1750 26380 1760
rect 26440 1800 26450 1810
rect 26530 1810 26610 1820
rect 26530 1800 26540 1810
rect 26440 1760 26540 1800
rect 26440 1750 26450 1760
rect 26370 1740 26450 1750
rect 26530 1750 26540 1760
rect 26600 1800 26610 1810
rect 26690 1810 26770 1820
rect 26690 1800 26700 1810
rect 26600 1760 26700 1800
rect 26600 1750 26610 1760
rect 26530 1740 26610 1750
rect 26690 1750 26700 1760
rect 26760 1800 26770 1810
rect 26850 1810 26930 1820
rect 26850 1800 26860 1810
rect 26760 1760 26860 1800
rect 26760 1750 26770 1760
rect 26690 1740 26770 1750
rect 26850 1750 26860 1760
rect 26920 1800 26930 1810
rect 27010 1810 27090 1820
rect 27010 1800 27020 1810
rect 26920 1760 27020 1800
rect 26920 1750 26930 1760
rect 26850 1740 26930 1750
rect 27010 1750 27020 1760
rect 27080 1800 27090 1810
rect 27170 1810 27250 1820
rect 27170 1800 27180 1810
rect 27080 1760 27180 1800
rect 27080 1750 27090 1760
rect 27010 1740 27090 1750
rect 27170 1750 27180 1760
rect 27240 1800 27250 1810
rect 27330 1810 27410 1820
rect 27330 1800 27340 1810
rect 27240 1760 27340 1800
rect 27240 1750 27250 1760
rect 27170 1740 27250 1750
rect 27330 1750 27340 1760
rect 27400 1800 27410 1810
rect 27490 1810 27570 1820
rect 27490 1800 27500 1810
rect 27400 1760 27500 1800
rect 27400 1750 27410 1760
rect 27330 1740 27410 1750
rect 27490 1750 27500 1760
rect 27560 1800 27570 1810
rect 27650 1810 27730 1820
rect 27650 1800 27660 1810
rect 27560 1760 27660 1800
rect 27560 1750 27570 1760
rect 27490 1740 27570 1750
rect 27650 1750 27660 1760
rect 27720 1800 27730 1810
rect 27810 1810 27890 1820
rect 27810 1800 27820 1810
rect 27720 1760 27820 1800
rect 27720 1750 27730 1760
rect 27650 1740 27730 1750
rect 27810 1750 27820 1760
rect 27880 1800 27890 1810
rect 27970 1810 28050 1820
rect 27970 1800 27980 1810
rect 27880 1760 27980 1800
rect 27880 1750 27890 1760
rect 27810 1740 27890 1750
rect 27970 1750 27980 1760
rect 28040 1750 28050 1810
rect 27970 1740 28050 1750
rect 28130 1810 28210 1820
rect 28130 1750 28140 1810
rect 28200 1800 28210 1810
rect 28290 1810 28370 1820
rect 28290 1800 28300 1810
rect 28200 1760 28300 1800
rect 28200 1750 28210 1760
rect 28130 1740 28210 1750
rect 28290 1750 28300 1760
rect 28360 1800 28370 1810
rect 28450 1810 28530 1820
rect 28450 1800 28460 1810
rect 28360 1760 28460 1800
rect 28360 1750 28370 1760
rect 28290 1740 28370 1750
rect 28450 1750 28460 1760
rect 28520 1800 28530 1810
rect 28610 1810 28690 1820
rect 28610 1800 28620 1810
rect 28520 1760 28620 1800
rect 28520 1750 28530 1760
rect 28450 1740 28530 1750
rect 28610 1750 28620 1760
rect 28680 1800 28690 1810
rect 28770 1810 28850 1820
rect 28770 1800 28780 1810
rect 28680 1760 28780 1800
rect 28680 1750 28690 1760
rect 28610 1740 28690 1750
rect 28770 1750 28780 1760
rect 28840 1800 28850 1810
rect 28930 1810 29010 1820
rect 28930 1800 28940 1810
rect 28840 1760 28940 1800
rect 28840 1750 28850 1760
rect 28770 1740 28850 1750
rect 28930 1750 28940 1760
rect 29000 1800 29010 1810
rect 29090 1810 29170 1820
rect 29090 1800 29100 1810
rect 29000 1760 29100 1800
rect 29000 1750 29010 1760
rect 28930 1740 29010 1750
rect 29090 1750 29100 1760
rect 29160 1800 29170 1810
rect 29250 1810 29330 1820
rect 29250 1800 29260 1810
rect 29160 1760 29260 1800
rect 29160 1750 29170 1760
rect 29090 1740 29170 1750
rect 29250 1750 29260 1760
rect 29320 1800 29330 1810
rect 29410 1810 29490 1820
rect 29410 1800 29420 1810
rect 29320 1760 29420 1800
rect 29320 1750 29330 1760
rect 29250 1740 29330 1750
rect 29410 1750 29420 1760
rect 29480 1800 29490 1810
rect 29570 1810 29650 1820
rect 29570 1800 29580 1810
rect 29480 1760 29580 1800
rect 29480 1750 29490 1760
rect 29410 1740 29490 1750
rect 29570 1750 29580 1760
rect 29640 1800 29650 1810
rect 29730 1810 29810 1820
rect 29730 1800 29740 1810
rect 29640 1760 29740 1800
rect 29640 1750 29650 1760
rect 29570 1740 29650 1750
rect 29730 1750 29740 1760
rect 29800 1800 29810 1810
rect 29890 1810 29970 1820
rect 29890 1800 29900 1810
rect 29800 1760 29900 1800
rect 29800 1750 29810 1760
rect 29730 1740 29810 1750
rect 29890 1750 29900 1760
rect 29960 1800 29970 1810
rect 30050 1810 30130 1820
rect 30050 1800 30060 1810
rect 29960 1760 30060 1800
rect 29960 1750 29970 1760
rect 29890 1740 29970 1750
rect 30050 1750 30060 1760
rect 30120 1750 30130 1810
rect 30050 1740 30130 1750
rect 25150 1640 25230 1650
rect 25150 1580 25160 1640
rect 25220 1630 25230 1640
rect 25970 1640 26050 1650
rect 25970 1630 25980 1640
rect 25220 1590 25980 1630
rect 25220 1580 25230 1590
rect 25150 1570 25230 1580
rect 25970 1580 25980 1590
rect 26040 1580 26050 1640
rect 25970 1570 26050 1580
rect 30370 1640 30450 1650
rect 30370 1580 30380 1640
rect 30440 1630 30450 1640
rect 31330 1640 31410 1650
rect 31330 1630 31340 1640
rect 30440 1590 31340 1630
rect 30440 1580 30450 1590
rect 30370 1570 30450 1580
rect 31330 1580 31340 1590
rect 31400 1580 31410 1640
rect 31330 1570 31410 1580
rect 25750 1260 25830 1270
rect 25750 1200 25760 1260
rect 25820 1250 25830 1260
rect 26110 1260 26190 1270
rect 26110 1250 26120 1260
rect 25820 1210 26120 1250
rect 25820 1200 25830 1210
rect 25750 1190 25830 1200
rect 26110 1200 26120 1210
rect 26180 1250 26190 1260
rect 26470 1260 26550 1270
rect 26470 1250 26480 1260
rect 26180 1210 26480 1250
rect 26180 1200 26190 1210
rect 26110 1190 26190 1200
rect 26470 1200 26480 1210
rect 26540 1250 26550 1260
rect 27590 1260 27670 1270
rect 27590 1250 27600 1260
rect 26540 1210 27600 1250
rect 26540 1200 26550 1210
rect 26470 1190 26550 1200
rect 27590 1200 27600 1210
rect 27660 1250 27670 1260
rect 27950 1260 28030 1270
rect 27950 1250 27960 1260
rect 27660 1210 27960 1250
rect 27660 1200 27670 1210
rect 27590 1190 27670 1200
rect 27950 1200 27960 1210
rect 28020 1250 28030 1260
rect 28310 1260 28390 1270
rect 28310 1250 28320 1260
rect 28020 1210 28320 1250
rect 28020 1200 28030 1210
rect 27950 1190 28030 1200
rect 28310 1200 28320 1210
rect 28380 1250 28390 1260
rect 28670 1260 28750 1270
rect 28670 1250 28680 1260
rect 28380 1210 28680 1250
rect 28380 1200 28390 1210
rect 28310 1190 28390 1200
rect 28670 1200 28680 1210
rect 28740 1250 28750 1260
rect 29750 1260 29830 1270
rect 29750 1250 29760 1260
rect 28740 1210 29760 1250
rect 28740 1200 28750 1210
rect 28670 1190 28750 1200
rect 29750 1200 29760 1210
rect 29820 1250 29830 1260
rect 30110 1260 30190 1270
rect 30110 1250 30120 1260
rect 29820 1210 30120 1250
rect 29820 1200 29830 1210
rect 29750 1190 29830 1200
rect 30110 1200 30120 1210
rect 30180 1250 30190 1260
rect 30470 1260 30550 1270
rect 30470 1250 30480 1260
rect 30180 1210 30480 1250
rect 30180 1200 30190 1210
rect 30110 1190 30190 1200
rect 30470 1200 30480 1210
rect 30540 1250 30550 1260
rect 31330 1260 31410 1270
rect 31330 1250 31340 1260
rect 30540 1210 31340 1250
rect 30540 1200 30550 1210
rect 31330 1200 31340 1210
rect 31400 1200 31410 1260
rect 30470 1190 30550 1200
rect 25570 920 25650 930
rect 25570 860 25580 920
rect 25640 910 25650 920
rect 26290 920 26370 930
rect 26290 910 26300 920
rect 25640 870 26300 910
rect 25640 860 25650 870
rect 25570 850 25650 860
rect 26290 860 26300 870
rect 26360 860 26370 920
rect 26290 850 26370 860
rect 28130 920 28210 930
rect 28130 860 28140 920
rect 28200 910 28210 920
rect 28490 920 28570 930
rect 28490 910 28500 920
rect 28200 870 28500 910
rect 28200 860 28210 870
rect 28130 850 28210 860
rect 28490 860 28500 870
rect 28560 910 28570 920
rect 28850 920 28930 930
rect 28850 910 28860 920
rect 28560 870 28860 910
rect 28560 860 28570 870
rect 28490 850 28570 860
rect 28850 860 28860 870
rect 28920 860 28930 920
rect 28850 850 28930 860
rect 29570 920 29650 930
rect 29570 860 29580 920
rect 29640 910 29650 920
rect 30290 920 30370 930
rect 30290 910 30300 920
rect 29640 870 30300 910
rect 29640 860 29650 870
rect 29570 850 29650 860
rect 30290 860 30300 870
rect 30360 860 30370 920
rect 30290 850 30370 860
rect 25930 810 26010 820
rect 25930 750 25940 810
rect 26000 800 26010 810
rect 26650 810 26730 820
rect 26650 800 26660 810
rect 26000 760 26660 800
rect 26000 750 26010 760
rect 25930 740 26010 750
rect 26650 750 26660 760
rect 26720 750 26730 810
rect 26650 740 26730 750
rect 29930 810 30010 820
rect 29930 750 29940 810
rect 30000 800 30010 810
rect 30650 810 30730 820
rect 30650 800 30660 810
rect 30000 760 30660 800
rect 30000 750 30010 760
rect 29930 740 30010 750
rect 30650 750 30660 760
rect 30720 750 30730 810
rect 30650 740 30730 750
rect 25060 720 25140 730
rect 25060 660 25070 720
rect 25130 710 25140 720
rect 27410 720 27490 730
rect 27410 710 27420 720
rect 25130 670 27420 710
rect 25130 660 25140 670
rect 25060 650 25140 660
rect 27410 660 27420 670
rect 27480 660 27490 720
rect 27410 650 27490 660
rect 19610 450 19690 460
rect 19610 390 19620 450
rect 19680 390 19690 450
rect 19610 380 19690 390
<< via2 >>
rect 19620 9920 19680 9980
rect 31510 9920 31570 9980
rect 19790 6990 19850 7050
rect 28890 6930 28950 6990
rect 31510 6930 31570 6990
rect 21890 6830 21950 6890
rect 23290 6830 23350 6890
rect 30290 6830 30350 6890
rect 25390 6720 25450 6780
rect 26790 6610 26850 6670
rect 19790 6220 19850 6280
rect 19790 5940 19850 6000
rect 19790 5760 19850 5820
rect 31510 5560 31570 5620
rect 31510 4160 31570 4220
rect 19790 2980 19850 3040
rect 31510 2730 31570 2790
rect 31340 2100 31400 2160
rect 31340 1580 31400 1640
rect 31340 1200 31400 1260
rect 19620 390 19680 450
<< metal3 >>
rect 19600 9990 19700 10000
rect 19600 9910 19610 9990
rect 19690 9910 19700 9990
rect 19600 9900 19700 9910
rect 31490 9990 31590 10000
rect 31490 9910 31500 9990
rect 31580 9910 31590 9990
rect 31490 9900 31590 9910
rect 19610 470 19690 9900
rect 19770 9820 19870 9830
rect 19770 9740 19780 9820
rect 19860 9740 19870 9820
rect 19770 9730 19870 9740
rect 31320 9820 31420 9830
rect 31320 9740 31330 9820
rect 31410 9740 31420 9820
rect 31320 9730 31420 9740
rect 19780 7050 19860 9730
rect 20290 9540 20750 9710
rect 20990 9540 21450 9710
rect 21690 9540 22150 9710
rect 22390 9540 22850 9710
rect 23090 9540 23550 9710
rect 20290 9440 23550 9540
rect 20290 9250 20750 9440
rect 20990 9250 21450 9440
rect 21690 9250 22150 9440
rect 22390 9250 22850 9440
rect 23090 9250 23550 9440
rect 23790 9540 24250 9710
rect 24490 9540 24950 9710
rect 25190 9540 25650 9710
rect 25890 9540 26350 9710
rect 26590 9540 27050 9710
rect 23790 9440 27050 9540
rect 23790 9250 24250 9440
rect 24490 9250 24950 9440
rect 25190 9250 25650 9440
rect 25890 9250 26350 9440
rect 26590 9250 27050 9440
rect 27290 9540 27750 9710
rect 27990 9540 28450 9710
rect 28690 9540 29150 9710
rect 29390 9540 29850 9710
rect 30090 9540 30550 9710
rect 27290 9440 30550 9540
rect 27290 9250 27750 9440
rect 27990 9250 28450 9440
rect 28690 9250 29150 9440
rect 29390 9250 29850 9440
rect 30090 9250 30550 9440
rect 21870 9010 21970 9250
rect 25370 9010 25470 9250
rect 28870 9010 28970 9250
rect 20290 8840 20750 9010
rect 20990 8840 21450 9010
rect 21690 8840 22150 9010
rect 22390 8840 22850 9010
rect 23090 8840 23550 9010
rect 20290 8740 23550 8840
rect 20290 8550 20750 8740
rect 20990 8550 21450 8740
rect 21690 8550 22150 8740
rect 22390 8550 22850 8740
rect 23090 8550 23550 8740
rect 23790 8840 24250 9010
rect 24490 8840 24950 9010
rect 25190 8840 25650 9010
rect 25890 8840 26350 9010
rect 26590 8840 27050 9010
rect 23790 8740 27050 8840
rect 23790 8550 24250 8740
rect 24490 8550 24950 8740
rect 25190 8550 25650 8740
rect 25890 8550 26350 8740
rect 26590 8550 27050 8740
rect 27290 8840 27750 9010
rect 27990 8840 28450 9010
rect 28690 8840 29150 9010
rect 29390 8840 29850 9010
rect 30090 8840 30550 9010
rect 27290 8740 30550 8840
rect 27290 8550 27750 8740
rect 27990 8550 28450 8740
rect 28690 8550 29150 8740
rect 29390 8550 29850 8740
rect 30090 8550 30550 8740
rect 21870 8310 21970 8550
rect 25370 8310 25470 8550
rect 28870 8310 28970 8550
rect 20290 8140 20750 8310
rect 20990 8140 21450 8310
rect 21690 8140 22150 8310
rect 22390 8140 22850 8310
rect 23090 8140 23550 8310
rect 20290 8040 23550 8140
rect 20290 7850 20750 8040
rect 20990 7850 21450 8040
rect 21690 7850 22150 8040
rect 22390 7850 22850 8040
rect 23090 7850 23550 8040
rect 23790 8140 24250 8310
rect 24490 8140 24950 8310
rect 25190 8140 25650 8310
rect 25890 8140 26350 8310
rect 26590 8140 27050 8310
rect 23790 8040 27050 8140
rect 23790 7850 24250 8040
rect 24490 7850 24950 8040
rect 25190 7850 25650 8040
rect 25890 7850 26350 8040
rect 26590 7850 27050 8040
rect 27290 8140 27750 8310
rect 27990 8140 28450 8310
rect 28690 8140 29150 8310
rect 29390 8140 29850 8310
rect 30090 8140 30550 8310
rect 27290 8040 30550 8140
rect 27290 7850 27750 8040
rect 27990 7850 28450 8040
rect 28690 7850 29150 8040
rect 29390 7850 29850 8040
rect 30090 7850 30550 8040
rect 21870 7610 21970 7850
rect 25370 7610 25470 7850
rect 28870 7610 28970 7850
rect 20290 7440 20750 7610
rect 20990 7440 21450 7610
rect 21690 7440 22150 7610
rect 22390 7440 22850 7610
rect 23090 7440 23550 7610
rect 20290 7340 23550 7440
rect 20290 7150 20750 7340
rect 20990 7150 21450 7340
rect 21690 7150 22150 7340
rect 22390 7150 22850 7340
rect 23090 7150 23550 7340
rect 23790 7440 24250 7610
rect 24490 7440 24950 7610
rect 25190 7440 25650 7610
rect 25890 7440 26350 7610
rect 26590 7440 27050 7610
rect 23790 7340 27050 7440
rect 23790 7150 24250 7340
rect 24490 7150 24950 7340
rect 25190 7150 25650 7340
rect 25890 7150 26350 7340
rect 26590 7150 27050 7340
rect 27290 7440 27750 7610
rect 27990 7440 28450 7610
rect 28690 7440 29150 7610
rect 29390 7440 29850 7610
rect 30090 7440 30550 7610
rect 27290 7340 30550 7440
rect 27290 7150 27750 7340
rect 27990 7150 28450 7340
rect 28690 7150 29150 7340
rect 29390 7150 29850 7340
rect 30090 7150 30550 7340
rect 19780 6990 19790 7050
rect 19850 6990 19860 7050
rect 19780 6280 19860 6990
rect 21880 6890 21960 7150
rect 21880 6830 21890 6890
rect 21950 6830 21960 6890
rect 21880 6820 21960 6830
rect 23270 6900 23370 6910
rect 23270 6820 23280 6900
rect 23360 6820 23370 6900
rect 23270 6810 23370 6820
rect 25380 6780 25460 7150
rect 28880 6990 28960 7150
rect 28880 6930 28890 6990
rect 28950 6930 28960 6990
rect 28880 6920 28960 6930
rect 30270 6900 30370 6910
rect 30270 6820 30280 6900
rect 30360 6820 30370 6900
rect 30270 6810 30370 6820
rect 25380 6720 25390 6780
rect 25450 6720 25460 6780
rect 25380 6710 25460 6720
rect 26770 6680 26870 6690
rect 26770 6600 26780 6680
rect 26860 6600 26870 6680
rect 26770 6590 26870 6600
rect 19780 6220 19790 6280
rect 19850 6220 19860 6280
rect 19780 6000 19860 6220
rect 19780 5940 19790 6000
rect 19850 5940 19860 6000
rect 19780 5820 19860 5940
rect 19780 5760 19790 5820
rect 19850 5760 19860 5820
rect 19780 3040 19860 5760
rect 19780 2980 19790 3040
rect 19850 2980 19860 3040
rect 19780 630 19860 2980
rect 31330 2160 31410 9730
rect 31330 2100 31340 2160
rect 31400 2100 31410 2160
rect 31330 1640 31410 2100
rect 31330 1580 31340 1640
rect 31400 1580 31410 1640
rect 31330 1260 31410 1580
rect 31330 1200 31340 1260
rect 31400 1200 31410 1260
rect 31330 630 31410 1200
rect 31500 6990 31580 9900
rect 31500 6930 31510 6990
rect 31570 6930 31580 6990
rect 31500 5620 31580 6930
rect 31500 5560 31510 5620
rect 31570 5560 31580 5620
rect 31500 4220 31580 5560
rect 31500 4160 31510 4220
rect 31570 4160 31580 4220
rect 31500 2790 31580 4160
rect 31500 2730 31510 2790
rect 31570 2730 31580 2790
rect 19770 620 19870 630
rect 19770 540 19780 620
rect 19860 540 19870 620
rect 19770 530 19870 540
rect 31320 620 31420 630
rect 31320 540 31330 620
rect 31410 540 31420 620
rect 31320 530 31420 540
rect 31500 470 31580 2730
rect 19600 460 19700 470
rect 19600 380 19610 460
rect 19690 380 19700 460
rect 19600 370 19700 380
rect 31490 460 31590 470
rect 31490 380 31500 460
rect 31580 380 31590 460
rect 31490 370 31590 380
<< via3 >>
rect 19610 9980 19690 9990
rect 19610 9920 19620 9980
rect 19620 9920 19680 9980
rect 19680 9920 19690 9980
rect 19610 9910 19690 9920
rect 31500 9980 31580 9990
rect 31500 9920 31510 9980
rect 31510 9920 31570 9980
rect 31570 9920 31580 9980
rect 31500 9910 31580 9920
rect 19780 9740 19860 9820
rect 31330 9740 31410 9820
rect 23280 6890 23360 6900
rect 23280 6830 23290 6890
rect 23290 6830 23350 6890
rect 23350 6830 23360 6890
rect 23280 6820 23360 6830
rect 30280 6890 30360 6900
rect 30280 6830 30290 6890
rect 30290 6830 30350 6890
rect 30350 6830 30360 6890
rect 30280 6820 30360 6830
rect 26780 6670 26860 6680
rect 26780 6610 26790 6670
rect 26790 6610 26850 6670
rect 26850 6610 26860 6670
rect 26780 6600 26860 6610
rect 19780 540 19860 620
rect 31330 540 31410 620
rect 19610 450 19690 460
rect 19610 390 19620 450
rect 19620 390 19680 450
rect 19680 390 19690 450
rect 19610 380 19690 390
rect 31500 380 31580 460
<< mimcap >>
rect 20320 9530 20720 9680
rect 20320 9450 20480 9530
rect 20560 9450 20720 9530
rect 20320 9280 20720 9450
rect 21020 9530 21420 9680
rect 21020 9450 21180 9530
rect 21260 9450 21420 9530
rect 21020 9280 21420 9450
rect 21720 9530 22120 9680
rect 21720 9450 21880 9530
rect 21960 9450 22120 9530
rect 21720 9280 22120 9450
rect 22420 9530 22820 9680
rect 22420 9450 22580 9530
rect 22660 9450 22820 9530
rect 22420 9280 22820 9450
rect 23120 9530 23520 9680
rect 23120 9450 23280 9530
rect 23360 9450 23520 9530
rect 23120 9280 23520 9450
rect 23820 9530 24220 9680
rect 23820 9450 23980 9530
rect 24060 9450 24220 9530
rect 23820 9280 24220 9450
rect 24520 9530 24920 9680
rect 24520 9450 24680 9530
rect 24760 9450 24920 9530
rect 24520 9280 24920 9450
rect 25220 9530 25620 9680
rect 25220 9450 25380 9530
rect 25460 9450 25620 9530
rect 25220 9280 25620 9450
rect 25920 9530 26320 9680
rect 25920 9450 26080 9530
rect 26160 9450 26320 9530
rect 25920 9280 26320 9450
rect 26620 9530 27020 9680
rect 26620 9450 26780 9530
rect 26860 9450 27020 9530
rect 26620 9280 27020 9450
rect 27320 9530 27720 9680
rect 27320 9450 27480 9530
rect 27560 9450 27720 9530
rect 27320 9280 27720 9450
rect 28020 9530 28420 9680
rect 28020 9450 28180 9530
rect 28260 9450 28420 9530
rect 28020 9280 28420 9450
rect 28720 9530 29120 9680
rect 28720 9450 28880 9530
rect 28960 9450 29120 9530
rect 28720 9280 29120 9450
rect 29420 9530 29820 9680
rect 29420 9450 29580 9530
rect 29660 9450 29820 9530
rect 29420 9280 29820 9450
rect 30120 9530 30520 9680
rect 30120 9450 30280 9530
rect 30360 9450 30520 9530
rect 30120 9280 30520 9450
rect 20320 8830 20720 8980
rect 20320 8750 20480 8830
rect 20560 8750 20720 8830
rect 20320 8580 20720 8750
rect 21020 8830 21420 8980
rect 21020 8750 21180 8830
rect 21260 8750 21420 8830
rect 21020 8580 21420 8750
rect 21720 8830 22120 8980
rect 21720 8750 21880 8830
rect 21960 8750 22120 8830
rect 21720 8580 22120 8750
rect 22420 8830 22820 8980
rect 22420 8750 22580 8830
rect 22660 8750 22820 8830
rect 22420 8580 22820 8750
rect 23120 8830 23520 8980
rect 23120 8750 23280 8830
rect 23360 8750 23520 8830
rect 23120 8580 23520 8750
rect 23820 8830 24220 8980
rect 23820 8750 23980 8830
rect 24060 8750 24220 8830
rect 23820 8580 24220 8750
rect 24520 8830 24920 8980
rect 24520 8750 24680 8830
rect 24760 8750 24920 8830
rect 24520 8580 24920 8750
rect 25220 8830 25620 8980
rect 25220 8750 25380 8830
rect 25460 8750 25620 8830
rect 25220 8580 25620 8750
rect 25920 8830 26320 8980
rect 25920 8750 26080 8830
rect 26160 8750 26320 8830
rect 25920 8580 26320 8750
rect 26620 8830 27020 8980
rect 26620 8750 26780 8830
rect 26860 8750 27020 8830
rect 26620 8580 27020 8750
rect 27320 8830 27720 8980
rect 27320 8750 27480 8830
rect 27560 8750 27720 8830
rect 27320 8580 27720 8750
rect 28020 8830 28420 8980
rect 28020 8750 28180 8830
rect 28260 8750 28420 8830
rect 28020 8580 28420 8750
rect 28720 8830 29120 8980
rect 28720 8750 28880 8830
rect 28960 8750 29120 8830
rect 28720 8580 29120 8750
rect 29420 8830 29820 8980
rect 29420 8750 29580 8830
rect 29660 8750 29820 8830
rect 29420 8580 29820 8750
rect 30120 8830 30520 8980
rect 30120 8750 30280 8830
rect 30360 8750 30520 8830
rect 30120 8580 30520 8750
rect 20320 8130 20720 8280
rect 20320 8050 20480 8130
rect 20560 8050 20720 8130
rect 20320 7880 20720 8050
rect 21020 8130 21420 8280
rect 21020 8050 21180 8130
rect 21260 8050 21420 8130
rect 21020 7880 21420 8050
rect 21720 8130 22120 8280
rect 21720 8050 21880 8130
rect 21960 8050 22120 8130
rect 21720 7880 22120 8050
rect 22420 8130 22820 8280
rect 22420 8050 22580 8130
rect 22660 8050 22820 8130
rect 22420 7880 22820 8050
rect 23120 8130 23520 8280
rect 23120 8050 23280 8130
rect 23360 8050 23520 8130
rect 23120 7880 23520 8050
rect 23820 8130 24220 8280
rect 23820 8050 23980 8130
rect 24060 8050 24220 8130
rect 23820 7880 24220 8050
rect 24520 8130 24920 8280
rect 24520 8050 24680 8130
rect 24760 8050 24920 8130
rect 24520 7880 24920 8050
rect 25220 8130 25620 8280
rect 25220 8050 25380 8130
rect 25460 8050 25620 8130
rect 25220 7880 25620 8050
rect 25920 8130 26320 8280
rect 25920 8050 26080 8130
rect 26160 8050 26320 8130
rect 25920 7880 26320 8050
rect 26620 8130 27020 8280
rect 26620 8050 26780 8130
rect 26860 8050 27020 8130
rect 26620 7880 27020 8050
rect 27320 8130 27720 8280
rect 27320 8050 27480 8130
rect 27560 8050 27720 8130
rect 27320 7880 27720 8050
rect 28020 8130 28420 8280
rect 28020 8050 28180 8130
rect 28260 8050 28420 8130
rect 28020 7880 28420 8050
rect 28720 8130 29120 8280
rect 28720 8050 28880 8130
rect 28960 8050 29120 8130
rect 28720 7880 29120 8050
rect 29420 8130 29820 8280
rect 29420 8050 29580 8130
rect 29660 8050 29820 8130
rect 29420 7880 29820 8050
rect 30120 8130 30520 8280
rect 30120 8050 30280 8130
rect 30360 8050 30520 8130
rect 30120 7880 30520 8050
rect 20320 7430 20720 7580
rect 20320 7350 20480 7430
rect 20560 7350 20720 7430
rect 20320 7180 20720 7350
rect 21020 7430 21420 7580
rect 21020 7350 21180 7430
rect 21260 7350 21420 7430
rect 21020 7180 21420 7350
rect 21720 7430 22120 7580
rect 21720 7350 21880 7430
rect 21960 7350 22120 7430
rect 21720 7180 22120 7350
rect 22420 7430 22820 7580
rect 22420 7350 22580 7430
rect 22660 7350 22820 7430
rect 22420 7180 22820 7350
rect 23120 7430 23520 7580
rect 23120 7350 23280 7430
rect 23360 7350 23520 7430
rect 23120 7180 23520 7350
rect 23820 7430 24220 7580
rect 23820 7350 23980 7430
rect 24060 7350 24220 7430
rect 23820 7180 24220 7350
rect 24520 7430 24920 7580
rect 24520 7350 24680 7430
rect 24760 7350 24920 7430
rect 24520 7180 24920 7350
rect 25220 7430 25620 7580
rect 25220 7350 25380 7430
rect 25460 7350 25620 7430
rect 25220 7180 25620 7350
rect 25920 7430 26320 7580
rect 25920 7350 26080 7430
rect 26160 7350 26320 7430
rect 25920 7180 26320 7350
rect 26620 7430 27020 7580
rect 26620 7350 26780 7430
rect 26860 7350 27020 7430
rect 26620 7180 27020 7350
rect 27320 7430 27720 7580
rect 27320 7350 27480 7430
rect 27560 7350 27720 7430
rect 27320 7180 27720 7350
rect 28020 7430 28420 7580
rect 28020 7350 28180 7430
rect 28260 7350 28420 7430
rect 28020 7180 28420 7350
rect 28720 7430 29120 7580
rect 28720 7350 28880 7430
rect 28960 7350 29120 7430
rect 28720 7180 29120 7350
rect 29420 7430 29820 7580
rect 29420 7350 29580 7430
rect 29660 7350 29820 7430
rect 29420 7180 29820 7350
rect 30120 7430 30520 7580
rect 30120 7350 30280 7430
rect 30360 7350 30520 7430
rect 30120 7180 30520 7350
<< mimcapcontact >>
rect 20480 9450 20560 9530
rect 21180 9450 21260 9530
rect 21880 9450 21960 9530
rect 22580 9450 22660 9530
rect 23280 9450 23360 9530
rect 23980 9450 24060 9530
rect 24680 9450 24760 9530
rect 25380 9450 25460 9530
rect 26080 9450 26160 9530
rect 26780 9450 26860 9530
rect 27480 9450 27560 9530
rect 28180 9450 28260 9530
rect 28880 9450 28960 9530
rect 29580 9450 29660 9530
rect 30280 9450 30360 9530
rect 20480 8750 20560 8830
rect 21180 8750 21260 8830
rect 21880 8750 21960 8830
rect 22580 8750 22660 8830
rect 23280 8750 23360 8830
rect 23980 8750 24060 8830
rect 24680 8750 24760 8830
rect 25380 8750 25460 8830
rect 26080 8750 26160 8830
rect 26780 8750 26860 8830
rect 27480 8750 27560 8830
rect 28180 8750 28260 8830
rect 28880 8750 28960 8830
rect 29580 8750 29660 8830
rect 30280 8750 30360 8830
rect 20480 8050 20560 8130
rect 21180 8050 21260 8130
rect 21880 8050 21960 8130
rect 22580 8050 22660 8130
rect 23280 8050 23360 8130
rect 23980 8050 24060 8130
rect 24680 8050 24760 8130
rect 25380 8050 25460 8130
rect 26080 8050 26160 8130
rect 26780 8050 26860 8130
rect 27480 8050 27560 8130
rect 28180 8050 28260 8130
rect 28880 8050 28960 8130
rect 29580 8050 29660 8130
rect 30280 8050 30360 8130
rect 20480 7350 20560 7430
rect 21180 7350 21260 7430
rect 21880 7350 21960 7430
rect 22580 7350 22660 7430
rect 23280 7350 23360 7430
rect 23980 7350 24060 7430
rect 24680 7350 24760 7430
rect 25380 7350 25460 7430
rect 26080 7350 26160 7430
rect 26780 7350 26860 7430
rect 27480 7350 27560 7430
rect 28180 7350 28260 7430
rect 28880 7350 28960 7430
rect 29580 7350 29660 7430
rect 30280 7350 30360 7430
<< metal4 >>
rect 19600 9990 31590 10000
rect 19600 9910 19610 9990
rect 19690 9910 31500 9990
rect 31580 9910 31590 9990
rect 19600 9900 31590 9910
rect 19770 9820 31420 9830
rect 19770 9740 19780 9820
rect 19860 9740 31330 9820
rect 31410 9740 31420 9820
rect 19770 9730 31420 9740
rect 20470 9530 23370 9540
rect 20470 9450 20480 9530
rect 20560 9450 21180 9530
rect 21260 9450 21880 9530
rect 21960 9450 22580 9530
rect 22660 9450 23280 9530
rect 23360 9450 23370 9530
rect 20470 9440 23370 9450
rect 23970 9530 26870 9540
rect 23970 9450 23980 9530
rect 24060 9450 24680 9530
rect 24760 9450 25380 9530
rect 25460 9450 26080 9530
rect 26160 9450 26780 9530
rect 26860 9450 26870 9530
rect 23970 9440 26870 9450
rect 27470 9530 30370 9540
rect 27470 9450 27480 9530
rect 27560 9450 28180 9530
rect 28260 9450 28880 9530
rect 28960 9450 29580 9530
rect 29660 9450 30280 9530
rect 30360 9450 30370 9530
rect 27470 9440 30370 9450
rect 21870 8840 21970 9440
rect 25370 8840 25470 9440
rect 28870 8840 28970 9440
rect 20470 8830 23370 8840
rect 20470 8750 20480 8830
rect 20560 8750 21180 8830
rect 21260 8750 21880 8830
rect 21960 8750 22580 8830
rect 22660 8750 23280 8830
rect 23360 8750 23370 8830
rect 20470 8740 23370 8750
rect 23970 8830 26870 8840
rect 23970 8750 23980 8830
rect 24060 8750 24680 8830
rect 24760 8750 25380 8830
rect 25460 8750 26080 8830
rect 26160 8750 26780 8830
rect 26860 8750 26870 8830
rect 23970 8740 26870 8750
rect 27470 8830 30370 8840
rect 27470 8750 27480 8830
rect 27560 8750 28180 8830
rect 28260 8750 28880 8830
rect 28960 8750 29580 8830
rect 29660 8750 30280 8830
rect 30360 8750 30370 8830
rect 27470 8740 30370 8750
rect 21870 8140 21970 8740
rect 25370 8140 25470 8740
rect 28870 8140 28970 8740
rect 20470 8130 23370 8140
rect 20470 8050 20480 8130
rect 20560 8050 21180 8130
rect 21260 8050 21880 8130
rect 21960 8050 22580 8130
rect 22660 8050 23280 8130
rect 23360 8050 23370 8130
rect 20470 8040 23370 8050
rect 23970 8130 26870 8140
rect 23970 8050 23980 8130
rect 24060 8050 24680 8130
rect 24760 8050 25380 8130
rect 25460 8050 26080 8130
rect 26160 8050 26780 8130
rect 26860 8050 26870 8130
rect 23970 8040 26870 8050
rect 27470 8130 30370 8140
rect 27470 8050 27480 8130
rect 27560 8050 28180 8130
rect 28260 8050 28880 8130
rect 28960 8050 29580 8130
rect 29660 8050 30280 8130
rect 30360 8050 30370 8130
rect 27470 8040 30370 8050
rect 21870 7440 21970 8040
rect 25370 7440 25470 8040
rect 28870 7440 28970 8040
rect 20470 7430 23370 7440
rect 20470 7350 20480 7430
rect 20560 7350 21180 7430
rect 21260 7350 21880 7430
rect 21960 7350 22580 7430
rect 22660 7350 23280 7430
rect 23360 7350 23370 7430
rect 20470 7340 23370 7350
rect 23970 7430 26870 7440
rect 23970 7350 23980 7430
rect 24060 7350 24680 7430
rect 24760 7350 25380 7430
rect 25460 7350 26080 7430
rect 26160 7350 26780 7430
rect 26860 7350 26870 7430
rect 23970 7340 26870 7350
rect 27470 7430 30370 7440
rect 27470 7350 27480 7430
rect 27560 7350 28180 7430
rect 28260 7350 28880 7430
rect 28960 7350 29580 7430
rect 29660 7350 30280 7430
rect 30360 7350 30370 7430
rect 27470 7340 30370 7350
rect 23270 6900 23370 7340
rect 23270 6820 23280 6900
rect 23360 6820 23370 6900
rect 23270 6810 23370 6820
rect 26770 6680 26870 7340
rect 30270 6900 30370 7340
rect 30270 6820 30280 6900
rect 30360 6820 30370 6900
rect 30270 6810 30370 6820
rect 26770 6600 26780 6680
rect 26860 6600 26870 6680
rect 26770 6590 26870 6600
rect 19770 620 31420 630
rect 19770 540 19780 620
rect 19860 540 31330 620
rect 31410 540 31420 620
rect 19770 530 31420 540
rect 19600 460 31590 470
rect 19600 380 19610 460
rect 19690 380 31500 460
rect 31580 380 31590 460
rect 19600 370 31590 380
<< labels >>
flabel metal2 20910 6880 20910 6880 1 FreeSans 800 0 0 80 cap_res1
flabel metal2 32560 6150 32560 6150 1 FreeSans 800 0 0 400 VB1_CUR_BIAS
port 1 n
flabel metal2 32600 6040 32600 6040 3 FreeSans 800 0 400 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 32560 5910 32560 5910 5 FreeSans 800 0 0 -400 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal3 31580 8800 31580 8800 3 FreeSans 1600 0 160 0 VDDA
port 4 e
flabel metal3 31410 8350 31410 8350 3 FreeSans 1600 0 160 0 GNDA
port 2 e
flabel metal1 26550 0 26550 0 7 FreeSans 800 0 -800 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 27650 -110 27650 -110 5 FreeSans 800 0 0 -400 VB2_CUR_BIAS
port 5 s
flabel metal1 28030 0 28030 0 3 FreeSans 800 0 400 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 29450 -110 29450 -110 5 FreeSans 800 0 0 -400 VB3_CUR_BIAS
port 6 s
flabel metal2 32600 3410 32600 3410 3 FreeSans 800 0 400 0 ERR_AMP_REF
port 3 e
flabel metal1 30130 1780 30130 1780 3 FreeSans 800 0 400 0 START_UP_NFET1
flabel metal2 27430 2960 27430 2960 3 FreeSans 800 0 80 0 V_p1
flabel poly 29430 4680 29430 4680 5 FreeSans 800 0 0 -80 V_TOP
flabel metal2 30430 3100 30430 3100 1 FreeSans 800 0 0 160 V_CUR_REF_REG
flabel metal2 28910 2960 28910 2960 7 FreeSans 800 0 -80 0 V_p2
flabel metal2 30530 3690 30530 3690 5 FreeSans 800 0 0 -80 V_mir2
flabel metal2 25810 3690 25810 3690 5 FreeSans 800 0 0 -80 V_mir1
flabel metal3 25460 6750 25460 6750 3 FreeSans 800 0 80 0 cap_res2
flabel metal1 25210 2210 25210 2210 3 FreeSans 800 0 400 0 START_UP
flabel metal1 25120 1290 25120 1290 3 FreeSans 800 0 80 0 NFET_GATE_10uA
flabel metal2 26100 3390 26100 3390 5 FreeSans 800 0 0 -160 Vin-
flabel metal2 26110 3100 26110 3100 1 FreeSans 800 0 0 160 Vin+
flabel locali s 22180 3422 22298 3462 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 22203 3572 22304 3621 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 22144 2946 22392 3050 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 22180 4782 22298 4822 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 22203 4932 22304 4981 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 22144 4306 22392 4410 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 22180 2062 22298 2102 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 22203 2212 22304 2261 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 22144 1586 22392 1690 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 20820 4782 20938 4822 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 20843 4932 20944 4981 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 20784 4306 21032 4410 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 20820 3422 20938 3462 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 20843 3572 20944 3621 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 20784 2946 21032 3050 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 20820 2062 20938 2102 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 20843 2212 20944 2261 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 20784 1586 21032 1690 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 23540 4782 23658 4822 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 23563 4932 23664 4981 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 23504 4306 23752 4410 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 23540 2062 23658 2102 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 23563 2212 23664 2261 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 23504 1586 23752 1690 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel locali s 23540 3422 23658 3462 0 FreeSans 400 0 0 0 Base
port 4 nsew
flabel locali s 23563 3572 23664 3621 0 FreeSans 400 0 0 0 Collector
port 3 nsew
flabel locali s 23504 2946 23752 3050 0 FreeSans 400 0 0 0 Emitter
port 2 nsew
flabel metal1 24360 1620 24360 1620 3 FreeSans 800 0 80 0 Vbe2
<< end >>
