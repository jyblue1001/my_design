* PEX produced on Fri Jul  4 08:03:05 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_7.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_7 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t299 bgr_0.V_TOP.t14 bgr_0.Vin-.t3 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA.t219 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 bgr_0.V_TOP.t15 VDDA.t297 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA.t311 GNDA.t313 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X5 two_stage_opamp_dummy_magic_0.VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t224 GNDA.t310 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_0.X.t13 GNDA.t15 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X8 two_stage_opamp_dummy_magic_0.VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 two_stage_opamp_dummy_magic_0.VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.t1 GNDA.t332 GNDA.t331 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X11 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 bgr_0.V_TOP.t16 VDDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 VDDA.t86 bgr_0.V_mir2.t12 bgr_0.V_mir2.t13 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X14 two_stage_opamp_dummy_magic_0.V_err_gate.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 two_stage_opamp_dummy_magic_0.VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 two_stage_opamp_dummy_magic_0.VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 a_8420_8490.t9 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD3.t26 two_stage_opamp_dummy_magic_0.VD3.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X18 VDDA.t453 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.VOUT+.t12 VDDA.t452 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X19 two_stage_opamp_dummy_magic_0.X.t11 GNDA.t307 GNDA.t309 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X20 two_stage_opamp_dummy_magic_0.VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 two_stage_opamp_dummy_magic_0.VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t195 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.VOUT+.t11 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X23 VDDA.t97 bgr_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X24 two_stage_opamp_dummy_magic_0.VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 a_14520_5068.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t108 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X26 bgr_0.V_TOP.t17 VDDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 two_stage_opamp_dummy_magic_0.VOUT-.t17 GNDA.t304 GNDA.t306 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X28 VDDA.t71 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X29 VDDA.t435 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t8 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X30 two_stage_opamp_dummy_magic_0.VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t129 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X32 two_stage_opamp_dummy_magic_0.VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_0.VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 two_stage_opamp_dummy_magic_0.VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 two_stage_opamp_dummy_magic_0.VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 two_stage_opamp_dummy_magic_0.VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 two_stage_opamp_dummy_magic_0.VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 two_stage_opamp_dummy_magic_0.V_p_mir.t2 bgr_0.TAIL_CUR_MIR_BIAS.t12 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X40 VDDA.t17 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.VOUT-.t2 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X41 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 two_stage_opamp_dummy_magic_0.Y.t15 VDDA.t213 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X42 two_stage_opamp_dummy_magic_0.VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 bgr_0.V_mir2.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 bgr_0.V_p_2.t5 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X44 bgr_0.Vin-.t4 bgr_0.V_TOP.t18 VDDA.t294 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X45 VDDA.t414 VDDA.t412 two_stage_opamp_dummy_magic_0.V_err_gate.t9 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 GNDA.t49 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X47 GNDA.t38 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X49 two_stage_opamp_dummy_magic_0.VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 two_stage_opamp_dummy_magic_0.VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 a_8420_8490.t8 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.VD3.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X52 two_stage_opamp_dummy_magic_0.V_err_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 two_stage_opamp_dummy_magic_0.Y.t10 GNDA.t301 GNDA.t303 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X54 two_stage_opamp_dummy_magic_0.Y.t11 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA.t314 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X55 two_stage_opamp_dummy_magic_0.VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 two_stage_opamp_dummy_magic_0.VOUT-.t4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X57 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 two_stage_opamp_dummy_magic_0.Y.t16 GNDA.t340 VDDA.t449 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X58 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X59 two_stage_opamp_dummy_magic_0.VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 GNDA.t61 bgr_0.TAIL_CUR_MIR_BIAS.t13 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X62 VDDA.t411 VDDA.t409 bgr_0.V_TOP.t11 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X63 GNDA.t116 bgr_0.TAIL_CUR_MIR_BIAS.t14 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X64 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_0.X.t15 VDDA.t18 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X65 two_stage_opamp_dummy_magic_0.VD1.t19 VIN-.t0 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X66 two_stage_opamp_dummy_magic_0.V_err_p.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X67 two_stage_opamp_dummy_magic_0.VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 GNDA.t40 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X69 GNDA.t300 GNDA.t298 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X70 VDDA.t444 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t9 VDDA.t443 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X71 two_stage_opamp_dummy_magic_0.VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 two_stage_opamp_dummy_magic_0.VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t215 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X74 two_stage_opamp_dummy_magic_0.VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 two_stage_opamp_dummy_magic_0.VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 two_stage_opamp_dummy_magic_0.VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 two_stage_opamp_dummy_magic_0.VD1.t3 VIN-.t1 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X78 two_stage_opamp_dummy_magic_0.VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 bgr_0.NFET_GATE_10uA.t0 bgr_0.PFET_GATE_10uA.t11 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X80 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t217 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X81 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VDDA.t32 bgr_0.PFET_GATE_10uA.t12 bgr_0.TAIL_CUR_MIR_BIAS.t7 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X83 two_stage_opamp_dummy_magic_0.VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VDDA.t408 VDDA.t406 bgr_0.NFET_GATE_10uA.t3 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X85 VDDA.t220 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.VOUT+.t10 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X86 VDDA.t26 bgr_0.1st_Vout_1.t14 bgr_0.V_TOP.t1 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X87 GNDA.t297 GNDA.t295 two_stage_opamp_dummy_magic_0.VD1.t16 GNDA.t296 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X88 two_stage_opamp_dummy_magic_0.VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 two_stage_opamp_dummy_magic_0.VD4.t36 VDDA.t403 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X90 two_stage_opamp_dummy_magic_0.VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 two_stage_opamp_dummy_magic_0.VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_0.VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 VDDA.t193 bgr_0.V_mir2.t10 bgr_0.V_mir2.t11 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X94 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.VD4.t3 a_10480_8490.t1 two_stage_opamp_dummy_magic_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X95 GNDA.t68 bgr_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X96 VDDA.t89 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t11 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X97 two_stage_opamp_dummy_magic_0.VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 two_stage_opamp_dummy_magic_0.Vb3.t4 bgr_0.NFET_GATE_10uA.t9 GNDA.t70 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X99 GNDA.t294 GNDA.t292 two_stage_opamp_dummy_magic_0.VD1.t15 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X100 VDDA.t207 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t7 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X101 two_stage_opamp_dummy_magic_0.VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 bgr_0.V_TOP.t6 bgr_0.cap_res1.t20 GNDA.t85 sky130_fd_pr__res_high_po_0p35 l=2.05
X103 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_0.Y.t18 VDDA.t98 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X104 two_stage_opamp_dummy_magic_0.V_p.t21 bgr_0.TAIL_CUR_MIR_BIAS.t15 GNDA.t342 GNDA.t341 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X105 a_11220_17410.t0 GNDA.t81 GNDA.t80 sky130_fd_pr__res_xhigh_po_0p35 l=6
X106 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_0.Y.t19 VDDA.t169 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X107 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X108 two_stage_opamp_dummy_magic_0.VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 two_stage_opamp_dummy_magic_0.Vb1.t1 bgr_0.PFET_GATE_10uA.t13 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X110 GNDA.t291 GNDA.t289 two_stage_opamp_dummy_magic_0.X.t10 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X111 two_stage_opamp_dummy_magic_0.VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 two_stage_opamp_dummy_magic_0.VOUT-.t18 a_5750_2276.t1 GNDA.t338 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X113 bgr_0.PFET_GATE_10uA.t3 bgr_0.1st_Vout_2.t13 VDDA.t179 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X114 two_stage_opamp_dummy_magic_0.VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 GNDA.t118 bgr_0.TAIL_CUR_MIR_BIAS.t16 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X116 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb3.t8 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 two_stage_opamp_dummy_magic_0.VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 two_stage_opamp_dummy_magic_0.VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 two_stage_opamp_dummy_magic_0.VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 two_stage_opamp_dummy_magic_0.VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 two_stage_opamp_dummy_magic_0.VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VDDA.t199 bgr_0.V_mir1.t10 bgr_0.V_mir1.t11 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X123 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_0.X.t16 VDDA.t190 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X124 two_stage_opamp_dummy_magic_0.VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 two_stage_opamp_dummy_magic_0.VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X127 two_stage_opamp_dummy_magic_0.VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VDDA.t211 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t6 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.Vb3.t9 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X131 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t123 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X132 bgr_0.V_TOP.t19 VDDA.t292 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.Vb2.t13 a_8420_8490.t7 two_stage_opamp_dummy_magic_0.VD3.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X134 two_stage_opamp_dummy_magic_0.VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 GNDA.t288 GNDA.t286 two_stage_opamp_dummy_magic_0.Y.t9 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X137 two_stage_opamp_dummy_magic_0.VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 a_14640_5068.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA.t72 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X139 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X140 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t283 GNDA.t285 GNDA.t284 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X141 two_stage_opamp_dummy_magic_0.VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 two_stage_opamp_dummy_magic_0.VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 two_stage_opamp_dummy_magic_0.V_p.t30 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 two_stage_opamp_dummy_magic_0.VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VDDA.t173 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t6 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X146 two_stage_opamp_dummy_magic_0.VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 two_stage_opamp_dummy_magic_0.VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 a_13730_17020.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t102 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X150 GNDA.t89 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X151 two_stage_opamp_dummy_magic_0.V_p.t27 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X152 two_stage_opamp_dummy_magic_0.VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 bgr_0.V_CUR_REF_REG.t1 VDDA.t400 VDDA.t402 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X154 a_11220_17410.t1 a_12828_17530.t0 GNDA.t80 sky130_fd_pr__res_xhigh_po_0p35 l=6
X155 two_stage_opamp_dummy_magic_0.VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VDDA.t117 two_stage_opamp_dummy_magic_0.X.t19 two_stage_opamp_dummy_magic_0.VOUT-.t8 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X157 two_stage_opamp_dummy_magic_0.VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 bgr_0.TAIL_CUR_MIR_BIAS.t6 bgr_0.PFET_GATE_10uA.t14 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X159 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_0.Y.t20 VDDA.t170 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X160 two_stage_opamp_dummy_magic_0.VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 two_stage_opamp_dummy_magic_0.VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 two_stage_opamp_dummy_magic_0.V_p.t19 bgr_0.TAIL_CUR_MIR_BIAS.t17 GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X163 VDDA.t155 bgr_0.PFET_GATE_10uA.t15 bgr_0.V_CUR_REF_REG.t0 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X164 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X165 two_stage_opamp_dummy_magic_0.VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 bgr_0.PFET_GATE_10uA.t4 bgr_0.cap_res2.t20 GNDA.t121 sky130_fd_pr__res_high_po_0p35 l=2.05
X167 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.Vb2.t14 a_8420_8490.t6 two_stage_opamp_dummy_magic_0.VD3.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X168 bgr_0.V_p_1.t9 bgr_0.Vin-.t8 bgr_0.V_mir1.t12 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X169 VDDA.t36 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 two_stage_opamp_dummy_magic_0.VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 two_stage_opamp_dummy_magic_0.VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 two_stage_opamp_dummy_magic_0.VD2.t3 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t0 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X173 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 two_stage_opamp_dummy_magic_0.VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 two_stage_opamp_dummy_magic_0.VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VDDA.t421 bgr_0.1st_Vout_1.t19 bgr_0.V_TOP.t9 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X177 VDDA.t291 bgr_0.V_TOP.t20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X178 two_stage_opamp_dummy_magic_0.VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 GNDA.t98 bgr_0.TAIL_CUR_MIR_BIAS.t18 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X180 two_stage_opamp_dummy_magic_0.VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 bgr_0.V_p_2.t0 bgr_0.V_CUR_REF_REG.t3 bgr_0.1st_Vout_2.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X182 two_stage_opamp_dummy_magic_0.VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 two_stage_opamp_dummy_magic_0.VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 two_stage_opamp_dummy_magic_0.VOUT-.t7 two_stage_opamp_dummy_magic_0.X.t20 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X185 two_stage_opamp_dummy_magic_0.VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 bgr_0.V_p_1.t8 bgr_0.Vin-.t9 bgr_0.V_mir1.t15 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X187 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 GNDA.t100 bgr_0.TAIL_CUR_MIR_BIAS.t19 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X189 bgr_0.V_TOP.t0 VDDA.t397 VDDA.t399 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X190 two_stage_opamp_dummy_magic_0.VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_0.Vin-.t0 bgr_0.START_UP.t6 bgr_0.V_TOP.t5 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X192 VDDA.t396 VDDA.t394 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X193 two_stage_opamp_dummy_magic_0.VD1.t12 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.Y.t2 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X194 two_stage_opamp_dummy_magic_0.VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 two_stage_opamp_dummy_magic_0.VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_0.V_TOP.t21 VDDA.t281 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X199 two_stage_opamp_dummy_magic_0.VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 two_stage_opamp_dummy_magic_0.VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VDDA.t205 two_stage_opamp_dummy_magic_0.Vb3.t11 two_stage_opamp_dummy_magic_0.VD4.t32 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X202 GNDA.t347 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 VDDA.t468 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X203 two_stage_opamp_dummy_magic_0.VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 two_stage_opamp_dummy_magic_0.V_p.t16 bgr_0.TAIL_CUR_MIR_BIAS.t20 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X205 a_13730_17020.t1 GNDA.t164 GNDA.t102 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X206 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 bgr_0.V_TOP.t22 VDDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.VD3.t30 a_8420_8490.t11 two_stage_opamp_dummy_magic_0.VD3.t31 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X209 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t391 VDDA.t393 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X210 a_11220_17290.t1 a_12828_17650.t0 GNDA.t80 sky130_fd_pr__res_xhigh_po_0p35 l=6
X211 VDDA.t20 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD3.t1 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X212 two_stage_opamp_dummy_magic_0.VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_0.VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 two_stage_opamp_dummy_magic_0.VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 two_stage_opamp_dummy_magic_0.VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 bgr_0.V_p_2.t10 bgr_0.V_CUR_REF_REG.t4 bgr_0.1st_Vout_2.t10 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X217 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 bgr_0.PFET_GATE_10uA.t16 VDDA.t425 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X218 two_stage_opamp_dummy_magic_0.VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VDDA.t30 bgr_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X220 two_stage_opamp_dummy_magic_0.V_p.t25 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X221 two_stage_opamp_dummy_magic_0.VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 GNDA.t29 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 two_stage_opamp_dummy_magic_0.VOUT+.t0 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X223 GNDA.t76 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X224 a_11220_17290.t0 GNDA.t124 GNDA.t80 sky130_fd_pr__res_xhigh_po_0p35 l=6
X225 two_stage_opamp_dummy_magic_0.V_p.t1 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X226 bgr_0.TAIL_CUR_MIR_BIAS.t11 GNDA.t281 GNDA.t282 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X227 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 two_stage_opamp_dummy_magic_0.VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 two_stage_opamp_dummy_magic_0.VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 bgr_0.START_UP.t5 bgr_0.V_TOP.t23 VDDA.t289 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X231 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t5 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X232 two_stage_opamp_dummy_magic_0.V_p.t15 bgr_0.TAIL_CUR_MIR_BIAS.t21 GNDA.t120 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X233 bgr_0.1st_Vout_2.t5 bgr_0.V_mir2.t18 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X234 bgr_0.V_TOP.t24 VDDA.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 two_stage_opamp_dummy_magic_0.VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 two_stage_opamp_dummy_magic_0.VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 two_stage_opamp_dummy_magic_0.VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 two_stage_opamp_dummy_magic_0.VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDDA.t112 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD4.t29 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X240 VDDA.t446 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t10 VDDA.t445 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X241 two_stage_opamp_dummy_magic_0.VOUT+.t9 two_stage_opamp_dummy_magic_0.Y.t22 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X242 two_stage_opamp_dummy_magic_0.VD2.t16 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t9 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X243 two_stage_opamp_dummy_magic_0.VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 two_stage_opamp_dummy_magic_0.VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 GNDA.t6 bgr_0.TAIL_CUR_MIR_BIAS.t22 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X247 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t9 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X248 GNDA.t280 GNDA.t278 two_stage_opamp_dummy_magic_0.VOUT+.t17 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X249 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 two_stage_opamp_dummy_magic_0.X.t22 VDDA.t231 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X250 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t388 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X251 two_stage_opamp_dummy_magic_0.VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 two_stage_opamp_dummy_magic_0.VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VDDA.t243 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.VD3.t35 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X254 two_stage_opamp_dummy_magic_0.VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 two_stage_opamp_dummy_magic_0.VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 two_stage_opamp_dummy_magic_0.VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 bgr_0.V_TOP.t25 VDDA.t286 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 GNDA.t224 GNDA.t264 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X259 two_stage_opamp_dummy_magic_0.VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 two_stage_opamp_dummy_magic_0.VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 two_stage_opamp_dummy_magic_0.VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VDDA.t230 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD4.t34 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X263 two_stage_opamp_dummy_magic_0.VOUT-.t13 two_stage_opamp_dummy_magic_0.X.t23 VDDA.t233 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X264 a_8420_8490.t5 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X265 two_stage_opamp_dummy_magic_0.VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 GNDA.t153 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X268 two_stage_opamp_dummy_magic_0.VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDDA.t166 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t10 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X270 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X271 two_stage_opamp_dummy_magic_0.VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 a_14640_5068.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X273 VDDA.t168 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X274 two_stage_opamp_dummy_magic_0.VD1.t11 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X275 two_stage_opamp_dummy_magic_0.VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X277 bgr_0.V_mir2.t9 bgr_0.V_mir2.t8 VDDA.t108 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X278 VDDA.t285 bgr_0.V_TOP.t26 bgr_0.Vin-.t5 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X279 GNDA.t109 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X280 VDDA.t387 VDDA.t385 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 bgr_0.PFET_GATE_10uA.t18 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X282 bgr_0.TAIL_CUR_MIR_BIAS.t8 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X283 two_stage_opamp_dummy_magic_0.V_p.t37 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t325 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X284 two_stage_opamp_dummy_magic_0.VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t382 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=1.28 ps=7.2 w=3.2 l=0.2
X286 VDDA.t234 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X287 two_stage_opamp_dummy_magic_0.VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 two_stage_opamp_dummy_magic_0.VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 bgr_0.Vin-.t7 a_12828_17650.t1 GNDA.t80 sky130_fd_pr__res_xhigh_po_0p35 l=6
X290 two_stage_opamp_dummy_magic_0.VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 two_stage_opamp_dummy_magic_0.VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 two_stage_opamp_dummy_magic_0.VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 GNDA.t224 GNDA.t277 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X294 two_stage_opamp_dummy_magic_0.V_p.t32 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X295 a_8420_8490.t4 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X296 VDDA.t228 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.VD4.t33 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X297 GNDA.t176 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X298 two_stage_opamp_dummy_magic_0.VD3.t37 VDDA.t379 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X299 GNDA.t96 two_stage_opamp_dummy_magic_0.X.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X300 two_stage_opamp_dummy_magic_0.VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 two_stage_opamp_dummy_magic_0.VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_0.VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 GNDA.t155 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X305 bgr_0.PFET_GATE_10uA.t0 bgr_0.1st_Vout_2.t19 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X306 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t10 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X307 two_stage_opamp_dummy_magic_0.VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 two_stage_opamp_dummy_magic_0.VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t274 GNDA.t276 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X310 GNDA.t273 GNDA.t271 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X311 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X312 two_stage_opamp_dummy_magic_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t12 GNDA.t149 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X313 bgr_0.START_UP.t1 bgr_0.START_UP.t0 bgr_0.START_UP_NFET1.t0 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X314 two_stage_opamp_dummy_magic_0.VOUT+.t8 two_stage_opamp_dummy_magic_0.Y.t24 VDDA.t464 VDDA.t463 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X315 two_stage_opamp_dummy_magic_0.VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 two_stage_opamp_dummy_magic_0.VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_0.VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 two_stage_opamp_dummy_magic_0.VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 two_stage_opamp_dummy_magic_0.VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 two_stage_opamp_dummy_magic_0.VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 two_stage_opamp_dummy_magic_0.VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 two_stage_opamp_dummy_magic_0.VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 GNDA.t151 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 bgr_0.V_p_1.t3 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t3 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X325 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t136 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X326 two_stage_opamp_dummy_magic_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t14 GNDA.t183 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X327 two_stage_opamp_dummy_magic_0.VOUT+.t16 GNDA.t268 GNDA.t270 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X328 two_stage_opamp_dummy_magic_0.Vb2.t2 bgr_0.NFET_GATE_10uA.t15 GNDA.t185 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X329 two_stage_opamp_dummy_magic_0.VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.Vb2.t17 a_10480_8490.t11 two_stage_opamp_dummy_magic_0.VD4.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X331 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 two_stage_opamp_dummy_magic_0.VOUT-.t10 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X333 two_stage_opamp_dummy_magic_0.VOUT-.t6 two_stage_opamp_dummy_magic_0.X.t28 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X334 VDDA.t67 two_stage_opamp_dummy_magic_0.Y.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X335 bgr_0.Vin+.t4 bgr_0.V_TOP.t27 VDDA.t283 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X336 two_stage_opamp_dummy_magic_0.VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 two_stage_opamp_dummy_magic_0.VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 two_stage_opamp_dummy_magic_0.VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VDDA.t138 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X340 two_stage_opamp_dummy_magic_0.VOUT-.t11 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA.t169 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X341 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.Vb3.t17 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X342 VDDA.t451 bgr_0.PFET_GATE_10uA.t19 bgr_0.TAIL_CUR_MIR_BIAS.t5 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X343 two_stage_opamp_dummy_magic_0.VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 bgr_0.TAIL_CUR_MIR_BIAS.t4 bgr_0.PFET_GATE_10uA.t20 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X345 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t14 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X346 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t211 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X347 two_stage_opamp_dummy_magic_0.VD1.t10 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.Y.t12 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X348 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t1 GNDA.t26 sky130_fd_pr__res_high_po_1p41 l=1.41
X349 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_p.t16 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X350 two_stage_opamp_dummy_magic_0.VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GNDA.t75 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X352 two_stage_opamp_dummy_magic_0.VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 two_stage_opamp_dummy_magic_0.VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 two_stage_opamp_dummy_magic_0.VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 bgr_0.V_TOP.t28 VDDA.t279 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 bgr_0.Vin+.t0 a_12828_17530.t1 GNDA.t80 sky130_fd_pr__res_xhigh_po_0p35 l=6
X357 two_stage_opamp_dummy_magic_0.V_p.t29 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X358 two_stage_opamp_dummy_magic_0.VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 GNDA.t267 GNDA.t265 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X360 two_stage_opamp_dummy_magic_0.VD3.t0 two_stage_opamp_dummy_magic_0.Vb3.t18 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X361 VDDA.t54 two_stage_opamp_dummy_magic_0.X.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X362 two_stage_opamp_dummy_magic_0.VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t261 GNDA.t263 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X365 GNDA.t260 GNDA.t258 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X366 two_stage_opamp_dummy_magic_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t16 GNDA.t145 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X367 GNDA.t147 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X368 two_stage_opamp_dummy_magic_0.V_p.t26 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X369 bgr_0.V_mir1.t7 bgr_0.V_mir1.t6 VDDA.t427 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X370 GNDA.t14 two_stage_opamp_dummy_magic_0.X.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X371 a_5230_5088.t0 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t101 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X372 two_stage_opamp_dummy_magic_0.VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 two_stage_opamp_dummy_magic_0.VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t4 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X375 two_stage_opamp_dummy_magic_0.VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 bgr_0.V_p_2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 bgr_0.V_mir2.t16 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X377 two_stage_opamp_dummy_magic_0.VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VDDA.t433 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.Vb1.t0 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X379 two_stage_opamp_dummy_magic_0.VD2.t8 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t5 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X380 two_stage_opamp_dummy_magic_0.VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 two_stage_opamp_dummy_magic_0.VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 two_stage_opamp_dummy_magic_0.VOUT+.t7 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t120 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X383 two_stage_opamp_dummy_magic_0.VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X385 bgr_0.V_p_1.t2 bgr_0.Vin+.t8 bgr_0.1st_Vout_1.t1 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X386 two_stage_opamp_dummy_magic_0.VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t278 bgr_0.V_TOP.t29 bgr_0.START_UP.t4 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X388 two_stage_opamp_dummy_magic_0.V_err_p.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t149 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X389 two_stage_opamp_dummy_magic_0.VOUT+.t2 a_14240_2276.t1 GNDA.t77 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X390 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.Vb2.t18 a_8420_8490.t3 two_stage_opamp_dummy_magic_0.VD3.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X391 two_stage_opamp_dummy_magic_0.VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X394 two_stage_opamp_dummy_magic_0.VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 two_stage_opamp_dummy_magic_0.VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X397 a_14520_5068.t0 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t79 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X398 bgr_0.V_p_2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 bgr_0.V_mir2.t14 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X399 two_stage_opamp_dummy_magic_0.VOUT-.t0 two_stage_opamp_dummy_magic_0.X.t31 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X400 two_stage_opamp_dummy_magic_0.VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VDDA.t76 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X402 two_stage_opamp_dummy_magic_0.VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VDDA.t151 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t8 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X405 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_0.V_err_p.t15 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X406 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA.t255 GNDA.t257 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X407 two_stage_opamp_dummy_magic_0.VD1.t9 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t8 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X408 two_stage_opamp_dummy_magic_0.VD1.t8 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X409 GNDA.t71 two_stage_opamp_dummy_magic_0.Y.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X410 two_stage_opamp_dummy_magic_0.VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 two_stage_opamp_dummy_magic_0.VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 VDDA.t224 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0.64 ps=3.6 w=3.2 l=0.2
X413 GNDA.t56 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X414 two_stage_opamp_dummy_magic_0.VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 two_stage_opamp_dummy_magic_0.V_p.t4 a_11120_2960# GNDA.t25 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X416 VDDA.t244 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X417 two_stage_opamp_dummy_magic_0.V_p.t40 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA.t348 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X418 bgr_0.1st_Vout_1.t4 bgr_0.V_mir1.t20 VDDA.t185 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X419 VDDA.t93 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t7 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X420 VDDA.t245 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X421 GNDA.t199 VDDA.t469 bgr_0.V_TOP.t2 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X422 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.Vb3.t21 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X423 two_stage_opamp_dummy_magic_0.VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 a_10480_8490.t0 two_stage_opamp_dummy_magic_0.VD4.t0 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X425 GNDA.t209 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X426 two_stage_opamp_dummy_magic_0.VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 two_stage_opamp_dummy_magic_0.VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 bgr_0.1st_Vout_2.t4 bgr_0.V_mir2.t19 VDDA.t62 VDDA.t61 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X429 two_stage_opamp_dummy_magic_0.VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 two_stage_opamp_dummy_magic_0.VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_0.VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 two_stage_opamp_dummy_magic_0.VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 GNDA.t31 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 two_stage_opamp_dummy_magic_0.VOUT-.t3 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X436 VDDA.t442 bgr_0.PFET_GATE_10uA.t22 bgr_0.TAIL_CUR_MIR_BIAS.t3 VDDA.t441 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X437 two_stage_opamp_dummy_magic_0.VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t95 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X439 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 two_stage_opamp_dummy_magic_0.VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 bgr_0.V_TOP.t30 VDDA.t276 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t7 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X443 two_stage_opamp_dummy_magic_0.VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 bgr_0.START_UP.t3 bgr_0.V_TOP.t31 VDDA.t275 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X445 two_stage_opamp_dummy_magic_0.VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 two_stage_opamp_dummy_magic_0.VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 two_stage_opamp_dummy_magic_0.VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 two_stage_opamp_dummy_magic_0.VOUT+.t6 two_stage_opamp_dummy_magic_0.Y.t31 VDDA.t466 VDDA.t465 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X449 two_stage_opamp_dummy_magic_0.VOUT+.t5 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t222 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X450 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 bgr_0.V_mir2.t7 bgr_0.V_mir2.t6 VDDA.t241 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X452 two_stage_opamp_dummy_magic_0.VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 two_stage_opamp_dummy_magic_0.VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 a_10480_8490.t10 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X455 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X457 two_stage_opamp_dummy_magic_0.VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 bgr_0.V_TOP.t10 bgr_0.1st_Vout_1.t27 VDDA.t423 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X459 two_stage_opamp_dummy_magic_0.VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 two_stage_opamp_dummy_magic_0.VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 two_stage_opamp_dummy_magic_0.VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 GNDA.t254 GNDA.t251 GNDA.t253 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X464 GNDA.t224 GNDA.t249 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X465 bgr_0.V_mir2.t5 bgr_0.V_mir2.t4 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X466 VDDA.t273 bgr_0.V_TOP.t32 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X467 GNDA.t63 bgr_0.TAIL_CUR_MIR_BIAS.t23 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X468 VDDA.t437 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t335 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X469 two_stage_opamp_dummy_magic_0.VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 two_stage_opamp_dummy_magic_0.VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VDDA.t378 VDDA.t376 bgr_0.V_TOP.t4 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X472 two_stage_opamp_dummy_magic_0.V_err_gate.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X473 two_stage_opamp_dummy_magic_0.VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VDDA.t164 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X475 two_stage_opamp_dummy_magic_0.VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 bgr_0.V_TOP.t33 VDDA.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 VDDA.t209 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.VD3.t33 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X478 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 VDDA.t373 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X479 GNDA.t196 VDDA.t370 VDDA.t372 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X480 two_stage_opamp_dummy_magic_0.V_p.t12 bgr_0.TAIL_CUR_MIR_BIAS.t24 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X481 two_stage_opamp_dummy_magic_0.VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 two_stage_opamp_dummy_magic_0.VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 two_stage_opamp_dummy_magic_0.VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 GNDA.t224 GNDA.t248 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X485 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 two_stage_opamp_dummy_magic_0.V_p.t2 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X487 bgr_0.V_TOP.t34 VDDA.t270 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VDDA.t113 two_stage_opamp_dummy_magic_0.X.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X489 two_stage_opamp_dummy_magic_0.VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 two_stage_opamp_dummy_magic_0.V_p.t31 two_stage_opamp_dummy_magic_0.Vb1.t2 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X491 two_stage_opamp_dummy_magic_0.VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t26 VDDA.t203 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X493 a_13790_17550.t1 bgr_0.V_CUR_REF_REG.t2 GNDA.t105 sky130_fd_pr__res_xhigh_po_0p35 l=6
X494 GNDA.t207 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X495 two_stage_opamp_dummy_magic_0.VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VDDA.t183 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X497 VDDA.t269 bgr_0.V_TOP.t35 bgr_0.Vin+.t3 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X498 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t367 VDDA.t369 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X499 a_5350_5088.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t42 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X500 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 two_stage_opamp_dummy_magic_0.VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 GNDA.t198 VDDA.t470 bgr_0.V_p_2.t6 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X503 two_stage_opamp_dummy_magic_0.VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 GNDA.t205 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X505 bgr_0.V_p_1.t7 bgr_0.Vin-.t10 bgr_0.V_mir1.t13 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X506 VDDA.t42 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD3.t4 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X507 a_10480_8490.t9 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X508 two_stage_opamp_dummy_magic_0.VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 two_stage_opamp_dummy_magic_0.VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 bgr_0.V_TOP.t12 bgr_0.1st_Vout_1.t30 VDDA.t459 VDDA.t458 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X511 two_stage_opamp_dummy_magic_0.VOUT+.t15 VDDA.t364 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X512 two_stage_opamp_dummy_magic_0.VD2.t11 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.X.t6 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X513 two_stage_opamp_dummy_magic_0.VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 bgr_0.V_TOP.t36 VDDA.t267 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 two_stage_opamp_dummy_magic_0.VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 GNDA.t224 GNDA.t250 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X517 two_stage_opamp_dummy_magic_0.VD1.t17 VIN-.t6 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X518 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_14240_2276.t0 GNDA.t64 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X519 bgr_0.1st_Vout_1.t5 bgr_0.V_mir1.t21 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X520 two_stage_opamp_dummy_magic_0.VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 two_stage_opamp_dummy_magic_0.VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 two_stage_opamp_dummy_magic_0.VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 two_stage_opamp_dummy_magic_0.VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 two_stage_opamp_dummy_magic_0.VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 two_stage_opamp_dummy_magic_0.VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 two_stage_opamp_dummy_magic_0.VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 bgr_0.Vin+.t2 bgr_0.V_TOP.t37 VDDA.t266 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X528 bgr_0.V_mir2.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t2 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X529 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X530 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 bgr_0.PFET_GATE_10uA.t9 VDDA.t471 GNDA.t195 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X532 two_stage_opamp_dummy_magic_0.VD1.t18 VIN-.t7 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X533 two_stage_opamp_dummy_magic_0.VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 two_stage_opamp_dummy_magic_0.VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 two_stage_opamp_dummy_magic_0.VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VDDA.t417 two_stage_opamp_dummy_magic_0.Y.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X538 two_stage_opamp_dummy_magic_0.VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 GNDA.t247 GNDA.t245 bgr_0.NFET_GATE_10uA.t4 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X540 two_stage_opamp_dummy_magic_0.VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 GNDA.t327 bgr_0.TAIL_CUR_MIR_BIAS.t25 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X542 two_stage_opamp_dummy_magic_0.V_err_gate.t0 bgr_0.NFET_GATE_10uA.t18 GNDA.t141 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X543 bgr_0.1st_Vout_1.t6 bgr_0.Vin+.t9 bgr_0.V_p_1.t1 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X544 VDDA.t456 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t343 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X545 VDDA.t363 VDDA.t361 VDDA.t363 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0 ps=0 w=3.2 l=0.2
X546 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t6 GNDA.t107 sky130_fd_pr__res_high_po_1p41 l=1.41
X547 bgr_0.V_TOP.t13 bgr_0.1st_Vout_1.t31 VDDA.t461 VDDA.t460 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X548 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X549 two_stage_opamp_dummy_magic_0.VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 two_stage_opamp_dummy_magic_0.VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 bgr_0.PFET_GATE_10uA.t24 VDDA.t431 VDDA.t430 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X552 two_stage_opamp_dummy_magic_0.VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_0.VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 bgr_0.Vin-.t6 bgr_0.V_TOP.t38 VDDA.t264 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X555 VDDA.t440 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 VDDA.t439 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X556 VDDA.t360 VDDA.t358 two_stage_opamp_dummy_magic_0.VD4.t35 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X557 two_stage_opamp_dummy_magic_0.VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 two_stage_opamp_dummy_magic_0.V_p.t10 bgr_0.TAIL_CUR_MIR_BIAS.t26 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X559 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.Vb2.t22 a_10480_8490.t8 two_stage_opamp_dummy_magic_0.VD4.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X560 two_stage_opamp_dummy_magic_0.VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 a_13790_17550.t0 GNDA.t106 GNDA.t105 sky130_fd_pr__res_xhigh_po_0p35 l=6
X562 two_stage_opamp_dummy_magic_0.VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 two_stage_opamp_dummy_magic_0.VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 bgr_0.V_TOP.t3 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X565 GNDA.t203 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X566 VDDA.t354 VDDA.t352 two_stage_opamp_dummy_magic_0.VD3.t36 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X567 two_stage_opamp_dummy_magic_0.VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 two_stage_opamp_dummy_magic_0.VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 two_stage_opamp_dummy_magic_0.VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 GNDA.t194 VDDA.t349 VDDA.t351 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X571 bgr_0.V_TOP.t39 VDDA.t262 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 two_stage_opamp_dummy_magic_0.VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 two_stage_opamp_dummy_magic_0.VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 bgr_0.NFET_GATE_10uA.t19 GNDA.t143 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X575 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 bgr_0.NFET_GATE_10uA.t20 GNDA.t137 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X576 two_stage_opamp_dummy_magic_0.VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 two_stage_opamp_dummy_magic_0.VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 VDDA.t64 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t3 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X580 VDDA.t348 VDDA.t346 two_stage_opamp_dummy_magic_0.err_amp_out.t5 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X581 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.VD1.t7 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X582 two_stage_opamp_dummy_magic_0.VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 bgr_0.V_TOP.t40 VDDA.t261 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 VDDA.t260 bgr_0.V_TOP.t41 bgr_0.Vin+.t1 VDDA.t259 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X585 VDDA.t345 VDDA.t343 GNDA.t193 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X586 two_stage_opamp_dummy_magic_0.VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 two_stage_opamp_dummy_magic_0.VD2.t20 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.X.t12 GNDA.t316 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X588 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.Vb2.t23 a_10480_8490.t7 two_stage_opamp_dummy_magic_0.VD4.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X589 bgr_0.V_mir1.t3 bgr_0.V_mir1.t2 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X590 two_stage_opamp_dummy_magic_0.VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 bgr_0.NFET_GATE_10uA.t21 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X592 a_8420_8490.t2 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X593 GNDA.t224 GNDA.t244 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X594 bgr_0.V_mir2.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 bgr_0.V_p_2.t1 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X595 bgr_0.PFET_GATE_10uA.t8 VDDA.t340 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X596 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 two_stage_opamp_dummy_magic_0.X.t35 GNDA.t88 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X597 two_stage_opamp_dummy_magic_0.VD2.t0 VIN+.t7 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X598 two_stage_opamp_dummy_magic_0.VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 two_stage_opamp_dummy_magic_0.VOUT-.t15 VDDA.t337 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X600 VDDA.t171 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X601 two_stage_opamp_dummy_magic_0.VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 GNDA.t157 bgr_0.TAIL_CUR_MIR_BIAS.t27 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X603 two_stage_opamp_dummy_magic_0.V_err_gate.t13 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X604 two_stage_opamp_dummy_magic_0.VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 VDDA.t336 VDDA.t334 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X606 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X607 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.Vb2.t25 a_10480_8490.t6 two_stage_opamp_dummy_magic_0.VD4.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X608 two_stage_opamp_dummy_magic_0.VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 bgr_0.V_TOP.t42 VDDA.t258 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 bgr_0.TAIL_CUR_MIR_BIAS.t2 bgr_0.PFET_GATE_10uA.t26 VDDA.t181 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X611 two_stage_opamp_dummy_magic_0.VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 two_stage_opamp_dummy_magic_0.VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X614 VDDA.t333 VDDA.t331 two_stage_opamp_dummy_magic_0.VOUT+.t14 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X615 two_stage_opamp_dummy_magic_0.VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 bgr_0.1st_Vout_2.t2 bgr_0.V_mir2.t21 VDDA.t58 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X617 two_stage_opamp_dummy_magic_0.VOUT+.t13 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t83 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X618 two_stage_opamp_dummy_magic_0.V_p.t8 bgr_0.TAIL_CUR_MIR_BIAS.t28 GNDA.t324 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X619 VDDA.t330 VDDA.t327 VDDA.t329 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X620 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 a_5350_5088.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X622 GNDA.t224 GNDA.t223 bgr_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X623 two_stage_opamp_dummy_magic_0.VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 GNDA.t133 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X625 two_stage_opamp_dummy_magic_0.VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_0.VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 VDDA.t10 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.VOUT-.t1 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X628 two_stage_opamp_dummy_magic_0.VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_0.VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 two_stage_opamp_dummy_magic_0.V_p.t7 bgr_0.TAIL_CUR_MIR_BIAS.t29 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X631 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 bgr_0.V_TOP.t43 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X632 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t324 VDDA.t326 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X634 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.Vb2.t26 a_10480_8490.t5 two_stage_opamp_dummy_magic_0.VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X635 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X636 two_stage_opamp_dummy_magic_0.V_err_p.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t132 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X637 two_stage_opamp_dummy_magic_0.VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 two_stage_opamp_dummy_magic_0.VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t6 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X640 two_stage_opamp_dummy_magic_0.VOUT+.t18 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA.t330 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X641 VDDA.t128 bgr_0.1st_Vout_2.t32 bgr_0.PFET_GATE_10uA.t2 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X642 VDDA.t323 VDDA.t321 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X643 two_stage_opamp_dummy_magic_0.VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t318 VDDA.t320 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X645 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X646 two_stage_opamp_dummy_magic_0.VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_0.Y.t36 GNDA.t336 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X648 two_stage_opamp_dummy_magic_0.VD2.t19 VIN+.t8 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X649 GNDA.t240 GNDA.t238 bgr_0.TAIL_CUR_MIR_BIAS.t10 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X650 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 two_stage_opamp_dummy_magic_0.VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 two_stage_opamp_dummy_magic_0.VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 two_stage_opamp_dummy_magic_0.VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 two_stage_opamp_dummy_magic_0.VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 bgr_0.V_mir1.t16 bgr_0.Vin-.t11 bgr_0.V_p_1.t6 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X657 two_stage_opamp_dummy_magic_0.VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 two_stage_opamp_dummy_magic_0.VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 two_stage_opamp_dummy_magic_0.VD2.t2 VIN+.t9 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X660 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t448 VDDA.t447 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X661 two_stage_opamp_dummy_magic_0.VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 two_stage_opamp_dummy_magic_0.X.t37 GNDA.t20 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X663 VDDA.t317 VDDA.t315 GNDA.t192 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X664 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 GNDA.t111 bgr_0.TAIL_CUR_MIR_BIAS.t30 two_stage_opamp_dummy_magic_0.V_p_mir.t1 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X666 two_stage_opamp_dummy_magic_0.V_err_gate.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X667 VDDA.t314 VDDA.t312 two_stage_opamp_dummy_magic_0.Vb2.t8 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X668 a_10480_8490.t4 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X669 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X670 VDDA.t455 two_stage_opamp_dummy_magic_0.Y.t37 two_stage_opamp_dummy_magic_0.VOUT+.t4 VDDA.t454 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X671 GNDA.t135 bgr_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X672 VDDA.t255 bgr_0.V_TOP.t44 bgr_0.START_UP.t2 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X673 two_stage_opamp_dummy_magic_0.VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.Vb2.t28 a_8420_8490.t1 two_stage_opamp_dummy_magic_0.VD3.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X675 two_stage_opamp_dummy_magic_0.VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 two_stage_opamp_dummy_magic_0.V_p.t6 bgr_0.TAIL_CUR_MIR_BIAS.t31 GNDA.t114 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X677 VDDA.t43 GNDA.t235 GNDA.t237 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X678 two_stage_opamp_dummy_magic_0.VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VDDA.t134 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X680 two_stage_opamp_dummy_magic_0.VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 GNDA.t224 GNDA.t234 bgr_0.Vbe2.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X682 two_stage_opamp_dummy_magic_0.VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 two_stage_opamp_dummy_magic_0.VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 VDDA.t122 two_stage_opamp_dummy_magic_0.X.t38 two_stage_opamp_dummy_magic_0.VOUT-.t9 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X685 VDDA.t311 VDDA.t309 two_stage_opamp_dummy_magic_0.VOUT-.t14 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X686 VDDA.t237 bgr_0.V_mir2.t2 bgr_0.V_mir2.t3 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X687 VDDA.t153 bgr_0.PFET_GATE_10uA.t27 bgr_0.TAIL_CUR_MIR_BIAS.t1 VDDA.t152 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X688 two_stage_opamp_dummy_magic_0.VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 GNDA.t233 GNDA.t231 VDDA.t218 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X691 bgr_0.TAIL_CUR_MIR_BIAS.t0 bgr_0.PFET_GATE_10uA.t28 VDDA.t429 VDDA.t428 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X692 two_stage_opamp_dummy_magic_0.VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 bgr_0.V_TOP.t45 VDDA.t253 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 two_stage_opamp_dummy_magic_0.V_err_p.t5 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t145 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X695 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t22 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X696 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X697 two_stage_opamp_dummy_magic_0.VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 two_stage_opamp_dummy_magic_0.V_err_p.t3 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X699 two_stage_opamp_dummy_magic_0.V_err_p.t19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X700 two_stage_opamp_dummy_magic_0.VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_0.Y.t38 GNDA.t345 VDDA.t462 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X702 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 bgr_0.1st_Vout_2.t8 bgr_0.V_CUR_REF_REG.t6 bgr_0.V_p_2.t8 GNDA.t318 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X704 bgr_0.V_TOP.t46 VDDA.t252 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.Vb2.t29 a_8420_8490.t0 two_stage_opamp_dummy_magic_0.VD3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X706 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_0.X.t39 VDDA.t123 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X707 two_stage_opamp_dummy_magic_0.V_p_mir.t3 VIN-.t8 bgr_0.TAIL_CUR_MIR_BIAS.t9 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X708 two_stage_opamp_dummy_magic_0.VD1.t1 VIN-.t9 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X709 two_stage_opamp_dummy_magic_0.VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 two_stage_opamp_dummy_magic_0.VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 two_stage_opamp_dummy_magic_0.VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 two_stage_opamp_dummy_magic_0.VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 bgr_0.V_p_1.t10 VDDA.t472 GNDA.t191 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X714 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 bgr_0.V_mir1.t14 bgr_0.Vin-.t12 bgr_0.V_p_1.t5 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X716 VDDA.t308 VDDA.t306 bgr_0.PFET_GATE_10uA.t7 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X717 two_stage_opamp_dummy_magic_0.VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 two_stage_opamp_dummy_magic_0.VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 GNDA.t172 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 two_stage_opamp_dummy_magic_0.VOUT-.t12 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X720 two_stage_opamp_dummy_magic_0.VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 two_stage_opamp_dummy_magic_0.VD1.t2 VIN-.t10 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X722 a_10480_8490.t3 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X723 bgr_0.V_TOP.t47 VDDA.t251 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VDDA.t226 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD3.t34 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X725 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 two_stage_opamp_dummy_magic_0.X.t40 GNDA.t43 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X726 VDDA.t130 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X727 two_stage_opamp_dummy_magic_0.VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 two_stage_opamp_dummy_magic_0.VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 GNDA.t54 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 two_stage_opamp_dummy_magic_0.VOUT+.t1 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X730 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 bgr_0.V_TOP.t48 VDDA.t250 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X731 bgr_0.V_TOP.t8 bgr_0.START_UP.t7 bgr_0.Vin-.t1 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X732 two_stage_opamp_dummy_magic_0.V_err_gate.t8 VDDA.t303 VDDA.t305 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X733 two_stage_opamp_dummy_magic_0.VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 bgr_0.1st_Vout_2.t7 bgr_0.V_CUR_REF_REG.t7 bgr_0.V_p_2.t7 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X735 two_stage_opamp_dummy_magic_0.V_err_gate.t12 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X736 two_stage_opamp_dummy_magic_0.VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VDDA.t100 bgr_0.1st_Vout_2.t36 bgr_0.PFET_GATE_10uA.t1 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X738 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X740 two_stage_opamp_dummy_magic_0.Vb2.t1 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X741 VDDA.t419 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.VOUT+.t3 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X742 two_stage_opamp_dummy_magic_0.VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 a_5230_5088.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t104 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X744 two_stage_opamp_dummy_magic_0.VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 two_stage_opamp_dummy_magic_0.VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 GNDA.t230 GNDA.t228 two_stage_opamp_dummy_magic_0.VOUT-.t16 GNDA.t229 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X747 two_stage_opamp_dummy_magic_0.VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_0.VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 two_stage_opamp_dummy_magic_0.VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 two_stage_opamp_dummy_magic_0.VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VDDA.t147 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t4 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X752 a_8420_8490.t10 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.VD3.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X753 two_stage_opamp_dummy_magic_0.VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_0.VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VDDA.t302 VDDA.t300 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X756 two_stage_opamp_dummy_magic_0.VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 bgr_0.PFET_GATE_10uA.t29 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X758 a_10480_8490.t2 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.VD4.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X759 two_stage_opamp_dummy_magic_0.VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VDDA.t60 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t1 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X761 VDDA.t51 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.VOUT-.t5 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X762 two_stage_opamp_dummy_magic_0.VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 two_stage_opamp_dummy_magic_0.VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 two_stage_opamp_dummy_magic_0.Y.t40 VDDA.t467 GNDA.t346 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X765 two_stage_opamp_dummy_magic_0.VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X767 two_stage_opamp_dummy_magic_0.VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 two_stage_opamp_dummy_magic_0.Y.t4 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD1.t4 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X769 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X770 GNDA.t201 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X771 two_stage_opamp_dummy_magic_0.VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_0.Y.t41 GNDA.t180 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X773 two_stage_opamp_dummy_magic_0.VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 two_stage_opamp_dummy_magic_0.VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 two_stage_opamp_dummy_magic_0.VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t42 GNDA.t163 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X777 two_stage_opamp_dummy_magic_0.VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 bgr_0.V_TOP.t49 VDDA.t248 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 bgr_0.1st_Vout_1.t0 bgr_0.Vin+.t10 bgr_0.V_p_1.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X780 GNDA.t334 two_stage_opamp_dummy_magic_0.err_amp_out.t12 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA.t333 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X781 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA.t225 GNDA.t227 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X782 two_stage_opamp_dummy_magic_0.VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 two_stage_opamp_dummy_magic_0.X.t42 VDDA.t2 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X784 GNDA.t222 GNDA.t220 VDDA.t247 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X785 two_stage_opamp_dummy_magic_0.VD2.t21 VIN+.t10 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA.t344 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X786 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_5750_2276.t0 GNDA.t337 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X787 bgr_0.Vin+.t5 bgr_0.Vbe2.t8 GNDA.t328 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X788 VDDA.t80 two_stage_opamp_dummy_magic_0.Vb3.t28 two_stage_opamp_dummy_magic_0.VD4.t8 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X789 two_stage_opamp_dummy_magic_0.VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.V_TOP.n0 bgr_0.V_TOP.t43 369.534
R1 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 339.961
R2 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 339.272
R3 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R4 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R5 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R6 bgr_0.V_TOP.n12 bgr_0.V_TOP.n8 334.772
R7 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R8 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R9 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R10 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R11 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R12 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R13 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R14 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R15 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R16 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R17 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R18 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R19 bgr_0.V_TOP bgr_0.V_TOP.t32 214.222
R20 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R21 bgr_0.V_TOP.n7 bgr_0.V_TOP.t6 176.114
R22 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R23 bgr_0.V_TOP.n27 bgr_0.V_TOP.t31 144.601
R24 bgr_0.V_TOP.n26 bgr_0.V_TOP.t44 144.601
R25 bgr_0.V_TOP.n25 bgr_0.V_TOP.t18 144.601
R26 bgr_0.V_TOP.n24 bgr_0.V_TOP.t26 144.601
R27 bgr_0.V_TOP.n23 bgr_0.V_TOP.t37 144.601
R28 bgr_0.V_TOP.n22 bgr_0.V_TOP.t35 144.601
R29 bgr_0.V_TOP.n21 bgr_0.V_TOP.t48 144.601
R30 bgr_0.V_TOP.n20 bgr_0.V_TOP.t20 144.601
R31 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 144.601
R32 bgr_0.V_TOP.n1 bgr_0.V_TOP.t23 144.601
R33 bgr_0.V_TOP.n2 bgr_0.V_TOP.t14 144.601
R34 bgr_0.V_TOP.n3 bgr_0.V_TOP.t38 144.601
R35 bgr_0.V_TOP.n4 bgr_0.V_TOP.t41 144.601
R36 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R37 bgr_0.V_TOP.n18 bgr_0.V_TOP.t2 95.4466
R38 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R39 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R40 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R41 bgr_0.V_TOP.n6 bgr_0.V_TOP.t11 39.4005
R42 bgr_0.V_TOP.n6 bgr_0.V_TOP.t12 39.4005
R43 bgr_0.V_TOP.n8 bgr_0.V_TOP.t1 39.4005
R44 bgr_0.V_TOP.n8 bgr_0.V_TOP.t13 39.4005
R45 bgr_0.V_TOP.n10 bgr_0.V_TOP.t5 39.4005
R46 bgr_0.V_TOP.n10 bgr_0.V_TOP.t0 39.4005
R47 bgr_0.V_TOP.n9 bgr_0.V_TOP.t4 39.4005
R48 bgr_0.V_TOP.n9 bgr_0.V_TOP.t8 39.4005
R49 bgr_0.V_TOP.n14 bgr_0.V_TOP.t9 39.4005
R50 bgr_0.V_TOP.n14 bgr_0.V_TOP.t10 39.4005
R51 bgr_0.V_TOP.n16 bgr_0.V_TOP.t7 39.4005
R52 bgr_0.V_TOP.n16 bgr_0.V_TOP.t3 39.4005
R53 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 8.313
R54 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R55 bgr_0.V_TOP.n28 bgr_0.V_TOP.t49 4.8295
R56 bgr_0.V_TOP.n29 bgr_0.V_TOP.t25 4.8295
R57 bgr_0.V_TOP.n31 bgr_0.V_TOP.t21 4.8295
R58 bgr_0.V_TOP.n32 bgr_0.V_TOP.t34 4.8295
R59 bgr_0.V_TOP.n34 bgr_0.V_TOP.t30 4.8295
R60 bgr_0.V_TOP.n35 bgr_0.V_TOP.t46 4.8295
R61 bgr_0.V_TOP.n37 bgr_0.V_TOP.t24 4.8295
R62 bgr_0.V_TOP.n28 bgr_0.V_TOP.t39 4.5005
R63 bgr_0.V_TOP.n30 bgr_0.V_TOP.t28 4.5005
R64 bgr_0.V_TOP.n29 bgr_0.V_TOP.t33 4.5005
R65 bgr_0.V_TOP.n31 bgr_0.V_TOP.t15 4.5005
R66 bgr_0.V_TOP.n33 bgr_0.V_TOP.t40 4.5005
R67 bgr_0.V_TOP.n32 bgr_0.V_TOP.t45 4.5005
R68 bgr_0.V_TOP.n34 bgr_0.V_TOP.t22 4.5005
R69 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 4.5005
R70 bgr_0.V_TOP.n35 bgr_0.V_TOP.t19 4.5005
R71 bgr_0.V_TOP.n37 bgr_0.V_TOP.t17 4.5005
R72 bgr_0.V_TOP.n38 bgr_0.V_TOP.t42 4.5005
R73 bgr_0.V_TOP.n39 bgr_0.V_TOP.t47 4.5005
R74 bgr_0.V_TOP.n40 bgr_0.V_TOP.t36 4.5005
R75 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R76 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R77 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R78 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R79 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R80 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R81 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R82 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R83 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R84 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R85 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R86 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R87 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R88 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R89 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R90 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R91 bgr_0.Vin-.n21 bgr_0.Vin-.n20 1850.93
R92 bgr_0.Vin-.n9 bgr_0.Vin-.t10 688.859
R93 bgr_0.Vin-.n11 bgr_0.Vin-.n10 514.134
R94 bgr_0.Vin-.n7 bgr_0.Vin-.n6 345.115
R95 bgr_0.Vin-.n13 bgr_0.Vin-.n12 214.713
R96 bgr_0.Vin-.n9 bgr_0.Vin-.t12 174.726
R97 bgr_0.Vin-.n10 bgr_0.Vin-.t8 174.726
R98 bgr_0.Vin-.n11 bgr_0.Vin-.t11 174.726
R99 bgr_0.Vin-.n12 bgr_0.Vin-.t9 174.726
R100 bgr_0.Vin-.n5 bgr_0.Vin-.n3 173.029
R101 bgr_0.Vin-.n5 bgr_0.Vin-.n4 168.654
R102 bgr_0.Vin-.n7 bgr_0.Vin-.t7 162.921
R103 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R104 bgr_0.Vin-.n12 bgr_0.Vin-.n11 128.534
R105 bgr_0.Vin-.n22 bgr_0.Vin-.n21 84.0884
R106 bgr_0.Vin-.n17 bgr_0.Vin-.n16 83.5719
R107 bgr_0.Vin-.n18 bgr_0.Vin-.n0 83.5719
R108 bgr_0.Vin-.n19 bgr_0.Vin-.n1 83.5719
R109 bgr_0.Vin-.n14 bgr_0.Vin-.t2 65.0299
R110 bgr_0.Vin-.n6 bgr_0.Vin-.t1 39.4005
R111 bgr_0.Vin-.n6 bgr_0.Vin-.t0 39.4005
R112 bgr_0.Vin-.n18 bgr_0.Vin-.n17 26.074
R113 bgr_0.Vin-.n19 bgr_0.Vin-.n18 26.074
R114 bgr_0.Vin-.n21 bgr_0.Vin-.n19 26.074
R115 bgr_0.Vin-.n23 bgr_0.Vin-.n13 17.526
R116 bgr_0.Vin-.n4 bgr_0.Vin-.t3 13.1338
R117 bgr_0.Vin-.n4 bgr_0.Vin-.t6 13.1338
R118 bgr_0.Vin-.n3 bgr_0.Vin-.t5 13.1338
R119 bgr_0.Vin-.n3 bgr_0.Vin-.t4 13.1338
R120 bgr_0.Vin-.n13 bgr_0.Vin-.n8 12.5317
R121 bgr_0.Vin-.n8 bgr_0.Vin-.n7 6.40675
R122 bgr_0.Vin-.n8 bgr_0.Vin-.n5 3.8755
R123 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56363
R124 bgr_0.Vin-.n23 bgr_0.Vin-.n22 1.5505
R125 bgr_0.Vin-.n25 bgr_0.Vin-.n24 1.5505
R126 bgr_0.Vin-.n15 bgr_0.Vin-.n2 1.5505
R127 bgr_0.Vin-.n22 bgr_0.Vin-.n1 1.14402
R128 bgr_0.Vin-.n15 bgr_0.Vin-.n0 0.885803
R129 bgr_0.Vin-.n16 bgr_0.Vin-.n15 0.77514
R130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.756696
R131 bgr_0.Vin-.n25 bgr_0.Vin-.n1 0.701365
R132 bgr_0.Vin-.n14 bgr_0.Vin-.n2 0.537712
R133 bgr_0.Vin-.n17 bgr_0.Vin-.t2 0.290206
R134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n25 0.203382
R135 bgr_0.Vin-.n24 bgr_0.Vin-.n2 0.0183571
R136 bgr_0.Vin-.n24 bgr_0.Vin-.n23 0.0183571
R137 VDDA.n376 VDDA.n343 6600
R138 VDDA.n378 VDDA.n343 6600
R139 VDDA.n378 VDDA.n344 6570
R140 VDDA.n376 VDDA.n344 6570
R141 VDDA.n331 VDDA.n266 4710
R142 VDDA.n331 VDDA.n267 4710
R143 VDDA.n333 VDDA.n266 4710
R144 VDDA.n333 VDDA.n267 4710
R145 VDDA.n289 VDDA.n288 4710
R146 VDDA.n291 VDDA.n288 4710
R147 VDDA.n289 VDDA.n282 4710
R148 VDDA.n291 VDDA.n282 4710
R149 VDDA.n143 VDDA.n129 4605
R150 VDDA.n145 VDDA.n129 4605
R151 VDDA.n69 VDDA.n65 4605
R152 VDDA.n69 VDDA.n66 4605
R153 VDDA.n179 VDDA.n175 4590
R154 VDDA.n179 VDDA.n176 4590
R155 VDDA.n181 VDDA.n176 4590
R156 VDDA.n181 VDDA.n175 4590
R157 VDDA.n143 VDDA.n130 4575
R158 VDDA.n145 VDDA.n130 4575
R159 VDDA.n71 VDDA.n65 4575
R160 VDDA.n71 VDDA.n66 4575
R161 VDDA.n205 VDDA.n198 4020
R162 VDDA.n207 VDDA.n198 4020
R163 VDDA.n205 VDDA.n204 4020
R164 VDDA.n207 VDDA.n204 4020
R165 VDDA.n93 VDDA.n86 4020
R166 VDDA.n95 VDDA.n86 4020
R167 VDDA.n93 VDDA.n92 4020
R168 VDDA.n95 VDDA.n92 4020
R169 VDDA.n442 VDDA.n410 3420
R170 VDDA.n442 VDDA.n411 3420
R171 VDDA.n122 VDDA.n115 3390
R172 VDDA.n124 VDDA.n115 3390
R173 VDDA.n122 VDDA.n121 3390
R174 VDDA.n124 VDDA.n121 3390
R175 VDDA.n49 VDDA.n42 3390
R176 VDDA.n51 VDDA.n42 3390
R177 VDDA.n49 VDDA.n48 3390
R178 VDDA.n51 VDDA.n48 3390
R179 VDDA.n23 VDDA.n17 2940
R180 VDDA.n25 VDDA.n17 2940
R181 VDDA.n25 VDDA.n22 2940
R182 VDDA.n23 VDDA.n22 2940
R183 VDDA.n31 VDDA.n12 2940
R184 VDDA.n33 VDDA.n12 2940
R185 VDDA.n33 VDDA.n30 2940
R186 VDDA.n31 VDDA.n30 2940
R187 VDDA.n444 VDDA.n410 2760
R188 VDDA.n444 VDDA.n411 2760
R189 VDDA.n235 VDDA.n224 2415
R190 VDDA.n235 VDDA.n225 2370
R191 VDDA.n232 VDDA.n225 2280
R192 VDDA.n232 VDDA.n224 2235
R193 VDDA.n458 VDDA.n404 2145
R194 VDDA.n458 VDDA.n405 2100
R195 VDDA.n455 VDDA.n405 2100
R196 VDDA.n423 VDDA.n416 2100
R197 VDDA.n425 VDDA.n416 2100
R198 VDDA.n425 VDDA.n417 2100
R199 VDDA.n423 VDDA.n417 2100
R200 VDDA.n455 VDDA.n404 2055
R201 VDDA.n391 VDDA.n389 1770
R202 VDDA.n393 VDDA.n389 1770
R203 VDDA.n391 VDDA.n386 1770
R204 VDDA.n393 VDDA.n386 1770
R205 VDDA.n352 VDDA.n350 1770
R206 VDDA.n354 VDDA.n350 1770
R207 VDDA.n352 VDDA.n347 1770
R208 VDDA.n354 VDDA.n347 1770
R209 VDDA.n247 VDDA.n220 1575
R210 VDDA.n246 VDDA.n220 1575
R211 VDDA.n246 VDDA.n219 1545
R212 VDDA.n247 VDDA.n219 1545
R213 VDDA.n140 VDDA.t331 1216.42
R214 VDDA.n148 VDDA.t364 1216.42
R215 VDDA.n63 VDDA.t337 1216.42
R216 VDDA.n74 VDDA.t309 1216.42
R217 VDDA.n375 VDDA.n342 704
R218 VDDA.n379 VDDA.n342 704
R219 VDDA.n19 VDDA.t348 689.4
R220 VDDA.n18 VDDA.t375 689.4
R221 VDDA.n14 VDDA.t414 689.4
R222 VDDA.n13 VDDA.t305 689.4
R223 VDDA.n172 VDDA.t390 663.801
R224 VDDA.n185 VDDA.t396 663.801
R225 VDDA.n201 VDDA.t352 660.109
R226 VDDA.n199 VDDA.t379 660.109
R227 VDDA.n89 VDDA.t358 660.109
R228 VDDA.n87 VDDA.t403 660.109
R229 VDDA.n242 VDDA.t314 647.54
R230 VDDA.n251 VDDA.t330 647.54
R231 VDDA.n216 VDDA.n215 633.361
R232 VDDA.n152 VDDA.n151 626.534
R233 VDDA.n155 VDDA.n154 626.534
R234 VDDA.n157 VDDA.n156 626.534
R235 VDDA.n159 VDDA.n158 626.534
R236 VDDA.n161 VDDA.n160 626.534
R237 VDDA.n163 VDDA.n162 626.534
R238 VDDA.n165 VDDA.n164 626.534
R239 VDDA.n167 VDDA.n166 626.534
R240 VDDA.n169 VDDA.n168 626.534
R241 VDDA.n171 VDDA.n170 626.534
R242 VDDA.n229 VDDA.t361 623.958
R243 VDDA.n238 VDDA.t382 623.958
R244 VDDA.t361 VDDA.n228 615.926
R245 VDDA.n118 VDDA.t343 573.75
R246 VDDA.n116 VDDA.t370 573.75
R247 VDDA.n45 VDDA.t315 573.75
R248 VDDA.n43 VDDA.t349 573.75
R249 VDDA.n374 VDDA.n341 518.4
R250 VDDA.n380 VDDA.n341 518.4
R251 VDDA.n293 VDDA.n292 496
R252 VDDA.n293 VDDA.n281 496
R253 VDDA.n146 VDDA.n128 491.2
R254 VDDA.n142 VDDA.n128 491.2
R255 VDDA.n68 VDDA.n40 491.2
R256 VDDA.n68 VDDA.n67 491.2
R257 VDDA.n178 VDDA.n153 489.601
R258 VDDA.n178 VDDA.n177 489.601
R259 VDDA.n209 VDDA.n208 428.8
R260 VDDA.n209 VDDA.n197 428.8
R261 VDDA.n97 VDDA.n96 428.8
R262 VDDA.n97 VDDA.n85 428.8
R263 VDDA.n387 VDDA.t318 419.108
R264 VDDA.n384 VDDA.t321 419.108
R265 VDDA.n348 VDDA.t397 413.084
R266 VDDA.n345 VDDA.t376 413.084
R267 VDDA.n452 VDDA.t385 409.067
R268 VDDA.n461 VDDA.t324 409.067
R269 VDDA.n439 VDDA.t406 409.067
R270 VDDA.n447 VDDA.t400 409.067
R271 VDDA.n420 VDDA.t300 409.067
R272 VDDA.n428 VDDA.t367 390.322
R273 VDDA.t395 VDDA.n175 389.375
R274 VDDA.t389 VDDA.n176 389.375
R275 VDDA.t413 VDDA.n30 389.375
R276 VDDA.t304 VDDA.n12 389.375
R277 VDDA.n387 VDDA.t320 389.185
R278 VDDA.n384 VDDA.t323 389.185
R279 VDDA.n183 VDDA.n182 387.2
R280 VDDA.n182 VDDA.n174 387.2
R281 VDDA.n439 VDDA.t408 387.051
R282 VDDA.n447 VDDA.t402 387.051
R283 VDDA.n264 VDDA.t342 384.918
R284 VDDA.n268 VDDA.t308 384.918
R285 VDDA.n283 VDDA.t357 384.918
R286 VDDA.n285 VDDA.t411 384.918
R287 VDDA.n348 VDDA.t399 384.918
R288 VDDA.n345 VDDA.t378 384.918
R289 VDDA.t347 VDDA.n22 384.168
R290 VDDA.t374 VDDA.n17 384.168
R291 VDDA.n270 VDDA.n269 384
R292 VDDA.n269 VDDA.n265 384
R293 VDDA.n287 VDDA.n286 384
R294 VDDA.n287 VDDA.n284 384
R295 VDDA.n420 VDDA.t302 370.728
R296 VDDA.n428 VDDA.t369 370.728
R297 VDDA.n452 VDDA.t387 370.3
R298 VDDA.n461 VDDA.t326 370.3
R299 VDDA.n441 VDDA.n409 364.8
R300 VDDA.n373 VDDA.t334 360.868
R301 VDDA.n381 VDDA.t391 360.868
R302 VDDA.n264 VDDA.t340 358.858
R303 VDDA.n268 VDDA.t306 358.858
R304 VDDA.n283 VDDA.t355 358.858
R305 VDDA.n285 VDDA.t409 358.858
R306 VDDA.n126 VDDA.n125 355.2
R307 VDDA.n126 VDDA.n114 355.2
R308 VDDA.n53 VDDA.n52 355.2
R309 VDDA.n53 VDDA.n41 355.2
R310 VDDA.t307 VDDA.n331 351.591
R311 VDDA.n333 VDDA.t341 351.591
R312 VDDA.t410 VDDA.n289 351.591
R313 VDDA.n291 VDDA.t356 351.591
R314 VDDA.t313 VDDA.n246 346.668
R315 VDDA.n247 VDDA.t328 346.668
R316 VDDA.n413 VDDA.n412 345.127
R317 VDDA.n419 VDDA.n418 345.127
R318 VDDA.n401 VDDA.n400 344.7
R319 VDDA.n450 VDDA.n449 344.7
R320 VDDA.t322 VDDA.n391 344.394
R321 VDDA.n393 VDDA.t319 344.394
R322 VDDA.t377 VDDA.n352 344.394
R323 VDDA.n354 VDDA.t398 344.394
R324 VDDA.t386 VDDA.n455 344.394
R325 VDDA.n458 VDDA.t325 344.394
R326 VDDA.n275 VDDA.n273 342.3
R327 VDDA.n303 VDDA.n302 341.675
R328 VDDA.n301 VDDA.n300 341.675
R329 VDDA.n299 VDDA.n298 341.675
R330 VDDA.n297 VDDA.n296 341.675
R331 VDDA.n279 VDDA.n278 341.675
R332 VDDA.n277 VDDA.n276 341.675
R333 VDDA.n275 VDDA.n274 341.675
R334 VDDA.t407 VDDA.n442 340.635
R335 VDDA.n444 VDDA.t401 340.635
R336 VDDA.t301 VDDA.n423 340.635
R337 VDDA.n425 VDDA.t368 340.635
R338 VDDA.n407 VDDA.n406 339.272
R339 VDDA.n431 VDDA.n430 339.272
R340 VDDA.n433 VDDA.n432 339.272
R341 VDDA.n435 VDDA.n434 339.272
R342 VDDA.n437 VDDA.n436 339.272
R343 VDDA.n336 VDDA.n260 337.175
R344 VDDA.n262 VDDA.n261 337.175
R345 VDDA.n312 VDDA.n311 337.175
R346 VDDA.n315 VDDA.n309 337.175
R347 VDDA.n307 VDDA.n306 337.175
R348 VDDA.n319 VDDA.n318 337.175
R349 VDDA.n322 VDDA.n305 337.175
R350 VDDA.n325 VDDA.n324 337.175
R351 VDDA.n328 VDDA.n272 337.175
R352 VDDA.n294 VDDA.n280 337.175
R353 VDDA.n397 VDDA.n383 335.022
R354 VDDA.n173 VDDA.t388 332.75
R355 VDDA.n184 VDDA.t394 332.75
R356 VDDA.n19 VDDA.t346 332.75
R357 VDDA.n18 VDDA.t373 332.75
R358 VDDA.n14 VDDA.t412 332.75
R359 VDDA.n13 VDDA.t303 332.75
R360 VDDA.n243 VDDA.t312 314.274
R361 VDDA.n250 VDDA.t327 314.274
R362 VDDA.n21 VDDA.n16 313.601
R363 VDDA.n28 VDDA.n16 307.2
R364 VDDA.n36 VDDA.n11 307.2
R365 VDDA.n29 VDDA.n11 307.2
R366 VDDA.n445 VDDA.n409 294.401
R367 VDDA.t344 VDDA.n122 285.815
R368 VDDA.n124 VDDA.t371 285.815
R369 VDDA.t316 VDDA.n49 285.815
R370 VDDA.n51 VDDA.t350 285.815
R371 VDDA.t335 VDDA.n376 278.95
R372 VDDA.n378 VDDA.t392 278.95
R373 VDDA.n118 VDDA.t345 277.916
R374 VDDA.n116 VDDA.t372 277.916
R375 VDDA.n45 VDDA.t317 277.916
R376 VDDA.n43 VDDA.t351 277.916
R377 VDDA.n147 VDDA.n146 276.8
R378 VDDA.n142 VDDA.n141 276.8
R379 VDDA.n73 VDDA.n40 276.8
R380 VDDA.n67 VDDA.n64 276.8
R381 VDDA.n373 VDDA.t336 270.705
R382 VDDA.n381 VDDA.t393 270.705
R383 VDDA.n236 VDDA.n223 257.601
R384 VDDA.n440 VDDA.n408 246.4
R385 VDDA.t353 VDDA.n205 239.915
R386 VDDA.n207 VDDA.t380 239.915
R387 VDDA.t359 VDDA.n93 239.915
R388 VDDA.n95 VDDA.t404 239.915
R389 VDDA.n231 VDDA.n223 238.4
R390 VDDA.n203 VDDA.n202 230.4
R391 VDDA.n203 VDDA.n200 230.4
R392 VDDA.n91 VDDA.n90 230.4
R393 VDDA.n91 VDDA.n88 230.4
R394 VDDA.n459 VDDA.n403 228.8
R395 VDDA.n422 VDDA.n415 224
R396 VDDA.n426 VDDA.n415 224
R397 VDDA.n454 VDDA.n403 219.201
R398 VDDA.n120 VDDA.n119 211.201
R399 VDDA.n120 VDDA.n117 211.201
R400 VDDA.n47 VDDA.n46 211.201
R401 VDDA.n47 VDDA.n44 211.201
R402 VDDA.n26 VDDA.n20 211.201
R403 VDDA.n27 VDDA.n26 211.201
R404 VDDA.n35 VDDA.n34 211.201
R405 VDDA.n141 VDDA.n127 204.8
R406 VDDA.n147 VDDA.n127 204.8
R407 VDDA.n73 VDDA.n72 204.8
R408 VDDA.n72 VDDA.n64 204.8
R409 VDDA.n34 VDDA.n15 202.971
R410 VDDA.n208 VDDA.n200 198.4
R411 VDDA.n202 VDDA.n197 198.4
R412 VDDA.n96 VDDA.n88 198.4
R413 VDDA.n90 VDDA.n85 198.4
R414 VDDA.n231 VDDA.n230 192
R415 VDDA.t68 VDDA.t313 190
R416 VDDA.t328 VDDA.t68 190
R417 VDDA.n237 VDDA.n236 188.8
R418 VDDA.n335 VDDA.n334 188.8
R419 VDDA.n330 VDDA.n329 188.8
R420 VDDA.n394 VDDA.n388 188.8
R421 VDDA.n390 VDDA.n388 188.8
R422 VDDA.n355 VDDA.n349 188.8
R423 VDDA.n351 VDDA.n349 188.8
R424 VDDA.t131 VDDA.t395 186.607
R425 VDDA.t167 VDDA.t131 186.607
R426 VDDA.t94 VDDA.t167 186.607
R427 VDDA.t165 VDDA.t94 186.607
R428 VDDA.t144 VDDA.t165 186.607
R429 VDDA.t137 VDDA.t144 186.607
R430 VDDA.t159 VDDA.t137 186.607
R431 VDDA.t150 VDDA.t159 186.607
R432 VDDA.t12 VDDA.t150 186.607
R433 VDDA.t163 VDDA.t12 186.607
R434 VDDA.t90 VDDA.t92 186.607
R435 VDDA.t92 VDDA.t14 186.607
R436 VDDA.t14 VDDA.t133 186.607
R437 VDDA.t133 VDDA.t135 186.607
R438 VDDA.t135 VDDA.t146 186.607
R439 VDDA.t146 VDDA.t148 186.607
R440 VDDA.t148 VDDA.t70 186.607
R441 VDDA.t70 VDDA.t161 186.607
R442 VDDA.t161 VDDA.t88 186.607
R443 VDDA.t88 VDDA.t389 186.607
R444 VDDA.t215 VDDA.t413 186.607
R445 VDDA.t416 VDDA.t215 186.607
R446 VDDA.t436 VDDA.t416 186.607
R447 VDDA.t216 VDDA.t436 186.607
R448 VDDA.t75 VDDA.t216 186.607
R449 VDDA.t212 VDDA.t457 186.607
R450 VDDA.t457 VDDA.t7 186.607
R451 VDDA.t7 VDDA.t46 186.607
R452 VDDA.t46 VDDA.t415 186.607
R453 VDDA.t415 VDDA.t304 186.607
R454 VDDA.t55 VDDA.t347 183.333
R455 VDDA.t87 VDDA.t55 183.333
R456 VDDA.t81 VDDA.t87 183.333
R457 VDDA.t82 VDDA.t81 183.333
R458 VDDA.t8 VDDA.t82 183.333
R459 VDDA.t102 VDDA.t139 183.333
R460 VDDA.t139 VDDA.t83 183.333
R461 VDDA.t83 VDDA.t118 183.333
R462 VDDA.t118 VDDA.t56 183.333
R463 VDDA.t56 VDDA.t374 183.333
R464 VDDA.n375 VDDA.n374 182.4
R465 VDDA.n380 VDDA.n379 182.4
R466 VDDA.n139 VDDA.t333 178.124
R467 VDDA.n149 VDDA.t366 178.124
R468 VDDA.n62 VDDA.t339 178.124
R469 VDDA.n75 VDDA.t311 178.124
R470 VDDA.n446 VDDA.n408 176
R471 VDDA.n226 VDDA.n221 174.393
R472 VDDA.t178 VDDA.t307 172.727
R473 VDDA.t63 VDDA.t178 172.727
R474 VDDA.t174 VDDA.t63 172.727
R475 VDDA.t236 VDDA.t174 172.727
R476 VDDA.t240 VDDA.t236 172.727
R477 VDDA.t127 VDDA.t240 172.727
R478 VDDA.t39 VDDA.t127 172.727
R479 VDDA.t59 VDDA.t39 172.727
R480 VDDA.t61 VDDA.t59 172.727
R481 VDDA.t107 VDDA.t192 172.727
R482 VDDA.t99 VDDA.t107 172.727
R483 VDDA.t202 VDDA.t99 172.727
R484 VDDA.t172 VDDA.t202 172.727
R485 VDDA.t57 VDDA.t172 172.727
R486 VDDA.t85 VDDA.t57 172.727
R487 VDDA.t238 VDDA.t85 172.727
R488 VDDA.t210 VDDA.t238 172.727
R489 VDDA.t341 VDDA.t210 172.727
R490 VDDA.t458 VDDA.t410 172.727
R491 VDDA.t35 VDDA.t458 172.727
R492 VDDA.t426 VDDA.t35 172.727
R493 VDDA.t434 VDDA.t426 172.727
R494 VDDA.t184 VDDA.t434 172.727
R495 VDDA.t25 VDDA.t184 172.727
R496 VDDA.t460 VDDA.t25 172.727
R497 VDDA.t129 VDDA.t460 172.727
R498 VDDA.t156 VDDA.t129 172.727
R499 VDDA.t186 VDDA.t443 172.727
R500 VDDA.t420 VDDA.t186 172.727
R501 VDDA.t422 VDDA.t420 172.727
R502 VDDA.t198 VDDA.t422 172.727
R503 VDDA.t142 VDDA.t198 172.727
R504 VDDA.t445 VDDA.t142 172.727
R505 VDDA.t109 VDDA.t445 172.727
R506 VDDA.t206 VDDA.t109 172.727
R507 VDDA.t356 VDDA.t206 172.727
R508 VDDA.t362 VDDA.n232 172.554
R509 VDDA.n235 VDDA.t383 172.554
R510 VDDA.n340 VDDA.n339 168.435
R511 VDDA.n359 VDDA.n358 168.435
R512 VDDA.n361 VDDA.n360 168.435
R513 VDDA.n363 VDDA.n362 168.435
R514 VDDA.n365 VDDA.n364 168.435
R515 VDDA.n367 VDDA.n366 168.435
R516 VDDA.n369 VDDA.n368 168.435
R517 VDDA.n371 VDDA.n370 168.435
R518 VDDA.n245 VDDA.n218 164.8
R519 VDDA.n248 VDDA.n218 164.8
R520 VDDA.t332 VDDA.n143 161.817
R521 VDDA.n145 VDDA.t365 161.817
R522 VDDA.t310 VDDA.n65 161.817
R523 VDDA.t338 VDDA.n66 161.817
R524 VDDA.n195 VDDA.n193 160.428
R525 VDDA.n192 VDDA.n190 160.428
R526 VDDA.n83 VDDA.n81 160.428
R527 VDDA.n80 VDDA.n78 160.428
R528 VDDA.t256 VDDA.t335 159.814
R529 VDDA.t277 VDDA.t256 159.814
R530 VDDA.t288 VDDA.t277 159.814
R531 VDDA.t298 VDDA.t288 159.814
R532 VDDA.t263 VDDA.t298 159.814
R533 VDDA.t259 VDDA.t263 159.814
R534 VDDA.t282 VDDA.t259 159.814
R535 VDDA.t290 VDDA.t282 159.814
R536 VDDA.t268 VDDA.t249 159.814
R537 VDDA.t265 VDDA.t268 159.814
R538 VDDA.t284 VDDA.t265 159.814
R539 VDDA.t293 VDDA.t284 159.814
R540 VDDA.t254 VDDA.t293 159.814
R541 VDDA.t274 VDDA.t254 159.814
R542 VDDA.t272 VDDA.t274 159.814
R543 VDDA.t392 VDDA.t272 159.814
R544 VDDA.n195 VDDA.n194 159.803
R545 VDDA.n192 VDDA.n191 159.803
R546 VDDA.n83 VDDA.n82 159.803
R547 VDDA.n80 VDDA.n79 159.803
R548 VDDA.t65 VDDA.t322 158.333
R549 VDDA.t319 VDDA.t432 158.333
R550 VDDA.t214 VDDA.t377 158.333
R551 VDDA.t398 VDDA.t103 158.333
R552 VDDA.t430 VDDA.t386 158.333
R553 VDDA.t96 VDDA.t430 158.333
R554 VDDA.t439 VDDA.t196 158.333
R555 VDDA.t325 VDDA.t439 158.333
R556 VDDA.t33 VDDA.t407 155.97
R557 VDDA.t450 VDDA.t33 155.97
R558 VDDA.t180 VDDA.t450 155.97
R559 VDDA.t31 VDDA.t180 155.97
R560 VDDA.t47 VDDA.t31 155.97
R561 VDDA.t152 VDDA.t47 155.97
R562 VDDA.t441 VDDA.t140 155.97
R563 VDDA.t428 VDDA.t441 155.97
R564 VDDA.t154 VDDA.t428 155.97
R565 VDDA.t401 VDDA.t154 155.97
R566 VDDA.t424 VDDA.t301 155.97
R567 VDDA.t182 VDDA.t424 155.97
R568 VDDA.t29 VDDA.t27 155.97
R569 VDDA.t368 VDDA.t29 155.97
R570 VDDA.n201 VDDA.t354 155.125
R571 VDDA.n199 VDDA.t381 155.125
R572 VDDA.n89 VDDA.t360 155.125
R573 VDDA.n87 VDDA.t405 155.125
R574 VDDA.n139 VDDA.n138 151.882
R575 VDDA.n62 VDDA.n61 151.882
R576 VDDA.n150 VDDA.n149 151.321
R577 VDDA.n76 VDDA.n75 151.321
R578 VDDA.n125 VDDA.n117 150.4
R579 VDDA.n119 VDDA.n114 150.4
R580 VDDA.n52 VDDA.n44 150.4
R581 VDDA.n46 VDDA.n41 150.4
R582 VDDA.n211 VDDA.n210 146.002
R583 VDDA.n99 VDDA.n98 146.002
R584 VDDA.n113 VDDA.n112 145.429
R585 VDDA.n132 VDDA.n131 145.429
R586 VDDA.n134 VDDA.n133 145.429
R587 VDDA.n136 VDDA.n135 145.429
R588 VDDA.n138 VDDA.n137 145.429
R589 VDDA.n39 VDDA.n38 145.429
R590 VDDA.n55 VDDA.n54 145.429
R591 VDDA.n57 VDDA.n56 145.429
R592 VDDA.n59 VDDA.n58 145.429
R593 VDDA.n61 VDDA.n60 145.429
R594 VDDA.n149 VDDA.n148 135.387
R595 VDDA.n140 VDDA.n139 135.387
R596 VDDA.n75 VDDA.n74 135.387
R597 VDDA.n63 VDDA.n62 135.387
R598 VDDA.t468 VDDA.t344 121.513
R599 VDDA.t438 VDDA.t468 121.513
R600 VDDA.t158 VDDA.t438 121.513
R601 VDDA.t462 VDDA.t158 121.513
R602 VDDA.t101 VDDA.t462 121.513
R603 VDDA.t74 VDDA.t217 121.513
R604 VDDA.t246 VDDA.t74 121.513
R605 VDDA.t84 VDDA.t246 121.513
R606 VDDA.t449 VDDA.t84 121.513
R607 VDDA.t371 VDDA.t449 121.513
R608 VDDA.t124 VDDA.t316 121.513
R609 VDDA.t49 VDDA.t124 121.513
R610 VDDA.t3 VDDA.t49 121.513
R611 VDDA.t6 VDDA.t3 121.513
R612 VDDA.t115 VDDA.t6 121.513
R613 VDDA.t106 VDDA.t114 121.513
R614 VDDA.t11 VDDA.t106 121.513
R615 VDDA.t235 VDDA.t11 121.513
R616 VDDA.t191 VDDA.t235 121.513
R617 VDDA.t350 VDDA.t191 121.513
R618 VDDA.n334 VDDA.n265 118.4
R619 VDDA.n330 VDDA.n270 118.4
R620 VDDA.n292 VDDA.n284 118.4
R621 VDDA.n286 VDDA.n281 118.4
R622 VDDA.n395 VDDA.n394 118.4
R623 VDDA.n390 VDDA.n385 118.4
R624 VDDA.n356 VDDA.n355 118.4
R625 VDDA.n351 VDDA.n346 118.4
R626 VDDA.n454 VDDA.n453 118.4
R627 VDDA.n460 VDDA.n459 118.4
R628 VDDA.n441 VDDA.n440 118.4
R629 VDDA.n446 VDDA.n445 118.4
R630 VDDA.n422 VDDA.n421 118.4
R631 VDDA.n427 VDDA.n426 118.4
R632 VDDA.n245 VDDA.n244 110.4
R633 VDDA.n249 VDDA.n248 110.4
R634 VDDA.n453 VDDA.n402 105.6
R635 VDDA.n460 VDDA.n402 105.6
R636 VDDA.n421 VDDA.n414 105.6
R637 VDDA.n427 VDDA.n414 105.6
R638 VDDA.t383 VDDA.t223 102.704
R639 VDDA.n183 VDDA.n153 102.4
R640 VDDA.n177 VDDA.n174 102.4
R641 VDDA.n21 VDDA.n20 102.4
R642 VDDA.n240 VDDA.n239 101.267
R643 VDDA.t21 VDDA.t353 98.2764
R644 VDDA.t41 VDDA.t21 98.2764
R645 VDDA.t23 VDDA.t41 98.2764
R646 VDDA.t242 VDDA.t23 98.2764
R647 VDDA.t77 VDDA.t242 98.2764
R648 VDDA.t44 VDDA.t225 98.2764
R649 VDDA.t208 VDDA.t44 98.2764
R650 VDDA.t0 VDDA.t208 98.2764
R651 VDDA.t19 VDDA.t0 98.2764
R652 VDDA.t380 VDDA.t19 98.2764
R653 VDDA.t188 VDDA.t359 98.2764
R654 VDDA.t227 VDDA.t188 98.2764
R655 VDDA.t72 VDDA.t227 98.2764
R656 VDDA.t111 VDDA.t72 98.2764
R657 VDDA.t200 VDDA.t111 98.2764
R658 VDDA.t447 VDDA.t79 98.2764
R659 VDDA.t229 VDDA.t447 98.2764
R660 VDDA.t37 VDDA.t229 98.2764
R661 VDDA.t204 VDDA.t37 98.2764
R662 VDDA.t404 VDDA.t204 98.2764
R663 VDDA.n103 VDDA.n101 97.4034
R664 VDDA.n2 VDDA.n0 97.4034
R665 VDDA.n111 VDDA.n110 96.8409
R666 VDDA.n109 VDDA.n108 96.8409
R667 VDDA.n107 VDDA.n106 96.8409
R668 VDDA.n105 VDDA.n104 96.8409
R669 VDDA.n103 VDDA.n102 96.8409
R670 VDDA.n10 VDDA.n9 96.8409
R671 VDDA.n8 VDDA.n7 96.8409
R672 VDDA.n6 VDDA.n5 96.8409
R673 VDDA.n4 VDDA.n3 96.8409
R674 VDDA.n2 VDDA.n1 96.8409
R675 VDDA.n28 VDDA.n27 96.0005
R676 VDDA.n29 VDDA.n15 96.0005
R677 VDDA.n36 VDDA.n35 96.0005
R678 VDDA.n180 VDDA.t163 93.3041
R679 VDDA.n180 VDDA.t90 93.3041
R680 VDDA.n32 VDDA.t75 93.3041
R681 VDDA.n32 VDDA.t212 93.3041
R682 VDDA.n219 VDDA.n218 92.5005
R683 VDDA.t68 VDDA.n219 92.5005
R684 VDDA.n220 VDDA.n217 92.5005
R685 VDDA.t68 VDDA.n220 92.5005
R686 VDDA.n224 VDDA.n223 92.5005
R687 VDDA.n233 VDDA.n224 92.5005
R688 VDDA.n225 VDDA.n222 92.5005
R689 VDDA.n234 VDDA.n225 92.5005
R690 VDDA.n208 VDDA.n207 92.5005
R691 VDDA.n204 VDDA.n203 92.5005
R692 VDDA.n206 VDDA.n204 92.5005
R693 VDDA.n205 VDDA.n197 92.5005
R694 VDDA.n209 VDDA.n198 92.5005
R695 VDDA.n206 VDDA.n198 92.5005
R696 VDDA.n175 VDDA.n153 92.5005
R697 VDDA.n179 VDDA.n178 92.5005
R698 VDDA.n180 VDDA.n179 92.5005
R699 VDDA.n177 VDDA.n176 92.5005
R700 VDDA.n182 VDDA.n181 92.5005
R701 VDDA.n181 VDDA.n180 92.5005
R702 VDDA.n125 VDDA.n124 92.5005
R703 VDDA.n121 VDDA.n120 92.5005
R704 VDDA.n123 VDDA.n121 92.5005
R705 VDDA.n122 VDDA.n114 92.5005
R706 VDDA.n126 VDDA.n115 92.5005
R707 VDDA.n123 VDDA.n115 92.5005
R708 VDDA.n130 VDDA.n127 92.5005
R709 VDDA.n144 VDDA.n130 92.5005
R710 VDDA.n129 VDDA.n128 92.5005
R711 VDDA.n144 VDDA.n129 92.5005
R712 VDDA.n96 VDDA.n95 92.5005
R713 VDDA.n92 VDDA.n91 92.5005
R714 VDDA.n94 VDDA.n92 92.5005
R715 VDDA.n93 VDDA.n85 92.5005
R716 VDDA.n97 VDDA.n86 92.5005
R717 VDDA.n94 VDDA.n86 92.5005
R718 VDDA.n52 VDDA.n51 92.5005
R719 VDDA.n48 VDDA.n47 92.5005
R720 VDDA.n50 VDDA.n48 92.5005
R721 VDDA.n49 VDDA.n41 92.5005
R722 VDDA.n53 VDDA.n42 92.5005
R723 VDDA.n50 VDDA.n42 92.5005
R724 VDDA.n72 VDDA.n71 92.5005
R725 VDDA.n71 VDDA.n70 92.5005
R726 VDDA.n69 VDDA.n68 92.5005
R727 VDDA.n70 VDDA.n69 92.5005
R728 VDDA.n23 VDDA.n16 92.5005
R729 VDDA.n24 VDDA.n23 92.5005
R730 VDDA.n22 VDDA.n21 92.5005
R731 VDDA.n26 VDDA.n25 92.5005
R732 VDDA.n25 VDDA.n24 92.5005
R733 VDDA.n28 VDDA.n17 92.5005
R734 VDDA.n31 VDDA.n11 92.5005
R735 VDDA.n32 VDDA.n31 92.5005
R736 VDDA.n30 VDDA.n29 92.5005
R737 VDDA.n34 VDDA.n33 92.5005
R738 VDDA.n33 VDDA.n32 92.5005
R739 VDDA.n36 VDDA.n12 92.5005
R740 VDDA.n317 VDDA.n267 92.5005
R741 VDDA.n332 VDDA.n267 92.5005
R742 VDDA.n334 VDDA.n333 92.5005
R743 VDDA.n269 VDDA.n266 92.5005
R744 VDDA.n332 VDDA.n266 92.5005
R745 VDDA.n331 VDDA.n330 92.5005
R746 VDDA.n292 VDDA.n291 92.5005
R747 VDDA.n288 VDDA.n287 92.5005
R748 VDDA.n290 VDDA.n288 92.5005
R749 VDDA.n289 VDDA.n281 92.5005
R750 VDDA.n293 VDDA.n282 92.5005
R751 VDDA.n290 VDDA.n282 92.5005
R752 VDDA.n394 VDDA.n393 92.5005
R753 VDDA.n389 VDDA.n388 92.5005
R754 VDDA.n392 VDDA.n389 92.5005
R755 VDDA.n391 VDDA.n390 92.5005
R756 VDDA.n396 VDDA.n386 92.5005
R757 VDDA.n392 VDDA.n386 92.5005
R758 VDDA.n376 VDDA.n375 92.5005
R759 VDDA.n343 VDDA.n342 92.5005
R760 VDDA.n377 VDDA.n343 92.5005
R761 VDDA.n379 VDDA.n378 92.5005
R762 VDDA.n344 VDDA.n341 92.5005
R763 VDDA.n377 VDDA.n344 92.5005
R764 VDDA.n355 VDDA.n354 92.5005
R765 VDDA.n350 VDDA.n349 92.5005
R766 VDDA.n353 VDDA.n350 92.5005
R767 VDDA.n352 VDDA.n351 92.5005
R768 VDDA.n357 VDDA.n347 92.5005
R769 VDDA.n353 VDDA.n347 92.5005
R770 VDDA.n455 VDDA.n454 92.5005
R771 VDDA.n404 VDDA.n403 92.5005
R772 VDDA.n456 VDDA.n404 92.5005
R773 VDDA.n459 VDDA.n458 92.5005
R774 VDDA.n405 VDDA.n402 92.5005
R775 VDDA.n457 VDDA.n405 92.5005
R776 VDDA.n442 VDDA.n441 92.5005
R777 VDDA.n410 VDDA.n409 92.5005
R778 VDDA.n443 VDDA.n410 92.5005
R779 VDDA.n445 VDDA.n444 92.5005
R780 VDDA.n411 VDDA.n408 92.5005
R781 VDDA.n443 VDDA.n411 92.5005
R782 VDDA.n423 VDDA.n422 92.5005
R783 VDDA.n416 VDDA.n415 92.5005
R784 VDDA.n424 VDDA.n416 92.5005
R785 VDDA.n426 VDDA.n425 92.5005
R786 VDDA.n417 VDDA.n414 92.5005
R787 VDDA.n424 VDDA.n417 92.5005
R788 VDDA.n24 VDDA.t8 91.6672
R789 VDDA.n24 VDDA.t102 91.6672
R790 VDDA.n228 VDDA.n227 87.4672
R791 VDDA.n332 VDDA.t61 86.3641
R792 VDDA.t192 VDDA.n332 86.3641
R793 VDDA.n290 VDDA.t156 86.3641
R794 VDDA.t443 VDDA.n290 86.3641
R795 VDDA.n227 VDDA.t363 85.438
R796 VDDA.n239 VDDA.t384 85.438
R797 VDDA.n233 VDDA.t362 81.3068
R798 VDDA.n239 VDDA.n238 81.0672
R799 VDDA.n229 VDDA.n227 81.0672
R800 VDDA.n377 VDDA.t290 79.907
R801 VDDA.t249 VDDA.n377 79.907
R802 VDDA.n392 VDDA.t65 79.1672
R803 VDDA.t432 VDDA.n392 79.1672
R804 VDDA.n353 VDDA.t214 79.1672
R805 VDDA.t103 VDDA.n353 79.1672
R806 VDDA.t196 VDDA.n457 79.1672
R807 VDDA.n151 VDDA.t132 78.8005
R808 VDDA.n151 VDDA.t168 78.8005
R809 VDDA.n154 VDDA.t95 78.8005
R810 VDDA.n154 VDDA.t166 78.8005
R811 VDDA.n156 VDDA.t145 78.8005
R812 VDDA.n156 VDDA.t138 78.8005
R813 VDDA.n158 VDDA.t160 78.8005
R814 VDDA.n158 VDDA.t151 78.8005
R815 VDDA.n160 VDDA.t13 78.8005
R816 VDDA.n160 VDDA.t164 78.8005
R817 VDDA.n162 VDDA.t91 78.8005
R818 VDDA.n162 VDDA.t93 78.8005
R819 VDDA.n164 VDDA.t15 78.8005
R820 VDDA.n164 VDDA.t134 78.8005
R821 VDDA.n166 VDDA.t136 78.8005
R822 VDDA.n166 VDDA.t147 78.8005
R823 VDDA.n168 VDDA.t149 78.8005
R824 VDDA.n168 VDDA.t71 78.8005
R825 VDDA.n170 VDDA.t162 78.8005
R826 VDDA.n170 VDDA.t89 78.8005
R827 VDDA.n443 VDDA.t152 77.9856
R828 VDDA.t140 VDDA.n443 77.9856
R829 VDDA.n424 VDDA.t182 77.9856
R830 VDDA.t27 VDDA.n424 77.9856
R831 VDDA.n237 VDDA.n222 64.0005
R832 VDDA.n329 VDDA.n271 64.0005
R833 VDDA.n321 VDDA.n271 64.0005
R834 VDDA.n321 VDDA.n320 64.0005
R835 VDDA.n320 VDDA.n317 64.0005
R836 VDDA.n317 VDDA.n316 64.0005
R837 VDDA.n316 VDDA.n308 64.0005
R838 VDDA.n308 VDDA.n263 64.0005
R839 VDDA.n335 VDDA.n263 64.0005
R840 VDDA.n357 VDDA.n356 64.0005
R841 VDDA.n357 VDDA.n346 64.0005
R842 VDDA.t176 VDDA.t332 62.9523
R843 VDDA.t454 VDDA.t176 62.9523
R844 VDDA.t463 VDDA.t454 62.9523
R845 VDDA.t418 VDDA.t463 62.9523
R846 VDDA.t119 VDDA.t418 62.9523
R847 VDDA.t221 VDDA.t194 62.9523
R848 VDDA.t452 VDDA.t221 62.9523
R849 VDDA.t465 VDDA.t452 62.9523
R850 VDDA.t219 VDDA.t465 62.9523
R851 VDDA.t365 VDDA.t219 62.9523
R852 VDDA.t52 VDDA.t310 62.9523
R853 VDDA.t50 VDDA.t52 62.9523
R854 VDDA.t4 VDDA.t50 62.9523
R855 VDDA.t16 VDDA.t4 62.9523
R856 VDDA.t104 VDDA.t16 62.9523
R857 VDDA.t9 VDDA.t232 62.9523
R858 VDDA.t232 VDDA.t121 62.9523
R859 VDDA.t121 VDDA.t125 62.9523
R860 VDDA.t125 VDDA.t116 62.9523
R861 VDDA.t116 VDDA.t338 62.9523
R862 VDDA.n396 VDDA.n395 62.7205
R863 VDDA.n396 VDDA.n385 62.7205
R864 VDDA.n215 VDDA.t69 62.5402
R865 VDDA.n215 VDDA.t329 62.5402
R866 VDDA.n246 VDDA.n245 61.6672
R867 VDDA.n248 VDDA.n247 61.6672
R868 VDDA.n146 VDDA.n145 61.6672
R869 VDDA.n143 VDDA.n142 61.6672
R870 VDDA.n65 VDDA.n40 61.6672
R871 VDDA.n67 VDDA.n66 61.6672
R872 VDDA.n123 VDDA.t101 60.7563
R873 VDDA.t217 VDDA.n123 60.7563
R874 VDDA.n50 VDDA.t115 60.7563
R875 VDDA.t114 VDDA.n50 60.7563
R876 VDDA.n256 VDDA.t471 59.5681
R877 VDDA.n255 VDDA.t469 59.5681
R878 VDDA.n244 VDDA.n217 57.6005
R879 VDDA.n249 VDDA.n217 57.6005
R880 VDDA.n456 VDDA.t96 57.5763
R881 VDDA.n255 VDDA.t472 51.8888
R882 VDDA.n230 VDDA.n222 51.2005
R883 VDDA.n206 VDDA.t77 49.1384
R884 VDDA.t225 VDDA.n206 49.1384
R885 VDDA.n94 VDDA.t200 49.1384
R886 VDDA.t79 VDDA.n94 49.1384
R887 VDDA.n257 VDDA.t470 48.9557
R888 VDDA.n252 VDDA.n251 48.3605
R889 VDDA.n242 VDDA.n241 43.8605
R890 VDDA.n172 VDDA.n171 42.0963
R891 VDDA.n186 VDDA.n185 41.5338
R892 VDDA.n260 VDDA.t239 39.4005
R893 VDDA.n260 VDDA.t211 39.4005
R894 VDDA.n261 VDDA.t58 39.4005
R895 VDDA.n261 VDDA.t86 39.4005
R896 VDDA.n311 VDDA.t203 39.4005
R897 VDDA.n311 VDDA.t173 39.4005
R898 VDDA.n309 VDDA.t108 39.4005
R899 VDDA.n309 VDDA.t100 39.4005
R900 VDDA.n306 VDDA.t62 39.4005
R901 VDDA.n306 VDDA.t193 39.4005
R902 VDDA.n318 VDDA.t40 39.4005
R903 VDDA.n318 VDDA.t60 39.4005
R904 VDDA.n305 VDDA.t241 39.4005
R905 VDDA.n305 VDDA.t128 39.4005
R906 VDDA.n324 VDDA.t175 39.4005
R907 VDDA.n324 VDDA.t237 39.4005
R908 VDDA.n272 VDDA.t179 39.4005
R909 VDDA.n272 VDDA.t64 39.4005
R910 VDDA.n302 VDDA.t110 39.4005
R911 VDDA.n302 VDDA.t207 39.4005
R912 VDDA.n300 VDDA.t143 39.4005
R913 VDDA.n300 VDDA.t446 39.4005
R914 VDDA.n298 VDDA.t423 39.4005
R915 VDDA.n298 VDDA.t199 39.4005
R916 VDDA.n296 VDDA.t187 39.4005
R917 VDDA.n296 VDDA.t421 39.4005
R918 VDDA.n280 VDDA.t157 39.4005
R919 VDDA.n280 VDDA.t444 39.4005
R920 VDDA.n278 VDDA.t461 39.4005
R921 VDDA.n278 VDDA.t130 39.4005
R922 VDDA.n276 VDDA.t185 39.4005
R923 VDDA.n276 VDDA.t26 39.4005
R924 VDDA.n274 VDDA.t427 39.4005
R925 VDDA.n274 VDDA.t435 39.4005
R926 VDDA.n273 VDDA.t459 39.4005
R927 VDDA.n273 VDDA.t36 39.4005
R928 VDDA.n383 VDDA.t66 39.4005
R929 VDDA.n383 VDDA.t433 39.4005
R930 VDDA.n400 VDDA.t197 39.4005
R931 VDDA.n400 VDDA.t440 39.4005
R932 VDDA.n449 VDDA.t431 39.4005
R933 VDDA.n449 VDDA.t97 39.4005
R934 VDDA.n406 VDDA.t429 39.4005
R935 VDDA.n406 VDDA.t155 39.4005
R936 VDDA.n430 VDDA.t141 39.4005
R937 VDDA.n430 VDDA.t442 39.4005
R938 VDDA.n432 VDDA.t48 39.4005
R939 VDDA.n432 VDDA.t153 39.4005
R940 VDDA.n434 VDDA.t181 39.4005
R941 VDDA.n434 VDDA.t32 39.4005
R942 VDDA.n436 VDDA.t34 39.4005
R943 VDDA.n436 VDDA.t451 39.4005
R944 VDDA.n412 VDDA.t28 39.4005
R945 VDDA.n412 VDDA.t30 39.4005
R946 VDDA.n418 VDDA.t425 39.4005
R947 VDDA.n418 VDDA.t183 39.4005
R948 VDDA.n144 VDDA.t119 31.4764
R949 VDDA.t194 VDDA.n144 31.4764
R950 VDDA.n70 VDDA.t104 31.4764
R951 VDDA.n70 VDDA.t9 31.4764
R952 VDDA.n29 VDDA.n28 28.663
R953 VDDA.n251 VDDA.n250 25.6005
R954 VDDA.n243 VDDA.n242 25.6005
R955 VDDA.n185 VDDA.n184 25.6005
R956 VDDA.n173 VDDA.n172 25.6005
R957 VDDA.n258 VDDA.n254 24.7453
R958 VDDA.n250 VDDA.n249 24.5338
R959 VDDA.n244 VDDA.n243 24.5338
R960 VDDA.n238 VDDA.n237 24.5338
R961 VDDA.n230 VDDA.n229 24.5338
R962 VDDA.n457 VDDA.n456 21.5914
R963 VDDA.n254 VDDA.n253 21.5392
R964 VDDA.n202 VDDA.n201 21.3338
R965 VDDA.n200 VDDA.n199 21.3338
R966 VDDA.n184 VDDA.n183 21.3338
R967 VDDA.n174 VDDA.n173 21.3338
R968 VDDA.n119 VDDA.n118 21.3338
R969 VDDA.n117 VDDA.n116 21.3338
R970 VDDA.n148 VDDA.n147 21.3338
R971 VDDA.n141 VDDA.n140 21.3338
R972 VDDA.n90 VDDA.n89 21.3338
R973 VDDA.n88 VDDA.n87 21.3338
R974 VDDA.n46 VDDA.n45 21.3338
R975 VDDA.n44 VDDA.n43 21.3338
R976 VDDA.n74 VDDA.n73 21.3338
R977 VDDA.n64 VDDA.n63 21.3338
R978 VDDA.n20 VDDA.n19 21.3338
R979 VDDA.n27 VDDA.n18 21.3338
R980 VDDA.n15 VDDA.n14 21.3338
R981 VDDA.n35 VDDA.n13 21.3338
R982 VDDA.n265 VDDA.n264 21.3338
R983 VDDA.n270 VDDA.n268 21.3338
R984 VDDA.n284 VDDA.n283 21.3338
R985 VDDA.n286 VDDA.n285 21.3338
R986 VDDA.n395 VDDA.n387 21.3338
R987 VDDA.n385 VDDA.n384 21.3338
R988 VDDA.n356 VDDA.n348 21.3338
R989 VDDA.n346 VDDA.n345 21.3338
R990 VDDA.n37 VDDA.n36 19.5505
R991 VDDA.n127 VDDA.n126 19.538
R992 VDDA.n72 VDDA.n53 19.538
R993 VDDA.n211 VDDA.n209 19.2005
R994 VDDA.n99 VDDA.n97 19.2005
R995 VDDA.n381 VDDA.n380 19.2005
R996 VDDA.n374 VDDA.n373 19.2005
R997 VDDA.n461 VDDA.n460 19.2005
R998 VDDA.n453 VDDA.n452 19.2005
R999 VDDA.n447 VDDA.n446 19.2005
R1000 VDDA.n440 VDDA.n439 19.2005
R1001 VDDA.n428 VDDA.n427 19.2005
R1002 VDDA.n421 VDDA.n420 19.2005
R1003 VDDA.n232 VDDA.n231 18.5005
R1004 VDDA.n236 VDDA.n235 18.5005
R1005 VDDA.t223 VDDA.n234 17.1176
R1006 VDDA.n188 VDDA.n111 16.8443
R1007 VDDA.n372 VDDA.n357 16.363
R1008 VDDA.n468 VDDA.t258 15.0181
R1009 VDDA.n420 VDDA.n419 14.363
R1010 VDDA.n228 VDDA.n221 14.0505
R1011 VDDA.n373 VDDA.n372 13.8005
R1012 VDDA.n382 VDDA.n381 13.8005
R1013 VDDA.n452 VDDA.n451 13.8005
R1014 VDDA.n439 VDDA.n438 13.8005
R1015 VDDA.n429 VDDA.n428 13.8005
R1016 VDDA.n448 VDDA.n447 13.8005
R1017 VDDA.n462 VDDA.n461 13.8005
R1018 VDDA.n37 VDDA.n10 13.6255
R1019 VDDA.n213 VDDA.n189 13.563
R1020 VDDA.n339 VDDA.t275 13.1338
R1021 VDDA.n339 VDDA.t273 13.1338
R1022 VDDA.n358 VDDA.t294 13.1338
R1023 VDDA.n358 VDDA.t255 13.1338
R1024 VDDA.n360 VDDA.t266 13.1338
R1025 VDDA.n360 VDDA.t285 13.1338
R1026 VDDA.n362 VDDA.t250 13.1338
R1027 VDDA.n362 VDDA.t269 13.1338
R1028 VDDA.n364 VDDA.t283 13.1338
R1029 VDDA.n364 VDDA.t291 13.1338
R1030 VDDA.n366 VDDA.t264 13.1338
R1031 VDDA.n366 VDDA.t260 13.1338
R1032 VDDA.n368 VDDA.t289 13.1338
R1033 VDDA.n368 VDDA.t299 13.1338
R1034 VDDA.n370 VDDA.t257 13.1338
R1035 VDDA.n370 VDDA.t278 13.1338
R1036 VDDA.t363 VDDA.n226 12.313
R1037 VDDA.n226 VDDA.t224 12.313
R1038 VDDA.n210 VDDA.t78 11.2576
R1039 VDDA.n210 VDDA.t226 11.2576
R1040 VDDA.n194 VDDA.t45 11.2576
R1041 VDDA.n194 VDDA.t209 11.2576
R1042 VDDA.n193 VDDA.t1 11.2576
R1043 VDDA.n193 VDDA.t20 11.2576
R1044 VDDA.n191 VDDA.t24 11.2576
R1045 VDDA.n191 VDDA.t243 11.2576
R1046 VDDA.n190 VDDA.t22 11.2576
R1047 VDDA.n190 VDDA.t42 11.2576
R1048 VDDA.n98 VDDA.t201 11.2576
R1049 VDDA.n98 VDDA.t80 11.2576
R1050 VDDA.n82 VDDA.t448 11.2576
R1051 VDDA.n82 VDDA.t230 11.2576
R1052 VDDA.n81 VDDA.t38 11.2576
R1053 VDDA.n81 VDDA.t205 11.2576
R1054 VDDA.n79 VDDA.t73 11.2576
R1055 VDDA.n79 VDDA.t112 11.2576
R1056 VDDA.n78 VDDA.t189 11.2576
R1057 VDDA.n78 VDDA.t228 11.2576
R1058 VDDA.n189 VDDA.n188 9.5005
R1059 VDDA.n212 VDDA.n211 9.3005
R1060 VDDA.n100 VDDA.n99 9.3005
R1061 VDDA.n325 VDDA.n271 9.3005
R1062 VDDA.n322 VDDA.n321 9.3005
R1063 VDDA.n320 VDDA.n319 9.3005
R1064 VDDA.n317 VDDA.n307 9.3005
R1065 VDDA.n316 VDDA.n315 9.3005
R1066 VDDA.n312 VDDA.n308 9.3005
R1067 VDDA.n263 VDDA.n262 9.3005
R1068 VDDA.n336 VDDA.n335 9.3005
R1069 VDDA.n329 VDDA.n328 9.3005
R1070 VDDA.n294 VDDA.n293 9.3005
R1071 VDDA.n397 VDDA.n396 9.3005
R1072 VDDA.n241 VDDA.n240 8.938
R1073 VDDA.n258 VDDA.n257 8.03219
R1074 VDDA.n110 VDDA.t170 8.0005
R1075 VDDA.n110 VDDA.t171 8.0005
R1076 VDDA.n108 VDDA.t98 8.0005
R1077 VDDA.n108 VDDA.t417 8.0005
R1078 VDDA.n106 VDDA.t169 8.0005
R1079 VDDA.n106 VDDA.t456 8.0005
R1080 VDDA.n104 VDDA.t213 8.0005
R1081 VDDA.n104 VDDA.t437 8.0005
R1082 VDDA.n102 VDDA.t467 8.0005
R1083 VDDA.n102 VDDA.t76 8.0005
R1084 VDDA.n101 VDDA.t218 8.0005
R1085 VDDA.n101 VDDA.t67 8.0005
R1086 VDDA.n9 VDDA.t247 8.0005
R1087 VDDA.n9 VDDA.t245 8.0005
R1088 VDDA.n7 VDDA.t18 8.0005
R1089 VDDA.n7 VDDA.t113 8.0005
R1090 VDDA.n5 VDDA.t190 8.0005
R1091 VDDA.n5 VDDA.t234 8.0005
R1092 VDDA.n3 VDDA.t123 8.0005
R1093 VDDA.n3 VDDA.t54 8.0005
R1094 VDDA.n1 VDDA.t2 8.0005
R1095 VDDA.n1 VDDA.t244 8.0005
R1096 VDDA.n0 VDDA.t231 8.0005
R1097 VDDA.n0 VDDA.t43 8.0005
R1098 VDDA.n213 VDDA.n212 7.8755
R1099 VDDA.n189 VDDA.n100 7.8755
R1100 VDDA.n463 VDDA.n462 7.44175
R1101 VDDA.n253 VDDA.n252 6.6255
R1102 VDDA.n112 VDDA.t466 6.56717
R1103 VDDA.n112 VDDA.t220 6.56717
R1104 VDDA.n131 VDDA.t222 6.56717
R1105 VDDA.n131 VDDA.t453 6.56717
R1106 VDDA.n133 VDDA.t120 6.56717
R1107 VDDA.n133 VDDA.t195 6.56717
R1108 VDDA.n135 VDDA.t464 6.56717
R1109 VDDA.n135 VDDA.t419 6.56717
R1110 VDDA.n137 VDDA.t177 6.56717
R1111 VDDA.n137 VDDA.t455 6.56717
R1112 VDDA.n38 VDDA.t53 6.56717
R1113 VDDA.n38 VDDA.t51 6.56717
R1114 VDDA.n54 VDDA.t5 6.56717
R1115 VDDA.n54 VDDA.t17 6.56717
R1116 VDDA.n56 VDDA.t105 6.56717
R1117 VDDA.n56 VDDA.t10 6.56717
R1118 VDDA.n58 VDDA.t233 6.56717
R1119 VDDA.n58 VDDA.t122 6.56717
R1120 VDDA.n60 VDDA.t126 6.56717
R1121 VDDA.n60 VDDA.t117 6.56717
R1122 VDDA.n399 VDDA.n398 6.13371
R1123 VDDA.n338 VDDA.n337 6.098
R1124 VDDA.n77 VDDA.n76 5.438
R1125 VDDA.n241 VDDA.n216 5.1255
R1126 VDDA.n214 VDDA.n77 5.0005
R1127 VDDA.n212 VDDA.n196 4.5005
R1128 VDDA.n188 VDDA.n187 4.5005
R1129 VDDA.n100 VDDA.n84 4.5005
R1130 VDDA.n214 VDDA.n213 4.5005
R1131 VDDA.n295 VDDA.n294 4.5005
R1132 VDDA.n328 VDDA.n327 4.5005
R1133 VDDA.n326 VDDA.n325 4.5005
R1134 VDDA.n323 VDDA.n322 4.5005
R1135 VDDA.n319 VDDA.n304 4.5005
R1136 VDDA.n310 VDDA.n307 4.5005
R1137 VDDA.n315 VDDA.n314 4.5005
R1138 VDDA.n313 VDDA.n312 4.5005
R1139 VDDA.n262 VDDA.n259 4.5005
R1140 VDDA.n337 VDDA.n336 4.5005
R1141 VDDA.n398 VDDA.n397 4.5005
R1142 VDDA.n234 VDDA.n233 4.27978
R1143 VDDA.n256 VDDA.n255 4.12334
R1144 VDDA.n469 VDDA 4.08025
R1145 VDDA.n327 VDDA.n303 3.3755
R1146 VDDA.n77 VDDA.n37 3.09425
R1147 VDDA.n187 VDDA.n186 2.938
R1148 VDDA.n257 VDDA.n256 2.93377
R1149 VDDA.n451 VDDA.n448 2.5005
R1150 VDDA.n398 VDDA.n382 2.47371
R1151 VDDA.n253 VDDA.n214 1.938
R1152 VDDA.n438 VDDA.n429 1.813
R1153 VDDA VDDA.n469 1.20605
R1154 VDDA VDDA.n468 1.0815
R1155 VDDA.n372 VDDA.n371 1.0005
R1156 VDDA.n371 VDDA.n369 1.0005
R1157 VDDA.n369 VDDA.n367 1.0005
R1158 VDDA.n367 VDDA.n365 1.0005
R1159 VDDA.n365 VDDA.n363 1.0005
R1160 VDDA.n363 VDDA.n361 1.0005
R1161 VDDA.n361 VDDA.n359 1.0005
R1162 VDDA.n359 VDDA.n340 1.0005
R1163 VDDA.n382 VDDA.n340 1.0005
R1164 VDDA.n187 VDDA.n150 0.938
R1165 VDDA.n338 VDDA.n258 0.840625
R1166 VDDA.n469 VDDA.n254 0.7948
R1167 VDDA.n399 VDDA.n338 0.74075
R1168 VDDA.n240 VDDA.n221 0.6255
R1169 VDDA.n196 VDDA.n195 0.6255
R1170 VDDA.n196 VDDA.n192 0.6255
R1171 VDDA.n84 VDDA.n83 0.6255
R1172 VDDA.n84 VDDA.n80 0.6255
R1173 VDDA.n277 VDDA.n275 0.6255
R1174 VDDA.n279 VDDA.n277 0.6255
R1175 VDDA.n295 VDDA.n279 0.6255
R1176 VDDA.n297 VDDA.n295 0.6255
R1177 VDDA.n299 VDDA.n297 0.6255
R1178 VDDA.n301 VDDA.n299 0.6255
R1179 VDDA.n303 VDDA.n301 0.6255
R1180 VDDA.n327 VDDA.n326 0.6255
R1181 VDDA.n326 VDDA.n323 0.6255
R1182 VDDA.n323 VDDA.n304 0.6255
R1183 VDDA.n310 VDDA.n304 0.6255
R1184 VDDA.n314 VDDA.n310 0.6255
R1185 VDDA.n314 VDDA.n313 0.6255
R1186 VDDA.n313 VDDA.n259 0.6255
R1187 VDDA.n337 VDDA.n259 0.6255
R1188 VDDA.n171 VDDA.n169 0.563
R1189 VDDA.n169 VDDA.n167 0.563
R1190 VDDA.n167 VDDA.n165 0.563
R1191 VDDA.n165 VDDA.n163 0.563
R1192 VDDA.n163 VDDA.n161 0.563
R1193 VDDA.n161 VDDA.n159 0.563
R1194 VDDA.n159 VDDA.n157 0.563
R1195 VDDA.n157 VDDA.n155 0.563
R1196 VDDA.n155 VDDA.n152 0.563
R1197 VDDA.n186 VDDA.n152 0.563
R1198 VDDA.n138 VDDA.n136 0.563
R1199 VDDA.n136 VDDA.n134 0.563
R1200 VDDA.n134 VDDA.n132 0.563
R1201 VDDA.n132 VDDA.n113 0.563
R1202 VDDA.n150 VDDA.n113 0.563
R1203 VDDA.n105 VDDA.n103 0.563
R1204 VDDA.n107 VDDA.n105 0.563
R1205 VDDA.n109 VDDA.n107 0.563
R1206 VDDA.n111 VDDA.n109 0.563
R1207 VDDA.n61 VDDA.n59 0.563
R1208 VDDA.n59 VDDA.n57 0.563
R1209 VDDA.n57 VDDA.n55 0.563
R1210 VDDA.n55 VDDA.n39 0.563
R1211 VDDA.n76 VDDA.n39 0.563
R1212 VDDA.n4 VDDA.n2 0.563
R1213 VDDA.n6 VDDA.n4 0.563
R1214 VDDA.n8 VDDA.n6 0.563
R1215 VDDA.n10 VDDA.n8 0.563
R1216 VDDA.n419 VDDA.n413 0.563
R1217 VDDA.n429 VDDA.n413 0.563
R1218 VDDA.n438 VDDA.n437 0.563
R1219 VDDA.n437 VDDA.n435 0.563
R1220 VDDA.n435 VDDA.n433 0.563
R1221 VDDA.n433 VDDA.n431 0.563
R1222 VDDA.n431 VDDA.n407 0.563
R1223 VDDA.n448 VDDA.n407 0.563
R1224 VDDA.n451 VDDA.n450 0.563
R1225 VDDA.n450 VDDA.n401 0.563
R1226 VDDA.n462 VDDA.n401 0.563
R1227 VDDA.n463 VDDA.n399 0.546875
R1228 VDDA.n468 VDDA.n463 0.370625
R1229 VDDA.n252 VDDA.n216 0.2505
R1230 VDDA.t251 VDDA.t267 0.1603
R1231 VDDA.t295 VDDA.t287 0.1603
R1232 VDDA.t292 VDDA.t252 0.1603
R1233 VDDA.t280 VDDA.t276 0.1603
R1234 VDDA.t253 VDDA.t270 0.1603
R1235 VDDA.t297 VDDA.t281 0.1603
R1236 VDDA.t271 VDDA.t286 0.1603
R1237 VDDA.t262 VDDA.t248 0.1603
R1238 VDDA.n465 VDDA.t279 0.159278
R1239 VDDA.n466 VDDA.t261 0.159278
R1240 VDDA.n467 VDDA.t296 0.159278
R1241 VDDA.n467 VDDA.t251 0.1368
R1242 VDDA.n467 VDDA.t295 0.1368
R1243 VDDA.n466 VDDA.t292 0.1368
R1244 VDDA.n466 VDDA.t280 0.1368
R1245 VDDA.n465 VDDA.t253 0.1368
R1246 VDDA.n465 VDDA.t297 0.1368
R1247 VDDA.n464 VDDA.t271 0.1368
R1248 VDDA.n464 VDDA.t262 0.1368
R1249 VDDA.t279 VDDA.n464 0.00152174
R1250 VDDA.t261 VDDA.n465 0.00152174
R1251 VDDA.t296 VDDA.n466 0.00152174
R1252 VDDA.t258 VDDA.n467 0.00152174
R1253 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 628.034
R1254 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 626.784
R1255 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 622.284
R1256 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 289.2
R1257 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 289.2
R1258 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 227.252
R1259 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 212.733
R1260 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 212.733
R1261 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 176.733
R1262 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 176.733
R1263 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R1264 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 176.733
R1265 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 176.733
R1266 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 152
R1267 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 152
R1268 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 112.468
R1269 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 112.468
R1270 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R1271 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R1272 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 112.468
R1273 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R1274 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R1275 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 112.468
R1276 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 78.8005
R1277 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 78.8005
R1278 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R1279 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R1280 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R1281 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 78.8005
R1282 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 48.0005
R1283 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R1284 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 48.0005
R1285 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 48.0005
R1286 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 48.0005
R1287 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R1288 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R1289 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 45.5227
R1290 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 45.5227
R1291 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 45.5227
R1292 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 15.488
R1293 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 14.238
R1294 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 6.1255
R1295 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 5.7505
R1296 GNDA.n209 GNDA.n29 227083
R1297 GNDA.n1394 GNDA.n213 33145.9
R1298 GNDA.n207 GNDA.n30 31003.1
R1299 GNDA.n2373 GNDA.n79 29344.6
R1300 GNDA.n210 GNDA.n207 28430.8
R1301 GNDA.n2373 GNDA.n92 28430.8
R1302 GNDA.n209 GNDA.n208 26656.2
R1303 GNDA.n1397 GNDA.n1396 26648.4
R1304 GNDA.n1397 GNDA.n214 26648.4
R1305 GNDA.n108 GNDA.n92 23523.1
R1306 GNDA.n210 GNDA.n108 23523.1
R1307 GNDA.n1394 GNDA.n212 21442.2
R1308 GNDA.n2336 GNDA.n108 19630.8
R1309 GNDA.n2337 GNDA.n107 19321
R1310 GNDA.n2338 GNDA.n92 17609.2
R1311 GNDA.n211 GNDA.n210 17609.2
R1312 GNDA.n2332 GNDA.n214 17265.8
R1313 GNDA.n214 GNDA.n213 15861.4
R1314 GNDA.n1395 GNDA.n1394 13428.1
R1315 GNDA.n1400 GNDA.n1399 12361.8
R1316 GNDA.n1401 GNDA.n1399 12312.5
R1317 GNDA.n2338 GNDA.n2337 12272.1
R1318 GNDA.n210 GNDA.n209 11934.7
R1319 GNDA.n1405 GNDA.n1400 11918.5
R1320 GNDA.n1405 GNDA.n1401 11869.2
R1321 GNDA.n1396 GNDA.n1395 11169.2
R1322 GNDA.n2336 GNDA.n2335 10879.5
R1323 GNDA.n2404 GNDA.n62 10835
R1324 GNDA.n2404 GNDA.n63 10835
R1325 GNDA.n62 GNDA.n61 10835
R1326 GNDA.n63 GNDA.n61 10835
R1327 GNDA.n1479 GNDA.n1397 10371.4
R1328 GNDA.n2339 GNDA.n2338 10311.6
R1329 GNDA.n2389 GNDA.n59 9308.25
R1330 GNDA.n2400 GNDA.n59 9308.25
R1331 GNDA.n2389 GNDA.n60 9308.25
R1332 GNDA.n2400 GNDA.n60 9308.25
R1333 GNDA.n2418 GNDA.n31 9259
R1334 GNDA.n2323 GNDA.n220 9062
R1335 GNDA.n2418 GNDA.n32 8914.25
R1336 GNDA.n249 GNDA.n246 8175.5
R1337 GNDA.n252 GNDA.n246 8126.25
R1338 GNDA.n1396 GNDA.n259 7953.85
R1339 GNDA.n2326 GNDA.n216 7880
R1340 GNDA.n2330 GNDA.n216 7880
R1341 GNDA.n1485 GNDA.n1390 7880
R1342 GNDA.n1481 GNDA.n1390 7880
R1343 GNDA.n2326 GNDA.n217 7830.75
R1344 GNDA.n2330 GNDA.n217 7830.75
R1345 GNDA.n1485 GNDA.n1391 7830.75
R1346 GNDA.n1481 GNDA.n1391 7830.75
R1347 GNDA.n146 GNDA.n134 7732.25
R1348 GNDA.n182 GNDA.n134 7732.25
R1349 GNDA.n146 GNDA.n135 7732.25
R1350 GNDA.n182 GNDA.n135 7732.25
R1351 GNDA.n87 GNDA.n81 7732.25
R1352 GNDA.n2384 GNDA.n81 7732.25
R1353 GNDA.n87 GNDA.n82 7732.25
R1354 GNDA.n2384 GNDA.n82 7732.25
R1355 GNDA.n249 GNDA.n245 7732.25
R1356 GNDA.n252 GNDA.n245 7683
R1357 GNDA.n2300 GNDA.n2297 6845.75
R1358 GNDA.n2304 GNDA.n2297 6845.75
R1359 GNDA.n2300 GNDA.n239 6796.5
R1360 GNDA.n2304 GNDA.n239 6796.5
R1361 GNDA.n236 GNDA.n234 6698
R1362 GNDA.n2307 GNDA.n236 6698
R1363 GNDA.n234 GNDA.n231 6648.75
R1364 GNDA.n2307 GNDA.n231 6648.75
R1365 GNDA.n2337 GNDA.n2336 6600
R1366 GNDA.n133 GNDA.n128 6057.75
R1367 GNDA.n185 GNDA.n128 6057.75
R1368 GNDA.n184 GNDA.n133 6057.75
R1369 GNDA.n185 GNDA.n184 6057.75
R1370 GNDA.n2371 GNDA.n94 6057.75
R1371 GNDA.n2365 GNDA.n94 6057.75
R1372 GNDA.n2371 GNDA.n96 6057.75
R1373 GNDA.n2365 GNDA.n96 6057.75
R1374 GNDA.n2411 GNDA.n31 5713
R1375 GNDA.n2413 GNDA.n32 5713
R1376 GNDA.n208 GNDA.n79 5446.53
R1377 GNDA.n189 GNDA.n124 5368.25
R1378 GNDA.n2357 GNDA.n102 5368.25
R1379 GNDA.n194 GNDA.n124 5319
R1380 GNDA.n193 GNDA.n189 5319
R1381 GNDA.n2359 GNDA.n102 5319
R1382 GNDA.n194 GNDA.n193 5269.75
R1383 GNDA.n2359 GNDA.n101 5269.75
R1384 GNDA.n206 GNDA.n111 5171.25
R1385 GNDA.n2374 GNDA.n90 5171.25
R1386 GNDA.n202 GNDA.n111 5122
R1387 GNDA.n2357 GNDA.n101 5122
R1388 GNDA.n2349 GNDA.n90 5122
R1389 GNDA.n2323 GNDA.n221 4974.25
R1390 GNDA.n1422 GNDA.n1418 4974.25
R1391 GNDA.n1426 GNDA.n1418 4974.25
R1392 GNDA.n206 GNDA.n112 4944.7
R1393 GNDA.n2374 GNDA.n91 4944.7
R1394 GNDA.n39 GNDA.n38 4925
R1395 GNDA.n40 GNDA.n38 4925
R1396 GNDA.n202 GNDA.n112 4895.45
R1397 GNDA.n2349 GNDA.n91 4895.45
R1398 GNDA.n58 GNDA.n39 4728
R1399 GNDA.n58 GNDA.n40 4728
R1400 GNDA.n2292 GNDA.n243 4678.75
R1401 GNDA.n2288 GNDA.n243 4629.5
R1402 GNDA.n2292 GNDA.n242 4629.5
R1403 GNDA.n2274 GNDA.n257 4580.25
R1404 GNDA.n2285 GNDA.n257 4580.25
R1405 GNDA.n2288 GNDA.n242 4580.25
R1406 GNDA.n2282 GNDA.n2281 4580.25
R1407 GNDA.n2281 GNDA.n2280 4580.25
R1408 GNDA.n1478 GNDA.n1406 4531
R1409 GNDA.n1478 GNDA.n1407 4531
R1410 GNDA.n1406 GNDA.n1398 4531
R1411 GNDA.n1407 GNDA.n1398 4531
R1412 GNDA.n1430 GNDA.n1422 4531
R1413 GNDA.n1430 GNDA.n1426 4531
R1414 GNDA.n2274 GNDA.n256 4481.75
R1415 GNDA.n2285 GNDA.n256 4481.75
R1416 GNDA.n2280 GNDA.n2279 4481.75
R1417 GNDA.n2282 GNDA.n2279 4481.75
R1418 GNDA.n2340 GNDA.n2339 4181.99
R1419 GNDA.n208 GNDA.n92 3964.58
R1420 GNDA.n2411 GNDA.n36 3595.25
R1421 GNDA.n2421 GNDA.n26 3349
R1422 GNDA.n2407 GNDA.n26 3299.75
R1423 GNDA.n2332 GNDA.n2331 3287.9
R1424 GNDA.n2413 GNDA.n36 3250.5
R1425 GNDA.n2421 GNDA.n27 3250.5
R1426 GNDA.n2407 GNDA.n27 3201.25
R1427 GNDA.n2333 GNDA.n213 3156.82
R1428 GNDA.n1395 GNDA.n1393 2871.88
R1429 GNDA.n119 GNDA.n116 2326.02
R1430 GNDA.n190 GNDA.n116 2326.02
R1431 GNDA.n2343 GNDA.n2342 2326.02
R1432 GNDA.n2345 GNDA.n2343 2326.02
R1433 GNDA.n1467 GNDA.n1441 2142.38
R1434 GNDA.n1419 GNDA.n1417 2142.38
R1435 GNDA.n1473 GNDA.n1441 1846.88
R1436 GNDA.n1417 GNDA.n1413 1846.88
R1437 GNDA.n2334 GNDA.n2333 1749.05
R1438 GNDA.n2388 GNDA.n79 1658.46
R1439 GNDA.t224 GNDA.n315 1378.22
R1440 GNDA.n2333 GNDA.n2332 1226.55
R1441 GNDA.n852 GNDA.n713 1214.72
R1442 GNDA.n846 GNDA.n713 1214.72
R1443 GNDA.n846 GNDA.n845 1214.72
R1444 GNDA.n845 GNDA.n844 1214.72
R1445 GNDA.n844 GNDA.n313 1214.72
R1446 GNDA.n837 GNDA.n312 1214.72
R1447 GNDA.n837 GNDA.n836 1214.72
R1448 GNDA.n836 GNDA.n835 1214.72
R1449 GNDA.n835 GNDA.n292 1214.72
R1450 GNDA.n2244 GNDA.n292 1214.72
R1451 GNDA.n1896 GNDA.n853 1214.72
R1452 GNDA.n1890 GNDA.n853 1214.72
R1453 GNDA.n1890 GNDA.n1889 1214.72
R1454 GNDA.n1889 GNDA.n1888 1214.72
R1455 GNDA.n1888 GNDA.n311 1214.72
R1456 GNDA.n1881 GNDA.n310 1214.72
R1457 GNDA.n1881 GNDA.n1880 1214.72
R1458 GNDA.n1880 GNDA.n1879 1214.72
R1459 GNDA.n1879 GNDA.n995 1214.72
R1460 GNDA.n995 GNDA.n309 1214.72
R1461 GNDA.n2335 GNDA.n2334 1163.28
R1462 GNDA.n199 GNDA.n116 1114.8
R1463 GNDA.n2352 GNDA.n2343 1114.8
R1464 GNDA.n2240 GNDA.n341 1097.06
R1465 GNDA.n1469 GNDA.n1441 991.841
R1466 GNDA.n1433 GNDA.n1417 991.841
R1467 GNDA.n211 GNDA.n109 971.551
R1468 GNDA.n2335 GNDA.n211 890.324
R1469 GNDA.n2388 GNDA.t287 863.077
R1470 GNDA.t308 GNDA.n30 863.077
R1471 GNDA.n2334 GNDA.n212 831.111
R1472 GNDA.t224 GNDA.n313 823.313
R1473 GNDA.t224 GNDA.n311 823.313
R1474 GNDA.n1402 GNDA.n224 803.201
R1475 GNDA.n1403 GNDA.n224 800
R1476 GNDA.n1404 GNDA.n1402 774.4
R1477 GNDA.n1404 GNDA.n1403 771.201
R1478 GNDA.n1847 GNDA.n308 735.866
R1479 GNDA.n125 GNDA.t235 734.418
R1480 GNDA.n129 GNDA.t220 734.418
R1481 GNDA.n2362 GNDA.t241 734.418
R1482 GNDA.n97 GNDA.t231 734.418
R1483 GNDA.t80 GNDA.n250 712.497
R1484 GNDA.n74 GNDA.n73 704
R1485 GNDA.n75 GNDA.n74 697.601
R1486 GNDA.n251 GNDA.n238 685.793
R1487 GNDA.n34 GNDA.t251 682.201
R1488 GNDA.n1599 GNDA.n1571 675.63
R1489 GNDA.n149 GNDA.t265 666.134
R1490 GNDA.t224 GNDA.n298 662.155
R1491 GNDA.n121 GNDA.n120 617.601
R1492 GNDA.n104 GNDA.n103 617.601
R1493 GNDA.n2417 GNDA.n33 601.601
R1494 GNDA.n2402 GNDA.n2390 598.4
R1495 GNDA.n2402 GNDA.n2401 598.4
R1496 GNDA.n1354 GNDA.n1353 585
R1497 GNDA.n1355 GNDA.n1198 585
R1498 GNDA.n1357 GNDA.n1356 585
R1499 GNDA.n1359 GNDA.n1197 585
R1500 GNDA.n1362 GNDA.n1361 585
R1501 GNDA.n1363 GNDA.n1196 585
R1502 GNDA.n1365 GNDA.n1364 585
R1503 GNDA.n1367 GNDA.n1195 585
R1504 GNDA.n1370 GNDA.n1369 585
R1505 GNDA.n1371 GNDA.n1194 585
R1506 GNDA.n1373 GNDA.n1372 585
R1507 GNDA.n1375 GNDA.n680 585
R1508 GNDA.n1335 GNDA.n1334 585
R1509 GNDA.n1337 GNDA.n1204 585
R1510 GNDA.n1339 GNDA.n1338 585
R1511 GNDA.n1340 GNDA.n1203 585
R1512 GNDA.n1342 GNDA.n1341 585
R1513 GNDA.n1344 GNDA.n1201 585
R1514 GNDA.n1346 GNDA.n1345 585
R1515 GNDA.n1347 GNDA.n1200 585
R1516 GNDA.n1349 GNDA.n1348 585
R1517 GNDA.n1351 GNDA.n1199 585
R1518 GNDA.n1544 GNDA.n1519 585
R1519 GNDA.n1543 GNDA.n1542 585
R1520 GNDA.n1541 GNDA.n1520 585
R1521 GNDA.n1539 GNDA.n1538 585
R1522 GNDA.n1537 GNDA.n1522 585
R1523 GNDA.n1536 GNDA.n1535 585
R1524 GNDA.n1534 GNDA.n1523 585
R1525 GNDA.n1532 GNDA.n1531 585
R1526 GNDA.n1530 GNDA.n1525 585
R1527 GNDA.n1529 GNDA.n1528 585
R1528 GNDA.n1527 GNDA.n1036 585
R1529 GNDA.n1693 GNDA.n1692 585
R1530 GNDA.n1546 GNDA.n1545 585
R1531 GNDA.n1548 GNDA.n1518 585
R1532 GNDA.n1551 GNDA.n1550 585
R1533 GNDA.n1552 GNDA.n1517 585
R1534 GNDA.n1554 GNDA.n1553 585
R1535 GNDA.n1556 GNDA.n1516 585
R1536 GNDA.n1559 GNDA.n1558 585
R1537 GNDA.n1560 GNDA.n1515 585
R1538 GNDA.n1562 GNDA.n1561 585
R1539 GNDA.n1564 GNDA.n1514 585
R1540 GNDA.n1773 GNDA.n1771 585
R1541 GNDA.n1773 GNDA.n1772 585
R1542 GNDA.n1775 GNDA.n1774 585
R1543 GNDA.n1774 GNDA.n300 585
R1544 GNDA.n1761 GNDA.n1758 585
R1545 GNDA.n1758 GNDA.n299 585
R1546 GNDA.n1782 GNDA.n1781 585
R1547 GNDA.n1783 GNDA.n1782 585
R1548 GNDA.n1759 GNDA.n1756 585
R1549 GNDA.n1784 GNDA.n1756 585
R1550 GNDA.n1787 GNDA.n1786 585
R1551 GNDA.n1786 GNDA.n1785 585
R1552 GNDA.n1755 GNDA.n1020 585
R1553 GNDA.n1757 GNDA.n1755 585
R1554 GNDA.n1754 GNDA.n1753 585
R1555 GNDA.n1754 GNDA.n298 585
R1556 GNDA.n2211 GNDA.n360 585
R1557 GNDA.n360 GNDA.n359 585
R1558 GNDA.n2214 GNDA.n2213 585
R1559 GNDA.n2215 GNDA.n2214 585
R1560 GNDA.n361 GNDA.n357 585
R1561 GNDA.n2216 GNDA.n357 585
R1562 GNDA.n2219 GNDA.n2218 585
R1563 GNDA.n2218 GNDA.n2217 585
R1564 GNDA.n356 GNDA.n354 585
R1565 GNDA.n358 GNDA.n356 585
R1566 GNDA.n350 GNDA.n349 585
R1567 GNDA.n349 GNDA.n296 585
R1568 GNDA.n2227 GNDA.n2226 585
R1569 GNDA.n2227 GNDA.n295 585
R1570 GNDA.n2230 GNDA.n2229 585
R1571 GNDA.n2229 GNDA.n2228 585
R1572 GNDA.n345 GNDA.n343 585
R1573 GNDA.n343 GNDA.n342 585
R1574 GNDA.n2237 GNDA.n2236 585
R1575 GNDA.n2238 GNDA.n2237 585
R1576 GNDA.n379 GNDA.n339 585
R1577 GNDA.n2239 GNDA.n339 585
R1578 GNDA.n2241 GNDA.n340 585
R1579 GNDA.n2241 GNDA.n2240 585
R1580 GNDA.n2210 GNDA.n2209 585
R1581 GNDA.n2209 GNDA.n297 585
R1582 GNDA.n1664 GNDA.n1387 585
R1583 GNDA.n1664 GNDA.n1663 585
R1584 GNDA.n1490 GNDA.n1388 585
R1585 GNDA.n1661 GNDA.n1388 585
R1586 GNDA.n1659 GNDA.n1658 585
R1587 GNDA.n1660 GNDA.n1659 585
R1588 GNDA.n1580 GNDA.n1488 585
R1589 GNDA.n1488 GNDA.n1487 585
R1590 GNDA.n1587 GNDA.n1585 585
R1591 GNDA.n1587 GNDA.n1586 585
R1592 GNDA.n1589 GNDA.n1588 585
R1593 GNDA.n1588 GNDA.n294 585
R1594 GNDA.n1575 GNDA.n1572 585
R1595 GNDA.n1572 GNDA.n293 585
R1596 GNDA.n1596 GNDA.n1595 585
R1597 GNDA.n1597 GNDA.n1596 585
R1598 GNDA.n1573 GNDA.n1512 585
R1599 GNDA.n1598 GNDA.n1512 585
R1600 GNDA.n1601 GNDA.n1600 585
R1601 GNDA.n1600 GNDA.n1599 585
R1602 GNDA.n1511 GNDA.n1509 585
R1603 GNDA.n1570 GNDA.n1569 585
R1604 GNDA.n1666 GNDA.n1665 585
R1605 GNDA.n1665 GNDA.n341 585
R1606 GNDA.n1565 GNDA.n303 585
R1607 GNDA.n1513 GNDA.n303 585
R1608 GNDA.n1696 GNDA.n1695 585
R1609 GNDA.n1699 GNDA.n1698 585
R1610 GNDA.n1700 GNDA.n1033 585
R1611 GNDA.n1033 GNDA.n319 585
R1612 GNDA.n1702 GNDA.n1701 585
R1613 GNDA.n1704 GNDA.n1032 585
R1614 GNDA.n1707 GNDA.n1706 585
R1615 GNDA.n1708 GNDA.n1031 585
R1616 GNDA.n1710 GNDA.n1709 585
R1617 GNDA.n1712 GNDA.n1030 585
R1618 GNDA.n1715 GNDA.n1714 585
R1619 GNDA.n1716 GNDA.n1029 585
R1620 GNDA.n1718 GNDA.n1717 585
R1621 GNDA.n1718 GNDA.n319 585
R1622 GNDA.n2243 GNDA.n2242 585
R1623 GNDA.n1672 GNDA.n1386 585
R1624 GNDA.n1673 GNDA.n1385 585
R1625 GNDA.n1676 GNDA.n1384 585
R1626 GNDA.n1677 GNDA.n1383 585
R1627 GNDA.n1680 GNDA.n1382 585
R1628 GNDA.n1681 GNDA.n1381 585
R1629 GNDA.n1684 GNDA.n1380 585
R1630 GNDA.n1685 GNDA.n1379 585
R1631 GNDA.n1688 GNDA.n1378 585
R1632 GNDA.n1689 GNDA.n332 585
R1633 GNDA.n2243 GNDA.n332 585
R1634 GNDA.n1691 GNDA.n1035 585
R1635 GNDA.n1691 GNDA.n1377 585
R1636 GNDA.n1690 GNDA.n1689 585
R1637 GNDA.n1688 GNDA.n1687 585
R1638 GNDA.n1686 GNDA.n1685 585
R1639 GNDA.n1684 GNDA.n1683 585
R1640 GNDA.n1682 GNDA.n1681 585
R1641 GNDA.n1680 GNDA.n1679 585
R1642 GNDA.n1678 GNDA.n1677 585
R1643 GNDA.n1676 GNDA.n1675 585
R1644 GNDA.n1674 GNDA.n1673 585
R1645 GNDA.n1672 GNDA.n1671 585
R1646 GNDA.n2102 GNDA.n490 585
R1647 GNDA.n2102 GNDA.n496 585
R1648 GNDA.n1175 GNDA.n1173 585
R1649 GNDA.n1176 GNDA.n1046 585
R1650 GNDA.n1179 GNDA.n1045 585
R1651 GNDA.n1180 GNDA.n1044 585
R1652 GNDA.n1183 GNDA.n1043 585
R1653 GNDA.n1184 GNDA.n1042 585
R1654 GNDA.n1187 GNDA.n1041 585
R1655 GNDA.n1188 GNDA.n1040 585
R1656 GNDA.n1191 GNDA.n1039 585
R1657 GNDA.n1192 GNDA.n683 585
R1658 GNDA.n1376 GNDA.n681 585
R1659 GNDA.n1377 GNDA.n1376 585
R1660 GNDA.n1193 GNDA.n1192 585
R1661 GNDA.n1191 GNDA.n1190 585
R1662 GNDA.n1189 GNDA.n1188 585
R1663 GNDA.n1187 GNDA.n1186 585
R1664 GNDA.n1185 GNDA.n1184 585
R1665 GNDA.n1183 GNDA.n1182 585
R1666 GNDA.n1181 GNDA.n1180 585
R1667 GNDA.n1179 GNDA.n1178 585
R1668 GNDA.n1177 GNDA.n1176 585
R1669 GNDA.n1175 GNDA.n1174 585
R1670 GNDA.n1946 GNDA.n1945 585
R1671 GNDA.n684 GNDA.n682 585
R1672 GNDA.n1941 GNDA.n1940 585
R1673 GNDA.n1939 GNDA.n689 585
R1674 GNDA.n1938 GNDA.n1937 585
R1675 GNDA.n1936 GNDA.n1935 585
R1676 GNDA.n1934 GNDA.n1933 585
R1677 GNDA.n1932 GNDA.n1931 585
R1678 GNDA.n1930 GNDA.n1929 585
R1679 GNDA.n1928 GNDA.n1927 585
R1680 GNDA.n1926 GNDA.n1925 585
R1681 GNDA.n1924 GNDA.n1923 585
R1682 GNDA.n1171 GNDA.n1047 585
R1683 GNDA.n1172 GNDA.n1171 585
R1684 GNDA.n1074 GNDA.n1073 585
R1685 GNDA.n1068 GNDA.n1067 585
R1686 GNDA.n1145 GNDA.n1144 585
R1687 GNDA.n1148 GNDA.n1147 585
R1688 GNDA.n1066 GNDA.n1063 585
R1689 GNDA.n1059 GNDA.n1058 585
R1690 GNDA.n1156 GNDA.n1155 585
R1691 GNDA.n1159 GNDA.n1158 585
R1692 GNDA.n1057 GNDA.n1054 585
R1693 GNDA.n1050 GNDA.n1049 585
R1694 GNDA.n1167 GNDA.n1166 585
R1695 GNDA.n1170 GNDA.n1169 585
R1696 GNDA.n1209 GNDA.n303 585
R1697 GNDA.n1206 GNDA.n303 585
R1698 GNDA.n1236 GNDA.n1235 585
R1699 GNDA.n1229 GNDA.n1228 585
R1700 GNDA.n1307 GNDA.n1306 585
R1701 GNDA.n1310 GNDA.n1309 585
R1702 GNDA.n1227 GNDA.n1224 585
R1703 GNDA.n1220 GNDA.n1219 585
R1704 GNDA.n1318 GNDA.n1317 585
R1705 GNDA.n1321 GNDA.n1320 585
R1706 GNDA.n1218 GNDA.n1215 585
R1707 GNDA.n1211 GNDA.n1210 585
R1708 GNDA.n1329 GNDA.n1328 585
R1709 GNDA.n1332 GNDA.n1331 585
R1710 GNDA.n1233 GNDA.n1038 585
R1711 GNDA.n1377 GNDA.n1038 585
R1712 GNDA.n2102 GNDA.n484 585
R1713 GNDA.n2102 GNDA.n497 585
R1714 GNDA.n1898 GNDA.n316 585
R1715 GNDA.n1903 GNDA.n705 585
R1716 GNDA.n1904 GNDA.n704 585
R1717 GNDA.n1907 GNDA.n702 585
R1718 GNDA.n1908 GNDA.n701 585
R1719 GNDA.n1911 GNDA.n699 585
R1720 GNDA.n1912 GNDA.n698 585
R1721 GNDA.n1915 GNDA.n696 585
R1722 GNDA.n1916 GNDA.n695 585
R1723 GNDA.n1919 GNDA.n693 585
R1724 GNDA.n1920 GNDA.n692 585
R1725 GNDA.n692 GNDA.n316 585
R1726 GNDA.n1022 GNDA.n316 585
R1727 GNDA.n1748 GNDA.n1747 585
R1728 GNDA.n1745 GNDA.n1024 585
R1729 GNDA.n1742 GNDA.n1741 585
R1730 GNDA.n1739 GNDA.n1738 585
R1731 GNDA.n1735 GNDA.n1734 585
R1732 GNDA.n1733 GNDA.n1026 585
R1733 GNDA.n1731 GNDA.n1730 585
R1734 GNDA.n1727 GNDA.n1027 585
R1735 GNDA.n1724 GNDA.n1723 585
R1736 GNDA.n1721 GNDA.n854 585
R1737 GNDA.n854 GNDA.n316 585
R1738 GNDA.n1072 GNDA.n1070 585
R1739 GNDA.n1072 GNDA.n690 585
R1740 GNDA.n1922 GNDA.n691 585
R1741 GNDA.n1922 GNDA.n690 585
R1742 GNDA.n1921 GNDA.n1920 585
R1743 GNDA.n1919 GNDA.n1918 585
R1744 GNDA.n1917 GNDA.n1916 585
R1745 GNDA.n1915 GNDA.n1914 585
R1746 GNDA.n1913 GNDA.n1912 585
R1747 GNDA.n1911 GNDA.n1910 585
R1748 GNDA.n1909 GNDA.n1908 585
R1749 GNDA.n1907 GNDA.n1906 585
R1750 GNDA.n1905 GNDA.n1904 585
R1751 GNDA.n1903 GNDA.n1902 585
R1752 GNDA.n2207 GNDA.n448 585
R1753 GNDA.n2207 GNDA.n454 585
R1754 GNDA.n1719 GNDA.n1028 585
R1755 GNDA.n1719 GNDA.n690 585
R1756 GNDA.n1721 GNDA.n1720 585
R1757 GNDA.n1725 GNDA.n1724 585
R1758 GNDA.n1727 GNDA.n1726 585
R1759 GNDA.n1730 GNDA.n1729 585
R1760 GNDA.n1728 GNDA.n1026 585
R1761 GNDA.n1736 GNDA.n1735 585
R1762 GNDA.n1738 GNDA.n1737 585
R1763 GNDA.n1743 GNDA.n1742 585
R1764 GNDA.n1745 GNDA.n1744 585
R1765 GNDA.n1747 GNDA.n1746 585
R1766 GNDA.n2207 GNDA.n442 585
R1767 GNDA.n2208 GNDA.n2207 585
R1768 GNDA.n2199 GNDA.n459 585
R1769 GNDA.n2197 GNDA.n2196 585
R1770 GNDA.n2193 GNDA.n462 585
R1771 GNDA.n2192 GNDA.n2189 585
R1772 GNDA.n2187 GNDA.n463 585
R1773 GNDA.n2185 GNDA.n2184 585
R1774 GNDA.n2181 GNDA.n464 585
R1775 GNDA.n2180 GNDA.n2177 585
R1776 GNDA.n2175 GNDA.n465 585
R1777 GNDA.n2173 GNDA.n2172 585
R1778 GNDA.n2172 GNDA.n2171 585
R1779 GNDA.n2178 GNDA.n465 585
R1780 GNDA.n2180 GNDA.n2179 585
R1781 GNDA.n2182 GNDA.n2181 585
R1782 GNDA.n2184 GNDA.n2183 585
R1783 GNDA.n2190 GNDA.n463 585
R1784 GNDA.n2192 GNDA.n2191 585
R1785 GNDA.n2194 GNDA.n2193 585
R1786 GNDA.n2196 GNDA.n2195 585
R1787 GNDA.n459 GNDA.n458 585
R1788 GNDA.n2095 GNDA.n1971 585
R1789 GNDA.n1969 GNDA.n1966 585
R1790 GNDA.n1965 GNDA.n1964 585
R1791 GNDA.n1963 GNDA.n1960 585
R1792 GNDA.n1959 GNDA.n1958 585
R1793 GNDA.n1957 GNDA.n1954 585
R1794 GNDA.n1953 GNDA.n1952 585
R1795 GNDA.n1951 GNDA.n1949 585
R1796 GNDA.n1948 GNDA.n476 585
R1797 GNDA.n2106 GNDA.n2105 585
R1798 GNDA.n2105 GNDA.n2104 585
R1799 GNDA.n478 GNDA.n476 585
R1800 GNDA.n1951 GNDA.n1950 585
R1801 GNDA.n1955 GNDA.n1952 585
R1802 GNDA.n1957 GNDA.n1956 585
R1803 GNDA.n1961 GNDA.n1958 585
R1804 GNDA.n1963 GNDA.n1962 585
R1805 GNDA.n1967 GNDA.n1964 585
R1806 GNDA.n1969 GNDA.n1968 585
R1807 GNDA.n1971 GNDA.n1970 585
R1808 GNDA.n576 GNDA.n522 585
R1809 GNDA.n574 GNDA.n573 585
R1810 GNDA.n572 GNDA.n523 585
R1811 GNDA.n571 GNDA.n570 585
R1812 GNDA.n568 GNDA.n524 585
R1813 GNDA.n566 GNDA.n565 585
R1814 GNDA.n564 GNDA.n525 585
R1815 GNDA.n563 GNDA.n562 585
R1816 GNDA.n560 GNDA.n526 585
R1817 GNDA.n558 GNDA.n557 585
R1818 GNDA.n2202 GNDA.n460 585
R1819 GNDA.n2202 GNDA.n2201 585
R1820 GNDA.n2097 GNDA.n1972 585
R1821 GNDA.n2097 GNDA.n2096 585
R1822 GNDA.n1998 GNDA.n1997 585
R1823 GNDA.n1994 GNDA.n1993 585
R1824 GNDA.n2069 GNDA.n2068 585
R1825 GNDA.n2072 GNDA.n2071 585
R1826 GNDA.n1992 GNDA.n1989 585
R1827 GNDA.n1985 GNDA.n1984 585
R1828 GNDA.n2080 GNDA.n2079 585
R1829 GNDA.n2083 GNDA.n2082 585
R1830 GNDA.n1983 GNDA.n1980 585
R1831 GNDA.n1976 GNDA.n1975 585
R1832 GNDA.n2091 GNDA.n2090 585
R1833 GNDA.n2094 GNDA.n2093 585
R1834 GNDA.n456 GNDA.n455 585
R1835 GNDA.n690 GNDA.n455 585
R1836 GNDA.n2207 GNDA.n436 585
R1837 GNDA.n2207 GNDA.n2206 585
R1838 GNDA.n521 GNDA.n303 585
R1839 GNDA.n577 GNDA.n303 585
R1840 GNDA.n678 GNDA.n677 585
R1841 GNDA.n675 GNDA.n674 585
R1842 GNDA.n501 GNDA.n500 585
R1843 GNDA.n596 GNDA.n595 585
R1844 GNDA.n603 GNDA.n602 585
R1845 GNDA.n606 GNDA.n605 585
R1846 GNDA.n593 GNDA.n590 585
R1847 GNDA.n586 GNDA.n585 585
R1848 GNDA.n614 GNDA.n613 585
R1849 GNDA.n617 GNDA.n616 585
R1850 GNDA.n584 GNDA.n519 585
R1851 GNDA.n582 GNDA.n581 585
R1852 GNDA.n679 GNDA.n498 585
R1853 GNDA.n1377 GNDA.n498 585
R1854 GNDA.n2102 GNDA.n479 585
R1855 GNDA.n2102 GNDA.n2101 585
R1856 GNDA.n2165 GNDA.n466 585
R1857 GNDA.n2164 GNDA.n2163 585
R1858 GNDA.n2161 GNDA.n2137 585
R1859 GNDA.n2159 GNDA.n2158 585
R1860 GNDA.n2157 GNDA.n2138 585
R1861 GNDA.n2156 GNDA.n2155 585
R1862 GNDA.n2153 GNDA.n2139 585
R1863 GNDA.n2151 GNDA.n2150 585
R1864 GNDA.n2149 GNDA.n2140 585
R1865 GNDA.n2148 GNDA.n2147 585
R1866 GNDA.n2145 GNDA.n2141 585
R1867 GNDA.n2143 GNDA.n2142 585
R1868 GNDA.n2126 GNDA.n2125 585
R1869 GNDA.n2125 GNDA.n2124 585
R1870 GNDA.n2122 GNDA.n2119 585
R1871 GNDA.n2123 GNDA.n2122 585
R1872 GNDA.n2121 GNDA.n2120 585
R1873 GNDA.n2121 GNDA.n315 585
R1874 GNDA.n2109 GNDA.n2108 585
R1875 GNDA.n2110 GNDA.n473 585
R1876 GNDA.n2112 GNDA.n2111 585
R1877 GNDA.n2114 GNDA.n472 585
R1878 GNDA.n2117 GNDA.n2116 585
R1879 GNDA.n2118 GNDA.n471 585
R1880 GNDA.n2129 GNDA.n2128 585
R1881 GNDA.n2131 GNDA.n470 585
R1882 GNDA.n2132 GNDA.n469 585
R1883 GNDA.n2135 GNDA.n2134 585
R1884 GNDA.n2136 GNDA.n468 585
R1885 GNDA.n468 GNDA.n314 585
R1886 GNDA.n2168 GNDA.n2167 585
R1887 GNDA.n2170 GNDA.n467 585
R1888 GNDA.n556 GNDA.n527 585
R1889 GNDA.n555 GNDA.n554 585
R1890 GNDA.n552 GNDA.n528 585
R1891 GNDA.n552 GNDA.n314 585
R1892 GNDA.n551 GNDA.n550 585
R1893 GNDA.n549 GNDA.n548 585
R1894 GNDA.n547 GNDA.n530 585
R1895 GNDA.n545 GNDA.n544 585
R1896 GNDA.n543 GNDA.n531 585
R1897 GNDA.n542 GNDA.n541 585
R1898 GNDA.n539 GNDA.n532 585
R1899 GNDA.n537 GNDA.n536 585
R1900 GNDA.n535 GNDA.n534 585
R1901 GNDA.n477 GNDA.n475 585
R1902 GNDA.n284 GNDA.n283 585
R1903 GNDA.n2244 GNDA.n284 585
R1904 GNDA.n727 GNDA.n725 585
R1905 GNDA.n725 GNDA.n292 585
R1906 GNDA.n830 GNDA.n829 585
R1907 GNDA.n835 GNDA.n830 585
R1908 GNDA.n754 GNDA.n724 585
R1909 GNDA.n836 GNDA.n724 585
R1910 GNDA.n759 GNDA.n723 585
R1911 GNDA.n837 GNDA.n723 585
R1912 GNDA.n763 GNDA.n762 585
R1913 GNDA.n762 GNDA.n312 585
R1914 GNDA.n761 GNDA.n753 585
R1915 GNDA.n761 GNDA.n313 585
R1916 GNDA.n749 GNDA.n719 585
R1917 GNDA.n844 GNDA.n719 585
R1918 GNDA.n770 GNDA.n718 585
R1919 GNDA.n845 GNDA.n718 585
R1920 GNDA.n772 GNDA.n717 585
R1921 GNDA.n846 GNDA.n717 585
R1922 GNDA.n748 GNDA.n747 585
R1923 GNDA.n747 GNDA.n713 585
R1924 GNDA.n712 GNDA.n461 585
R1925 GNDA.n852 GNDA.n712 585
R1926 GNDA.n851 GNDA.n850 585
R1927 GNDA.n852 GNDA.n851 585
R1928 GNDA.n849 GNDA.n714 585
R1929 GNDA.n714 GNDA.n713 585
R1930 GNDA.n848 GNDA.n847 585
R1931 GNDA.n847 GNDA.n846 585
R1932 GNDA.n716 GNDA.n715 585
R1933 GNDA.n845 GNDA.n716 585
R1934 GNDA.n843 GNDA.n842 585
R1935 GNDA.n844 GNDA.n843 585
R1936 GNDA.n841 GNDA.n720 585
R1937 GNDA.n720 GNDA.n313 585
R1938 GNDA.n840 GNDA.n839 585
R1939 GNDA.n839 GNDA.n312 585
R1940 GNDA.n838 GNDA.n721 585
R1941 GNDA.n838 GNDA.n837 585
R1942 GNDA.n831 GNDA.n722 585
R1943 GNDA.n836 GNDA.n722 585
R1944 GNDA.n834 GNDA.n833 585
R1945 GNDA.n835 GNDA.n834 585
R1946 GNDA.n832 GNDA.n290 585
R1947 GNDA.n292 GNDA.n290 585
R1948 GNDA.n2245 GNDA.n291 585
R1949 GNDA.n2245 GNDA.n2244 585
R1950 GNDA.n991 GNDA.n867 585
R1951 GNDA.n867 GNDA.n309 585
R1952 GNDA.n994 GNDA.n993 585
R1953 GNDA.n995 GNDA.n994 585
R1954 GNDA.n894 GNDA.n866 585
R1955 GNDA.n1879 GNDA.n866 585
R1956 GNDA.n892 GNDA.n865 585
R1957 GNDA.n1880 GNDA.n865 585
R1958 GNDA.n900 GNDA.n864 585
R1959 GNDA.n1881 GNDA.n864 585
R1960 GNDA.n904 GNDA.n903 585
R1961 GNDA.n903 GNDA.n310 585
R1962 GNDA.n902 GNDA.n891 585
R1963 GNDA.n902 GNDA.n311 585
R1964 GNDA.n887 GNDA.n860 585
R1965 GNDA.n1888 GNDA.n860 585
R1966 GNDA.n911 GNDA.n859 585
R1967 GNDA.n1889 GNDA.n859 585
R1968 GNDA.n913 GNDA.n858 585
R1969 GNDA.n1890 GNDA.n858 585
R1970 GNDA.n886 GNDA.n711 585
R1971 GNDA.n853 GNDA.n711 585
R1972 GNDA.n1897 GNDA.n709 585
R1973 GNDA.n1897 GNDA.n1896 585
R1974 GNDA.n1895 GNDA.n1894 585
R1975 GNDA.n1896 GNDA.n1895 585
R1976 GNDA.n1893 GNDA.n855 585
R1977 GNDA.n855 GNDA.n853 585
R1978 GNDA.n1892 GNDA.n1891 585
R1979 GNDA.n1891 GNDA.n1890 585
R1980 GNDA.n857 GNDA.n856 585
R1981 GNDA.n1889 GNDA.n857 585
R1982 GNDA.n1887 GNDA.n1886 585
R1983 GNDA.n1888 GNDA.n1887 585
R1984 GNDA.n1885 GNDA.n861 585
R1985 GNDA.n861 GNDA.n311 585
R1986 GNDA.n1884 GNDA.n1883 585
R1987 GNDA.n1883 GNDA.n310 585
R1988 GNDA.n1882 GNDA.n862 585
R1989 GNDA.n1882 GNDA.n1881 585
R1990 GNDA.n997 GNDA.n863 585
R1991 GNDA.n1880 GNDA.n863 585
R1992 GNDA.n1878 GNDA.n1877 585
R1993 GNDA.n1879 GNDA.n1878 585
R1994 GNDA.n1876 GNDA.n996 585
R1995 GNDA.n996 GNDA.n995 585
R1996 GNDA.n1875 GNDA.n1874 585
R1997 GNDA.n1874 GNDA.n309 585
R1998 GNDA.n1850 GNDA.n1849 585
R1999 GNDA.n1002 GNDA.n999 585
R2000 GNDA.n1845 GNDA.n1844 585
R2001 GNDA.n1766 GNDA.n1000 585
R2002 GNDA.n2249 GNDA.n2248 585
R2003 GNDA.n2248 GNDA.n2247 585
R2004 GNDA.n282 GNDA.n281 585
R2005 GNDA.n2247 GNDA.n281 585
R2006 GNDA.n2269 GNDA.n2268 585
R2007 GNDA.n2267 GNDA.n280 585
R2008 GNDA.n2266 GNDA.n279 585
R2009 GNDA.n2271 GNDA.n279 585
R2010 GNDA.n2265 GNDA.n2264 585
R2011 GNDA.n2263 GNDA.n2262 585
R2012 GNDA.n2261 GNDA.n2260 585
R2013 GNDA.n2259 GNDA.n2258 585
R2014 GNDA.n2257 GNDA.n2256 585
R2015 GNDA.n2255 GNDA.n2254 585
R2016 GNDA.n2253 GNDA.n2252 585
R2017 GNDA.n2271 GNDA.n264 585
R2018 GNDA.n990 GNDA.n285 585
R2019 GNDA.n2247 GNDA.n285 585
R2020 GNDA.n2246 GNDA.n289 585
R2021 GNDA.n2247 GNDA.n2246 585
R2022 GNDA.n970 GNDA.n278 585
R2023 GNDA.n2271 GNDA.n278 585
R2024 GNDA.n972 GNDA.n971 585
R2025 GNDA.n974 GNDA.n973 585
R2026 GNDA.n976 GNDA.n975 585
R2027 GNDA.n978 GNDA.n977 585
R2028 GNDA.n980 GNDA.n979 585
R2029 GNDA.n982 GNDA.n981 585
R2030 GNDA.n984 GNDA.n983 585
R2031 GNDA.n986 GNDA.n985 585
R2032 GNDA.n988 GNDA.n987 585
R2033 GNDA.n2271 GNDA.n270 585
R2034 GNDA.n1851 GNDA.n286 585
R2035 GNDA.n2247 GNDA.n286 585
R2036 GNDA.n1873 GNDA.n288 585
R2037 GNDA.n2247 GNDA.n288 585
R2038 GNDA.n1872 GNDA.n277 585
R2039 GNDA.n2271 GNDA.n277 585
R2040 GNDA.n1871 GNDA.n1870 585
R2041 GNDA.n1869 GNDA.n1868 585
R2042 GNDA.n1867 GNDA.n1866 585
R2043 GNDA.n1865 GNDA.n1864 585
R2044 GNDA.n1863 GNDA.n1862 585
R2045 GNDA.n1861 GNDA.n1860 585
R2046 GNDA.n1859 GNDA.n1858 585
R2047 GNDA.n1857 GNDA.n1856 585
R2048 GNDA.n1855 GNDA.n1854 585
R2049 GNDA.n2271 GNDA.n276 585
R2050 GNDA.n1662 GNDA.n1486 556.322
R2051 GNDA.n136 GNDA.t304 535.191
R2052 GNDA.n138 GNDA.t228 535.191
R2053 GNDA.n85 GNDA.t278 535.191
R2054 GNDA.n83 GNDA.t268 535.191
R2055 GNDA.n248 GNDA.n244 531.201
R2056 GNDA.n253 GNDA.n244 528
R2057 GNDA.n2244 GNDA.t224 512.884
R2058 GNDA.t224 GNDA.n309 512.884
R2059 GNDA.n2329 GNDA.n218 512
R2060 GNDA.n2327 GNDA.n218 512
R2061 GNDA.n1482 GNDA.n1392 512
R2062 GNDA.n1484 GNDA.n1392 512
R2063 GNDA.n1393 GNDA.n212 511.39
R2064 GNDA.n2329 GNDA.n2328 508.8
R2065 GNDA.n2328 GNDA.n2327 508.8
R2066 GNDA.n1483 GNDA.n1482 508.8
R2067 GNDA.n1484 GNDA.n1483 508.8
R2068 GNDA.n248 GNDA.n247 499.2
R2069 GNDA.n180 GNDA.n147 496
R2070 GNDA.n2383 GNDA.n2382 496
R2071 GNDA.n64 GNDA.t238 493.418
R2072 GNDA.n70 GNDA.t225 493.418
R2073 GNDA.n69 GNDA.t295 493.418
R2074 GNDA.n68 GNDA.t311 493.418
R2075 GNDA.n67 GNDA.t292 493.418
R2076 GNDA.n66 GNDA.t281 493.418
R2077 GNDA.n2391 GNDA.t307 493.418
R2078 GNDA.n2392 GNDA.t289 493.418
R2079 GNDA.n2393 GNDA.t301 493.418
R2080 GNDA.n2394 GNDA.t286 493.418
R2081 GNDA.n181 GNDA.n180 489.601
R2082 GNDA.n2382 GNDA.n2377 489.601
R2083 GNDA.n253 GNDA.n232 486.401
R2084 GNDA.t102 GNDA.n237 451.531
R2085 GNDA.n2303 GNDA.n2302 444.8
R2086 GNDA.n2302 GNDA.n2301 444.8
R2087 GNDA.n2303 GNDA.n2298 441.601
R2088 GNDA.n2301 GNDA.n2299 438.401
R2089 GNDA.n235 GNDA.n230 435.2
R2090 GNDA.t224 GNDA.n297 434.906
R2091 GNDA.n2416 GNDA.n2415 428.8
R2092 GNDA.n2309 GNDA.n230 425.601
R2093 GNDA.n77 GNDA.n76 422.401
R2094 GNDA.n72 GNDA.n71 422.401
R2095 GNDA.n2396 GNDA.n2395 422.401
R2096 GNDA.n2399 GNDA.n2398 422.401
R2097 GNDA.n2308 GNDA.n233 422.401
R2098 GNDA.n2309 GNDA.n2308 419.2
R2099 GNDA.n1411 GNDA.t283 413.084
R2100 GNDA.n1414 GNDA.t298 413.084
R2101 GNDA.n1410 GNDA.t261 413.084
R2102 GNDA.n1408 GNDA.t245 413.084
R2103 GNDA.n1443 GNDA.t274 413.084
R2104 GNDA.n1438 GNDA.t271 413.084
R2105 GNDA.n2386 GNDA.n2385 396.17
R2106 GNDA.n145 GNDA.n142 396.17
R2107 GNDA.t224 GNDA.n312 391.411
R2108 GNDA.t224 GNDA.n310 391.411
R2109 GNDA.n132 GNDA.n127 387.2
R2110 GNDA.n2369 GNDA.n2366 387.2
R2111 GNDA.n222 GNDA.n220 383.118
R2112 GNDA.n186 GNDA.n127 380.8
R2113 GNDA.n2370 GNDA.n2369 380.8
R2114 GNDA.t287 GNDA.t65 372.308
R2115 GNDA.t23 GNDA.t65 372.308
R2116 GNDA.t23 GNDA.t314 372.308
R2117 GNDA.t314 GNDA.t44 372.308
R2118 GNDA.t44 GNDA.t166 372.308
R2119 GNDA.t126 GNDA.t131 372.308
R2120 GNDA.t131 GNDA.t316 372.308
R2121 GNDA.t57 GNDA.t94 372.308
R2122 GNDA.t94 GNDA.t308 372.308
R2123 GNDA.n2410 GNDA.n33 371.2
R2124 GNDA.n2415 GNDA.n2414 371.2
R2125 GNDA.t224 GNDA.n303 72.949
R2126 GNDA.t32 GNDA.n37 355.385
R2127 GNDA.t59 GNDA.n28 355.385
R2128 GNDA.t316 GNDA.n29 355.385
R2129 GNDA.n1421 GNDA.n1389 354.024
R2130 GNDA.n1599 GNDA.n1598 352.627
R2131 GNDA.n1598 GNDA.n1597 352.627
R2132 GNDA.n1597 GNDA.n293 352.627
R2133 GNDA.n1586 GNDA.n294 352.627
R2134 GNDA.n1586 GNDA.n1487 352.627
R2135 GNDA.n1660 GNDA.n1487 352.627
R2136 GNDA.n1661 GNDA.n1660 352.627
R2137 GNDA.n1663 GNDA.n341 352.627
R2138 GNDA.n2240 GNDA.n2239 352.627
R2139 GNDA.n2239 GNDA.n2238 352.627
R2140 GNDA.n2238 GNDA.n342 352.627
R2141 GNDA.n2228 GNDA.n342 352.627
R2142 GNDA.n2228 GNDA.n295 352.627
R2143 GNDA.n358 GNDA.n296 352.627
R2144 GNDA.n2217 GNDA.n358 352.627
R2145 GNDA.n2217 GNDA.n2216 352.627
R2146 GNDA.n2216 GNDA.n2215 352.627
R2147 GNDA.n2215 GNDA.n359 352.627
R2148 GNDA.n359 GNDA.n297 352.627
R2149 GNDA.n1757 GNDA.n298 352.627
R2150 GNDA.n1785 GNDA.n1757 352.627
R2151 GNDA.n1785 GNDA.n1784 352.627
R2152 GNDA.n1784 GNDA.n1783 352.627
R2153 GNDA.n1783 GNDA.n299 352.627
R2154 GNDA.n1772 GNDA.n300 352.627
R2155 GNDA.n188 GNDA.n122 348.8
R2156 GNDA.n2356 GNDA.n99 348.8
R2157 GNDA.n195 GNDA.n123 342.401
R2158 GNDA.n2360 GNDA.n100 342.401
R2159 GNDA.n1442 GNDA.n215 341.38
R2160 GNDA.n203 GNDA.n114 332.8
R2161 GNDA.n2348 GNDA.n88 332.8
R2162 GNDA.n51 GNDA.t255 332.75
R2163 GNDA.n52 GNDA.t258 332.75
R2164 GNDA.t224 GNDA.n301 172.876
R2165 GNDA.t224 GNDA.n304 172.876
R2166 GNDA.t224 GNDA.n302 172.615
R2167 GNDA.t224 GNDA.n305 172.615
R2168 GNDA.n1428 GNDA.n1427 323.2
R2169 GNDA.n222 GNDA.n221 322.861
R2170 GNDA.n205 GNDA.n204 321.281
R2171 GNDA.n2375 GNDA.n89 321.281
R2172 GNDA.n196 GNDA.n195 320
R2173 GNDA.n2355 GNDA.n100 320
R2174 GNDA.n2294 GNDA.n106 318.622
R2175 GNDA.n204 GNDA.n203 318.08
R2176 GNDA.n2348 GNDA.n89 318.08
R2177 GNDA.n1427 GNDA.n223 316.8
R2178 GNDA.n147 GNDA.n141 310.401
R2179 GNDA.n2383 GNDA.n84 310.401
R2180 GNDA.n181 GNDA.n137 304
R2181 GNDA.n2291 GNDA.n2290 304
R2182 GNDA.n2377 GNDA.n86 304
R2183 GNDA.n57 GNDA.n41 300.8
R2184 GNDA.n57 GNDA.n56 300.8
R2185 GNDA.n114 GNDA.n113 300.8
R2186 GNDA.n2290 GNDA.n2289 300.8
R2187 GNDA.n2291 GNDA.n254 300.8
R2188 GNDA.n2376 GNDA.n88 300.8
R2189 GNDA.n1393 GNDA.n107 299.781
R2190 GNDA.n2289 GNDA.n254 297.601
R2191 GNDA.n2276 GNDA.n2275 297.601
R2192 GNDA.n2284 GNDA.n2276 297.601
R2193 GNDA.n2283 GNDA.n2278 297.601
R2194 GNDA.n2278 GNDA.n229 297.601
R2195 GNDA.n198 GNDA.n120 296
R2196 GNDA.n2353 GNDA.n104 296
R2197 GNDA.n1437 GNDA.n1436 294.401
R2198 GNDA.n1475 GNDA.n1437 294.401
R2199 GNDA.n1429 GNDA.n1428 294.401
R2200 GNDA.n203 GNDA.n202 292.5
R2201 GNDA.n202 GNDA.n201 292.5
R2202 GNDA.n204 GNDA.n112 292.5
R2203 GNDA.n117 GNDA.n112 292.5
R2204 GNDA.n114 GNDA.n111 292.5
R2205 GNDA.n117 GNDA.n111 292.5
R2206 GNDA.n195 GNDA.n194 292.5
R2207 GNDA.n194 GNDA.n109 292.5
R2208 GNDA.n193 GNDA.n123 292.5
R2209 GNDA.n193 GNDA.n192 292.5
R2210 GNDA.n189 GNDA.n188 292.5
R2211 GNDA.n189 GNDA.n115 292.5
R2212 GNDA.n124 GNDA.n122 292.5
R2213 GNDA.n192 GNDA.n124 292.5
R2214 GNDA.n199 GNDA.n198 292.5
R2215 GNDA.n200 GNDA.n199 292.5
R2216 GNDA.n1426 GNDA.n223 292.5
R2217 GNDA.n1426 GNDA.n1425 292.5
R2218 GNDA.n1427 GNDA.n1418 292.5
R2219 GNDA.n1431 GNDA.n1418 292.5
R2220 GNDA.n1428 GNDA.n1422 292.5
R2221 GNDA.n1422 GNDA.n1421 292.5
R2222 GNDA.n1430 GNDA.n1429 292.5
R2223 GNDA.n1431 GNDA.n1430 292.5
R2224 GNDA.n1442 GNDA.n220 292.5
R2225 GNDA.n1471 GNDA.n221 292.5
R2226 GNDA.n2323 GNDA.n2322 292.5
R2227 GNDA.n2324 GNDA.n2323 292.5
R2228 GNDA.n1482 GNDA.n1481 292.5
R2229 GNDA.n1481 GNDA.n1480 292.5
R2230 GNDA.n1483 GNDA.n1391 292.5
R2231 GNDA.n1431 GNDA.n1391 292.5
R2232 GNDA.n1485 GNDA.n1484 292.5
R2233 GNDA.n1486 GNDA.n1485 292.5
R2234 GNDA.n1392 GNDA.n1390 292.5
R2235 GNDA.n1431 GNDA.n1390 292.5
R2236 GNDA.n2330 GNDA.n2329 292.5
R2237 GNDA.n2331 GNDA.n2330 292.5
R2238 GNDA.n2328 GNDA.n217 292.5
R2239 GNDA.n1471 GNDA.n217 292.5
R2240 GNDA.n2327 GNDA.n2326 292.5
R2241 GNDA.n2326 GNDA.n2325 292.5
R2242 GNDA.n218 GNDA.n216 292.5
R2243 GNDA.n1471 GNDA.n216 292.5
R2244 GNDA.n1403 GNDA.n1401 292.5
R2245 GNDA.n1401 GNDA.n215 292.5
R2246 GNDA.n1399 GNDA.n224 292.5
R2247 GNDA.n1479 GNDA.n1399 292.5
R2248 GNDA.n1402 GNDA.n1400 292.5
R2249 GNDA.n1400 GNDA.n1389 292.5
R2250 GNDA.n1405 GNDA.n1404 292.5
R2251 GNDA.n1479 GNDA.n1405 292.5
R2252 GNDA.n1435 GNDA.n1413 292.5
R2253 GNDA.n1423 GNDA.n1413 292.5
R2254 GNDA.n1434 GNDA.n1433 292.5
R2255 GNDA.n1433 GNDA.n1432 292.5
R2256 GNDA.n1419 GNDA.n1416 292.5
R2257 GNDA.n1420 GNDA.n1419 292.5
R2258 GNDA.n1475 GNDA.n1407 292.5
R2259 GNDA.n1407 GNDA.n219 292.5
R2260 GNDA.n1437 GNDA.n1398 292.5
R2261 GNDA.n1479 GNDA.n1398 292.5
R2262 GNDA.n1436 GNDA.n1406 292.5
R2263 GNDA.n1424 GNDA.n1406 292.5
R2264 GNDA.n1478 GNDA.n1477 292.5
R2265 GNDA.n1479 GNDA.n1478 292.5
R2266 GNDA.n1467 GNDA.n1466 292.5
R2267 GNDA.n1468 GNDA.n1467 292.5
R2268 GNDA.n1469 GNDA.n1440 292.5
R2269 GNDA.n1470 GNDA.n1469 292.5
R2270 GNDA.n1474 GNDA.n1473 292.5
R2271 GNDA.n1473 GNDA.n1472 292.5
R2272 GNDA.n2283 GNDA.n2282 292.5
R2273 GNDA.n2282 GNDA.n241 292.5
R2274 GNDA.n2290 GNDA.n243 292.5
R2275 GNDA.n255 GNDA.n243 292.5
R2276 GNDA.n2292 GNDA.n2291 292.5
R2277 GNDA.n2293 GNDA.n2292 292.5
R2278 GNDA.n254 GNDA.n242 292.5
R2279 GNDA.n255 GNDA.n242 292.5
R2280 GNDA.n2289 GNDA.n2288 292.5
R2281 GNDA.n2288 GNDA.n2287 292.5
R2282 GNDA.n2276 GNDA.n257 292.5
R2283 GNDA.n2272 GNDA.n257 292.5
R2284 GNDA.n2285 GNDA.n2284 292.5
R2285 GNDA.n2286 GNDA.n2285 292.5
R2286 GNDA.n258 GNDA.n256 292.5
R2287 GNDA.n2272 GNDA.n256 292.5
R2288 GNDA.n2275 GNDA.n2274 292.5
R2289 GNDA.n2274 GNDA.n2273 292.5
R2290 GNDA.n2304 GNDA.n2303 292.5
R2291 GNDA.n2305 GNDA.n2304 292.5
R2292 GNDA.n2302 GNDA.n2297 292.5
R2293 GNDA.n2297 GNDA.n2296 292.5
R2294 GNDA.n2301 GNDA.n2300 292.5
R2295 GNDA.n2300 GNDA.n105 292.5
R2296 GNDA.n2298 GNDA.n239 292.5
R2297 GNDA.n2296 GNDA.n239 292.5
R2298 GNDA.n2308 GNDA.n2307 292.5
R2299 GNDA.n2307 GNDA.n2306 292.5
R2300 GNDA.n236 GNDA.n235 292.5
R2301 GNDA.n240 GNDA.n236 292.5
R2302 GNDA.n234 GNDA.n230 292.5
R2303 GNDA.n234 GNDA.n105 292.5
R2304 GNDA.n2309 GNDA.n231 292.5
R2305 GNDA.n240 GNDA.n231 292.5
R2306 GNDA.n246 GNDA.n244 292.5
R2307 GNDA.n250 GNDA.n246 292.5
R2308 GNDA.n249 GNDA.n248 292.5
R2309 GNDA.n251 GNDA.n249 292.5
R2310 GNDA.n247 GNDA.n245 292.5
R2311 GNDA.n245 GNDA.n238 292.5
R2312 GNDA.n253 GNDA.n252 292.5
R2313 GNDA.n252 GNDA.n251 292.5
R2314 GNDA.n2281 GNDA.n2278 292.5
R2315 GNDA.n2281 GNDA.n237 292.5
R2316 GNDA.n2280 GNDA.n229 292.5
R2317 GNDA.n2280 GNDA.n240 292.5
R2318 GNDA.n2279 GNDA.n2277 292.5
R2319 GNDA.n2279 GNDA.n106 292.5
R2320 GNDA.n2375 GNDA.n2374 292.5
R2321 GNDA.n2374 GNDA.n2373 292.5
R2322 GNDA.n91 GNDA.n89 292.5
R2323 GNDA.n2344 GNDA.n91 292.5
R2324 GNDA.n2349 GNDA.n2348 292.5
R2325 GNDA.n2350 GNDA.n2349 292.5
R2326 GNDA.n90 GNDA.n88 292.5
R2327 GNDA.n2344 GNDA.n90 292.5
R2328 GNDA.n2357 GNDA.n2356 292.5
R2329 GNDA.n2358 GNDA.n2357 292.5
R2330 GNDA.n102 GNDA.n99 292.5
R2331 GNDA.n2347 GNDA.n102 292.5
R2332 GNDA.n2360 GNDA.n2359 292.5
R2333 GNDA.n2359 GNDA.n2358 292.5
R2334 GNDA.n101 GNDA.n100 292.5
R2335 GNDA.n2340 GNDA.n101 292.5
R2336 GNDA.n2353 GNDA.n2352 292.5
R2337 GNDA.n2352 GNDA.n2351 292.5
R2338 GNDA.n2401 GNDA.n2400 292.5
R2339 GNDA.n2400 GNDA.n30 292.5
R2340 GNDA.n2390 GNDA.n2389 292.5
R2341 GNDA.n2389 GNDA.n2388 292.5
R2342 GNDA.n2397 GNDA.n59 292.5
R2343 GNDA.n2405 GNDA.n59 292.5
R2344 GNDA.n56 GNDA.n40 292.5
R2345 GNDA.n40 GNDA.n28 292.5
R2346 GNDA.n58 GNDA.n57 292.5
R2347 GNDA.n2405 GNDA.n58 292.5
R2348 GNDA.n41 GNDA.n39 292.5
R2349 GNDA.n39 GNDA.n37 292.5
R2350 GNDA.n54 GNDA.n38 292.5
R2351 GNDA.n2405 GNDA.n38 292.5
R2352 GNDA.n2418 GNDA.n2417 292.5
R2353 GNDA.n2419 GNDA.n2418 292.5
R2354 GNDA.n2415 GNDA.n32 292.5
R2355 GNDA.n2405 GNDA.n32 292.5
R2356 GNDA.n2414 GNDA.n2413 292.5
R2357 GNDA.n2413 GNDA.n2412 292.5
R2358 GNDA.n2409 GNDA.n36 292.5
R2359 GNDA.n2387 GNDA.n36 292.5
R2360 GNDA.n2411 GNDA.n2410 292.5
R2361 GNDA.n2412 GNDA.n2411 292.5
R2362 GNDA.n33 GNDA.n31 292.5
R2363 GNDA.n2405 GNDA.n31 292.5
R2364 GNDA.n2384 GNDA.n2383 292.5
R2365 GNDA.n2385 GNDA.n2384 292.5
R2366 GNDA.n2382 GNDA.n82 292.5
R2367 GNDA.n95 GNDA.n82 292.5
R2368 GNDA.n2377 GNDA.n87 292.5
R2369 GNDA.n93 GNDA.n87 292.5
R2370 GNDA.n2367 GNDA.n81 292.5
R2371 GNDA.n95 GNDA.n81 292.5
R2372 GNDA.n206 GNDA.n205 292.5
R2373 GNDA.n207 GNDA.n206 292.5
R2374 GNDA.n182 GNDA.n181 292.5
R2375 GNDA.n183 GNDA.n182 292.5
R2376 GNDA.n180 GNDA.n135 292.5
R2377 GNDA.n143 GNDA.n135 292.5
R2378 GNDA.n147 GNDA.n146 292.5
R2379 GNDA.n146 GNDA.n145 292.5
R2380 GNDA.n140 GNDA.n134 292.5
R2381 GNDA.n143 GNDA.n134 292.5
R2382 GNDA.n75 GNDA.n63 292.5
R2383 GNDA.n142 GNDA.n63 292.5
R2384 GNDA.n74 GNDA.n61 292.5
R2385 GNDA.n2405 GNDA.n61 292.5
R2386 GNDA.n73 GNDA.n62 292.5
R2387 GNDA.n2386 GNDA.n62 292.5
R2388 GNDA.n2404 GNDA.n2403 292.5
R2389 GNDA.n2405 GNDA.n2404 292.5
R2390 GNDA.n2366 GNDA.n2365 292.5
R2391 GNDA.n2365 GNDA.n80 292.5
R2392 GNDA.n2369 GNDA.n96 292.5
R2393 GNDA.n96 GNDA.t28 292.5
R2394 GNDA.n2371 GNDA.n2370 292.5
R2395 GNDA.n2372 GNDA.n2371 292.5
R2396 GNDA.n2363 GNDA.n94 292.5
R2397 GNDA.t28 GNDA.n94 292.5
R2398 GNDA.n186 GNDA.n185 292.5
R2399 GNDA.n185 GNDA.n110 292.5
R2400 GNDA.n184 GNDA.n127 292.5
R2401 GNDA.n184 GNDA.t33 292.5
R2402 GNDA.n133 GNDA.n132 292.5
R2403 GNDA.n144 GNDA.n133 292.5
R2404 GNDA.n130 GNDA.n128 292.5
R2405 GNDA.t33 GNDA.n128 292.5
R2406 GNDA.n2402 GNDA.n60 292.5
R2407 GNDA.n2405 GNDA.n60 292.5
R2408 GNDA.n2422 GNDA.n2421 292.5
R2409 GNDA.n2421 GNDA.n2420 292.5
R2410 GNDA.n26 GNDA.n25 292.5
R2411 GNDA.n2405 GNDA.n26 292.5
R2412 GNDA.n2407 GNDA.n2406 292.5
R2413 GNDA.n2408 GNDA.n2407 292.5
R2414 GNDA.n27 GNDA.n24 292.5
R2415 GNDA.n2405 GNDA.n27 292.5
R2416 GNDA.n2275 GNDA.n258 291.2
R2417 GNDA.n2284 GNDA.n258 291.2
R2418 GNDA.n2283 GNDA.n2277 291.2
R2419 GNDA.n2277 GNDA.n229 291.2
R2420 GNDA.n1429 GNDA.n223 288
R2421 GNDA.n1415 GNDA.n1412 281.601
R2422 GNDA.n1444 GNDA.n1439 281.601
R2423 GNDA.n1434 GNDA.n1416 278.401
R2424 GNDA.n1466 GNDA.n1440 278.401
R2425 GNDA.n250 GNDA.n107 267.034
R2426 GNDA.n2331 GNDA.n215 265.517
R2427 GNDA.n533 GNDA.n314 264.301
R2428 GNDA.n2169 GNDA.n314 264.301
R2429 GNDA.n582 GNDA.n521 259.416
R2430 GNDA.n2093 GNDA.n1972 259.416
R2431 GNDA.n1898 GNDA.n1897 259.416
R2432 GNDA.n2242 GNDA.n2241 259.416
R2433 GNDA.n1754 GNDA.n1022 259.416
R2434 GNDA.n1331 GNDA.n1209 259.416
R2435 GNDA.n1570 GNDA.n1513 259.416
R2436 GNDA.n1169 GNDA.n1047 259.416
R2437 GNDA.n712 GNDA.n460 259.416
R2438 GNDA.n51 GNDA.t257 258.601
R2439 GNDA.n52 GNDA.t260 258.601
R2440 GNDA.n1567 GNDA.n1566 254.494
R2441 GNDA.n1333 GNDA.n1207 254.392
R2442 GNDA.n579 GNDA.n578 254.392
R2443 GNDA.n1352 GNDA.n302 254.34
R2444 GNDA.n1358 GNDA.n302 254.34
R2445 GNDA.n1360 GNDA.n302 254.34
R2446 GNDA.n1366 GNDA.n302 254.34
R2447 GNDA.n1368 GNDA.n302 254.34
R2448 GNDA.n1374 GNDA.n302 254.34
R2449 GNDA.n1336 GNDA.n303 254.34
R2450 GNDA.n1205 GNDA.n303 254.34
R2451 GNDA.n1343 GNDA.n303 254.34
R2452 GNDA.n1202 GNDA.n303 254.34
R2453 GNDA.n1350 GNDA.n303 254.34
R2454 GNDA.n1521 GNDA.n305 254.34
R2455 GNDA.n1540 GNDA.n305 254.34
R2456 GNDA.n1524 GNDA.n305 254.34
R2457 GNDA.n1533 GNDA.n305 254.34
R2458 GNDA.n1526 GNDA.n305 254.34
R2459 GNDA.n1037 GNDA.n305 254.34
R2460 GNDA.n1547 GNDA.n303 254.34
R2461 GNDA.n1549 GNDA.n303 254.34
R2462 GNDA.n1555 GNDA.n303 254.34
R2463 GNDA.n1557 GNDA.n303 254.34
R2464 GNDA.n1563 GNDA.n303 254.34
R2465 GNDA.n1697 GNDA.n319 254.34
R2466 GNDA.n1703 GNDA.n319 254.34
R2467 GNDA.n1705 GNDA.n319 254.34
R2468 GNDA.n1711 GNDA.n319 254.34
R2469 GNDA.n1713 GNDA.n319 254.34
R2470 GNDA.n1669 GNDA.n338 254.34
R2471 GNDA.n2243 GNDA.n337 254.34
R2472 GNDA.n2243 GNDA.n336 254.34
R2473 GNDA.n2243 GNDA.n335 254.34
R2474 GNDA.n2243 GNDA.n334 254.34
R2475 GNDA.n2243 GNDA.n333 254.34
R2476 GNDA.n2102 GNDA.n495 254.34
R2477 GNDA.n2102 GNDA.n494 254.34
R2478 GNDA.n2102 GNDA.n493 254.34
R2479 GNDA.n2102 GNDA.n492 254.34
R2480 GNDA.n2102 GNDA.n491 254.34
R2481 GNDA.n1668 GNDA.n1667 254.34
R2482 GNDA.n2243 GNDA.n331 254.34
R2483 GNDA.n2243 GNDA.n330 254.34
R2484 GNDA.n2243 GNDA.n329 254.34
R2485 GNDA.n2243 GNDA.n328 254.34
R2486 GNDA.n2243 GNDA.n327 254.34
R2487 GNDA.n2102 GNDA.n489 254.34
R2488 GNDA.n2102 GNDA.n488 254.34
R2489 GNDA.n2102 GNDA.n487 254.34
R2490 GNDA.n2102 GNDA.n486 254.34
R2491 GNDA.n2102 GNDA.n485 254.34
R2492 GNDA.n1944 GNDA.n1943 254.34
R2493 GNDA.n1943 GNDA.n1942 254.34
R2494 GNDA.n1943 GNDA.n688 254.34
R2495 GNDA.n1943 GNDA.n687 254.34
R2496 GNDA.n1943 GNDA.n686 254.34
R2497 GNDA.n1943 GNDA.n685 254.34
R2498 GNDA.n2243 GNDA.n326 254.34
R2499 GNDA.n1071 GNDA.n307 254.34
R2500 GNDA.n1146 GNDA.n307 254.34
R2501 GNDA.n1065 GNDA.n307 254.34
R2502 GNDA.n1157 GNDA.n307 254.34
R2503 GNDA.n1056 GNDA.n307 254.34
R2504 GNDA.n1168 GNDA.n307 254.34
R2505 GNDA.n1234 GNDA.n304 254.34
R2506 GNDA.n1308 GNDA.n304 254.34
R2507 GNDA.n1226 GNDA.n304 254.34
R2508 GNDA.n1319 GNDA.n304 254.34
R2509 GNDA.n1217 GNDA.n304 254.34
R2510 GNDA.n1330 GNDA.n304 254.34
R2511 GNDA.n1232 GNDA.n1231 254.34
R2512 GNDA.n1900 GNDA.n1899 254.34
R2513 GNDA.n710 GNDA.n316 254.34
R2514 GNDA.n703 GNDA.n316 254.34
R2515 GNDA.n700 GNDA.n316 254.34
R2516 GNDA.n697 GNDA.n316 254.34
R2517 GNDA.n694 GNDA.n316 254.34
R2518 GNDA.n1751 GNDA.n1750 254.34
R2519 GNDA.n1749 GNDA.n316 254.34
R2520 GNDA.n1740 GNDA.n316 254.34
R2521 GNDA.n1025 GNDA.n316 254.34
R2522 GNDA.n1732 GNDA.n316 254.34
R2523 GNDA.n1722 GNDA.n316 254.34
R2524 GNDA.n2207 GNDA.n453 254.34
R2525 GNDA.n2207 GNDA.n452 254.34
R2526 GNDA.n2207 GNDA.n451 254.34
R2527 GNDA.n2207 GNDA.n450 254.34
R2528 GNDA.n2207 GNDA.n449 254.34
R2529 GNDA.n708 GNDA.n707 254.34
R2530 GNDA.n2207 GNDA.n447 254.34
R2531 GNDA.n2207 GNDA.n446 254.34
R2532 GNDA.n2207 GNDA.n445 254.34
R2533 GNDA.n2207 GNDA.n444 254.34
R2534 GNDA.n2207 GNDA.n443 254.34
R2535 GNDA.n435 GNDA.n434 254.34
R2536 GNDA.n2198 GNDA.n316 254.34
R2537 GNDA.n2188 GNDA.n316 254.34
R2538 GNDA.n2186 GNDA.n316 254.34
R2539 GNDA.n2176 GNDA.n316 254.34
R2540 GNDA.n2174 GNDA.n316 254.34
R2541 GNDA.n2207 GNDA.n441 254.34
R2542 GNDA.n2207 GNDA.n440 254.34
R2543 GNDA.n2207 GNDA.n439 254.34
R2544 GNDA.n2207 GNDA.n438 254.34
R2545 GNDA.n2207 GNDA.n437 254.34
R2546 GNDA.n2243 GNDA.n325 254.34
R2547 GNDA.n2243 GNDA.n324 254.34
R2548 GNDA.n2243 GNDA.n323 254.34
R2549 GNDA.n2243 GNDA.n322 254.34
R2550 GNDA.n2243 GNDA.n321 254.34
R2551 GNDA.n2103 GNDA.n2102 254.34
R2552 GNDA.n2102 GNDA.n483 254.34
R2553 GNDA.n2102 GNDA.n482 254.34
R2554 GNDA.n2102 GNDA.n481 254.34
R2555 GNDA.n2102 GNDA.n480 254.34
R2556 GNDA.n575 GNDA.n303 254.34
R2557 GNDA.n569 GNDA.n303 254.34
R2558 GNDA.n567 GNDA.n303 254.34
R2559 GNDA.n561 GNDA.n303 254.34
R2560 GNDA.n559 GNDA.n303 254.34
R2561 GNDA.n2200 GNDA.n316 254.34
R2562 GNDA.n2243 GNDA.n320 254.34
R2563 GNDA.n1996 GNDA.n1974 254.34
R2564 GNDA.n2070 GNDA.n1974 254.34
R2565 GNDA.n1991 GNDA.n1974 254.34
R2566 GNDA.n2081 GNDA.n1974 254.34
R2567 GNDA.n1982 GNDA.n1974 254.34
R2568 GNDA.n2092 GNDA.n1974 254.34
R2569 GNDA.n2205 GNDA.n2204 254.34
R2570 GNDA.n676 GNDA.n301 254.34
R2571 GNDA.n594 GNDA.n301 254.34
R2572 GNDA.n604 GNDA.n301 254.34
R2573 GNDA.n592 GNDA.n301 254.34
R2574 GNDA.n615 GNDA.n301 254.34
R2575 GNDA.n583 GNDA.n301 254.34
R2576 GNDA.n2100 GNDA.n2099 254.34
R2577 GNDA.n2162 GNDA.n314 254.34
R2578 GNDA.n2160 GNDA.n314 254.34
R2579 GNDA.n2154 GNDA.n314 254.34
R2580 GNDA.n2152 GNDA.n314 254.34
R2581 GNDA.n2146 GNDA.n314 254.34
R2582 GNDA.n2144 GNDA.n314 254.34
R2583 GNDA.n2107 GNDA.n314 254.34
R2584 GNDA.n2113 GNDA.n314 254.34
R2585 GNDA.n2115 GNDA.n314 254.34
R2586 GNDA.n2130 GNDA.n314 254.34
R2587 GNDA.n2133 GNDA.n314 254.34
R2588 GNDA.n553 GNDA.n314 254.34
R2589 GNDA.n529 GNDA.n314 254.34
R2590 GNDA.n546 GNDA.n314 254.34
R2591 GNDA.n540 GNDA.n314 254.34
R2592 GNDA.n538 GNDA.n314 254.34
R2593 GNDA.n1848 GNDA.n1847 254.34
R2594 GNDA.n1847 GNDA.n1846 254.34
R2595 GNDA.n2271 GNDA.n2270 254.34
R2596 GNDA.n2271 GNDA.n260 254.34
R2597 GNDA.n2271 GNDA.n261 254.34
R2598 GNDA.n2271 GNDA.n262 254.34
R2599 GNDA.n2271 GNDA.n263 254.34
R2600 GNDA.n2251 GNDA.n2250 254.34
R2601 GNDA.n2271 GNDA.n265 254.34
R2602 GNDA.n2271 GNDA.n266 254.34
R2603 GNDA.n2271 GNDA.n267 254.34
R2604 GNDA.n2271 GNDA.n268 254.34
R2605 GNDA.n2271 GNDA.n269 254.34
R2606 GNDA.n989 GNDA.n969 254.34
R2607 GNDA.n2271 GNDA.n271 254.34
R2608 GNDA.n2271 GNDA.n272 254.34
R2609 GNDA.n2271 GNDA.n273 254.34
R2610 GNDA.n2271 GNDA.n274 254.34
R2611 GNDA.n2271 GNDA.n275 254.34
R2612 GNDA.n1853 GNDA.n1852 254.34
R2613 GNDA.n1486 GNDA.n1389 252.875
R2614 GNDA.n558 GNDA.n527 249.663
R2615 GNDA.n851 GNDA.n692 249.663
R2616 GNDA.n1696 GNDA.n332 249.663
R2617 GNDA.n1895 GNDA.n854 249.663
R2618 GNDA.n1353 GNDA.n1351 249.663
R2619 GNDA.n1546 GNDA.n1519 249.663
R2620 GNDA.n1945 GNDA.n683 249.663
R2621 GNDA.n2173 GNDA.n466 249.663
R2622 GNDA.n2108 GNDA.n2106 249.663
R2623 GNDA.n187 GNDA.n123 246.4
R2624 GNDA.n2361 GNDA.n2360 246.4
R2625 GNDA.n1435 GNDA.n1434 240
R2626 GNDA.n1474 GNDA.n1440 240
R2627 GNDA.t224 GNDA.n293 239.004
R2628 GNDA.n1662 GNDA.n1661 239.004
R2629 GNDA.t224 GNDA.n295 239.004
R2630 GNDA.t224 GNDA.n299 239.004
R2631 GNDA.n197 GNDA.n121 238.4
R2632 GNDA.n2354 GNDA.n103 238.4
R2633 GNDA.t32 GNDA.t259 236.923
R2634 GNDA.t46 GNDA.t218 236.923
R2635 GNDA.t339 GNDA.t208 236.923
R2636 GNDA.t50 GNDA.t214 236.923
R2637 GNDA.t170 GNDA.t206 236.923
R2638 GNDA.t302 GNDA.t212 236.923
R2639 GNDA.t290 GNDA.t202 236.923
R2640 GNDA.t173 GNDA.t216 236.923
R2641 GNDA.t12 GNDA.t204 236.923
R2642 GNDA.t210 GNDA.t73 236.923
R2643 GNDA.t181 GNDA.t200 236.923
R2644 GNDA.t59 GNDA.t256 236.923
R2645 GNDA.n2410 GNDA.n2409 233.601
R2646 GNDA.n2339 GNDA.n105 227.587
R2647 GNDA.n47 GNDA.n45 227.096
R2648 GNDA.n44 GNDA.n42 227.096
R2649 GNDA.n47 GNDA.n46 226.534
R2650 GNDA.n44 GNDA.n43 226.534
R2651 GNDA.n2306 GNDA.n237 224.553
R2652 GNDA.n136 GNDA.t306 224.525
R2653 GNDA.n138 GNDA.t230 224.525
R2654 GNDA.n85 GNDA.t280 224.525
R2655 GNDA.n83 GNDA.t270 224.525
R2656 GNDA.n50 GNDA.n49 222.034
R2657 GNDA.n1287 GNDA.n1286 221.667
R2658 GNDA.n1125 GNDA.n1124 221.667
R2659 GNDA.n953 GNDA.n875 221.667
R2660 GNDA.n1639 GNDA.n1638 221.667
R2661 GNDA.n418 GNDA.n370 221.667
R2662 GNDA.n1825 GNDA.n1824 221.667
R2663 GNDA.n655 GNDA.n654 221.667
R2664 GNDA.n2049 GNDA.n2048 221.667
R2665 GNDA.n810 GNDA.n809 221.667
R2666 GNDA.n2422 GNDA.n25 217.601
R2667 GNDA.t296 GNDA.n2386 214.944
R2668 GNDA.n142 GNDA.t312 214.944
R2669 GNDA.n2406 GNDA.n25 214.4
R2670 GNDA.n54 GNDA.n53 211.201
R2671 GNDA.n55 GNDA.n54 211.201
R2672 GNDA.n131 GNDA.n130 211.201
R2673 GNDA.n130 GNDA.n126 211.201
R2674 GNDA.n2363 GNDA.n98 211.201
R2675 GNDA.n2364 GNDA.n2363 211.201
R2676 GNDA.n14 GNDA.n12 206.052
R2677 GNDA.n3 GNDA.n1 206.052
R2678 GNDA.n22 GNDA.n21 205.488
R2679 GNDA.n20 GNDA.n19 205.488
R2680 GNDA.n18 GNDA.n17 205.488
R2681 GNDA.n16 GNDA.n15 205.488
R2682 GNDA.n14 GNDA.n13 205.488
R2683 GNDA.n11 GNDA.n10 205.488
R2684 GNDA.n9 GNDA.n8 205.488
R2685 GNDA.n7 GNDA.n6 205.488
R2686 GNDA.n5 GNDA.n4 205.488
R2687 GNDA.n3 GNDA.n2 205.488
R2688 GNDA.n2406 GNDA.n24 203.201
R2689 GNDA.n2423 GNDA.n2422 201.601
R2690 GNDA.n2122 GNDA.n2121 197
R2691 GNDA.n2125 GNDA.n2122 197
R2692 GNDA.n2101 GNDA.n498 197
R2693 GNDA.n285 GNDA.n270 197
R2694 GNDA.n2209 GNDA.n2208 197
R2695 GNDA.n286 GNDA.n276 197
R2696 GNDA.n1038 GNDA.n497 197
R2697 GNDA.n1665 GNDA.n496 197
R2698 GNDA.n1072 GNDA.n454 197
R2699 GNDA.n2248 GNDA.n264 197
R2700 GNDA.n2206 GNDA.n455 197
R2701 GNDA.n190 GNDA.n121 195
R2702 GNDA.n191 GNDA.n190 195
R2703 GNDA.n120 GNDA.n119 195
R2704 GNDA.n119 GNDA.n118 195
R2705 GNDA.n2345 GNDA.n104 195
R2706 GNDA.n2346 GNDA.n2345 195
R2707 GNDA.n2342 GNDA.n103 195
R2708 GNDA.n2342 GNDA.n2341 195
R2709 GNDA.n141 GNDA.n140 192
R2710 GNDA.n2367 GNDA.n84 192
R2711 GNDA.n2104 GNDA.n477 187.249
R2712 GNDA.n2246 GNDA.n278 187.249
R2713 GNDA.n1720 GNDA.n1719 187.249
R2714 GNDA.n288 GNDA.n277 187.249
R2715 GNDA.n1376 GNDA.n1193 187.249
R2716 GNDA.n1691 GNDA.n1690 187.249
R2717 GNDA.n1922 GNDA.n1921 187.249
R2718 GNDA.n2269 GNDA.n281 187.249
R2719 GNDA.n2171 GNDA.n2170 187.249
R2720 GNDA.n1772 GNDA.n308 186.451
R2721 GNDA.n2405 GNDA.t212 186.155
R2722 GNDA.n2405 GNDA.t202 186.155
R2723 GNDA.n1253 GNDA.n1252 185
R2724 GNDA.n1254 GNDA.n1251 185
R2725 GNDA.n1254 GNDA.t244 185
R2726 GNDA.n1257 GNDA.n1256 185
R2727 GNDA.n1258 GNDA.n1250 185
R2728 GNDA.n1260 GNDA.n1259 185
R2729 GNDA.n1262 GNDA.n1249 185
R2730 GNDA.n1265 GNDA.n1264 185
R2731 GNDA.n1266 GNDA.n1248 185
R2732 GNDA.n1268 GNDA.n1267 185
R2733 GNDA.n1270 GNDA.n1247 185
R2734 GNDA.n1273 GNDA.n1272 185
R2735 GNDA.n1274 GNDA.n1246 185
R2736 GNDA.n1276 GNDA.n1275 185
R2737 GNDA.n1278 GNDA.n1245 185
R2738 GNDA.n1281 GNDA.n1280 185
R2739 GNDA.n1282 GNDA.n1244 185
R2740 GNDA.n1284 GNDA.n1283 185
R2741 GNDA.n1286 GNDA.n1243 185
R2742 GNDA.n1303 GNDA.n1238 185
R2743 GNDA.n1301 GNDA.n1300 185
R2744 GNDA.n1299 GNDA.n1239 185
R2745 GNDA.n1298 GNDA.n1297 185
R2746 GNDA.n1295 GNDA.n1240 185
R2747 GNDA.n1293 GNDA.n1292 185
R2748 GNDA.n1291 GNDA.n1241 185
R2749 GNDA.n1241 GNDA.t244 185
R2750 GNDA.n1290 GNDA.n1289 185
R2751 GNDA.n1287 GNDA.n1242 185
R2752 GNDA.n1091 GNDA.n1090 185
R2753 GNDA.n1092 GNDA.n1089 185
R2754 GNDA.n1092 GNDA.t223 185
R2755 GNDA.n1095 GNDA.n1094 185
R2756 GNDA.n1096 GNDA.n1088 185
R2757 GNDA.n1098 GNDA.n1097 185
R2758 GNDA.n1100 GNDA.n1087 185
R2759 GNDA.n1103 GNDA.n1102 185
R2760 GNDA.n1104 GNDA.n1086 185
R2761 GNDA.n1106 GNDA.n1105 185
R2762 GNDA.n1108 GNDA.n1085 185
R2763 GNDA.n1111 GNDA.n1110 185
R2764 GNDA.n1112 GNDA.n1084 185
R2765 GNDA.n1114 GNDA.n1113 185
R2766 GNDA.n1116 GNDA.n1083 185
R2767 GNDA.n1119 GNDA.n1118 185
R2768 GNDA.n1120 GNDA.n1082 185
R2769 GNDA.n1122 GNDA.n1121 185
R2770 GNDA.n1124 GNDA.n1081 185
R2771 GNDA.n1141 GNDA.n1076 185
R2772 GNDA.n1139 GNDA.n1138 185
R2773 GNDA.n1137 GNDA.n1077 185
R2774 GNDA.n1136 GNDA.n1135 185
R2775 GNDA.n1133 GNDA.n1078 185
R2776 GNDA.n1131 GNDA.n1130 185
R2777 GNDA.n1129 GNDA.n1079 185
R2778 GNDA.n1079 GNDA.t223 185
R2779 GNDA.n1128 GNDA.n1127 185
R2780 GNDA.n1125 GNDA.n1080 185
R2781 GNDA.n918 GNDA.n917 185
R2782 GNDA.n919 GNDA.n883 185
R2783 GNDA.n883 GNDA.t310 185
R2784 GNDA.n921 GNDA.n920 185
R2785 GNDA.n923 GNDA.n882 185
R2786 GNDA.n926 GNDA.n925 185
R2787 GNDA.n927 GNDA.n881 185
R2788 GNDA.n929 GNDA.n928 185
R2789 GNDA.n931 GNDA.n880 185
R2790 GNDA.n934 GNDA.n933 185
R2791 GNDA.n935 GNDA.n879 185
R2792 GNDA.n937 GNDA.n936 185
R2793 GNDA.n939 GNDA.n878 185
R2794 GNDA.n942 GNDA.n941 185
R2795 GNDA.n943 GNDA.n877 185
R2796 GNDA.n945 GNDA.n944 185
R2797 GNDA.n947 GNDA.n876 185
R2798 GNDA.n950 GNDA.n949 185
R2799 GNDA.n951 GNDA.n875 185
R2800 GNDA.n968 GNDA.n967 185
R2801 GNDA.n965 GNDA.n869 185
R2802 GNDA.n964 GNDA.n871 185
R2803 GNDA.n962 GNDA.n961 185
R2804 GNDA.n960 GNDA.n872 185
R2805 GNDA.n959 GNDA.n958 185
R2806 GNDA.n956 GNDA.n873 185
R2807 GNDA.n956 GNDA.t310 185
R2808 GNDA.n955 GNDA.n874 185
R2809 GNDA.n953 GNDA.n952 185
R2810 GNDA.n1605 GNDA.n1507 185
R2811 GNDA.n1606 GNDA.n1506 185
R2812 GNDA.n1606 GNDA.t248 185
R2813 GNDA.n1609 GNDA.n1608 185
R2814 GNDA.n1610 GNDA.n1505 185
R2815 GNDA.n1612 GNDA.n1611 185
R2816 GNDA.n1614 GNDA.n1504 185
R2817 GNDA.n1617 GNDA.n1616 185
R2818 GNDA.n1618 GNDA.n1503 185
R2819 GNDA.n1620 GNDA.n1619 185
R2820 GNDA.n1622 GNDA.n1502 185
R2821 GNDA.n1625 GNDA.n1624 185
R2822 GNDA.n1626 GNDA.n1501 185
R2823 GNDA.n1628 GNDA.n1627 185
R2824 GNDA.n1630 GNDA.n1500 185
R2825 GNDA.n1633 GNDA.n1632 185
R2826 GNDA.n1634 GNDA.n1499 185
R2827 GNDA.n1636 GNDA.n1635 185
R2828 GNDA.n1638 GNDA.n1498 185
R2829 GNDA.n1655 GNDA.n1493 185
R2830 GNDA.n1653 GNDA.n1652 185
R2831 GNDA.n1651 GNDA.n1494 185
R2832 GNDA.n1650 GNDA.n1649 185
R2833 GNDA.n1647 GNDA.n1495 185
R2834 GNDA.n1645 GNDA.n1644 185
R2835 GNDA.n1643 GNDA.n1496 185
R2836 GNDA.n1496 GNDA.t248 185
R2837 GNDA.n1642 GNDA.n1641 185
R2838 GNDA.n1639 GNDA.n1497 185
R2839 GNDA.n383 GNDA.n382 185
R2840 GNDA.n384 GNDA.n378 185
R2841 GNDA.n378 GNDA.t250 185
R2842 GNDA.n386 GNDA.n385 185
R2843 GNDA.n388 GNDA.n377 185
R2844 GNDA.n391 GNDA.n390 185
R2845 GNDA.n392 GNDA.n376 185
R2846 GNDA.n394 GNDA.n393 185
R2847 GNDA.n396 GNDA.n375 185
R2848 GNDA.n399 GNDA.n398 185
R2849 GNDA.n400 GNDA.n374 185
R2850 GNDA.n402 GNDA.n401 185
R2851 GNDA.n404 GNDA.n373 185
R2852 GNDA.n407 GNDA.n406 185
R2853 GNDA.n408 GNDA.n372 185
R2854 GNDA.n410 GNDA.n409 185
R2855 GNDA.n412 GNDA.n371 185
R2856 GNDA.n415 GNDA.n414 185
R2857 GNDA.n416 GNDA.n370 185
R2858 GNDA.n433 GNDA.n432 185
R2859 GNDA.n430 GNDA.n363 185
R2860 GNDA.n429 GNDA.n366 185
R2861 GNDA.n427 GNDA.n426 185
R2862 GNDA.n425 GNDA.n367 185
R2863 GNDA.n424 GNDA.n423 185
R2864 GNDA.n421 GNDA.n368 185
R2865 GNDA.n421 GNDA.t250 185
R2866 GNDA.n420 GNDA.n369 185
R2867 GNDA.n418 GNDA.n417 185
R2868 GNDA.n1791 GNDA.n1018 185
R2869 GNDA.n1792 GNDA.n1017 185
R2870 GNDA.n1792 GNDA.t234 185
R2871 GNDA.n1795 GNDA.n1794 185
R2872 GNDA.n1796 GNDA.n1016 185
R2873 GNDA.n1798 GNDA.n1797 185
R2874 GNDA.n1800 GNDA.n1015 185
R2875 GNDA.n1803 GNDA.n1802 185
R2876 GNDA.n1804 GNDA.n1014 185
R2877 GNDA.n1806 GNDA.n1805 185
R2878 GNDA.n1808 GNDA.n1013 185
R2879 GNDA.n1811 GNDA.n1810 185
R2880 GNDA.n1812 GNDA.n1012 185
R2881 GNDA.n1814 GNDA.n1813 185
R2882 GNDA.n1816 GNDA.n1011 185
R2883 GNDA.n1819 GNDA.n1818 185
R2884 GNDA.n1820 GNDA.n1010 185
R2885 GNDA.n1822 GNDA.n1821 185
R2886 GNDA.n1824 GNDA.n1009 185
R2887 GNDA.n1841 GNDA.n1004 185
R2888 GNDA.n1839 GNDA.n1838 185
R2889 GNDA.n1837 GNDA.n1005 185
R2890 GNDA.n1836 GNDA.n1835 185
R2891 GNDA.n1833 GNDA.n1006 185
R2892 GNDA.n1831 GNDA.n1830 185
R2893 GNDA.n1829 GNDA.n1007 185
R2894 GNDA.n1007 GNDA.t234 185
R2895 GNDA.n1828 GNDA.n1827 185
R2896 GNDA.n1825 GNDA.n1008 185
R2897 GNDA.n1843 GNDA.n1842 185
R2898 GNDA.n1768 GNDA.n1001 185
R2899 GNDA.n1770 GNDA.n1769 185
R2900 GNDA.n1765 GNDA.n1764 185
R2901 GNDA.n1777 GNDA.n1776 185
R2902 GNDA.n1780 GNDA.n1779 185
R2903 GNDA.n1763 GNDA.n1760 185
R2904 GNDA.n1021 GNDA.n1019 185
R2905 GNDA.n1789 GNDA.n1788 185
R2906 GNDA.n365 GNDA.n362 185
R2907 GNDA.n355 GNDA.n353 185
R2908 GNDA.n2221 GNDA.n2220 185
R2909 GNDA.n2223 GNDA.n352 185
R2910 GNDA.n2225 GNDA.n2224 185
R2911 GNDA.n348 GNDA.n347 185
R2912 GNDA.n2232 GNDA.n2231 185
R2913 GNDA.n2235 GNDA.n2234 185
R2914 GNDA.n346 GNDA.n344 185
R2915 GNDA.n1657 GNDA.n1656 185
R2916 GNDA.n1582 GNDA.n1489 185
R2917 GNDA.n1584 GNDA.n1583 185
R2918 GNDA.n1579 GNDA.n1578 185
R2919 GNDA.n1591 GNDA.n1590 185
R2920 GNDA.n1594 GNDA.n1593 185
R2921 GNDA.n1577 GNDA.n1574 185
R2922 GNDA.n1510 GNDA.n1508 185
R2923 GNDA.n1603 GNDA.n1602 185
R2924 GNDA.n870 GNDA.n868 185
R2925 GNDA.n897 GNDA.n895 185
R2926 GNDA.n899 GNDA.n898 185
R2927 GNDA.n901 GNDA.n890 185
R2928 GNDA.n906 GNDA.n905 185
R2929 GNDA.n908 GNDA.n889 185
R2930 GNDA.n910 GNDA.n909 185
R2931 GNDA.n912 GNDA.n885 185
R2932 GNDA.n915 GNDA.n914 185
R2933 GNDA.n1143 GNDA.n1142 185
R2934 GNDA.n1064 GNDA.n1062 185
R2935 GNDA.n1150 GNDA.n1149 185
R2936 GNDA.n1152 GNDA.n1061 185
R2937 GNDA.n1154 GNDA.n1153 185
R2938 GNDA.n1055 GNDA.n1053 185
R2939 GNDA.n1161 GNDA.n1160 185
R2940 GNDA.n1163 GNDA.n1052 185
R2941 GNDA.n1165 GNDA.n1164 185
R2942 GNDA.n1305 GNDA.n1304 185
R2943 GNDA.n1225 GNDA.n1223 185
R2944 GNDA.n1312 GNDA.n1311 185
R2945 GNDA.n1314 GNDA.n1222 185
R2946 GNDA.n1316 GNDA.n1315 185
R2947 GNDA.n1216 GNDA.n1214 185
R2948 GNDA.n1323 GNDA.n1322 185
R2949 GNDA.n1325 GNDA.n1213 185
R2950 GNDA.n1327 GNDA.n1326 185
R2951 GNDA.n621 GNDA.n517 185
R2952 GNDA.n622 GNDA.n516 185
R2953 GNDA.n622 GNDA.t264 185
R2954 GNDA.n625 GNDA.n624 185
R2955 GNDA.n626 GNDA.n515 185
R2956 GNDA.n628 GNDA.n627 185
R2957 GNDA.n630 GNDA.n514 185
R2958 GNDA.n633 GNDA.n632 185
R2959 GNDA.n634 GNDA.n513 185
R2960 GNDA.n636 GNDA.n635 185
R2961 GNDA.n638 GNDA.n512 185
R2962 GNDA.n641 GNDA.n640 185
R2963 GNDA.n642 GNDA.n511 185
R2964 GNDA.n644 GNDA.n643 185
R2965 GNDA.n646 GNDA.n510 185
R2966 GNDA.n649 GNDA.n648 185
R2967 GNDA.n650 GNDA.n509 185
R2968 GNDA.n652 GNDA.n651 185
R2969 GNDA.n654 GNDA.n508 185
R2970 GNDA.n671 GNDA.n503 185
R2971 GNDA.n669 GNDA.n668 185
R2972 GNDA.n667 GNDA.n504 185
R2973 GNDA.n666 GNDA.n665 185
R2974 GNDA.n663 GNDA.n505 185
R2975 GNDA.n661 GNDA.n660 185
R2976 GNDA.n659 GNDA.n506 185
R2977 GNDA.n506 GNDA.t264 185
R2978 GNDA.n658 GNDA.n657 185
R2979 GNDA.n655 GNDA.n507 185
R2980 GNDA.n2015 GNDA.n2014 185
R2981 GNDA.n2016 GNDA.n2013 185
R2982 GNDA.n2016 GNDA.t277 185
R2983 GNDA.n2019 GNDA.n2018 185
R2984 GNDA.n2020 GNDA.n2012 185
R2985 GNDA.n2022 GNDA.n2021 185
R2986 GNDA.n2024 GNDA.n2011 185
R2987 GNDA.n2027 GNDA.n2026 185
R2988 GNDA.n2028 GNDA.n2010 185
R2989 GNDA.n2030 GNDA.n2029 185
R2990 GNDA.n2032 GNDA.n2009 185
R2991 GNDA.n2035 GNDA.n2034 185
R2992 GNDA.n2036 GNDA.n2008 185
R2993 GNDA.n2038 GNDA.n2037 185
R2994 GNDA.n2040 GNDA.n2007 185
R2995 GNDA.n2043 GNDA.n2042 185
R2996 GNDA.n2044 GNDA.n2006 185
R2997 GNDA.n2046 GNDA.n2045 185
R2998 GNDA.n2048 GNDA.n2005 185
R2999 GNDA.n2065 GNDA.n2000 185
R3000 GNDA.n2063 GNDA.n2062 185
R3001 GNDA.n2061 GNDA.n2001 185
R3002 GNDA.n2060 GNDA.n2059 185
R3003 GNDA.n2057 GNDA.n2002 185
R3004 GNDA.n2055 GNDA.n2054 185
R3005 GNDA.n2053 GNDA.n2003 185
R3006 GNDA.n2003 GNDA.t277 185
R3007 GNDA.n2052 GNDA.n2051 185
R3008 GNDA.n2049 GNDA.n2004 185
R3009 GNDA.n776 GNDA.n744 185
R3010 GNDA.n777 GNDA.n743 185
R3011 GNDA.n777 GNDA.t249 185
R3012 GNDA.n780 GNDA.n779 185
R3013 GNDA.n781 GNDA.n742 185
R3014 GNDA.n783 GNDA.n782 185
R3015 GNDA.n785 GNDA.n741 185
R3016 GNDA.n788 GNDA.n787 185
R3017 GNDA.n789 GNDA.n740 185
R3018 GNDA.n791 GNDA.n790 185
R3019 GNDA.n793 GNDA.n739 185
R3020 GNDA.n796 GNDA.n795 185
R3021 GNDA.n797 GNDA.n738 185
R3022 GNDA.n799 GNDA.n798 185
R3023 GNDA.n801 GNDA.n737 185
R3024 GNDA.n804 GNDA.n803 185
R3025 GNDA.n805 GNDA.n736 185
R3026 GNDA.n807 GNDA.n806 185
R3027 GNDA.n809 GNDA.n735 185
R3028 GNDA.n826 GNDA.n730 185
R3029 GNDA.n824 GNDA.n823 185
R3030 GNDA.n822 GNDA.n731 185
R3031 GNDA.n821 GNDA.n820 185
R3032 GNDA.n818 GNDA.n732 185
R3033 GNDA.n816 GNDA.n815 185
R3034 GNDA.n814 GNDA.n733 185
R3035 GNDA.n733 GNDA.t249 185
R3036 GNDA.n813 GNDA.n812 185
R3037 GNDA.n810 GNDA.n734 185
R3038 GNDA.n828 GNDA.n827 185
R3039 GNDA.n756 GNDA.n726 185
R3040 GNDA.n758 GNDA.n757 185
R3041 GNDA.n760 GNDA.n752 185
R3042 GNDA.n765 GNDA.n764 185
R3043 GNDA.n767 GNDA.n751 185
R3044 GNDA.n769 GNDA.n768 185
R3045 GNDA.n771 GNDA.n745 185
R3046 GNDA.n774 GNDA.n773 185
R3047 GNDA.n2067 GNDA.n2066 185
R3048 GNDA.n1990 GNDA.n1988 185
R3049 GNDA.n2074 GNDA.n2073 185
R3050 GNDA.n2076 GNDA.n1987 185
R3051 GNDA.n2078 GNDA.n2077 185
R3052 GNDA.n1981 GNDA.n1979 185
R3053 GNDA.n2085 GNDA.n2084 185
R3054 GNDA.n2087 GNDA.n1978 185
R3055 GNDA.n2089 GNDA.n2088 185
R3056 GNDA.n673 GNDA.n672 185
R3057 GNDA.n599 GNDA.n598 185
R3058 GNDA.n601 GNDA.n600 185
R3059 GNDA.n591 GNDA.n589 185
R3060 GNDA.n608 GNDA.n607 185
R3061 GNDA.n610 GNDA.n588 185
R3062 GNDA.n612 GNDA.n611 185
R3063 GNDA.n520 GNDA.n518 185
R3064 GNDA.n619 GNDA.n618 185
R3065 GNDA.n132 GNDA.n131 182.4
R3066 GNDA.n2366 GNDA.n2364 182.4
R3067 GNDA.n2322 GNDA.n222 179.917
R3068 GNDA.n186 GNDA.n126 176
R3069 GNDA.n1477 GNDA.n1409 176
R3070 GNDA.n1477 GNDA.n1476 176
R3071 GNDA.n2370 GNDA.n98 176
R3072 GNDA.n616 GNDA.n584 175.546
R3073 GNDA.n614 GNDA.n585 175.546
R3074 GNDA.n605 GNDA.n593 175.546
R3075 GNDA.n603 GNDA.n595 175.546
R3076 GNDA.n675 GNDA.n500 175.546
R3077 GNDA.n554 GNDA.n552 175.546
R3078 GNDA.n552 GNDA.n551 175.546
R3079 GNDA.n548 GNDA.n547 175.546
R3080 GNDA.n545 GNDA.n531 175.546
R3081 GNDA.n541 GNDA.n539 175.546
R3082 GNDA.n537 GNDA.n534 175.546
R3083 GNDA.n562 GNDA.n560 175.546
R3084 GNDA.n566 GNDA.n525 175.546
R3085 GNDA.n570 GNDA.n568 175.546
R3086 GNDA.n574 GNDA.n523 175.546
R3087 GNDA.n577 GNDA.n576 175.546
R3088 GNDA.n1950 GNDA.n478 175.546
R3089 GNDA.n1956 GNDA.n1955 175.546
R3090 GNDA.n1962 GNDA.n1961 175.546
R3091 GNDA.n1968 GNDA.n1967 175.546
R3092 GNDA.n1970 GNDA.n479 175.546
R3093 GNDA.n2091 GNDA.n1975 175.546
R3094 GNDA.n2082 GNDA.n1983 175.546
R3095 GNDA.n2080 GNDA.n1984 175.546
R3096 GNDA.n2071 GNDA.n1992 175.546
R3097 GNDA.n2069 GNDA.n1993 175.546
R3098 GNDA.n1897 GNDA.n711 175.546
R3099 GNDA.n858 GNDA.n711 175.546
R3100 GNDA.n859 GNDA.n858 175.546
R3101 GNDA.n860 GNDA.n859 175.546
R3102 GNDA.n902 GNDA.n860 175.546
R3103 GNDA.n903 GNDA.n902 175.546
R3104 GNDA.n903 GNDA.n864 175.546
R3105 GNDA.n865 GNDA.n864 175.546
R3106 GNDA.n866 GNDA.n865 175.546
R3107 GNDA.n994 GNDA.n866 175.546
R3108 GNDA.n994 GNDA.n867 175.546
R3109 GNDA.n971 GNDA.n278 175.546
R3110 GNDA.n975 GNDA.n974 175.546
R3111 GNDA.n979 GNDA.n978 175.546
R3112 GNDA.n983 GNDA.n982 175.546
R3113 GNDA.n987 GNDA.n986 175.546
R3114 GNDA.n851 GNDA.n714 175.546
R3115 GNDA.n847 GNDA.n714 175.546
R3116 GNDA.n847 GNDA.n716 175.546
R3117 GNDA.n843 GNDA.n716 175.546
R3118 GNDA.n843 GNDA.n720 175.546
R3119 GNDA.n839 GNDA.n720 175.546
R3120 GNDA.n839 GNDA.n838 175.546
R3121 GNDA.n838 GNDA.n722 175.546
R3122 GNDA.n834 GNDA.n722 175.546
R3123 GNDA.n834 GNDA.n290 175.546
R3124 GNDA.n2245 GNDA.n290 175.546
R3125 GNDA.n693 GNDA.n692 175.546
R3126 GNDA.n696 GNDA.n695 175.546
R3127 GNDA.n699 GNDA.n698 175.546
R3128 GNDA.n702 GNDA.n701 175.546
R3129 GNDA.n705 GNDA.n704 175.546
R3130 GNDA.n1698 GNDA.n1033 175.546
R3131 GNDA.n1702 GNDA.n1033 175.546
R3132 GNDA.n1706 GNDA.n1704 175.546
R3133 GNDA.n1710 GNDA.n1031 175.546
R3134 GNDA.n1714 GNDA.n1712 175.546
R3135 GNDA.n1718 GNDA.n1029 175.546
R3136 GNDA.n1378 GNDA.n332 175.546
R3137 GNDA.n1380 GNDA.n1379 175.546
R3138 GNDA.n1382 GNDA.n1381 175.546
R3139 GNDA.n1384 GNDA.n1383 175.546
R3140 GNDA.n1386 GNDA.n1385 175.546
R3141 GNDA.n1726 GNDA.n1725 175.546
R3142 GNDA.n1729 GNDA.n1728 175.546
R3143 GNDA.n1737 GNDA.n1736 175.546
R3144 GNDA.n1744 GNDA.n1743 175.546
R3145 GNDA.n1746 GNDA.n442 175.546
R3146 GNDA.n2241 GNDA.n339 175.546
R3147 GNDA.n2237 GNDA.n339 175.546
R3148 GNDA.n2237 GNDA.n343 175.546
R3149 GNDA.n2229 GNDA.n343 175.546
R3150 GNDA.n2229 GNDA.n2227 175.546
R3151 GNDA.n2227 GNDA.n349 175.546
R3152 GNDA.n356 GNDA.n349 175.546
R3153 GNDA.n2218 GNDA.n356 175.546
R3154 GNDA.n2218 GNDA.n357 175.546
R3155 GNDA.n2214 GNDA.n357 175.546
R3156 GNDA.n2214 GNDA.n360 175.546
R3157 GNDA.n1895 GNDA.n855 175.546
R3158 GNDA.n1891 GNDA.n855 175.546
R3159 GNDA.n1891 GNDA.n857 175.546
R3160 GNDA.n1887 GNDA.n857 175.546
R3161 GNDA.n1887 GNDA.n861 175.546
R3162 GNDA.n1883 GNDA.n861 175.546
R3163 GNDA.n1883 GNDA.n1882 175.546
R3164 GNDA.n1882 GNDA.n863 175.546
R3165 GNDA.n1878 GNDA.n863 175.546
R3166 GNDA.n1878 GNDA.n996 175.546
R3167 GNDA.n1874 GNDA.n996 175.546
R3168 GNDA.n1723 GNDA.n854 175.546
R3169 GNDA.n1731 GNDA.n1027 175.546
R3170 GNDA.n1734 GNDA.n1733 175.546
R3171 GNDA.n1741 GNDA.n1739 175.546
R3172 GNDA.n1748 GNDA.n1024 175.546
R3173 GNDA.n1870 GNDA.n277 175.546
R3174 GNDA.n1868 GNDA.n1867 175.546
R3175 GNDA.n1864 GNDA.n1863 175.546
R3176 GNDA.n1860 GNDA.n1859 175.546
R3177 GNDA.n1856 GNDA.n1855 175.546
R3178 GNDA.n1755 GNDA.n1754 175.546
R3179 GNDA.n1786 GNDA.n1755 175.546
R3180 GNDA.n1786 GNDA.n1756 175.546
R3181 GNDA.n1782 GNDA.n1756 175.546
R3182 GNDA.n1782 GNDA.n1758 175.546
R3183 GNDA.n1774 GNDA.n1758 175.546
R3184 GNDA.n1774 GNDA.n1773 175.546
R3185 GNDA.n1773 GNDA.n1000 175.546
R3186 GNDA.n1845 GNDA.n999 175.546
R3187 GNDA.n1329 GNDA.n1210 175.546
R3188 GNDA.n1320 GNDA.n1218 175.546
R3189 GNDA.n1318 GNDA.n1219 175.546
R3190 GNDA.n1309 GNDA.n1227 175.546
R3191 GNDA.n1307 GNDA.n1228 175.546
R3192 GNDA.n1349 GNDA.n1200 175.546
R3193 GNDA.n1345 GNDA.n1344 175.546
R3194 GNDA.n1342 GNDA.n1203 175.546
R3195 GNDA.n1338 GNDA.n1337 175.546
R3196 GNDA.n1335 GNDA.n1206 175.546
R3197 GNDA.n1190 GNDA.n1189 175.546
R3198 GNDA.n1186 GNDA.n1185 175.546
R3199 GNDA.n1182 GNDA.n1181 175.546
R3200 GNDA.n1178 GNDA.n1177 175.546
R3201 GNDA.n1174 GNDA.n484 175.546
R3202 GNDA.n1357 GNDA.n1198 175.546
R3203 GNDA.n1361 GNDA.n1359 175.546
R3204 GNDA.n1365 GNDA.n1196 175.546
R3205 GNDA.n1369 GNDA.n1367 175.546
R3206 GNDA.n1373 GNDA.n1194 175.546
R3207 GNDA.n1600 GNDA.n1511 175.546
R3208 GNDA.n1600 GNDA.n1512 175.546
R3209 GNDA.n1596 GNDA.n1512 175.546
R3210 GNDA.n1596 GNDA.n1572 175.546
R3211 GNDA.n1588 GNDA.n1572 175.546
R3212 GNDA.n1588 GNDA.n1587 175.546
R3213 GNDA.n1587 GNDA.n1488 175.546
R3214 GNDA.n1659 GNDA.n1488 175.546
R3215 GNDA.n1659 GNDA.n1388 175.546
R3216 GNDA.n1664 GNDA.n1388 175.546
R3217 GNDA.n1550 GNDA.n1548 175.546
R3218 GNDA.n1554 GNDA.n1517 175.546
R3219 GNDA.n1558 GNDA.n1556 175.546
R3220 GNDA.n1562 GNDA.n1515 175.546
R3221 GNDA.n1565 GNDA.n1564 175.546
R3222 GNDA.n1687 GNDA.n1686 175.546
R3223 GNDA.n1683 GNDA.n1682 175.546
R3224 GNDA.n1679 GNDA.n1678 175.546
R3225 GNDA.n1675 GNDA.n1674 175.546
R3226 GNDA.n1671 GNDA.n490 175.546
R3227 GNDA.n1542 GNDA.n1541 175.546
R3228 GNDA.n1539 GNDA.n1522 175.546
R3229 GNDA.n1535 GNDA.n1534 175.546
R3230 GNDA.n1532 GNDA.n1525 175.546
R3231 GNDA.n1528 GNDA.n1527 175.546
R3232 GNDA.n1167 GNDA.n1049 175.546
R3233 GNDA.n1158 GNDA.n1057 175.546
R3234 GNDA.n1156 GNDA.n1058 175.546
R3235 GNDA.n1147 GNDA.n1066 175.546
R3236 GNDA.n1145 GNDA.n1067 175.546
R3237 GNDA.n1918 GNDA.n1917 175.546
R3238 GNDA.n1914 GNDA.n1913 175.546
R3239 GNDA.n1910 GNDA.n1909 175.546
R3240 GNDA.n1906 GNDA.n1905 175.546
R3241 GNDA.n1902 GNDA.n448 175.546
R3242 GNDA.n1941 GNDA.n684 175.546
R3243 GNDA.n1937 GNDA.n689 175.546
R3244 GNDA.n1935 GNDA.n1934 175.546
R3245 GNDA.n1931 GNDA.n1930 175.546
R3246 GNDA.n1927 GNDA.n1926 175.546
R3247 GNDA.n1040 GNDA.n1039 175.546
R3248 GNDA.n1042 GNDA.n1041 175.546
R3249 GNDA.n1044 GNDA.n1043 175.546
R3250 GNDA.n1046 GNDA.n1045 175.546
R3251 GNDA.n1173 GNDA.n1172 175.546
R3252 GNDA.n747 GNDA.n712 175.546
R3253 GNDA.n747 GNDA.n717 175.546
R3254 GNDA.n718 GNDA.n717 175.546
R3255 GNDA.n719 GNDA.n718 175.546
R3256 GNDA.n761 GNDA.n719 175.546
R3257 GNDA.n762 GNDA.n761 175.546
R3258 GNDA.n762 GNDA.n723 175.546
R3259 GNDA.n724 GNDA.n723 175.546
R3260 GNDA.n830 GNDA.n724 175.546
R3261 GNDA.n830 GNDA.n725 175.546
R3262 GNDA.n725 GNDA.n284 175.546
R3263 GNDA.n280 GNDA.n279 175.546
R3264 GNDA.n2264 GNDA.n279 175.546
R3265 GNDA.n2262 GNDA.n2261 175.546
R3266 GNDA.n2258 GNDA.n2257 175.546
R3267 GNDA.n2254 GNDA.n2253 175.546
R3268 GNDA.n2163 GNDA.n2161 175.546
R3269 GNDA.n2159 GNDA.n2138 175.546
R3270 GNDA.n2155 GNDA.n2153 175.546
R3271 GNDA.n2151 GNDA.n2140 175.546
R3272 GNDA.n2147 GNDA.n2145 175.546
R3273 GNDA.n2177 GNDA.n2175 175.546
R3274 GNDA.n2185 GNDA.n464 175.546
R3275 GNDA.n2189 GNDA.n2187 175.546
R3276 GNDA.n2197 GNDA.n462 175.546
R3277 GNDA.n2201 GNDA.n2199 175.546
R3278 GNDA.n2179 GNDA.n2178 175.546
R3279 GNDA.n2183 GNDA.n2182 175.546
R3280 GNDA.n2191 GNDA.n2190 175.546
R3281 GNDA.n2195 GNDA.n2194 175.546
R3282 GNDA.n458 GNDA.n436 175.546
R3283 GNDA.n2112 GNDA.n473 175.546
R3284 GNDA.n2116 GNDA.n2114 175.546
R3285 GNDA.n2129 GNDA.n471 175.546
R3286 GNDA.n2132 GNDA.n2131 175.546
R3287 GNDA.n2134 GNDA.n468 175.546
R3288 GNDA.n2168 GNDA.n468 175.546
R3289 GNDA.n1949 GNDA.n1948 175.546
R3290 GNDA.n1954 GNDA.n1953 175.546
R3291 GNDA.n1960 GNDA.n1959 175.546
R3292 GNDA.n1966 GNDA.n1965 175.546
R3293 GNDA.n2096 GNDA.n2095 175.546
R3294 GNDA.n1974 GNDA.n306 173.881
R3295 GNDA.t224 GNDA.n307 172.876
R3296 GNDA.t224 GNDA.n319 172.615
R3297 GNDA.n1943 GNDA.n306 171.624
R3298 GNDA.n1425 GNDA.n1424 164.369
R3299 GNDA.n2324 GNDA.n219 164.369
R3300 GNDA.n1304 GNDA.n1303 163.333
R3301 GNDA.n1142 GNDA.n1141 163.333
R3302 GNDA.n967 GNDA.n870 163.333
R3303 GNDA.n1656 GNDA.n1655 163.333
R3304 GNDA.n432 GNDA.n365 163.333
R3305 GNDA.n1842 GNDA.n1841 163.333
R3306 GNDA.n672 GNDA.n671 163.333
R3307 GNDA.n2066 GNDA.n2065 163.333
R3308 GNDA.n827 GNDA.n826 163.333
R3309 GNDA.n1411 GNDA.t285 160.725
R3310 GNDA.n1414 GNDA.t300 160.725
R3311 GNDA.n1410 GNDA.t263 160.725
R3312 GNDA.n1408 GNDA.t247 160.725
R3313 GNDA.n1443 GNDA.t276 160.725
R3314 GNDA.n1438 GNDA.t273 160.725
R3315 GNDA.n73 GNDA.n72 160
R3316 GNDA.n2395 GNDA.n2390 160
R3317 GNDA.n2401 GNDA.n2399 160
R3318 GNDA.n2311 GNDA.t106 157.555
R3319 GNDA.n2312 GNDA.t164 157.555
R3320 GNDA.n2409 GNDA.n35 156.8
R3321 GNDA.n76 GNDA.n75 153.601
R3322 GNDA.n139 GNDA.n137 153.601
R3323 GNDA.n2368 GNDA.n86 153.601
R3324 GNDA.n227 GNDA.t129 153.294
R3325 GNDA.n125 GNDA.t237 152.994
R3326 GNDA.n129 GNDA.t222 152.994
R3327 GNDA.n2362 GNDA.t243 152.994
R3328 GNDA.n97 GNDA.t233 152.994
R3329 GNDA.n969 GNDA.n269 152.643
R3330 GNDA.n1899 GNDA.n710 152.643
R3331 GNDA.n338 GNDA.n337 152.643
R3332 GNDA.n1750 GNDA.n1749 152.643
R3333 GNDA.n1852 GNDA.n275 152.643
R3334 GNDA.n2250 GNDA.n263 152.643
R3335 GNDA.n2124 GNDA.n314 152.596
R3336 GNDA.n2417 GNDA.n2416 150.4
R3337 GNDA.n1326 GNDA.n1325 150
R3338 GNDA.n1323 GNDA.n1214 150
R3339 GNDA.n1315 GNDA.n1314 150
R3340 GNDA.n1312 GNDA.n1223 150
R3341 GNDA.n1289 GNDA.n1241 150
R3342 GNDA.n1293 GNDA.n1241 150
R3343 GNDA.n1297 GNDA.n1295 150
R3344 GNDA.n1301 GNDA.n1239 150
R3345 GNDA.n1272 GNDA.n1270 150
R3346 GNDA.n1276 GNDA.n1246 150
R3347 GNDA.n1280 GNDA.n1278 150
R3348 GNDA.n1284 GNDA.n1244 150
R3349 GNDA.n1268 GNDA.n1248 150
R3350 GNDA.n1264 GNDA.n1262 150
R3351 GNDA.n1260 GNDA.n1250 150
R3352 GNDA.n1256 GNDA.n1254 150
R3353 GNDA.n1254 GNDA.n1253 150
R3354 GNDA.n1164 GNDA.n1163 150
R3355 GNDA.n1161 GNDA.n1053 150
R3356 GNDA.n1153 GNDA.n1152 150
R3357 GNDA.n1150 GNDA.n1062 150
R3358 GNDA.n1127 GNDA.n1079 150
R3359 GNDA.n1131 GNDA.n1079 150
R3360 GNDA.n1135 GNDA.n1133 150
R3361 GNDA.n1139 GNDA.n1077 150
R3362 GNDA.n1110 GNDA.n1108 150
R3363 GNDA.n1114 GNDA.n1084 150
R3364 GNDA.n1118 GNDA.n1116 150
R3365 GNDA.n1122 GNDA.n1082 150
R3366 GNDA.n1106 GNDA.n1086 150
R3367 GNDA.n1102 GNDA.n1100 150
R3368 GNDA.n1098 GNDA.n1088 150
R3369 GNDA.n1094 GNDA.n1092 150
R3370 GNDA.n1092 GNDA.n1091 150
R3371 GNDA.n915 GNDA.n885 150
R3372 GNDA.n909 GNDA.n908 150
R3373 GNDA.n906 GNDA.n890 150
R3374 GNDA.n898 GNDA.n897 150
R3375 GNDA.n956 GNDA.n955 150
R3376 GNDA.n958 GNDA.n956 150
R3377 GNDA.n962 GNDA.n872 150
R3378 GNDA.n965 GNDA.n964 150
R3379 GNDA.n937 GNDA.n879 150
R3380 GNDA.n941 GNDA.n939 150
R3381 GNDA.n945 GNDA.n877 150
R3382 GNDA.n949 GNDA.n947 150
R3383 GNDA.n933 GNDA.n931 150
R3384 GNDA.n929 GNDA.n881 150
R3385 GNDA.n925 GNDA.n923 150
R3386 GNDA.n921 GNDA.n883 150
R3387 GNDA.n917 GNDA.n883 150
R3388 GNDA.n1603 GNDA.n1508 150
R3389 GNDA.n1593 GNDA.n1577 150
R3390 GNDA.n1591 GNDA.n1578 150
R3391 GNDA.n1583 GNDA.n1582 150
R3392 GNDA.n1641 GNDA.n1496 150
R3393 GNDA.n1645 GNDA.n1496 150
R3394 GNDA.n1649 GNDA.n1647 150
R3395 GNDA.n1653 GNDA.n1494 150
R3396 GNDA.n1624 GNDA.n1622 150
R3397 GNDA.n1628 GNDA.n1501 150
R3398 GNDA.n1632 GNDA.n1630 150
R3399 GNDA.n1636 GNDA.n1499 150
R3400 GNDA.n1620 GNDA.n1503 150
R3401 GNDA.n1616 GNDA.n1614 150
R3402 GNDA.n1612 GNDA.n1505 150
R3403 GNDA.n1608 GNDA.n1606 150
R3404 GNDA.n1606 GNDA.n1605 150
R3405 GNDA.n2234 GNDA.n346 150
R3406 GNDA.n2232 GNDA.n347 150
R3407 GNDA.n2224 GNDA.n2223 150
R3408 GNDA.n2221 GNDA.n353 150
R3409 GNDA.n421 GNDA.n420 150
R3410 GNDA.n423 GNDA.n421 150
R3411 GNDA.n427 GNDA.n367 150
R3412 GNDA.n430 GNDA.n429 150
R3413 GNDA.n402 GNDA.n374 150
R3414 GNDA.n406 GNDA.n404 150
R3415 GNDA.n410 GNDA.n372 150
R3416 GNDA.n414 GNDA.n412 150
R3417 GNDA.n398 GNDA.n396 150
R3418 GNDA.n394 GNDA.n376 150
R3419 GNDA.n390 GNDA.n388 150
R3420 GNDA.n386 GNDA.n378 150
R3421 GNDA.n382 GNDA.n378 150
R3422 GNDA.n1789 GNDA.n1019 150
R3423 GNDA.n1779 GNDA.n1763 150
R3424 GNDA.n1777 GNDA.n1764 150
R3425 GNDA.n1769 GNDA.n1768 150
R3426 GNDA.n1827 GNDA.n1007 150
R3427 GNDA.n1831 GNDA.n1007 150
R3428 GNDA.n1835 GNDA.n1833 150
R3429 GNDA.n1839 GNDA.n1005 150
R3430 GNDA.n1810 GNDA.n1808 150
R3431 GNDA.n1814 GNDA.n1012 150
R3432 GNDA.n1818 GNDA.n1816 150
R3433 GNDA.n1822 GNDA.n1010 150
R3434 GNDA.n1806 GNDA.n1014 150
R3435 GNDA.n1802 GNDA.n1800 150
R3436 GNDA.n1798 GNDA.n1016 150
R3437 GNDA.n1794 GNDA.n1792 150
R3438 GNDA.n1792 GNDA.n1791 150
R3439 GNDA.n619 GNDA.n518 150
R3440 GNDA.n611 GNDA.n610 150
R3441 GNDA.n608 GNDA.n589 150
R3442 GNDA.n600 GNDA.n599 150
R3443 GNDA.n657 GNDA.n506 150
R3444 GNDA.n661 GNDA.n506 150
R3445 GNDA.n665 GNDA.n663 150
R3446 GNDA.n669 GNDA.n504 150
R3447 GNDA.n640 GNDA.n638 150
R3448 GNDA.n644 GNDA.n511 150
R3449 GNDA.n648 GNDA.n646 150
R3450 GNDA.n652 GNDA.n509 150
R3451 GNDA.n636 GNDA.n513 150
R3452 GNDA.n632 GNDA.n630 150
R3453 GNDA.n628 GNDA.n515 150
R3454 GNDA.n624 GNDA.n622 150
R3455 GNDA.n622 GNDA.n621 150
R3456 GNDA.n2088 GNDA.n2087 150
R3457 GNDA.n2085 GNDA.n1979 150
R3458 GNDA.n2077 GNDA.n2076 150
R3459 GNDA.n2074 GNDA.n1988 150
R3460 GNDA.n2051 GNDA.n2003 150
R3461 GNDA.n2055 GNDA.n2003 150
R3462 GNDA.n2059 GNDA.n2057 150
R3463 GNDA.n2063 GNDA.n2001 150
R3464 GNDA.n2034 GNDA.n2032 150
R3465 GNDA.n2038 GNDA.n2008 150
R3466 GNDA.n2042 GNDA.n2040 150
R3467 GNDA.n2046 GNDA.n2006 150
R3468 GNDA.n2030 GNDA.n2010 150
R3469 GNDA.n2026 GNDA.n2024 150
R3470 GNDA.n2022 GNDA.n2012 150
R3471 GNDA.n2018 GNDA.n2016 150
R3472 GNDA.n2016 GNDA.n2015 150
R3473 GNDA.n774 GNDA.n745 150
R3474 GNDA.n768 GNDA.n767 150
R3475 GNDA.n765 GNDA.n752 150
R3476 GNDA.n757 GNDA.n756 150
R3477 GNDA.n812 GNDA.n733 150
R3478 GNDA.n816 GNDA.n733 150
R3479 GNDA.n820 GNDA.n818 150
R3480 GNDA.n824 GNDA.n731 150
R3481 GNDA.n795 GNDA.n793 150
R3482 GNDA.n799 GNDA.n738 150
R3483 GNDA.n803 GNDA.n801 150
R3484 GNDA.n807 GNDA.n736 150
R3485 GNDA.n791 GNDA.n740 150
R3486 GNDA.n787 GNDA.n785 150
R3487 GNDA.n783 GNDA.n742 150
R3488 GNDA.n779 GNDA.n777 150
R3489 GNDA.n777 GNDA.n776 150
R3490 GNDA.n2313 GNDA.t81 148.906
R3491 GNDA.n2313 GNDA.t124 148.653
R3492 GNDA.t242 GNDA.n80 147.511
R3493 GNDA.n144 GNDA.t221 147.511
R3494 GNDA.t165 GNDA.t284 145.403
R3495 GNDA.t1 GNDA.t272 145.403
R3496 GNDA.n1447 GNDA.n1445 139.638
R3497 GNDA.t246 GNDA.t331 139.081
R3498 GNDA.t331 GNDA.t152 139.081
R3499 GNDA.t152 GNDA.t140 139.081
R3500 GNDA.t132 GNDA.t69 139.081
R3501 GNDA.t69 GNDA.t146 139.081
R3502 GNDA.t146 GNDA.t262 139.081
R3503 GNDA.n1463 GNDA.n1462 139.077
R3504 GNDA.n1461 GNDA.n1460 139.077
R3505 GNDA.n1459 GNDA.n1458 139.077
R3506 GNDA.n1457 GNDA.n1456 139.077
R3507 GNDA.n1455 GNDA.n1454 139.077
R3508 GNDA.n1453 GNDA.n1452 139.077
R3509 GNDA.n1451 GNDA.n1450 139.077
R3510 GNDA.n1449 GNDA.n1448 139.077
R3511 GNDA.n1447 GNDA.n1446 139.077
R3512 GNDA.t46 GNDA.t259 135.386
R3513 GNDA.t339 GNDA.t218 135.386
R3514 GNDA.t50 GNDA.t208 135.386
R3515 GNDA.t170 GNDA.t214 135.386
R3516 GNDA.t302 GNDA.t206 135.386
R3517 GNDA.t290 GNDA.t216 135.386
R3518 GNDA.t173 GNDA.t204 135.386
R3519 GNDA.t12 GNDA.t210 135.386
R3520 GNDA.t200 GNDA.t73 135.386
R3521 GNDA.t181 GNDA.t256 135.386
R3522 GNDA.n2372 GNDA.n93 134.867
R3523 GNDA.n183 GNDA.n110 134.867
R3524 GNDA.n1480 GNDA.t140 132.76
R3525 GNDA.n2325 GNDA.t132 132.76
R3526 GNDA.n1420 GNDA.t130 126.438
R3527 GNDA.t197 GNDA.n1468 126.438
R3528 GNDA.n677 GNDA.n498 124.832
R3529 GNDA.n1997 GNDA.n455 124.832
R3530 GNDA.n867 GNDA.n285 124.832
R3531 GNDA.n2246 GNDA.n2245 124.832
R3532 GNDA.n1719 GNDA.n1718 124.832
R3533 GNDA.n2209 GNDA.n360 124.832
R3534 GNDA.n1874 GNDA.n288 124.832
R3535 GNDA.n1849 GNDA.n286 124.832
R3536 GNDA.n1235 GNDA.n1038 124.832
R3537 GNDA.n1376 GNDA.n1375 124.832
R3538 GNDA.n1665 GNDA.n1664 124.832
R3539 GNDA.n1692 GNDA.n1691 124.832
R3540 GNDA.n1073 GNDA.n1072 124.832
R3541 GNDA.n1923 GNDA.n1922 124.832
R3542 GNDA.n2248 GNDA.n284 124.832
R3543 GNDA.n2143 GNDA.n281 124.832
R3544 GNDA.t186 GNDA.t182 120.115
R3545 GNDA.t90 GNDA.t37 120.115
R3546 GNDA.n1416 GNDA.n1415 118.4
R3547 GNDA.n1435 GNDA.n1412 118.4
R3548 GNDA.n1436 GNDA.n1409 118.4
R3549 GNDA.n1476 GNDA.n1475 118.4
R3550 GNDA.n1474 GNDA.n1439 118.4
R3551 GNDA.n1466 GNDA.n1444 118.4
R3552 GNDA.n2305 GNDA.n238 115.311
R3553 GNDA.n64 GNDA.t240 113.974
R3554 GNDA.n70 GNDA.t227 113.974
R3555 GNDA.n69 GNDA.t297 113.974
R3556 GNDA.n68 GNDA.t313 113.974
R3557 GNDA.n67 GNDA.t294 113.974
R3558 GNDA.n66 GNDA.t282 113.974
R3559 GNDA.n2391 GNDA.t309 113.974
R3560 GNDA.n2392 GNDA.t291 113.974
R3561 GNDA.n2393 GNDA.t303 113.974
R3562 GNDA.n2394 GNDA.t288 113.974
R3563 GNDA.t224 GNDA.n294 113.624
R3564 GNDA.n1663 GNDA.n1662 113.624
R3565 GNDA.t224 GNDA.n296 113.624
R3566 GNDA.t224 GNDA.n300 113.624
R3567 GNDA.n53 GNDA.n41 108.8
R3568 GNDA.n56 GNDA.n55 108.8
R3569 GNDA.n1421 GNDA.n1420 101.15
R3570 GNDA.t21 GNDA.t167 101.15
R3571 GNDA.t317 GNDA.t128 101.15
R3572 GNDA.n1468 GNDA.n1442 101.15
R3573 GNDA.t224 GNDA.n316 47.6748
R3574 GNDA.n151 GNDA.n150 99.0842
R3575 GNDA.n153 GNDA.n152 99.0842
R3576 GNDA.n155 GNDA.n154 99.0842
R3577 GNDA.n157 GNDA.n156 99.0842
R3578 GNDA.n159 GNDA.n158 99.0842
R3579 GNDA.n161 GNDA.n160 99.0842
R3580 GNDA.n163 GNDA.n162 99.0842
R3581 GNDA.n165 GNDA.n164 99.0842
R3582 GNDA.n167 GNDA.n166 99.0842
R3583 GNDA.n169 GNDA.n168 99.0842
R3584 GNDA.n171 GNDA.n170 99.0842
R3585 GNDA.n173 GNDA.n172 99.0842
R3586 GNDA.n2123 GNDA.n315 97.1951
R3587 GNDA.n2124 GNDA.n2123 97.1951
R3588 GNDA.n1571 GNDA.n1570 96.926
R3589 GNDA.n179 GNDA.n178 95.101
R3590 GNDA.n2381 GNDA.n2378 95.101
R3591 GNDA.t267 GNDA.n149 94.8842
R3592 GNDA.n34 GNDA.t254 94.8842
R3593 GNDA.t130 GNDA.t299 94.8281
R3594 GNDA.t138 GNDA.t10 94.8281
R3595 GNDA.t319 GNDA.t154 94.8281
R3596 GNDA.t275 GNDA.t197 94.8281
R3597 GNDA.n177 GNDA.n176 94.601
R3598 GNDA.n2380 GNDA.n2379 94.601
R3599 GNDA.t55 GNDA.t232 92.7208
R3600 GNDA.t58 GNDA.t346 92.7208
R3601 GNDA.t335 GNDA.t160 92.7208
R3602 GNDA.t74 GNDA.t323 92.7208
R3603 GNDA.t320 GNDA.t296 92.7208
R3604 GNDA.t312 GNDA.t103 92.7208
R3605 GNDA.t22 GNDA.t87 92.7208
R3606 GNDA.t95 GNDA.t45 92.7208
R3607 GNDA.t13 GNDA.t178 92.7208
R3608 GNDA.t174 GNDA.t236 92.7208
R3609 GNDA.t113 GNDA.t269 88.5063
R3610 GNDA.t229 GNDA.t179 88.5063
R3611 GNDA.n188 GNDA.n187 86.4005
R3612 GNDA.n2361 GNDA.n99 86.4005
R3613 GNDA.n2317 GNDA.n2316 85.2845
R3614 GNDA.n226 GNDA.n225 85.2845
R3615 GNDA.t189 GNDA.t184 82.1844
R3616 GNDA.t150 GNDA.t93 82.1844
R3617 GNDA.t318 GNDA.t142 82.1844
R3618 GNDA.t48 GNDA.t47 82.1844
R3619 GNDA.n2273 GNDA.n2272 81.7659
R3620 GNDA.t224 GNDA.n852 80.9821
R3621 GNDA.n1896 GNDA.t224 80.9821
R3622 GNDA.n2273 GNDA.n2271 80.7438
R3623 GNDA.t279 GNDA.t55 80.0771
R3624 GNDA.t53 GNDA.t113 80.0771
R3625 GNDA.n2419 GNDA.t103 80.0771
R3626 GNDA.t179 GNDA.t168 80.0771
R3627 GNDA.t305 GNDA.t174 80.0771
R3628 GNDA.t224 GNDA.n306 76.3879
R3629 GNDA.n584 GNDA.n583 76.3222
R3630 GNDA.n615 GNDA.n614 76.3222
R3631 GNDA.n593 GNDA.n592 76.3222
R3632 GNDA.n604 GNDA.n603 76.3222
R3633 GNDA.n594 GNDA.n500 76.3222
R3634 GNDA.n677 GNDA.n676 76.3222
R3635 GNDA.n553 GNDA.n527 76.3222
R3636 GNDA.n551 GNDA.n529 76.3222
R3637 GNDA.n547 GNDA.n546 76.3222
R3638 GNDA.n540 GNDA.n531 76.3222
R3639 GNDA.n539 GNDA.n538 76.3222
R3640 GNDA.n560 GNDA.n559 76.3222
R3641 GNDA.n561 GNDA.n525 76.3222
R3642 GNDA.n568 GNDA.n567 76.3222
R3643 GNDA.n569 GNDA.n523 76.3222
R3644 GNDA.n576 GNDA.n575 76.3222
R3645 GNDA.n578 GNDA.n521 76.3222
R3646 GNDA.n2104 GNDA.n2103 76.3222
R3647 GNDA.n1950 GNDA.n483 76.3222
R3648 GNDA.n1956 GNDA.n482 76.3222
R3649 GNDA.n1962 GNDA.n481 76.3222
R3650 GNDA.n1968 GNDA.n480 76.3222
R3651 GNDA.n2100 GNDA.n479 76.3222
R3652 GNDA.n2092 GNDA.n2091 76.3222
R3653 GNDA.n1983 GNDA.n1982 76.3222
R3654 GNDA.n2081 GNDA.n2080 76.3222
R3655 GNDA.n1992 GNDA.n1991 76.3222
R3656 GNDA.n2070 GNDA.n2069 76.3222
R3657 GNDA.n1997 GNDA.n1996 76.3222
R3658 GNDA.n971 GNDA.n265 76.3222
R3659 GNDA.n975 GNDA.n266 76.3222
R3660 GNDA.n979 GNDA.n267 76.3222
R3661 GNDA.n983 GNDA.n268 76.3222
R3662 GNDA.n987 GNDA.n269 76.3222
R3663 GNDA.n695 GNDA.n694 76.3222
R3664 GNDA.n698 GNDA.n697 76.3222
R3665 GNDA.n701 GNDA.n700 76.3222
R3666 GNDA.n704 GNDA.n703 76.3222
R3667 GNDA.n1899 GNDA.n1898 76.3222
R3668 GNDA.n1697 GNDA.n1696 76.3222
R3669 GNDA.n1703 GNDA.n1702 76.3222
R3670 GNDA.n1706 GNDA.n1705 76.3222
R3671 GNDA.n1711 GNDA.n1710 76.3222
R3672 GNDA.n1714 GNDA.n1713 76.3222
R3673 GNDA.n1379 GNDA.n333 76.3222
R3674 GNDA.n1381 GNDA.n334 76.3222
R3675 GNDA.n1383 GNDA.n335 76.3222
R3676 GNDA.n1385 GNDA.n336 76.3222
R3677 GNDA.n2242 GNDA.n338 76.3222
R3678 GNDA.n1720 GNDA.n447 76.3222
R3679 GNDA.n1726 GNDA.n446 76.3222
R3680 GNDA.n1728 GNDA.n445 76.3222
R3681 GNDA.n1737 GNDA.n444 76.3222
R3682 GNDA.n1744 GNDA.n443 76.3222
R3683 GNDA.n442 GNDA.n435 76.3222
R3684 GNDA.n1722 GNDA.n1027 76.3222
R3685 GNDA.n1733 GNDA.n1732 76.3222
R3686 GNDA.n1739 GNDA.n1025 76.3222
R3687 GNDA.n1740 GNDA.n1024 76.3222
R3688 GNDA.n1750 GNDA.n1022 76.3222
R3689 GNDA.n1870 GNDA.n271 76.3222
R3690 GNDA.n1867 GNDA.n272 76.3222
R3691 GNDA.n1863 GNDA.n273 76.3222
R3692 GNDA.n1859 GNDA.n274 76.3222
R3693 GNDA.n1855 GNDA.n275 76.3222
R3694 GNDA.n1846 GNDA.n1845 76.3222
R3695 GNDA.n1849 GNDA.n1848 76.3222
R3696 GNDA.n1330 GNDA.n1329 76.3222
R3697 GNDA.n1218 GNDA.n1217 76.3222
R3698 GNDA.n1319 GNDA.n1318 76.3222
R3699 GNDA.n1227 GNDA.n1226 76.3222
R3700 GNDA.n1308 GNDA.n1307 76.3222
R3701 GNDA.n1235 GNDA.n1234 76.3222
R3702 GNDA.n1350 GNDA.n1349 76.3222
R3703 GNDA.n1345 GNDA.n1202 76.3222
R3704 GNDA.n1343 GNDA.n1342 76.3222
R3705 GNDA.n1338 GNDA.n1205 76.3222
R3706 GNDA.n1336 GNDA.n1335 76.3222
R3707 GNDA.n1209 GNDA.n1207 76.3222
R3708 GNDA.n1193 GNDA.n489 76.3222
R3709 GNDA.n1189 GNDA.n488 76.3222
R3710 GNDA.n1185 GNDA.n487 76.3222
R3711 GNDA.n1181 GNDA.n486 76.3222
R3712 GNDA.n1177 GNDA.n485 76.3222
R3713 GNDA.n1231 GNDA.n484 76.3222
R3714 GNDA.n1352 GNDA.n1198 76.3222
R3715 GNDA.n1359 GNDA.n1358 76.3222
R3716 GNDA.n1360 GNDA.n1196 76.3222
R3717 GNDA.n1367 GNDA.n1366 76.3222
R3718 GNDA.n1368 GNDA.n1194 76.3222
R3719 GNDA.n1375 GNDA.n1374 76.3222
R3720 GNDA.n1353 GNDA.n1352 76.3222
R3721 GNDA.n1358 GNDA.n1357 76.3222
R3722 GNDA.n1361 GNDA.n1360 76.3222
R3723 GNDA.n1366 GNDA.n1365 76.3222
R3724 GNDA.n1369 GNDA.n1368 76.3222
R3725 GNDA.n1374 GNDA.n1373 76.3222
R3726 GNDA.n1337 GNDA.n1336 76.3222
R3727 GNDA.n1205 GNDA.n1203 76.3222
R3728 GNDA.n1344 GNDA.n1343 76.3222
R3729 GNDA.n1202 GNDA.n1200 76.3222
R3730 GNDA.n1351 GNDA.n1350 76.3222
R3731 GNDA.n1547 GNDA.n1546 76.3222
R3732 GNDA.n1550 GNDA.n1549 76.3222
R3733 GNDA.n1555 GNDA.n1554 76.3222
R3734 GNDA.n1558 GNDA.n1557 76.3222
R3735 GNDA.n1563 GNDA.n1562 76.3222
R3736 GNDA.n1566 GNDA.n1565 76.3222
R3737 GNDA.n1690 GNDA.n495 76.3222
R3738 GNDA.n1686 GNDA.n494 76.3222
R3739 GNDA.n1682 GNDA.n493 76.3222
R3740 GNDA.n1678 GNDA.n492 76.3222
R3741 GNDA.n1674 GNDA.n491 76.3222
R3742 GNDA.n1667 GNDA.n490 76.3222
R3743 GNDA.n1542 GNDA.n1521 76.3222
R3744 GNDA.n1540 GNDA.n1539 76.3222
R3745 GNDA.n1535 GNDA.n1524 76.3222
R3746 GNDA.n1533 GNDA.n1532 76.3222
R3747 GNDA.n1528 GNDA.n1526 76.3222
R3748 GNDA.n1692 GNDA.n1037 76.3222
R3749 GNDA.n1521 GNDA.n1519 76.3222
R3750 GNDA.n1541 GNDA.n1540 76.3222
R3751 GNDA.n1524 GNDA.n1522 76.3222
R3752 GNDA.n1534 GNDA.n1533 76.3222
R3753 GNDA.n1526 GNDA.n1525 76.3222
R3754 GNDA.n1527 GNDA.n1037 76.3222
R3755 GNDA.n1548 GNDA.n1547 76.3222
R3756 GNDA.n1549 GNDA.n1517 76.3222
R3757 GNDA.n1556 GNDA.n1555 76.3222
R3758 GNDA.n1557 GNDA.n1515 76.3222
R3759 GNDA.n1564 GNDA.n1563 76.3222
R3760 GNDA.n1566 GNDA.n1513 76.3222
R3761 GNDA.n1698 GNDA.n1697 76.3222
R3762 GNDA.n1704 GNDA.n1703 76.3222
R3763 GNDA.n1705 GNDA.n1031 76.3222
R3764 GNDA.n1712 GNDA.n1711 76.3222
R3765 GNDA.n1713 GNDA.n1029 76.3222
R3766 GNDA.n1386 GNDA.n337 76.3222
R3767 GNDA.n1384 GNDA.n336 76.3222
R3768 GNDA.n1382 GNDA.n335 76.3222
R3769 GNDA.n1380 GNDA.n334 76.3222
R3770 GNDA.n1378 GNDA.n333 76.3222
R3771 GNDA.n1687 GNDA.n495 76.3222
R3772 GNDA.n1683 GNDA.n494 76.3222
R3773 GNDA.n1679 GNDA.n493 76.3222
R3774 GNDA.n1675 GNDA.n492 76.3222
R3775 GNDA.n1671 GNDA.n491 76.3222
R3776 GNDA.n1667 GNDA.n496 76.3222
R3777 GNDA.n1168 GNDA.n1167 76.3222
R3778 GNDA.n1057 GNDA.n1056 76.3222
R3779 GNDA.n1157 GNDA.n1156 76.3222
R3780 GNDA.n1066 GNDA.n1065 76.3222
R3781 GNDA.n1146 GNDA.n1145 76.3222
R3782 GNDA.n1073 GNDA.n1071 76.3222
R3783 GNDA.n1921 GNDA.n453 76.3222
R3784 GNDA.n1917 GNDA.n452 76.3222
R3785 GNDA.n1913 GNDA.n451 76.3222
R3786 GNDA.n1909 GNDA.n450 76.3222
R3787 GNDA.n1905 GNDA.n449 76.3222
R3788 GNDA.n707 GNDA.n448 76.3222
R3789 GNDA.n1945 GNDA.n1944 76.3222
R3790 GNDA.n1942 GNDA.n1941 76.3222
R3791 GNDA.n1937 GNDA.n688 76.3222
R3792 GNDA.n1934 GNDA.n687 76.3222
R3793 GNDA.n1930 GNDA.n686 76.3222
R3794 GNDA.n1926 GNDA.n685 76.3222
R3795 GNDA.n683 GNDA.n327 76.3222
R3796 GNDA.n1040 GNDA.n328 76.3222
R3797 GNDA.n1042 GNDA.n329 76.3222
R3798 GNDA.n1044 GNDA.n330 76.3222
R3799 GNDA.n1046 GNDA.n331 76.3222
R3800 GNDA.n1172 GNDA.n326 76.3222
R3801 GNDA.n1173 GNDA.n331 76.3222
R3802 GNDA.n1045 GNDA.n330 76.3222
R3803 GNDA.n1043 GNDA.n329 76.3222
R3804 GNDA.n1041 GNDA.n328 76.3222
R3805 GNDA.n1039 GNDA.n327 76.3222
R3806 GNDA.n1190 GNDA.n489 76.3222
R3807 GNDA.n1186 GNDA.n488 76.3222
R3808 GNDA.n1182 GNDA.n487 76.3222
R3809 GNDA.n1178 GNDA.n486 76.3222
R3810 GNDA.n1174 GNDA.n485 76.3222
R3811 GNDA.n1944 GNDA.n684 76.3222
R3812 GNDA.n1942 GNDA.n689 76.3222
R3813 GNDA.n1935 GNDA.n688 76.3222
R3814 GNDA.n1931 GNDA.n687 76.3222
R3815 GNDA.n1927 GNDA.n686 76.3222
R3816 GNDA.n1923 GNDA.n685 76.3222
R3817 GNDA.n1047 GNDA.n326 76.3222
R3818 GNDA.n1071 GNDA.n1067 76.3222
R3819 GNDA.n1147 GNDA.n1146 76.3222
R3820 GNDA.n1065 GNDA.n1058 76.3222
R3821 GNDA.n1158 GNDA.n1157 76.3222
R3822 GNDA.n1056 GNDA.n1049 76.3222
R3823 GNDA.n1169 GNDA.n1168 76.3222
R3824 GNDA.n1207 GNDA.n1206 76.3222
R3825 GNDA.n1234 GNDA.n1228 76.3222
R3826 GNDA.n1309 GNDA.n1308 76.3222
R3827 GNDA.n1226 GNDA.n1219 76.3222
R3828 GNDA.n1320 GNDA.n1319 76.3222
R3829 GNDA.n1217 GNDA.n1210 76.3222
R3830 GNDA.n1331 GNDA.n1330 76.3222
R3831 GNDA.n1231 GNDA.n497 76.3222
R3832 GNDA.n710 GNDA.n705 76.3222
R3833 GNDA.n703 GNDA.n702 76.3222
R3834 GNDA.n700 GNDA.n699 76.3222
R3835 GNDA.n697 GNDA.n696 76.3222
R3836 GNDA.n694 GNDA.n693 76.3222
R3837 GNDA.n1749 GNDA.n1748 76.3222
R3838 GNDA.n1741 GNDA.n1740 76.3222
R3839 GNDA.n1734 GNDA.n1025 76.3222
R3840 GNDA.n1732 GNDA.n1731 76.3222
R3841 GNDA.n1723 GNDA.n1722 76.3222
R3842 GNDA.n1918 GNDA.n453 76.3222
R3843 GNDA.n1914 GNDA.n452 76.3222
R3844 GNDA.n1910 GNDA.n451 76.3222
R3845 GNDA.n1906 GNDA.n450 76.3222
R3846 GNDA.n1902 GNDA.n449 76.3222
R3847 GNDA.n707 GNDA.n454 76.3222
R3848 GNDA.n1725 GNDA.n447 76.3222
R3849 GNDA.n1729 GNDA.n446 76.3222
R3850 GNDA.n1736 GNDA.n445 76.3222
R3851 GNDA.n1743 GNDA.n444 76.3222
R3852 GNDA.n1746 GNDA.n443 76.3222
R3853 GNDA.n2208 GNDA.n435 76.3222
R3854 GNDA.n2270 GNDA.n2269 76.3222
R3855 GNDA.n2264 GNDA.n260 76.3222
R3856 GNDA.n2261 GNDA.n261 76.3222
R3857 GNDA.n2257 GNDA.n262 76.3222
R3858 GNDA.n2253 GNDA.n263 76.3222
R3859 GNDA.n2162 GNDA.n466 76.3222
R3860 GNDA.n2161 GNDA.n2160 76.3222
R3861 GNDA.n2154 GNDA.n2138 76.3222
R3862 GNDA.n2153 GNDA.n2152 76.3222
R3863 GNDA.n2146 GNDA.n2140 76.3222
R3864 GNDA.n2145 GNDA.n2144 76.3222
R3865 GNDA.n2174 GNDA.n2173 76.3222
R3866 GNDA.n2177 GNDA.n2176 76.3222
R3867 GNDA.n2186 GNDA.n2185 76.3222
R3868 GNDA.n2189 GNDA.n2188 76.3222
R3869 GNDA.n2198 GNDA.n2197 76.3222
R3870 GNDA.n2201 GNDA.n2200 76.3222
R3871 GNDA.n2199 GNDA.n2198 76.3222
R3872 GNDA.n2188 GNDA.n462 76.3222
R3873 GNDA.n2187 GNDA.n2186 76.3222
R3874 GNDA.n2176 GNDA.n464 76.3222
R3875 GNDA.n2175 GNDA.n2174 76.3222
R3876 GNDA.n2171 GNDA.n441 76.3222
R3877 GNDA.n2179 GNDA.n440 76.3222
R3878 GNDA.n2183 GNDA.n439 76.3222
R3879 GNDA.n2191 GNDA.n438 76.3222
R3880 GNDA.n2195 GNDA.n437 76.3222
R3881 GNDA.n2205 GNDA.n436 76.3222
R3882 GNDA.n2178 GNDA.n441 76.3222
R3883 GNDA.n2182 GNDA.n440 76.3222
R3884 GNDA.n2190 GNDA.n439 76.3222
R3885 GNDA.n2194 GNDA.n438 76.3222
R3886 GNDA.n458 GNDA.n437 76.3222
R3887 GNDA.n2108 GNDA.n2107 76.3222
R3888 GNDA.n2113 GNDA.n2112 76.3222
R3889 GNDA.n2116 GNDA.n2115 76.3222
R3890 GNDA.n2130 GNDA.n2129 76.3222
R3891 GNDA.n2133 GNDA.n2132 76.3222
R3892 GNDA.n2106 GNDA.n321 76.3222
R3893 GNDA.n1949 GNDA.n322 76.3222
R3894 GNDA.n1954 GNDA.n323 76.3222
R3895 GNDA.n1960 GNDA.n324 76.3222
R3896 GNDA.n1966 GNDA.n325 76.3222
R3897 GNDA.n2096 GNDA.n320 76.3222
R3898 GNDA.n2095 GNDA.n325 76.3222
R3899 GNDA.n1965 GNDA.n324 76.3222
R3900 GNDA.n1959 GNDA.n323 76.3222
R3901 GNDA.n1953 GNDA.n322 76.3222
R3902 GNDA.n1948 GNDA.n321 76.3222
R3903 GNDA.n2103 GNDA.n478 76.3222
R3904 GNDA.n1955 GNDA.n483 76.3222
R3905 GNDA.n1961 GNDA.n482 76.3222
R3906 GNDA.n1967 GNDA.n481 76.3222
R3907 GNDA.n1970 GNDA.n480 76.3222
R3908 GNDA.n575 GNDA.n574 76.3222
R3909 GNDA.n570 GNDA.n569 76.3222
R3910 GNDA.n567 GNDA.n566 76.3222
R3911 GNDA.n562 GNDA.n561 76.3222
R3912 GNDA.n559 GNDA.n558 76.3222
R3913 GNDA.n2200 GNDA.n460 76.3222
R3914 GNDA.n1972 GNDA.n320 76.3222
R3915 GNDA.n1996 GNDA.n1993 76.3222
R3916 GNDA.n2071 GNDA.n2070 76.3222
R3917 GNDA.n1991 GNDA.n1984 76.3222
R3918 GNDA.n2082 GNDA.n2081 76.3222
R3919 GNDA.n1982 GNDA.n1975 76.3222
R3920 GNDA.n2093 GNDA.n2092 76.3222
R3921 GNDA.n2206 GNDA.n2205 76.3222
R3922 GNDA.n578 GNDA.n577 76.3222
R3923 GNDA.n676 GNDA.n675 76.3222
R3924 GNDA.n595 GNDA.n594 76.3222
R3925 GNDA.n605 GNDA.n604 76.3222
R3926 GNDA.n592 GNDA.n585 76.3222
R3927 GNDA.n616 GNDA.n615 76.3222
R3928 GNDA.n583 GNDA.n582 76.3222
R3929 GNDA.n2101 GNDA.n2100 76.3222
R3930 GNDA.n2163 GNDA.n2162 76.3222
R3931 GNDA.n2160 GNDA.n2159 76.3222
R3932 GNDA.n2155 GNDA.n2154 76.3222
R3933 GNDA.n2152 GNDA.n2151 76.3222
R3934 GNDA.n2147 GNDA.n2146 76.3222
R3935 GNDA.n2144 GNDA.n2143 76.3222
R3936 GNDA.n2107 GNDA.n473 76.3222
R3937 GNDA.n2114 GNDA.n2113 76.3222
R3938 GNDA.n2115 GNDA.n471 76.3222
R3939 GNDA.n2131 GNDA.n2130 76.3222
R3940 GNDA.n2134 GNDA.n2133 76.3222
R3941 GNDA.n554 GNDA.n553 76.3222
R3942 GNDA.n548 GNDA.n529 76.3222
R3943 GNDA.n546 GNDA.n545 76.3222
R3944 GNDA.n541 GNDA.n540 76.3222
R3945 GNDA.n538 GNDA.n537 76.3222
R3946 GNDA.n1848 GNDA.n999 76.3222
R3947 GNDA.n1846 GNDA.n1000 76.3222
R3948 GNDA.n2270 GNDA.n280 76.3222
R3949 GNDA.n2262 GNDA.n260 76.3222
R3950 GNDA.n2258 GNDA.n261 76.3222
R3951 GNDA.n2254 GNDA.n262 76.3222
R3952 GNDA.n2250 GNDA.n264 76.3222
R3953 GNDA.n974 GNDA.n265 76.3222
R3954 GNDA.n978 GNDA.n266 76.3222
R3955 GNDA.n982 GNDA.n267 76.3222
R3956 GNDA.n986 GNDA.n268 76.3222
R3957 GNDA.n969 GNDA.n270 76.3222
R3958 GNDA.n1868 GNDA.n271 76.3222
R3959 GNDA.n1864 GNDA.n272 76.3222
R3960 GNDA.n1860 GNDA.n273 76.3222
R3961 GNDA.n1856 GNDA.n274 76.3222
R3962 GNDA.n1852 GNDA.n276 76.3222
R3963 GNDA.n1270 GNDA.n1269 76.062
R3964 GNDA.n1269 GNDA.n1268 76.062
R3965 GNDA.n1108 GNDA.n1107 76.062
R3966 GNDA.n1107 GNDA.n1106 76.062
R3967 GNDA.n932 GNDA.n879 76.062
R3968 GNDA.n933 GNDA.n932 76.062
R3969 GNDA.n1622 GNDA.n1621 76.062
R3970 GNDA.n1621 GNDA.n1620 76.062
R3971 GNDA.n397 GNDA.n374 76.062
R3972 GNDA.n398 GNDA.n397 76.062
R3973 GNDA.n1808 GNDA.n1807 76.062
R3974 GNDA.n1807 GNDA.n1806 76.062
R3975 GNDA.n638 GNDA.n637 76.062
R3976 GNDA.n637 GNDA.n636 76.062
R3977 GNDA.n2032 GNDA.n2031 76.062
R3978 GNDA.n2031 GNDA.n2030 76.062
R3979 GNDA.n793 GNDA.n792 76.062
R3980 GNDA.n792 GNDA.n791 76.062
R3981 GNDA.n1431 GNDA.t190 75.8626
R3982 GNDA.n1423 GNDA.t165 75.8626
R3983 GNDA.t188 GNDA.n1423 75.8626
R3984 GNDA.n1472 GNDA.t161 75.8626
R3985 GNDA.n1472 GNDA.t1 75.8626
R3986 GNDA.t41 GNDA.n1471 75.8626
R3987 GNDA.t287 GNDA.t159 75.8626
R3988 GNDA.t308 GNDA.t78 75.8626
R3989 GNDA.n1326 GNDA.n1212 74.5978
R3990 GNDA.n1253 GNDA.n1212 74.5978
R3991 GNDA.n1164 GNDA.n1051 74.5978
R3992 GNDA.n1091 GNDA.n1051 74.5978
R3993 GNDA.n916 GNDA.n915 74.5978
R3994 GNDA.n917 GNDA.n916 74.5978
R3995 GNDA.n1604 GNDA.n1603 74.5978
R3996 GNDA.n1605 GNDA.n1604 74.5978
R3997 GNDA.n381 GNDA.n346 74.5978
R3998 GNDA.n382 GNDA.n381 74.5978
R3999 GNDA.n1790 GNDA.n1789 74.5978
R4000 GNDA.n1791 GNDA.n1790 74.5978
R4001 GNDA.n620 GNDA.n619 74.5978
R4002 GNDA.n621 GNDA.n620 74.5978
R4003 GNDA.n2088 GNDA.n1977 74.5978
R4004 GNDA.n2015 GNDA.n1977 74.5978
R4005 GNDA.n775 GNDA.n774 74.5978
R4006 GNDA.n776 GNDA.n775 74.5978
R4007 GNDA.t224 GNDA.n314 73.8684
R4008 GNDA.n207 GNDA.t338 72.3996
R4009 GNDA.t101 GNDA.n109 72.3996
R4010 GNDA.t79 GNDA.n2340 72.3996
R4011 GNDA.n2373 GNDA.t77 72.3996
R4012 GNDA.n2387 GNDA.t320 71.648
R4013 GNDA.n201 GNDA.n115 70.0642
R4014 GNDA.n2350 GNDA.n2347 70.0642
R4015 GNDA.t184 GNDA.t187 69.5407
R4016 GNDA.t187 GNDA.t150 69.5407
R4017 GNDA.t67 GNDA.n1479 69.5407
R4018 GNDA.n1479 GNDA.t144 69.5407
R4019 GNDA.t142 GNDA.t162 69.5407
R4020 GNDA.t162 GNDA.t48 69.5407
R4021 GNDA.n1255 GNDA.t244 65.8183
R4022 GNDA.n1261 GNDA.t244 65.8183
R4023 GNDA.n1263 GNDA.t244 65.8183
R4024 GNDA.n1271 GNDA.t244 65.8183
R4025 GNDA.n1277 GNDA.t244 65.8183
R4026 GNDA.n1279 GNDA.t244 65.8183
R4027 GNDA.n1285 GNDA.t244 65.8183
R4028 GNDA.n1302 GNDA.t244 65.8183
R4029 GNDA.n1296 GNDA.t244 65.8183
R4030 GNDA.n1294 GNDA.t244 65.8183
R4031 GNDA.n1288 GNDA.t244 65.8183
R4032 GNDA.n1093 GNDA.t223 65.8183
R4033 GNDA.n1099 GNDA.t223 65.8183
R4034 GNDA.n1101 GNDA.t223 65.8183
R4035 GNDA.n1109 GNDA.t223 65.8183
R4036 GNDA.n1115 GNDA.t223 65.8183
R4037 GNDA.n1117 GNDA.t223 65.8183
R4038 GNDA.n1123 GNDA.t223 65.8183
R4039 GNDA.n1140 GNDA.t223 65.8183
R4040 GNDA.n1134 GNDA.t223 65.8183
R4041 GNDA.n1132 GNDA.t223 65.8183
R4042 GNDA.n1126 GNDA.t223 65.8183
R4043 GNDA.n922 GNDA.t310 65.8183
R4044 GNDA.n924 GNDA.t310 65.8183
R4045 GNDA.n930 GNDA.t310 65.8183
R4046 GNDA.n938 GNDA.t310 65.8183
R4047 GNDA.n940 GNDA.t310 65.8183
R4048 GNDA.n946 GNDA.t310 65.8183
R4049 GNDA.n948 GNDA.t310 65.8183
R4050 GNDA.n966 GNDA.t310 65.8183
R4051 GNDA.n963 GNDA.t310 65.8183
R4052 GNDA.n957 GNDA.t310 65.8183
R4053 GNDA.n954 GNDA.t310 65.8183
R4054 GNDA.n1607 GNDA.t248 65.8183
R4055 GNDA.n1613 GNDA.t248 65.8183
R4056 GNDA.n1615 GNDA.t248 65.8183
R4057 GNDA.n1623 GNDA.t248 65.8183
R4058 GNDA.n1629 GNDA.t248 65.8183
R4059 GNDA.n1631 GNDA.t248 65.8183
R4060 GNDA.n1637 GNDA.t248 65.8183
R4061 GNDA.n1654 GNDA.t248 65.8183
R4062 GNDA.n1648 GNDA.t248 65.8183
R4063 GNDA.n1646 GNDA.t248 65.8183
R4064 GNDA.n1640 GNDA.t248 65.8183
R4065 GNDA.n387 GNDA.t250 65.8183
R4066 GNDA.n389 GNDA.t250 65.8183
R4067 GNDA.n395 GNDA.t250 65.8183
R4068 GNDA.n403 GNDA.t250 65.8183
R4069 GNDA.n405 GNDA.t250 65.8183
R4070 GNDA.n411 GNDA.t250 65.8183
R4071 GNDA.n413 GNDA.t250 65.8183
R4072 GNDA.n431 GNDA.t250 65.8183
R4073 GNDA.n428 GNDA.t250 65.8183
R4074 GNDA.n422 GNDA.t250 65.8183
R4075 GNDA.n419 GNDA.t250 65.8183
R4076 GNDA.n1793 GNDA.t234 65.8183
R4077 GNDA.n1799 GNDA.t234 65.8183
R4078 GNDA.n1801 GNDA.t234 65.8183
R4079 GNDA.n1809 GNDA.t234 65.8183
R4080 GNDA.n1815 GNDA.t234 65.8183
R4081 GNDA.n1817 GNDA.t234 65.8183
R4082 GNDA.n1823 GNDA.t234 65.8183
R4083 GNDA.n1840 GNDA.t234 65.8183
R4084 GNDA.n1834 GNDA.t234 65.8183
R4085 GNDA.n1832 GNDA.t234 65.8183
R4086 GNDA.n1826 GNDA.t234 65.8183
R4087 GNDA.t234 GNDA.n1003 65.8183
R4088 GNDA.n1767 GNDA.t234 65.8183
R4089 GNDA.n1778 GNDA.t234 65.8183
R4090 GNDA.n1762 GNDA.t234 65.8183
R4091 GNDA.n364 GNDA.t250 65.8183
R4092 GNDA.n2222 GNDA.t250 65.8183
R4093 GNDA.n351 GNDA.t250 65.8183
R4094 GNDA.n2233 GNDA.t250 65.8183
R4095 GNDA.t248 GNDA.n1491 65.8183
R4096 GNDA.n1581 GNDA.t248 65.8183
R4097 GNDA.n1592 GNDA.t248 65.8183
R4098 GNDA.n1576 GNDA.t248 65.8183
R4099 GNDA.n896 GNDA.t310 65.8183
R4100 GNDA.n893 GNDA.t310 65.8183
R4101 GNDA.n907 GNDA.t310 65.8183
R4102 GNDA.n888 GNDA.t310 65.8183
R4103 GNDA.n1069 GNDA.t223 65.8183
R4104 GNDA.n1151 GNDA.t223 65.8183
R4105 GNDA.n1060 GNDA.t223 65.8183
R4106 GNDA.n1162 GNDA.t223 65.8183
R4107 GNDA.n1230 GNDA.t244 65.8183
R4108 GNDA.n1313 GNDA.t244 65.8183
R4109 GNDA.n1221 GNDA.t244 65.8183
R4110 GNDA.n1324 GNDA.t244 65.8183
R4111 GNDA.n623 GNDA.t264 65.8183
R4112 GNDA.n629 GNDA.t264 65.8183
R4113 GNDA.n631 GNDA.t264 65.8183
R4114 GNDA.n639 GNDA.t264 65.8183
R4115 GNDA.n645 GNDA.t264 65.8183
R4116 GNDA.n647 GNDA.t264 65.8183
R4117 GNDA.n653 GNDA.t264 65.8183
R4118 GNDA.n670 GNDA.t264 65.8183
R4119 GNDA.n664 GNDA.t264 65.8183
R4120 GNDA.n662 GNDA.t264 65.8183
R4121 GNDA.n656 GNDA.t264 65.8183
R4122 GNDA.n2017 GNDA.t277 65.8183
R4123 GNDA.n2023 GNDA.t277 65.8183
R4124 GNDA.n2025 GNDA.t277 65.8183
R4125 GNDA.n2033 GNDA.t277 65.8183
R4126 GNDA.n2039 GNDA.t277 65.8183
R4127 GNDA.n2041 GNDA.t277 65.8183
R4128 GNDA.n2047 GNDA.t277 65.8183
R4129 GNDA.n2064 GNDA.t277 65.8183
R4130 GNDA.n2058 GNDA.t277 65.8183
R4131 GNDA.n2056 GNDA.t277 65.8183
R4132 GNDA.n2050 GNDA.t277 65.8183
R4133 GNDA.n778 GNDA.t249 65.8183
R4134 GNDA.n784 GNDA.t249 65.8183
R4135 GNDA.n786 GNDA.t249 65.8183
R4136 GNDA.n794 GNDA.t249 65.8183
R4137 GNDA.n800 GNDA.t249 65.8183
R4138 GNDA.n802 GNDA.t249 65.8183
R4139 GNDA.n808 GNDA.t249 65.8183
R4140 GNDA.n825 GNDA.t249 65.8183
R4141 GNDA.n819 GNDA.t249 65.8183
R4142 GNDA.n817 GNDA.t249 65.8183
R4143 GNDA.n811 GNDA.t249 65.8183
R4144 GNDA.t249 GNDA.n728 65.8183
R4145 GNDA.n755 GNDA.t249 65.8183
R4146 GNDA.n766 GNDA.t249 65.8183
R4147 GNDA.n750 GNDA.t249 65.8183
R4148 GNDA.n1995 GNDA.t277 65.8183
R4149 GNDA.n2075 GNDA.t277 65.8183
R4150 GNDA.n1986 GNDA.t277 65.8183
R4151 GNDA.n2086 GNDA.t277 65.8183
R4152 GNDA.t264 GNDA.n502 65.8183
R4153 GNDA.n597 GNDA.t264 65.8183
R4154 GNDA.n609 GNDA.t264 65.8183
R4155 GNDA.n587 GNDA.t264 65.8183
R4156 GNDA.n2403 GNDA.n78 64.0005
R4157 GNDA.n2403 GNDA.n65 64.0005
R4158 GNDA.n1424 GNDA.t188 63.2189
R4159 GNDA.t161 GNDA.n219 63.2189
R4160 GNDA.t329 GNDA.t58 63.2189
R4161 GNDA.t82 GNDA.t74 63.2189
R4162 GNDA.t87 GNDA.t171 63.2189
R4163 GNDA.t30 GNDA.t13 63.2189
R4164 GNDA.n1571 GNDA.n1511 60.474
R4165 GNDA.t50 GNDA.t97 59.0043
R4166 GNDA.t170 GNDA.t239 59.0043
R4167 GNDA.t302 GNDA.t5 59.0043
R4168 GNDA.t86 GNDA.t290 59.0043
R4169 GNDA.t99 GNDA.t173 59.0043
R4170 GNDA.t3 GNDA.t12 59.0043
R4171 GNDA.t299 GNDA.t189 56.897
R4172 GNDA.t93 GNDA.t138 56.897
R4173 GNDA.n1425 GNDA.t246 56.897
R4174 GNDA.t262 GNDA.n2324 56.897
R4175 GNDA.t154 GNDA.t318 56.897
R4176 GNDA.t47 GNDA.t275 56.897
R4177 GNDA.n534 GNDA.n533 56.3995
R4178 GNDA.n533 GNDA.n477 56.3995
R4179 GNDA.n2169 GNDA.n2168 56.3995
R4180 GNDA.n2170 GNDA.n2169 56.3995
R4181 GNDA.n2287 GNDA.n2286 56.2142
R4182 GNDA.n1790 GNDA.t234 55.2026
R4183 GNDA.n381 GNDA.t250 55.2026
R4184 GNDA.n1604 GNDA.t248 55.2026
R4185 GNDA.n916 GNDA.t310 55.2026
R4186 GNDA.t223 GNDA.n1051 55.2026
R4187 GNDA.t244 GNDA.n1212 55.2026
R4188 GNDA.n775 GNDA.t249 55.2026
R4189 GNDA.t277 GNDA.n1977 55.2026
R4190 GNDA.n620 GNDA.t264 55.2026
R4191 GNDA.n95 GNDA.t343 54.7898
R4192 GNDA.t122 GNDA.n143 54.7898
R4193 GNDA.n1269 GNDA.t244 54.4705
R4194 GNDA.n1107 GNDA.t223 54.4705
R4195 GNDA.n932 GNDA.t310 54.4705
R4196 GNDA.n1621 GNDA.t248 54.4705
R4197 GNDA.n397 GNDA.t250 54.4705
R4198 GNDA.n1807 GNDA.t234 54.4705
R4199 GNDA.n637 GNDA.t264 54.4705
R4200 GNDA.n2031 GNDA.t277 54.4705
R4201 GNDA.n792 GNDA.t249 54.4705
R4202 GNDA.n2414 GNDA.n35 54.4005
R4203 GNDA.n1324 GNDA.n1323 53.3664
R4204 GNDA.n1315 GNDA.n1221 53.3664
R4205 GNDA.n1313 GNDA.n1312 53.3664
R4206 GNDA.n1304 GNDA.n1230 53.3664
R4207 GNDA.n1288 GNDA.n1287 53.3664
R4208 GNDA.n1294 GNDA.n1293 53.3664
R4209 GNDA.n1297 GNDA.n1296 53.3664
R4210 GNDA.n1302 GNDA.n1301 53.3664
R4211 GNDA.n1272 GNDA.n1271 53.3664
R4212 GNDA.n1277 GNDA.n1276 53.3664
R4213 GNDA.n1280 GNDA.n1279 53.3664
R4214 GNDA.n1285 GNDA.n1284 53.3664
R4215 GNDA.n1263 GNDA.n1248 53.3664
R4216 GNDA.n1262 GNDA.n1261 53.3664
R4217 GNDA.n1255 GNDA.n1250 53.3664
R4218 GNDA.n1256 GNDA.n1255 53.3664
R4219 GNDA.n1261 GNDA.n1260 53.3664
R4220 GNDA.n1264 GNDA.n1263 53.3664
R4221 GNDA.n1271 GNDA.n1246 53.3664
R4222 GNDA.n1278 GNDA.n1277 53.3664
R4223 GNDA.n1279 GNDA.n1244 53.3664
R4224 GNDA.n1286 GNDA.n1285 53.3664
R4225 GNDA.n1303 GNDA.n1302 53.3664
R4226 GNDA.n1296 GNDA.n1239 53.3664
R4227 GNDA.n1295 GNDA.n1294 53.3664
R4228 GNDA.n1289 GNDA.n1288 53.3664
R4229 GNDA.n1162 GNDA.n1161 53.3664
R4230 GNDA.n1153 GNDA.n1060 53.3664
R4231 GNDA.n1151 GNDA.n1150 53.3664
R4232 GNDA.n1142 GNDA.n1069 53.3664
R4233 GNDA.n1126 GNDA.n1125 53.3664
R4234 GNDA.n1132 GNDA.n1131 53.3664
R4235 GNDA.n1135 GNDA.n1134 53.3664
R4236 GNDA.n1140 GNDA.n1139 53.3664
R4237 GNDA.n1110 GNDA.n1109 53.3664
R4238 GNDA.n1115 GNDA.n1114 53.3664
R4239 GNDA.n1118 GNDA.n1117 53.3664
R4240 GNDA.n1123 GNDA.n1122 53.3664
R4241 GNDA.n1101 GNDA.n1086 53.3664
R4242 GNDA.n1100 GNDA.n1099 53.3664
R4243 GNDA.n1093 GNDA.n1088 53.3664
R4244 GNDA.n1094 GNDA.n1093 53.3664
R4245 GNDA.n1099 GNDA.n1098 53.3664
R4246 GNDA.n1102 GNDA.n1101 53.3664
R4247 GNDA.n1109 GNDA.n1084 53.3664
R4248 GNDA.n1116 GNDA.n1115 53.3664
R4249 GNDA.n1117 GNDA.n1082 53.3664
R4250 GNDA.n1124 GNDA.n1123 53.3664
R4251 GNDA.n1141 GNDA.n1140 53.3664
R4252 GNDA.n1134 GNDA.n1077 53.3664
R4253 GNDA.n1133 GNDA.n1132 53.3664
R4254 GNDA.n1127 GNDA.n1126 53.3664
R4255 GNDA.n909 GNDA.n888 53.3664
R4256 GNDA.n907 GNDA.n906 53.3664
R4257 GNDA.n898 GNDA.n893 53.3664
R4258 GNDA.n896 GNDA.n870 53.3664
R4259 GNDA.n954 GNDA.n953 53.3664
R4260 GNDA.n958 GNDA.n957 53.3664
R4261 GNDA.n963 GNDA.n962 53.3664
R4262 GNDA.n966 GNDA.n965 53.3664
R4263 GNDA.n938 GNDA.n937 53.3664
R4264 GNDA.n941 GNDA.n940 53.3664
R4265 GNDA.n946 GNDA.n945 53.3664
R4266 GNDA.n949 GNDA.n948 53.3664
R4267 GNDA.n931 GNDA.n930 53.3664
R4268 GNDA.n924 GNDA.n881 53.3664
R4269 GNDA.n923 GNDA.n922 53.3664
R4270 GNDA.n922 GNDA.n921 53.3664
R4271 GNDA.n925 GNDA.n924 53.3664
R4272 GNDA.n930 GNDA.n929 53.3664
R4273 GNDA.n939 GNDA.n938 53.3664
R4274 GNDA.n940 GNDA.n877 53.3664
R4275 GNDA.n947 GNDA.n946 53.3664
R4276 GNDA.n948 GNDA.n875 53.3664
R4277 GNDA.n967 GNDA.n966 53.3664
R4278 GNDA.n964 GNDA.n963 53.3664
R4279 GNDA.n957 GNDA.n872 53.3664
R4280 GNDA.n955 GNDA.n954 53.3664
R4281 GNDA.n1577 GNDA.n1576 53.3664
R4282 GNDA.n1592 GNDA.n1591 53.3664
R4283 GNDA.n1583 GNDA.n1581 53.3664
R4284 GNDA.n1656 GNDA.n1491 53.3664
R4285 GNDA.n1640 GNDA.n1639 53.3664
R4286 GNDA.n1646 GNDA.n1645 53.3664
R4287 GNDA.n1649 GNDA.n1648 53.3664
R4288 GNDA.n1654 GNDA.n1653 53.3664
R4289 GNDA.n1624 GNDA.n1623 53.3664
R4290 GNDA.n1629 GNDA.n1628 53.3664
R4291 GNDA.n1632 GNDA.n1631 53.3664
R4292 GNDA.n1637 GNDA.n1636 53.3664
R4293 GNDA.n1615 GNDA.n1503 53.3664
R4294 GNDA.n1614 GNDA.n1613 53.3664
R4295 GNDA.n1607 GNDA.n1505 53.3664
R4296 GNDA.n1608 GNDA.n1607 53.3664
R4297 GNDA.n1613 GNDA.n1612 53.3664
R4298 GNDA.n1616 GNDA.n1615 53.3664
R4299 GNDA.n1623 GNDA.n1501 53.3664
R4300 GNDA.n1630 GNDA.n1629 53.3664
R4301 GNDA.n1631 GNDA.n1499 53.3664
R4302 GNDA.n1638 GNDA.n1637 53.3664
R4303 GNDA.n1655 GNDA.n1654 53.3664
R4304 GNDA.n1648 GNDA.n1494 53.3664
R4305 GNDA.n1647 GNDA.n1646 53.3664
R4306 GNDA.n1641 GNDA.n1640 53.3664
R4307 GNDA.n2233 GNDA.n2232 53.3664
R4308 GNDA.n2224 GNDA.n351 53.3664
R4309 GNDA.n2222 GNDA.n2221 53.3664
R4310 GNDA.n365 GNDA.n364 53.3664
R4311 GNDA.n419 GNDA.n418 53.3664
R4312 GNDA.n423 GNDA.n422 53.3664
R4313 GNDA.n428 GNDA.n427 53.3664
R4314 GNDA.n431 GNDA.n430 53.3664
R4315 GNDA.n403 GNDA.n402 53.3664
R4316 GNDA.n406 GNDA.n405 53.3664
R4317 GNDA.n411 GNDA.n410 53.3664
R4318 GNDA.n414 GNDA.n413 53.3664
R4319 GNDA.n396 GNDA.n395 53.3664
R4320 GNDA.n389 GNDA.n376 53.3664
R4321 GNDA.n388 GNDA.n387 53.3664
R4322 GNDA.n387 GNDA.n386 53.3664
R4323 GNDA.n390 GNDA.n389 53.3664
R4324 GNDA.n395 GNDA.n394 53.3664
R4325 GNDA.n404 GNDA.n403 53.3664
R4326 GNDA.n405 GNDA.n372 53.3664
R4327 GNDA.n412 GNDA.n411 53.3664
R4328 GNDA.n413 GNDA.n370 53.3664
R4329 GNDA.n432 GNDA.n431 53.3664
R4330 GNDA.n429 GNDA.n428 53.3664
R4331 GNDA.n422 GNDA.n367 53.3664
R4332 GNDA.n420 GNDA.n419 53.3664
R4333 GNDA.n1763 GNDA.n1762 53.3664
R4334 GNDA.n1778 GNDA.n1777 53.3664
R4335 GNDA.n1769 GNDA.n1767 53.3664
R4336 GNDA.n1842 GNDA.n1003 53.3664
R4337 GNDA.n1826 GNDA.n1825 53.3664
R4338 GNDA.n1832 GNDA.n1831 53.3664
R4339 GNDA.n1835 GNDA.n1834 53.3664
R4340 GNDA.n1840 GNDA.n1839 53.3664
R4341 GNDA.n1810 GNDA.n1809 53.3664
R4342 GNDA.n1815 GNDA.n1814 53.3664
R4343 GNDA.n1818 GNDA.n1817 53.3664
R4344 GNDA.n1823 GNDA.n1822 53.3664
R4345 GNDA.n1801 GNDA.n1014 53.3664
R4346 GNDA.n1800 GNDA.n1799 53.3664
R4347 GNDA.n1793 GNDA.n1016 53.3664
R4348 GNDA.n1794 GNDA.n1793 53.3664
R4349 GNDA.n1799 GNDA.n1798 53.3664
R4350 GNDA.n1802 GNDA.n1801 53.3664
R4351 GNDA.n1809 GNDA.n1012 53.3664
R4352 GNDA.n1816 GNDA.n1815 53.3664
R4353 GNDA.n1817 GNDA.n1010 53.3664
R4354 GNDA.n1824 GNDA.n1823 53.3664
R4355 GNDA.n1841 GNDA.n1840 53.3664
R4356 GNDA.n1834 GNDA.n1005 53.3664
R4357 GNDA.n1833 GNDA.n1832 53.3664
R4358 GNDA.n1827 GNDA.n1826 53.3664
R4359 GNDA.n1768 GNDA.n1003 53.3664
R4360 GNDA.n1767 GNDA.n1764 53.3664
R4361 GNDA.n1779 GNDA.n1778 53.3664
R4362 GNDA.n1762 GNDA.n1019 53.3664
R4363 GNDA.n364 GNDA.n353 53.3664
R4364 GNDA.n2223 GNDA.n2222 53.3664
R4365 GNDA.n351 GNDA.n347 53.3664
R4366 GNDA.n2234 GNDA.n2233 53.3664
R4367 GNDA.n1582 GNDA.n1491 53.3664
R4368 GNDA.n1581 GNDA.n1578 53.3664
R4369 GNDA.n1593 GNDA.n1592 53.3664
R4370 GNDA.n1576 GNDA.n1508 53.3664
R4371 GNDA.n897 GNDA.n896 53.3664
R4372 GNDA.n893 GNDA.n890 53.3664
R4373 GNDA.n908 GNDA.n907 53.3664
R4374 GNDA.n888 GNDA.n885 53.3664
R4375 GNDA.n1069 GNDA.n1062 53.3664
R4376 GNDA.n1152 GNDA.n1151 53.3664
R4377 GNDA.n1060 GNDA.n1053 53.3664
R4378 GNDA.n1163 GNDA.n1162 53.3664
R4379 GNDA.n1230 GNDA.n1223 53.3664
R4380 GNDA.n1314 GNDA.n1313 53.3664
R4381 GNDA.n1221 GNDA.n1214 53.3664
R4382 GNDA.n1325 GNDA.n1324 53.3664
R4383 GNDA.n611 GNDA.n587 53.3664
R4384 GNDA.n609 GNDA.n608 53.3664
R4385 GNDA.n600 GNDA.n597 53.3664
R4386 GNDA.n672 GNDA.n502 53.3664
R4387 GNDA.n656 GNDA.n655 53.3664
R4388 GNDA.n662 GNDA.n661 53.3664
R4389 GNDA.n665 GNDA.n664 53.3664
R4390 GNDA.n670 GNDA.n669 53.3664
R4391 GNDA.n640 GNDA.n639 53.3664
R4392 GNDA.n645 GNDA.n644 53.3664
R4393 GNDA.n648 GNDA.n647 53.3664
R4394 GNDA.n653 GNDA.n652 53.3664
R4395 GNDA.n631 GNDA.n513 53.3664
R4396 GNDA.n630 GNDA.n629 53.3664
R4397 GNDA.n623 GNDA.n515 53.3664
R4398 GNDA.n624 GNDA.n623 53.3664
R4399 GNDA.n629 GNDA.n628 53.3664
R4400 GNDA.n632 GNDA.n631 53.3664
R4401 GNDA.n639 GNDA.n511 53.3664
R4402 GNDA.n646 GNDA.n645 53.3664
R4403 GNDA.n647 GNDA.n509 53.3664
R4404 GNDA.n654 GNDA.n653 53.3664
R4405 GNDA.n671 GNDA.n670 53.3664
R4406 GNDA.n664 GNDA.n504 53.3664
R4407 GNDA.n663 GNDA.n662 53.3664
R4408 GNDA.n657 GNDA.n656 53.3664
R4409 GNDA.n2086 GNDA.n2085 53.3664
R4410 GNDA.n2077 GNDA.n1986 53.3664
R4411 GNDA.n2075 GNDA.n2074 53.3664
R4412 GNDA.n2066 GNDA.n1995 53.3664
R4413 GNDA.n2050 GNDA.n2049 53.3664
R4414 GNDA.n2056 GNDA.n2055 53.3664
R4415 GNDA.n2059 GNDA.n2058 53.3664
R4416 GNDA.n2064 GNDA.n2063 53.3664
R4417 GNDA.n2034 GNDA.n2033 53.3664
R4418 GNDA.n2039 GNDA.n2038 53.3664
R4419 GNDA.n2042 GNDA.n2041 53.3664
R4420 GNDA.n2047 GNDA.n2046 53.3664
R4421 GNDA.n2025 GNDA.n2010 53.3664
R4422 GNDA.n2024 GNDA.n2023 53.3664
R4423 GNDA.n2017 GNDA.n2012 53.3664
R4424 GNDA.n2018 GNDA.n2017 53.3664
R4425 GNDA.n2023 GNDA.n2022 53.3664
R4426 GNDA.n2026 GNDA.n2025 53.3664
R4427 GNDA.n2033 GNDA.n2008 53.3664
R4428 GNDA.n2040 GNDA.n2039 53.3664
R4429 GNDA.n2041 GNDA.n2006 53.3664
R4430 GNDA.n2048 GNDA.n2047 53.3664
R4431 GNDA.n2065 GNDA.n2064 53.3664
R4432 GNDA.n2058 GNDA.n2001 53.3664
R4433 GNDA.n2057 GNDA.n2056 53.3664
R4434 GNDA.n2051 GNDA.n2050 53.3664
R4435 GNDA.n768 GNDA.n750 53.3664
R4436 GNDA.n766 GNDA.n765 53.3664
R4437 GNDA.n757 GNDA.n755 53.3664
R4438 GNDA.n827 GNDA.n728 53.3664
R4439 GNDA.n811 GNDA.n810 53.3664
R4440 GNDA.n817 GNDA.n816 53.3664
R4441 GNDA.n820 GNDA.n819 53.3664
R4442 GNDA.n825 GNDA.n824 53.3664
R4443 GNDA.n795 GNDA.n794 53.3664
R4444 GNDA.n800 GNDA.n799 53.3664
R4445 GNDA.n803 GNDA.n802 53.3664
R4446 GNDA.n808 GNDA.n807 53.3664
R4447 GNDA.n786 GNDA.n740 53.3664
R4448 GNDA.n785 GNDA.n784 53.3664
R4449 GNDA.n778 GNDA.n742 53.3664
R4450 GNDA.n779 GNDA.n778 53.3664
R4451 GNDA.n784 GNDA.n783 53.3664
R4452 GNDA.n787 GNDA.n786 53.3664
R4453 GNDA.n794 GNDA.n738 53.3664
R4454 GNDA.n801 GNDA.n800 53.3664
R4455 GNDA.n802 GNDA.n736 53.3664
R4456 GNDA.n809 GNDA.n808 53.3664
R4457 GNDA.n826 GNDA.n825 53.3664
R4458 GNDA.n819 GNDA.n731 53.3664
R4459 GNDA.n818 GNDA.n817 53.3664
R4460 GNDA.n812 GNDA.n811 53.3664
R4461 GNDA.n756 GNDA.n728 53.3664
R4462 GNDA.n755 GNDA.n752 53.3664
R4463 GNDA.n767 GNDA.n766 53.3664
R4464 GNDA.n750 GNDA.n745 53.3664
R4465 GNDA.n1995 GNDA.n1988 53.3664
R4466 GNDA.n2076 GNDA.n2075 53.3664
R4467 GNDA.n1986 GNDA.n1979 53.3664
R4468 GNDA.n2087 GNDA.n2086 53.3664
R4469 GNDA.n599 GNDA.n502 53.3664
R4470 GNDA.n597 GNDA.n589 53.3664
R4471 GNDA.n610 GNDA.n609 53.3664
R4472 GNDA.n587 GNDA.n518 53.3664
R4473 GNDA.n78 GNDA.n77 51.2005
R4474 GNDA.n71 GNDA.n65 51.2005
R4475 GNDA.n2293 GNDA.n241 51.1039
R4476 GNDA.n2373 GNDA.n2372 50.5752
R4477 GNDA.n207 GNDA.n110 50.5752
R4478 GNDA.t42 GNDA.n191 49.0451
R4479 GNDA.n2341 GNDA.t9 49.0451
R4480 GNDA.n49 GNDA.t213 48.0005
R4481 GNDA.n49 GNDA.t203 48.0005
R4482 GNDA.n46 GNDA.t217 48.0005
R4483 GNDA.n46 GNDA.t205 48.0005
R4484 GNDA.n45 GNDA.t211 48.0005
R4485 GNDA.n45 GNDA.t201 48.0005
R4486 GNDA.n43 GNDA.t215 48.0005
R4487 GNDA.n43 GNDA.t207 48.0005
R4488 GNDA.n42 GNDA.t219 48.0005
R4489 GNDA.n42 GNDA.t209 48.0005
R4490 GNDA.t224 GNDA.n2243 47.6748
R4491 GNDA.t28 GNDA.t335 46.3607
R4492 GNDA.t28 GNDA.t112 46.3607
R4493 GNDA.t5 GNDA.n2405 46.3607
R4494 GNDA.t33 GNDA.t175 46.3607
R4495 GNDA.t33 GNDA.t95 46.3607
R4496 GNDA.n198 GNDA.n197 44.8005
R4497 GNDA.n2354 GNDA.n2353 44.8005
R4498 GNDA.t10 GNDA.t39 44.2534
R4499 GNDA.t148 GNDA.t319 44.2534
R4500 GNDA.t344 GNDA.t266 42.1461
R4501 GNDA.t322 GNDA.t24 42.1461
R4502 GNDA.t7 GNDA.t115 42.1461
R4503 GNDA.t315 GNDA.t16 42.1461
R4504 GNDA.t325 GNDA.t60 42.1461
R4505 GNDA.t27 GNDA.t18 42.1461
R4506 GNDA.t158 GNDA.t117 42.1461
R4507 GNDA.t226 GNDA.t35 42.1461
R4508 GNDA.t62 GNDA.t293 42.1461
R4509 GNDA.t341 GNDA.t321 42.1461
R4510 GNDA.t326 GNDA.t125 42.1461
R4511 GNDA.t91 GNDA.t0 42.1461
R4512 GNDA.t156 GNDA.t2 42.1461
R4513 GNDA.t119 GNDA.t127 42.1461
R4514 GNDA.t110 GNDA.t84 42.1461
R4515 GNDA.t51 GNDA.t8 42.1461
R4516 GNDA.t252 GNDA.t177 42.1461
R4517 GNDA.t104 GNDA.n200 39.7033
R4518 GNDA.n2351 GNDA.t108 39.7033
R4519 GNDA.t112 GNDA.n95 37.9315
R4520 GNDA.n2412 GNDA.t348 37.9315
R4521 GNDA.t11 GNDA.t86 37.9315
R4522 GNDA.n143 GNDA.t175 37.9315
R4523 GNDA.n2306 GNDA.n2305 36.4143
R4524 GNDA.n23 GNDA.n22 34.813
R4525 GNDA.n2425 GNDA.n11 34.813
R4526 GNDA.n2385 GNDA.n80 33.717
R4527 GNDA.t266 GNDA.t65 33.717
R4528 GNDA.t333 GNDA.t23 33.717
R4529 GNDA.t24 GNDA.t314 33.717
R4530 GNDA.t115 GNDA.t44 33.717
R4531 GNDA.t16 GNDA.t166 33.717
R4532 GNDA.t60 GNDA.t32 33.717
R4533 GNDA.t18 GNDA.t46 33.717
R4534 GNDA.t117 GNDA.t339 33.717
R4535 GNDA.t35 GNDA.t50 33.717
R4536 GNDA.t97 GNDA.t170 33.717
R4537 GNDA.t239 GNDA.t302 33.717
R4538 GNDA.t290 GNDA.t99 33.717
R4539 GNDA.t173 GNDA.t3 33.717
R4540 GNDA.t12 GNDA.t62 33.717
R4541 GNDA.t181 GNDA.t326 33.717
R4542 GNDA.t59 GNDA.t91 33.717
R4543 GNDA.t126 GNDA.t156 33.717
R4544 GNDA.t131 GNDA.t119 33.717
R4545 GNDA.t316 GNDA.t110 33.717
R4546 GNDA.t57 GNDA.t51 33.717
R4547 GNDA.t94 GNDA.t252 33.717
R4548 GNDA.n145 GNDA.n144 33.717
R4549 GNDA.t224 GNDA.n318 32.9056
R4550 GNDA.t224 GNDA.n317 32.9056
R4551 GNDA.t182 GNDA.t190 31.6097
R4552 GNDA.t167 GNDA.t134 31.6097
R4553 GNDA.t128 GNDA.t136 31.6097
R4554 GNDA.t37 GNDA.t41 31.6097
R4555 GNDA.n117 GNDA.t338 30.3614
R4556 GNDA.n192 GNDA.t66 30.3614
R4557 GNDA.n2358 GNDA.t72 30.3614
R4558 GNDA.n2344 GNDA.t77 30.3614
R4559 GNDA.t160 GNDA.t329 29.5024
R4560 GNDA.t343 GNDA.t82 29.5024
R4561 GNDA.n2420 GNDA.t341 29.5024
R4562 GNDA.t171 GNDA.t122 29.5024
R4563 GNDA.t45 GNDA.t30 29.5024
R4564 GNDA.n187 GNDA.n186 28.413
R4565 GNDA.n2370 GNDA.n2361 28.413
R4566 GNDA.n2308 GNDA.n232 28.1318
R4567 GNDA.t328 GNDA.n241 28.1074
R4568 GNDA.n181 GNDA.n113 28.038
R4569 GNDA.n2377 GNDA.n2376 28.038
R4570 GNDA.n251 GNDA.t80 27.9177
R4571 GNDA.n1436 GNDA.n1435 27.8193
R4572 GNDA.n1475 GNDA.n1474 27.8193
R4573 GNDA.n1267 GNDA.n1247 27.5561
R4574 GNDA.n1105 GNDA.n1085 27.5561
R4575 GNDA.n935 GNDA.n934 27.5561
R4576 GNDA.n1619 GNDA.n1502 27.5561
R4577 GNDA.n400 GNDA.n399 27.5561
R4578 GNDA.n1805 GNDA.n1013 27.5561
R4579 GNDA.n635 GNDA.n512 27.5561
R4580 GNDA.n2029 GNDA.n2009 27.5561
R4581 GNDA.n790 GNDA.n739 27.5561
R4582 GNDA.t224 GNDA.n287 26.4365
R4583 GNDA.n192 GNDA.t42 25.6905
R4584 GNDA.n2358 GNDA.t9 25.6905
R4585 GNDA.n140 GNDA.n139 25.6005
R4586 GNDA.n2368 GNDA.n2367 25.6005
R4587 GNDA.n1432 GNDA.n1431 25.2879
R4588 GNDA.n1471 GNDA.n1470 25.2879
R4589 GNDA.n1462 GNDA.t143 24.0005
R4590 GNDA.n1462 GNDA.t49 24.0005
R4591 GNDA.n1460 GNDA.t149 24.0005
R4592 GNDA.n1460 GNDA.t155 24.0005
R4593 GNDA.n1458 GNDA.t137 24.0005
R4594 GNDA.n1458 GNDA.t38 24.0005
R4595 GNDA.n1456 GNDA.t70 24.0005
R4596 GNDA.n1456 GNDA.t147 24.0005
R4597 GNDA.n1454 GNDA.t145 24.0005
R4598 GNDA.n1454 GNDA.t133 24.0005
R4599 GNDA.n1452 GNDA.t141 24.0005
R4600 GNDA.n1452 GNDA.t68 24.0005
R4601 GNDA.n1450 GNDA.t332 24.0005
R4602 GNDA.n1450 GNDA.t153 24.0005
R4603 GNDA.n1448 GNDA.t183 24.0005
R4604 GNDA.n1448 GNDA.t135 24.0005
R4605 GNDA.n1446 GNDA.t139 24.0005
R4606 GNDA.n1446 GNDA.t40 24.0005
R4607 GNDA.n1445 GNDA.t185 24.0005
R4608 GNDA.n1445 GNDA.t151 24.0005
R4609 GNDA.n1243 GNDA.n1242 23.6449
R4610 GNDA.n1081 GNDA.n1080 23.6449
R4611 GNDA.n952 GNDA.n951 23.6449
R4612 GNDA.n1498 GNDA.n1497 23.6449
R4613 GNDA.n417 GNDA.n416 23.6449
R4614 GNDA.n1009 GNDA.n1008 23.6449
R4615 GNDA.n508 GNDA.n507 23.6449
R4616 GNDA.n2005 GNDA.n2004 23.6449
R4617 GNDA.n735 GNDA.n734 23.6449
R4618 GNDA.n2287 GNDA.t85 22.997
R4619 GNDA.t224 GNDA.n308 22.7597
R4620 GNDA.n149 GNDA.n35 22.4005
R4621 GNDA.n2416 GNDA.n34 22.4005
R4622 GNDA.n2397 GNDA.n2396 22.4005
R4623 GNDA.n2398 GNDA.n2397 22.4005
R4624 GNDA.n205 GNDA.n113 22.4005
R4625 GNDA.n2376 GNDA.n2375 22.4005
R4626 GNDA GNDA.n2426 22.3396
R4627 GNDA.n2310 GNDA.n2309 21.4917
R4628 GNDA.n55 GNDA.n51 21.3338
R4629 GNDA.n53 GNDA.n52 21.3338
R4630 GNDA.n65 GNDA.n64 21.3338
R4631 GNDA.n71 GNDA.n70 21.3338
R4632 GNDA.n72 GNDA.n69 21.3338
R4633 GNDA.n76 GNDA.n68 21.3338
R4634 GNDA.n77 GNDA.n67 21.3338
R4635 GNDA.n78 GNDA.n66 21.3338
R4636 GNDA.n2399 GNDA.n2391 21.3338
R4637 GNDA.n2398 GNDA.n2392 21.3338
R4638 GNDA.n2396 GNDA.n2393 21.3338
R4639 GNDA.n2395 GNDA.n2394 21.3338
R4640 GNDA.n126 GNDA.n125 21.3338
R4641 GNDA.n131 GNDA.n129 21.3338
R4642 GNDA.n137 GNDA.n136 21.3338
R4643 GNDA.n141 GNDA.n138 21.3338
R4644 GNDA.n1412 GNDA.n1411 21.3338
R4645 GNDA.n1415 GNDA.n1414 21.3338
R4646 GNDA.n1476 GNDA.n1410 21.3338
R4647 GNDA.n1409 GNDA.n1408 21.3338
R4648 GNDA.n1444 GNDA.n1443 21.3338
R4649 GNDA.n1439 GNDA.n1438 21.3338
R4650 GNDA.n2364 GNDA.n2362 21.3338
R4651 GNDA.n98 GNDA.n97 21.3338
R4652 GNDA.n86 GNDA.n85 21.3338
R4653 GNDA.n84 GNDA.n83 21.3338
R4654 GNDA.n1466 GNDA.n1465 21.1792
R4655 GNDA.t159 GNDA.n2387 21.0733
R4656 GNDA.n197 GNDA.n196 20.6005
R4657 GNDA.n2355 GNDA.n2354 20.6005
R4658 GNDA.n2286 GNDA.n255 20.4418
R4659 GNDA.n2294 GNDA.n2293 20.4418
R4660 GNDA.n21 GNDA.t123 19.7005
R4661 GNDA.n21 GNDA.t194 19.7005
R4662 GNDA.n19 GNDA.t20 19.7005
R4663 GNDA.n19 GNDA.t176 19.7005
R4664 GNDA.n17 GNDA.t88 19.7005
R4665 GNDA.n17 GNDA.t76 19.7005
R4666 GNDA.n15 GNDA.t15 19.7005
R4667 GNDA.n15 GNDA.t89 19.7005
R4668 GNDA.n13 GNDA.t43 19.7005
R4669 GNDA.n13 GNDA.t14 19.7005
R4670 GNDA.n12 GNDA.t192 19.7005
R4671 GNDA.n12 GNDA.t96 19.7005
R4672 GNDA.n10 GNDA.t193 19.7005
R4673 GNDA.n10 GNDA.t347 19.7005
R4674 GNDA.n8 GNDA.t336 19.7005
R4675 GNDA.n8 GNDA.t109 19.7005
R4676 GNDA.n6 GNDA.t345 19.7005
R4677 GNDA.n6 GNDA.t75 19.7005
R4678 GNDA.n4 GNDA.t163 19.7005
R4679 GNDA.n4 GNDA.t56 19.7005
R4680 GNDA.n2 GNDA.t180 19.7005
R4681 GNDA.n2 GNDA.t71 19.7005
R4682 GNDA.n1 GNDA.t340 19.7005
R4683 GNDA.n1 GNDA.t196 19.7005
R4684 GNDA.n2314 GNDA.n2313 19.4279
R4685 GNDA.n2403 GNDA.n2402 19.288
R4686 GNDA.n2291 GNDA.n253 19.2005
R4687 GNDA.n2284 GNDA.n2283 19.2005
R4688 GNDA.n2317 GNDA.n218 19.2005
R4689 GNDA.n2309 GNDA.n229 19.2005
R4690 GNDA.n2299 GNDA.n233 19.2005
R4691 GNDA.n1392 GNDA.n226 19.2005
R4692 GNDA.n139 GNDA.n127 19.1005
R4693 GNDA.n2369 GNDA.n2368 19.1005
R4694 GNDA.t134 GNDA.t186 18.966
R4695 GNDA.t136 GNDA.t90 18.966
R4696 GNDA.n118 GNDA.n117 18.6842
R4697 GNDA.n2346 GNDA.n2344 18.6842
R4698 GNDA.n2319 GNDA.n226 17.613
R4699 GNDA.n2120 GNDA.n228 17.4917
R4700 GNDA.n2127 GNDA.n2126 16.9605
R4701 GNDA.n1354 GNDA.n1199 16.9379
R4702 GNDA.n1545 GNDA.n1544 16.9379
R4703 GNDA.n557 GNDA.n556 16.9379
R4704 GNDA.t166 GNDA.n37 16.9236
R4705 GNDA.t126 GNDA.n28 16.9236
R4706 GNDA.t57 GNDA.n29 16.9236
R4707 GNDA.t287 GNDA.t344 16.8587
R4708 GNDA.t65 GNDA.t348 16.8587
R4709 GNDA.t23 GNDA.t322 16.8587
R4710 GNDA.t314 GNDA.t7 16.8587
R4711 GNDA.t44 GNDA.t315 16.8587
R4712 GNDA.t166 GNDA.t325 16.8587
R4713 GNDA.t32 GNDA.t27 16.8587
R4714 GNDA.t46 GNDA.t158 16.8587
R4715 GNDA.t293 GNDA.t73 16.8587
R4716 GNDA.t321 GNDA.t181 16.8587
R4717 GNDA.t125 GNDA.t59 16.8587
R4718 GNDA.t0 GNDA.t126 16.8587
R4719 GNDA.t2 GNDA.t131 16.8587
R4720 GNDA.t127 GNDA.t316 16.8587
R4721 GNDA.t84 GNDA.t57 16.8587
R4722 GNDA.t8 GNDA.t94 16.8587
R4723 GNDA.t177 GNDA.t308 16.8587
R4724 GNDA.n1267 GNDA.n1266 16.0005
R4725 GNDA.n1266 GNDA.n1265 16.0005
R4726 GNDA.n1265 GNDA.n1249 16.0005
R4727 GNDA.n1259 GNDA.n1249 16.0005
R4728 GNDA.n1259 GNDA.n1258 16.0005
R4729 GNDA.n1258 GNDA.n1257 16.0005
R4730 GNDA.n1257 GNDA.n1251 16.0005
R4731 GNDA.n1252 GNDA.n1251 16.0005
R4732 GNDA.n1273 GNDA.n1247 16.0005
R4733 GNDA.n1274 GNDA.n1273 16.0005
R4734 GNDA.n1275 GNDA.n1274 16.0005
R4735 GNDA.n1275 GNDA.n1245 16.0005
R4736 GNDA.n1281 GNDA.n1245 16.0005
R4737 GNDA.n1282 GNDA.n1281 16.0005
R4738 GNDA.n1283 GNDA.n1282 16.0005
R4739 GNDA.n1283 GNDA.n1243 16.0005
R4740 GNDA.n1290 GNDA.n1242 16.0005
R4741 GNDA.n1291 GNDA.n1290 16.0005
R4742 GNDA.n1292 GNDA.n1291 16.0005
R4743 GNDA.n1292 GNDA.n1240 16.0005
R4744 GNDA.n1299 GNDA.n1298 16.0005
R4745 GNDA.n1300 GNDA.n1299 16.0005
R4746 GNDA.n1300 GNDA.n1238 16.0005
R4747 GNDA.n1105 GNDA.n1104 16.0005
R4748 GNDA.n1104 GNDA.n1103 16.0005
R4749 GNDA.n1103 GNDA.n1087 16.0005
R4750 GNDA.n1097 GNDA.n1087 16.0005
R4751 GNDA.n1097 GNDA.n1096 16.0005
R4752 GNDA.n1096 GNDA.n1095 16.0005
R4753 GNDA.n1095 GNDA.n1089 16.0005
R4754 GNDA.n1090 GNDA.n1089 16.0005
R4755 GNDA.n1111 GNDA.n1085 16.0005
R4756 GNDA.n1112 GNDA.n1111 16.0005
R4757 GNDA.n1113 GNDA.n1112 16.0005
R4758 GNDA.n1113 GNDA.n1083 16.0005
R4759 GNDA.n1119 GNDA.n1083 16.0005
R4760 GNDA.n1120 GNDA.n1119 16.0005
R4761 GNDA.n1121 GNDA.n1120 16.0005
R4762 GNDA.n1121 GNDA.n1081 16.0005
R4763 GNDA.n1128 GNDA.n1080 16.0005
R4764 GNDA.n1129 GNDA.n1128 16.0005
R4765 GNDA.n1130 GNDA.n1129 16.0005
R4766 GNDA.n1130 GNDA.n1078 16.0005
R4767 GNDA.n1137 GNDA.n1136 16.0005
R4768 GNDA.n1138 GNDA.n1137 16.0005
R4769 GNDA.n1138 GNDA.n1076 16.0005
R4770 GNDA.n934 GNDA.n880 16.0005
R4771 GNDA.n928 GNDA.n880 16.0005
R4772 GNDA.n928 GNDA.n927 16.0005
R4773 GNDA.n927 GNDA.n926 16.0005
R4774 GNDA.n926 GNDA.n882 16.0005
R4775 GNDA.n920 GNDA.n882 16.0005
R4776 GNDA.n920 GNDA.n919 16.0005
R4777 GNDA.n919 GNDA.n918 16.0005
R4778 GNDA.n936 GNDA.n935 16.0005
R4779 GNDA.n936 GNDA.n878 16.0005
R4780 GNDA.n942 GNDA.n878 16.0005
R4781 GNDA.n943 GNDA.n942 16.0005
R4782 GNDA.n944 GNDA.n943 16.0005
R4783 GNDA.n944 GNDA.n876 16.0005
R4784 GNDA.n950 GNDA.n876 16.0005
R4785 GNDA.n951 GNDA.n950 16.0005
R4786 GNDA.n952 GNDA.n874 16.0005
R4787 GNDA.n874 GNDA.n873 16.0005
R4788 GNDA.n959 GNDA.n873 16.0005
R4789 GNDA.n960 GNDA.n959 16.0005
R4790 GNDA.n961 GNDA.n871 16.0005
R4791 GNDA.n871 GNDA.n869 16.0005
R4792 GNDA.n968 GNDA.n869 16.0005
R4793 GNDA.n2120 GNDA.n2119 16.0005
R4794 GNDA.n2126 GNDA.n2119 16.0005
R4795 GNDA.n1619 GNDA.n1618 16.0005
R4796 GNDA.n1618 GNDA.n1617 16.0005
R4797 GNDA.n1617 GNDA.n1504 16.0005
R4798 GNDA.n1611 GNDA.n1504 16.0005
R4799 GNDA.n1611 GNDA.n1610 16.0005
R4800 GNDA.n1610 GNDA.n1609 16.0005
R4801 GNDA.n1609 GNDA.n1506 16.0005
R4802 GNDA.n1507 GNDA.n1506 16.0005
R4803 GNDA.n1625 GNDA.n1502 16.0005
R4804 GNDA.n1626 GNDA.n1625 16.0005
R4805 GNDA.n1627 GNDA.n1626 16.0005
R4806 GNDA.n1627 GNDA.n1500 16.0005
R4807 GNDA.n1633 GNDA.n1500 16.0005
R4808 GNDA.n1634 GNDA.n1633 16.0005
R4809 GNDA.n1635 GNDA.n1634 16.0005
R4810 GNDA.n1635 GNDA.n1498 16.0005
R4811 GNDA.n1642 GNDA.n1497 16.0005
R4812 GNDA.n1643 GNDA.n1642 16.0005
R4813 GNDA.n1644 GNDA.n1643 16.0005
R4814 GNDA.n1644 GNDA.n1495 16.0005
R4815 GNDA.n1651 GNDA.n1650 16.0005
R4816 GNDA.n1652 GNDA.n1651 16.0005
R4817 GNDA.n1652 GNDA.n1493 16.0005
R4818 GNDA.n399 GNDA.n375 16.0005
R4819 GNDA.n393 GNDA.n375 16.0005
R4820 GNDA.n393 GNDA.n392 16.0005
R4821 GNDA.n392 GNDA.n391 16.0005
R4822 GNDA.n391 GNDA.n377 16.0005
R4823 GNDA.n385 GNDA.n377 16.0005
R4824 GNDA.n385 GNDA.n384 16.0005
R4825 GNDA.n384 GNDA.n383 16.0005
R4826 GNDA.n401 GNDA.n400 16.0005
R4827 GNDA.n401 GNDA.n373 16.0005
R4828 GNDA.n407 GNDA.n373 16.0005
R4829 GNDA.n408 GNDA.n407 16.0005
R4830 GNDA.n409 GNDA.n408 16.0005
R4831 GNDA.n409 GNDA.n371 16.0005
R4832 GNDA.n415 GNDA.n371 16.0005
R4833 GNDA.n416 GNDA.n415 16.0005
R4834 GNDA.n417 GNDA.n369 16.0005
R4835 GNDA.n369 GNDA.n368 16.0005
R4836 GNDA.n424 GNDA.n368 16.0005
R4837 GNDA.n425 GNDA.n424 16.0005
R4838 GNDA.n426 GNDA.n366 16.0005
R4839 GNDA.n366 GNDA.n363 16.0005
R4840 GNDA.n433 GNDA.n363 16.0005
R4841 GNDA.n1805 GNDA.n1804 16.0005
R4842 GNDA.n1804 GNDA.n1803 16.0005
R4843 GNDA.n1803 GNDA.n1015 16.0005
R4844 GNDA.n1797 GNDA.n1015 16.0005
R4845 GNDA.n1797 GNDA.n1796 16.0005
R4846 GNDA.n1796 GNDA.n1795 16.0005
R4847 GNDA.n1795 GNDA.n1017 16.0005
R4848 GNDA.n1018 GNDA.n1017 16.0005
R4849 GNDA.n1811 GNDA.n1013 16.0005
R4850 GNDA.n1812 GNDA.n1811 16.0005
R4851 GNDA.n1813 GNDA.n1812 16.0005
R4852 GNDA.n1813 GNDA.n1011 16.0005
R4853 GNDA.n1819 GNDA.n1011 16.0005
R4854 GNDA.n1820 GNDA.n1819 16.0005
R4855 GNDA.n1821 GNDA.n1820 16.0005
R4856 GNDA.n1821 GNDA.n1009 16.0005
R4857 GNDA.n1828 GNDA.n1008 16.0005
R4858 GNDA.n1829 GNDA.n1828 16.0005
R4859 GNDA.n1830 GNDA.n1829 16.0005
R4860 GNDA.n1830 GNDA.n1006 16.0005
R4861 GNDA.n1837 GNDA.n1836 16.0005
R4862 GNDA.n1838 GNDA.n1837 16.0005
R4863 GNDA.n1838 GNDA.n1004 16.0005
R4864 GNDA.n635 GNDA.n634 16.0005
R4865 GNDA.n634 GNDA.n633 16.0005
R4866 GNDA.n633 GNDA.n514 16.0005
R4867 GNDA.n627 GNDA.n514 16.0005
R4868 GNDA.n627 GNDA.n626 16.0005
R4869 GNDA.n626 GNDA.n625 16.0005
R4870 GNDA.n625 GNDA.n516 16.0005
R4871 GNDA.n517 GNDA.n516 16.0005
R4872 GNDA.n641 GNDA.n512 16.0005
R4873 GNDA.n642 GNDA.n641 16.0005
R4874 GNDA.n643 GNDA.n642 16.0005
R4875 GNDA.n643 GNDA.n510 16.0005
R4876 GNDA.n649 GNDA.n510 16.0005
R4877 GNDA.n650 GNDA.n649 16.0005
R4878 GNDA.n651 GNDA.n650 16.0005
R4879 GNDA.n651 GNDA.n508 16.0005
R4880 GNDA.n658 GNDA.n507 16.0005
R4881 GNDA.n659 GNDA.n658 16.0005
R4882 GNDA.n660 GNDA.n659 16.0005
R4883 GNDA.n660 GNDA.n505 16.0005
R4884 GNDA.n667 GNDA.n666 16.0005
R4885 GNDA.n668 GNDA.n667 16.0005
R4886 GNDA.n668 GNDA.n503 16.0005
R4887 GNDA.n2029 GNDA.n2028 16.0005
R4888 GNDA.n2028 GNDA.n2027 16.0005
R4889 GNDA.n2027 GNDA.n2011 16.0005
R4890 GNDA.n2021 GNDA.n2011 16.0005
R4891 GNDA.n2021 GNDA.n2020 16.0005
R4892 GNDA.n2020 GNDA.n2019 16.0005
R4893 GNDA.n2019 GNDA.n2013 16.0005
R4894 GNDA.n2014 GNDA.n2013 16.0005
R4895 GNDA.n2035 GNDA.n2009 16.0005
R4896 GNDA.n2036 GNDA.n2035 16.0005
R4897 GNDA.n2037 GNDA.n2036 16.0005
R4898 GNDA.n2037 GNDA.n2007 16.0005
R4899 GNDA.n2043 GNDA.n2007 16.0005
R4900 GNDA.n2044 GNDA.n2043 16.0005
R4901 GNDA.n2045 GNDA.n2044 16.0005
R4902 GNDA.n2045 GNDA.n2005 16.0005
R4903 GNDA.n2052 GNDA.n2004 16.0005
R4904 GNDA.n2053 GNDA.n2052 16.0005
R4905 GNDA.n2054 GNDA.n2053 16.0005
R4906 GNDA.n2054 GNDA.n2002 16.0005
R4907 GNDA.n2061 GNDA.n2060 16.0005
R4908 GNDA.n2062 GNDA.n2061 16.0005
R4909 GNDA.n2062 GNDA.n2000 16.0005
R4910 GNDA.n790 GNDA.n789 16.0005
R4911 GNDA.n789 GNDA.n788 16.0005
R4912 GNDA.n788 GNDA.n741 16.0005
R4913 GNDA.n782 GNDA.n741 16.0005
R4914 GNDA.n782 GNDA.n781 16.0005
R4915 GNDA.n781 GNDA.n780 16.0005
R4916 GNDA.n780 GNDA.n743 16.0005
R4917 GNDA.n744 GNDA.n743 16.0005
R4918 GNDA.n796 GNDA.n739 16.0005
R4919 GNDA.n797 GNDA.n796 16.0005
R4920 GNDA.n798 GNDA.n797 16.0005
R4921 GNDA.n798 GNDA.n737 16.0005
R4922 GNDA.n804 GNDA.n737 16.0005
R4923 GNDA.n805 GNDA.n804 16.0005
R4924 GNDA.n806 GNDA.n805 16.0005
R4925 GNDA.n806 GNDA.n735 16.0005
R4926 GNDA.n813 GNDA.n734 16.0005
R4927 GNDA.n814 GNDA.n813 16.0005
R4928 GNDA.n815 GNDA.n814 16.0005
R4929 GNDA.n815 GNDA.n732 16.0005
R4930 GNDA.n822 GNDA.n821 16.0005
R4931 GNDA.n823 GNDA.n822 16.0005
R4932 GNDA.n823 GNDA.n730 16.0005
R4933 GNDA.t66 GNDA.t26 15.8816
R4934 GNDA.t107 GNDA.t72 15.8816
R4935 GNDA.n2322 GNDA.n2321 15.363
R4936 GNDA.n2321 GNDA.n223 15.363
R4937 GNDA GNDA.n2314 14.6989
R4938 GNDA.n2102 GNDA.n318 14.555
R4939 GNDA.n2207 GNDA.n317 14.555
R4940 GNDA.n180 GNDA.n179 14.0505
R4941 GNDA.n2382 GNDA.n2381 14.0505
R4942 GNDA.n1298 GNDA 14.0449
R4943 GNDA.n1136 GNDA 14.0449
R4944 GNDA.n961 GNDA 14.0449
R4945 GNDA.n1650 GNDA 14.0449
R4946 GNDA.n426 GNDA 14.0449
R4947 GNDA.n1836 GNDA 14.0449
R4948 GNDA.n666 GNDA 14.0449
R4949 GNDA.n2060 GNDA 14.0449
R4950 GNDA.n821 GNDA 14.0449
R4951 GNDA.n2424 GNDA.n2423 14.0193
R4952 GNDA.n2318 GNDA.n2317 13.8005
R4953 GNDA.n174 GNDA.n34 13.8005
R4954 GNDA.n149 GNDA.n148 13.8005
R4955 GNDA.n1465 GNDA.n228 13.7706
R4956 GNDA.n1694 GNDA.n1034 12.9309
R4957 GNDA.n1901 GNDA.n706 12.9309
R4958 GNDA.n2098 GNDA.n1947 12.9309
R4959 GNDA.n2203 GNDA.n457 12.9309
R4960 GNDA.n196 GNDA.n122 12.8005
R4961 GNDA.n2356 GNDA.n2355 12.8005
R4962 GNDA.t232 GNDA.n93 12.6442
R4963 GNDA.t346 GNDA.t279 12.6442
R4964 GNDA.t323 GNDA.t53 12.6442
R4965 GNDA.n2408 GNDA.t226 12.6442
R4966 GNDA.t78 GNDA.n2419 12.6442
R4967 GNDA.t168 GNDA.t22 12.6442
R4968 GNDA.t178 GNDA.t305 12.6442
R4969 GNDA.t236 GNDA.n183 12.6442
R4970 GNDA.n1873 GNDA.n1872 12.4126
R4971 GNDA.n970 GNDA.n289 12.4126
R4972 GNDA.n2268 GNDA.n282 12.4126
R4973 GNDA.n2110 GNDA.n2109 11.6369
R4974 GNDA.n2111 GNDA.n2110 11.6369
R4975 GNDA.n2111 GNDA.n472 11.6369
R4976 GNDA.n2117 GNDA.n472 11.6369
R4977 GNDA.n2118 GNDA.n2117 11.6369
R4978 GNDA.n2128 GNDA.n470 11.6369
R4979 GNDA.n470 GNDA.n469 11.6369
R4980 GNDA.n2135 GNDA.n469 11.6369
R4981 GNDA.n2136 GNDA.n2135 11.6369
R4982 GNDA.n2167 GNDA.n2136 11.6369
R4983 GNDA.n1894 GNDA.n1893 11.6369
R4984 GNDA.n1893 GNDA.n1892 11.6369
R4985 GNDA.n1892 GNDA.n856 11.6369
R4986 GNDA.n1886 GNDA.n856 11.6369
R4987 GNDA.n1886 GNDA.n1885 11.6369
R4988 GNDA.n1885 GNDA.n1884 11.6369
R4989 GNDA.n1884 GNDA.n862 11.6369
R4990 GNDA.n997 GNDA.n862 11.6369
R4991 GNDA.n1877 GNDA.n997 11.6369
R4992 GNDA.n1877 GNDA.n1876 11.6369
R4993 GNDA.n1876 GNDA.n1875 11.6369
R4994 GNDA.n1872 GNDA.n1871 11.6369
R4995 GNDA.n1871 GNDA.n1869 11.6369
R4996 GNDA.n1869 GNDA.n1866 11.6369
R4997 GNDA.n1866 GNDA.n1865 11.6369
R4998 GNDA.n1865 GNDA.n1862 11.6369
R4999 GNDA.n1862 GNDA.n1861 11.6369
R5000 GNDA.n1858 GNDA.n1857 11.6369
R5001 GNDA.n1857 GNDA.n1854 11.6369
R5002 GNDA.n1355 GNDA.n1354 11.6369
R5003 GNDA.n1356 GNDA.n1355 11.6369
R5004 GNDA.n1356 GNDA.n1197 11.6369
R5005 GNDA.n1362 GNDA.n1197 11.6369
R5006 GNDA.n1363 GNDA.n1362 11.6369
R5007 GNDA.n1364 GNDA.n1363 11.6369
R5008 GNDA.n1364 GNDA.n1195 11.6369
R5009 GNDA.n1370 GNDA.n1195 11.6369
R5010 GNDA.n1371 GNDA.n1370 11.6369
R5011 GNDA.n1372 GNDA.n1371 11.6369
R5012 GNDA.n1372 GNDA.n680 11.6369
R5013 GNDA.n1348 GNDA.n1199 11.6369
R5014 GNDA.n1348 GNDA.n1347 11.6369
R5015 GNDA.n1347 GNDA.n1346 11.6369
R5016 GNDA.n1346 GNDA.n1201 11.6369
R5017 GNDA.n1341 GNDA.n1201 11.6369
R5018 GNDA.n1341 GNDA.n1340 11.6369
R5019 GNDA.n1340 GNDA.n1339 11.6369
R5020 GNDA.n1339 GNDA.n1204 11.6369
R5021 GNDA.n1334 GNDA.n1204 11.6369
R5022 GNDA.n1544 GNDA.n1543 11.6369
R5023 GNDA.n1543 GNDA.n1520 11.6369
R5024 GNDA.n1538 GNDA.n1520 11.6369
R5025 GNDA.n1538 GNDA.n1537 11.6369
R5026 GNDA.n1537 GNDA.n1536 11.6369
R5027 GNDA.n1536 GNDA.n1523 11.6369
R5028 GNDA.n1531 GNDA.n1523 11.6369
R5029 GNDA.n1531 GNDA.n1530 11.6369
R5030 GNDA.n1530 GNDA.n1529 11.6369
R5031 GNDA.n1529 GNDA.n1036 11.6369
R5032 GNDA.n1693 GNDA.n1036 11.6369
R5033 GNDA.n1545 GNDA.n1518 11.6369
R5034 GNDA.n1551 GNDA.n1518 11.6369
R5035 GNDA.n1552 GNDA.n1551 11.6369
R5036 GNDA.n1553 GNDA.n1552 11.6369
R5037 GNDA.n1553 GNDA.n1516 11.6369
R5038 GNDA.n1559 GNDA.n1516 11.6369
R5039 GNDA.n1560 GNDA.n1559 11.6369
R5040 GNDA.n1561 GNDA.n1560 11.6369
R5041 GNDA.n1561 GNDA.n1514 11.6369
R5042 GNDA.n1699 GNDA.n1695 11.6369
R5043 GNDA.n1700 GNDA.n1699 11.6369
R5044 GNDA.n1701 GNDA.n1700 11.6369
R5045 GNDA.n1701 GNDA.n1032 11.6369
R5046 GNDA.n1707 GNDA.n1032 11.6369
R5047 GNDA.n1708 GNDA.n1707 11.6369
R5048 GNDA.n1709 GNDA.n1708 11.6369
R5049 GNDA.n1709 GNDA.n1030 11.6369
R5050 GNDA.n1715 GNDA.n1030 11.6369
R5051 GNDA.n1716 GNDA.n1715 11.6369
R5052 GNDA.n1717 GNDA.n1716 11.6369
R5053 GNDA.n1946 GNDA.n682 11.6369
R5054 GNDA.n1940 GNDA.n682 11.6369
R5055 GNDA.n1940 GNDA.n1939 11.6369
R5056 GNDA.n1939 GNDA.n1938 11.6369
R5057 GNDA.n1938 GNDA.n1936 11.6369
R5058 GNDA.n1936 GNDA.n1933 11.6369
R5059 GNDA.n1933 GNDA.n1932 11.6369
R5060 GNDA.n1932 GNDA.n1929 11.6369
R5061 GNDA.n1929 GNDA.n1928 11.6369
R5062 GNDA.n1928 GNDA.n1925 11.6369
R5063 GNDA.n1925 GNDA.n1924 11.6369
R5064 GNDA.n850 GNDA.n849 11.6369
R5065 GNDA.n849 GNDA.n848 11.6369
R5066 GNDA.n848 GNDA.n715 11.6369
R5067 GNDA.n842 GNDA.n715 11.6369
R5068 GNDA.n842 GNDA.n841 11.6369
R5069 GNDA.n841 GNDA.n840 11.6369
R5070 GNDA.n840 GNDA.n721 11.6369
R5071 GNDA.n831 GNDA.n721 11.6369
R5072 GNDA.n833 GNDA.n831 11.6369
R5073 GNDA.n833 GNDA.n832 11.6369
R5074 GNDA.n832 GNDA.n291 11.6369
R5075 GNDA.n972 GNDA.n970 11.6369
R5076 GNDA.n973 GNDA.n972 11.6369
R5077 GNDA.n976 GNDA.n973 11.6369
R5078 GNDA.n977 GNDA.n976 11.6369
R5079 GNDA.n980 GNDA.n977 11.6369
R5080 GNDA.n981 GNDA.n980 11.6369
R5081 GNDA.n985 GNDA.n984 11.6369
R5082 GNDA.n988 GNDA.n985 11.6369
R5083 GNDA.n556 GNDA.n555 11.6369
R5084 GNDA.n555 GNDA.n528 11.6369
R5085 GNDA.n550 GNDA.n528 11.6369
R5086 GNDA.n550 GNDA.n549 11.6369
R5087 GNDA.n549 GNDA.n530 11.6369
R5088 GNDA.n544 GNDA.n530 11.6369
R5089 GNDA.n544 GNDA.n543 11.6369
R5090 GNDA.n543 GNDA.n542 11.6369
R5091 GNDA.n542 GNDA.n532 11.6369
R5092 GNDA.n536 GNDA.n532 11.6369
R5093 GNDA.n536 GNDA.n535 11.6369
R5094 GNDA.n557 GNDA.n526 11.6369
R5095 GNDA.n563 GNDA.n526 11.6369
R5096 GNDA.n564 GNDA.n563 11.6369
R5097 GNDA.n565 GNDA.n564 11.6369
R5098 GNDA.n565 GNDA.n524 11.6369
R5099 GNDA.n571 GNDA.n524 11.6369
R5100 GNDA.n572 GNDA.n571 11.6369
R5101 GNDA.n573 GNDA.n572 11.6369
R5102 GNDA.n573 GNDA.n522 11.6369
R5103 GNDA.n2268 GNDA.n2267 11.6369
R5104 GNDA.n2267 GNDA.n2266 11.6369
R5105 GNDA.n2266 GNDA.n2265 11.6369
R5106 GNDA.n2265 GNDA.n2263 11.6369
R5107 GNDA.n2263 GNDA.n2260 11.6369
R5108 GNDA.n2260 GNDA.n2259 11.6369
R5109 GNDA.n2256 GNDA.n2255 11.6369
R5110 GNDA.n2255 GNDA.n2252 11.6369
R5111 GNDA.n2165 GNDA.n2164 11.6369
R5112 GNDA.n2164 GNDA.n2137 11.6369
R5113 GNDA.n2158 GNDA.n2137 11.6369
R5114 GNDA.n2158 GNDA.n2157 11.6369
R5115 GNDA.n2157 GNDA.n2156 11.6369
R5116 GNDA.n2156 GNDA.n2139 11.6369
R5117 GNDA.n2150 GNDA.n2139 11.6369
R5118 GNDA.n2150 GNDA.n2149 11.6369
R5119 GNDA.n2149 GNDA.n2148 11.6369
R5120 GNDA.n2148 GNDA.n2141 11.6369
R5121 GNDA.n2142 GNDA.n2141 11.6369
R5122 GNDA.n1858 GNDA 11.5076
R5123 GNDA.n984 GNDA 11.5076
R5124 GNDA.n2256 GNDA 11.5076
R5125 GNDA.n1854 GNDA.n1853 11.4026
R5126 GNDA.n989 GNDA.n988 11.4026
R5127 GNDA.n2252 GNDA.n2251 11.4026
R5128 GNDA.n2295 GNDA.n2294 11.381
R5129 GNDA.n1334 GNDA.n1333 11.249
R5130 GNDA.n1567 GNDA.n1514 11.249
R5131 GNDA.n579 GNDA.n522 11.249
R5132 GNDA.n2127 GNDA.n2118 10.4732
R5133 GNDA.n2320 GNDA.n224 9.78488
R5134 GNDA.n2296 GNDA.t102 9.71084
R5135 GNDA.n150 GNDA.t267 9.6005
R5136 GNDA.n150 GNDA.t334 9.6005
R5137 GNDA.n152 GNDA.t25 9.6005
R5138 GNDA.n152 GNDA.t116 9.6005
R5139 GNDA.n154 GNDA.t17 9.6005
R5140 GNDA.n154 GNDA.t61 9.6005
R5141 GNDA.n156 GNDA.t19 9.6005
R5142 GNDA.n156 GNDA.t118 9.6005
R5143 GNDA.n158 GNDA.t36 9.6005
R5144 GNDA.n158 GNDA.t98 9.6005
R5145 GNDA.n160 GNDA.t324 9.6005
R5146 GNDA.n160 GNDA.t6 9.6005
R5147 GNDA.n162 GNDA.t114 9.6005
R5148 GNDA.n162 GNDA.t100 9.6005
R5149 GNDA.n164 GNDA.t4 9.6005
R5150 GNDA.n164 GNDA.t63 9.6005
R5151 GNDA.n166 GNDA.t342 9.6005
R5152 GNDA.n166 GNDA.t327 9.6005
R5153 GNDA.n168 GNDA.t92 9.6005
R5154 GNDA.n168 GNDA.t157 9.6005
R5155 GNDA.n170 GNDA.t120 9.6005
R5156 GNDA.n170 GNDA.t111 9.6005
R5157 GNDA.n172 GNDA.t52 9.6005
R5158 GNDA.n172 GNDA.t253 9.6005
R5159 GNDA.n2316 GNDA.t195 9.6005
R5160 GNDA.n2316 GNDA.t198 9.6005
R5161 GNDA.n225 GNDA.t191 9.6005
R5162 GNDA.n225 GNDA.t199 9.6005
R5163 GNDA.n57 GNDA.n50 9.5505
R5164 GNDA.n2318 GNDA.n2315 9.37925
R5165 GNDA.n2339 GNDA.n106 9.10395
R5166 GNDA.n175 GNDA.n174 9.0005
R5167 GNDA.n148 GNDA.n0 8.96925
R5168 GNDA.n1875 GNDA.n1873 8.66313
R5169 GNDA.n291 GNDA.n289 8.66313
R5170 GNDA.n2142 GNDA.n282 8.66313
R5171 GNDA.n1377 GNDA.n318 8.60107
R5172 GNDA.n690 GNDA.n317 8.60107
R5173 GNDA.n2167 GNDA.n2166 8.53383
R5174 GNDA.n1947 GNDA.n680 8.53383
R5175 GNDA.n1694 GNDA.n1693 8.53383
R5176 GNDA.n1717 GNDA.n706 8.53383
R5177 GNDA.n1924 GNDA.n457 8.53383
R5178 GNDA.n535 GNDA.n474 8.53383
R5179 GNDA.n2296 GNDA.t105 8.49705
R5180 GNDA.n1464 GNDA.n1463 8.44175
R5181 GNDA.n2405 GNDA.t11 8.42962
R5182 GNDA.n1252 GNDA.n1208 8.35606
R5183 GNDA.n1090 GNDA.n1048 8.35606
R5184 GNDA.n918 GNDA.n884 8.35606
R5185 GNDA.n1568 GNDA.n1507 8.35606
R5186 GNDA.n383 GNDA.n380 8.35606
R5187 GNDA.n1752 GNDA.n1018 8.35606
R5188 GNDA.n580 GNDA.n517 8.35606
R5189 GNDA.n2014 GNDA.n1973 8.35606
R5190 GNDA.n746 GNDA.n744 8.35606
R5191 GNDA.n2321 GNDA.n2320 7.71925
R5192 GNDA.n287 GNDA.n259 7.62664
R5193 GNDA.n118 GNDA.t337 7.00687
R5194 GNDA.n191 GNDA.t101 7.00687
R5195 GNDA.n2341 GNDA.t79 7.00687
R5196 GNDA.t64 GNDA.n2346 7.00687
R5197 GNDA.n2425 GNDA.n2424 6.7505
R5198 GNDA.n2424 GNDA.n23 6.688
R5199 GNDA.n177 GNDA.n175 6.563
R5200 GNDA.n2380 GNDA.n0 6.563
R5201 GNDA.n235 GNDA.n233 6.4005
R5202 GNDA.n1432 GNDA.t39 6.32234
R5203 GNDA.t284 GNDA.t21 6.32234
R5204 GNDA.n1480 GNDA.t67 6.32234
R5205 GNDA.n2325 GNDA.t144 6.32234
R5206 GNDA.t272 GNDA.t317 6.32234
R5207 GNDA.n1470 GNDA.t148 6.32234
R5208 GNDA.n175 GNDA.n23 5.03175
R5209 GNDA.n2295 GNDA.n240 4.8663
R5210 GNDA.n1666 GNDA.n1387 4.6085
R5211 GNDA.n2211 GNDA.n2210 4.6085
R5212 GNDA.n1851 GNDA.n1850 4.6085
R5213 GNDA.n1236 GNDA.n1233 4.6085
R5214 GNDA.n1074 GNDA.n1070 4.6085
R5215 GNDA.n991 GNDA.n990 4.6085
R5216 GNDA.n679 GNDA.n678 4.6085
R5217 GNDA.n1998 GNDA.n456 4.6085
R5218 GNDA.n2249 GNDA.n283 4.6085
R5219 GNDA.n1689 GNDA.n1035 4.55161
R5220 GNDA.n1721 GNDA.n1028 4.55161
R5221 GNDA.n1192 GNDA.n681 4.55161
R5222 GNDA.n1920 GNDA.n691 4.55161
R5223 GNDA.n2172 GNDA.n467 4.55161
R5224 GNDA.n2105 GNDA.n475 4.55161
R5225 GNDA.n1670 GNDA.n1668 4.5061
R5226 GNDA.n1023 GNDA.n434 4.5061
R5227 GNDA.n1232 GNDA.n1034 4.5061
R5228 GNDA.n1901 GNDA.n708 4.5061
R5229 GNDA.n2099 GNDA.n2098 4.5061
R5230 GNDA.n2204 GNDA.n2203 4.5061
R5231 GNDA.n50 GNDA.n48 4.5005
R5232 GNDA.n2320 GNDA.n2319 4.5005
R5233 GNDA.n2426 GNDA.n2425 4.5005
R5234 GNDA.n2109 GNDA.n474 4.39646
R5235 GNDA.n1894 GNDA.n706 4.39646
R5236 GNDA.n1695 GNDA.n1694 4.39646
R5237 GNDA.n1947 GNDA.n1946 4.39646
R5238 GNDA.n850 GNDA.n457 4.39646
R5239 GNDA.n2166 GNDA.n2165 4.39646
R5240 GNDA.n1670 GNDA.n1669 4.3525
R5241 GNDA.n1751 GNDA.n1023 4.3525
R5242 GNDA.n1171 GNDA.n1034 4.3525
R5243 GNDA.n1901 GNDA.n1900 4.3525
R5244 GNDA.n2098 GNDA.n2097 4.3525
R5245 GNDA.n2203 GNDA.n2202 4.3525
R5246 GNDA.n1669 GNDA.n340 4.3013
R5247 GNDA.n1753 GNDA.n1751 4.3013
R5248 GNDA.n1171 GNDA.n1170 4.3013
R5249 GNDA.n1900 GNDA.n709 4.3013
R5250 GNDA.n2097 GNDA.n2094 4.3013
R5251 GNDA.n2202 GNDA.n461 4.3013
R5252 GNDA.n1689 GNDA.n1688 4.26717
R5253 GNDA.n1688 GNDA.n1685 4.26717
R5254 GNDA.n1685 GNDA.n1684 4.26717
R5255 GNDA.n1684 GNDA.n1681 4.26717
R5256 GNDA.n1681 GNDA.n1680 4.26717
R5257 GNDA.n1680 GNDA.n1677 4.26717
R5258 GNDA.n1676 GNDA.n1673 4.26717
R5259 GNDA.n1673 GNDA.n1672 4.26717
R5260 GNDA.n1724 GNDA.n1721 4.26717
R5261 GNDA.n1727 GNDA.n1724 4.26717
R5262 GNDA.n1730 GNDA.n1727 4.26717
R5263 GNDA.n1730 GNDA.n1026 4.26717
R5264 GNDA.n1735 GNDA.n1026 4.26717
R5265 GNDA.n1738 GNDA.n1735 4.26717
R5266 GNDA.n1745 GNDA.n1742 4.26717
R5267 GNDA.n1747 GNDA.n1745 4.26717
R5268 GNDA.n1192 GNDA.n1191 4.26717
R5269 GNDA.n1191 GNDA.n1188 4.26717
R5270 GNDA.n1188 GNDA.n1187 4.26717
R5271 GNDA.n1187 GNDA.n1184 4.26717
R5272 GNDA.n1184 GNDA.n1183 4.26717
R5273 GNDA.n1183 GNDA.n1180 4.26717
R5274 GNDA.n1179 GNDA.n1176 4.26717
R5275 GNDA.n1176 GNDA.n1175 4.26717
R5276 GNDA.n1920 GNDA.n1919 4.26717
R5277 GNDA.n1919 GNDA.n1916 4.26717
R5278 GNDA.n1916 GNDA.n1915 4.26717
R5279 GNDA.n1915 GNDA.n1912 4.26717
R5280 GNDA.n1912 GNDA.n1911 4.26717
R5281 GNDA.n1911 GNDA.n1908 4.26717
R5282 GNDA.n1907 GNDA.n1904 4.26717
R5283 GNDA.n1904 GNDA.n1903 4.26717
R5284 GNDA.n2172 GNDA.n465 4.26717
R5285 GNDA.n2180 GNDA.n465 4.26717
R5286 GNDA.n2181 GNDA.n2180 4.26717
R5287 GNDA.n2184 GNDA.n2181 4.26717
R5288 GNDA.n2184 GNDA.n463 4.26717
R5289 GNDA.n2192 GNDA.n463 4.26717
R5290 GNDA.n2196 GNDA.n2193 4.26717
R5291 GNDA.n2196 GNDA.n459 4.26717
R5292 GNDA.n2105 GNDA.n476 4.26717
R5293 GNDA.n1951 GNDA.n476 4.26717
R5294 GNDA.n1952 GNDA.n1951 4.26717
R5295 GNDA.n1957 GNDA.n1952 4.26717
R5296 GNDA.n1958 GNDA.n1957 4.26717
R5297 GNDA.n1963 GNDA.n1958 4.26717
R5298 GNDA.n1969 GNDA.n1964 4.26717
R5299 GNDA.n1971 GNDA.n1969 4.26717
R5300 GNDA.n1333 GNDA.n1332 4.2501
R5301 GNDA.n581 GNDA.n579 4.2501
R5302 GNDA.t105 GNDA.t121 4.24878
R5303 GNDA GNDA.n1676 4.21976
R5304 GNDA.n1742 GNDA 4.21976
R5305 GNDA GNDA.n1179 4.21976
R5306 GNDA GNDA.n1907 4.21976
R5307 GNDA.n2193 GNDA 4.21976
R5308 GNDA.n1964 GNDA 4.21976
R5309 GNDA.t269 GNDA.t242 4.21506
R5310 GNDA.n2412 GNDA.t333 4.21506
R5311 GNDA.t339 GNDA.n2408 4.21506
R5312 GNDA.n2420 GNDA.t73 4.21506
R5313 GNDA.t221 GNDA.t229 4.21506
R5314 GNDA.n1569 GNDA.n1567 4.1477
R5315 GNDA.n1672 GNDA.n1670 4.12494
R5316 GNDA.n1747 GNDA.n1023 4.12494
R5317 GNDA.n1175 GNDA.n1034 4.12494
R5318 GNDA.n1903 GNDA.n1901 4.12494
R5319 GNDA.n2203 GNDA.n459 4.12494
R5320 GNDA.n2098 GNDA.n1971 4.12494
R5321 GNDA.n2271 GNDA.n259 4.08877
R5322 GNDA.n2319 GNDA.n2318 3.813
R5323 GNDA.n2315 GNDA 3.68412
R5324 GNDA.n1602 GNDA.n1509 3.5845
R5325 GNDA.n1601 GNDA.n1510 3.5845
R5326 GNDA.n1574 GNDA.n1573 3.5845
R5327 GNDA.n1595 GNDA.n1594 3.5845
R5328 GNDA.n1590 GNDA.n1575 3.5845
R5329 GNDA.n1589 GNDA.n1579 3.5845
R5330 GNDA.n1585 GNDA.n1584 3.5845
R5331 GNDA.n1580 GNDA.n1489 3.5845
R5332 GNDA.n1658 GNDA.n1657 3.5845
R5333 GNDA.n379 GNDA.n344 3.5845
R5334 GNDA.n2236 GNDA.n2235 3.5845
R5335 GNDA.n2231 GNDA.n345 3.5845
R5336 GNDA.n2230 GNDA.n348 3.5845
R5337 GNDA.n2226 GNDA.n2225 3.5845
R5338 GNDA.n352 GNDA.n350 3.5845
R5339 GNDA.n2220 GNDA.n354 3.5845
R5340 GNDA.n2219 GNDA.n355 3.5845
R5341 GNDA.n362 GNDA.n361 3.5845
R5342 GNDA.n1788 GNDA.n1020 3.5845
R5343 GNDA.n1787 GNDA.n1021 3.5845
R5344 GNDA.n1760 GNDA.n1759 3.5845
R5345 GNDA.n1781 GNDA.n1780 3.5845
R5346 GNDA.n1776 GNDA.n1761 3.5845
R5347 GNDA.n1775 GNDA.n1765 3.5845
R5348 GNDA.n1771 GNDA.n1770 3.5845
R5349 GNDA.n1766 GNDA.n1001 3.5845
R5350 GNDA.n1844 GNDA.n1843 3.5845
R5351 GNDA.n1328 GNDA.n1327 3.5845
R5352 GNDA.n1213 GNDA.n1211 3.5845
R5353 GNDA.n1322 GNDA.n1215 3.5845
R5354 GNDA.n1321 GNDA.n1216 3.5845
R5355 GNDA.n1317 GNDA.n1316 3.5845
R5356 GNDA.n1222 GNDA.n1220 3.5845
R5357 GNDA.n1311 GNDA.n1224 3.5845
R5358 GNDA.n1310 GNDA.n1225 3.5845
R5359 GNDA.n1306 GNDA.n1305 3.5845
R5360 GNDA.n1166 GNDA.n1165 3.5845
R5361 GNDA.n1052 GNDA.n1050 3.5845
R5362 GNDA.n1160 GNDA.n1054 3.5845
R5363 GNDA.n1159 GNDA.n1055 3.5845
R5364 GNDA.n1155 GNDA.n1154 3.5845
R5365 GNDA.n1061 GNDA.n1059 3.5845
R5366 GNDA.n1149 GNDA.n1063 3.5845
R5367 GNDA.n1148 GNDA.n1064 3.5845
R5368 GNDA.n1144 GNDA.n1143 3.5845
R5369 GNDA.n914 GNDA.n886 3.5845
R5370 GNDA.n913 GNDA.n912 3.5845
R5371 GNDA.n911 GNDA.n910 3.5845
R5372 GNDA.n889 GNDA.n887 3.5845
R5373 GNDA.n905 GNDA.n891 3.5845
R5374 GNDA.n904 GNDA.n901 3.5845
R5375 GNDA.n900 GNDA.n899 3.5845
R5376 GNDA.n895 GNDA.n892 3.5845
R5377 GNDA.n894 GNDA.n868 3.5845
R5378 GNDA.n618 GNDA.n519 3.5845
R5379 GNDA.n617 GNDA.n520 3.5845
R5380 GNDA.n613 GNDA.n612 3.5845
R5381 GNDA.n588 GNDA.n586 3.5845
R5382 GNDA.n607 GNDA.n590 3.5845
R5383 GNDA.n606 GNDA.n591 3.5845
R5384 GNDA.n602 GNDA.n601 3.5845
R5385 GNDA.n598 GNDA.n596 3.5845
R5386 GNDA.n673 GNDA.n501 3.5845
R5387 GNDA.n2090 GNDA.n2089 3.5845
R5388 GNDA.n1978 GNDA.n1976 3.5845
R5389 GNDA.n2084 GNDA.n1980 3.5845
R5390 GNDA.n2083 GNDA.n1981 3.5845
R5391 GNDA.n2079 GNDA.n2078 3.5845
R5392 GNDA.n1987 GNDA.n1985 3.5845
R5393 GNDA.n2073 GNDA.n1989 3.5845
R5394 GNDA.n2072 GNDA.n1990 3.5845
R5395 GNDA.n2068 GNDA.n2067 3.5845
R5396 GNDA.n773 GNDA.n748 3.5845
R5397 GNDA.n772 GNDA.n771 3.5845
R5398 GNDA.n770 GNDA.n769 3.5845
R5399 GNDA.n751 GNDA.n749 3.5845
R5400 GNDA.n764 GNDA.n753 3.5845
R5401 GNDA.n763 GNDA.n760 3.5845
R5402 GNDA.n759 GNDA.n758 3.5845
R5403 GNDA.n754 GNDA.n726 3.5845
R5404 GNDA.n829 GNDA.n828 3.5845
R5405 GNDA.n178 GNDA.t34 3.42907
R5406 GNDA.n178 GNDA.t31 3.42907
R5407 GNDA.n176 GNDA.t169 3.42907
R5408 GNDA.n176 GNDA.t172 3.42907
R5409 GNDA.n2379 GNDA.t83 3.42907
R5410 GNDA.n2379 GNDA.t54 3.42907
R5411 GNDA.n2378 GNDA.t330 3.42907
R5412 GNDA.n2378 GNDA.t29 3.42907
R5413 GNDA.n1569 GNDA.n1568 3.3797
R5414 GNDA.n380 GNDA.n340 3.3797
R5415 GNDA.n1753 GNDA.n1752 3.3797
R5416 GNDA.n1332 GNDA.n1208 3.3797
R5417 GNDA.n1170 GNDA.n1048 3.3797
R5418 GNDA.n884 GNDA.n709 3.3797
R5419 GNDA.n581 GNDA.n580 3.3797
R5420 GNDA.n2094 GNDA.n1973 3.3797
R5421 GNDA.n746 GNDA.n461 3.3797
R5422 GNDA.n247 GNDA.n232 3.2005
R5423 GNDA.n2299 GNDA.n2298 3.2005
R5424 GNDA.n1492 GNDA.n1490 2.8677
R5425 GNDA.n2213 GNDA.n2212 2.8677
R5426 GNDA.n1002 GNDA.n998 2.8677
R5427 GNDA.n1237 GNDA.n1229 2.8677
R5428 GNDA.n1075 GNDA.n1068 2.8677
R5429 GNDA.n993 GNDA.n992 2.8677
R5430 GNDA.n674 GNDA.n499 2.8677
R5431 GNDA.n1999 GNDA.n1994 2.8677
R5432 GNDA.n729 GNDA.n727 2.8677
R5433 GNDA.n2272 GNDA.t85 2.55567
R5434 GNDA.n255 GNDA.t328 2.55567
R5435 GNDA.n1451 GNDA.n1449 2.34425
R5436 GNDA.n1459 GNDA.n1457 2.34425
R5437 GNDA.t337 GNDA.n115 2.33596
R5438 GNDA.n201 GNDA.t104 2.33596
R5439 GNDA.t108 GNDA.n2350 2.33596
R5440 GNDA.n2347 GNDA.t64 2.33596
R5441 GNDA.n1238 GNDA.n1237 2.31161
R5442 GNDA.n1076 GNDA.n1075 2.31161
R5443 GNDA.n992 GNDA.n968 2.31161
R5444 GNDA.n1493 GNDA.n1492 2.31161
R5445 GNDA.n2212 GNDA.n433 2.31161
R5446 GNDA.n1004 GNDA.n998 2.31161
R5447 GNDA.n503 GNDA.n499 2.31161
R5448 GNDA.n2000 GNDA.n1999 2.31161
R5449 GNDA.n730 GNDA.n729 2.31161
R5450 GNDA.n1240 GNDA 1.95606
R5451 GNDA.n1078 GNDA 1.95606
R5452 GNDA GNDA.n960 1.95606
R5453 GNDA.n1495 GNDA 1.95606
R5454 GNDA GNDA.n425 1.95606
R5455 GNDA.n1006 GNDA 1.95606
R5456 GNDA.n505 GNDA 1.95606
R5457 GNDA.n2002 GNDA 1.95606
R5458 GNDA.n732 GNDA 1.95606
R5459 GNDA.n1492 GNDA.n1387 1.7413
R5460 GNDA.n2212 GNDA.n2211 1.7413
R5461 GNDA.n1850 GNDA.n998 1.7413
R5462 GNDA.n1237 GNDA.n1236 1.7413
R5463 GNDA.n1075 GNDA.n1074 1.7413
R5464 GNDA.n992 GNDA.n991 1.7413
R5465 GNDA.n678 GNDA.n499 1.7413
R5466 GNDA.n1999 GNDA.n1998 1.7413
R5467 GNDA.n729 GNDA.n283 1.7413
R5468 GNDA.n2310 GNDA.n228 1.73362
R5469 GNDA.n2423 GNDA.n24 1.6005
R5470 GNDA.n1568 GNDA.n1509 1.2293
R5471 GNDA.n380 GNDA.n379 1.2293
R5472 GNDA.n1752 GNDA.n1020 1.2293
R5473 GNDA.n1328 GNDA.n1208 1.2293
R5474 GNDA.n1166 GNDA.n1048 1.2293
R5475 GNDA.n886 GNDA.n884 1.2293
R5476 GNDA.n580 GNDA.n519 1.2293
R5477 GNDA.n2090 GNDA.n1973 1.2293
R5478 GNDA.n748 GNDA.n746 1.2293
R5479 GNDA.n1668 GNDA.n1666 1.1781
R5480 GNDA.n2210 GNDA.n434 1.1781
R5481 GNDA.n1853 GNDA.n1851 1.1781
R5482 GNDA.n1233 GNDA.n1232 1.1781
R5483 GNDA.n1070 GNDA.n708 1.1781
R5484 GNDA.n990 GNDA.n989 1.1781
R5485 GNDA.n2099 GNDA.n679 1.1781
R5486 GNDA.n2204 GNDA.n456 1.1781
R5487 GNDA.n2251 GNDA.n2249 1.1781
R5488 GNDA.n2128 GNDA.n2127 1.16414
R5489 GNDA.n1602 GNDA.n1601 1.0245
R5490 GNDA.n1573 GNDA.n1510 1.0245
R5491 GNDA.n1595 GNDA.n1574 1.0245
R5492 GNDA.n1594 GNDA.n1575 1.0245
R5493 GNDA.n1590 GNDA.n1589 1.0245
R5494 GNDA.n1585 GNDA.n1579 1.0245
R5495 GNDA.n1584 GNDA.n1580 1.0245
R5496 GNDA.n1658 GNDA.n1489 1.0245
R5497 GNDA.n1657 GNDA.n1490 1.0245
R5498 GNDA.n2236 GNDA.n344 1.0245
R5499 GNDA.n2235 GNDA.n345 1.0245
R5500 GNDA.n2231 GNDA.n2230 1.0245
R5501 GNDA.n2226 GNDA.n348 1.0245
R5502 GNDA.n2225 GNDA.n350 1.0245
R5503 GNDA.n354 GNDA.n352 1.0245
R5504 GNDA.n2220 GNDA.n2219 1.0245
R5505 GNDA.n361 GNDA.n355 1.0245
R5506 GNDA.n2213 GNDA.n362 1.0245
R5507 GNDA.n1788 GNDA.n1787 1.0245
R5508 GNDA.n1759 GNDA.n1021 1.0245
R5509 GNDA.n1781 GNDA.n1760 1.0245
R5510 GNDA.n1780 GNDA.n1761 1.0245
R5511 GNDA.n1776 GNDA.n1775 1.0245
R5512 GNDA.n1771 GNDA.n1765 1.0245
R5513 GNDA.n1770 GNDA.n1766 1.0245
R5514 GNDA.n1844 GNDA.n1001 1.0245
R5515 GNDA.n1843 GNDA.n1002 1.0245
R5516 GNDA.n1327 GNDA.n1211 1.0245
R5517 GNDA.n1215 GNDA.n1213 1.0245
R5518 GNDA.n1322 GNDA.n1321 1.0245
R5519 GNDA.n1317 GNDA.n1216 1.0245
R5520 GNDA.n1316 GNDA.n1220 1.0245
R5521 GNDA.n1224 GNDA.n1222 1.0245
R5522 GNDA.n1311 GNDA.n1310 1.0245
R5523 GNDA.n1306 GNDA.n1225 1.0245
R5524 GNDA.n1305 GNDA.n1229 1.0245
R5525 GNDA.n1165 GNDA.n1050 1.0245
R5526 GNDA.n1054 GNDA.n1052 1.0245
R5527 GNDA.n1160 GNDA.n1159 1.0245
R5528 GNDA.n1155 GNDA.n1055 1.0245
R5529 GNDA.n1154 GNDA.n1059 1.0245
R5530 GNDA.n1063 GNDA.n1061 1.0245
R5531 GNDA.n1149 GNDA.n1148 1.0245
R5532 GNDA.n1144 GNDA.n1064 1.0245
R5533 GNDA.n1143 GNDA.n1068 1.0245
R5534 GNDA.n914 GNDA.n913 1.0245
R5535 GNDA.n912 GNDA.n911 1.0245
R5536 GNDA.n910 GNDA.n887 1.0245
R5537 GNDA.n891 GNDA.n889 1.0245
R5538 GNDA.n905 GNDA.n904 1.0245
R5539 GNDA.n901 GNDA.n900 1.0245
R5540 GNDA.n899 GNDA.n892 1.0245
R5541 GNDA.n895 GNDA.n894 1.0245
R5542 GNDA.n993 GNDA.n868 1.0245
R5543 GNDA.n618 GNDA.n617 1.0245
R5544 GNDA.n613 GNDA.n520 1.0245
R5545 GNDA.n612 GNDA.n586 1.0245
R5546 GNDA.n590 GNDA.n588 1.0245
R5547 GNDA.n607 GNDA.n606 1.0245
R5548 GNDA.n602 GNDA.n591 1.0245
R5549 GNDA.n601 GNDA.n596 1.0245
R5550 GNDA.n598 GNDA.n501 1.0245
R5551 GNDA.n674 GNDA.n673 1.0245
R5552 GNDA.n2089 GNDA.n1976 1.0245
R5553 GNDA.n1980 GNDA.n1978 1.0245
R5554 GNDA.n2084 GNDA.n2083 1.0245
R5555 GNDA.n2079 GNDA.n1981 1.0245
R5556 GNDA.n2078 GNDA.n1985 1.0245
R5557 GNDA.n1989 GNDA.n1987 1.0245
R5558 GNDA.n2073 GNDA.n2072 1.0245
R5559 GNDA.n2068 GNDA.n1990 1.0245
R5560 GNDA.n2067 GNDA.n1994 1.0245
R5561 GNDA.n773 GNDA.n772 1.0245
R5562 GNDA.n771 GNDA.n770 1.0245
R5563 GNDA.n769 GNDA.n749 1.0245
R5564 GNDA.n753 GNDA.n751 1.0245
R5565 GNDA.n764 GNDA.n763 1.0245
R5566 GNDA.n760 GNDA.n759 1.0245
R5567 GNDA.n758 GNDA.n754 1.0245
R5568 GNDA.n829 GNDA.n726 1.0245
R5569 GNDA.n828 GNDA.n727 1.0245
R5570 GNDA.n16 GNDA.n14 0.563
R5571 GNDA.n18 GNDA.n16 0.563
R5572 GNDA.n20 GNDA.n18 0.563
R5573 GNDA.n22 GNDA.n20 0.563
R5574 GNDA.n48 GNDA.n47 0.563
R5575 GNDA.n48 GNDA.n44 0.563
R5576 GNDA.n1449 GNDA.n1447 0.563
R5577 GNDA.n1453 GNDA.n1451 0.563
R5578 GNDA.n1455 GNDA.n1453 0.563
R5579 GNDA.n1457 GNDA.n1455 0.563
R5580 GNDA.n1461 GNDA.n1459 0.563
R5581 GNDA.n1463 GNDA.n1461 0.563
R5582 GNDA.n5 GNDA.n3 0.563
R5583 GNDA.n7 GNDA.n5 0.563
R5584 GNDA.n9 GNDA.n7 0.563
R5585 GNDA.n11 GNDA.n9 0.563
R5586 GNDA.n173 GNDA.n171 0.563
R5587 GNDA.n171 GNDA.n169 0.563
R5588 GNDA.n169 GNDA.n167 0.563
R5589 GNDA.n167 GNDA.n165 0.563
R5590 GNDA.n165 GNDA.n163 0.563
R5591 GNDA.n163 GNDA.n161 0.563
R5592 GNDA.n161 GNDA.n159 0.563
R5593 GNDA.n159 GNDA.n157 0.563
R5594 GNDA.n157 GNDA.n155 0.563
R5595 GNDA.n155 GNDA.n153 0.563
R5596 GNDA.n153 GNDA.n151 0.563
R5597 GNDA.n2426 GNDA.n0 0.53175
R5598 GNDA.n179 GNDA.n177 0.5005
R5599 GNDA.n2381 GNDA.n2380 0.5005
R5600 GNDA.n200 GNDA.t26 0.467591
R5601 GNDA.n2351 GNDA.t107 0.467591
R5602 GNDA.t121 GNDA.n2295 0.419041
R5603 GNDA.n2314 GNDA.n2312 0.41175
R5604 GNDA.n2312 GNDA.n2311 0.311875
R5605 GNDA.n174 GNDA.n173 0.28175
R5606 GNDA.n2315 GNDA.n227 0.276625
R5607 GNDA.n151 GNDA.n148 0.2505
R5608 GNDA.n1464 GNDA.n227 0.22375
R5609 GNDA.n1861 GNDA 0.129793
R5610 GNDA.n981 GNDA 0.129793
R5611 GNDA.n2259 GNDA 0.129793
R5612 GNDA.n1465 GNDA.n1464 0.100375
R5613 GNDA.n2311 GNDA.n2310 0.076875
R5614 GNDA.n1694 GNDA.n1035 0.0479074
R5615 GNDA.n1677 GNDA 0.0479074
R5616 GNDA.n1028 GNDA.n706 0.0479074
R5617 GNDA.n1738 GNDA 0.0479074
R5618 GNDA.n1947 GNDA.n681 0.0479074
R5619 GNDA.n1180 GNDA 0.0479074
R5620 GNDA.n691 GNDA.n457 0.0479074
R5621 GNDA.n1908 GNDA 0.0479074
R5622 GNDA.n2166 GNDA.n467 0.0479074
R5623 GNDA GNDA.n2192 0.0479074
R5624 GNDA.n475 GNDA.n474 0.0479074
R5625 GNDA GNDA.n1963 0.0479074
R5626 GNDA.n2247 GNDA.n287 0.0319432
R5627 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t15 354.854
R5628 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t30 346.8
R5629 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 339.522
R5630 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n4 339.522
R5631 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n9 335.022
R5632 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t6 275.909
R5633 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 227.909
R5634 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 222.034
R5635 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t27 184.097
R5636 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t19 184.097
R5637 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t31 184.097
R5638 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t14 184.097
R5639 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 166.05
R5640 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 166.05
R5641 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t3 48.0005
R5642 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t0 48.0005
R5643 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t1 48.0005
R5644 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t7 48.0005
R5645 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t9 39.4005
R5646 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t5 39.4005
R5647 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t8 39.4005
R5648 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t4 39.4005
R5649 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t10 39.4005
R5650 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t2 39.4005
R5651 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n2 33.1711
R5652 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n0 5.6255
R5653 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 5.28175
R5654 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R5655 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t29 4.8295
R5656 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t25 4.8295
R5657 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t35 4.8295
R5658 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t33 4.8295
R5659 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t17 4.8295
R5660 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t28 4.8295
R5661 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n7 4.5005
R5662 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t11 4.5005
R5663 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t32 4.5005
R5664 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t34 4.5005
R5665 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t21 4.5005
R5666 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t12 4.5005
R5667 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t16 4.5005
R5668 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t26 4.5005
R5669 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t22 4.5005
R5670 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.5005
R5671 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.5005
R5672 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t13 4.5005
R5673 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t18 4.5005
R5674 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t36 4.5005
R5675 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.8075
R5676 bgr_0.cap_res1.t20 bgr_0.cap_res1.t17 178.633
R5677 bgr_0.cap_res1.t14 bgr_0.cap_res1.t0 0.1603
R5678 bgr_0.cap_res1.t10 bgr_0.cap_res1.t6 0.1603
R5679 bgr_0.cap_res1.t9 bgr_0.cap_res1.t15 0.1603
R5680 bgr_0.cap_res1.t7 bgr_0.cap_res1.t3 0.1603
R5681 bgr_0.cap_res1.t16 bgr_0.cap_res1.t1 0.1603
R5682 bgr_0.cap_res1.t12 bgr_0.cap_res1.t8 0.1603
R5683 bgr_0.cap_res1.t2 bgr_0.cap_res1.t5 0.1603
R5684 bgr_0.cap_res1.t19 bgr_0.cap_res1.t13 0.1603
R5685 bgr_0.cap_res1.n1 bgr_0.cap_res1.t4 0.159278
R5686 bgr_0.cap_res1.n2 bgr_0.cap_res1.t18 0.159278
R5687 bgr_0.cap_res1.n3 bgr_0.cap_res1.t11 0.159278
R5688 bgr_0.cap_res1.n3 bgr_0.cap_res1.t14 0.1368
R5689 bgr_0.cap_res1.n3 bgr_0.cap_res1.t10 0.1368
R5690 bgr_0.cap_res1.n2 bgr_0.cap_res1.t9 0.1368
R5691 bgr_0.cap_res1.n2 bgr_0.cap_res1.t7 0.1368
R5692 bgr_0.cap_res1.n1 bgr_0.cap_res1.t16 0.1368
R5693 bgr_0.cap_res1.n1 bgr_0.cap_res1.t12 0.1368
R5694 bgr_0.cap_res1.n0 bgr_0.cap_res1.t2 0.1368
R5695 bgr_0.cap_res1.n0 bgr_0.cap_res1.t19 0.1368
R5696 bgr_0.cap_res1.t4 bgr_0.cap_res1.n0 0.00152174
R5697 bgr_0.cap_res1.t18 bgr_0.cap_res1.n1 0.00152174
R5698 bgr_0.cap_res1.t11 bgr_0.cap_res1.n2 0.00152174
R5699 bgr_0.cap_res1.t17 bgr_0.cap_res1.n3 0.00152174
R5700 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 114.719
R5701 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5702 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5703 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 114.156
R5704 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5705 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5706 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5707 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5708 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5709 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5710 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5711 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5712 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5713 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5714 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5715 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5716 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5717 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5718 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5719 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5720 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5721 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5722 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5723 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5724 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5725 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5726 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5727 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5728 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5729 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5730 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5731 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5732 two_stage_opamp_dummy_magic_0.VD2.t18 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5733 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5734 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5735 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5736 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5737 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5738 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5739 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5740 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n8 0.563
R5741 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.n5 145.989
R5742 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n6 145.989
R5743 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n11 145.427
R5744 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n9 145.427
R5745 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n7 145.427
R5746 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n14 140.927
R5747 two_stage_opamp_dummy_magic_0.VOUT-.t18 two_stage_opamp_dummy_magic_0.VOUT-.n96 113.192
R5748 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n0 95.7303
R5749 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n3 94.6053
R5750 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n1 94.6053
R5751 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.n15 20.688
R5752 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.n94 11.7059
R5753 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n95 10.438
R5754 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t5 6.56717
R5755 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t0 6.56717
R5756 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t2 6.56717
R5757 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t7 6.56717
R5758 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t1 6.56717
R5759 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t13 6.56717
R5760 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t9 6.56717
R5761 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t10 6.56717
R5762 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.t8 6.56717
R5763 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.t15 6.56717
R5764 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t14 6.56717
R5765 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t6 6.56717
R5766 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t85 4.8295
R5767 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t131 4.8295
R5768 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t31 4.8295
R5769 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t62 4.8295
R5770 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t114 4.8295
R5771 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t40 4.8295
R5772 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t34 4.8295
R5773 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t136 4.8295
R5774 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t70 4.8295
R5775 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t36 4.8295
R5776 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.t95 4.8295
R5777 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t66 4.8295
R5778 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.t55 4.8295
R5779 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t29 4.8295
R5780 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.t91 4.8295
R5781 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t58 4.8295
R5782 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.t49 4.8295
R5783 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t20 4.8295
R5784 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.t148 4.8295
R5785 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t122 4.8295
R5786 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.t44 4.8295
R5787 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t152 4.8295
R5788 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.t142 4.8295
R5789 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t116 4.8295
R5790 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t108 4.8295
R5791 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t28 4.8295
R5792 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t24 4.8295
R5793 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t129 4.8295
R5794 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t61 4.8295
R5795 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t32 4.8295
R5796 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t100 4.8295
R5797 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t71 4.8295
R5798 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t69 4.8295
R5799 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t35 4.8295
R5800 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t77 4.8295
R5801 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t26 4.8154
R5802 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t59 4.8154
R5803 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t37 4.8154
R5804 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t81 4.8154
R5805 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t132 4.806
R5806 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t115 4.806
R5807 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t146 4.806
R5808 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.t46 4.806
R5809 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t87 4.806
R5810 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t65 4.806
R5811 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t102 4.806
R5812 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t134 4.806
R5813 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t120 4.806
R5814 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t155 4.806
R5815 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t48 4.806
R5816 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t92 4.806
R5817 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t42 4.806
R5818 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t130 4.806
R5819 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t84 4.806
R5820 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t125 4.806
R5821 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t74 4.806
R5822 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t23 4.806
R5823 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t64 4.806
R5824 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t150 4.806
R5825 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.t96 4.5005
R5826 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t57 4.5005
R5827 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t104 4.5005
R5828 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.t73 4.5005
R5829 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t138 4.5005
R5830 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.t107 4.5005
R5831 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t41 4.5005
R5832 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.t143 4.5005
R5833 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t21 4.5005
R5834 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.t126 4.5005
R5835 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t119 4.5005
R5836 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t82 4.5005
R5837 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t97 4.5005
R5838 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t63 4.5005
R5839 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t27 4.5005
R5840 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t45 4.5005
R5841 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.t144 4.5005
R5842 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t112 4.5005
R5843 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t76 4.5005
R5844 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t93 4.5005
R5845 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.t56 4.5005
R5846 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t19 4.5005
R5847 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t52 4.5005
R5848 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.t156 4.5005
R5849 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t121 4.5005
R5850 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t89 4.5005
R5851 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.t50 4.5005
R5852 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t151 4.5005
R5853 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.t43 4.5005
R5854 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.t145 4.5005
R5855 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t118 4.5005
R5856 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.t141 4.5005
R5857 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.t111 4.5005
R5858 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t80 4.5005
R5859 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.t39 4.5005
R5860 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.t139 4.5005
R5861 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t109 4.5005
R5862 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.t135 4.5005
R5863 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.t103 4.5005
R5864 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t72 4.5005
R5865 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.t99 4.5005
R5866 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.t68 4.5005
R5867 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t33 4.5005
R5868 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.t133 4.5005
R5869 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.t98 4.5005
R5870 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t67 4.5005
R5871 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.t94 4.5005
R5872 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.t60 4.5005
R5873 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t30 4.5005
R5874 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.t101 4.5005
R5875 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t149 4.5005
R5876 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t88 4.5005
R5877 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t51 4.5005
R5878 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t137 4.5005
R5879 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t106 4.5005
R5880 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t75 4.5005
R5881 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t25 4.5005
R5882 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t128 4.5005
R5883 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t90 4.5005
R5884 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t54 4.5005
R5885 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t140 4.5005
R5886 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.t110 4.5005
R5887 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t79 4.5005
R5888 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t113 4.5005
R5889 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.t78 4.5005
R5890 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t38 4.5005
R5891 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t147 4.5005
R5892 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.t117 4.5005
R5893 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t83 4.5005
R5894 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t47 4.5005
R5895 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.t153 4.5005
R5896 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t123 4.5005
R5897 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t154 4.5005
R5898 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.t124 4.5005
R5899 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t86 4.5005
R5900 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.t105 4.5005
R5901 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.t53 4.5005
R5902 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.t22 4.5005
R5903 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t127 4.5005
R5904 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n13 4.5005
R5905 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t3 3.42907
R5906 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t17 3.42907
R5907 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t12 3.42907
R5908 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t4 3.42907
R5909 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t16 3.42907
R5910 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t11 3.42907
R5911 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n4 2.03175
R5912 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n2 1.1255
R5913 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n8 0.563
R5914 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n10 0.563
R5915 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.n12 0.563
R5916 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.n42 0.3295
R5917 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.n44 0.3295
R5918 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.n46 0.3295
R5919 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.n48 0.3295
R5920 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.n50 0.3295
R5921 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.n52 0.3295
R5922 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.n53 0.3295
R5923 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.n54 0.3295
R5924 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.n55 0.3295
R5925 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.n56 0.3295
R5926 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n57 0.3295
R5927 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.n58 0.3295
R5928 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.n59 0.3295
R5929 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.n60 0.3295
R5930 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n61 0.3295
R5931 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n62 0.3295
R5932 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n64 0.3295
R5933 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n65 0.3295
R5934 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.n67 0.3295
R5935 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.n68 0.3295
R5936 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.n70 0.3295
R5937 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.n71 0.3295
R5938 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.n73 0.3295
R5939 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.n74 0.3295
R5940 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.n76 0.3295
R5941 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.n77 0.3295
R5942 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.n79 0.3295
R5943 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.n80 0.3295
R5944 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.n82 0.3295
R5945 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.n83 0.3295
R5946 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n85 0.3295
R5947 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n86 0.3295
R5948 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n88 0.3295
R5949 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n89 0.3295
R5950 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.n16 0.3295
R5951 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.n18 0.3295
R5952 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.n19 0.3295
R5953 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.n20 0.3295
R5954 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.n21 0.3295
R5955 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.n22 0.3295
R5956 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.n23 0.3295
R5957 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.n24 0.3295
R5958 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.n25 0.3295
R5959 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.n26 0.3295
R5960 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n27 0.3295
R5961 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n28 0.3295
R5962 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n30 0.3295
R5963 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n31 0.3295
R5964 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n33 0.3295
R5965 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n34 0.3295
R5966 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n36 0.3295
R5967 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n37 0.3295
R5968 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n39 0.3295
R5969 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n40 0.3295
R5970 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.n93 0.3295
R5971 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.n92 0.3295
R5972 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.n91 0.3295
R5973 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.n45 0.306
R5974 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n47 0.306
R5975 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.n49 0.306
R5976 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.n51 0.306
R5977 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n43 0.2825
R5978 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n63 0.2825
R5979 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.n66 0.2825
R5980 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.n69 0.2825
R5981 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.n72 0.2825
R5982 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.n75 0.2825
R5983 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.n78 0.2825
R5984 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.n81 0.2825
R5985 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n84 0.2825
R5986 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n87 0.2825
R5987 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n17 0.2825
R5988 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n29 0.2825
R5989 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n32 0.2825
R5990 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n35 0.2825
R5991 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n38 0.2825
R5992 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.n41 0.2825
R5993 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.n90 0.2825
R5994 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.083
R5995 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.922875
R5996 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1603
R5997 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.1603
R5998 two_stage_opamp_dummy_magic_0.cap_res_X.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R5999 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R6000 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R6001 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1603
R6002 two_stage_opamp_dummy_magic_0.cap_res_X.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R6003 two_stage_opamp_dummy_magic_0.cap_res_X.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.1603
R6004 two_stage_opamp_dummy_magic_0.cap_res_X.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R6005 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.1603
R6006 two_stage_opamp_dummy_magic_0.cap_res_X.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.1603
R6007 two_stage_opamp_dummy_magic_0.cap_res_X.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R6008 two_stage_opamp_dummy_magic_0.cap_res_X.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R6009 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1603
R6010 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1603
R6011 two_stage_opamp_dummy_magic_0.cap_res_X.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1603
R6012 two_stage_opamp_dummy_magic_0.cap_res_X.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1603
R6013 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R6014 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.1603
R6015 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1603
R6016 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.1603
R6017 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.1603
R6018 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R6019 two_stage_opamp_dummy_magic_0.cap_res_X.t3 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R6020 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R6021 two_stage_opamp_dummy_magic_0.cap_res_X.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1603
R6022 two_stage_opamp_dummy_magic_0.cap_res_X.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R6023 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.1603
R6024 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1603
R6025 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1603
R6026 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R6027 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.1603
R6028 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R6029 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R6030 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R6031 two_stage_opamp_dummy_magic_0.cap_res_X.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R6032 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1603
R6033 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1603
R6034 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1603
R6035 two_stage_opamp_dummy_magic_0.cap_res_X.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1603
R6036 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1603
R6037 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1603
R6038 two_stage_opamp_dummy_magic_0.cap_res_X.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R6039 two_stage_opamp_dummy_magic_0.cap_res_X.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R6040 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1603
R6041 two_stage_opamp_dummy_magic_0.cap_res_X.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1603
R6042 two_stage_opamp_dummy_magic_0.cap_res_X.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1603
R6043 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R6044 two_stage_opamp_dummy_magic_0.cap_res_X.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R6045 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.1603
R6046 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R6047 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1603
R6048 two_stage_opamp_dummy_magic_0.cap_res_X.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R6049 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R6050 two_stage_opamp_dummy_magic_0.cap_res_X.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R6051 two_stage_opamp_dummy_magic_0.cap_res_X.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R6052 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R6053 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R6054 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.159278
R6055 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R6056 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R6057 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R6058 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R6059 two_stage_opamp_dummy_magic_0.cap_res_X.t33 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R6060 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R6061 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R6062 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R6063 two_stage_opamp_dummy_magic_0.cap_res_X.t89 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R6064 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R6065 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.159278
R6066 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.159278
R6067 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.159278
R6068 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.159278
R6069 two_stage_opamp_dummy_magic_0.cap_res_X.t1 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.159278
R6070 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.159278
R6071 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.159278
R6072 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.159278
R6073 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.159278
R6074 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.159278
R6075 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.159278
R6076 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.159278
R6077 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.159278
R6078 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.159278
R6079 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.159278
R6080 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.159278
R6081 two_stage_opamp_dummy_magic_0.cap_res_X.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.137822
R6082 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1368
R6083 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1368
R6084 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R6085 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1368
R6086 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R6087 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1368
R6088 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1368
R6089 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1368
R6090 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R6091 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1368
R6092 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1368
R6093 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1368
R6094 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R6095 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R6096 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1368
R6097 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1368
R6098 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R6099 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R6100 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1368
R6101 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.1368
R6102 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.1368
R6103 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.1368
R6104 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1368
R6105 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.1368
R6106 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1368
R6107 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1368
R6108 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1368
R6109 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R6110 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1368
R6111 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R6112 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R6113 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.114322
R6114 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R6115 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R6116 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R6117 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.1133
R6118 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.1133
R6119 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.1133
R6120 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.1133
R6121 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.1133
R6122 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.1133
R6123 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R6124 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R6125 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R6126 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R6127 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R6128 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R6129 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R6130 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R6131 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R6132 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R6133 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.00152174
R6134 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.00152174
R6135 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.00152174
R6136 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R6137 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R6138 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R6139 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.00152174
R6140 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.00152174
R6141 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R6142 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.00152174
R6143 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R6144 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.00152174
R6145 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.00152174
R6146 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R6147 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.00152174
R6148 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.00152174
R6149 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.00152174
R6150 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.00152174
R6151 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.00152174
R6152 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.00152174
R6153 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R6154 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R6155 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R6156 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.00152174
R6157 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R6158 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.00152174
R6159 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.00152174
R6160 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.00152174
R6161 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.00152174
R6162 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.00152174
R6163 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.00152174
R6164 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R6165 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.00152174
R6166 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R6167 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.00152174
R6168 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R6169 bgr_0.Vbe2.n145 bgr_0.Vbe2.n144 413.99
R6170 bgr_0.Vbe2.n136 bgr_0.Vbe2.t8 162.458
R6171 bgr_0.Vbe2.n146 bgr_0.Vbe2.n145 84.0884
R6172 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 83.5719
R6173 bgr_0.Vbe2.n55 bgr_0.Vbe2.n48 83.5719
R6174 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 83.5719
R6175 bgr_0.Vbe2.n127 bgr_0.Vbe2.n6 83.5719
R6176 bgr_0.Vbe2.n122 bgr_0.Vbe2.n7 83.5719
R6177 bgr_0.Vbe2.n45 bgr_0.Vbe2.n44 83.5719
R6178 bgr_0.Vbe2.n43 bgr_0.Vbe2.n42 83.5719
R6179 bgr_0.Vbe2.n41 bgr_0.Vbe2.n40 83.5719
R6180 bgr_0.Vbe2.n78 bgr_0.Vbe2.n77 83.5719
R6181 bgr_0.Vbe2.n76 bgr_0.Vbe2.n75 83.5719
R6182 bgr_0.Vbe2.n27 bgr_0.Vbe2.n26 83.5719
R6183 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 83.5719
R6184 bgr_0.Vbe2.n22 bgr_0.Vbe2.n20 83.5719
R6185 bgr_0.Vbe2.n91 bgr_0.Vbe2.n19 83.5719
R6186 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 83.5719
R6187 bgr_0.Vbe2.n17 bgr_0.Vbe2.n16 83.5719
R6188 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 83.5719
R6189 bgr_0.Vbe2.n112 bgr_0.Vbe2.n111 83.5719
R6190 bgr_0.Vbe2.n110 bgr_0.Vbe2.n109 83.5719
R6191 bgr_0.Vbe2.n143 bgr_0.Vbe2.n1 83.5719
R6192 bgr_0.Vbe2.n142 bgr_0.Vbe2.n0 83.5719
R6193 bgr_0.Vbe2.n141 bgr_0.Vbe2.n140 83.5719
R6194 bgr_0.Vbe2.n132 bgr_0.Vbe2.n4 83.5719
R6195 bgr_0.Vbe2.n72 bgr_0.Vbe2.n26 73.8495
R6196 bgr_0.Vbe2.n59 bgr_0.Vbe2.n58 73.3165
R6197 bgr_0.Vbe2.n129 bgr_0.Vbe2.n6 73.3165
R6198 bgr_0.Vbe2.n44 bgr_0.Vbe2.n36 73.3165
R6199 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 73.3165
R6200 bgr_0.Vbe2.n98 bgr_0.Vbe2.n97 73.3165
R6201 bgr_0.Vbe2.n115 bgr_0.Vbe2.n114 73.3165
R6202 bgr_0.Vbe2.n54 bgr_0.Vbe2.n49 73.19
R6203 bgr_0.Vbe2.n41 bgr_0.Vbe2.n39 73.19
R6204 bgr_0.Vbe2.n77 bgr_0.Vbe2.n23 73.19
R6205 bgr_0.Vbe2.n93 bgr_0.Vbe2.n19 73.19
R6206 bgr_0.Vbe2.n110 bgr_0.Vbe2.n13 73.19
R6207 bgr_0.Vbe2.n133 bgr_0.Vbe2.n132 73.19
R6208 bgr_0.Vbe2.n123 bgr_0.Vbe2.t4 65.0299
R6209 bgr_0.Vbe2.t6 bgr_0.Vbe2.n14 65.0299
R6210 bgr_0.Vbe2.n59 bgr_0.Vbe2.n55 26.074
R6211 bgr_0.Vbe2.n122 bgr_0.Vbe2.n6 26.074
R6212 bgr_0.Vbe2.n44 bgr_0.Vbe2.n43 26.074
R6213 bgr_0.Vbe2.n76 bgr_0.Vbe2.n26 26.074
R6214 bgr_0.Vbe2.n85 bgr_0.Vbe2.n22 26.074
R6215 bgr_0.Vbe2.n98 bgr_0.Vbe2.n17 26.074
R6216 bgr_0.Vbe2.n114 bgr_0.Vbe2.n112 26.074
R6217 bgr_0.Vbe2.n142 bgr_0.Vbe2.n141 26.074
R6218 bgr_0.Vbe2.n143 bgr_0.Vbe2.n142 26.074
R6219 bgr_0.Vbe2.n145 bgr_0.Vbe2.n143 26.074
R6220 bgr_0.Vbe2.t0 bgr_0.Vbe2.n54 25.7843
R6221 bgr_0.Vbe2.t2 bgr_0.Vbe2.n41 25.7843
R6222 bgr_0.Vbe2.n77 bgr_0.Vbe2.t3 25.7843
R6223 bgr_0.Vbe2.t1 bgr_0.Vbe2.n19 25.7843
R6224 bgr_0.Vbe2.t5 bgr_0.Vbe2.n110 25.7843
R6225 bgr_0.Vbe2.n132 bgr_0.Vbe2.t7 25.7843
R6226 bgr_0.Vbe2.n116 bgr_0.Vbe2.n104 9.3005
R6227 bgr_0.Vbe2.n104 bgr_0.Vbe2.n11 9.3005
R6228 bgr_0.Vbe2.n104 bgr_0.Vbe2.n12 9.3005
R6229 bgr_0.Vbe2.n120 bgr_0.Vbe2.n104 9.3005
R6230 bgr_0.Vbe2.n106 bgr_0.Vbe2.n11 9.3005
R6231 bgr_0.Vbe2.n106 bgr_0.Vbe2.n12 9.3005
R6232 bgr_0.Vbe2.n106 bgr_0.Vbe2.n9 9.3005
R6233 bgr_0.Vbe2.n120 bgr_0.Vbe2.n106 9.3005
R6234 bgr_0.Vbe2.n121 bgr_0.Vbe2.n11 9.3005
R6235 bgr_0.Vbe2.n121 bgr_0.Vbe2.n10 9.3005
R6236 bgr_0.Vbe2.n121 bgr_0.Vbe2.n12 9.3005
R6237 bgr_0.Vbe2.n121 bgr_0.Vbe2.n9 9.3005
R6238 bgr_0.Vbe2.n121 bgr_0.Vbe2.n120 9.3005
R6239 bgr_0.Vbe2.n120 bgr_0.Vbe2.n108 9.3005
R6240 bgr_0.Vbe2.n108 bgr_0.Vbe2.n9 9.3005
R6241 bgr_0.Vbe2.n108 bgr_0.Vbe2.n12 9.3005
R6242 bgr_0.Vbe2.n108 bgr_0.Vbe2.n10 9.3005
R6243 bgr_0.Vbe2.n120 bgr_0.Vbe2.n103 9.3005
R6244 bgr_0.Vbe2.n103 bgr_0.Vbe2.n9 9.3005
R6245 bgr_0.Vbe2.n103 bgr_0.Vbe2.n12 9.3005
R6246 bgr_0.Vbe2.n103 bgr_0.Vbe2.n10 9.3005
R6247 bgr_0.Vbe2.n116 bgr_0.Vbe2.n103 9.3005
R6248 bgr_0.Vbe2.n119 bgr_0.Vbe2.n11 9.3005
R6249 bgr_0.Vbe2.n119 bgr_0.Vbe2.n10 9.3005
R6250 bgr_0.Vbe2.n119 bgr_0.Vbe2.n12 9.3005
R6251 bgr_0.Vbe2.n120 bgr_0.Vbe2.n119 9.3005
R6252 bgr_0.Vbe2.n69 bgr_0.Vbe2.n68 9.3005
R6253 bgr_0.Vbe2.n68 bgr_0.Vbe2.n67 9.3005
R6254 bgr_0.Vbe2.n68 bgr_0.Vbe2.n29 9.3005
R6255 bgr_0.Vbe2.n68 bgr_0.Vbe2.n30 9.3005
R6256 bgr_0.Vbe2.n67 bgr_0.Vbe2.n65 9.3005
R6257 bgr_0.Vbe2.n65 bgr_0.Vbe2.n29 9.3005
R6258 bgr_0.Vbe2.n65 bgr_0.Vbe2.n31 9.3005
R6259 bgr_0.Vbe2.n65 bgr_0.Vbe2.n30 9.3005
R6260 bgr_0.Vbe2.n67 bgr_0.Vbe2.n64 9.3005
R6261 bgr_0.Vbe2.n64 bgr_0.Vbe2.n32 9.3005
R6262 bgr_0.Vbe2.n64 bgr_0.Vbe2.n29 9.3005
R6263 bgr_0.Vbe2.n64 bgr_0.Vbe2.n31 9.3005
R6264 bgr_0.Vbe2.n64 bgr_0.Vbe2.n30 9.3005
R6265 bgr_0.Vbe2.n33 bgr_0.Vbe2.n30 9.3005
R6266 bgr_0.Vbe2.n33 bgr_0.Vbe2.n31 9.3005
R6267 bgr_0.Vbe2.n33 bgr_0.Vbe2.n29 9.3005
R6268 bgr_0.Vbe2.n33 bgr_0.Vbe2.n32 9.3005
R6269 bgr_0.Vbe2.n70 bgr_0.Vbe2.n30 9.3005
R6270 bgr_0.Vbe2.n70 bgr_0.Vbe2.n31 9.3005
R6271 bgr_0.Vbe2.n70 bgr_0.Vbe2.n29 9.3005
R6272 bgr_0.Vbe2.n70 bgr_0.Vbe2.n32 9.3005
R6273 bgr_0.Vbe2.n70 bgr_0.Vbe2.n69 9.3005
R6274 bgr_0.Vbe2.n67 bgr_0.Vbe2.n66 9.3005
R6275 bgr_0.Vbe2.n66 bgr_0.Vbe2.n32 9.3005
R6276 bgr_0.Vbe2.n66 bgr_0.Vbe2.n29 9.3005
R6277 bgr_0.Vbe2.n66 bgr_0.Vbe2.n30 9.3005
R6278 bgr_0.Vbe2.n118 bgr_0.Vbe2.n9 4.64654
R6279 bgr_0.Vbe2.n105 bgr_0.Vbe2.n10 4.64654
R6280 bgr_0.Vbe2.n116 bgr_0.Vbe2.n8 4.64654
R6281 bgr_0.Vbe2.n107 bgr_0.Vbe2.n11 4.64654
R6282 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 4.64654
R6283 bgr_0.Vbe2.n37 bgr_0.Vbe2.n31 4.64654
R6284 bgr_0.Vbe2.n38 bgr_0.Vbe2.n32 4.64654
R6285 bgr_0.Vbe2.n69 bgr_0.Vbe2.n35 4.64654
R6286 bgr_0.Vbe2.n67 bgr_0.Vbe2.n28 4.64654
R6287 bgr_0.Vbe2.n69 bgr_0.Vbe2.n34 4.64654
R6288 bgr_0.Vbe2.n49 bgr_0.Vbe2.n3 2.36206
R6289 bgr_0.Vbe2.n81 bgr_0.Vbe2.n23 2.36206
R6290 bgr_0.Vbe2.n94 bgr_0.Vbe2.n93 2.36206
R6291 bgr_0.Vbe2.n133 bgr_0.Vbe2.n131 2.36206
R6292 bgr_0.Vbe2.n58 bgr_0.Vbe2.n56 2.19742
R6293 bgr_0.Vbe2.n130 bgr_0.Vbe2.n129 2.19742
R6294 bgr_0.Vbe2.n84 bgr_0.Vbe2.n82 2.19742
R6295 bgr_0.Vbe2.n97 bgr_0.Vbe2.n95 2.19742
R6296 bgr_0.Vbe2.n123 bgr_0.Vbe2.n7 1.56363
R6297 bgr_0.Vbe2.n16 bgr_0.Vbe2.n14 1.56363
R6298 bgr_0.Vbe2.n96 bgr_0.Vbe2.n15 1.5505
R6299 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 1.5505
R6300 bgr_0.Vbe2.n83 bgr_0.Vbe2.n21 1.5505
R6301 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 1.5505
R6302 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 1.5505
R6303 bgr_0.Vbe2.n92 bgr_0.Vbe2.n18 1.5505
R6304 bgr_0.Vbe2.n74 bgr_0.Vbe2.n73 1.5505
R6305 bgr_0.Vbe2.n80 bgr_0.Vbe2.n79 1.5505
R6306 bgr_0.Vbe2.n25 bgr_0.Vbe2.n24 1.5505
R6307 bgr_0.Vbe2.n128 bgr_0.Vbe2.n5 1.5505
R6308 bgr_0.Vbe2.n126 bgr_0.Vbe2.n125 1.5505
R6309 bgr_0.Vbe2.n57 bgr_0.Vbe2.n47 1.5505
R6310 bgr_0.Vbe2.n62 bgr_0.Vbe2.n61 1.5505
R6311 bgr_0.Vbe2.n52 bgr_0.Vbe2.n46 1.5505
R6312 bgr_0.Vbe2.n51 bgr_0.Vbe2.n50 1.5505
R6313 bgr_0.Vbe2.n147 bgr_0.Vbe2.n146 1.5505
R6314 bgr_0.Vbe2.n149 bgr_0.Vbe2.n148 1.5505
R6315 bgr_0.Vbe2.n139 bgr_0.Vbe2.n2 1.5505
R6316 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 1.5505
R6317 bgr_0.Vbe2.n135 bgr_0.Vbe2.n134 1.5505
R6318 bgr_0.Vbe2.n53 bgr_0.Vbe2.n51 1.25468
R6319 bgr_0.Vbe2.n40 bgr_0.Vbe2.n31 1.25468
R6320 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 1.25468
R6321 bgr_0.Vbe2.n92 bgr_0.Vbe2.n91 1.25468
R6322 bgr_0.Vbe2.n109 bgr_0.Vbe2.n9 1.25468
R6323 bgr_0.Vbe2.n134 bgr_0.Vbe2.n4 1.25468
R6324 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 1.19225
R6325 bgr_0.Vbe2.n129 bgr_0.Vbe2.n128 1.19225
R6326 bgr_0.Vbe2.n67 bgr_0.Vbe2.n36 1.19225
R6327 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 1.19225
R6328 bgr_0.Vbe2.n97 bgr_0.Vbe2.n96 1.19225
R6329 bgr_0.Vbe2.n115 bgr_0.Vbe2.n11 1.19225
R6330 bgr_0.Vbe2.n146 bgr_0.Vbe2.n1 1.14402
R6331 bgr_0.Vbe2.n52 bgr_0.Vbe2.n48 1.07024
R6332 bgr_0.Vbe2.n42 bgr_0.Vbe2.n29 1.07024
R6333 bgr_0.Vbe2.n75 bgr_0.Vbe2.n25 1.07024
R6334 bgr_0.Vbe2.n90 bgr_0.Vbe2.n20 1.07024
R6335 bgr_0.Vbe2.n111 bgr_0.Vbe2.n12 1.07024
R6336 bgr_0.Vbe2.n140 bgr_0.Vbe2.n138 1.07024
R6337 bgr_0.Vbe2.n51 bgr_0.Vbe2.n49 1.0237
R6338 bgr_0.Vbe2.n39 bgr_0.Vbe2.n31 1.0237
R6339 bgr_0.Vbe2.n79 bgr_0.Vbe2.n23 1.0237
R6340 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 1.0237
R6341 bgr_0.Vbe2.n13 bgr_0.Vbe2.n9 1.0237
R6342 bgr_0.Vbe2.n134 bgr_0.Vbe2.n133 1.0237
R6343 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 0.885803
R6344 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 0.885803
R6345 bgr_0.Vbe2.n45 bgr_0.Vbe2.n32 0.885803
R6346 bgr_0.Vbe2.n74 bgr_0.Vbe2.n27 0.885803
R6347 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 0.885803
R6348 bgr_0.Vbe2.n100 bgr_0.Vbe2.n99 0.885803
R6349 bgr_0.Vbe2.n113 bgr_0.Vbe2.n10 0.885803
R6350 bgr_0.Vbe2.n139 bgr_0.Vbe2.n0 0.885803
R6351 bgr_0.Vbe2.n39 bgr_0.Vbe2.n30 0.812055
R6352 bgr_0.Vbe2.n120 bgr_0.Vbe2.n13 0.812055
R6353 bgr_0.Vbe2.n61 bgr_0.Vbe2.n48 0.77514
R6354 bgr_0.Vbe2.n126 bgr_0.Vbe2.n7 0.77514
R6355 bgr_0.Vbe2.n42 bgr_0.Vbe2.n32 0.77514
R6356 bgr_0.Vbe2.n75 bgr_0.Vbe2.n74 0.77514
R6357 bgr_0.Vbe2.n87 bgr_0.Vbe2.n20 0.77514
R6358 bgr_0.Vbe2.n100 bgr_0.Vbe2.n16 0.77514
R6359 bgr_0.Vbe2.n111 bgr_0.Vbe2.n10 0.77514
R6360 bgr_0.Vbe2.n140 bgr_0.Vbe2.n139 0.77514
R6361 bgr_0.Vbe2.n60 bgr_0.Vbe2 0.756696
R6362 bgr_0.Vbe2 bgr_0.Vbe2.n127 0.756696
R6363 bgr_0.Vbe2 bgr_0.Vbe2.n45 0.756696
R6364 bgr_0.Vbe2 bgr_0.Vbe2.n27 0.756696
R6365 bgr_0.Vbe2.n86 bgr_0.Vbe2 0.756696
R6366 bgr_0.Vbe2.n99 bgr_0.Vbe2 0.756696
R6367 bgr_0.Vbe2.n113 bgr_0.Vbe2 0.756696
R6368 bgr_0.Vbe2 bgr_0.Vbe2.n0 0.756696
R6369 bgr_0.Vbe2.n73 bgr_0.Vbe2.n72 0.711459
R6370 bgr_0.Vbe2.n149 bgr_0.Vbe2.n1 0.701365
R6371 bgr_0.Vbe2.n69 bgr_0.Vbe2.n36 0.647417
R6372 bgr_0.Vbe2.n116 bgr_0.Vbe2.n115 0.647417
R6373 bgr_0.Vbe2.n53 bgr_0.Vbe2.n52 0.590702
R6374 bgr_0.Vbe2.n40 bgr_0.Vbe2.n29 0.590702
R6375 bgr_0.Vbe2.n78 bgr_0.Vbe2.n25 0.590702
R6376 bgr_0.Vbe2.n91 bgr_0.Vbe2.n90 0.590702
R6377 bgr_0.Vbe2.n109 bgr_0.Vbe2.n12 0.590702
R6378 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 0.590702
R6379 bgr_0.Vbe2.n72 bgr_0.Vbe2 0.576566
R6380 bgr_0.Vbe2.n102 bgr_0.Vbe2.n14 0.530034
R6381 bgr_0.Vbe2.n124 bgr_0.Vbe2.n123 0.530034
R6382 bgr_0.Vbe2.n55 bgr_0.Vbe2.t0 0.290206
R6383 bgr_0.Vbe2.t4 bgr_0.Vbe2.n122 0.290206
R6384 bgr_0.Vbe2.n43 bgr_0.Vbe2.t2 0.290206
R6385 bgr_0.Vbe2.t3 bgr_0.Vbe2.n76 0.290206
R6386 bgr_0.Vbe2.n22 bgr_0.Vbe2.t1 0.290206
R6387 bgr_0.Vbe2.n17 bgr_0.Vbe2.t6 0.290206
R6388 bgr_0.Vbe2.n112 bgr_0.Vbe2.t5 0.290206
R6389 bgr_0.Vbe2.n141 bgr_0.Vbe2.t7 0.290206
R6390 bgr_0.Vbe2.n57 bgr_0.Vbe2 0.203382
R6391 bgr_0.Vbe2.n128 bgr_0.Vbe2 0.203382
R6392 bgr_0.Vbe2.n67 bgr_0.Vbe2 0.203382
R6393 bgr_0.Vbe2.n83 bgr_0.Vbe2 0.203382
R6394 bgr_0.Vbe2.n96 bgr_0.Vbe2 0.203382
R6395 bgr_0.Vbe2 bgr_0.Vbe2.n11 0.203382
R6396 bgr_0.Vbe2 bgr_0.Vbe2.n149 0.203382
R6397 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.154071
R6398 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 0.154071
R6399 bgr_0.Vbe2.n131 bgr_0.Vbe2.n130 0.154071
R6400 bgr_0.Vbe2.n147 bgr_0.Vbe2.n3 0.154071
R6401 bgr_0.Vbe2.n124 bgr_0.Vbe2.n121 0.137464
R6402 bgr_0.Vbe2.n64 bgr_0.Vbe2.n63 0.137464
R6403 bgr_0.Vbe2.n103 bgr_0.Vbe2.n102 0.134964
R6404 bgr_0.Vbe2.n71 bgr_0.Vbe2.n70 0.134964
R6405 bgr_0.Vbe2.n56 bgr_0.Vbe2 0.0196071
R6406 bgr_0.Vbe2.n101 bgr_0.Vbe2.n15 0.0183571
R6407 bgr_0.Vbe2.n95 bgr_0.Vbe2.n15 0.0183571
R6408 bgr_0.Vbe2.n94 bgr_0.Vbe2.n18 0.0183571
R6409 bgr_0.Vbe2.n89 bgr_0.Vbe2.n18 0.0183571
R6410 bgr_0.Vbe2.n89 bgr_0.Vbe2.n88 0.0183571
R6411 bgr_0.Vbe2.n88 bgr_0.Vbe2.n21 0.0183571
R6412 bgr_0.Vbe2.n82 bgr_0.Vbe2.n21 0.0183571
R6413 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 0.0183571
R6414 bgr_0.Vbe2.n80 bgr_0.Vbe2.n24 0.0183571
R6415 bgr_0.Vbe2.n125 bgr_0.Vbe2.n5 0.0183571
R6416 bgr_0.Vbe2.n130 bgr_0.Vbe2.n5 0.0183571
R6417 bgr_0.Vbe2.n135 bgr_0.Vbe2.n131 0.0183571
R6418 bgr_0.Vbe2.n137 bgr_0.Vbe2.n135 0.0183571
R6419 bgr_0.Vbe2.n148 bgr_0.Vbe2.n2 0.0183571
R6420 bgr_0.Vbe2.n148 bgr_0.Vbe2.n147 0.0183571
R6421 bgr_0.Vbe2.n50 bgr_0.Vbe2.n3 0.0183571
R6422 bgr_0.Vbe2.n50 bgr_0.Vbe2.n46 0.0183571
R6423 bgr_0.Vbe2.n62 bgr_0.Vbe2.n47 0.0183571
R6424 bgr_0.Vbe2.n56 bgr_0.Vbe2.n47 0.0183571
R6425 bgr_0.Vbe2.n71 bgr_0.Vbe2.n24 0.0106786
R6426 bgr_0.Vbe2.n63 bgr_0.Vbe2.n46 0.0106786
R6427 bgr_0.Vbe2.n136 bgr_0.Vbe2.n2 0.00996429
R6428 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 0.00992001
R6429 bgr_0.Vbe2.n119 bgr_0.Vbe2.n117 0.00992001
R6430 bgr_0.Vbe2.n118 bgr_0.Vbe2.n104 0.00992001
R6431 bgr_0.Vbe2.n106 bgr_0.Vbe2.n105 0.00992001
R6432 bgr_0.Vbe2.n121 bgr_0.Vbe2.n8 0.00992001
R6433 bgr_0.Vbe2.n105 bgr_0.Vbe2.n104 0.00992001
R6434 bgr_0.Vbe2.n106 bgr_0.Vbe2.n8 0.00992001
R6435 bgr_0.Vbe2.n117 bgr_0.Vbe2.n108 0.00992001
R6436 bgr_0.Vbe2.n107 bgr_0.Vbe2.n103 0.00992001
R6437 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 0.00992001
R6438 bgr_0.Vbe2.n33 bgr_0.Vbe2.n28 0.00992001
R6439 bgr_0.Vbe2.n66 bgr_0.Vbe2.n34 0.00992001
R6440 bgr_0.Vbe2.n68 bgr_0.Vbe2.n37 0.00992001
R6441 bgr_0.Vbe2.n65 bgr_0.Vbe2.n38 0.00992001
R6442 bgr_0.Vbe2.n64 bgr_0.Vbe2.n35 0.00992001
R6443 bgr_0.Vbe2.n68 bgr_0.Vbe2.n38 0.00992001
R6444 bgr_0.Vbe2.n65 bgr_0.Vbe2.n35 0.00992001
R6445 bgr_0.Vbe2.n34 bgr_0.Vbe2.n33 0.00992001
R6446 bgr_0.Vbe2.n70 bgr_0.Vbe2.n28 0.00992001
R6447 bgr_0.Vbe2.n66 bgr_0.Vbe2.n37 0.00992001
R6448 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 0.00889286
R6449 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 0.00817857
R6450 bgr_0.Vbe2.n73 bgr_0.Vbe2.n71 0.00817857
R6451 bgr_0.Vbe2.n125 bgr_0.Vbe2.n124 0.00817857
R6452 bgr_0.Vbe2.n63 bgr_0.Vbe2.n62 0.00817857
R6453 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t19 1172.87
R6454 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.t28 1172.87
R6455 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t38 996.134
R6456 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t27 996.134
R6457 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.t41 996.134
R6458 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t31 996.134
R6459 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t14 996.134
R6460 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t20 996.134
R6461 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t36 996.134
R6462 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t23 996.134
R6463 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t22 690.867
R6464 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t33 690.867
R6465 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t17 530.201
R6466 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t26 530.201
R6467 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t32 514.134
R6468 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t42 514.134
R6469 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t29 514.134
R6470 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t39 514.134
R6471 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t24 514.134
R6472 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t16 514.134
R6473 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t34 514.134
R6474 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t15 514.134
R6475 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t30 353.467
R6476 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.t13 353.467
R6477 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t18 353.467
R6478 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.t35 353.467
R6479 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t21 353.467
R6480 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6481 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t25 353.467
R6482 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t40 353.467
R6483 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6484 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.n31 176.733
R6485 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 176.733
R6486 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6487 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6488 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6489 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n17 176.733
R6490 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 176.733
R6491 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.n15 176.733
R6492 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 176.733
R6493 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n13 176.733
R6494 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.n12 176.733
R6495 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R6496 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6497 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6498 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.n23 176.733
R6499 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 176.733
R6500 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 176.733
R6501 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 166.436
R6502 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n19 161.843
R6503 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 161.718
R6504 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.n1 114.689
R6505 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n8 114.126
R6506 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.n6 114.126
R6507 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.n4 114.126
R6508 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.n2 114.126
R6509 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n0 109.626
R6510 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 51.9494
R6511 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n36 51.9494
R6512 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 51.9494
R6513 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n11 51.9494
R6514 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 51.9494
R6515 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n20 51.9494
R6516 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.X.n40 49.3036
R6517 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 18.4693
R6518 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.t12 16.0005
R6519 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.t2 16.0005
R6520 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.t6 16.0005
R6521 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.t7 16.0005
R6522 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.t9 16.0005
R6523 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R6524 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t0 16.0005
R6525 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t4 16.0005
R6526 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t10 16.0005
R6527 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t8 16.0005
R6528 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t5 16.0005
R6529 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t11 16.0005
R6530 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n10 9.28175
R6531 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 5.063
R6532 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n30 3.40675
R6533 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.n3 0.563
R6534 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.n5 0.563
R6535 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n7 0.563
R6536 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R6537 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R6538 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R6539 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 206.052
R6540 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 205.488
R6541 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 205.488
R6542 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 205.488
R6543 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 205.488
R6544 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 122.504
R6545 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 71.2813
R6546 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 54.5005
R6547 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R6548 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 39.4005
R6549 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R6550 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 39.4005
R6551 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 39.4005
R6552 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 39.4005
R6553 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R6554 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R6555 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R6556 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R6557 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 19.7005
R6558 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R6559 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 19.7005
R6560 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 19.7005
R6561 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R6562 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R6563 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 19.7005
R6564 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 6.09425
R6565 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 1.15675
R6566 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R6567 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R6568 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R6569 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t1 384.967
R6570 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t5 369.534
R6571 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t20 369.534
R6572 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t23 369.534
R6573 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t15 369.534
R6574 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t17 369.534
R6575 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.n18 369.534
R6576 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 365.491
R6577 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t12 192.8
R6578 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t11 192.8
R6579 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t19 192.8
R6580 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t6 192.8
R6581 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t14 192.8
R6582 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t13 192.8
R6583 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t21 192.8
R6584 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t7 192.8
R6585 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t16 192.8
R6586 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t22 192.8
R6587 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t9 192.8
R6588 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t10 192.8
R6589 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t18 192.8
R6590 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t8 192.8
R6591 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R6592 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R6593 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R6594 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R6595 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R6596 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R6597 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R6598 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R6599 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R6600 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R6601 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R6602 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R6603 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R6604 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R6605 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R6606 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R6607 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R6608 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R6609 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t3 39.4005
R6610 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t0 39.4005
R6611 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 28.6755
R6612 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t4 24.0005
R6613 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t2 24.0005
R6614 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R6615 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R6616 bgr_0.V_mir2.n4 bgr_0.V_mir2.n3 325.473
R6617 bgr_0.V_mir2.n16 bgr_0.V_mir2.t17 310.488
R6618 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R6619 bgr_0.V_mir2.n0 bgr_0.V_mir2.t20 310.488
R6620 bgr_0.V_mir2.n7 bgr_0.V_mir2.t15 278.312
R6621 bgr_0.V_mir2.n7 bgr_0.V_mir2.n6 228.939
R6622 bgr_0.V_mir2.n8 bgr_0.V_mir2.n5 224.439
R6623 bgr_0.V_mir2.n18 bgr_0.V_mir2.t4 184.097
R6624 bgr_0.V_mir2.n11 bgr_0.V_mir2.t8 184.097
R6625 bgr_0.V_mir2.n2 bgr_0.V_mir2.t6 184.097
R6626 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R6627 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R6628 bgr_0.V_mir2.n1 bgr_0.V_mir2.n0 167.094
R6629 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R6630 bgr_0.V_mir2.n4 bgr_0.V_mir2.n2 152
R6631 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R6632 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 120.501
R6633 bgr_0.V_mir2.n17 bgr_0.V_mir2.t12 120.501
R6634 bgr_0.V_mir2.n9 bgr_0.V_mir2.t19 120.501
R6635 bgr_0.V_mir2.n10 bgr_0.V_mir2.t10 120.501
R6636 bgr_0.V_mir2.n0 bgr_0.V_mir2.t18 120.501
R6637 bgr_0.V_mir2.n1 bgr_0.V_mir2.t2 120.501
R6638 bgr_0.V_mir2.n6 bgr_0.V_mir2.t14 48.0005
R6639 bgr_0.V_mir2.n6 bgr_0.V_mir2.t0 48.0005
R6640 bgr_0.V_mir2.n5 bgr_0.V_mir2.t16 48.0005
R6641 bgr_0.V_mir2.n5 bgr_0.V_mir2.t1 48.0005
R6642 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R6643 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R6644 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 40.7027
R6645 bgr_0.V_mir2.n12 bgr_0.V_mir2.t11 39.4005
R6646 bgr_0.V_mir2.n12 bgr_0.V_mir2.t9 39.4005
R6647 bgr_0.V_mir2.n3 bgr_0.V_mir2.t3 39.4005
R6648 bgr_0.V_mir2.n3 bgr_0.V_mir2.t7 39.4005
R6649 bgr_0.V_mir2.t13 bgr_0.V_mir2.n20 39.4005
R6650 bgr_0.V_mir2.n20 bgr_0.V_mir2.t5 39.4005
R6651 bgr_0.V_mir2.n15 bgr_0.V_mir2.n4 15.8005
R6652 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 15.8005
R6653 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 9.3005
R6654 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 5.8755
R6655 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R6656 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 0.78175
R6657 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6658 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 514.134
R6659 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 323.491
R6660 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 322.692
R6661 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6662 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6663 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 270.591
R6664 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 270.591
R6665 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 233.374
R6666 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 233.374
R6667 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 233.374
R6668 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 233.374
R6669 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 208.838
R6670 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 197.964
R6671 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 174.726
R6672 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 174.726
R6673 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 174.726
R6674 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6675 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 169.216
R6676 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 169.216
R6677 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 169.216
R6678 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 129.24
R6679 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 129.24
R6680 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6681 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6682 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 128.534
R6683 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 128.534
R6684 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 16.8443
R6685 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6686 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6687 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6688 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6689 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6690 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6691 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 4.3755
R6692 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 4.3755
R6693 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 3.688
R6694 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 3.1255
R6695 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 2.0005
R6696 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 1.2755
R6697 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 1.2755
R6698 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 0.8005
R6699 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 632.186
R6700 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 630.264
R6701 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6702 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6703 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 628.003
R6704 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 628.003
R6705 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 626.753
R6706 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 626.753
R6707 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 625.756
R6708 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 622.231
R6709 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6710 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6711 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6712 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6713 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6714 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6715 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6716 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6717 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6718 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6719 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6720 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6721 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6722 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6723 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6724 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6725 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6726 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6727 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6728 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6729 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 8.22272
R6730 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 6.188
R6731 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 630.264
R6732 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n2 627.316
R6733 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 626.784
R6734 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n3 626.784
R6735 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 626.784
R6736 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.n24 585
R6737 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6738 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6739 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.n21 176.733
R6740 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R6741 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6742 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6743 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6744 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6745 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6746 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6747 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6748 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6749 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6750 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6751 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6752 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6753 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6754 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6755 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n23 162.494
R6756 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 135.81
R6757 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n1 131.392
R6758 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6759 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6760 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6761 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6762 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6763 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6764 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6765 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6766 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6767 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6768 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6769 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6770 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6771 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6772 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6773 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6774 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6775 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6776 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6777 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6778 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R6779 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6780 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6781 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R6782 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6783 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6784 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6785 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6786 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6787 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R6788 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 49.8072
R6789 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n20 49.8072
R6790 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n25 41.7838
R6791 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6792 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t1 24.0005
R6793 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t0 24.0005
R6794 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 2.313
R6795 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t19 673.034
R6796 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 619.134
R6797 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t28 611.739
R6798 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t16 611.739
R6799 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R6800 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t31 611.739
R6801 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R6802 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R6803 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R6804 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t18 421.75
R6805 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R6806 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t12 421.75
R6807 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R6808 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t24 421.75
R6809 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t27 421.75
R6810 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R6811 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R6812 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R6813 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R6814 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R6815 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R6816 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R6817 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t0 288.166
R6818 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n10 169.311
R6819 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 168.936
R6820 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R6821 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R6822 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R6823 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R6824 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R6825 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R6826 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R6827 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R6828 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R6829 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R6830 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.n3 167.094
R6831 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R6832 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n23 140.547
R6833 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n26 140.546
R6834 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 139.297
R6835 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 139.297
R6836 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n22 109.312
R6837 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t8 62.5402
R6838 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t1 62.5402
R6839 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n18 47.1294
R6840 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n14 47.1294
R6841 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 47.1294
R6842 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n5 47.1294
R6843 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R6844 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R6845 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R6846 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R6847 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t10 24.0005
R6848 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R6849 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R6850 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R6851 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n1 18.0505
R6852 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 13.0943
R6853 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 5.6255
R6854 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 4.34425
R6855 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n25 3.71925
R6856 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 3.71925
R6857 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n4 4020
R6858 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n4 4020
R6859 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n10 4020
R6860 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n10 4020
R6861 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t30 660.109
R6862 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t27 660.109
R6863 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n14 428.8
R6864 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n3 428.8
R6865 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.VD3.n11 239.915
R6866 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.t28 239.915
R6867 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n8 230.4
R6868 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n6 230.4
R6869 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.n6 198.4
R6870 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n3 198.4
R6871 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 160.428
R6872 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n23 160.427
R6873 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 159.804
R6874 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.n19 159.803
R6875 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n21 159.803
R6876 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 159.802
R6877 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 159.802
R6878 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n28 159.802
R6879 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n26 159.802
R6880 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 159.802
R6881 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t32 155.125
R6882 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t29 155.125
R6883 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n16 146.002
R6884 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.VD3.t31 98.2764
R6885 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.t15 98.2764
R6886 two_stage_opamp_dummy_magic_0.VD3.t23 two_stage_opamp_dummy_magic_0.VD3.t19 98.2764
R6887 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.VD3.t23 98.2764
R6888 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.VD3.t7 98.2764
R6889 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t13 98.2764
R6890 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.VD3.t17 98.2764
R6891 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.VD3.t21 98.2764
R6892 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.VD3.t25 98.2764
R6893 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.VD3.t9 98.2764
R6894 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.n13 92.5005
R6895 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 92.5005
R6896 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n10 92.5005
R6897 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n3 92.5005
R6898 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n4 92.5005
R6899 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n4 92.5005
R6900 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t11 49.1384
R6901 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.VD3.n12 49.1384
R6902 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 21.3338
R6903 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 21.3338
R6904 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 19.2005
R6905 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.n17 13.8005
R6906 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t12 11.2576
R6907 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t14 11.2576
R6908 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.t18 11.2576
R6909 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R6910 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.t26 11.2576
R6911 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.t10 11.2576
R6912 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t36 11.2576
R6913 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t2 11.2576
R6914 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t4 11.2576
R6915 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R6916 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t35 11.2576
R6917 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t6 11.2576
R6918 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t34 11.2576
R6919 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R6920 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t33 11.2576
R6921 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t0 11.2576
R6922 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R6923 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R6924 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t16 11.2576
R6925 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R6926 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R6927 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t8 11.2576
R6928 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n33 8.3755
R6929 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n22 6.063
R6930 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n25 0.6255
R6931 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n27 0.6255
R6932 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n29 0.6255
R6933 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n31 0.6255
R6934 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.n18 0.6255
R6935 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R6936 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n20 0.5005
R6937 a_8420_8490.n8 a_8420_8490.n7 160.427
R6938 a_8420_8490.n2 a_8420_8490.n0 160.427
R6939 a_8420_8490.n6 a_8420_8490.n5 159.802
R6940 a_8420_8490.n4 a_8420_8490.n3 159.802
R6941 a_8420_8490.n2 a_8420_8490.n1 159.802
R6942 a_8420_8490.n9 a_8420_8490.n8 159.798
R6943 a_8420_8490.n7 a_8420_8490.t1 11.2576
R6944 a_8420_8490.n7 a_8420_8490.t10 11.2576
R6945 a_8420_8490.n5 a_8420_8490.t3 11.2576
R6946 a_8420_8490.n5 a_8420_8490.t5 11.2576
R6947 a_8420_8490.n3 a_8420_8490.t0 11.2576
R6948 a_8420_8490.n3 a_8420_8490.t2 11.2576
R6949 a_8420_8490.n1 a_8420_8490.t6 11.2576
R6950 a_8420_8490.n1 a_8420_8490.t8 11.2576
R6951 a_8420_8490.n0 a_8420_8490.t11 11.2576
R6952 a_8420_8490.n0 a_8420_8490.t4 11.2576
R6953 a_8420_8490.n9 a_8420_8490.t7 11.2576
R6954 a_8420_8490.t9 a_8420_8490.n9 11.2576
R6955 a_8420_8490.n4 a_8420_8490.n2 0.6255
R6956 a_8420_8490.n6 a_8420_8490.n4 0.6255
R6957 a_8420_8490.n8 a_8420_8490.n6 0.6255
R6958 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t17 1172.87
R6959 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t22 1172.87
R6960 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t39 996.134
R6961 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t27 996.134
R6962 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t14 996.134
R6963 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6964 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t13 996.134
R6965 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t31 996.134
R6966 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t37 996.134
R6967 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t24 996.134
R6968 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t20 690.867
R6969 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.t25 690.867
R6970 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t16 530.201
R6971 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.t21 530.201
R6972 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t34 514.134
R6973 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t18 514.134
R6974 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t35 514.134
R6975 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t19 514.134
R6976 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R6977 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t15 514.134
R6978 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t28 514.134
R6979 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.t40 514.134
R6980 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t29 353.467
R6981 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.t36 353.467
R6982 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t23 353.467
R6983 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t38 353.467
R6984 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t26 353.467
R6985 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t42 353.467
R6986 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t30 353.467
R6987 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R6988 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 176.733
R6989 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 176.733
R6990 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n15 176.733
R6991 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 176.733
R6992 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 176.733
R6993 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.n11 176.733
R6994 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.n21 176.733
R6995 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R6996 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6997 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6998 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6999 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R7000 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.n30 176.733
R7001 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R7002 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R7003 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R7004 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R7005 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R7006 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 166.436
R7007 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n29 161.843
R7008 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 161.718
R7009 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n1 114.689
R7010 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n8 114.126
R7011 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n6 114.126
R7012 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n4 114.126
R7013 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n2 114.126
R7014 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n0 109.626
R7015 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 51.9494
R7016 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n12 51.9494
R7017 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n28 51.9494
R7018 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n27 51.9494
R7019 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 51.9494
R7020 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n36 51.9494
R7021 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t6 49.3037
R7022 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 18.3443
R7023 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t0 16.0005
R7024 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R7025 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t2 16.0005
R7026 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t7 16.0005
R7027 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R7028 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t3 16.0005
R7029 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t12 16.0005
R7030 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R7031 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t8 16.0005
R7032 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t10 16.0005
R7033 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R7034 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R7035 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 7.6255
R7036 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 5.063
R7037 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n20 3.28175
R7038 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n10 1.71925
R7039 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n3 0.563
R7040 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n5 0.563
R7041 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n7 0.563
R7042 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n41 0.063
R7043 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n0 145.989
R7044 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n7 145.989
R7045 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.n5 145.427
R7046 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n3 145.427
R7047 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n1 145.427
R7048 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n9 140.927
R7049 two_stage_opamp_dummy_magic_0.VOUT+.t2 two_stage_opamp_dummy_magic_0.VOUT+.n96 113.192
R7050 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.n91 95.7303
R7051 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.n94 94.6053
R7052 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.n92 94.6053
R7053 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n10 20.688
R7054 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n89 11.7059
R7055 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.n90 10.438
R7056 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t12 6.56717
R7057 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t6 6.56717
R7058 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t10 6.56717
R7059 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t15 6.56717
R7060 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t11 6.56717
R7061 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t5 6.56717
R7062 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t3 6.56717
R7063 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t7 6.56717
R7064 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t4 6.56717
R7065 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t8 6.56717
R7066 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t14 6.56717
R7067 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t9 6.56717
R7068 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t108 4.8295
R7069 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t65 4.8295
R7070 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t118 4.8295
R7071 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t151 4.8295
R7072 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t44 4.8295
R7073 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t67 4.8295
R7074 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t27 4.8295
R7075 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t76 4.8295
R7076 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t62 4.8295
R7077 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t112 4.8295
R7078 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t114 4.8295
R7079 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t99 4.8295
R7080 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t74 4.8295
R7081 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t55 4.8295
R7082 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t109 4.8295
R7083 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t91 4.8295
R7084 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t68 4.8295
R7085 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t52 4.8295
R7086 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t29 4.8295
R7087 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t153 4.8295
R7088 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t63 4.8295
R7089 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t46 4.8295
R7090 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t22 4.8295
R7091 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t146 4.8295
R7092 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t117 4.8295
R7093 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.t72 4.8295
R7094 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t37 4.8295
R7095 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t20 4.8295
R7096 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t79 4.8295
R7097 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t60 4.8295
R7098 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t121 4.8295
R7099 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t104 4.8295
R7100 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t84 4.8295
R7101 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t66 4.8295
R7102 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t123 4.8295
R7103 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t95 4.8154
R7104 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t70 4.8154
R7105 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t110 4.8154
R7106 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t145 4.8154
R7107 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t32 4.806
R7108 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t150 4.806
R7109 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t50 4.806
R7110 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t87 4.806
R7111 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t125 4.806
R7112 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t105 4.806
R7113 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t140 4.806
R7114 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t36 4.806
R7115 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t156 4.806
R7116 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t53 4.806
R7117 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t73 4.806
R7118 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.t116 4.806
R7119 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t64 4.806
R7120 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t154 4.806
R7121 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t106 4.806
R7122 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t143 4.806
R7123 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t96 4.806
R7124 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t42 4.806
R7125 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t86 4.806
R7126 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t34 4.806
R7127 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t69 4.5005
R7128 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.t90 4.5005
R7129 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t80 4.5005
R7130 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.t43 4.5005
R7131 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t56 4.5005
R7132 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.t21 4.5005
R7133 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t98 4.5005
R7134 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.t59 4.5005
R7135 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t136 4.5005
R7136 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.t101 4.5005
R7137 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t30 4.5005
R7138 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.t51 4.5005
R7139 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t155 4.5005
R7140 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t119 4.5005
R7141 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t139 4.5005
R7142 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t102 4.5005
R7143 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t61 4.5005
R7144 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t85 4.5005
R7145 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t45 4.5005
R7146 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t147 4.5005
R7147 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t111 4.5005
R7148 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t134 4.5005
R7149 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t130 4.5005
R7150 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.t152 4.5005
R7151 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t115 4.5005
R7152 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t23 4.5005
R7153 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.t47 4.5005
R7154 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t148 4.5005
R7155 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t78 4.5005
R7156 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.t26 4.5005
R7157 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t132 4.5005
R7158 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t39 4.5005
R7159 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.t128 4.5005
R7160 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t92 4.5005
R7161 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t71 4.5005
R7162 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.t19 4.5005
R7163 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t126 4.5005
R7164 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t33 4.5005
R7165 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.t122 4.5005
R7166 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t88 4.5005
R7167 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t135 4.5005
R7168 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.t82 4.5005
R7169 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t48 4.5005
R7170 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t28 4.5005
R7171 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.t120 4.5005
R7172 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t81 4.5005
R7173 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t129 4.5005
R7174 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.t77 4.5005
R7175 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t40 4.5005
R7176 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t25 4.5005
R7177 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.t124 4.5005
R7178 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.t38 4.5005
R7179 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.t127 4.5005
R7180 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t94 4.5005
R7181 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t54 4.5005
R7182 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t144 4.5005
R7183 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t113 4.5005
R7184 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t75 4.5005
R7185 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t24 4.5005
R7186 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t131 4.5005
R7187 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t97 4.5005
R7188 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.t58 4.5005
R7189 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t149 4.5005
R7190 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t142 4.5005
R7191 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.t93 4.5005
R7192 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t57 4.5005
R7193 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t41 4.5005
R7194 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.t133 4.5005
R7195 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t100 4.5005
R7196 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t83 4.5005
R7197 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.t31 4.5005
R7198 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t137 4.5005
R7199 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t49 4.5005
R7200 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.t138 4.5005
R7201 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t103 4.5005
R7202 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t89 4.5005
R7203 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.t35 4.5005
R7204 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.t141 4.5005
R7205 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.t107 4.5005
R7206 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n8 4.5005
R7207 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.t17 3.42907
R7208 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.t18 3.42907
R7209 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.t0 3.42907
R7210 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.t13 3.42907
R7211 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t1 3.42907
R7212 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t16 3.42907
R7213 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.n95 2.03175
R7214 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.n93 1.1255
R7215 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n2 0.563
R7216 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.n4 0.563
R7217 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n6 0.563
R7218 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.n37 0.3295
R7219 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.n46 0.3295
R7220 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.n44 0.3295
R7221 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.n42 0.3295
R7222 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.n40 0.3295
R7223 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n39 0.3295
R7224 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n57 0.3295
R7225 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.n56 0.3295
R7226 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.n55 0.3295
R7227 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.n54 0.3295
R7228 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.n53 0.3295
R7229 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.n52 0.3295
R7230 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.n51 0.3295
R7231 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.n50 0.3295
R7232 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.n49 0.3295
R7233 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.n48 0.3295
R7234 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n59 0.3295
R7235 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n60 0.3295
R7236 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n62 0.3295
R7237 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n63 0.3295
R7238 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.n65 0.3295
R7239 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.n66 0.3295
R7240 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.n68 0.3295
R7241 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.n69 0.3295
R7242 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.n71 0.3295
R7243 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.n72 0.3295
R7244 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.n74 0.3295
R7245 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.n75 0.3295
R7246 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.n77 0.3295
R7247 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.n78 0.3295
R7248 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.n80 0.3295
R7249 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.n81 0.3295
R7250 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.n83 0.3295
R7251 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.n84 0.3295
R7252 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.n11 0.3295
R7253 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n13 0.3295
R7254 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n23 0.3295
R7255 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.n22 0.3295
R7256 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.n21 0.3295
R7257 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.n20 0.3295
R7258 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.n19 0.3295
R7259 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.n18 0.3295
R7260 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.n17 0.3295
R7261 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.n16 0.3295
R7262 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.n15 0.3295
R7263 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.n14 0.3295
R7264 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n25 0.3295
R7265 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n26 0.3295
R7266 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n28 0.3295
R7267 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n29 0.3295
R7268 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n31 0.3295
R7269 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n32 0.3295
R7270 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n34 0.3295
R7271 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n35 0.3295
R7272 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n86 0.3295
R7273 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.n87 0.3295
R7274 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.n88 0.3295
R7275 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.n47 0.306
R7276 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.n45 0.306
R7277 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.n43 0.306
R7278 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.n41 0.306
R7279 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n38 0.2825
R7280 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n58 0.2825
R7281 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n61 0.2825
R7282 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.n64 0.2825
R7283 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.n67 0.2825
R7284 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.n70 0.2825
R7285 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.n73 0.2825
R7286 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.n76 0.2825
R7287 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.n79 0.2825
R7288 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.n82 0.2825
R7289 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n12 0.2825
R7290 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n24 0.2825
R7291 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n27 0.2825
R7292 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n30 0.2825
R7293 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n33 0.2825
R7294 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n36 0.2825
R7295 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n85 0.2825
R7296 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t25 369.534
R7297 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t24 369.534
R7298 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t15 369.534
R7299 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t11 369.534
R7300 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t17 369.534
R7301 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t16 369.534
R7302 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7303 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7304 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7305 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7306 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t21 238.322
R7307 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t13 238.322
R7308 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t4 194.895
R7309 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t18 192.8
R7310 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t10 192.8
R7311 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t14 192.8
R7312 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t22 192.8
R7313 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t28 192.8
R7314 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t19 192.8
R7315 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t26 192.8
R7316 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t12 192.8
R7317 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t20 192.8
R7318 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t27 192.8
R7319 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t29 192.8
R7320 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t23 192.8
R7321 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7322 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7323 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7324 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7325 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7326 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7327 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7328 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 169.394
R7329 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7330 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7331 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t9 100.635
R7332 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7333 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7334 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7335 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7336 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7337 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7338 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t7 39.4005
R7339 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t3 39.4005
R7340 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t2 39.4005
R7341 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t0 39.4005
R7342 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t1 39.4005
R7343 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t5 39.4005
R7344 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t6 39.4005
R7345 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t8 39.4005
R7346 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 26.9067
R7347 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 5.15675
R7348 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7349 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n14 4.188
R7350 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 3.03175
R7351 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7352 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7353 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R7354 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 344.7
R7355 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R7356 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 206.052
R7357 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 205.488
R7358 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 205.488
R7359 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 205.488
R7360 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 205.488
R7361 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 122.474
R7362 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 83.3443
R7363 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 39.4005
R7364 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R7365 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 39.4005
R7366 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 39.4005
R7367 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 39.4005
R7368 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 39.4005
R7369 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 19.7005
R7370 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R7371 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 19.7005
R7372 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R7373 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R7374 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R7375 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R7376 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R7377 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R7378 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 19.7005
R7379 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 6.15675
R7380 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 6.1255
R7381 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R7382 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R7383 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R7384 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R7385 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 0.21925
R7386 a_14520_5068.t0 a_14520_5068.t1 294.339
R7387 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 144.827
R7388 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 134.577
R7389 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 120.629
R7390 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 114.501
R7391 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 97.4009
R7392 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 96.8384
R7393 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 96.8384
R7394 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 96.8384
R7395 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 96.8384
R7396 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 24.0005
R7397 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R7398 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R7399 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 24.0005
R7400 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R7401 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 8.0005
R7402 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R7403 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 8.0005
R7404 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R7405 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R7406 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R7407 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 8.0005
R7408 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R7409 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R7410 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 5.84425
R7411 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 1.46925
R7412 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 0.563
R7413 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 0.563
R7414 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 0.563
R7415 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7416 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7417 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7418 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 310.488
R7419 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7420 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7421 bgr_0.V_mir1.n7 bgr_0.V_mir1.t13 278.312
R7422 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7423 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7424 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R7425 bgr_0.V_mir1.n11 bgr_0.V_mir1.t0 184.097
R7426 bgr_0.V_mir1.n2 bgr_0.V_mir1.t8 184.097
R7427 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7428 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7429 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7430 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7431 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7432 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7433 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 120.501
R7434 bgr_0.V_mir1.n17 bgr_0.V_mir1.t2 120.501
R7435 bgr_0.V_mir1.n9 bgr_0.V_mir1.t18 120.501
R7436 bgr_0.V_mir1.n10 bgr_0.V_mir1.t4 120.501
R7437 bgr_0.V_mir1.n0 bgr_0.V_mir1.t17 120.501
R7438 bgr_0.V_mir1.n1 bgr_0.V_mir1.t6 120.501
R7439 bgr_0.V_mir1.n6 bgr_0.V_mir1.t12 48.0005
R7440 bgr_0.V_mir1.n6 bgr_0.V_mir1.t14 48.0005
R7441 bgr_0.V_mir1.n5 bgr_0.V_mir1.t15 48.0005
R7442 bgr_0.V_mir1.n5 bgr_0.V_mir1.t16 48.0005
R7443 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7444 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7445 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7446 bgr_0.V_mir1.n12 bgr_0.V_mir1.t1 39.4005
R7447 bgr_0.V_mir1.n12 bgr_0.V_mir1.t5 39.4005
R7448 bgr_0.V_mir1.n3 bgr_0.V_mir1.t9 39.4005
R7449 bgr_0.V_mir1.n3 bgr_0.V_mir1.t7 39.4005
R7450 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7451 bgr_0.V_mir1.n20 bgr_0.V_mir1.t3 39.4005
R7452 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7453 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7454 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7455 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7456 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7457 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7458 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 50.0055
R7459 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1603
R7460 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R7461 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1603
R7462 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R7463 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R7464 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1603
R7465 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1603
R7466 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R7467 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R7468 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R7469 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R7470 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R7471 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.1603
R7472 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.1603
R7473 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.1603
R7474 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R7475 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1603
R7476 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1603
R7477 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.1603
R7478 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R7479 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1603
R7480 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R7481 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.1603
R7482 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R7483 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1603
R7484 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R7485 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.1603
R7486 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.1603
R7487 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1603
R7488 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R7489 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R7490 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1603
R7491 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R7492 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1603
R7493 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1603
R7494 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1603
R7495 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R7496 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1603
R7497 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R7498 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R7499 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R7500 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1603
R7501 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R7502 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1603
R7503 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1603
R7504 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R7505 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.1603
R7506 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R7507 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1603
R7508 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1603
R7509 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1603
R7510 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R7511 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R7512 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1603
R7513 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1603
R7514 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R7515 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1603
R7516 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.1603
R7517 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.159278
R7518 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.159278
R7519 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.159278
R7520 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.159278
R7521 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.159278
R7522 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.159278
R7523 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.159278
R7524 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.159278
R7525 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.159278
R7526 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.159278
R7527 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.159278
R7528 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.159278
R7529 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.159278
R7530 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R7531 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R7532 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R7533 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7534 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7535 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7536 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7537 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7538 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7539 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7540 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.159278
R7541 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.159278
R7542 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.159278
R7543 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.159278
R7544 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.137822
R7545 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1368
R7546 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1368
R7547 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1368
R7548 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1368
R7549 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1368
R7550 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.1368
R7551 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.1368
R7552 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1368
R7553 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R7554 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1368
R7555 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1368
R7556 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.1368
R7557 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1368
R7558 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1368
R7559 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.1368
R7560 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1368
R7561 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1368
R7562 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7563 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.1368
R7564 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.1368
R7565 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1368
R7566 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.1368
R7567 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1368
R7568 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1368
R7569 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.1368
R7570 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R7571 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1368
R7572 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1368
R7573 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R7574 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1368
R7575 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.1368
R7576 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.114322
R7577 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.1133
R7578 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.1133
R7579 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7580 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7581 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7582 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7583 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7584 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7585 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7586 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7587 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7588 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7589 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7590 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7591 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.1133
R7592 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.1133
R7593 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.1133
R7594 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.1133
R7595 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R7596 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.00152174
R7597 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R7598 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.00152174
R7599 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.00152174
R7600 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.00152174
R7601 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.00152174
R7602 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.00152174
R7603 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R7604 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.00152174
R7605 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.00152174
R7606 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.00152174
R7607 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R7608 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.00152174
R7609 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.00152174
R7610 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.00152174
R7611 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.00152174
R7612 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.00152174
R7613 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.00152174
R7614 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.00152174
R7615 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.00152174
R7616 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R7617 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.00152174
R7618 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.00152174
R7619 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R7620 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.00152174
R7621 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.00152174
R7622 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.00152174
R7623 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R7624 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.00152174
R7625 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.00152174
R7626 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.00152174
R7627 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R7628 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.00152174
R7629 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R7630 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R7631 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R7632 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R7633 bgr_0.TAIL_CUR_MIR_BIAS.n17 bgr_0.TAIL_CUR_MIR_BIAS.t12 610.534
R7634 bgr_0.TAIL_CUR_MIR_BIAS.n8 bgr_0.TAIL_CUR_MIR_BIAS.t14 610.534
R7635 bgr_0.TAIL_CUR_MIR_BIAS.n17 bgr_0.TAIL_CUR_MIR_BIAS.t30 433.8
R7636 bgr_0.TAIL_CUR_MIR_BIAS.n18 bgr_0.TAIL_CUR_MIR_BIAS.t21 433.8
R7637 bgr_0.TAIL_CUR_MIR_BIAS.n19 bgr_0.TAIL_CUR_MIR_BIAS.t27 433.8
R7638 bgr_0.TAIL_CUR_MIR_BIAS.n20 bgr_0.TAIL_CUR_MIR_BIAS.t17 433.8
R7639 bgr_0.TAIL_CUR_MIR_BIAS.n21 bgr_0.TAIL_CUR_MIR_BIAS.t25 433.8
R7640 bgr_0.TAIL_CUR_MIR_BIAS.n22 bgr_0.TAIL_CUR_MIR_BIAS.t15 433.8
R7641 bgr_0.TAIL_CUR_MIR_BIAS.n23 bgr_0.TAIL_CUR_MIR_BIAS.t23 433.8
R7642 bgr_0.TAIL_CUR_MIR_BIAS.n24 bgr_0.TAIL_CUR_MIR_BIAS.t29 433.8
R7643 bgr_0.TAIL_CUR_MIR_BIAS.n25 bgr_0.TAIL_CUR_MIR_BIAS.t19 433.8
R7644 bgr_0.TAIL_CUR_MIR_BIAS.n16 bgr_0.TAIL_CUR_MIR_BIAS.t31 433.8
R7645 bgr_0.TAIL_CUR_MIR_BIAS.n15 bgr_0.TAIL_CUR_MIR_BIAS.t22 433.8
R7646 bgr_0.TAIL_CUR_MIR_BIAS.n14 bgr_0.TAIL_CUR_MIR_BIAS.t28 433.8
R7647 bgr_0.TAIL_CUR_MIR_BIAS.n13 bgr_0.TAIL_CUR_MIR_BIAS.t18 433.8
R7648 bgr_0.TAIL_CUR_MIR_BIAS.n12 bgr_0.TAIL_CUR_MIR_BIAS.t26 433.8
R7649 bgr_0.TAIL_CUR_MIR_BIAS.n11 bgr_0.TAIL_CUR_MIR_BIAS.t16 433.8
R7650 bgr_0.TAIL_CUR_MIR_BIAS.n10 bgr_0.TAIL_CUR_MIR_BIAS.t24 433.8
R7651 bgr_0.TAIL_CUR_MIR_BIAS.n9 bgr_0.TAIL_CUR_MIR_BIAS.t13 433.8
R7652 bgr_0.TAIL_CUR_MIR_BIAS.n8 bgr_0.TAIL_CUR_MIR_BIAS.t20 433.8
R7653 bgr_0.TAIL_CUR_MIR_BIAS.n3 bgr_0.TAIL_CUR_MIR_BIAS.n1 339.836
R7654 bgr_0.TAIL_CUR_MIR_BIAS.n5 bgr_0.TAIL_CUR_MIR_BIAS.n4 339.834
R7655 bgr_0.TAIL_CUR_MIR_BIAS.n3 bgr_0.TAIL_CUR_MIR_BIAS.n2 339.272
R7656 bgr_0.TAIL_CUR_MIR_BIAS.n6 bgr_0.TAIL_CUR_MIR_BIAS.n0 334.772
R7657 bgr_0.TAIL_CUR_MIR_BIAS.n28 bgr_0.TAIL_CUR_MIR_BIAS.n26 221.293
R7658 bgr_0.TAIL_CUR_MIR_BIAS.n25 bgr_0.TAIL_CUR_MIR_BIAS.n24 176.733
R7659 bgr_0.TAIL_CUR_MIR_BIAS.n24 bgr_0.TAIL_CUR_MIR_BIAS.n23 176.733
R7660 bgr_0.TAIL_CUR_MIR_BIAS.n23 bgr_0.TAIL_CUR_MIR_BIAS.n22 176.733
R7661 bgr_0.TAIL_CUR_MIR_BIAS.n22 bgr_0.TAIL_CUR_MIR_BIAS.n21 176.733
R7662 bgr_0.TAIL_CUR_MIR_BIAS.n21 bgr_0.TAIL_CUR_MIR_BIAS.n20 176.733
R7663 bgr_0.TAIL_CUR_MIR_BIAS.n20 bgr_0.TAIL_CUR_MIR_BIAS.n19 176.733
R7664 bgr_0.TAIL_CUR_MIR_BIAS.n19 bgr_0.TAIL_CUR_MIR_BIAS.n18 176.733
R7665 bgr_0.TAIL_CUR_MIR_BIAS.n18 bgr_0.TAIL_CUR_MIR_BIAS.n17 176.733
R7666 bgr_0.TAIL_CUR_MIR_BIAS.n9 bgr_0.TAIL_CUR_MIR_BIAS.n8 176.733
R7667 bgr_0.TAIL_CUR_MIR_BIAS.n10 bgr_0.TAIL_CUR_MIR_BIAS.n9 176.733
R7668 bgr_0.TAIL_CUR_MIR_BIAS.n11 bgr_0.TAIL_CUR_MIR_BIAS.n10 176.733
R7669 bgr_0.TAIL_CUR_MIR_BIAS.n12 bgr_0.TAIL_CUR_MIR_BIAS.n11 176.733
R7670 bgr_0.TAIL_CUR_MIR_BIAS.n13 bgr_0.TAIL_CUR_MIR_BIAS.n12 176.733
R7671 bgr_0.TAIL_CUR_MIR_BIAS.n14 bgr_0.TAIL_CUR_MIR_BIAS.n13 176.733
R7672 bgr_0.TAIL_CUR_MIR_BIAS.n15 bgr_0.TAIL_CUR_MIR_BIAS.n14 176.733
R7673 bgr_0.TAIL_CUR_MIR_BIAS.n16 bgr_0.TAIL_CUR_MIR_BIAS.n15 176.733
R7674 bgr_0.TAIL_CUR_MIR_BIAS.n29 bgr_0.TAIL_CUR_MIR_BIAS.n7 118.45
R7675 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.TAIL_CUR_MIR_BIAS.n29 86.7036
R7676 bgr_0.TAIL_CUR_MIR_BIAS.n29 bgr_0.TAIL_CUR_MIR_BIAS.n28 64.5795
R7677 bgr_0.TAIL_CUR_MIR_BIAS.n26 bgr_0.TAIL_CUR_MIR_BIAS.n25 56.2338
R7678 bgr_0.TAIL_CUR_MIR_BIAS.n26 bgr_0.TAIL_CUR_MIR_BIAS.n16 56.2338
R7679 bgr_0.TAIL_CUR_MIR_BIAS.n28 bgr_0.TAIL_CUR_MIR_BIAS.n27 53.2453
R7680 bgr_0.TAIL_CUR_MIR_BIAS.n0 bgr_0.TAIL_CUR_MIR_BIAS.t1 39.4005
R7681 bgr_0.TAIL_CUR_MIR_BIAS.n0 bgr_0.TAIL_CUR_MIR_BIAS.t6 39.4005
R7682 bgr_0.TAIL_CUR_MIR_BIAS.n4 bgr_0.TAIL_CUR_MIR_BIAS.t3 39.4005
R7683 bgr_0.TAIL_CUR_MIR_BIAS.n4 bgr_0.TAIL_CUR_MIR_BIAS.t0 39.4005
R7684 bgr_0.TAIL_CUR_MIR_BIAS.n1 bgr_0.TAIL_CUR_MIR_BIAS.t5 39.4005
R7685 bgr_0.TAIL_CUR_MIR_BIAS.n1 bgr_0.TAIL_CUR_MIR_BIAS.t2 39.4005
R7686 bgr_0.TAIL_CUR_MIR_BIAS.n2 bgr_0.TAIL_CUR_MIR_BIAS.t7 39.4005
R7687 bgr_0.TAIL_CUR_MIR_BIAS.n2 bgr_0.TAIL_CUR_MIR_BIAS.t4 39.4005
R7688 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.TAIL_CUR_MIR_BIAS.n6 18.3599
R7689 bgr_0.TAIL_CUR_MIR_BIAS.n27 bgr_0.TAIL_CUR_MIR_BIAS.t9 16.0005
R7690 bgr_0.TAIL_CUR_MIR_BIAS.n27 bgr_0.TAIL_CUR_MIR_BIAS.t11 16.0005
R7691 bgr_0.TAIL_CUR_MIR_BIAS.n7 bgr_0.TAIL_CUR_MIR_BIAS.t10 16.0005
R7692 bgr_0.TAIL_CUR_MIR_BIAS.n7 bgr_0.TAIL_CUR_MIR_BIAS.t8 16.0005
R7693 bgr_0.TAIL_CUR_MIR_BIAS.n6 bgr_0.TAIL_CUR_MIR_BIAS.n5 4.5005
R7694 bgr_0.TAIL_CUR_MIR_BIAS.n5 bgr_0.TAIL_CUR_MIR_BIAS.n3 0.563
R7695 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 219.928
R7696 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R7697 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R7698 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t1 9.6005
R7699 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R7700 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 229.562
R7701 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7702 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7703 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7704 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7705 bgr_0.V_p_2.n1 bgr_0.V_p_2.t6 98.2279
R7706 bgr_0.V_p_2.n5 bgr_0.V_p_2.t8 48.0005
R7707 bgr_0.V_p_2.n5 bgr_0.V_p_2.t4 48.0005
R7708 bgr_0.V_p_2.n4 bgr_0.V_p_2.t1 48.0005
R7709 bgr_0.V_p_2.n4 bgr_0.V_p_2.t9 48.0005
R7710 bgr_0.V_p_2.n3 bgr_0.V_p_2.t7 48.0005
R7711 bgr_0.V_p_2.n3 bgr_0.V_p_2.t3 48.0005
R7712 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R7713 bgr_0.V_p_2.n2 bgr_0.V_p_2.t0 48.0005
R7714 bgr_0.V_p_2.t5 bgr_0.V_p_2.n6 48.0005
R7715 bgr_0.V_p_2.n6 bgr_0.V_p_2.t10 48.0005
R7716 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7717 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7718 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7719 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7720 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7721 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7722 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7723 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7724 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7725 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7726 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7727 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7728 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7729 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7730 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7731 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7732 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7733 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7734 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7735 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7736 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7737 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7738 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7739 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7740 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7741 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7742 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7743 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7744 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7745 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7746 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7747 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7748 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7749 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7750 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7751 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7752 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.60845
R7753 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R7754 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R7755 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R7756 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7757 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7758 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R7759 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R7760 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R7761 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R7762 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 167.05
R7763 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R7764 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R7765 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R7766 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R7767 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R7768 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R7769 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R7770 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R7771 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R7772 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t1 117.591
R7773 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 117.591
R7774 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t2 108.424
R7775 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 108.424
R7776 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n0 35.9871
R7777 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 35.9246
R7778 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 10.6255
R7779 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 1.8755
R7780 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n4 1.31612
R7781 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.26612
R7782 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 1.15363
R7783 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7784 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7785 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t14 449.868
R7786 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t18 449.868
R7787 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R7788 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R7789 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7790 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7791 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7792 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R7793 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7794 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7795 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7796 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7797 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7798 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7799 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7800 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7801 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R7802 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7803 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7804 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7805 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t3 184.625
R7806 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R7807 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R7808 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R7809 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 176.733
R7810 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R7811 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7812 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R7813 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R7814 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R7815 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R7816 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R7817 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7818 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n11 170.269
R7819 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 165.8
R7820 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 99.2817
R7821 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t2 61.1914
R7822 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 56.2338
R7823 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n15 56.2338
R7824 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 56.2338
R7825 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n6 56.2338
R7826 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7827 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7828 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7829 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t1 39.4005
R7830 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n21 17.8599
R7831 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 14.3735
R7832 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 4.46925
R7833 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n7 114.719
R7834 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7835 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.n8 114.156
R7836 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7837 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7838 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7839 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7840 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7841 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7842 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7843 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7844 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7845 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7846 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7847 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7848 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7849 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7850 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7851 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7852 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7853 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7854 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7855 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7856 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7857 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7858 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7859 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7860 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7861 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7862 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7863 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7864 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7865 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7866 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7867 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7868 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7869 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7870 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7871 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7872 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 0.563
R7873 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7874 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7875 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 525.38
R7876 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 525.38
R7877 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 366.856
R7878 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 366.856
R7879 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 281.168
R7880 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 281.168
R7881 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 281.168
R7882 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 281.168
R7883 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7884 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7885 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7886 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7887 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7888 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7889 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7890 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7891 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 17.688
R7892 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7893 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7894 bgr_0.Vin+.n0 bgr_0.Vin+.t6 303.259
R7895 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R7896 bgr_0.Vin+.n0 bgr_0.Vin+.t8 174.726
R7897 bgr_0.Vin+.n1 bgr_0.Vin+.t10 174.726
R7898 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R7899 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R7900 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R7901 bgr_0.Vin+.n8 bgr_0.Vin+.t5 158.796
R7902 bgr_0.Vin+.t0 bgr_0.Vin+.n8 147.981
R7903 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7904 bgr_0.Vin+.n3 bgr_0.Vin+.t9 96.4005
R7905 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R7906 bgr_0.Vin+.n5 bgr_0.Vin+.t1 13.1338
R7907 bgr_0.Vin+.n5 bgr_0.Vin+.t4 13.1338
R7908 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R7909 bgr_0.Vin+.n4 bgr_0.Vin+.t2 13.1338
R7910 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R7911 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 229.562
R7912 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R7913 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R7914 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R7915 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R7916 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.2279
R7917 bgr_0.V_p_1.n5 bgr_0.V_p_1.t5 48.0005
R7918 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R7919 bgr_0.V_p_1.n4 bgr_0.V_p_1.t0 48.0005
R7920 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R7921 bgr_0.V_p_1.n3 bgr_0.V_p_1.t6 48.0005
R7922 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R7923 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R7924 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R7925 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R7926 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R7927 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R7928 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t13 355.293
R7929 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.t14 346.8
R7930 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.n20 339.522
R7931 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 339.522
R7932 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n14 335.022
R7933 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t10 275.909
R7934 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 227.909
R7935 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 222.034
R7936 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t26 184.097
R7937 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t36 184.097
R7938 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t19 184.097
R7939 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t32 184.097
R7940 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n17 166.05
R7941 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n8 166.05
R7942 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n4 57.7228
R7943 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t9 48.0005
R7944 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t8 48.0005
R7945 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t0 48.0005
R7946 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t7 48.0005
R7947 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t1 39.4005
R7948 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t4 39.4005
R7949 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t3 39.4005
R7950 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t5 39.4005
R7951 bgr_0.1st_Vout_2.t6 bgr_0.1st_Vout_2.n21 39.4005
R7952 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.t2 39.4005
R7953 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t17 4.8295
R7954 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t16 4.8295
R7955 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t27 4.8295
R7956 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t23 4.8295
R7957 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t35 4.8295
R7958 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t34 4.8295
R7959 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t28 4.8295
R7960 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R7961 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t15 4.5005
R7962 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t12 4.5005
R7963 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t30 4.5005
R7964 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t22 4.5005
R7965 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t18 4.5005
R7966 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t11 4.5005
R7967 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R7968 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t29 4.5005
R7969 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.5005
R7970 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t24 4.5005
R7971 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R7972 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.5005
R7973 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n11 4.5005
R7974 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n15 4.5005
R7975 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n7 1.3755
R7976 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n16 1.3755
R7977 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 1.188
R7978 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 0.9405
R7979 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n0 0.8935
R7980 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n13 0.78175
R7981 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 0.6585
R7982 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n3 0.6585
R7983 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n1 0.6585
R7984 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n9 0.6255
R7985 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n18 0.6255
R7986 bgr_0.cap_res2 bgr_0.cap_res2.t20 188.315
R7987 bgr_0.cap_res2 bgr_0.cap_res2.t9 0.259
R7988 bgr_0.cap_res2.t13 bgr_0.cap_res2.t8 0.1603
R7989 bgr_0.cap_res2.t2 bgr_0.cap_res2.t6 0.1603
R7990 bgr_0.cap_res2.t5 bgr_0.cap_res2.t1 0.1603
R7991 bgr_0.cap_res2.t19 bgr_0.cap_res2.t0 0.1603
R7992 bgr_0.cap_res2.t14 bgr_0.cap_res2.t10 0.1603
R7993 bgr_0.cap_res2.t4 bgr_0.cap_res2.t7 0.1603
R7994 bgr_0.cap_res2.t18 bgr_0.cap_res2.t16 0.1603
R7995 bgr_0.cap_res2.t12 bgr_0.cap_res2.t15 0.1603
R7996 bgr_0.cap_res2.n1 bgr_0.cap_res2.t17 0.159278
R7997 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.159278
R7998 bgr_0.cap_res2.n3 bgr_0.cap_res2.t3 0.159278
R7999 bgr_0.cap_res2.n3 bgr_0.cap_res2.t13 0.1368
R8000 bgr_0.cap_res2.n3 bgr_0.cap_res2.t2 0.1368
R8001 bgr_0.cap_res2.n2 bgr_0.cap_res2.t5 0.1368
R8002 bgr_0.cap_res2.n2 bgr_0.cap_res2.t19 0.1368
R8003 bgr_0.cap_res2.n1 bgr_0.cap_res2.t14 0.1368
R8004 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R8005 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R8006 bgr_0.cap_res2.n0 bgr_0.cap_res2.t12 0.1368
R8007 bgr_0.cap_res2.t17 bgr_0.cap_res2.n0 0.00152174
R8008 bgr_0.cap_res2.t11 bgr_0.cap_res2.n1 0.00152174
R8009 bgr_0.cap_res2.t3 bgr_0.cap_res2.n2 0.00152174
R8010 bgr_0.cap_res2.t9 bgr_0.cap_res2.n3 0.00152174
R8011 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.t31 206.407
R8012 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n26 118.168
R8013 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n19 117.831
R8014 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n33 117.269
R8015 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n31 117.269
R8016 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n29 117.269
R8017 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n27 117.269
R8018 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n24 117.269
R8019 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n22 117.269
R8020 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n20 117.269
R8021 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n18 113.136
R8022 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n3 99.647
R8023 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n0 99.5532
R8024 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n15 99.0845
R8025 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.n13 99.0845
R8026 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.n11 99.0845
R8027 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n6 99.0845
R8028 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n4 99.0845
R8029 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n1 99.0845
R8030 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.n37 94.5857
R8031 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.n8 94.5845
R8032 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.t35 16.0005
R8033 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.t27 16.0005
R8034 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t0 16.0005
R8035 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t1 16.0005
R8036 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t28 16.0005
R8037 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t25 16.0005
R8038 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t3 16.0005
R8039 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t32 16.0005
R8040 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t24 16.0005
R8041 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t26 16.0005
R8042 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t33 16.0005
R8043 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t37 16.0005
R8044 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t36 16.0005
R8045 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t2 16.0005
R8046 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t39 16.0005
R8047 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t40 16.0005
R8048 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t34 16.0005
R8049 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t30 16.0005
R8050 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.t5 16.0005
R8051 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.t29 16.0005
R8052 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t20 9.6005
R8053 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t10 9.6005
R8054 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t18 9.6005
R8055 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t8 9.6005
R8056 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.t14 9.6005
R8057 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.t6 9.6005
R8058 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t17 9.6005
R8059 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t7 9.6005
R8060 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t13 9.6005
R8061 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t21 9.6005
R8062 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t11 9.6005
R8063 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t19 9.6005
R8064 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t9 9.6005
R8065 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t15 9.6005
R8066 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t22 9.6005
R8067 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t16 9.6005
R8068 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t38 9.6005
R8069 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t4 9.6005
R8070 two_stage_opamp_dummy_magic_0.V_p.t23 two_stage_opamp_dummy_magic_0.V_p.n38 9.6005
R8071 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.t12 9.6005
R8072 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.n9 4.5005
R8073 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n35 4.5005
R8074 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n17 4.5005
R8075 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.n34 3.65675
R8076 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n36 1.28175
R8077 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n5 0.563
R8078 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.n7 0.563
R8079 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.n10 0.563
R8080 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.n12 0.563
R8081 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n14 0.563
R8082 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n16 0.563
R8083 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n2 0.563
R8084 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n28 0.563
R8085 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n30 0.563
R8086 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n32 0.563
R8087 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n21 0.563
R8088 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n23 0.563
R8089 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.n25 0.53175
R8090 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 144.827
R8091 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 134.577
R8092 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 120.66
R8093 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 98.063
R8094 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 97.4009
R8095 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 96.8384
R8096 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 96.8384
R8097 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 96.8384
R8098 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 96.8384
R8099 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 24.0005
R8100 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 24.0005
R8101 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 24.0005
R8102 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R8103 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R8104 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R8105 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R8106 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 8.0005
R8107 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R8108 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R8109 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R8110 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R8111 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R8112 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R8113 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 5.813
R8114 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 1.46925
R8115 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 0.563
R8116 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 0.563
R8117 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 0.563
R8118 VIN-.n4 VIN-.t8 485.021
R8119 VIN-.n1 VIN-.t6 484.159
R8120 VIN-.n5 VIN-.t7 483.358
R8121 VIN-.n8 VIN-.t10 431.536
R8122 VIN-.n2 VIN-.t9 431.536
R8123 VIN-.n6 VIN-.t1 431.257
R8124 VIN-.n0 VIN-.t0 431.257
R8125 VIN-.n6 VIN-.t2 289.908
R8126 VIN-.n0 VIN-.t5 289.908
R8127 VIN-.n8 VIN-.t4 279.183
R8128 VIN-.n2 VIN-.t3 279.183
R8129 VIN-.n7 VIN-.n6 233.374
R8130 VIN-.n1 VIN-.n0 233.374
R8131 VIN-.n9 VIN-.n8 188.989
R8132 VIN-.n3 VIN-.n2 188.989
R8133 VIN-.n4 VIN-.n3 2.463
R8134 VIN- VIN-.n9 2.03175
R8135 VIN-.n5 VIN-.n4 1.563
R8136 VIN-.n3 VIN-.n1 1.2755
R8137 VIN-.n9 VIN-.n7 1.2755
R8138 VIN-.n7 VIN-.n5 0.8005
R8139 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t12 668.604
R8140 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 631.982
R8141 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n3 627.128
R8142 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 627.128
R8143 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 226.534
R8144 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 226.534
R8145 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n4 222.034
R8146 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8147 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R8148 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R8149 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R8150 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t5 78.8005
R8151 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t4 78.8005
R8152 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R8153 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R8154 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R8155 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t11 48.0005
R8156 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R8157 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t10 48.0005
R8158 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 8.938
R8159 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 5.7505
R8160 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.313
R8161 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 1.2505
R8162 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.n23 4020
R8163 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n23 4020
R8164 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n24 4020
R8165 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.n24 4020
R8166 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.t0 660.109
R8167 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.t3 660.109
R8168 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n22 428.8
R8169 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n22 428.8
R8170 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.VD4.n28 239.915
R8171 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t1 239.915
R8172 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.n0 230.4
R8173 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n0 230.4
R8174 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 198.4
R8175 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 198.4
R8176 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n17 160.428
R8177 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.n2 160.427
R8178 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 159.803
R8179 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.n15 159.803
R8180 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n13 159.803
R8181 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 159.802
R8182 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n9 159.802
R8183 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 159.802
R8184 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 159.802
R8185 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.n3 159.802
R8186 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.t5 155.125
R8187 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.VD4.n33 155.125
R8188 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n1 146.002
R8189 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.VD4.t4 98.2764
R8190 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.VD4.t9 98.2764
R8191 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.VD4.t15 98.2764
R8192 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t23 98.2764
R8193 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.VD4.t19 98.2764
R8194 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.VD4.t27 98.2764
R8195 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t11 98.2764
R8196 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.t17 98.2764
R8197 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.t13 98.2764
R8198 two_stage_opamp_dummy_magic_0.VD4.t1 two_stage_opamp_dummy_magic_0.VD4.t21 98.2764
R8199 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.n27 92.5005
R8200 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.n22 92.5005
R8201 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n23 92.5005
R8202 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 92.5005
R8203 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.n0 92.5005
R8204 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n24 92.5005
R8205 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.t25 49.1384
R8206 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.VD4.n29 49.1384
R8207 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.n25 21.3338
R8208 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 21.3338
R8209 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 19.2005
R8210 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n12 14.438
R8211 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 13.8005
R8212 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t12 11.2576
R8213 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.t18 11.2576
R8214 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.t14 11.2576
R8215 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.t22 11.2576
R8216 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t24 11.2576
R8217 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.t20 11.2576
R8218 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R8219 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t16 11.2576
R8220 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.t32 11.2576
R8221 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.t36 11.2576
R8222 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t34 11.2576
R8223 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R8224 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R8225 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t37 11.2576
R8226 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R8227 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R8228 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.t33 11.2576
R8229 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8230 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t35 11.2576
R8231 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.t30 11.2576
R8232 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t26 11.2576
R8233 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t28 11.2576
R8234 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n19 0.6255
R8235 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n4 0.6255
R8236 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n6 0.6255
R8237 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n8 0.6255
R8238 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n10 0.6255
R8239 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n16 0.6255
R8240 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.n14 0.5005
R8241 a_10480_8490.n5 a_10480_8490.n3 160.427
R8242 a_10480_8490.n2 a_10480_8490.n0 160.427
R8243 a_10480_8490.n7 a_10480_8490.n6 159.802
R8244 a_10480_8490.n5 a_10480_8490.n4 159.802
R8245 a_10480_8490.n2 a_10480_8490.n1 159.802
R8246 a_10480_8490.n9 a_10480_8490.n8 159.798
R8247 a_10480_8490.n6 a_10480_8490.t11 11.2576
R8248 a_10480_8490.n6 a_10480_8490.t3 11.2576
R8249 a_10480_8490.n4 a_10480_8490.t6 11.2576
R8250 a_10480_8490.n4 a_10480_8490.t4 11.2576
R8251 a_10480_8490.n3 a_10480_8490.t8 11.2576
R8252 a_10480_8490.n3 a_10480_8490.t0 11.2576
R8253 a_10480_8490.n1 a_10480_8490.t5 11.2576
R8254 a_10480_8490.n1 a_10480_8490.t9 11.2576
R8255 a_10480_8490.n0 a_10480_8490.t1 11.2576
R8256 a_10480_8490.n0 a_10480_8490.t2 11.2576
R8257 a_10480_8490.n9 a_10480_8490.t7 11.2576
R8258 a_10480_8490.t10 a_10480_8490.n9 11.2576
R8259 a_10480_8490.n7 a_10480_8490.n5 0.6255
R8260 a_10480_8490.n8 a_10480_8490.n7 0.6255
R8261 a_10480_8490.n8 a_10480_8490.n2 0.6255
R8262 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.t20 619.201
R8263 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t12 611.739
R8264 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t25 611.739
R8265 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R8266 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t21 611.739
R8267 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R8268 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R8269 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R8270 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R8271 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R8272 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R8273 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R8274 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R8275 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R8276 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R8277 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t26 421.75
R8278 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R8279 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R8280 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R8281 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R8282 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R8283 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 176.155
R8284 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n13 175.79
R8285 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 172.667
R8286 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R8287 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R8288 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R8289 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R8290 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R8291 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R8292 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R8293 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R8294 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R8295 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R8296 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R8297 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R8298 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n1 139.639
R8299 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 139.638
R8300 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n0 134.577
R8301 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 106.891
R8302 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 47.1294
R8303 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n17 47.1294
R8304 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 47.1294
R8305 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n8 47.1294
R8306 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R8307 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R8308 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R8309 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R8310 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R8311 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R8312 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t6 10.9449
R8313 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t0 10.9449
R8314 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 9.5005
R8315 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n24 8.79738
R8316 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 4.5005
R8317 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 0.96925
R8318 a_11220_17410.t0 a_11220_17410.t1 258.591
R8319 a_5750_2276.t0 a_5750_2276.t1 169.905
R8320 a_14640_5068.t0 a_14640_5068.t1 169.905
R8321 VIN+.n9 VIN+.t5 485.127
R8322 VIN+.n4 VIN+.t3 485.127
R8323 VIN+.n3 VIN+.t4 485.127
R8324 VIN+.n7 VIN+.t9 318.656
R8325 VIN+.n7 VIN+.t2 318.656
R8326 VIN+.n5 VIN+.t7 318.656
R8327 VIN+.n5 VIN+.t1 318.656
R8328 VIN+.n1 VIN+.t8 318.656
R8329 VIN+.n1 VIN+.t6 318.656
R8330 VIN+.n0 VIN+.t10 318.656
R8331 VIN+.n0 VIN+.t0 318.656
R8332 VIN+.n2 VIN+.n0 167.05
R8333 VIN+.n8 VIN+.n7 165.8
R8334 VIN+.n6 VIN+.n5 165.8
R8335 VIN+.n2 VIN+.n1 165.8
R8336 VIN+.n6 VIN+.n4 2.34425
R8337 VIN+.n4 VIN+.n3 1.3005
R8338 VIN+.n8 VIN+.n6 1.2505
R8339 VIN+ VIN+.n9 1.213
R8340 VIN+.n3 VIN+.n2 1.15675
R8341 VIN+.n9 VIN+.n8 1.15675
R8342 a_13730_17020.t0 a_13730_17020.t1 258.591
R8343 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R8344 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R8345 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t3 303.259
R8346 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R8347 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R8348 bgr_0.V_CUR_REF_REG.t2 bgr_0.V_CUR_REF_REG.n5 245.284
R8349 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t7 174.726
R8350 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 174.726
R8351 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R8352 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R8353 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 96.4005
R8354 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t0 39.4005
R8355 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t1 39.4005
R8356 a_12828_17530.t0 a_12828_17530.t1 376.99
R8357 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8358 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8359 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8360 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8361 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8362 bgr_0.START_UP.n0 bgr_0.START_UP.t1 130.001
R8363 bgr_0.START_UP.n0 bgr_0.START_UP.t0 81.7074
R8364 bgr_0.START_UP bgr_0.START_UP.n0 38.2614
R8365 bgr_0.START_UP bgr_0.START_UP.n5 14.7817
R8366 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8367 bgr_0.START_UP.n1 bgr_0.START_UP.t3 13.1338
R8368 bgr_0.START_UP.n2 bgr_0.START_UP.t4 13.1338
R8369 bgr_0.START_UP.n2 bgr_0.START_UP.t5 13.1338
R8370 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8371 a_11220_17290.t0 a_11220_17290.t1 376.99
R8372 a_12828_17650.t0 a_12828_17650.t1 258.591
R8373 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8374 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2595
R8375 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2280
R8376 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2250
R8377 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 672.159
R8378 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 672.159
R8379 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 276.8
R8380 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 240
R8381 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 206.4
R8382 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 204.8
R8383 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 180.904
R8384 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 170.3
R8385 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 160.517
R8386 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 160.517
R8387 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 110.425
R8388 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 110.05
R8389 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 95.7988
R8390 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8391 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8392 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8393 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8394 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8395 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8396 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 76.8005
R8397 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 75.9449
R8398 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 75.9449
R8399 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 47.8997
R8400 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 47.8997
R8401 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 38.4005
R8402 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 24.5338
R8403 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 24.5338
R8404 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 16.8187
R8405 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 16.8187
R8406 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 12.313
R8407 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 12.313
R8408 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 10.9449
R8409 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 10.9449
R8410 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8411 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8412 a_5230_5088.t0 a_5230_5088.t1 294.339
R8413 a_14240_2276.t0 a_14240_2276.t1 169.905
R8414 a_13790_17550.t0 a_13790_17550.t1 258.591
R8415 a_5350_5088.t0 a_5350_5088.t1 169.905
C0 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.VD1 0.921543f
C1 VDDA two_stage_opamp_dummy_magic_0.VD3 4.36025f
C2 VDDA bgr_0.Vbe2 0.016701f
C3 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.err_amp_out 0.011225f
C4 VDDA two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.875085f
C5 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.551434f
C6 two_stage_opamp_dummy_magic_0.err_amp_out a_11120_2960# 0.012f
C7 bgr_0.1st_Vout_1 li_12710_16610# 0.020439f
C8 bgr_0.PFET_GATE_10uA m2_7180_19780# 0.012f
C9 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_gate 1.37399f
C10 li_7110_16510# VDDA 0.021911f
C11 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.318695f
C12 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 2.47368f
C13 bgr_0.V_TOP m2_8540_19780# 0.012f
C14 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.START_UP 2.09763f
C15 bgr_0.PFET_GATE_10uA bgr_0.1st_Vout_1 0.035393f
C16 bgr_0.1st_Vout_1 m2_8540_19780# 0.075543f
C17 bgr_0.PFET_GATE_10uA VDDA 10.3925f
C18 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.V_TOP 0.036996f
C19 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.VD3 0.036146f
C20 m2_8540_19780# VDDA 0.010446f
C21 bgr_0.NFET_GATE_10uA bgr_0.Vbe2 0.021455f
C22 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_gate 0.253351f
C23 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.528215f
C24 VIN- VIN+ 0.559567f
C25 bgr_0.TAIL_CUR_MIR_BIAS VDDA 5.87048f
C26 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.VD1 0.020203f
C27 bgr_0.cap_res2 bgr_0.1st_Vout_1 0.822981f
C28 bgr_0.cap_res2 VDDA 0.58582f
C29 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.VD1 1.05292f
C30 bgr_0.PFET_GATE_10uA bgr_0.NFET_GATE_10uA 0.050552f
C31 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.13839f
C32 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.err_amp_out 0.398657f
C33 bgr_0.V_TOP bgr_0.START_UP 0.815644f
C34 bgr_0.PFET_GATE_10uA bgr_0.Vbe2 0.242909f
C35 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.NFET_GATE_10uA 0.064423f
C36 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.cap_res_X 0.442088f
C37 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.1st_Vout_1 0.477103f
C38 bgr_0.TAIL_CUR_MIR_BIAS VIN- 0.315502f
C39 VDDA two_stage_opamp_dummy_magic_0.V_err_gate 5.03252f
C40 two_stage_opamp_dummy_magic_0.V_err_amp_ref VDDA 4.37237f
C41 bgr_0.cap_res2 li_10610_16720# 0.020538f
C42 bgr_0.1st_Vout_1 bgr_0.START_UP 0.030647f
C43 bgr_0.V_TOP li_5710_16610# 0.020062f
C44 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.VD3 0.397633f
C45 VDDA bgr_0.START_UP 1.37392f
C46 bgr_0.TAIL_CUR_MIR_BIAS VIN+ 0.111501f
C47 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.cap_res_X 0.048779f
C48 two_stage_opamp_dummy_magic_0.err_amp_out VDDA 1.20093f
C49 two_stage_opamp_dummy_magic_0.Y VDDA 3.98802f
C50 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 0.136183f
C51 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.NFET_GATE_10uA 0.559544f
C52 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.790473f
C53 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C54 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.PFET_GATE_10uA 0.213841f
C55 m2_7180_19780# VDDA 0.010446f
C56 bgr_0.NFET_GATE_10uA bgr_0.START_UP 0.518732f
C57 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.V_err_gate 0.013177f
C58 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.VD3 0.10263f
C59 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.Vbe2 0.014154f
C60 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.V_err_gate 0.065464f
C61 bgr_0.START_UP bgr_0.Vbe2 0.193132f
C62 bgr_0.V_TOP bgr_0.1st_Vout_1 0.925484f
C63 VIN- two_stage_opamp_dummy_magic_0.VD1 0.881219f
C64 bgr_0.TAIL_CUR_MIR_BIAS a_11120_2960# 0.012f
C65 bgr_0.V_TOP VDDA 16.1354f
C66 bgr_0.1st_Vout_1 VDDA 2.06087f
C67 bgr_0.cap_res2 bgr_0.PFET_GATE_10uA 0.018633f
C68 VIN+ two_stage_opamp_dummy_magic_0.VD1 0.057219f
C69 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.46518f
C70 bgr_0.PFET_GATE_10uA bgr_0.START_UP 0.166283f
C71 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_err_gate 0.039198f
C72 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_err_amp_ref 3.74826f
C73 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.080353f
C74 VDDA bgr_0.START_UP_NFET1 0.150608f
C75 bgr_0.1st_Vout_1 bgr_0.NFET_GATE_10uA 1.02268f
C76 bgr_0.V_TOP bgr_0.Vbe2 0.285619f
C77 VDDA bgr_0.NFET_GATE_10uA 1.04958f
C78 two_stage_opamp_dummy_magic_0.cap_res_X VDDA 0.921518f
C79 VOUT+ GNDA 0.038145f
C80 VOUT- GNDA 0.038151f
C81 VIN+ GNDA 2.09073f
C82 VIN- GNDA 2.163072f
C83 VDDA GNDA 0.150347p
C84 li_7110_16510# GNDA 0.050654f $ **FLOATING
C85 li_14110_16610# GNDA 0.050514f $ **FLOATING
C86 li_12710_16610# GNDA 0.049721f $ **FLOATING
C87 li_5710_16610# GNDA 0.047034f $ **FLOATING
C88 li_10610_16720# GNDA 0.049096f $ **FLOATING
C89 li_9210_16720# GNDA 0.043891f $ **FLOATING
C90 a_11120_2960# GNDA 0.110549f
C91 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.40894f
C92 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.718996f
C93 two_stage_opamp_dummy_magic_0.Y GNDA 5.187405f
C94 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 33.15933f
C95 bgr_0.cap_res2 GNDA 7.936877f
C96 bgr_0.TAIL_CUR_MIR_BIAS GNDA 10.99875f
C97 bgr_0.1st_Vout_1 GNDA 4.986571f
C98 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 15.223141f
C99 bgr_0.V_TOP GNDA 6.838887f
C100 bgr_0.PFET_GATE_10uA GNDA 5.13254f
C101 bgr_0.Vbe2 GNDA 17.0659f
C102 bgr_0.START_UP GNDA 7.190383f
C103 bgr_0.START_UP_NFET1 GNDA 5.28339f
C104 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 15.074302f
C105 bgr_0.NFET_GATE_10uA GNDA 7.08898f
C106 two_stage_opamp_dummy_magic_0.VD3 GNDA 6.496819f
C107 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.6041f
C108 bgr_0.START_UP.t0 GNDA 1.6623f
C109 bgr_0.START_UP.t1 GNDA 0.043697f
C110 bgr_0.START_UP.n0 GNDA 1.12862f
C111 bgr_0.START_UP.t2 GNDA 0.041701f
C112 bgr_0.START_UP.t3 GNDA 0.041701f
C113 bgr_0.START_UP.n1 GNDA 0.151283f
C114 bgr_0.START_UP.t4 GNDA 0.041701f
C115 bgr_0.START_UP.t5 GNDA 0.041701f
C116 bgr_0.START_UP.n2 GNDA 0.139173f
C117 bgr_0.START_UP.n3 GNDA 0.720787f
C118 bgr_0.START_UP.t7 GNDA 0.01567f
C119 bgr_0.START_UP.t6 GNDA 0.01567f
C120 bgr_0.START_UP.n4 GNDA 0.044238f
C121 bgr_0.START_UP.n5 GNDA 0.445182f
C122 bgr_0.V_CUR_REF_REG.t3 GNDA 0.014208f
C123 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C124 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C125 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C126 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C127 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C128 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C129 bgr_0.V_CUR_REF_REG.t2 GNDA 0.42777f
C130 VIN+.t0 GNDA 0.041803f
C131 VIN+.t10 GNDA 0.041803f
C132 VIN+.n0 GNDA 0.086391f
C133 VIN+.t6 GNDA 0.041803f
C134 VIN+.t8 GNDA 0.041803f
C135 VIN+.n1 GNDA 0.085194f
C136 VIN+.n2 GNDA 0.359761f
C137 VIN+.t4 GNDA 0.058811f
C138 VIN+.n3 GNDA 0.215335f
C139 VIN+.t3 GNDA 0.058811f
C140 VIN+.n4 GNDA 0.262589f
C141 VIN+.t1 GNDA 0.041803f
C142 VIN+.t7 GNDA 0.041803f
C143 VIN+.n5 GNDA 0.085194f
C144 VIN+.n6 GNDA 0.248358f
C145 VIN+.t2 GNDA 0.041803f
C146 VIN+.t9 GNDA 0.041803f
C147 VIN+.n7 GNDA 0.085194f
C148 VIN+.n8 GNDA 0.200956f
C149 VIN+.t5 GNDA 0.058811f
C150 VIN+.n9 GNDA 0.211601f
C151 bgr_0.VB3_CUR_BIAS GNDA 4.60549f
C152 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.031172f
C153 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.031172f
C154 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.094152f
C155 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.031172f
C156 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.031172f
C157 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.100408f
C158 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.031172f
C159 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.031172f
C160 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.100408f
C161 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.553544f
C162 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.206656f
C163 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.177535f
C164 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.154301f
C165 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.154301f
C166 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.154301f
C167 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.154301f
C168 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.178062f
C169 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.144567f
C170 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.08884f
C171 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.08884f
C172 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.083186f
C173 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.154301f
C174 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.154301f
C175 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.154301f
C176 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.154301f
C177 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.178062f
C178 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.144567f
C179 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.08884f
C180 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.08884f
C181 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.083186f
C182 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.086286f
C183 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.154301f
C184 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.154301f
C185 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.154301f
C186 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.154301f
C187 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.178062f
C188 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.144567f
C189 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.08884f
C190 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.08884f
C191 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.083186f
C192 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.154301f
C193 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.154301f
C194 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.154301f
C195 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.154301f
C196 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.178062f
C197 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.144567f
C198 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.08884f
C199 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.08884f
C200 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.083186f
C201 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.089524f
C202 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 2.44739f
C203 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.682611f
C204 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.112219f
C205 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.112219f
C206 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.401639f
C207 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 4.9401f
C208 a_10480_8490.t7 GNDA 0.066432f
C209 a_10480_8490.t1 GNDA 0.066432f
C210 a_10480_8490.t2 GNDA 0.066432f
C211 a_10480_8490.n0 GNDA 0.231036f
C212 a_10480_8490.t5 GNDA 0.066432f
C213 a_10480_8490.t9 GNDA 0.066432f
C214 a_10480_8490.n1 GNDA 0.230217f
C215 a_10480_8490.n2 GNDA 0.434626f
C216 a_10480_8490.t8 GNDA 0.066432f
C217 a_10480_8490.t0 GNDA 0.066432f
C218 a_10480_8490.n3 GNDA 0.231035f
C219 a_10480_8490.t6 GNDA 0.066432f
C220 a_10480_8490.t4 GNDA 0.066432f
C221 a_10480_8490.n4 GNDA 0.230217f
C222 a_10480_8490.n5 GNDA 0.434627f
C223 a_10480_8490.t11 GNDA 0.066432f
C224 a_10480_8490.t3 GNDA 0.066432f
C225 a_10480_8490.n6 GNDA 0.230217f
C226 a_10480_8490.n7 GNDA 0.225315f
C227 a_10480_8490.n8 GNDA 0.225315f
C228 a_10480_8490.n9 GNDA 0.230216f
C229 a_10480_8490.t10 GNDA 0.066432f
C230 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.053617f
C231 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.026064f
C232 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.026064f
C233 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.08498f
C234 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.026064f
C235 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.026064f
C236 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.090645f
C237 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.026064f
C238 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.026064f
C239 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.090324f
C240 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.170523f
C241 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.026064f
C242 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.026064f
C243 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.090324f
C244 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.088401f
C245 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.026064f
C246 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.026064f
C247 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.090324f
C248 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.088401f
C249 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.026064f
C250 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.026064f
C251 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.090324f
C252 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.088401f
C253 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.026064f
C254 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.026064f
C255 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.090324f
C256 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.168088f
C257 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.026064f
C258 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.026064f
C259 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.090324f
C260 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.162118f
C261 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.026064f
C262 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.026064f
C263 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.090324f
C264 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.085422f
C265 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.026064f
C266 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.026064f
C267 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.090645f
C268 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.026064f
C269 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.026064f
C270 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.090324f
C271 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.170523f
C272 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.03186f
C273 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.061885f
C274 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.103878f
C275 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.100899f
C276 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.100899f
C277 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.128579f
C278 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.045386f
C279 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.083882f
C280 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.054074f
C281 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.074201f
C282 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.300697f
C283 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.448835f
C284 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.259151f
C285 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.259151f
C286 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.259151f
C287 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.259151f
C288 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.194363f
C289 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.129575f
C290 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.194363f
C291 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.259151f
C292 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.259151f
C293 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.259151f
C294 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.259151f
C295 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.448835f
C296 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.300697f
C297 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.074201f
C298 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.054074f
C299 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.045386f
C300 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.083882f
C301 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.128579f
C302 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.017507f
C303 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.017316f
C304 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.345034f
C305 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.017316f
C306 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.019333f
C307 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.068944f
C308 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 0.020653f
C309 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 1.01255f
C310 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.020653f
C311 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.181418f
C312 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.176738f
C313 VIN-.t6 GNDA 0.050642f
C314 VIN-.t5 GNDA 0.033412f
C315 VIN-.t0 GNDA 0.041251f
C316 VIN-.n0 GNDA 0.059274f
C317 VIN-.n1 GNDA 0.280478f
C318 VIN-.t3 GNDA 0.032863f
C319 VIN-.t9 GNDA 0.041265f
C320 VIN-.n2 GNDA 0.064892f
C321 VIN-.n3 GNDA 0.200879f
C322 VIN-.t8 GNDA 0.050078f
C323 VIN-.n4 GNDA 0.236241f
C324 VIN-.t7 GNDA 0.050425f
C325 VIN-.n5 GNDA 0.180621f
C326 VIN-.t2 GNDA 0.033412f
C327 VIN-.t1 GNDA 0.041251f
C328 VIN-.n6 GNDA 0.059274f
C329 VIN-.n7 GNDA 0.149629f
C330 VIN-.t4 GNDA 0.032863f
C331 VIN-.t10 GNDA 0.041265f
C332 VIN-.n8 GNDA 0.064892f
C333 VIN-.n9 GNDA 0.186141f
C334 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.425414f
C335 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.102505f
C336 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.102505f
C337 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.423897f
C338 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.102505f
C339 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.102505f
C340 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.422271f
C341 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.585479f
C342 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.102505f
C343 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.102505f
C344 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.422271f
C345 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.305512f
C346 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.102505f
C347 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.102505f
C348 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.422271f
C349 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.305512f
C350 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.102505f
C351 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.102505f
C352 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.422271f
C353 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.439098f
C354 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 5.50033f
C355 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.034168f
C356 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.034168f
C357 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.124192f
C358 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.034168f
C359 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.034168f
C360 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.103202f
C361 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.645167f
C362 bgr_0.V_CMFB_S2 GNDA 4.4914f
C363 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA 0.024537f
C364 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA 0.024537f
C365 two_stage_opamp_dummy_magic_0.V_p.t4 GNDA 0.024537f
C366 two_stage_opamp_dummy_magic_0.V_p.n0 GNDA 0.097795f
C367 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA 0.024537f
C368 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA 0.024537f
C369 two_stage_opamp_dummy_magic_0.V_p.n1 GNDA 0.097424f
C370 two_stage_opamp_dummy_magic_0.V_p.n2 GNDA 0.164007f
C371 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA 0.024537f
C372 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA 0.024537f
C373 two_stage_opamp_dummy_magic_0.V_p.n3 GNDA 0.097877f
C374 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA 0.024537f
C375 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA 0.024537f
C376 two_stage_opamp_dummy_magic_0.V_p.n4 GNDA 0.097424f
C377 two_stage_opamp_dummy_magic_0.V_p.n5 GNDA 0.166869f
C378 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA 0.024537f
C379 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA 0.024537f
C380 two_stage_opamp_dummy_magic_0.V_p.n6 GNDA 0.097424f
C381 two_stage_opamp_dummy_magic_0.V_p.n7 GNDA 0.087096f
C382 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA 0.102522f
C383 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA 0.024537f
C384 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA 0.024537f
C385 two_stage_opamp_dummy_magic_0.V_p.n8 GNDA 0.094681f
C386 two_stage_opamp_dummy_magic_0.V_p.n9 GNDA 0.675343f
C387 two_stage_opamp_dummy_magic_0.V_p.n10 GNDA 0.029445f
C388 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA 0.024537f
C389 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA 0.024537f
C390 two_stage_opamp_dummy_magic_0.V_p.n11 GNDA 0.097424f
C391 two_stage_opamp_dummy_magic_0.V_p.n12 GNDA 0.087096f
C392 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA 0.024537f
C393 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA 0.024537f
C394 two_stage_opamp_dummy_magic_0.V_p.n13 GNDA 0.097424f
C395 two_stage_opamp_dummy_magic_0.V_p.n14 GNDA 0.087096f
C396 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA 0.024537f
C397 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA 0.024537f
C398 two_stage_opamp_dummy_magic_0.V_p.n15 GNDA 0.097424f
C399 two_stage_opamp_dummy_magic_0.V_p.n16 GNDA 0.087096f
C400 two_stage_opamp_dummy_magic_0.V_p.n17 GNDA 0.029445f
C401 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA 0.014722f
C402 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA 0.014722f
C403 two_stage_opamp_dummy_magic_0.V_p.n18 GNDA 0.050019f
C404 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA 0.014722f
C405 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA 0.014722f
C406 two_stage_opamp_dummy_magic_0.V_p.n19 GNDA 0.052892f
C407 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA 0.014722f
C408 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA 0.014722f
C409 two_stage_opamp_dummy_magic_0.V_p.n20 GNDA 0.052484f
C410 two_stage_opamp_dummy_magic_0.V_p.n21 GNDA 0.17749f
C411 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA 0.014722f
C412 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA 0.014722f
C413 two_stage_opamp_dummy_magic_0.V_p.n22 GNDA 0.052484f
C414 two_stage_opamp_dummy_magic_0.V_p.n23 GNDA 0.092385f
C415 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA 0.014722f
C416 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA 0.014722f
C417 two_stage_opamp_dummy_magic_0.V_p.n24 GNDA 0.052484f
C418 two_stage_opamp_dummy_magic_0.V_p.n25 GNDA 0.091894f
C419 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA 0.014722f
C420 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA 0.014722f
C421 two_stage_opamp_dummy_magic_0.V_p.n26 GNDA 0.052869f
C422 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA 0.014722f
C423 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA 0.014722f
C424 two_stage_opamp_dummy_magic_0.V_p.n27 GNDA 0.052484f
C425 two_stage_opamp_dummy_magic_0.V_p.n28 GNDA 0.175746f
C426 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA 0.014722f
C427 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA 0.014722f
C428 two_stage_opamp_dummy_magic_0.V_p.n29 GNDA 0.052484f
C429 two_stage_opamp_dummy_magic_0.V_p.n30 GNDA 0.092385f
C430 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA 0.014722f
C431 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA 0.014722f
C432 two_stage_opamp_dummy_magic_0.V_p.n31 GNDA 0.052484f
C433 two_stage_opamp_dummy_magic_0.V_p.n32 GNDA 0.092385f
C434 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA 0.014722f
C435 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA 0.014722f
C436 two_stage_opamp_dummy_magic_0.V_p.n33 GNDA 0.052484f
C437 two_stage_opamp_dummy_magic_0.V_p.n34 GNDA 0.140968f
C438 two_stage_opamp_dummy_magic_0.V_p.n35 GNDA 0.077538f
C439 two_stage_opamp_dummy_magic_0.V_p.n36 GNDA 0.082969f
C440 two_stage_opamp_dummy_magic_0.V_p.n37 GNDA 0.082287f
C441 two_stage_opamp_dummy_magic_0.V_p.n38 GNDA 0.094681f
C442 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA 0.024537f
C443 bgr_0.cap_res2.t6 GNDA 0.406156f
C444 bgr_0.cap_res2.t2 GNDA 0.407628f
C445 bgr_0.cap_res2.t8 GNDA 0.406156f
C446 bgr_0.cap_res2.t13 GNDA 0.407628f
C447 bgr_0.cap_res2.t0 GNDA 0.406156f
C448 bgr_0.cap_res2.t19 GNDA 0.407628f
C449 bgr_0.cap_res2.t1 GNDA 0.406156f
C450 bgr_0.cap_res2.t5 GNDA 0.407628f
C451 bgr_0.cap_res2.t7 GNDA 0.406156f
C452 bgr_0.cap_res2.t4 GNDA 0.407628f
C453 bgr_0.cap_res2.t10 GNDA 0.406156f
C454 bgr_0.cap_res2.t14 GNDA 0.407628f
C455 bgr_0.cap_res2.t15 GNDA 0.406156f
C456 bgr_0.cap_res2.t12 GNDA 0.407628f
C457 bgr_0.cap_res2.t16 GNDA 0.406156f
C458 bgr_0.cap_res2.t18 GNDA 0.407628f
C459 bgr_0.cap_res2.n0 GNDA 0.272247f
C460 bgr_0.cap_res2.t17 GNDA 0.216805f
C461 bgr_0.cap_res2.n1 GNDA 0.295394f
C462 bgr_0.cap_res2.t11 GNDA 0.216805f
C463 bgr_0.cap_res2.n2 GNDA 0.295394f
C464 bgr_0.cap_res2.t3 GNDA 0.216805f
C465 bgr_0.cap_res2.n3 GNDA 0.295394f
C466 bgr_0.cap_res2.t9 GNDA 0.214043f
C467 bgr_0.cap_res2.t20 GNDA 0.133038f
C468 bgr_0.1st_Vout_2.n0 GNDA 0.995956f
C469 bgr_0.1st_Vout_2.n1 GNDA 0.240335f
C470 bgr_0.1st_Vout_2.n2 GNDA 0.995956f
C471 bgr_0.1st_Vout_2.n3 GNDA 0.240335f
C472 bgr_0.1st_Vout_2.n4 GNDA 0.805677f
C473 bgr_0.1st_Vout_2.n5 GNDA 0.240335f
C474 bgr_0.1st_Vout_2.t13 GNDA 0.021508f
C475 bgr_0.1st_Vout_2.n6 GNDA 0.02259f
C476 bgr_0.1st_Vout_2.n7 GNDA 0.171874f
C477 bgr_0.1st_Vout_2.t32 GNDA 0.013652f
C478 bgr_0.1st_Vout_2.t19 GNDA 0.013652f
C479 bgr_0.1st_Vout_2.n8 GNDA 0.03037f
C480 bgr_0.1st_Vout_2.n9 GNDA 0.083918f
C481 bgr_0.1st_Vout_2.n10 GNDA 0.012945f
C482 bgr_0.1st_Vout_2.t10 GNDA 0.018875f
C483 bgr_0.1st_Vout_2.n11 GNDA 0.195802f
C484 bgr_0.1st_Vout_2.n12 GNDA 0.011712f
C485 bgr_0.1st_Vout_2.n13 GNDA 0.049674f
C486 bgr_0.1st_Vout_2.n14 GNDA 0.021654f
C487 bgr_0.1st_Vout_2.n15 GNDA 0.080059f
C488 bgr_0.1st_Vout_2.n16 GNDA 0.03943f
C489 bgr_0.1st_Vout_2.t36 GNDA 0.013652f
C490 bgr_0.1st_Vout_2.t26 GNDA 0.013652f
C491 bgr_0.1st_Vout_2.n17 GNDA 0.03037f
C492 bgr_0.1st_Vout_2.n18 GNDA 0.083918f
C493 bgr_0.1st_Vout_2.t17 GNDA 0.364565f
C494 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C495 bgr_0.1st_Vout_2.t15 GNDA 0.358459f
C496 bgr_0.1st_Vout_2.t16 GNDA 0.364565f
C497 bgr_0.1st_Vout_2.t12 GNDA 0.358459f
C498 bgr_0.1st_Vout_2.t27 GNDA 0.364565f
C499 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C500 bgr_0.1st_Vout_2.t22 GNDA 0.358459f
C501 bgr_0.1st_Vout_2.t23 GNDA 0.364565f
C502 bgr_0.1st_Vout_2.t18 GNDA 0.358459f
C503 bgr_0.1st_Vout_2.t35 GNDA 0.364565f
C504 bgr_0.1st_Vout_2.t11 GNDA 0.358459f
C505 bgr_0.1st_Vout_2.t31 GNDA 0.358459f
C506 bgr_0.1st_Vout_2.t34 GNDA 0.364565f
C507 bgr_0.1st_Vout_2.t29 GNDA 0.358459f
C508 bgr_0.1st_Vout_2.t28 GNDA 0.364565f
C509 bgr_0.1st_Vout_2.t33 GNDA 0.358459f
C510 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C511 bgr_0.1st_Vout_2.t20 GNDA 0.358459f
C512 bgr_0.1st_Vout_2.t25 GNDA 0.358459f
C513 bgr_0.1st_Vout_2.t14 GNDA 0.023417f
C514 bgr_0.1st_Vout_2.n19 GNDA 0.516024f
C515 bgr_0.1st_Vout_2.n20 GNDA 0.106455f
C516 bgr_0.1st_Vout_2.n21 GNDA 0.02259f
C517 bgr_0.Vin+.t6 GNDA 0.020459f
C518 bgr_0.Vin+.t8 GNDA 0.013299f
C519 bgr_0.Vin+.n0 GNDA 0.04388f
C520 bgr_0.Vin+.t10 GNDA 0.013299f
C521 bgr_0.Vin+.n1 GNDA 0.034146f
C522 bgr_0.Vin+.t7 GNDA 0.013299f
C523 bgr_0.Vin+.n2 GNDA 0.034607f
C524 bgr_0.Vin+.n3 GNDA 0.074523f
C525 bgr_0.Vin+.t3 GNDA 0.043132f
C526 bgr_0.Vin+.t2 GNDA 0.043132f
C527 bgr_0.Vin+.n4 GNDA 0.144858f
C528 bgr_0.Vin+.t1 GNDA 0.043132f
C529 bgr_0.Vin+.t4 GNDA 0.043132f
C530 bgr_0.Vin+.n5 GNDA 0.142495f
C531 bgr_0.Vin+.n6 GNDA 0.656763f
C532 bgr_0.Vin+.n7 GNDA 0.71769f
C533 bgr_0.Vin+.t5 GNDA 0.137433f
C534 bgr_0.Vin+.n8 GNDA 0.446219f
C535 bgr_0.Vin+.t0 GNDA 0.125873f
C536 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.174475f
C537 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.475245f
C538 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.435852f
C539 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.435852f
C540 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.517289f
C541 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.273228f
C542 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.17292f
C543 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.159805f
C544 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.805323f
C545 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.435852f
C546 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.435852f
C547 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.517289f
C548 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.273228f
C549 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.17292f
C550 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.475245f
C551 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.159805f
C552 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.805344f
C553 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.174475f
C554 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.175672f
C555 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.187155f
C556 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.175672f
C557 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.867885f
C558 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.041343f
C559 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.040593f
C560 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.225382f
C561 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.021075f
C562 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.123074f
C563 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.021216f
C564 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.034546f
C565 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.202018f
C566 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.040593f
C567 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.144283f
C568 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.160783f
C569 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 1.41037f
C570 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.867065f
C571 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.187134f
C572 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.021118f
C573 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020212f
C574 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020262f
C575 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021093f
C576 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.020966f
C577 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.297859f
C578 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.020966f
C579 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.155369f
C580 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.020966f
C581 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.189616f
C582 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.160506f
C583 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.14076f
C584 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.241198f
C585 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.021118f
C586 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020826f
C587 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.326026f
C588 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020826f
C589 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.179554f
C590 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.179554f
C591 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020826f
C592 bgr_0.TAIL_CUR_MIR_BIAS.t1 GNDA 0.03008f
C593 bgr_0.TAIL_CUR_MIR_BIAS.t6 GNDA 0.03008f
C594 bgr_0.TAIL_CUR_MIR_BIAS.n0 GNDA 0.072545f
C595 bgr_0.TAIL_CUR_MIR_BIAS.t5 GNDA 0.03008f
C596 bgr_0.TAIL_CUR_MIR_BIAS.t2 GNDA 0.03008f
C597 bgr_0.TAIL_CUR_MIR_BIAS.n1 GNDA 0.075298f
C598 bgr_0.TAIL_CUR_MIR_BIAS.t7 GNDA 0.03008f
C599 bgr_0.TAIL_CUR_MIR_BIAS.t4 GNDA 0.03008f
C600 bgr_0.TAIL_CUR_MIR_BIAS.n2 GNDA 0.074895f
C601 bgr_0.TAIL_CUR_MIR_BIAS.n3 GNDA 0.50855f
C602 bgr_0.TAIL_CUR_MIR_BIAS.t3 GNDA 0.03008f
C603 bgr_0.TAIL_CUR_MIR_BIAS.t0 GNDA 0.03008f
C604 bgr_0.TAIL_CUR_MIR_BIAS.n4 GNDA 0.075298f
C605 bgr_0.TAIL_CUR_MIR_BIAS.n5 GNDA 0.333784f
C606 bgr_0.TAIL_CUR_MIR_BIAS.n6 GNDA 0.774051f
C607 bgr_0.TAIL_CUR_MIR_BIAS.t10 GNDA 0.045119f
C608 bgr_0.TAIL_CUR_MIR_BIAS.t8 GNDA 0.045119f
C609 bgr_0.TAIL_CUR_MIR_BIAS.n7 GNDA 0.163283f
C610 bgr_0.TAIL_CUR_MIR_BIAS.t31 GNDA 0.080087f
C611 bgr_0.TAIL_CUR_MIR_BIAS.t22 GNDA 0.080087f
C612 bgr_0.TAIL_CUR_MIR_BIAS.t28 GNDA 0.080087f
C613 bgr_0.TAIL_CUR_MIR_BIAS.t18 GNDA 0.080087f
C614 bgr_0.TAIL_CUR_MIR_BIAS.t26 GNDA 0.080087f
C615 bgr_0.TAIL_CUR_MIR_BIAS.t16 GNDA 0.080087f
C616 bgr_0.TAIL_CUR_MIR_BIAS.t24 GNDA 0.080087f
C617 bgr_0.TAIL_CUR_MIR_BIAS.t13 GNDA 0.080087f
C618 bgr_0.TAIL_CUR_MIR_BIAS.t20 GNDA 0.080087f
C619 bgr_0.TAIL_CUR_MIR_BIAS.t14 GNDA 0.093474f
C620 bgr_0.TAIL_CUR_MIR_BIAS.n8 GNDA 0.088131f
C621 bgr_0.TAIL_CUR_MIR_BIAS.n9 GNDA 0.055271f
C622 bgr_0.TAIL_CUR_MIR_BIAS.n10 GNDA 0.055271f
C623 bgr_0.TAIL_CUR_MIR_BIAS.n11 GNDA 0.055271f
C624 bgr_0.TAIL_CUR_MIR_BIAS.n12 GNDA 0.055271f
C625 bgr_0.TAIL_CUR_MIR_BIAS.n13 GNDA 0.055271f
C626 bgr_0.TAIL_CUR_MIR_BIAS.n14 GNDA 0.055271f
C627 bgr_0.TAIL_CUR_MIR_BIAS.n15 GNDA 0.055271f
C628 bgr_0.TAIL_CUR_MIR_BIAS.n16 GNDA 0.04939f
C629 bgr_0.TAIL_CUR_MIR_BIAS.t19 GNDA 0.080087f
C630 bgr_0.TAIL_CUR_MIR_BIAS.t29 GNDA 0.080087f
C631 bgr_0.TAIL_CUR_MIR_BIAS.t23 GNDA 0.080087f
C632 bgr_0.TAIL_CUR_MIR_BIAS.t15 GNDA 0.080087f
C633 bgr_0.TAIL_CUR_MIR_BIAS.t25 GNDA 0.080087f
C634 bgr_0.TAIL_CUR_MIR_BIAS.t17 GNDA 0.080087f
C635 bgr_0.TAIL_CUR_MIR_BIAS.t27 GNDA 0.080087f
C636 bgr_0.TAIL_CUR_MIR_BIAS.t21 GNDA 0.080087f
C637 bgr_0.TAIL_CUR_MIR_BIAS.t30 GNDA 0.080087f
C638 bgr_0.TAIL_CUR_MIR_BIAS.t12 GNDA 0.093474f
C639 bgr_0.TAIL_CUR_MIR_BIAS.n17 GNDA 0.088131f
C640 bgr_0.TAIL_CUR_MIR_BIAS.n18 GNDA 0.055271f
C641 bgr_0.TAIL_CUR_MIR_BIAS.n19 GNDA 0.055271f
C642 bgr_0.TAIL_CUR_MIR_BIAS.n20 GNDA 0.055271f
C643 bgr_0.TAIL_CUR_MIR_BIAS.n21 GNDA 0.055271f
C644 bgr_0.TAIL_CUR_MIR_BIAS.n22 GNDA 0.055271f
C645 bgr_0.TAIL_CUR_MIR_BIAS.n23 GNDA 0.055271f
C646 bgr_0.TAIL_CUR_MIR_BIAS.n24 GNDA 0.055271f
C647 bgr_0.TAIL_CUR_MIR_BIAS.n25 GNDA 0.04939f
C648 bgr_0.TAIL_CUR_MIR_BIAS.n26 GNDA 0.12343f
C649 bgr_0.TAIL_CUR_MIR_BIAS.t9 GNDA 0.045119f
C650 bgr_0.TAIL_CUR_MIR_BIAS.t11 GNDA 0.045119f
C651 bgr_0.TAIL_CUR_MIR_BIAS.n27 GNDA 0.090239f
C652 bgr_0.TAIL_CUR_MIR_BIAS.n28 GNDA 0.349784f
C653 bgr_0.TAIL_CUR_MIR_BIAS.n29 GNDA 3.57484f
C654 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.344645f
C655 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.345894f
C656 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.344645f
C657 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.347347f
C658 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.37779f
C659 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.344645f
C660 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.345894f
C661 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.344645f
C662 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.345894f
C663 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.344645f
C664 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.345894f
C665 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.344645f
C666 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.345894f
C667 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.344645f
C668 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.345894f
C669 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.344645f
C670 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.345894f
C671 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.344645f
C672 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.345894f
C673 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.344645f
C674 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.345894f
C675 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.344645f
C676 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.345894f
C677 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.344645f
C678 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.345894f
C679 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.344645f
C680 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.345894f
C681 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.344645f
C682 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.345894f
C683 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.344645f
C684 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.345894f
C685 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.344645f
C686 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.345894f
C687 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.344645f
C688 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.345894f
C689 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.344645f
C690 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.345894f
C691 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.344645f
C692 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.345894f
C693 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.344645f
C694 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.345894f
C695 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.344645f
C696 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.345894f
C697 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.344645f
C698 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.345894f
C699 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.344645f
C700 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.345894f
C701 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.344645f
C702 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.345894f
C703 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.344645f
C704 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.345894f
C705 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.344645f
C706 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.345894f
C707 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.344645f
C708 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.345894f
C709 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.344645f
C710 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.345894f
C711 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.344645f
C712 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.345894f
C713 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.344645f
C714 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.345894f
C715 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.344645f
C716 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.345894f
C717 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.344645f
C718 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.361543f
C719 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.344645f
C720 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.185116f
C721 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.19812f
C722 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.344645f
C723 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.185116f
C724 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.196522f
C725 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.344645f
C726 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.185116f
C727 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.196522f
C728 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.344645f
C729 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.185116f
C730 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.196522f
C731 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.344645f
C732 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.185116f
C733 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.196522f
C734 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.344645f
C735 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.185116f
C736 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.196522f
C737 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.344645f
C738 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.185116f
C739 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.196522f
C740 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.344645f
C741 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.185116f
C742 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196522f
C743 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.344645f
C744 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.185116f
C745 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196522f
C746 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.344645f
C747 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.345894f
C748 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.166619f
C749 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.214914f
C750 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.18397f
C751 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.23341f
C752 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.18397f
C753 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.250658f
C754 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.18397f
C755 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.250658f
C756 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.18397f
C757 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.250658f
C758 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.18397f
C759 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.250658f
C760 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.18397f
C761 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.250658f
C762 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.18397f
C763 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.250658f
C764 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.18397f
C765 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250658f
C766 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.18397f
C767 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250658f
C768 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.18397f
C769 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250658f
C770 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.18397f
C771 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250658f
C772 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.18397f
C773 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250658f
C774 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.18397f
C775 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250658f
C776 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.18397f
C777 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250658f
C778 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.18397f
C779 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250658f
C780 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.18397f
C781 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.23341f
C782 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.343499f
C783 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.166619f
C784 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.216163f
C785 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.343499f
C786 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.166619f
C787 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.216163f
C788 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.343499f
C789 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.344645f
C790 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.363141f
C791 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.363141f
C792 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.185116f
C793 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.216163f
C794 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.343499f
C795 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.344645f
C796 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.185116f
C797 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.197667f
C798 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.343499f
C799 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.344645f
C800 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.185116f
C801 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.216163f
C802 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.343499f
C803 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.344645f
C804 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.185116f
C805 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.216163f
C806 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.343499f
C807 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.344645f
C808 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.185116f
C809 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216163f
C810 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.343499f
C811 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.344645f
C812 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.363141f
C813 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.363141f
C814 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.185116f
C815 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216163f
C816 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.343499f
C817 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.344645f
C818 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.363141f
C819 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.363141f
C820 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.185116f
C821 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216163f
C822 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.343499f
C823 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216163f
C824 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.185116f
C825 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.363141f
C826 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.363141f
C827 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.764814f
C828 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.3034f
C829 bgr_0.V_mir1.t8 GNDA 0.053881f
C830 bgr_0.V_mir1.t6 GNDA 0.042444f
C831 bgr_0.V_mir1.t17 GNDA 0.042444f
C832 bgr_0.V_mir1.t20 GNDA 0.06851f
C833 bgr_0.V_mir1.n0 GNDA 0.076506f
C834 bgr_0.V_mir1.n1 GNDA 0.052264f
C835 bgr_0.V_mir1.n2 GNDA 0.081315f
C836 bgr_0.V_mir1.t9 GNDA 0.03537f
C837 bgr_0.V_mir1.t7 GNDA 0.03537f
C838 bgr_0.V_mir1.n3 GNDA 0.08097f
C839 bgr_0.V_mir1.n4 GNDA 0.203577f
C840 bgr_0.V_mir1.t15 GNDA 0.017685f
C841 bgr_0.V_mir1.t16 GNDA 0.017685f
C842 bgr_0.V_mir1.n5 GNDA 0.046242f
C843 bgr_0.V_mir1.t13 GNDA 0.075466f
C844 bgr_0.V_mir1.t12 GNDA 0.017685f
C845 bgr_0.V_mir1.t14 GNDA 0.017685f
C846 bgr_0.V_mir1.n6 GNDA 0.050199f
C847 bgr_0.V_mir1.n7 GNDA 0.827814f
C848 bgr_0.V_mir1.n8 GNDA 0.268286f
C849 bgr_0.V_mir1.t0 GNDA 0.053881f
C850 bgr_0.V_mir1.t4 GNDA 0.042444f
C851 bgr_0.V_mir1.t18 GNDA 0.042444f
C852 bgr_0.V_mir1.t21 GNDA 0.06851f
C853 bgr_0.V_mir1.n9 GNDA 0.076506f
C854 bgr_0.V_mir1.n10 GNDA 0.052264f
C855 bgr_0.V_mir1.n11 GNDA 0.081315f
C856 bgr_0.V_mir1.t1 GNDA 0.03537f
C857 bgr_0.V_mir1.t5 GNDA 0.03537f
C858 bgr_0.V_mir1.n12 GNDA 0.08097f
C859 bgr_0.V_mir1.n13 GNDA 0.156007f
C860 bgr_0.V_mir1.n14 GNDA 0.09373f
C861 bgr_0.V_mir1.n15 GNDA 0.699157f
C862 bgr_0.V_mir1.t10 GNDA 0.053881f
C863 bgr_0.V_mir1.t2 GNDA 0.042444f
C864 bgr_0.V_mir1.t19 GNDA 0.042444f
C865 bgr_0.V_mir1.t22 GNDA 0.06851f
C866 bgr_0.V_mir1.n16 GNDA 0.076506f
C867 bgr_0.V_mir1.n17 GNDA 0.052264f
C868 bgr_0.V_mir1.n18 GNDA 0.081315f
C869 bgr_0.V_mir1.n19 GNDA 0.201563f
C870 bgr_0.V_mir1.t3 GNDA 0.03537f
C871 bgr_0.V_mir1.n20 GNDA 0.08097f
C872 bgr_0.V_mir1.t11 GNDA 0.03537f
C873 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.477162f
C874 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.115051f
C875 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.115051f
C876 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.47578f
C877 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.115051f
C878 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.115051f
C879 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.473954f
C880 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.657139f
C881 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.115051f
C882 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.115051f
C883 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.473954f
C884 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.342905f
C885 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.115051f
C886 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.115051f
C887 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.473954f
C888 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.342905f
C889 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.115051f
C890 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.115051f
C891 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.473954f
C892 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.49568f
C893 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 7.289f
C894 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.03835f
C895 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.03835f
C896 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.139392f
C897 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.03835f
C898 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.03835f
C899 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.115834f
C900 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.724132f
C901 bgr_0.V_CMFB_S4 GNDA 5.94035f
C902 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.033671f
C903 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.033671f
C904 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.084438f
C905 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.033671f
C906 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.033671f
C907 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.083993f
C908 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.568968f
C909 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.033671f
C910 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.033671f
C911 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.083993f
C912 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.597848f
C913 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.430908f
C914 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.067342f
C915 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.067342f
C916 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.19758f
C917 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.067342f
C918 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.067342f
C919 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.196683f
C920 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.679849f
C921 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.067342f
C922 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.067342f
C923 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.196683f
C924 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.352158f
C925 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.067342f
C926 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.067342f
C927 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.196683f
C928 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.352158f
C929 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.067342f
C930 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.067342f
C931 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.196683f
C932 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.508351f
C933 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 5.05557f
C934 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 GNDA 4.02733f
C935 bgr_0.V_CMFB_S3 GNDA 0.014671f
C936 bgr_0.PFET_GATE_10uA.t23 GNDA 0.039179f
C937 bgr_0.PFET_GATE_10uA.t16 GNDA 0.057916f
C938 bgr_0.PFET_GATE_10uA.n0 GNDA 0.063817f
C939 bgr_0.PFET_GATE_10uA.t29 GNDA 0.039179f
C940 bgr_0.PFET_GATE_10uA.t17 GNDA 0.057916f
C941 bgr_0.PFET_GATE_10uA.n1 GNDA 0.063817f
C942 bgr_0.PFET_GATE_10uA.n2 GNDA 0.076791f
C943 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039179f
C944 bgr_0.PFET_GATE_10uA.t24 GNDA 0.057916f
C945 bgr_0.PFET_GATE_10uA.n3 GNDA 0.063817f
C946 bgr_0.PFET_GATE_10uA.t18 GNDA 0.039179f
C947 bgr_0.PFET_GATE_10uA.t25 GNDA 0.057916f
C948 bgr_0.PFET_GATE_10uA.n4 GNDA 0.063817f
C949 bgr_0.PFET_GATE_10uA.n5 GNDA 0.064022f
C950 bgr_0.PFET_GATE_10uA.t4 GNDA 0.781422f
C951 bgr_0.PFET_GATE_10uA.t9 GNDA 0.586977f
C952 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040183f
C953 bgr_0.PFET_GATE_10uA.t8 GNDA 0.040183f
C954 bgr_0.PFET_GATE_10uA.n6 GNDA 0.102705f
C955 bgr_0.PFET_GATE_10uA.t1 GNDA 0.040183f
C956 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040183f
C957 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100051f
C958 bgr_0.PFET_GATE_10uA.n8 GNDA 0.978629f
C959 bgr_0.PFET_GATE_10uA.t2 GNDA 0.040183f
C960 bgr_0.PFET_GATE_10uA.t0 GNDA 0.040183f
C961 bgr_0.PFET_GATE_10uA.n9 GNDA 0.100051f
C962 bgr_0.PFET_GATE_10uA.n10 GNDA 0.554934f
C963 bgr_0.PFET_GATE_10uA.n11 GNDA 1.13286f
C964 bgr_0.PFET_GATE_10uA.t7 GNDA 0.040183f
C965 bgr_0.PFET_GATE_10uA.t3 GNDA 0.040183f
C966 bgr_0.PFET_GATE_10uA.n12 GNDA 0.096913f
C967 bgr_0.PFET_GATE_10uA.n13 GNDA 0.356682f
C968 bgr_0.PFET_GATE_10uA.n14 GNDA 3.84996f
C969 bgr_0.PFET_GATE_10uA.t13 GNDA 0.045299f
C970 bgr_0.PFET_GATE_10uA.t21 GNDA 0.045299f
C971 bgr_0.PFET_GATE_10uA.n15 GNDA 0.137138f
C972 bgr_0.PFET_GATE_10uA.n16 GNDA 1.78858f
C973 bgr_0.PFET_GATE_10uA.n17 GNDA 1.41725f
C974 bgr_0.PFET_GATE_10uA.t27 GNDA 0.039179f
C975 bgr_0.PFET_GATE_10uA.t20 GNDA 0.039179f
C976 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039179f
C977 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039179f
C978 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039179f
C979 bgr_0.PFET_GATE_10uA.t11 GNDA 0.057916f
C980 bgr_0.PFET_GATE_10uA.n18 GNDA 0.071675f
C981 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051234f
C982 bgr_0.PFET_GATE_10uA.n20 GNDA 0.051234f
C983 bgr_0.PFET_GATE_10uA.n21 GNDA 0.051234f
C984 bgr_0.PFET_GATE_10uA.n22 GNDA 0.043376f
C985 bgr_0.PFET_GATE_10uA.t14 GNDA 0.039179f
C986 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039179f
C987 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039179f
C988 bgr_0.PFET_GATE_10uA.t15 GNDA 0.057916f
C989 bgr_0.PFET_GATE_10uA.n23 GNDA 0.071675f
C990 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051234f
C991 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043376f
C992 bgr_0.PFET_GATE_10uA.n26 GNDA 0.05954f
C993 two_stage_opamp_dummy_magic_0.VOUT+.t14 GNDA 0.043632f
C994 two_stage_opamp_dummy_magic_0.VOUT+.t9 GNDA 0.043632f
C995 two_stage_opamp_dummy_magic_0.VOUT+.n0 GNDA 0.175369f
C996 two_stage_opamp_dummy_magic_0.VOUT+.t4 GNDA 0.043632f
C997 two_stage_opamp_dummy_magic_0.VOUT+.t8 GNDA 0.043632f
C998 two_stage_opamp_dummy_magic_0.VOUT+.n1 GNDA 0.175046f
C999 two_stage_opamp_dummy_magic_0.VOUT+.n2 GNDA 0.17244f
C1000 two_stage_opamp_dummy_magic_0.VOUT+.t3 GNDA 0.043632f
C1001 two_stage_opamp_dummy_magic_0.VOUT+.t7 GNDA 0.043632f
C1002 two_stage_opamp_dummy_magic_0.VOUT+.n3 GNDA 0.175046f
C1003 two_stage_opamp_dummy_magic_0.VOUT+.n4 GNDA 0.088927f
C1004 two_stage_opamp_dummy_magic_0.VOUT+.t11 GNDA 0.043632f
C1005 two_stage_opamp_dummy_magic_0.VOUT+.t5 GNDA 0.043632f
C1006 two_stage_opamp_dummy_magic_0.VOUT+.n5 GNDA 0.175046f
C1007 two_stage_opamp_dummy_magic_0.VOUT+.n6 GNDA 0.088927f
C1008 two_stage_opamp_dummy_magic_0.VOUT+.t10 GNDA 0.043632f
C1009 two_stage_opamp_dummy_magic_0.VOUT+.t15 GNDA 0.043632f
C1010 two_stage_opamp_dummy_magic_0.VOUT+.n7 GNDA 0.175368f
C1011 two_stage_opamp_dummy_magic_0.VOUT+.n8 GNDA 0.10533f
C1012 two_stage_opamp_dummy_magic_0.VOUT+.t12 GNDA 0.043632f
C1013 two_stage_opamp_dummy_magic_0.VOUT+.t6 GNDA 0.043632f
C1014 two_stage_opamp_dummy_magic_0.VOUT+.n9 GNDA 0.172903f
C1015 two_stage_opamp_dummy_magic_0.VOUT+.n10 GNDA 0.212302f
C1016 two_stage_opamp_dummy_magic_0.VOUT+.t117 GNDA 0.295834f
C1017 two_stage_opamp_dummy_magic_0.VOUT+.t25 GNDA 0.290879f
C1018 two_stage_opamp_dummy_magic_0.VOUT+.n11 GNDA 0.195025f
C1019 two_stage_opamp_dummy_magic_0.VOUT+.t124 GNDA 0.290879f
C1020 two_stage_opamp_dummy_magic_0.VOUT+.n12 GNDA 0.12726f
C1021 two_stage_opamp_dummy_magic_0.VOUT+.t72 GNDA 0.295834f
C1022 two_stage_opamp_dummy_magic_0.VOUT+.t38 GNDA 0.290879f
C1023 two_stage_opamp_dummy_magic_0.VOUT+.n13 GNDA 0.195025f
C1024 two_stage_opamp_dummy_magic_0.VOUT+.t127 GNDA 0.290879f
C1025 two_stage_opamp_dummy_magic_0.VOUT+.t34 GNDA 0.295213f
C1026 two_stage_opamp_dummy_magic_0.VOUT+.t86 GNDA 0.295213f
C1027 two_stage_opamp_dummy_magic_0.VOUT+.t42 GNDA 0.295213f
C1028 two_stage_opamp_dummy_magic_0.VOUT+.t96 GNDA 0.295213f
C1029 two_stage_opamp_dummy_magic_0.VOUT+.t143 GNDA 0.295213f
C1030 two_stage_opamp_dummy_magic_0.VOUT+.t106 GNDA 0.295213f
C1031 two_stage_opamp_dummy_magic_0.VOUT+.t154 GNDA 0.295213f
C1032 two_stage_opamp_dummy_magic_0.VOUT+.t64 GNDA 0.295213f
C1033 two_stage_opamp_dummy_magic_0.VOUT+.t116 GNDA 0.295213f
C1034 two_stage_opamp_dummy_magic_0.VOUT+.t73 GNDA 0.295213f
C1035 two_stage_opamp_dummy_magic_0.VOUT+.t149 GNDA 0.290879f
C1036 two_stage_opamp_dummy_magic_0.VOUT+.n14 GNDA 0.195645f
C1037 two_stage_opamp_dummy_magic_0.VOUT+.t58 GNDA 0.290879f
C1038 two_stage_opamp_dummy_magic_0.VOUT+.n15 GNDA 0.250185f
C1039 two_stage_opamp_dummy_magic_0.VOUT+.t97 GNDA 0.290879f
C1040 two_stage_opamp_dummy_magic_0.VOUT+.n16 GNDA 0.250185f
C1041 two_stage_opamp_dummy_magic_0.VOUT+.t131 GNDA 0.290879f
C1042 two_stage_opamp_dummy_magic_0.VOUT+.n17 GNDA 0.250185f
C1043 two_stage_opamp_dummy_magic_0.VOUT+.t24 GNDA 0.290879f
C1044 two_stage_opamp_dummy_magic_0.VOUT+.n18 GNDA 0.250185f
C1045 two_stage_opamp_dummy_magic_0.VOUT+.t75 GNDA 0.290879f
C1046 two_stage_opamp_dummy_magic_0.VOUT+.n19 GNDA 0.250185f
C1047 two_stage_opamp_dummy_magic_0.VOUT+.t113 GNDA 0.290879f
C1048 two_stage_opamp_dummy_magic_0.VOUT+.n20 GNDA 0.250185f
C1049 two_stage_opamp_dummy_magic_0.VOUT+.t144 GNDA 0.290879f
C1050 two_stage_opamp_dummy_magic_0.VOUT+.n21 GNDA 0.250185f
C1051 two_stage_opamp_dummy_magic_0.VOUT+.t54 GNDA 0.290879f
C1052 two_stage_opamp_dummy_magic_0.VOUT+.n22 GNDA 0.250185f
C1053 two_stage_opamp_dummy_magic_0.VOUT+.t94 GNDA 0.290879f
C1054 two_stage_opamp_dummy_magic_0.VOUT+.n23 GNDA 0.250185f
C1055 two_stage_opamp_dummy_magic_0.VOUT+.n24 GNDA 0.236339f
C1056 two_stage_opamp_dummy_magic_0.VOUT+.t37 GNDA 0.295834f
C1057 two_stage_opamp_dummy_magic_0.VOUT+.t142 GNDA 0.290879f
C1058 two_stage_opamp_dummy_magic_0.VOUT+.n25 GNDA 0.195025f
C1059 two_stage_opamp_dummy_magic_0.VOUT+.t93 GNDA 0.290879f
C1060 two_stage_opamp_dummy_magic_0.VOUT+.t20 GNDA 0.295834f
C1061 two_stage_opamp_dummy_magic_0.VOUT+.t57 GNDA 0.290879f
C1062 two_stage_opamp_dummy_magic_0.VOUT+.n26 GNDA 0.195025f
C1063 two_stage_opamp_dummy_magic_0.VOUT+.n27 GNDA 0.236339f
C1064 two_stage_opamp_dummy_magic_0.VOUT+.t79 GNDA 0.295834f
C1065 two_stage_opamp_dummy_magic_0.VOUT+.t41 GNDA 0.290879f
C1066 two_stage_opamp_dummy_magic_0.VOUT+.n28 GNDA 0.195025f
C1067 two_stage_opamp_dummy_magic_0.VOUT+.t133 GNDA 0.290879f
C1068 two_stage_opamp_dummy_magic_0.VOUT+.t60 GNDA 0.295834f
C1069 two_stage_opamp_dummy_magic_0.VOUT+.t100 GNDA 0.290879f
C1070 two_stage_opamp_dummy_magic_0.VOUT+.n29 GNDA 0.195025f
C1071 two_stage_opamp_dummy_magic_0.VOUT+.n30 GNDA 0.236339f
C1072 two_stage_opamp_dummy_magic_0.VOUT+.t121 GNDA 0.295834f
C1073 two_stage_opamp_dummy_magic_0.VOUT+.t83 GNDA 0.290879f
C1074 two_stage_opamp_dummy_magic_0.VOUT+.n31 GNDA 0.195025f
C1075 two_stage_opamp_dummy_magic_0.VOUT+.t31 GNDA 0.290879f
C1076 two_stage_opamp_dummy_magic_0.VOUT+.t104 GNDA 0.295834f
C1077 two_stage_opamp_dummy_magic_0.VOUT+.t137 GNDA 0.290879f
C1078 two_stage_opamp_dummy_magic_0.VOUT+.n32 GNDA 0.195025f
C1079 two_stage_opamp_dummy_magic_0.VOUT+.n33 GNDA 0.236339f
C1080 two_stage_opamp_dummy_magic_0.VOUT+.t84 GNDA 0.295834f
C1081 two_stage_opamp_dummy_magic_0.VOUT+.t49 GNDA 0.290879f
C1082 two_stage_opamp_dummy_magic_0.VOUT+.n34 GNDA 0.195025f
C1083 two_stage_opamp_dummy_magic_0.VOUT+.t138 GNDA 0.290879f
C1084 two_stage_opamp_dummy_magic_0.VOUT+.t66 GNDA 0.295834f
C1085 two_stage_opamp_dummy_magic_0.VOUT+.t103 GNDA 0.290879f
C1086 two_stage_opamp_dummy_magic_0.VOUT+.n35 GNDA 0.195025f
C1087 two_stage_opamp_dummy_magic_0.VOUT+.n36 GNDA 0.236339f
C1088 two_stage_opamp_dummy_magic_0.VOUT+.t108 GNDA 0.295834f
C1089 two_stage_opamp_dummy_magic_0.VOUT+.t69 GNDA 0.290879f
C1090 two_stage_opamp_dummy_magic_0.VOUT+.n37 GNDA 0.195025f
C1091 two_stage_opamp_dummy_magic_0.VOUT+.t90 GNDA 0.290879f
C1092 two_stage_opamp_dummy_magic_0.VOUT+.n38 GNDA 0.12726f
C1093 two_stage_opamp_dummy_magic_0.VOUT+.t67 GNDA 0.295834f
C1094 two_stage_opamp_dummy_magic_0.VOUT+.t30 GNDA 0.290879f
C1095 two_stage_opamp_dummy_magic_0.VOUT+.n39 GNDA 0.195025f
C1096 two_stage_opamp_dummy_magic_0.VOUT+.t51 GNDA 0.290879f
C1097 two_stage_opamp_dummy_magic_0.VOUT+.t53 GNDA 0.295213f
C1098 two_stage_opamp_dummy_magic_0.VOUT+.t156 GNDA 0.295213f
C1099 two_stage_opamp_dummy_magic_0.VOUT+.t44 GNDA 0.295834f
C1100 two_stage_opamp_dummy_magic_0.VOUT+.t136 GNDA 0.290879f
C1101 two_stage_opamp_dummy_magic_0.VOUT+.n40 GNDA 0.195025f
C1102 two_stage_opamp_dummy_magic_0.VOUT+.t101 GNDA 0.290879f
C1103 two_stage_opamp_dummy_magic_0.VOUT+.n41 GNDA 0.122715f
C1104 two_stage_opamp_dummy_magic_0.VOUT+.t36 GNDA 0.295213f
C1105 two_stage_opamp_dummy_magic_0.VOUT+.t151 GNDA 0.295834f
C1106 two_stage_opamp_dummy_magic_0.VOUT+.t98 GNDA 0.290879f
C1107 two_stage_opamp_dummy_magic_0.VOUT+.n42 GNDA 0.195025f
C1108 two_stage_opamp_dummy_magic_0.VOUT+.t59 GNDA 0.290879f
C1109 two_stage_opamp_dummy_magic_0.VOUT+.n43 GNDA 0.122715f
C1110 two_stage_opamp_dummy_magic_0.VOUT+.t140 GNDA 0.295213f
C1111 two_stage_opamp_dummy_magic_0.VOUT+.t118 GNDA 0.295834f
C1112 two_stage_opamp_dummy_magic_0.VOUT+.t56 GNDA 0.290879f
C1113 two_stage_opamp_dummy_magic_0.VOUT+.n44 GNDA 0.195025f
C1114 two_stage_opamp_dummy_magic_0.VOUT+.t21 GNDA 0.290879f
C1115 two_stage_opamp_dummy_magic_0.VOUT+.n45 GNDA 0.122715f
C1116 two_stage_opamp_dummy_magic_0.VOUT+.t105 GNDA 0.295213f
C1117 two_stage_opamp_dummy_magic_0.VOUT+.t65 GNDA 0.295834f
C1118 two_stage_opamp_dummy_magic_0.VOUT+.t80 GNDA 0.290879f
C1119 two_stage_opamp_dummy_magic_0.VOUT+.n46 GNDA 0.195025f
C1120 two_stage_opamp_dummy_magic_0.VOUT+.t43 GNDA 0.290879f
C1121 two_stage_opamp_dummy_magic_0.VOUT+.n47 GNDA 0.122715f
C1122 two_stage_opamp_dummy_magic_0.VOUT+.t125 GNDA 0.295213f
C1123 two_stage_opamp_dummy_magic_0.VOUT+.t145 GNDA 0.295457f
C1124 two_stage_opamp_dummy_magic_0.VOUT+.t87 GNDA 0.295213f
C1125 two_stage_opamp_dummy_magic_0.VOUT+.t110 GNDA 0.295457f
C1126 two_stage_opamp_dummy_magic_0.VOUT+.t50 GNDA 0.295213f
C1127 two_stage_opamp_dummy_magic_0.VOUT+.t70 GNDA 0.295457f
C1128 two_stage_opamp_dummy_magic_0.VOUT+.t150 GNDA 0.295213f
C1129 two_stage_opamp_dummy_magic_0.VOUT+.t95 GNDA 0.295457f
C1130 two_stage_opamp_dummy_magic_0.VOUT+.t32 GNDA 0.295213f
C1131 two_stage_opamp_dummy_magic_0.VOUT+.t134 GNDA 0.290879f
C1132 two_stage_opamp_dummy_magic_0.VOUT+.n48 GNDA 0.321963f
C1133 two_stage_opamp_dummy_magic_0.VOUT+.t111 GNDA 0.290879f
C1134 two_stage_opamp_dummy_magic_0.VOUT+.n49 GNDA 0.376503f
C1135 two_stage_opamp_dummy_magic_0.VOUT+.t147 GNDA 0.290879f
C1136 two_stage_opamp_dummy_magic_0.VOUT+.n50 GNDA 0.376503f
C1137 two_stage_opamp_dummy_magic_0.VOUT+.t45 GNDA 0.290879f
C1138 two_stage_opamp_dummy_magic_0.VOUT+.n51 GNDA 0.376503f
C1139 two_stage_opamp_dummy_magic_0.VOUT+.t85 GNDA 0.290879f
C1140 two_stage_opamp_dummy_magic_0.VOUT+.n52 GNDA 0.30927f
C1141 two_stage_opamp_dummy_magic_0.VOUT+.t61 GNDA 0.290879f
C1142 two_stage_opamp_dummy_magic_0.VOUT+.n53 GNDA 0.30927f
C1143 two_stage_opamp_dummy_magic_0.VOUT+.t102 GNDA 0.290879f
C1144 two_stage_opamp_dummy_magic_0.VOUT+.n54 GNDA 0.30927f
C1145 two_stage_opamp_dummy_magic_0.VOUT+.t139 GNDA 0.290879f
C1146 two_stage_opamp_dummy_magic_0.VOUT+.n55 GNDA 0.30927f
C1147 two_stage_opamp_dummy_magic_0.VOUT+.t119 GNDA 0.290879f
C1148 two_stage_opamp_dummy_magic_0.VOUT+.n56 GNDA 0.250185f
C1149 two_stage_opamp_dummy_magic_0.VOUT+.t155 GNDA 0.290879f
C1150 two_stage_opamp_dummy_magic_0.VOUT+.n57 GNDA 0.250185f
C1151 two_stage_opamp_dummy_magic_0.VOUT+.n58 GNDA 0.236339f
C1152 two_stage_opamp_dummy_magic_0.VOUT+.t27 GNDA 0.295834f
C1153 two_stage_opamp_dummy_magic_0.VOUT+.t130 GNDA 0.290879f
C1154 two_stage_opamp_dummy_magic_0.VOUT+.n59 GNDA 0.195025f
C1155 two_stage_opamp_dummy_magic_0.VOUT+.t152 GNDA 0.290879f
C1156 two_stage_opamp_dummy_magic_0.VOUT+.t76 GNDA 0.295834f
C1157 two_stage_opamp_dummy_magic_0.VOUT+.t115 GNDA 0.290879f
C1158 two_stage_opamp_dummy_magic_0.VOUT+.n60 GNDA 0.195025f
C1159 two_stage_opamp_dummy_magic_0.VOUT+.n61 GNDA 0.236339f
C1160 two_stage_opamp_dummy_magic_0.VOUT+.t62 GNDA 0.295834f
C1161 two_stage_opamp_dummy_magic_0.VOUT+.t23 GNDA 0.290879f
C1162 two_stage_opamp_dummy_magic_0.VOUT+.n62 GNDA 0.195025f
C1163 two_stage_opamp_dummy_magic_0.VOUT+.t47 GNDA 0.290879f
C1164 two_stage_opamp_dummy_magic_0.VOUT+.t112 GNDA 0.295834f
C1165 two_stage_opamp_dummy_magic_0.VOUT+.t148 GNDA 0.290879f
C1166 two_stage_opamp_dummy_magic_0.VOUT+.n63 GNDA 0.195025f
C1167 two_stage_opamp_dummy_magic_0.VOUT+.n64 GNDA 0.236339f
C1168 two_stage_opamp_dummy_magic_0.VOUT+.t114 GNDA 0.295834f
C1169 two_stage_opamp_dummy_magic_0.VOUT+.t78 GNDA 0.290879f
C1170 two_stage_opamp_dummy_magic_0.VOUT+.n65 GNDA 0.195025f
C1171 two_stage_opamp_dummy_magic_0.VOUT+.t26 GNDA 0.290879f
C1172 two_stage_opamp_dummy_magic_0.VOUT+.t99 GNDA 0.295834f
C1173 two_stage_opamp_dummy_magic_0.VOUT+.t132 GNDA 0.290879f
C1174 two_stage_opamp_dummy_magic_0.VOUT+.n66 GNDA 0.195025f
C1175 two_stage_opamp_dummy_magic_0.VOUT+.n67 GNDA 0.236339f
C1176 two_stage_opamp_dummy_magic_0.VOUT+.t74 GNDA 0.295834f
C1177 two_stage_opamp_dummy_magic_0.VOUT+.t39 GNDA 0.290879f
C1178 two_stage_opamp_dummy_magic_0.VOUT+.n68 GNDA 0.195025f
C1179 two_stage_opamp_dummy_magic_0.VOUT+.t128 GNDA 0.290879f
C1180 two_stage_opamp_dummy_magic_0.VOUT+.t55 GNDA 0.295834f
C1181 two_stage_opamp_dummy_magic_0.VOUT+.t92 GNDA 0.290879f
C1182 two_stage_opamp_dummy_magic_0.VOUT+.n69 GNDA 0.195025f
C1183 two_stage_opamp_dummy_magic_0.VOUT+.n70 GNDA 0.236339f
C1184 two_stage_opamp_dummy_magic_0.VOUT+.t109 GNDA 0.295834f
C1185 two_stage_opamp_dummy_magic_0.VOUT+.t71 GNDA 0.290879f
C1186 two_stage_opamp_dummy_magic_0.VOUT+.n71 GNDA 0.195025f
C1187 two_stage_opamp_dummy_magic_0.VOUT+.t19 GNDA 0.290879f
C1188 two_stage_opamp_dummy_magic_0.VOUT+.t91 GNDA 0.295834f
C1189 two_stage_opamp_dummy_magic_0.VOUT+.t126 GNDA 0.290879f
C1190 two_stage_opamp_dummy_magic_0.VOUT+.n72 GNDA 0.195025f
C1191 two_stage_opamp_dummy_magic_0.VOUT+.n73 GNDA 0.236339f
C1192 two_stage_opamp_dummy_magic_0.VOUT+.t68 GNDA 0.295834f
C1193 two_stage_opamp_dummy_magic_0.VOUT+.t33 GNDA 0.290879f
C1194 two_stage_opamp_dummy_magic_0.VOUT+.n74 GNDA 0.195025f
C1195 two_stage_opamp_dummy_magic_0.VOUT+.t122 GNDA 0.290879f
C1196 two_stage_opamp_dummy_magic_0.VOUT+.t52 GNDA 0.295834f
C1197 two_stage_opamp_dummy_magic_0.VOUT+.t88 GNDA 0.290879f
C1198 two_stage_opamp_dummy_magic_0.VOUT+.n75 GNDA 0.195025f
C1199 two_stage_opamp_dummy_magic_0.VOUT+.n76 GNDA 0.236339f
C1200 two_stage_opamp_dummy_magic_0.VOUT+.t29 GNDA 0.295834f
C1201 two_stage_opamp_dummy_magic_0.VOUT+.t135 GNDA 0.290879f
C1202 two_stage_opamp_dummy_magic_0.VOUT+.n77 GNDA 0.195025f
C1203 two_stage_opamp_dummy_magic_0.VOUT+.t82 GNDA 0.290879f
C1204 two_stage_opamp_dummy_magic_0.VOUT+.t153 GNDA 0.295834f
C1205 two_stage_opamp_dummy_magic_0.VOUT+.t48 GNDA 0.290879f
C1206 two_stage_opamp_dummy_magic_0.VOUT+.n78 GNDA 0.195025f
C1207 two_stage_opamp_dummy_magic_0.VOUT+.n79 GNDA 0.236339f
C1208 two_stage_opamp_dummy_magic_0.VOUT+.t63 GNDA 0.295834f
C1209 two_stage_opamp_dummy_magic_0.VOUT+.t28 GNDA 0.290879f
C1210 two_stage_opamp_dummy_magic_0.VOUT+.n80 GNDA 0.195025f
C1211 two_stage_opamp_dummy_magic_0.VOUT+.t120 GNDA 0.290879f
C1212 two_stage_opamp_dummy_magic_0.VOUT+.t46 GNDA 0.295834f
C1213 two_stage_opamp_dummy_magic_0.VOUT+.t81 GNDA 0.290879f
C1214 two_stage_opamp_dummy_magic_0.VOUT+.n81 GNDA 0.195025f
C1215 two_stage_opamp_dummy_magic_0.VOUT+.n82 GNDA 0.236339f
C1216 two_stage_opamp_dummy_magic_0.VOUT+.t22 GNDA 0.295834f
C1217 two_stage_opamp_dummy_magic_0.VOUT+.t129 GNDA 0.290879f
C1218 two_stage_opamp_dummy_magic_0.VOUT+.n83 GNDA 0.195025f
C1219 two_stage_opamp_dummy_magic_0.VOUT+.t77 GNDA 0.290879f
C1220 two_stage_opamp_dummy_magic_0.VOUT+.t146 GNDA 0.295834f
C1221 two_stage_opamp_dummy_magic_0.VOUT+.t40 GNDA 0.290879f
C1222 two_stage_opamp_dummy_magic_0.VOUT+.n84 GNDA 0.195025f
C1223 two_stage_opamp_dummy_magic_0.VOUT+.n85 GNDA 0.236339f
C1224 two_stage_opamp_dummy_magic_0.VOUT+.t123 GNDA 0.295834f
C1225 two_stage_opamp_dummy_magic_0.VOUT+.t89 GNDA 0.290879f
C1226 two_stage_opamp_dummy_magic_0.VOUT+.n86 GNDA 0.195025f
C1227 two_stage_opamp_dummy_magic_0.VOUT+.t35 GNDA 0.290879f
C1228 two_stage_opamp_dummy_magic_0.VOUT+.n87 GNDA 0.236339f
C1229 two_stage_opamp_dummy_magic_0.VOUT+.t141 GNDA 0.290879f
C1230 two_stage_opamp_dummy_magic_0.VOUT+.n88 GNDA 0.12726f
C1231 two_stage_opamp_dummy_magic_0.VOUT+.t107 GNDA 0.290879f
C1232 two_stage_opamp_dummy_magic_0.VOUT+.n89 GNDA 0.238316f
C1233 two_stage_opamp_dummy_magic_0.VOUT+.n90 GNDA 0.291354f
C1234 two_stage_opamp_dummy_magic_0.VOUT+.t1 GNDA 0.050904f
C1235 two_stage_opamp_dummy_magic_0.VOUT+.t16 GNDA 0.050904f
C1236 two_stage_opamp_dummy_magic_0.VOUT+.n91 GNDA 0.235484f
C1237 two_stage_opamp_dummy_magic_0.VOUT+.t0 GNDA 0.050904f
C1238 two_stage_opamp_dummy_magic_0.VOUT+.t13 GNDA 0.050904f
C1239 two_stage_opamp_dummy_magic_0.VOUT+.n92 GNDA 0.234695f
C1240 two_stage_opamp_dummy_magic_0.VOUT+.n93 GNDA 0.14503f
C1241 two_stage_opamp_dummy_magic_0.VOUT+.t17 GNDA 0.050904f
C1242 two_stage_opamp_dummy_magic_0.VOUT+.t18 GNDA 0.050904f
C1243 two_stage_opamp_dummy_magic_0.VOUT+.n94 GNDA 0.234695f
C1244 two_stage_opamp_dummy_magic_0.VOUT+.n95 GNDA 0.089271f
C1245 two_stage_opamp_dummy_magic_0.VOUT+.n96 GNDA 0.165389f
C1246 two_stage_opamp_dummy_magic_0.VOUT+.t2 GNDA 0.084162f
C1247 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.019819f
C1248 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.019819f
C1249 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.066913f
C1250 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.019819f
C1251 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.019819f
C1252 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.071516f
C1253 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.019819f
C1254 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.019819f
C1255 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.070891f
C1256 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.26322f
C1257 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.019819f
C1258 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.019819f
C1259 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.070891f
C1260 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.136547f
C1261 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.019819f
C1262 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.019819f
C1263 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.070891f
C1264 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.136547f
C1265 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.019819f
C1266 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.019819f
C1267 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.070891f
C1268 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.163559f
C1269 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.137812f
C1270 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.645498f
C1271 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.087203f
C1272 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.087203f
C1273 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.092877f
C1274 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.073601f
C1275 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.039346f
C1276 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.087203f
C1277 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.087203f
C1278 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.087203f
C1279 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.087203f
C1280 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.087203f
C1281 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.087203f
C1282 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.092877f
C1283 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.073601f
C1284 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.04162f
C1285 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.04162f
C1286 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.04162f
C1287 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.04162f
C1288 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.039346f
C1289 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.02132f
C1290 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.765352f
C1291 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.027747f
C1292 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.027747f
C1293 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.027747f
C1294 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.027747f
C1295 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.027747f
C1296 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.027747f
C1297 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.027747f
C1298 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.033692f
C1299 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.033692f
C1300 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.021801f
C1301 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.021801f
C1302 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.021801f
C1303 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.021801f
C1304 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.021801f
C1305 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.019527f
C1306 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.027747f
C1307 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.033692f
C1308 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.031419f
C1309 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.019205f
C1310 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.042611f
C1311 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.042611f
C1312 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.042611f
C1313 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.042611f
C1314 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.042611f
C1315 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.042611f
C1316 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.042611f
C1317 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.048441f
C1318 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.043717f
C1319 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.026756f
C1320 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.026756f
C1321 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.026756f
C1322 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.026756f
C1323 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.026756f
C1324 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.024482f
C1325 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.042611f
C1326 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.048441f
C1327 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.041443f
C1328 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.019165f
C1329 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.251975f
C1330 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.347762f
C1331 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.08699f
C1332 a_8420_8490.t7 GNDA 0.066432f
C1333 a_8420_8490.t11 GNDA 0.066432f
C1334 a_8420_8490.t4 GNDA 0.066432f
C1335 a_8420_8490.n0 GNDA 0.231036f
C1336 a_8420_8490.t6 GNDA 0.066432f
C1337 a_8420_8490.t8 GNDA 0.066432f
C1338 a_8420_8490.n1 GNDA 0.230217f
C1339 a_8420_8490.n2 GNDA 0.434626f
C1340 a_8420_8490.t0 GNDA 0.066432f
C1341 a_8420_8490.t2 GNDA 0.066432f
C1342 a_8420_8490.n3 GNDA 0.230217f
C1343 a_8420_8490.n4 GNDA 0.225315f
C1344 a_8420_8490.t3 GNDA 0.066432f
C1345 a_8420_8490.t5 GNDA 0.066432f
C1346 a_8420_8490.n5 GNDA 0.230217f
C1347 a_8420_8490.n6 GNDA 0.225315f
C1348 a_8420_8490.t1 GNDA 0.066432f
C1349 a_8420_8490.t10 GNDA 0.066432f
C1350 a_8420_8490.n7 GNDA 0.231035f
C1351 a_8420_8490.n8 GNDA 0.434627f
C1352 a_8420_8490.n9 GNDA 0.230216f
C1353 a_8420_8490.t9 GNDA 0.066432f
C1354 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.026064f
C1355 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.026064f
C1356 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.090645f
C1357 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.026064f
C1358 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.026064f
C1359 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.090324f
C1360 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.170523f
C1361 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.074201f
C1362 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.100899f
C1363 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.128579f
C1364 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.045386f
C1365 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.083882f
C1366 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.054074f
C1367 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.128579f
C1368 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.045386f
C1369 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.083882f
C1370 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.054074f
C1371 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.053617f
C1372 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.100899f
C1373 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.300697f
C1374 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.448835f
C1375 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.259151f
C1376 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.259151f
C1377 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.259151f
C1378 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.259151f
C1379 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.194363f
C1380 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.129575f
C1381 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.194363f
C1382 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.259151f
C1383 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.259151f
C1384 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.259151f
C1385 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.259151f
C1386 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.448835f
C1387 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.300697f
C1388 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.074201f
C1389 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.103878f
C1390 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.026064f
C1391 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.026064f
C1392 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.08498f
C1393 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.061885f
C1394 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.03186f
C1395 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.026064f
C1396 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.026064f
C1397 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.090324f
C1398 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.085422f
C1399 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.026064f
C1400 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.026064f
C1401 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.090324f
C1402 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.11501f
C1403 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.026064f
C1404 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.026064f
C1405 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.090645f
C1406 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.026064f
C1407 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.026064f
C1408 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.090324f
C1409 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.170523f
C1410 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.026064f
C1411 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.026064f
C1412 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.090324f
C1413 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.088401f
C1414 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.026064f
C1415 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.026064f
C1416 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.090324f
C1417 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.088401f
C1418 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.026064f
C1419 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.026064f
C1420 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.090324f
C1421 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.088401f
C1422 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.026064f
C1423 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.026064f
C1424 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.090324f
C1425 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.133988f
C1426 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.012583f
C1427 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.012583f
C1428 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.027269f
C1429 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.03908f
C1430 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.168132f
C1431 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.09887f
C1432 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.09887f
C1433 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.09887f
C1434 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.09887f
C1435 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.114095f
C1436 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.092633f
C1437 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.056925f
C1438 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.056925f
C1439 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.053303f
C1440 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.09887f
C1441 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.09887f
C1442 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.09887f
C1443 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.09887f
C1444 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.114095f
C1445 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.092633f
C1446 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.056925f
C1447 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.056925f
C1448 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.053303f
C1449 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.036003f
C1450 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.09887f
C1451 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.09887f
C1452 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.09887f
C1453 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.09887f
C1454 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.114095f
C1455 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.092633f
C1456 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.056925f
C1457 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.056925f
C1458 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.053303f
C1459 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.09887f
C1460 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.09887f
C1461 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.09887f
C1462 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.09887f
C1463 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.114095f
C1464 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.092633f
C1465 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.056925f
C1466 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.056925f
C1467 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.053303f
C1468 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.035316f
C1469 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.802639f
C1470 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.604613f
C1471 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.119293f
C1472 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 3.15867f
C1473 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.019974f
C1474 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.019974f
C1475 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.066969f
C1476 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.019974f
C1477 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.019974f
C1478 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.065132f
C1479 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.526032f
C1480 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.019974f
C1481 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.019974f
C1482 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.066969f
C1483 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.019974f
C1484 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.019974f
C1485 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.065132f
C1486 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.526032f
C1487 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.274372f
C1488 bgr_0.VB2_CUR_BIAS GNDA 3.05596f
C1489 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.7726f
C1490 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 8.91394f
C1491 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.024917f
C1492 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.024917f
C1493 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.058161f
C1494 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.024917f
C1495 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.024917f
C1496 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.057785f
C1497 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.024917f
C1498 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.024917f
C1499 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.057785f
C1500 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.020556f
C1501 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.020556f
C1502 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.020556f
C1503 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.020556f
C1504 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.020556f
C1505 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.020556f
C1506 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.020556f
C1507 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.020556f
C1508 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.020556f
C1509 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.020556f
C1510 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.020556f
C1511 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.020556f
C1512 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.020556f
C1513 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.020556f
C1514 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.020556f
C1515 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.020556f
C1516 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.044539f
C1517 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.069456f
C1518 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.054194f
C1519 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.054194f
C1520 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.054194f
C1521 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.054194f
C1522 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.054194f
C1523 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.054194f
C1524 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.054194f
C1525 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.054194f
C1526 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.054194f
C1527 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.054194f
C1528 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.054194f
C1529 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.054194f
C1530 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.054194f
C1531 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.054194f
C1532 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.046376f
C1533 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.020556f
C1534 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.020556f
C1535 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.044539f
C1536 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.069456f
C1537 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.046376f
C1538 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.075239f
C1539 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.024917f
C1540 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.024917f
C1541 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.049834f
C1542 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.148444f
C1543 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.024917f
C1544 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.024917f
C1545 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.057785f
C1546 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.024917f
C1547 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.024917f
C1548 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.057355f
C1549 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.049834f
C1550 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.049834f
C1551 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.153708f
C1552 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.074255f
C1553 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.027767f
C1554 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.087091f
C1555 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.027767f
C1556 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.071293f
C1557 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.027767f
C1558 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.071293f
C1559 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.027767f
C1560 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.109376f
C1561 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.709082f
C1562 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.090054f
C1563 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.090054f
C1564 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.301772f
C1565 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 3.40029f
C1566 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.090054f
C1567 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.090054f
C1568 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.301772f
C1569 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.814897f
C1570 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.090054f
C1571 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.090054f
C1572 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.301772f
C1573 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 1.16504f
C1574 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 1.01344f
C1575 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.043395f
C1576 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.013631f
C1577 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.025436f
C1578 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.060728f
C1579 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.379723f
C1580 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.013631f
C1581 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.025436f
C1582 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.060728f
C1583 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.350774f
C1584 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.042979f
C1585 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.341551f
C1586 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.013631f
C1587 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.025436f
C1588 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.060728f
C1589 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.212091f
C1590 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.013631f
C1591 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.025436f
C1592 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.060728f
C1593 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.269546f
C1594 bgr_0.V_mir2.t2 GNDA 0.042444f
C1595 bgr_0.V_mir2.t18 GNDA 0.042444f
C1596 bgr_0.V_mir2.t20 GNDA 0.06851f
C1597 bgr_0.V_mir2.n0 GNDA 0.076506f
C1598 bgr_0.V_mir2.n1 GNDA 0.052264f
C1599 bgr_0.V_mir2.t6 GNDA 0.053881f
C1600 bgr_0.V_mir2.n2 GNDA 0.081315f
C1601 bgr_0.V_mir2.t3 GNDA 0.03537f
C1602 bgr_0.V_mir2.t7 GNDA 0.03537f
C1603 bgr_0.V_mir2.n3 GNDA 0.08097f
C1604 bgr_0.V_mir2.n4 GNDA 0.201563f
C1605 bgr_0.V_mir2.t16 GNDA 0.017685f
C1606 bgr_0.V_mir2.t1 GNDA 0.017685f
C1607 bgr_0.V_mir2.n5 GNDA 0.046242f
C1608 bgr_0.V_mir2.t15 GNDA 0.075466f
C1609 bgr_0.V_mir2.t14 GNDA 0.017685f
C1610 bgr_0.V_mir2.t0 GNDA 0.017685f
C1611 bgr_0.V_mir2.n6 GNDA 0.050199f
C1612 bgr_0.V_mir2.n7 GNDA 0.827814f
C1613 bgr_0.V_mir2.n8 GNDA 0.268286f
C1614 bgr_0.V_mir2.t10 GNDA 0.042444f
C1615 bgr_0.V_mir2.t19 GNDA 0.042444f
C1616 bgr_0.V_mir2.t22 GNDA 0.06851f
C1617 bgr_0.V_mir2.n9 GNDA 0.076506f
C1618 bgr_0.V_mir2.n10 GNDA 0.052264f
C1619 bgr_0.V_mir2.t8 GNDA 0.053881f
C1620 bgr_0.V_mir2.n11 GNDA 0.081315f
C1621 bgr_0.V_mir2.t11 GNDA 0.03537f
C1622 bgr_0.V_mir2.t9 GNDA 0.03537f
C1623 bgr_0.V_mir2.n12 GNDA 0.08097f
C1624 bgr_0.V_mir2.n13 GNDA 0.156007f
C1625 bgr_0.V_mir2.n14 GNDA 0.09373f
C1626 bgr_0.V_mir2.n15 GNDA 0.699157f
C1627 bgr_0.V_mir2.t12 GNDA 0.042444f
C1628 bgr_0.V_mir2.t21 GNDA 0.042444f
C1629 bgr_0.V_mir2.t17 GNDA 0.06851f
C1630 bgr_0.V_mir2.n16 GNDA 0.076506f
C1631 bgr_0.V_mir2.n17 GNDA 0.052264f
C1632 bgr_0.V_mir2.t4 GNDA 0.053881f
C1633 bgr_0.V_mir2.n18 GNDA 0.081315f
C1634 bgr_0.V_mir2.n19 GNDA 0.203577f
C1635 bgr_0.V_mir2.t5 GNDA 0.03537f
C1636 bgr_0.V_mir2.n20 GNDA 0.08097f
C1637 bgr_0.V_mir2.t13 GNDA 0.03537f
C1638 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.03109f
C1639 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.03109f
C1640 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.077932f
C1641 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.03109f
C1642 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.03109f
C1643 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.077521f
C1644 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.689005f
C1645 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.03109f
C1646 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.03109f
C1647 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.06218f
C1648 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.347514f
C1649 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.398172f
C1650 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.06218f
C1651 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.06218f
C1652 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.182434f
C1653 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.06218f
C1654 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.06218f
C1655 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.181606f
C1656 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.627735f
C1657 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.06218f
C1658 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.06218f
C1659 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.181606f
C1660 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.325163f
C1661 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.06218f
C1662 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.06218f
C1663 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.181606f
C1664 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.325163f
C1665 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.06218f
C1666 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.06218f
C1667 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.181606f
C1668 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.467149f
C1669 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 3.26646f
C1670 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 3.56079f
C1671 bgr_0.V_CMFB_S1 GNDA 0.058021f
C1672 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.020126f
C1673 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.020126f
C1674 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.067951f
C1675 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.020126f
C1676 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.020126f
C1677 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.072625f
C1678 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.020126f
C1679 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.020126f
C1680 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.071991f
C1681 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.267304f
C1682 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.020126f
C1683 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.020126f
C1684 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.071991f
C1685 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.138665f
C1686 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.020126f
C1687 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.020126f
C1688 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.071991f
C1689 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.138665f
C1690 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.020126f
C1691 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.020126f
C1692 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.071991f
C1693 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.166097f
C1694 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.214408f
C1695 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.028177f
C1696 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.034215f
C1697 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.031906f
C1698 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.028177f
C1699 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.028177f
C1700 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.028177f
C1701 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.028177f
C1702 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.028177f
C1703 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.028177f
C1704 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.028177f
C1705 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.034215f
C1706 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.034215f
C1707 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.022139f
C1708 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.022139f
C1709 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.022139f
C1710 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.022139f
C1711 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.022139f
C1712 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.01983f
C1713 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.019503f
C1714 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.043272f
C1715 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.049193f
C1716 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.042086f
C1717 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.043272f
C1718 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.043272f
C1719 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.043272f
C1720 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.043272f
C1721 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.043272f
C1722 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.043272f
C1723 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.043272f
C1724 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.049193f
C1725 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.044395f
C1726 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.027171f
C1727 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.027171f
C1728 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.027171f
C1729 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.027171f
C1730 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.027171f
C1731 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.024862f
C1732 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.019462f
C1733 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.259144f
C1734 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.37183f
C1735 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.088556f
C1736 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.088556f
C1737 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.088556f
C1738 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.088556f
C1739 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.088556f
C1740 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.088556f
C1741 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.094318f
C1742 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.074743f
C1743 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.042265f
C1744 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.042265f
C1745 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.042265f
C1746 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.042265f
C1747 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.039957f
C1748 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.088556f
C1749 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.088556f
C1750 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.094318f
C1751 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.074743f
C1752 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.039957f
C1753 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.021651f
C1754 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.77991f
C1755 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.655511f
C1756 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.343499f
C1757 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.344645f
C1758 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.185116f
C1759 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.197667f
C1760 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.343499f
C1761 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.344645f
C1762 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.185116f
C1763 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.216163f
C1764 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.343499f
C1765 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.344645f
C1766 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.185116f
C1767 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.216163f
C1768 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.343499f
C1769 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.344645f
C1770 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.185116f
C1771 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.216163f
C1772 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.343499f
C1773 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C1774 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.363141f
C1775 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.363141f
C1776 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.185116f
C1777 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.216163f
C1778 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.343499f
C1779 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.344645f
C1780 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.363141f
C1781 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.363141f
C1782 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.185116f
C1783 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.216163f
C1784 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.344645f
C1785 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.345894f
C1786 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344645f
C1787 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.347347f
C1788 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.377789f
C1789 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.344645f
C1790 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.345894f
C1791 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.344645f
C1792 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.345894f
C1793 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.344645f
C1794 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345894f
C1795 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.344645f
C1796 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.345894f
C1797 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.344645f
C1798 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.345894f
C1799 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.344645f
C1800 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.345894f
C1801 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.344645f
C1802 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.345894f
C1803 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.344645f
C1804 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.345894f
C1805 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.344645f
C1806 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345894f
C1807 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.344645f
C1808 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.345894f
C1809 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.344645f
C1810 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.345894f
C1811 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.344645f
C1812 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.345894f
C1813 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.344645f
C1814 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.345894f
C1815 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.344645f
C1816 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.345894f
C1817 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.344645f
C1818 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.345894f
C1819 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.344645f
C1820 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.345894f
C1821 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.344645f
C1822 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.345894f
C1823 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.344645f
C1824 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.345894f
C1825 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.344645f
C1826 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.345894f
C1827 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.344645f
C1828 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.345894f
C1829 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.344645f
C1830 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.345894f
C1831 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.344645f
C1832 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.345894f
C1833 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.344645f
C1834 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.345894f
C1835 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.344645f
C1836 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.345894f
C1837 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.344645f
C1838 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.345894f
C1839 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.344645f
C1840 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345894f
C1841 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.344645f
C1842 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.345894f
C1843 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.344645f
C1844 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.345894f
C1845 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.344645f
C1846 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.361543f
C1847 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.344645f
C1848 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.185116f
C1849 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.19812f
C1850 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.344645f
C1851 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.185116f
C1852 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.196521f
C1853 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.344645f
C1854 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.185116f
C1855 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.196521f
C1856 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.344645f
C1857 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.185116f
C1858 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.196521f
C1859 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.344645f
C1860 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185116f
C1861 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.196521f
C1862 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.344645f
C1863 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.185116f
C1864 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.196521f
C1865 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.344645f
C1866 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.185116f
C1867 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.196521f
C1868 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.344645f
C1869 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.185116f
C1870 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.196521f
C1871 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.344645f
C1872 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185116f
C1873 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.196521f
C1874 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.344645f
C1875 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.345894f
C1876 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.344645f
C1877 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.345894f
C1878 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.166619f
C1879 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.214914f
C1880 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.18397f
C1881 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.23341f
C1882 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.18397f
C1883 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.250658f
C1884 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.18397f
C1885 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.250658f
C1886 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.18397f
C1887 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.250658f
C1888 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.18397f
C1889 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.250658f
C1890 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.18397f
C1891 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.250658f
C1892 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.18397f
C1893 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.250658f
C1894 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.18397f
C1895 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.250658f
C1896 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.18397f
C1897 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.250658f
C1898 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.18397f
C1899 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.250658f
C1900 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.18397f
C1901 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.250658f
C1902 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.18397f
C1903 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.250658f
C1904 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.18397f
C1905 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.250658f
C1906 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.18397f
C1907 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.250658f
C1908 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.18397f
C1909 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.250658f
C1910 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.18397f
C1911 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.23341f
C1912 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.343499f
C1913 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.166619f
C1914 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216163f
C1915 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.343499f
C1916 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.166619f
C1917 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216163f
C1918 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.343499f
C1919 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.344645f
C1920 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.363141f
C1921 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.363141f
C1922 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.185116f
C1923 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216163f
C1924 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.343499f
C1925 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216163f
C1926 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185116f
C1927 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.363141f
C1928 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.363141f
C1929 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.434494f
C1930 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.297192f
C1931 two_stage_opamp_dummy_magic_0.VOUT-.t16 GNDA 0.050904f
C1932 two_stage_opamp_dummy_magic_0.VOUT-.t11 GNDA 0.050904f
C1933 two_stage_opamp_dummy_magic_0.VOUT-.n0 GNDA 0.235484f
C1934 two_stage_opamp_dummy_magic_0.VOUT-.t12 GNDA 0.050904f
C1935 two_stage_opamp_dummy_magic_0.VOUT-.t4 GNDA 0.050904f
C1936 two_stage_opamp_dummy_magic_0.VOUT-.n1 GNDA 0.234695f
C1937 two_stage_opamp_dummy_magic_0.VOUT-.n2 GNDA 0.14503f
C1938 two_stage_opamp_dummy_magic_0.VOUT-.t3 GNDA 0.050904f
C1939 two_stage_opamp_dummy_magic_0.VOUT-.t17 GNDA 0.050904f
C1940 two_stage_opamp_dummy_magic_0.VOUT-.n3 GNDA 0.234695f
C1941 two_stage_opamp_dummy_magic_0.VOUT-.n4 GNDA 0.089271f
C1942 two_stage_opamp_dummy_magic_0.VOUT-.t14 GNDA 0.043632f
C1943 two_stage_opamp_dummy_magic_0.VOUT-.t6 GNDA 0.043632f
C1944 two_stage_opamp_dummy_magic_0.VOUT-.n5 GNDA 0.175369f
C1945 two_stage_opamp_dummy_magic_0.VOUT-.t8 GNDA 0.043632f
C1946 two_stage_opamp_dummy_magic_0.VOUT-.t15 GNDA 0.043632f
C1947 two_stage_opamp_dummy_magic_0.VOUT-.n6 GNDA 0.175368f
C1948 two_stage_opamp_dummy_magic_0.VOUT-.t9 GNDA 0.043632f
C1949 two_stage_opamp_dummy_magic_0.VOUT-.t10 GNDA 0.043632f
C1950 two_stage_opamp_dummy_magic_0.VOUT-.n7 GNDA 0.175046f
C1951 two_stage_opamp_dummy_magic_0.VOUT-.n8 GNDA 0.172441f
C1952 two_stage_opamp_dummy_magic_0.VOUT-.t1 GNDA 0.043632f
C1953 two_stage_opamp_dummy_magic_0.VOUT-.t13 GNDA 0.043632f
C1954 two_stage_opamp_dummy_magic_0.VOUT-.n9 GNDA 0.175046f
C1955 two_stage_opamp_dummy_magic_0.VOUT-.n10 GNDA 0.088927f
C1956 two_stage_opamp_dummy_magic_0.VOUT-.t2 GNDA 0.043632f
C1957 two_stage_opamp_dummy_magic_0.VOUT-.t7 GNDA 0.043632f
C1958 two_stage_opamp_dummy_magic_0.VOUT-.n11 GNDA 0.175046f
C1959 two_stage_opamp_dummy_magic_0.VOUT-.n12 GNDA 0.088927f
C1960 two_stage_opamp_dummy_magic_0.VOUT-.n13 GNDA 0.105329f
C1961 two_stage_opamp_dummy_magic_0.VOUT-.t5 GNDA 0.043632f
C1962 two_stage_opamp_dummy_magic_0.VOUT-.t0 GNDA 0.043632f
C1963 two_stage_opamp_dummy_magic_0.VOUT-.n14 GNDA 0.172903f
C1964 two_stage_opamp_dummy_magic_0.VOUT-.n15 GNDA 0.212301f
C1965 two_stage_opamp_dummy_magic_0.VOUT-.t101 GNDA 0.290879f
C1966 two_stage_opamp_dummy_magic_0.VOUT-.t108 GNDA 0.295834f
C1967 two_stage_opamp_dummy_magic_0.VOUT-.t149 GNDA 0.290879f
C1968 two_stage_opamp_dummy_magic_0.VOUT-.n16 GNDA 0.195025f
C1969 two_stage_opamp_dummy_magic_0.VOUT-.n17 GNDA 0.12726f
C1970 two_stage_opamp_dummy_magic_0.VOUT-.t48 GNDA 0.295213f
C1971 two_stage_opamp_dummy_magic_0.VOUT-.t92 GNDA 0.295213f
C1972 two_stage_opamp_dummy_magic_0.VOUT-.t42 GNDA 0.295213f
C1973 two_stage_opamp_dummy_magic_0.VOUT-.t130 GNDA 0.295213f
C1974 two_stage_opamp_dummy_magic_0.VOUT-.t84 GNDA 0.295213f
C1975 two_stage_opamp_dummy_magic_0.VOUT-.t125 GNDA 0.295213f
C1976 two_stage_opamp_dummy_magic_0.VOUT-.t74 GNDA 0.295213f
C1977 two_stage_opamp_dummy_magic_0.VOUT-.t23 GNDA 0.295213f
C1978 two_stage_opamp_dummy_magic_0.VOUT-.t64 GNDA 0.295213f
C1979 two_stage_opamp_dummy_magic_0.VOUT-.t150 GNDA 0.295213f
C1980 two_stage_opamp_dummy_magic_0.VOUT-.t88 GNDA 0.290879f
C1981 two_stage_opamp_dummy_magic_0.VOUT-.n18 GNDA 0.195645f
C1982 two_stage_opamp_dummy_magic_0.VOUT-.t51 GNDA 0.290879f
C1983 two_stage_opamp_dummy_magic_0.VOUT-.n19 GNDA 0.250185f
C1984 two_stage_opamp_dummy_magic_0.VOUT-.t137 GNDA 0.290879f
C1985 two_stage_opamp_dummy_magic_0.VOUT-.n20 GNDA 0.250185f
C1986 two_stage_opamp_dummy_magic_0.VOUT-.t106 GNDA 0.290879f
C1987 two_stage_opamp_dummy_magic_0.VOUT-.n21 GNDA 0.250185f
C1988 two_stage_opamp_dummy_magic_0.VOUT-.t75 GNDA 0.290879f
C1989 two_stage_opamp_dummy_magic_0.VOUT-.n22 GNDA 0.250185f
C1990 two_stage_opamp_dummy_magic_0.VOUT-.t25 GNDA 0.290879f
C1991 two_stage_opamp_dummy_magic_0.VOUT-.n23 GNDA 0.250185f
C1992 two_stage_opamp_dummy_magic_0.VOUT-.t128 GNDA 0.290879f
C1993 two_stage_opamp_dummy_magic_0.VOUT-.n24 GNDA 0.250185f
C1994 two_stage_opamp_dummy_magic_0.VOUT-.t90 GNDA 0.290879f
C1995 two_stage_opamp_dummy_magic_0.VOUT-.n25 GNDA 0.250185f
C1996 two_stage_opamp_dummy_magic_0.VOUT-.t54 GNDA 0.290879f
C1997 two_stage_opamp_dummy_magic_0.VOUT-.n26 GNDA 0.250185f
C1998 two_stage_opamp_dummy_magic_0.VOUT-.t140 GNDA 0.290879f
C1999 two_stage_opamp_dummy_magic_0.VOUT-.n27 GNDA 0.250185f
C2000 two_stage_opamp_dummy_magic_0.VOUT-.t110 GNDA 0.290879f
C2001 two_stage_opamp_dummy_magic_0.VOUT-.t28 GNDA 0.295834f
C2002 two_stage_opamp_dummy_magic_0.VOUT-.t79 GNDA 0.290879f
C2003 two_stage_opamp_dummy_magic_0.VOUT-.n28 GNDA 0.195025f
C2004 two_stage_opamp_dummy_magic_0.VOUT-.n29 GNDA 0.236339f
C2005 two_stage_opamp_dummy_magic_0.VOUT-.t24 GNDA 0.295834f
C2006 two_stage_opamp_dummy_magic_0.VOUT-.t113 GNDA 0.290879f
C2007 two_stage_opamp_dummy_magic_0.VOUT-.n30 GNDA 0.195025f
C2008 two_stage_opamp_dummy_magic_0.VOUT-.t78 GNDA 0.290879f
C2009 two_stage_opamp_dummy_magic_0.VOUT-.t129 GNDA 0.295834f
C2010 two_stage_opamp_dummy_magic_0.VOUT-.t38 GNDA 0.290879f
C2011 two_stage_opamp_dummy_magic_0.VOUT-.n31 GNDA 0.195025f
C2012 two_stage_opamp_dummy_magic_0.VOUT-.n32 GNDA 0.236339f
C2013 two_stage_opamp_dummy_magic_0.VOUT-.t61 GNDA 0.295834f
C2014 two_stage_opamp_dummy_magic_0.VOUT-.t147 GNDA 0.290879f
C2015 two_stage_opamp_dummy_magic_0.VOUT-.n33 GNDA 0.195025f
C2016 two_stage_opamp_dummy_magic_0.VOUT-.t117 GNDA 0.290879f
C2017 two_stage_opamp_dummy_magic_0.VOUT-.t32 GNDA 0.295834f
C2018 two_stage_opamp_dummy_magic_0.VOUT-.t83 GNDA 0.290879f
C2019 two_stage_opamp_dummy_magic_0.VOUT-.n34 GNDA 0.195025f
C2020 two_stage_opamp_dummy_magic_0.VOUT-.n35 GNDA 0.236339f
C2021 two_stage_opamp_dummy_magic_0.VOUT-.t100 GNDA 0.295834f
C2022 two_stage_opamp_dummy_magic_0.VOUT-.t47 GNDA 0.290879f
C2023 two_stage_opamp_dummy_magic_0.VOUT-.n36 GNDA 0.195025f
C2024 two_stage_opamp_dummy_magic_0.VOUT-.t153 GNDA 0.290879f
C2025 two_stage_opamp_dummy_magic_0.VOUT-.t71 GNDA 0.295834f
C2026 two_stage_opamp_dummy_magic_0.VOUT-.t123 GNDA 0.290879f
C2027 two_stage_opamp_dummy_magic_0.VOUT-.n37 GNDA 0.195025f
C2028 two_stage_opamp_dummy_magic_0.VOUT-.n38 GNDA 0.236339f
C2029 two_stage_opamp_dummy_magic_0.VOUT-.t69 GNDA 0.295834f
C2030 two_stage_opamp_dummy_magic_0.VOUT-.t154 GNDA 0.290879f
C2031 two_stage_opamp_dummy_magic_0.VOUT-.n39 GNDA 0.195025f
C2032 two_stage_opamp_dummy_magic_0.VOUT-.t124 GNDA 0.290879f
C2033 two_stage_opamp_dummy_magic_0.VOUT-.t35 GNDA 0.295834f
C2034 two_stage_opamp_dummy_magic_0.VOUT-.t86 GNDA 0.290879f
C2035 two_stage_opamp_dummy_magic_0.VOUT-.n40 GNDA 0.195025f
C2036 two_stage_opamp_dummy_magic_0.VOUT-.n41 GNDA 0.236339f
C2037 two_stage_opamp_dummy_magic_0.VOUT-.t96 GNDA 0.290879f
C2038 two_stage_opamp_dummy_magic_0.VOUT-.t85 GNDA 0.295834f
C2039 two_stage_opamp_dummy_magic_0.VOUT-.t57 GNDA 0.290879f
C2040 two_stage_opamp_dummy_magic_0.VOUT-.n42 GNDA 0.195025f
C2041 two_stage_opamp_dummy_magic_0.VOUT-.n43 GNDA 0.12726f
C2042 two_stage_opamp_dummy_magic_0.VOUT-.t132 GNDA 0.295213f
C2043 two_stage_opamp_dummy_magic_0.VOUT-.t115 GNDA 0.295213f
C2044 two_stage_opamp_dummy_magic_0.VOUT-.t131 GNDA 0.295834f
C2045 two_stage_opamp_dummy_magic_0.VOUT-.t104 GNDA 0.290879f
C2046 two_stage_opamp_dummy_magic_0.VOUT-.n44 GNDA 0.195025f
C2047 two_stage_opamp_dummy_magic_0.VOUT-.t73 GNDA 0.290879f
C2048 two_stage_opamp_dummy_magic_0.VOUT-.n45 GNDA 0.122715f
C2049 two_stage_opamp_dummy_magic_0.VOUT-.t146 GNDA 0.295213f
C2050 two_stage_opamp_dummy_magic_0.VOUT-.t31 GNDA 0.295834f
C2051 two_stage_opamp_dummy_magic_0.VOUT-.t138 GNDA 0.290879f
C2052 two_stage_opamp_dummy_magic_0.VOUT-.n46 GNDA 0.195025f
C2053 two_stage_opamp_dummy_magic_0.VOUT-.t107 GNDA 0.290879f
C2054 two_stage_opamp_dummy_magic_0.VOUT-.n47 GNDA 0.122715f
C2055 two_stage_opamp_dummy_magic_0.VOUT-.t46 GNDA 0.295213f
C2056 two_stage_opamp_dummy_magic_0.VOUT-.t62 GNDA 0.295834f
C2057 two_stage_opamp_dummy_magic_0.VOUT-.t41 GNDA 0.290879f
C2058 two_stage_opamp_dummy_magic_0.VOUT-.n48 GNDA 0.195025f
C2059 two_stage_opamp_dummy_magic_0.VOUT-.t143 GNDA 0.290879f
C2060 two_stage_opamp_dummy_magic_0.VOUT-.n49 GNDA 0.122715f
C2061 two_stage_opamp_dummy_magic_0.VOUT-.t87 GNDA 0.295213f
C2062 two_stage_opamp_dummy_magic_0.VOUT-.t114 GNDA 0.295834f
C2063 two_stage_opamp_dummy_magic_0.VOUT-.t21 GNDA 0.290879f
C2064 two_stage_opamp_dummy_magic_0.VOUT-.n50 GNDA 0.195025f
C2065 two_stage_opamp_dummy_magic_0.VOUT-.t126 GNDA 0.290879f
C2066 two_stage_opamp_dummy_magic_0.VOUT-.n51 GNDA 0.122715f
C2067 two_stage_opamp_dummy_magic_0.VOUT-.t65 GNDA 0.295213f
C2068 two_stage_opamp_dummy_magic_0.VOUT-.t26 GNDA 0.295457f
C2069 two_stage_opamp_dummy_magic_0.VOUT-.t102 GNDA 0.295213f
C2070 two_stage_opamp_dummy_magic_0.VOUT-.t59 GNDA 0.295457f
C2071 two_stage_opamp_dummy_magic_0.VOUT-.t134 GNDA 0.295213f
C2072 two_stage_opamp_dummy_magic_0.VOUT-.t37 GNDA 0.295457f
C2073 two_stage_opamp_dummy_magic_0.VOUT-.t120 GNDA 0.295213f
C2074 two_stage_opamp_dummy_magic_0.VOUT-.t81 GNDA 0.295457f
C2075 two_stage_opamp_dummy_magic_0.VOUT-.t155 GNDA 0.295213f
C2076 two_stage_opamp_dummy_magic_0.VOUT-.t119 GNDA 0.290879f
C2077 two_stage_opamp_dummy_magic_0.VOUT-.n52 GNDA 0.321963f
C2078 two_stage_opamp_dummy_magic_0.VOUT-.t82 GNDA 0.290879f
C2079 two_stage_opamp_dummy_magic_0.VOUT-.n53 GNDA 0.376503f
C2080 two_stage_opamp_dummy_magic_0.VOUT-.t97 GNDA 0.290879f
C2081 two_stage_opamp_dummy_magic_0.VOUT-.n54 GNDA 0.376503f
C2082 two_stage_opamp_dummy_magic_0.VOUT-.t63 GNDA 0.290879f
C2083 two_stage_opamp_dummy_magic_0.VOUT-.n55 GNDA 0.376503f
C2084 two_stage_opamp_dummy_magic_0.VOUT-.t27 GNDA 0.290879f
C2085 two_stage_opamp_dummy_magic_0.VOUT-.n56 GNDA 0.30927f
C2086 two_stage_opamp_dummy_magic_0.VOUT-.t45 GNDA 0.290879f
C2087 two_stage_opamp_dummy_magic_0.VOUT-.n57 GNDA 0.30927f
C2088 two_stage_opamp_dummy_magic_0.VOUT-.t144 GNDA 0.290879f
C2089 two_stage_opamp_dummy_magic_0.VOUT-.n58 GNDA 0.30927f
C2090 two_stage_opamp_dummy_magic_0.VOUT-.t112 GNDA 0.290879f
C2091 two_stage_opamp_dummy_magic_0.VOUT-.n59 GNDA 0.30927f
C2092 two_stage_opamp_dummy_magic_0.VOUT-.t76 GNDA 0.290879f
C2093 two_stage_opamp_dummy_magic_0.VOUT-.n60 GNDA 0.250185f
C2094 two_stage_opamp_dummy_magic_0.VOUT-.t93 GNDA 0.290879f
C2095 two_stage_opamp_dummy_magic_0.VOUT-.n61 GNDA 0.250185f
C2096 two_stage_opamp_dummy_magic_0.VOUT-.t56 GNDA 0.290879f
C2097 two_stage_opamp_dummy_magic_0.VOUT-.t40 GNDA 0.295834f
C2098 two_stage_opamp_dummy_magic_0.VOUT-.t19 GNDA 0.290879f
C2099 two_stage_opamp_dummy_magic_0.VOUT-.n62 GNDA 0.195025f
C2100 two_stage_opamp_dummy_magic_0.VOUT-.n63 GNDA 0.236339f
C2101 two_stage_opamp_dummy_magic_0.VOUT-.t34 GNDA 0.295834f
C2102 two_stage_opamp_dummy_magic_0.VOUT-.t52 GNDA 0.290879f
C2103 two_stage_opamp_dummy_magic_0.VOUT-.n64 GNDA 0.195025f
C2104 two_stage_opamp_dummy_magic_0.VOUT-.t156 GNDA 0.290879f
C2105 two_stage_opamp_dummy_magic_0.VOUT-.t136 GNDA 0.295834f
C2106 two_stage_opamp_dummy_magic_0.VOUT-.t121 GNDA 0.290879f
C2107 two_stage_opamp_dummy_magic_0.VOUT-.n65 GNDA 0.195025f
C2108 two_stage_opamp_dummy_magic_0.VOUT-.n66 GNDA 0.236339f
C2109 two_stage_opamp_dummy_magic_0.VOUT-.t70 GNDA 0.295834f
C2110 two_stage_opamp_dummy_magic_0.VOUT-.t89 GNDA 0.290879f
C2111 two_stage_opamp_dummy_magic_0.VOUT-.n67 GNDA 0.195025f
C2112 two_stage_opamp_dummy_magic_0.VOUT-.t50 GNDA 0.290879f
C2113 two_stage_opamp_dummy_magic_0.VOUT-.t36 GNDA 0.295834f
C2114 two_stage_opamp_dummy_magic_0.VOUT-.t151 GNDA 0.290879f
C2115 two_stage_opamp_dummy_magic_0.VOUT-.n68 GNDA 0.195025f
C2116 two_stage_opamp_dummy_magic_0.VOUT-.n69 GNDA 0.236339f
C2117 two_stage_opamp_dummy_magic_0.VOUT-.t95 GNDA 0.295834f
C2118 two_stage_opamp_dummy_magic_0.VOUT-.t43 GNDA 0.290879f
C2119 two_stage_opamp_dummy_magic_0.VOUT-.n70 GNDA 0.195025f
C2120 two_stage_opamp_dummy_magic_0.VOUT-.t145 GNDA 0.290879f
C2121 two_stage_opamp_dummy_magic_0.VOUT-.t66 GNDA 0.295834f
C2122 two_stage_opamp_dummy_magic_0.VOUT-.t118 GNDA 0.290879f
C2123 two_stage_opamp_dummy_magic_0.VOUT-.n71 GNDA 0.195025f
C2124 two_stage_opamp_dummy_magic_0.VOUT-.n72 GNDA 0.236339f
C2125 two_stage_opamp_dummy_magic_0.VOUT-.t55 GNDA 0.295834f
C2126 two_stage_opamp_dummy_magic_0.VOUT-.t141 GNDA 0.290879f
C2127 two_stage_opamp_dummy_magic_0.VOUT-.n73 GNDA 0.195025f
C2128 two_stage_opamp_dummy_magic_0.VOUT-.t111 GNDA 0.290879f
C2129 two_stage_opamp_dummy_magic_0.VOUT-.t29 GNDA 0.295834f
C2130 two_stage_opamp_dummy_magic_0.VOUT-.t80 GNDA 0.290879f
C2131 two_stage_opamp_dummy_magic_0.VOUT-.n74 GNDA 0.195025f
C2132 two_stage_opamp_dummy_magic_0.VOUT-.n75 GNDA 0.236339f
C2133 two_stage_opamp_dummy_magic_0.VOUT-.t91 GNDA 0.295834f
C2134 two_stage_opamp_dummy_magic_0.VOUT-.t39 GNDA 0.290879f
C2135 two_stage_opamp_dummy_magic_0.VOUT-.n76 GNDA 0.195025f
C2136 two_stage_opamp_dummy_magic_0.VOUT-.t139 GNDA 0.290879f
C2137 two_stage_opamp_dummy_magic_0.VOUT-.t58 GNDA 0.295834f
C2138 two_stage_opamp_dummy_magic_0.VOUT-.t109 GNDA 0.290879f
C2139 two_stage_opamp_dummy_magic_0.VOUT-.n77 GNDA 0.195025f
C2140 two_stage_opamp_dummy_magic_0.VOUT-.n78 GNDA 0.236339f
C2141 two_stage_opamp_dummy_magic_0.VOUT-.t49 GNDA 0.295834f
C2142 two_stage_opamp_dummy_magic_0.VOUT-.t135 GNDA 0.290879f
C2143 two_stage_opamp_dummy_magic_0.VOUT-.n79 GNDA 0.195025f
C2144 two_stage_opamp_dummy_magic_0.VOUT-.t103 GNDA 0.290879f
C2145 two_stage_opamp_dummy_magic_0.VOUT-.t20 GNDA 0.295834f
C2146 two_stage_opamp_dummy_magic_0.VOUT-.t72 GNDA 0.290879f
C2147 two_stage_opamp_dummy_magic_0.VOUT-.n80 GNDA 0.195025f
C2148 two_stage_opamp_dummy_magic_0.VOUT-.n81 GNDA 0.236339f
C2149 two_stage_opamp_dummy_magic_0.VOUT-.t148 GNDA 0.295834f
C2150 two_stage_opamp_dummy_magic_0.VOUT-.t99 GNDA 0.290879f
C2151 two_stage_opamp_dummy_magic_0.VOUT-.n82 GNDA 0.195025f
C2152 two_stage_opamp_dummy_magic_0.VOUT-.t68 GNDA 0.290879f
C2153 two_stage_opamp_dummy_magic_0.VOUT-.t122 GNDA 0.295834f
C2154 two_stage_opamp_dummy_magic_0.VOUT-.t33 GNDA 0.290879f
C2155 two_stage_opamp_dummy_magic_0.VOUT-.n83 GNDA 0.195025f
C2156 two_stage_opamp_dummy_magic_0.VOUT-.n84 GNDA 0.236339f
C2157 two_stage_opamp_dummy_magic_0.VOUT-.t44 GNDA 0.295834f
C2158 two_stage_opamp_dummy_magic_0.VOUT-.t133 GNDA 0.290879f
C2159 two_stage_opamp_dummy_magic_0.VOUT-.n85 GNDA 0.195025f
C2160 two_stage_opamp_dummy_magic_0.VOUT-.t98 GNDA 0.290879f
C2161 two_stage_opamp_dummy_magic_0.VOUT-.t152 GNDA 0.295834f
C2162 two_stage_opamp_dummy_magic_0.VOUT-.t67 GNDA 0.290879f
C2163 two_stage_opamp_dummy_magic_0.VOUT-.n86 GNDA 0.195025f
C2164 two_stage_opamp_dummy_magic_0.VOUT-.n87 GNDA 0.236339f
C2165 two_stage_opamp_dummy_magic_0.VOUT-.t142 GNDA 0.295834f
C2166 two_stage_opamp_dummy_magic_0.VOUT-.t94 GNDA 0.290879f
C2167 two_stage_opamp_dummy_magic_0.VOUT-.n88 GNDA 0.195025f
C2168 two_stage_opamp_dummy_magic_0.VOUT-.t60 GNDA 0.290879f
C2169 two_stage_opamp_dummy_magic_0.VOUT-.t116 GNDA 0.295834f
C2170 two_stage_opamp_dummy_magic_0.VOUT-.t30 GNDA 0.290879f
C2171 two_stage_opamp_dummy_magic_0.VOUT-.n89 GNDA 0.195025f
C2172 two_stage_opamp_dummy_magic_0.VOUT-.n90 GNDA 0.236339f
C2173 two_stage_opamp_dummy_magic_0.VOUT-.t77 GNDA 0.295834f
C2174 two_stage_opamp_dummy_magic_0.VOUT-.t127 GNDA 0.290879f
C2175 two_stage_opamp_dummy_magic_0.VOUT-.n91 GNDA 0.195025f
C2176 two_stage_opamp_dummy_magic_0.VOUT-.t22 GNDA 0.290879f
C2177 two_stage_opamp_dummy_magic_0.VOUT-.n92 GNDA 0.236339f
C2178 two_stage_opamp_dummy_magic_0.VOUT-.t53 GNDA 0.290879f
C2179 two_stage_opamp_dummy_magic_0.VOUT-.n93 GNDA 0.12726f
C2180 two_stage_opamp_dummy_magic_0.VOUT-.t105 GNDA 0.290879f
C2181 two_stage_opamp_dummy_magic_0.VOUT-.n94 GNDA 0.238316f
C2182 two_stage_opamp_dummy_magic_0.VOUT-.n95 GNDA 0.291354f
C2183 two_stage_opamp_dummy_magic_0.VOUT-.n96 GNDA 0.165389f
C2184 two_stage_opamp_dummy_magic_0.VOUT-.t18 GNDA 0.084162f
C2185 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2186 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2187 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2188 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2189 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2190 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2191 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2192 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2193 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2194 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2195 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2196 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2197 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2198 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2199 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2200 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2201 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2202 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2203 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2204 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2205 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.04969f
C2206 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.186051f
C2207 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2208 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2209 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.050131f
C2210 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2211 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2212 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2213 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.186051f
C2214 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.027755f
C2215 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2216 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2217 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2218 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2219 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2220 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2221 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2222 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2223 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2224 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2225 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2226 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2227 bgr_0.cap_res1.t6 GNDA 0.417173f
C2228 bgr_0.cap_res1.t10 GNDA 0.418684f
C2229 bgr_0.cap_res1.t0 GNDA 0.417173f
C2230 bgr_0.cap_res1.t14 GNDA 0.418684f
C2231 bgr_0.cap_res1.t3 GNDA 0.417173f
C2232 bgr_0.cap_res1.t7 GNDA 0.418684f
C2233 bgr_0.cap_res1.t15 GNDA 0.417173f
C2234 bgr_0.cap_res1.t9 GNDA 0.418684f
C2235 bgr_0.cap_res1.t8 GNDA 0.417173f
C2236 bgr_0.cap_res1.t12 GNDA 0.418684f
C2237 bgr_0.cap_res1.t1 GNDA 0.417173f
C2238 bgr_0.cap_res1.t16 GNDA 0.418684f
C2239 bgr_0.cap_res1.t13 GNDA 0.417173f
C2240 bgr_0.cap_res1.t19 GNDA 0.418684f
C2241 bgr_0.cap_res1.t5 GNDA 0.417173f
C2242 bgr_0.cap_res1.t2 GNDA 0.418684f
C2243 bgr_0.cap_res1.n0 GNDA 0.279631f
C2244 bgr_0.cap_res1.t4 GNDA 0.222685f
C2245 bgr_0.cap_res1.n1 GNDA 0.303406f
C2246 bgr_0.cap_res1.t18 GNDA 0.222685f
C2247 bgr_0.cap_res1.n2 GNDA 0.303406f
C2248 bgr_0.cap_res1.t11 GNDA 0.222685f
C2249 bgr_0.cap_res1.n3 GNDA 0.303406f
C2250 bgr_0.cap_res1.t17 GNDA 0.649059f
C2251 bgr_0.cap_res1.t20 GNDA 0.10618f
C2252 bgr_0.1st_Vout_1.n0 GNDA 0.573726f
C2253 bgr_0.1st_Vout_1.n1 GNDA 1.42916f
C2254 bgr_0.1st_Vout_1.n2 GNDA 1.78489f
C2255 bgr_0.1st_Vout_1.n3 GNDA 0.125562f
C2256 bgr_0.1st_Vout_1.t20 GNDA 0.352846f
C2257 bgr_0.1st_Vout_1.t11 GNDA 0.346937f
C2258 bgr_0.1st_Vout_1.t32 GNDA 0.346937f
C2259 bgr_0.1st_Vout_1.t29 GNDA 0.352846f
C2260 bgr_0.1st_Vout_1.t34 GNDA 0.346937f
C2261 bgr_0.1st_Vout_1.t25 GNDA 0.352846f
C2262 bgr_0.1st_Vout_1.t21 GNDA 0.346937f
C2263 bgr_0.1st_Vout_1.t12 GNDA 0.346937f
C2264 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C2265 bgr_0.1st_Vout_1.t16 GNDA 0.346937f
C2266 bgr_0.1st_Vout_1.t33 GNDA 0.352846f
C2267 bgr_0.1st_Vout_1.t26 GNDA 0.346937f
C2268 bgr_0.1st_Vout_1.t22 GNDA 0.346937f
C2269 bgr_0.1st_Vout_1.t17 GNDA 0.352846f
C2270 bgr_0.1st_Vout_1.t24 GNDA 0.346937f
C2271 bgr_0.1st_Vout_1.t28 GNDA 0.352846f
C2272 bgr_0.1st_Vout_1.t23 GNDA 0.346937f
C2273 bgr_0.1st_Vout_1.t13 GNDA 0.346937f
C2274 bgr_0.1st_Vout_1.t18 GNDA 0.346937f
C2275 bgr_0.1st_Vout_1.t36 GNDA 0.346937f
C2276 bgr_0.1st_Vout_1.t30 GNDA 0.022665f
C2277 bgr_0.1st_Vout_1.n4 GNDA 0.021864f
C2278 bgr_0.1st_Vout_1.t14 GNDA 0.013213f
C2279 bgr_0.1st_Vout_1.t31 GNDA 0.013213f
C2280 bgr_0.1st_Vout_1.n5 GNDA 0.029393f
C2281 bgr_0.1st_Vout_1.t6 GNDA 0.018268f
C2282 bgr_0.1st_Vout_1.n6 GNDA 0.012529f
C2283 bgr_0.1st_Vout_1.n7 GNDA 0.189508f
C2284 bgr_0.1st_Vout_1.n8 GNDA 0.011336f
C2285 bgr_0.1st_Vout_1.n9 GNDA 0.020958f
C2286 bgr_0.1st_Vout_1.t19 GNDA 0.013213f
C2287 bgr_0.1st_Vout_1.t27 GNDA 0.013213f
C2288 bgr_0.1st_Vout_1.n10 GNDA 0.029393f
C2289 bgr_0.1st_Vout_1.n11 GNDA 0.021864f
C2290 bgr_0.1st_Vout_1.t15 GNDA 0.020738f
C2291 VDDA.t231 GNDA 0.020165f
C2292 VDDA.t43 GNDA 0.020165f
C2293 VDDA.n0 GNDA 0.083391f
C2294 VDDA.t2 GNDA 0.020165f
C2295 VDDA.t244 GNDA 0.020165f
C2296 VDDA.n1 GNDA 0.083071f
C2297 VDDA.n2 GNDA 0.115173f
C2298 VDDA.t123 GNDA 0.020165f
C2299 VDDA.t54 GNDA 0.020165f
C2300 VDDA.n3 GNDA 0.083071f
C2301 VDDA.n4 GNDA 0.060099f
C2302 VDDA.t190 GNDA 0.020165f
C2303 VDDA.t234 GNDA 0.020165f
C2304 VDDA.n5 GNDA 0.083071f
C2305 VDDA.n6 GNDA 0.060099f
C2306 VDDA.t18 GNDA 0.020165f
C2307 VDDA.t113 GNDA 0.020165f
C2308 VDDA.n7 GNDA 0.083071f
C2309 VDDA.n8 GNDA 0.060099f
C2310 VDDA.t247 GNDA 0.020165f
C2311 VDDA.t245 GNDA 0.020165f
C2312 VDDA.n9 GNDA 0.083071f
C2313 VDDA.n10 GNDA 0.142818f
C2314 VDDA.n11 GNDA 0.065115f
C2315 VDDA.n12 GNDA 0.173839f
C2316 VDDA.t305 GNDA 0.012665f
C2317 VDDA.n13 GNDA 0.026949f
C2318 VDDA.t414 GNDA 0.012665f
C2319 VDDA.n14 GNDA 0.026949f
C2320 VDDA.n15 GNDA 0.039129f
C2321 VDDA.n16 GNDA 0.065768f
C2322 VDDA.n17 GNDA 0.175274f
C2323 VDDA.t375 GNDA 0.012665f
C2324 VDDA.n18 GNDA 0.026949f
C2325 VDDA.t348 GNDA 0.012665f
C2326 VDDA.n19 GNDA 0.026949f
C2327 VDDA.n20 GNDA 0.036465f
C2328 VDDA.n21 GNDA 0.045265f
C2329 VDDA.n22 GNDA 0.175274f
C2330 VDDA.t347 GNDA 0.170508f
C2331 VDDA.t55 GNDA 0.105361f
C2332 VDDA.t87 GNDA 0.105361f
C2333 VDDA.t81 GNDA 0.105361f
C2334 VDDA.t82 GNDA 0.105361f
C2335 VDDA.t8 GNDA 0.079021f
C2336 VDDA.t374 GNDA 0.170508f
C2337 VDDA.t56 GNDA 0.105361f
C2338 VDDA.t118 GNDA 0.105361f
C2339 VDDA.t83 GNDA 0.105361f
C2340 VDDA.t139 GNDA 0.105361f
C2341 VDDA.t102 GNDA 0.079021f
C2342 VDDA.n23 GNDA 0.06642f
C2343 VDDA.n24 GNDA 0.05268f
C2344 VDDA.n25 GNDA 0.06642f
C2345 VDDA.n26 GNDA 0.044363f
C2346 VDDA.n27 GNDA 0.035893f
C2347 VDDA.n28 GNDA 0.083457f
C2348 VDDA.n29 GNDA 0.083457f
C2349 VDDA.n30 GNDA 0.173839f
C2350 VDDA.t413 GNDA 0.16707f
C2351 VDDA.t215 GNDA 0.103513f
C2352 VDDA.t416 GNDA 0.103513f
C2353 VDDA.t436 GNDA 0.103513f
C2354 VDDA.t216 GNDA 0.103513f
C2355 VDDA.t75 GNDA 0.077634f
C2356 VDDA.t304 GNDA 0.16707f
C2357 VDDA.t415 GNDA 0.103513f
C2358 VDDA.t46 GNDA 0.103513f
C2359 VDDA.t7 GNDA 0.103513f
C2360 VDDA.t457 GNDA 0.103513f
C2361 VDDA.t212 GNDA 0.077634f
C2362 VDDA.n31 GNDA 0.06642f
C2363 VDDA.n32 GNDA 0.051756f
C2364 VDDA.n33 GNDA 0.06642f
C2365 VDDA.n34 GNDA 0.044151f
C2366 VDDA.n35 GNDA 0.035893f
C2367 VDDA.n36 GNDA 0.069486f
C2368 VDDA.n37 GNDA 0.206502f
C2369 VDDA.t53 GNDA 0.04033f
C2370 VDDA.t51 GNDA 0.04033f
C2371 VDDA.n38 GNDA 0.161797f
C2372 VDDA.n39 GNDA 0.082197f
C2373 VDDA.t311 GNDA 0.040175f
C2374 VDDA.n40 GNDA 0.081529f
C2375 VDDA.n41 GNDA 0.054401f
C2376 VDDA.n42 GNDA 0.076787f
C2377 VDDA.t351 GNDA 0.044619f
C2378 VDDA.t349 GNDA 0.019539f
C2379 VDDA.n43 GNDA 0.070778f
C2380 VDDA.n44 GNDA 0.041667f
C2381 VDDA.t317 GNDA 0.044619f
C2382 VDDA.t315 GNDA 0.019539f
C2383 VDDA.n45 GNDA 0.070778f
C2384 VDDA.n46 GNDA 0.041667f
C2385 VDDA.n47 GNDA 0.044363f
C2386 VDDA.n48 GNDA 0.076787f
C2387 VDDA.n49 GNDA 0.221983f
C2388 VDDA.t316 GNDA 0.274919f
C2389 VDDA.t124 GNDA 0.158966f
C2390 VDDA.t49 GNDA 0.158966f
C2391 VDDA.t3 GNDA 0.158966f
C2392 VDDA.t6 GNDA 0.158966f
C2393 VDDA.t115 GNDA 0.119224f
C2394 VDDA.n50 GNDA 0.079483f
C2395 VDDA.t114 GNDA 0.119224f
C2396 VDDA.t106 GNDA 0.158966f
C2397 VDDA.t11 GNDA 0.158966f
C2398 VDDA.t235 GNDA 0.158966f
C2399 VDDA.t191 GNDA 0.158966f
C2400 VDDA.t350 GNDA 0.274919f
C2401 VDDA.n51 GNDA 0.221983f
C2402 VDDA.n52 GNDA 0.054401f
C2403 VDDA.n53 GNDA 0.102943f
C2404 VDDA.t339 GNDA 0.040175f
C2405 VDDA.t5 GNDA 0.04033f
C2406 VDDA.t17 GNDA 0.04033f
C2407 VDDA.n54 GNDA 0.161797f
C2408 VDDA.n55 GNDA 0.082197f
C2409 VDDA.t105 GNDA 0.04033f
C2410 VDDA.t10 GNDA 0.04033f
C2411 VDDA.n56 GNDA 0.161797f
C2412 VDDA.n57 GNDA 0.082197f
C2413 VDDA.t233 GNDA 0.04033f
C2414 VDDA.t122 GNDA 0.04033f
C2415 VDDA.n58 GNDA 0.161797f
C2416 VDDA.n59 GNDA 0.082197f
C2417 VDDA.t126 GNDA 0.04033f
C2418 VDDA.t117 GNDA 0.04033f
C2419 VDDA.n60 GNDA 0.161797f
C2420 VDDA.n61 GNDA 0.172725f
C2421 VDDA.n62 GNDA 0.130411f
C2422 VDDA.t337 GNDA 0.048747f
C2423 VDDA.n63 GNDA 0.093268f
C2424 VDDA.n64 GNDA 0.054489f
C2425 VDDA.n65 GNDA 0.35886f
C2426 VDDA.n66 GNDA 0.35886f
C2427 VDDA.t310 GNDA 0.554296f
C2428 VDDA.t52 GNDA 0.306841f
C2429 VDDA.t50 GNDA 0.306841f
C2430 VDDA.t4 GNDA 0.306841f
C2431 VDDA.t16 GNDA 0.306841f
C2432 VDDA.t104 GNDA 0.230131f
C2433 VDDA.n67 GNDA 0.081529f
C2434 VDDA.n68 GNDA 0.104499f
C2435 VDDA.n69 GNDA 0.104499f
C2436 VDDA.t338 GNDA 0.554296f
C2437 VDDA.t116 GNDA 0.306841f
C2438 VDDA.t125 GNDA 0.306841f
C2439 VDDA.t121 GNDA 0.306841f
C2440 VDDA.t232 GNDA 0.306841f
C2441 VDDA.t9 GNDA 0.230131f
C2442 VDDA.n70 GNDA 0.153421f
C2443 VDDA.n71 GNDA 0.103818f
C2444 VDDA.n72 GNDA 0.070451f
C2445 VDDA.n73 GNDA 0.054489f
C2446 VDDA.t309 GNDA 0.048747f
C2447 VDDA.n74 GNDA 0.093268f
C2448 VDDA.n75 GNDA 0.130074f
C2449 VDDA.n76 GNDA 0.115735f
C2450 VDDA.n77 GNDA 0.098471f
C2451 VDDA.t189 GNDA 0.023526f
C2452 VDDA.t228 GNDA 0.023526f
C2453 VDDA.n78 GNDA 0.081817f
C2454 VDDA.t73 GNDA 0.023526f
C2455 VDDA.t112 GNDA 0.023526f
C2456 VDDA.n79 GNDA 0.081527f
C2457 VDDA.n80 GNDA 0.153915f
C2458 VDDA.t38 GNDA 0.023526f
C2459 VDDA.t205 GNDA 0.023526f
C2460 VDDA.n81 GNDA 0.081817f
C2461 VDDA.t448 GNDA 0.023526f
C2462 VDDA.t230 GNDA 0.023526f
C2463 VDDA.n82 GNDA 0.081527f
C2464 VDDA.n83 GNDA 0.153915f
C2465 VDDA.n84 GNDA 0.021509f
C2466 VDDA.n85 GNDA 0.066975f
C2467 VDDA.n86 GNDA 0.091073f
C2468 VDDA.t405 GNDA 0.116057f
C2469 VDDA.t403 GNDA 0.040966f
C2470 VDDA.n87 GNDA 0.075712f
C2471 VDDA.n88 GNDA 0.048807f
C2472 VDDA.t360 GNDA 0.116057f
C2473 VDDA.t358 GNDA 0.040966f
C2474 VDDA.n89 GNDA 0.075712f
C2475 VDDA.n90 GNDA 0.048807f
C2476 VDDA.n91 GNDA 0.048395f
C2477 VDDA.n92 GNDA 0.091073f
C2478 VDDA.n93 GNDA 0.271412f
C2479 VDDA.t359 GNDA 0.405122f
C2480 VDDA.t188 GNDA 0.233912f
C2481 VDDA.t227 GNDA 0.233912f
C2482 VDDA.t72 GNDA 0.233912f
C2483 VDDA.t111 GNDA 0.233912f
C2484 VDDA.t200 GNDA 0.175434f
C2485 VDDA.n94 GNDA 0.116956f
C2486 VDDA.t79 GNDA 0.175434f
C2487 VDDA.t447 GNDA 0.233912f
C2488 VDDA.t229 GNDA 0.233912f
C2489 VDDA.t37 GNDA 0.233912f
C2490 VDDA.t204 GNDA 0.233912f
C2491 VDDA.t404 GNDA 0.405122f
C2492 VDDA.n95 GNDA 0.271412f
C2493 VDDA.n96 GNDA 0.066975f
C2494 VDDA.n97 GNDA 0.093761f
C2495 VDDA.t201 GNDA 0.023526f
C2496 VDDA.t80 GNDA 0.023526f
C2497 VDDA.n98 GNDA 0.076703f
C2498 VDDA.n99 GNDA 0.052351f
C2499 VDDA.n100 GNDA 0.043979f
C2500 VDDA.t218 GNDA 0.020165f
C2501 VDDA.t67 GNDA 0.020165f
C2502 VDDA.n101 GNDA 0.083391f
C2503 VDDA.t467 GNDA 0.020165f
C2504 VDDA.t76 GNDA 0.020165f
C2505 VDDA.n102 GNDA 0.083071f
C2506 VDDA.n103 GNDA 0.115173f
C2507 VDDA.t213 GNDA 0.020165f
C2508 VDDA.t437 GNDA 0.020165f
C2509 VDDA.n104 GNDA 0.083071f
C2510 VDDA.n105 GNDA 0.060099f
C2511 VDDA.t169 GNDA 0.020165f
C2512 VDDA.t456 GNDA 0.020165f
C2513 VDDA.n106 GNDA 0.083071f
C2514 VDDA.n107 GNDA 0.060099f
C2515 VDDA.t98 GNDA 0.020165f
C2516 VDDA.t417 GNDA 0.020165f
C2517 VDDA.n108 GNDA 0.083071f
C2518 VDDA.n109 GNDA 0.060099f
C2519 VDDA.t170 GNDA 0.020165f
C2520 VDDA.t171 GNDA 0.020165f
C2521 VDDA.n110 GNDA 0.083071f
C2522 VDDA.n111 GNDA 0.173573f
C2523 VDDA.t466 GNDA 0.04033f
C2524 VDDA.t220 GNDA 0.04033f
C2525 VDDA.n112 GNDA 0.161797f
C2526 VDDA.n113 GNDA 0.082197f
C2527 VDDA.t366 GNDA 0.040175f
C2528 VDDA.n114 GNDA 0.054401f
C2529 VDDA.n115 GNDA 0.076787f
C2530 VDDA.t372 GNDA 0.044619f
C2531 VDDA.t370 GNDA 0.019539f
C2532 VDDA.n116 GNDA 0.070778f
C2533 VDDA.n117 GNDA 0.041667f
C2534 VDDA.t345 GNDA 0.044619f
C2535 VDDA.t343 GNDA 0.019539f
C2536 VDDA.n118 GNDA 0.070778f
C2537 VDDA.n119 GNDA 0.041667f
C2538 VDDA.n120 GNDA 0.044363f
C2539 VDDA.n121 GNDA 0.076787f
C2540 VDDA.n122 GNDA 0.221983f
C2541 VDDA.t344 GNDA 0.274919f
C2542 VDDA.t468 GNDA 0.158966f
C2543 VDDA.t438 GNDA 0.158966f
C2544 VDDA.t158 GNDA 0.158966f
C2545 VDDA.t462 GNDA 0.158966f
C2546 VDDA.t101 GNDA 0.119224f
C2547 VDDA.n123 GNDA 0.079483f
C2548 VDDA.t217 GNDA 0.119224f
C2549 VDDA.t74 GNDA 0.158966f
C2550 VDDA.t246 GNDA 0.158966f
C2551 VDDA.t84 GNDA 0.158966f
C2552 VDDA.t449 GNDA 0.158966f
C2553 VDDA.t371 GNDA 0.274919f
C2554 VDDA.n124 GNDA 0.221983f
C2555 VDDA.n125 GNDA 0.054401f
C2556 VDDA.n126 GNDA 0.102943f
C2557 VDDA.n127 GNDA 0.070451f
C2558 VDDA.n128 GNDA 0.104499f
C2559 VDDA.n129 GNDA 0.104499f
C2560 VDDA.n130 GNDA 0.103818f
C2561 VDDA.t333 GNDA 0.040175f
C2562 VDDA.t222 GNDA 0.04033f
C2563 VDDA.t453 GNDA 0.04033f
C2564 VDDA.n131 GNDA 0.161797f
C2565 VDDA.n132 GNDA 0.082197f
C2566 VDDA.t120 GNDA 0.04033f
C2567 VDDA.t195 GNDA 0.04033f
C2568 VDDA.n133 GNDA 0.161797f
C2569 VDDA.n134 GNDA 0.082197f
C2570 VDDA.t464 GNDA 0.04033f
C2571 VDDA.t419 GNDA 0.04033f
C2572 VDDA.n135 GNDA 0.161797f
C2573 VDDA.n136 GNDA 0.082197f
C2574 VDDA.t177 GNDA 0.04033f
C2575 VDDA.t455 GNDA 0.04033f
C2576 VDDA.n137 GNDA 0.161797f
C2577 VDDA.n138 GNDA 0.172725f
C2578 VDDA.n139 GNDA 0.130411f
C2579 VDDA.t331 GNDA 0.048747f
C2580 VDDA.n140 GNDA 0.093268f
C2581 VDDA.n141 GNDA 0.054489f
C2582 VDDA.n142 GNDA 0.081529f
C2583 VDDA.n143 GNDA 0.35886f
C2584 VDDA.t332 GNDA 0.554296f
C2585 VDDA.t176 GNDA 0.306841f
C2586 VDDA.t454 GNDA 0.306841f
C2587 VDDA.t463 GNDA 0.306841f
C2588 VDDA.t418 GNDA 0.306841f
C2589 VDDA.t119 GNDA 0.230131f
C2590 VDDA.n144 GNDA 0.153421f
C2591 VDDA.t194 GNDA 0.230131f
C2592 VDDA.t221 GNDA 0.306841f
C2593 VDDA.t452 GNDA 0.306841f
C2594 VDDA.t465 GNDA 0.306841f
C2595 VDDA.t219 GNDA 0.306841f
C2596 VDDA.t365 GNDA 0.554296f
C2597 VDDA.n145 GNDA 0.35886f
C2598 VDDA.n146 GNDA 0.081529f
C2599 VDDA.n147 GNDA 0.054489f
C2600 VDDA.t364 GNDA 0.048747f
C2601 VDDA.n148 GNDA 0.093268f
C2602 VDDA.n149 GNDA 0.130074f
C2603 VDDA.n150 GNDA 0.099603f
C2604 VDDA.n152 GNDA 0.051466f
C2605 VDDA.n153 GNDA 0.063847f
C2606 VDDA.n155 GNDA 0.051466f
C2607 VDDA.n157 GNDA 0.051466f
C2608 VDDA.n159 GNDA 0.051466f
C2609 VDDA.n161 GNDA 0.051466f
C2610 VDDA.n163 GNDA 0.051466f
C2611 VDDA.n165 GNDA 0.051466f
C2612 VDDA.n167 GNDA 0.051466f
C2613 VDDA.n169 GNDA 0.051466f
C2614 VDDA.n171 GNDA 0.084219f
C2615 VDDA.t390 GNDA 0.012246f
C2616 VDDA.n172 GNDA 0.018183f
C2617 VDDA.n173 GNDA 0.016089f
C2618 VDDA.n174 GNDA 0.054949f
C2619 VDDA.n175 GNDA 0.211005f
C2620 VDDA.n176 GNDA 0.211005f
C2621 VDDA.t395 GNDA 0.16707f
C2622 VDDA.t131 GNDA 0.103513f
C2623 VDDA.t167 GNDA 0.103513f
C2624 VDDA.t94 GNDA 0.103513f
C2625 VDDA.t165 GNDA 0.103513f
C2626 VDDA.t144 GNDA 0.103513f
C2627 VDDA.t137 GNDA 0.103513f
C2628 VDDA.t159 GNDA 0.103513f
C2629 VDDA.t150 GNDA 0.103513f
C2630 VDDA.t12 GNDA 0.103513f
C2631 VDDA.t163 GNDA 0.077634f
C2632 VDDA.t389 GNDA 0.16707f
C2633 VDDA.t88 GNDA 0.103513f
C2634 VDDA.t161 GNDA 0.103513f
C2635 VDDA.t70 GNDA 0.103513f
C2636 VDDA.t148 GNDA 0.103513f
C2637 VDDA.t146 GNDA 0.103513f
C2638 VDDA.t135 GNDA 0.103513f
C2639 VDDA.t133 GNDA 0.103513f
C2640 VDDA.t14 GNDA 0.103513f
C2641 VDDA.t92 GNDA 0.103513f
C2642 VDDA.t90 GNDA 0.077634f
C2643 VDDA.n177 GNDA 0.063847f
C2644 VDDA.n178 GNDA 0.103192f
C2645 VDDA.n179 GNDA 0.103192f
C2646 VDDA.n180 GNDA 0.051756f
C2647 VDDA.n181 GNDA 0.103192f
C2648 VDDA.n182 GNDA 0.081331f
C2649 VDDA.n183 GNDA 0.054949f
C2650 VDDA.n184 GNDA 0.016089f
C2651 VDDA.t396 GNDA 0.012246f
C2652 VDDA.n185 GNDA 0.01774f
C2653 VDDA.n186 GNDA 0.063444f
C2654 VDDA.n187 GNDA 0.04974f
C2655 VDDA.n188 GNDA 0.256568f
C2656 VDDA.n189 GNDA 0.244024f
C2657 VDDA.t22 GNDA 0.023526f
C2658 VDDA.t42 GNDA 0.023526f
C2659 VDDA.n190 GNDA 0.081817f
C2660 VDDA.t24 GNDA 0.023526f
C2661 VDDA.t243 GNDA 0.023526f
C2662 VDDA.n191 GNDA 0.081527f
C2663 VDDA.n192 GNDA 0.153915f
C2664 VDDA.t1 GNDA 0.023526f
C2665 VDDA.t20 GNDA 0.023526f
C2666 VDDA.n193 GNDA 0.081817f
C2667 VDDA.t45 GNDA 0.023526f
C2668 VDDA.t209 GNDA 0.023526f
C2669 VDDA.n194 GNDA 0.081527f
C2670 VDDA.n195 GNDA 0.153915f
C2671 VDDA.n196 GNDA 0.021509f
C2672 VDDA.n197 GNDA 0.066975f
C2673 VDDA.n198 GNDA 0.091073f
C2674 VDDA.t381 GNDA 0.116057f
C2675 VDDA.t379 GNDA 0.040966f
C2676 VDDA.n199 GNDA 0.075712f
C2677 VDDA.n200 GNDA 0.048807f
C2678 VDDA.t354 GNDA 0.116057f
C2679 VDDA.t352 GNDA 0.040966f
C2680 VDDA.n201 GNDA 0.075712f
C2681 VDDA.n202 GNDA 0.048807f
C2682 VDDA.n203 GNDA 0.048395f
C2683 VDDA.n204 GNDA 0.091073f
C2684 VDDA.n205 GNDA 0.271412f
C2685 VDDA.t353 GNDA 0.405122f
C2686 VDDA.t21 GNDA 0.233912f
C2687 VDDA.t41 GNDA 0.233912f
C2688 VDDA.t23 GNDA 0.233912f
C2689 VDDA.t242 GNDA 0.233912f
C2690 VDDA.t77 GNDA 0.175434f
C2691 VDDA.n206 GNDA 0.116956f
C2692 VDDA.t225 GNDA 0.175434f
C2693 VDDA.t44 GNDA 0.233912f
C2694 VDDA.t208 GNDA 0.233912f
C2695 VDDA.t0 GNDA 0.233912f
C2696 VDDA.t19 GNDA 0.233912f
C2697 VDDA.t380 GNDA 0.405122f
C2698 VDDA.n207 GNDA 0.271412f
C2699 VDDA.n208 GNDA 0.066975f
C2700 VDDA.n209 GNDA 0.093761f
C2701 VDDA.t78 GNDA 0.023526f
C2702 VDDA.t226 GNDA 0.023526f
C2703 VDDA.n210 GNDA 0.076703f
C2704 VDDA.n211 GNDA 0.052351f
C2705 VDDA.n212 GNDA 0.043979f
C2706 VDDA.n213 GNDA 0.21077f
C2707 VDDA.n214 GNDA 0.082676f
C2708 VDDA.n216 GNDA 0.065587f
C2709 VDDA.n217 GNDA 0.012099f
C2710 VDDA.n218 GNDA 0.035739f
C2711 VDDA.n219 GNDA 0.035739f
C2712 VDDA.n220 GNDA 0.036441f
C2713 VDDA.n221 GNDA 0.091565f
C2714 VDDA.n222 GNDA 0.012099f
C2715 VDDA.n223 GNDA 0.053742f
C2716 VDDA.n224 GNDA 0.053742f
C2717 VDDA.n225 GNDA 0.053741f
C2718 VDDA.t224 GNDA 0.021509f
C2719 VDDA.n226 GNDA 0.07464f
C2720 VDDA.t363 GNDA 0.098246f
C2721 VDDA.n227 GNDA 0.048719f
C2722 VDDA.n228 GNDA 0.04677f
C2723 VDDA.t361 GNDA 0.037331f
C2724 VDDA.n229 GNDA 0.039523f
C2725 VDDA.n230 GNDA 0.029584f
C2726 VDDA.n231 GNDA 0.045968f
C2727 VDDA.n232 GNDA 0.301361f
C2728 VDDA.t362 GNDA 0.286468f
C2729 VDDA.n233 GNDA 0.093262f
C2730 VDDA.n234 GNDA 0.023316f
C2731 VDDA.t223 GNDA 0.130567f
C2732 VDDA.t383 GNDA 0.309783f
C2733 VDDA.n235 GNDA 0.304482f
C2734 VDDA.n236 GNDA 0.047699f
C2735 VDDA.n237 GNDA 0.030588f
C2736 VDDA.t382 GNDA 0.038002f
C2737 VDDA.n238 GNDA 0.039523f
C2738 VDDA.t384 GNDA 0.076737f
C2739 VDDA.n239 GNDA 0.052664f
C2740 VDDA.n240 GNDA 0.110717f
C2741 VDDA.n241 GNDA 0.072542f
C2742 VDDA.t314 GNDA 0.015711f
C2743 VDDA.n242 GNDA 0.017069f
C2744 VDDA.t312 GNDA 0.013181f
C2745 VDDA.n243 GNDA 0.016688f
C2746 VDDA.n244 GNDA 0.021487f
C2747 VDDA.n245 GNDA 0.030154f
C2748 VDDA.n246 GNDA 0.160837f
C2749 VDDA.t313 GNDA 0.178139f
C2750 VDDA.t68 GNDA 0.120989f
C2751 VDDA.t328 GNDA 0.178139f
C2752 VDDA.n247 GNDA 0.160837f
C2753 VDDA.n248 GNDA 0.030154f
C2754 VDDA.n249 GNDA 0.021487f
C2755 VDDA.t327 GNDA 0.013181f
C2756 VDDA.n250 GNDA 0.016688f
C2757 VDDA.t330 GNDA 0.015711f
C2758 VDDA.n251 GNDA 0.019053f
C2759 VDDA.n252 GNDA 0.074867f
C2760 VDDA.n253 GNDA 0.21792f
C2761 VDDA.n254 GNDA 4.448f
C2762 VDDA.t470 GNDA 0.743101f
C2763 VDDA.t471 GNDA 0.792003f
C2764 VDDA.t469 GNDA 0.792003f
C2765 VDDA.t472 GNDA 0.759459f
C2766 VDDA.n255 GNDA 0.530883f
C2767 VDDA.n256 GNDA 0.257742f
C2768 VDDA.n257 GNDA 0.330442f
C2769 VDDA.n258 GNDA 2.36084f
C2770 VDDA.n259 GNDA 0.021509f
C2771 VDDA.n260 GNDA 0.01628f
C2772 VDDA.n261 GNDA 0.01628f
C2773 VDDA.n262 GNDA 0.047576f
C2774 VDDA.n263 GNDA 0.021509f
C2775 VDDA.t342 GNDA 0.02525f
C2776 VDDA.t340 GNDA 0.016638f
C2777 VDDA.n264 GNDA 0.039611f
C2778 VDDA.n265 GNDA 0.056362f
C2779 VDDA.n266 GNDA 0.105957f
C2780 VDDA.n267 GNDA 0.105957f
C2781 VDDA.t308 GNDA 0.02525f
C2782 VDDA.t306 GNDA 0.016638f
C2783 VDDA.n268 GNDA 0.039611f
C2784 VDDA.n269 GNDA 0.080659f
C2785 VDDA.n270 GNDA 0.056362f
C2786 VDDA.n271 GNDA 0.021509f
C2787 VDDA.n272 GNDA 0.01628f
C2788 VDDA.n273 GNDA 0.017021f
C2789 VDDA.n274 GNDA 0.016906f
C2790 VDDA.n275 GNDA 0.131424f
C2791 VDDA.n276 GNDA 0.016906f
C2792 VDDA.n277 GNDA 0.068458f
C2793 VDDA.n278 GNDA 0.016906f
C2794 VDDA.n279 GNDA 0.068458f
C2795 VDDA.n280 GNDA 0.01628f
C2796 VDDA.n281 GNDA 0.066117f
C2797 VDDA.n282 GNDA 0.105957f
C2798 VDDA.t357 GNDA 0.02525f
C2799 VDDA.t355 GNDA 0.016638f
C2800 VDDA.n283 GNDA 0.039611f
C2801 VDDA.n284 GNDA 0.056362f
C2802 VDDA.t411 GNDA 0.02525f
C2803 VDDA.t409 GNDA 0.016638f
C2804 VDDA.n285 GNDA 0.039611f
C2805 VDDA.n286 GNDA 0.056362f
C2806 VDDA.n287 GNDA 0.080659f
C2807 VDDA.n288 GNDA 0.105957f
C2808 VDDA.n289 GNDA 0.230382f
C2809 VDDA.t410 GNDA 0.210127f
C2810 VDDA.t458 GNDA 0.133088f
C2811 VDDA.t35 GNDA 0.133088f
C2812 VDDA.t426 GNDA 0.133088f
C2813 VDDA.t434 GNDA 0.133088f
C2814 VDDA.t184 GNDA 0.133088f
C2815 VDDA.t25 GNDA 0.133088f
C2816 VDDA.t460 GNDA 0.133088f
C2817 VDDA.t129 GNDA 0.133088f
C2818 VDDA.t156 GNDA 0.099816f
C2819 VDDA.n290 GNDA 0.066544f
C2820 VDDA.t443 GNDA 0.099816f
C2821 VDDA.t186 GNDA 0.133088f
C2822 VDDA.t420 GNDA 0.133088f
C2823 VDDA.t422 GNDA 0.133088f
C2824 VDDA.t198 GNDA 0.133088f
C2825 VDDA.t142 GNDA 0.133088f
C2826 VDDA.t445 GNDA 0.133088f
C2827 VDDA.t109 GNDA 0.133088f
C2828 VDDA.t206 GNDA 0.133088f
C2829 VDDA.t356 GNDA 0.210127f
C2830 VDDA.n291 GNDA 0.230382f
C2831 VDDA.n292 GNDA 0.066117f
C2832 VDDA.n293 GNDA 0.112632f
C2833 VDDA.n294 GNDA 0.047576f
C2834 VDDA.n295 GNDA 0.021509f
C2835 VDDA.n296 GNDA 0.016906f
C2836 VDDA.n297 GNDA 0.068458f
C2837 VDDA.n298 GNDA 0.016906f
C2838 VDDA.n299 GNDA 0.068458f
C2839 VDDA.n300 GNDA 0.016906f
C2840 VDDA.n301 GNDA 0.068458f
C2841 VDDA.n302 GNDA 0.016906f
C2842 VDDA.n303 GNDA 0.098033f
C2843 VDDA.n304 GNDA 0.021509f
C2844 VDDA.n305 GNDA 0.01628f
C2845 VDDA.n306 GNDA 0.01628f
C2846 VDDA.n307 GNDA 0.047576f
C2847 VDDA.n308 GNDA 0.021509f
C2848 VDDA.n309 GNDA 0.01628f
C2849 VDDA.n310 GNDA 0.021509f
C2850 VDDA.n311 GNDA 0.01628f
C2851 VDDA.n312 GNDA 0.047576f
C2852 VDDA.n313 GNDA 0.021509f
C2853 VDDA.n314 GNDA 0.021509f
C2854 VDDA.n315 GNDA 0.047576f
C2855 VDDA.n316 GNDA 0.021509f
C2856 VDDA.n317 GNDA 0.021509f
C2857 VDDA.n318 GNDA 0.01628f
C2858 VDDA.n319 GNDA 0.047576f
C2859 VDDA.n320 GNDA 0.021509f
C2860 VDDA.n321 GNDA 0.021509f
C2861 VDDA.n322 GNDA 0.047576f
C2862 VDDA.n323 GNDA 0.021509f
C2863 VDDA.n324 GNDA 0.01628f
C2864 VDDA.n325 GNDA 0.047576f
C2865 VDDA.n326 GNDA 0.021509f
C2866 VDDA.n327 GNDA 0.051084f
C2867 VDDA.n328 GNDA 0.047576f
C2868 VDDA.n329 GNDA 0.035117f
C2869 VDDA.n330 GNDA 0.033543f
C2870 VDDA.n331 GNDA 0.230382f
C2871 VDDA.t307 GNDA 0.210127f
C2872 VDDA.t178 GNDA 0.133088f
C2873 VDDA.t63 GNDA 0.133088f
C2874 VDDA.t174 GNDA 0.133088f
C2875 VDDA.t236 GNDA 0.133088f
C2876 VDDA.t240 GNDA 0.133088f
C2877 VDDA.t127 GNDA 0.133088f
C2878 VDDA.t39 GNDA 0.133088f
C2879 VDDA.t59 GNDA 0.133088f
C2880 VDDA.t61 GNDA 0.099816f
C2881 VDDA.n332 GNDA 0.066544f
C2882 VDDA.t192 GNDA 0.099816f
C2883 VDDA.t107 GNDA 0.133088f
C2884 VDDA.t99 GNDA 0.133088f
C2885 VDDA.t202 GNDA 0.133088f
C2886 VDDA.t172 GNDA 0.133088f
C2887 VDDA.t57 GNDA 0.133088f
C2888 VDDA.t85 GNDA 0.133088f
C2889 VDDA.t238 GNDA 0.133088f
C2890 VDDA.t210 GNDA 0.133088f
C2891 VDDA.t341 GNDA 0.210127f
C2892 VDDA.n333 GNDA 0.230382f
C2893 VDDA.n334 GNDA 0.033543f
C2894 VDDA.n335 GNDA 0.035117f
C2895 VDDA.n336 GNDA 0.047576f
C2896 VDDA.n337 GNDA 0.065117f
C2897 VDDA.n338 GNDA 0.197698f
C2898 VDDA.t275 GNDA 0.020165f
C2899 VDDA.t273 GNDA 0.020165f
C2900 VDDA.n339 GNDA 0.066618f
C2901 VDDA.n340 GNDA 0.085962f
C2902 VDDA.t393 GNDA 0.061797f
C2903 VDDA.n341 GNDA 0.10889f
C2904 VDDA.n342 GNDA 0.148437f
C2905 VDDA.n343 GNDA 0.148437f
C2906 VDDA.n344 GNDA 0.147756f
C2907 VDDA.t336 GNDA 0.061797f
C2908 VDDA.t334 GNDA 0.096154f
C2909 VDDA.t378 GNDA 0.02525f
C2910 VDDA.t376 GNDA 0.012743f
C2911 VDDA.n345 GNDA 0.03981f
C2912 VDDA.n346 GNDA 0.022955f
C2913 VDDA.n347 GNDA 0.040797f
C2914 VDDA.t399 GNDA 0.02525f
C2915 VDDA.t397 GNDA 0.012743f
C2916 VDDA.n348 GNDA 0.03981f
C2917 VDDA.n349 GNDA 0.040797f
C2918 VDDA.n350 GNDA 0.040797f
C2919 VDDA.n351 GNDA 0.033474f
C2920 VDDA.n352 GNDA 0.160856f
C2921 VDDA.t377 GNDA 0.201979f
C2922 VDDA.t214 GNDA 0.091498f
C2923 VDDA.n353 GNDA 0.060999f
C2924 VDDA.t103 GNDA 0.091498f
C2925 VDDA.t398 GNDA 0.204958f
C2926 VDDA.n354 GNDA 0.168968f
C2927 VDDA.n355 GNDA 0.033474f
C2928 VDDA.n356 GNDA 0.022955f
C2929 VDDA.n357 GNDA 0.032249f
C2930 VDDA.t294 GNDA 0.020165f
C2931 VDDA.t255 GNDA 0.020165f
C2932 VDDA.n358 GNDA 0.066618f
C2933 VDDA.n359 GNDA 0.085962f
C2934 VDDA.t266 GNDA 0.020165f
C2935 VDDA.t285 GNDA 0.020165f
C2936 VDDA.n360 GNDA 0.066618f
C2937 VDDA.n361 GNDA 0.085962f
C2938 VDDA.t250 GNDA 0.020165f
C2939 VDDA.t269 GNDA 0.020165f
C2940 VDDA.n362 GNDA 0.066618f
C2941 VDDA.n363 GNDA 0.085962f
C2942 VDDA.t283 GNDA 0.020165f
C2943 VDDA.t291 GNDA 0.020165f
C2944 VDDA.n364 GNDA 0.066618f
C2945 VDDA.n365 GNDA 0.085962f
C2946 VDDA.t264 GNDA 0.020165f
C2947 VDDA.t260 GNDA 0.020165f
C2948 VDDA.n366 GNDA 0.066618f
C2949 VDDA.n367 GNDA 0.085962f
C2950 VDDA.t289 GNDA 0.020165f
C2951 VDDA.t299 GNDA 0.020165f
C2952 VDDA.n368 GNDA 0.066618f
C2953 VDDA.n369 GNDA 0.085962f
C2954 VDDA.t257 GNDA 0.020165f
C2955 VDDA.t278 GNDA 0.020165f
C2956 VDDA.n370 GNDA 0.066618f
C2957 VDDA.n371 GNDA 0.085962f
C2958 VDDA.n372 GNDA 0.094912f
C2959 VDDA.n373 GNDA 0.114756f
C2960 VDDA.n374 GNDA 0.077351f
C2961 VDDA.n375 GNDA 0.09444f
C2962 VDDA.n376 GNDA 0.347967f
C2963 VDDA.t335 GNDA 0.448994f
C2964 VDDA.t256 GNDA 0.323645f
C2965 VDDA.t277 GNDA 0.323645f
C2966 VDDA.t288 GNDA 0.323645f
C2967 VDDA.t298 GNDA 0.323645f
C2968 VDDA.t263 GNDA 0.323645f
C2969 VDDA.t259 GNDA 0.323645f
C2970 VDDA.t282 GNDA 0.323645f
C2971 VDDA.t290 GNDA 0.242734f
C2972 VDDA.n377 GNDA 0.161823f
C2973 VDDA.t249 GNDA 0.242734f
C2974 VDDA.t268 GNDA 0.323645f
C2975 VDDA.t265 GNDA 0.323645f
C2976 VDDA.t284 GNDA 0.323645f
C2977 VDDA.t293 GNDA 0.323645f
C2978 VDDA.t254 GNDA 0.323645f
C2979 VDDA.t274 GNDA 0.323645f
C2980 VDDA.t272 GNDA 0.323645f
C2981 VDDA.t392 GNDA 0.448994f
C2982 VDDA.n378 GNDA 0.347967f
C2983 VDDA.n379 GNDA 0.09444f
C2984 VDDA.n380 GNDA 0.077351f
C2985 VDDA.t391 GNDA 0.096154f
C2986 VDDA.n381 GNDA 0.114756f
C2987 VDDA.n382 GNDA 0.052678f
C2988 VDDA.n383 GNDA 0.016233f
C2989 VDDA.t323 GNDA 0.025438f
C2990 VDDA.t321 GNDA 0.012413f
C2991 VDDA.n384 GNDA 0.038104f
C2992 VDDA.n385 GNDA 0.02285f
C2993 VDDA.n386 GNDA 0.040797f
C2994 VDDA.t320 GNDA 0.025438f
C2995 VDDA.t318 GNDA 0.012413f
C2996 VDDA.n387 GNDA 0.038104f
C2997 VDDA.n388 GNDA 0.040797f
C2998 VDDA.n389 GNDA 0.040797f
C2999 VDDA.n390 GNDA 0.033474f
C3000 VDDA.n391 GNDA 0.160856f
C3001 VDDA.t322 GNDA 0.201979f
C3002 VDDA.t65 GNDA 0.091498f
C3003 VDDA.n392 GNDA 0.060999f
C3004 VDDA.t432 GNDA 0.091498f
C3005 VDDA.t319 GNDA 0.201979f
C3006 VDDA.n393 GNDA 0.160856f
C3007 VDDA.n394 GNDA 0.033474f
C3008 VDDA.n395 GNDA 0.02285f
C3009 VDDA.n396 GNDA 0.024006f
C3010 VDDA.n397 GNDA 0.044933f
C3011 VDDA.n398 GNDA 0.094669f
C3012 VDDA.n399 GNDA 0.16439f
C3013 VDDA.n400 GNDA 0.016767f
C3014 VDDA.n401 GNDA 0.059187f
C3015 VDDA.t326 GNDA 0.026527f
C3016 VDDA.n402 GNDA 0.022181f
C3017 VDDA.n403 GNDA 0.048012f
C3018 VDDA.n404 GNDA 0.048012f
C3019 VDDA.n405 GNDA 0.048011f
C3020 VDDA.t387 GNDA 0.026527f
C3021 VDDA.t385 GNDA 0.013237f
C3022 VDDA.n406 GNDA 0.016736f
C3023 VDDA.n407 GNDA 0.059218f
C3024 VDDA.t402 GNDA 0.025315f
C3025 VDDA.n408 GNDA 0.044363f
C3026 VDDA.n409 GNDA 0.069893f
C3027 VDDA.n410 GNDA 0.069893f
C3028 VDDA.n411 GNDA 0.069893f
C3029 VDDA.t408 GNDA 0.025315f
C3030 VDDA.t406 GNDA 0.013237f
C3031 VDDA.n412 GNDA 0.016774f
C3032 VDDA.n413 GNDA 0.05918f
C3033 VDDA.t369 GNDA 0.026538f
C3034 VDDA.n414 GNDA 0.022181f
C3035 VDDA.n415 GNDA 0.048011f
C3036 VDDA.n416 GNDA 0.048011f
C3037 VDDA.n417 GNDA 0.048011f
C3038 VDDA.t302 GNDA 0.026538f
C3039 VDDA.t300 GNDA 0.013237f
C3040 VDDA.n418 GNDA 0.016774f
C3041 VDDA.n419 GNDA 0.080998f
C3042 VDDA.n420 GNDA 0.045449f
C3043 VDDA.n421 GNDA 0.027123f
C3044 VDDA.n422 GNDA 0.037261f
C3045 VDDA.n423 GNDA 0.16975f
C3046 VDDA.t301 GNDA 0.205532f
C3047 VDDA.t424 GNDA 0.123846f
C3048 VDDA.t182 GNDA 0.092884f
C3049 VDDA.n424 GNDA 0.061923f
C3050 VDDA.t27 GNDA 0.092884f
C3051 VDDA.t29 GNDA 0.123846f
C3052 VDDA.t368 GNDA 0.205532f
C3053 VDDA.n425 GNDA 0.16975f
C3054 VDDA.n426 GNDA 0.037261f
C3055 VDDA.n427 GNDA 0.027123f
C3056 VDDA.t367 GNDA 0.013657f
C3057 VDDA.n428 GNDA 0.04498f
C3058 VDDA.n429 GNDA 0.040856f
C3059 VDDA.n430 GNDA 0.016736f
C3060 VDDA.n431 GNDA 0.059218f
C3061 VDDA.n432 GNDA 0.016736f
C3062 VDDA.n433 GNDA 0.059218f
C3063 VDDA.n434 GNDA 0.016736f
C3064 VDDA.n435 GNDA 0.059218f
C3065 VDDA.n436 GNDA 0.016736f
C3066 VDDA.n437 GNDA 0.059218f
C3067 VDDA.n438 GNDA 0.040856f
C3068 VDDA.n439 GNDA 0.045782f
C3069 VDDA.n440 GNDA 0.04191f
C3070 VDDA.n441 GNDA 0.052234f
C3071 VDDA.n442 GNDA 0.199695f
C3072 VDDA.t407 GNDA 0.205532f
C3073 VDDA.t33 GNDA 0.123846f
C3074 VDDA.t450 GNDA 0.123846f
C3075 VDDA.t180 GNDA 0.123846f
C3076 VDDA.t31 GNDA 0.123846f
C3077 VDDA.t47 GNDA 0.123846f
C3078 VDDA.t152 GNDA 0.092884f
C3079 VDDA.n443 GNDA 0.061923f
C3080 VDDA.t140 GNDA 0.092884f
C3081 VDDA.t441 GNDA 0.123846f
C3082 VDDA.t428 GNDA 0.123846f
C3083 VDDA.t154 GNDA 0.123846f
C3084 VDDA.t401 GNDA 0.205532f
C3085 VDDA.n444 GNDA 0.184767f
C3086 VDDA.n445 GNDA 0.044769f
C3087 VDDA.n446 GNDA 0.034516f
C3088 VDDA.t400 GNDA 0.013237f
C3089 VDDA.n447 GNDA 0.045782f
C3090 VDDA.n448 GNDA 0.048249f
C3091 VDDA.n449 GNDA 0.016767f
C3092 VDDA.n450 GNDA 0.059187f
C3093 VDDA.n451 GNDA 0.048249f
C3094 VDDA.n452 GNDA 0.04457f
C3095 VDDA.n453 GNDA 0.027123f
C3096 VDDA.n454 GNDA 0.036746f
C3097 VDDA.n455 GNDA 0.167915f
C3098 VDDA.t386 GNDA 0.201979f
C3099 VDDA.t430 GNDA 0.121997f
C3100 VDDA.t96 GNDA 0.08318f
C3101 VDDA.n456 GNDA 0.030499f
C3102 VDDA.n457 GNDA 0.038817f
C3103 VDDA.t196 GNDA 0.091498f
C3104 VDDA.t439 GNDA 0.121997f
C3105 VDDA.t325 GNDA 0.201979f
C3106 VDDA.n458 GNDA 0.168943f
C3107 VDDA.n459 GNDA 0.037775f
C3108 VDDA.n460 GNDA 0.027123f
C3109 VDDA.t324 GNDA 0.013237f
C3110 VDDA.n461 GNDA 0.04457f
C3111 VDDA.n462 GNDA 0.088897f
C3112 VDDA.n463 GNDA 0.133442f
C3113 VDDA.t287 GNDA 0.375738f
C3114 VDDA.t295 GNDA 0.377099f
C3115 VDDA.t267 GNDA 0.375738f
C3116 VDDA.t251 GNDA 0.377099f
C3117 VDDA.t276 GNDA 0.375738f
C3118 VDDA.t280 GNDA 0.377099f
C3119 VDDA.t252 GNDA 0.375738f
C3120 VDDA.t292 GNDA 0.377099f
C3121 VDDA.t281 GNDA 0.375738f
C3122 VDDA.t297 GNDA 0.377099f
C3123 VDDA.t270 GNDA 0.375738f
C3124 VDDA.t253 GNDA 0.377099f
C3125 VDDA.t248 GNDA 0.375738f
C3126 VDDA.t262 GNDA 0.377099f
C3127 VDDA.t286 GNDA 0.375738f
C3128 VDDA.t271 GNDA 0.377099f
C3129 VDDA.n464 GNDA 0.251857f
C3130 VDDA.t279 GNDA 0.200567f
C3131 VDDA.n465 GNDA 0.273271f
C3132 VDDA.t261 GNDA 0.200567f
C3133 VDDA.n466 GNDA 0.273271f
C3134 VDDA.t296 GNDA 0.200567f
C3135 VDDA.n467 GNDA 0.273271f
C3136 VDDA.t258 GNDA 0.299287f
C3137 VDDA.n468 GNDA 0.260791f
C3138 VDDA.n469 GNDA 0.810475f
C3139 bgr_0.Vin-.n0 GNDA 0.073641f
C3140 bgr_0.Vin-.n1 GNDA 0.082742f
C3141 bgr_0.Vin-.n2 GNDA 0.998979f
C3142 bgr_0.Vin-.t5 GNDA 0.028614f
C3143 bgr_0.Vin-.t4 GNDA 0.028614f
C3144 bgr_0.Vin-.n3 GNDA 0.099613f
C3145 bgr_0.Vin-.t3 GNDA 0.028614f
C3146 bgr_0.Vin-.t6 GNDA 0.028614f
C3147 bgr_0.Vin-.n4 GNDA 0.095121f
C3148 bgr_0.Vin-.n5 GNDA 0.408067f
C3149 bgr_0.Vin-.t7 GNDA 0.098662f
C3150 bgr_0.Vin-.n6 GNDA 0.025702f
C3151 bgr_0.Vin-.n7 GNDA 0.469862f
C3152 bgr_0.Vin-.n8 GNDA 0.222852f
C3153 bgr_0.Vin-.t10 GNDA 0.023594f
C3154 bgr_0.Vin-.n9 GNDA 0.027673f
C3155 bgr_0.Vin-.n10 GNDA 0.022653f
C3156 bgr_0.Vin-.n11 GNDA 0.022653f
C3157 bgr_0.Vin-.n12 GNDA 0.040466f
C3158 bgr_0.Vin-.n13 GNDA 0.524007f
C3159 bgr_0.Vin-.t2 GNDA 0.276208f
C3160 bgr_0.Vin-.n14 GNDA 0.510829f
C3161 bgr_0.Vin-.n15 GNDA 0.074468f
C3162 bgr_0.Vin-.n16 GNDA 0.126176f
C3163 bgr_0.Vin-.n17 GNDA 0.073776f
C3164 bgr_0.Vin-.n18 GNDA 0.145931f
C3165 bgr_0.Vin-.n19 GNDA 0.145931f
C3166 bgr_0.Vin-.n20 GNDA -5.06787f
C3167 bgr_0.Vin-.n21 GNDA 5.25363f
C3168 bgr_0.Vin-.n22 GNDA 0.222489f
C3169 bgr_0.Vin-.n23 GNDA 0.382836f
C3170 bgr_0.Vin-.n24 GNDA 0.166915f
C3171 bgr_0.Vin-.n25 GNDA 0.040544f
C3172 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.043026f
C3173 bgr_0.V_TOP.t31 GNDA 0.115045f
C3174 bgr_0.V_TOP.t44 GNDA 0.115045f
C3175 bgr_0.V_TOP.t18 GNDA 0.115045f
C3176 bgr_0.V_TOP.t26 GNDA 0.115045f
C3177 bgr_0.V_TOP.t37 GNDA 0.115045f
C3178 bgr_0.V_TOP.t35 GNDA 0.115045f
C3179 bgr_0.V_TOP.t48 GNDA 0.115045f
C3180 bgr_0.V_TOP.t20 GNDA 0.115045f
C3181 bgr_0.V_TOP.t27 GNDA 0.115045f
C3182 bgr_0.V_TOP.t41 GNDA 0.115045f
C3183 bgr_0.V_TOP.t38 GNDA 0.115045f
C3184 bgr_0.V_TOP.t14 GNDA 0.115045f
C3185 bgr_0.V_TOP.t23 GNDA 0.115045f
C3186 bgr_0.V_TOP.t29 GNDA 0.115045f
C3187 bgr_0.V_TOP.t43 GNDA 0.150392f
C3188 bgr_0.V_TOP.n0 GNDA 0.084081f
C3189 bgr_0.V_TOP.n1 GNDA 0.061357f
C3190 bgr_0.V_TOP.n2 GNDA 0.061357f
C3191 bgr_0.V_TOP.n3 GNDA 0.061357f
C3192 bgr_0.V_TOP.n4 GNDA 0.061357f
C3193 bgr_0.V_TOP.n5 GNDA 0.057217f
C3194 bgr_0.V_TOP.t2 GNDA 0.147947f
C3195 bgr_0.V_TOP.t6 GNDA 0.155772f
C3196 bgr_0.V_TOP.t11 GNDA 0.010957f
C3197 bgr_0.V_TOP.t12 GNDA 0.010957f
C3198 bgr_0.V_TOP.n6 GNDA 0.027281f
C3199 bgr_0.V_TOP.n7 GNDA 0.726844f
C3200 bgr_0.V_TOP.t1 GNDA 0.010957f
C3201 bgr_0.V_TOP.t13 GNDA 0.010957f
C3202 bgr_0.V_TOP.n8 GNDA 0.026425f
C3203 bgr_0.V_TOP.t4 GNDA 0.010957f
C3204 bgr_0.V_TOP.t8 GNDA 0.010957f
C3205 bgr_0.V_TOP.n9 GNDA 0.027465f
C3206 bgr_0.V_TOP.t5 GNDA 0.010957f
C3207 bgr_0.V_TOP.t0 GNDA 0.010957f
C3208 bgr_0.V_TOP.n10 GNDA 0.027281f
C3209 bgr_0.V_TOP.n11 GNDA 0.252824f
C3210 bgr_0.V_TOP.n12 GNDA 0.153577f
C3211 bgr_0.V_TOP.n13 GNDA 0.087653f
C3212 bgr_0.V_TOP.t9 GNDA 0.010957f
C3213 bgr_0.V_TOP.t10 GNDA 0.010957f
C3214 bgr_0.V_TOP.n14 GNDA 0.027281f
C3215 bgr_0.V_TOP.n15 GNDA 0.151313f
C3216 bgr_0.V_TOP.t7 GNDA 0.010957f
C3217 bgr_0.V_TOP.t3 GNDA 0.010957f
C3218 bgr_0.V_TOP.n16 GNDA 0.027281f
C3219 bgr_0.V_TOP.n17 GNDA 0.149874f
C3220 bgr_0.V_TOP.n18 GNDA 0.329448f
C3221 bgr_0.V_TOP.n19 GNDA 0.023183f
C3222 bgr_0.V_TOP.n20 GNDA 0.057217f
C3223 bgr_0.V_TOP.n21 GNDA 0.061357f
C3224 bgr_0.V_TOP.n22 GNDA 0.061357f
C3225 bgr_0.V_TOP.n23 GNDA 0.061357f
C3226 bgr_0.V_TOP.n24 GNDA 0.061357f
C3227 bgr_0.V_TOP.n25 GNDA 0.061357f
C3228 bgr_0.V_TOP.n26 GNDA 0.061357f
C3229 bgr_0.V_TOP.n27 GNDA 0.057217f
C3230 bgr_0.V_TOP.t32 GNDA 0.132572f
C3231 bgr_0.V_TOP.t49 GNDA 0.445732f
C3232 bgr_0.V_TOP.t39 GNDA 0.438267f
C3233 bgr_0.V_TOP.n28 GNDA 0.293844f
C3234 bgr_0.V_TOP.t28 GNDA 0.438267f
C3235 bgr_0.V_TOP.t25 GNDA 0.445732f
C3236 bgr_0.V_TOP.t33 GNDA 0.438267f
C3237 bgr_0.V_TOP.n29 GNDA 0.293844f
C3238 bgr_0.V_TOP.n30 GNDA 0.273917f
C3239 bgr_0.V_TOP.t21 GNDA 0.445732f
C3240 bgr_0.V_TOP.t15 GNDA 0.438267f
C3241 bgr_0.V_TOP.n31 GNDA 0.293844f
C3242 bgr_0.V_TOP.t40 GNDA 0.438267f
C3243 bgr_0.V_TOP.t34 GNDA 0.445732f
C3244 bgr_0.V_TOP.t45 GNDA 0.438267f
C3245 bgr_0.V_TOP.n32 GNDA 0.293844f
C3246 bgr_0.V_TOP.n33 GNDA 0.356092f
C3247 bgr_0.V_TOP.t30 GNDA 0.445732f
C3248 bgr_0.V_TOP.t22 GNDA 0.438267f
C3249 bgr_0.V_TOP.n34 GNDA 0.293844f
C3250 bgr_0.V_TOP.t16 GNDA 0.438267f
C3251 bgr_0.V_TOP.t46 GNDA 0.445732f
C3252 bgr_0.V_TOP.t19 GNDA 0.438267f
C3253 bgr_0.V_TOP.n35 GNDA 0.293844f
C3254 bgr_0.V_TOP.n36 GNDA 0.356092f
C3255 bgr_0.V_TOP.t24 GNDA 0.445732f
C3256 bgr_0.V_TOP.t17 GNDA 0.438267f
C3257 bgr_0.V_TOP.n37 GNDA 0.293844f
C3258 bgr_0.V_TOP.t42 GNDA 0.438267f
C3259 bgr_0.V_TOP.n38 GNDA 0.273917f
C3260 bgr_0.V_TOP.t47 GNDA 0.438267f
C3261 bgr_0.V_TOP.n39 GNDA 0.191742f
C3262 bgr_0.V_TOP.t36 GNDA 0.438267f
C3263 bgr_0.V_TOP.n40 GNDA 0.893239f
.ends

