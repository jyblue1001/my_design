* PEX produced on Sun Jul  6 07:26:22 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t311 bgr_0.V_TOP.t14 bgr_0.Vin-.t3 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 bgr_0.V_TOP.t15 VDDA.t309 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 a_14710_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t165 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X4 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t310 GNDA.t312 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X5 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t40 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X7 GNDA.t230 GNDA.t309 bgr_0.Vbe2.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_0.Y.t25 GNDA.t162 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X9 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.t1 GNDA.t325 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X12 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 two_stage_opamp_dummy_magic_0.V_err_gate.t11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X14 bgr_0.V_TOP.t16 VDDA.t308 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VDDA.t125 bgr_0.V_mir2.t15 bgr_0.V_mir2.t16 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X16 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 two_stage_opamp_dummy_magic_0.Y.t4 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.VD4.t21 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X19 VDDA.t139 two_stage_opamp_dummy_magic_0.X.t25 VOUT+.t11 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X20 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t137 two_stage_opamp_dummy_magic_0.X.t26 VOUT+.t10 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X23 VDDA.t116 bgr_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X24 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 VOUT+.t18 GNDA.t306 GNDA.t308 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X26 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD1.t10 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X27 bgr_0.V_TOP.t17 VDDA.t307 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VDDA.t80 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X29 a_5160_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t180 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X30 VDDA.t156 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X31 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t126 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X33 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VDDA.t44 two_stage_opamp_dummy_magic_0.X.t27 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X36 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VOUT-.t6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X42 VDDA.t198 two_stage_opamp_dummy_magic_0.Y.t26 VOUT-.t7 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X43 VDDA.t426 VDDA.t424 two_stage_opamp_dummy_magic_0.V_err_gate.t13 VDDA.t425 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X44 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 bgr_0.V_mir2.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 bgr_0.V_p_2.t8 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X46 bgr_0.Vin-.t4 bgr_0.V_TOP.t18 VDDA.t306 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X47 GNDA.t28 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 GNDA.t168 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X49 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t252 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X50 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 two_stage_opamp_dummy_magic_0.V_err_p.t4 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 VDDA.t447 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 two_stage_opamp_dummy_magic_0.Y.t19 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X54 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VDDA.t194 two_stage_opamp_dummy_magic_0.Y.t27 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X56 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 two_stage_opamp_dummy_magic_0.X.t28 GNDA.t19 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X57 bgr_0.1st_Vout_1.t2 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X58 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VDDA.t423 VDDA.t421 bgr_0.V_TOP.t0 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X61 two_stage_opamp_dummy_magic_0.VD1.t21 VIN-.t0 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X62 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X63 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 GNDA.t170 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X65 GNDA.t305 GNDA.t303 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X66 VDDA.t160 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t6 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X67 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X70 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 GNDA.t164 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X74 two_stage_opamp_dummy_magic_0.VD1.t19 VIN-.t1 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA.t322 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X75 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 bgr_0.NFET_GATE_10uA.t0 bgr_0.PFET_GATE_10uA.t11 VDDA.t74 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X77 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 VDDA.t49 bgr_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X79 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VDDA.t420 VDDA.t418 bgr_0.NFET_GATE_10uA.t3 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X81 VDDA.t12 two_stage_opamp_dummy_magic_0.X.t29 VOUT+.t9 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X82 GNDA.t42 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X83 VDDA.t67 bgr_0.1st_Vout_1.t14 bgr_0.V_TOP.t3 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X84 GNDA.t302 GNDA.t300 two_stage_opamp_dummy_magic_0.VD1.t18 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X85 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 two_stage_opamp_dummy_magic_0.VD3.t30 VDDA.t415 VDDA.t417 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X87 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT+.t14 a_14240_2076.t0 GNDA.t150 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X89 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VDDA.t39 bgr_0.V_mir2.t13 bgr_0.V_mir2.t14 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X92 two_stage_opamp_dummy_magic_0.Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X93 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.VD1.t9 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X94 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.X.t19 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X95 GNDA.t176 bgr_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X96 VDDA.t63 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X97 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 two_stage_opamp_dummy_magic_0.Vb3.t5 bgr_0.NFET_GATE_10uA.t9 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X99 GNDA.t299 GNDA.t297 two_stage_opamp_dummy_magic_0.VD1.t17 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X100 VDDA.t90 two_stage_opamp_dummy_magic_0.X.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X101 VDDA.t65 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t2 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X102 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 bgr_0.V_TOP.t13 bgr_0.cap_res1.t20 GNDA.t148 sky130_fd_pr__res_high_po_0p35 l=2.05
X104 a_11220_17410.t0 GNDA.t22 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=6
X105 VDDA.t23 two_stage_opamp_dummy_magic_0.Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=0.71 ps=3.95 w=3.55 l=0.2
X106 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t466 VDDA.t465 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X107 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 two_stage_opamp_dummy_magic_0.V_source.t27 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA.t187 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X109 two_stage_opamp_dummy_magic_0.Vb1.t1 bgr_0.PFET_GATE_10uA.t13 VDDA.t107 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X110 VDDA.t195 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X111 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VDDA.t255 two_stage_opamp_dummy_magic_0.Y.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t200 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X113 bgr_0.PFET_GATE_10uA.t2 bgr_0.1st_Vout_2.t13 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X114 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 two_stage_opamp_dummy_magic_0.V_source.t8 two_stage_opamp_dummy_magic_0.Vb1.t2 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X116 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.Vb3.t9 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VDDA.t53 bgr_0.V_mir1.t10 bgr_0.V_mir1.t11 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X123 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 a_14590_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t344 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X125 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X126 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 GNDA.t327 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 VOUT-.t18 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X128 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VDDA.t47 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t0 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X131 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X132 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_0.Y.t30 GNDA.t201 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X133 bgr_0.V_TOP.t19 VDDA.t304 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 GNDA.t36 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X135 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.VD4.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X136 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.X.t20 GNDA.t153 sky130_fd_pr__res_high_po_1p41 l=1.41
X139 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t294 GNDA.t296 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X141 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 two_stage_opamp_dummy_magic_0.V_source.t13 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VDDA.t207 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t10 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X146 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 two_stage_opamp_dummy_magic_0.X.t22 GNDA.t291 GNDA.t293 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X149 GNDA.t290 GNDA.t287 GNDA.t289 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X150 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 GNDA.t93 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X152 a_13730_17020.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X153 GNDA.t202 two_stage_opamp_dummy_magic_0.Y.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X154 two_stage_opamp_dummy_magic_0.V_source.t37 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t332 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X155 VDDA.t460 two_stage_opamp_dummy_magic_0.X.t31 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA.t347 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X156 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 bgr_0.V_CUR_REF_REG.t2 VDDA.t412 VDDA.t414 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X158 a_11220_17410.t1 a_12828_17530.t0 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=6
X159 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VDDA.t259 two_stage_opamp_dummy_magic_0.Y.t32 VOUT-.t13 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X161 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t14 VDDA.t95 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X163 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VDDA.t92 bgr_0.PFET_GATE_10uA.t15 bgr_0.V_CUR_REF_REG.t0 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X166 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.Vb3.t11 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X167 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 bgr_0.PFET_GATE_10uA.t4 bgr_0.cap_res2.t20 GNDA.t148 sky130_fd_pr__res_high_po_0p35 l=2.05
X169 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X170 bgr_0.V_p_1.t9 bgr_0.Vin-.t8 bgr_0.V_mir1.t14 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X171 VDDA.t57 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X172 two_stage_opamp_dummy_magic_0.V_source.t0 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X173 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VDDA.t101 bgr_0.1st_Vout_1.t19 bgr_0.V_TOP.t5 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X179 VDDA.t303 bgr_0.V_TOP.t20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X180 VDDA.t246 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X181 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 bgr_0.V_p_2.t2 bgr_0.V_CUR_REF_REG.t3 bgr_0.1st_Vout_2.t2 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X184 two_stage_opamp_dummy_magic_0.Y.t6 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X185 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 VOUT-.t12 two_stage_opamp_dummy_magic_0.Y.t34 VDDA.t248 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X188 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 bgr_0.V_p_1.t8 bgr_0.Vin-.t9 bgr_0.V_mir1.t12 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X190 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_0.V_TOP.t9 VDDA.t409 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X192 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 bgr_0.Vin-.t7 bgr_0.START_UP.t6 bgr_0.V_TOP.t12 VDDA.t430 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X194 VDDA.t408 VDDA.t406 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X195 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t19 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X199 bgr_0.V_TOP.t21 VDDA.t293 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_2076.t1 GNDA.t179 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X203 VDDA.t21 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD3.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X204 GNDA.t96 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X205 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X207 a_13730_17020.t1 GNDA.t334 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X208 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 bgr_0.V_TOP.t22 VDDA.t292 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.VD4.t35 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X211 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t387 VDDA.t389 VDDA.t388 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X212 a_11220_17290.t1 a_12828_17650.t1 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=6
X213 VDDA.t173 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD4.t24 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X214 two_stage_opamp_dummy_magic_0.X.t16 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.VD1.t8 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X215 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 GNDA.t14 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X220 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t4 bgr_0.1st_Vout_2.t4 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X221 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 bgr_0.PFET_GATE_10uA.t16 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X222 VDDA.t185 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X223 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 VDDA.t114 bgr_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X225 two_stage_opamp_dummy_magic_0.V_source.t38 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t335 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X226 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VDDA.t405 VDDA.t403 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=0 ps=0 w=3.55 l=0.2
X228 GNDA.t191 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X229 VDDA.t448 two_stage_opamp_dummy_magic_0.X.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X230 a_11220_17290.t0 GNDA.t321 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=6
X231 two_stage_opamp_dummy_magic_0.V_source.t22 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X232 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t284 GNDA.t286 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X233 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t10 VDDA.t253 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X236 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 bgr_0.START_UP.t5 bgr_0.V_TOP.t23 VDDA.t301 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X238 bgr_0.1st_Vout_2.t9 bgr_0.V_mir2.t18 VDDA.t209 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X239 bgr_0.V_TOP.t24 VDDA.t299 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 two_stage_opamp_dummy_magic_0.V_source.t39 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA.t341 GNDA.t340 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X243 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VDDA.t227 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.VD3.t26 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X246 VDDA.t162 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t7 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X247 VOUT+.t8 two_stage_opamp_dummy_magic_0.X.t35 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X248 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 bgr_0.V_p_2.t3 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t3 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X252 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t400 VDDA.t402 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X253 GNDA.t283 GNDA.t281 two_stage_opamp_dummy_magic_0.X.t21 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X254 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 VDDA.t33 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD4.t2 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X257 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 two_stage_opamp_dummy_magic_0.Y.t21 GNDA.t278 GNDA.t280 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X259 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 bgr_0.V_TOP.t25 VDDA.t298 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 GNDA.t234 GNDA.t277 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X263 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VDDA.t2 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.VD3.t0 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X267 VOUT-.t11 two_stage_opamp_dummy_magic_0.Y.t36 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X268 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X269 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 GNDA.t133 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X272 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 VDDA.t29 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t11 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X274 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 VDDA.t211 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X276 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X278 bgr_0.V_mir2.t12 bgr_0.V_mir2.t11 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X279 VDDA.t297 bgr_0.V_TOP.t26 bgr_0.Vin-.t5 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X280 GNDA.t336 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X281 VDDA.t399 VDDA.t397 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 bgr_0.PFET_GATE_10uA.t18 VDDA.t450 VDDA.t449 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X283 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X284 two_stage_opamp_dummy_magic_0.V_source.t21 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X285 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 bgr_0.Vin-.t1 a_12828_17650.t0 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=6
X289 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 GNDA.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X293 GNDA.t236 GNDA.t276 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X294 VDDA.t176 GNDA.t273 GNDA.t275 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.15
X295 two_stage_opamp_dummy_magic_0.V_source.t20 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X296 two_stage_opamp_dummy_magic_0.Y.t11 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X297 VDDA.t233 two_stage_opamp_dummy_magic_0.Vb3.t17 two_stage_opamp_dummy_magic_0.VD3.t28 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X298 GNDA.t189 two_stage_opamp_dummy_magic_0.Y.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X299 two_stage_opamp_dummy_magic_0.VD4.t30 VDDA.t394 VDDA.t396 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X300 GNDA.t190 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X301 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t4 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X304 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 GNDA.t195 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X307 bgr_0.PFET_GATE_10uA.t3 bgr_0.1st_Vout_2.t19 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X308 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t3 VDDA.t452 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X309 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t270 GNDA.t272 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X312 GNDA.t269 GNDA.t267 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X313 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 bgr_0.NFET_GATE_10uA.t12 GNDA.t83 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X314 bgr_0.START_UP.t1 bgr_0.START_UP.t0 bgr_0.START_UP_NFET1.t0 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X315 two_stage_opamp_dummy_magic_0.V_source.t5 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X316 VDDA.t393 VDDA.t390 VDDA.t392 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.24 pd=2 as=0 ps=0 w=0.6 l=0.2
X317 VOUT+.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA.t53 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X318 VOUT+.t7 two_stage_opamp_dummy_magic_0.X.t37 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X319 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 GNDA.t137 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X328 bgr_0.V_p_1.t3 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t1 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X329 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t213 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X330 two_stage_opamp_dummy_magic_0.Vb2.t5 bgr_0.NFET_GATE_10uA.t14 GNDA.t129 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X331 two_stage_opamp_dummy_magic_0.VD1.t7 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.X.t15 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X332 two_stage_opamp_dummy_magic_0.V_source.t9 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA.t62 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X333 two_stage_opamp_dummy_magic_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t15 GNDA.t115 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X334 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X336 two_stage_opamp_dummy_magic_0.VD3.t23 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.VD3.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X337 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 VOUT-.t9 two_stage_opamp_dummy_magic_0.Y.t39 VDDA.t238 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X339 VOUT-.t10 two_stage_opamp_dummy_magic_0.Y.t40 VDDA.t240 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X340 bgr_0.Vin+.t5 bgr_0.V_TOP.t27 VDDA.t295 VDDA.t294 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X341 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VOUT+.t13 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t135 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X344 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VDDA.t220 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X346 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.Vb3.t18 VDDA.t440 VDDA.t439 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X347 VDDA.t455 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 VDDA.t454 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X348 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t2 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X349 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 bgr_0.PFET_GATE_10uA.t20 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X351 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_p.t18 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X352 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 GNDA.t177 two_stage_opamp_dummy_magic_0.X.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X354 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 GNDA.t38 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X356 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 bgr_0.V_TOP.t28 VDDA.t291 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 bgr_0.Vin+.t1 a_12828_17530.t1 GNDA.t21 sky130_fd_pr__res_xhigh_po_0p35 l=6
X360 two_stage_opamp_dummy_magic_0.V_source.t25 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X361 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t118 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X363 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t264 GNDA.t266 GNDA.t265 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X366 GNDA.t263 GNDA.t261 two_stage_opamp_dummy_magic_0.Y.t20 GNDA.t262 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X367 two_stage_opamp_dummy_magic_0.Vb3.t4 bgr_0.NFET_GATE_10uA.t16 GNDA.t174 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X368 GNDA.t60 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_p_mir.t2 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X369 GNDA.t197 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA.t196 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X370 VDDA.t386 VDDA.t384 two_stage_opamp_dummy_magic_0.Vb2.t8 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=0.24 pd=2 as=0.12 ps=1 w=0.6 l=0.2
X371 two_stage_opamp_dummy_magic_0.V_source.t31 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA.t314 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X372 bgr_0.V_mir1.t7 bgr_0.V_mir1.t6 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X373 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t68 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X374 GNDA.t188 two_stage_opamp_dummy_magic_0.Y.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X375 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t9 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X378 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 bgr_0.V_p_2.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 bgr_0.V_mir2.t1 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X380 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 two_stage_opamp_dummy_magic_0.V_source.t10 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X382 VDDA.t446 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.Vb1.t0 VDDA.t445 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X383 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VOUT+.t6 two_stage_opamp_dummy_magic_0.X.t39 VDDA.t167 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X386 VDDA.t444 GNDA.t258 GNDA.t260 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=1.6 ps=8.8 w=4 l=0.15
X387 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.Vb3.t20 VDDA.t457 VDDA.t456 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X389 bgr_0.V_p_1.t2 bgr_0.Vin+.t8 bgr_0.1st_Vout_1.t10 GNDA.t343 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X390 two_stage_opamp_dummy_magic_0.VD1.t6 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.X.t1 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X391 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 VDDA.t290 bgr_0.V_TOP.t29 bgr_0.START_UP.t4 VDDA.t289 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X393 two_stage_opamp_dummy_magic_0.V_err_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X394 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Y.t24 two_stage_opamp_dummy_magic_0.VD4.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X395 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 GNDA.t257 GNDA.t255 VDDA.t110 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.15
X398 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X399 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 bgr_0.V_p_2.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 bgr_0.V_mir2.t3 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X402 VOUT-.t8 two_stage_opamp_dummy_magic_0.Y.t42 VDDA.t236 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X403 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VDDA.t87 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X407 two_stage_opamp_dummy_magic_0.err_amp_out.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X408 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t43 VDDA.t84 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X409 GNDA.t75 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X410 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 GNDA.t319 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 VDDA.t435 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X413 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 two_stage_opamp_dummy_magic_0.V_source.t19 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t12 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X415 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t20 VDDA.t146 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X416 VDDA.t224 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t8 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X417 GNDA.t51 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 VOUT-.t3 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X418 GNDA.t216 VDDA.t469 bgr_0.V_TOP.t7 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X419 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.Vb3.t21 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X420 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X422 two_stage_opamp_dummy_magic_0.VD2.t1 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X423 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 bgr_0.1st_Vout_2.t8 bgr_0.V_mir2.t19 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X426 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 GNDA.t70 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 VOUT+.t1 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X431 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_0.err_amp_out.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA.t64 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X433 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VDDA.t17 bgr_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X435 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 two_stage_opamp_dummy_magic_0.Vb2.t1 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.12 pd=1 as=0.12 ps=1 w=0.6 l=0.2
X437 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t432 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X438 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 bgr_0.V_TOP.t30 VDDA.t288 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X442 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 bgr_0.START_UP.t3 bgr_0.V_TOP.t31 VDDA.t287 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X444 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 GNDA.t254 GNDA.t252 VOUT-.t17 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X448 VOUT+.t5 two_stage_opamp_dummy_magic_0.X.t42 VDDA.t442 VDDA.t441 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X449 two_stage_opamp_dummy_magic_0.err_amp_out.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 GNDA.t66 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X450 VOUT+.t4 two_stage_opamp_dummy_magic_0.X.t43 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X451 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 bgr_0.V_mir2.t10 bgr_0.V_mir2.t9 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X453 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 two_stage_opamp_dummy_magic_0.VD1.t5 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.X.t24 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X455 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.VD3.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X457 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t464 VDDA.t463 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X459 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 bgr_0.V_TOP.t6 bgr_0.1st_Vout_1.t27 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X461 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 two_stage_opamp_dummy_magic_0.X.t44 VDDA.t177 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X463 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 GNDA.t230 GNDA.t251 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X467 bgr_0.V_mir2.t8 bgr_0.V_mir2.t7 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X468 VDDA.t285 bgr_0.V_TOP.t32 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X469 two_stage_opamp_dummy_magic_0.V_err_gate.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X470 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VDDA.t383 VDDA.t381 bgr_0.V_TOP.t8 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X473 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VDDA.t468 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X475 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 bgr_0.V_TOP.t33 VDDA.t283 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 GNDA.t250 GNDA.t248 two_stage_opamp_dummy_magic_0.V_source.t30 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X478 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 VDDA.t378 VDDA.t380 VDDA.t379 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X479 VDDA.t231 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.VD4.t28 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X480 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_0.Y.t44 VDDA.t85 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X481 GNDA.t247 GNDA.t245 VDDA.t103 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=1.6 pd=8.8 as=0.8 ps=4.4 w=4 l=0.15
X482 GNDA.t215 VDDA.t375 VDDA.t377 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X483 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5750_2076.t1 GNDA.t149 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X484 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 GNDA.t234 GNDA.t244 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X488 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 two_stage_opamp_dummy_magic_0.V_source.t29 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X490 bgr_0.V_TOP.t34 VDDA.t282 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t26 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X494 a_13790_17550.t0 bgr_0.V_CUR_REF_REG.t1 GNDA.t88 sky130_fd_pr__res_xhigh_po_0p35 l=6
X495 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VDDA.t72 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X497 VDDA.t281 bgr_0.V_TOP.t35 bgr_0.Vin+.t4 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X498 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 VDDA.t372 VDDA.t374 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X499 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X502 GNDA.t214 VDDA.t470 bgr_0.V_p_2.t10 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X503 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 bgr_0.V_p_1.t7 bgr_0.Vin-.t10 bgr_0.V_mir1.t15 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X505 VDDA.t19 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD4.t1 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X506 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X507 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 bgr_0.V_TOP.t1 bgr_0.1st_Vout_1.t30 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X510 VOUT+.t16 VDDA.t369 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X511 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 bgr_0.V_TOP.t36 VDDA.t277 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 VOUT-.t16 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X515 GNDA.t236 GNDA.t240 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X516 two_stage_opamp_dummy_magic_0.VD1.t16 VIN-.t6 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X517 bgr_0.1st_Vout_1.t4 bgr_0.V_mir1.t21 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X518 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 two_stage_opamp_dummy_magic_0.VD1.t4 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X525 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 two_stage_opamp_dummy_magic_0.V_p_mir.t1 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t26 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X527 bgr_0.Vin+.t3 bgr_0.V_TOP.t37 VDDA.t279 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X528 bgr_0.V_mir2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t5 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X529 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 bgr_0.PFET_GATE_10uA.t8 VDDA.t471 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X531 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_0.X.t45 VDDA.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X532 two_stage_opamp_dummy_magic_0.VD1.t11 VIN-.t7 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X533 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 GNDA.t239 GNDA.t237 bgr_0.NFET_GATE_10uA.t4 GNDA.t238 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X539 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 two_stage_opamp_dummy_magic_0.V_err_gate.t5 bgr_0.NFET_GATE_10uA.t18 GNDA.t142 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X541 bgr_0.1st_Vout_1.t0 bgr_0.Vin+.t9 bgr_0.V_p_1.t1 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X542 VOUT-.t1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X543 GNDA.t145 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X544 GNDA.t184 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_0.V_source.t28 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X545 bgr_0.V_TOP.t4 bgr_0.1st_Vout_1.t31 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X546 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 two_stage_opamp_dummy_magic_0.Y.t45 VDDA.t131 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X549 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 bgr_0.PFET_GATE_10uA.t24 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X550 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 bgr_0.Vin-.t2 bgr_0.V_TOP.t38 VDDA.t276 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X553 VDDA.t205 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X554 VDDA.t368 VDDA.t366 two_stage_opamp_dummy_magic_0.VD3.t29 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X555 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X557 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 a_13790_17550.t1 GNDA.t139 GNDA.t88 sky130_fd_pr__res_xhigh_po_0p35 l=6
X559 two_stage_opamp_dummy_magic_0.VD2.t5 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.Y.t9 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X560 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 bgr_0.V_TOP.t10 VDDA.t363 VDDA.t365 VDDA.t364 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X563 VDDA.t362 VDDA.t360 two_stage_opamp_dummy_magic_0.VD4.t29 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X564 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 GNDA.t211 VDDA.t357 VDDA.t359 VDDA.t358 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X568 bgr_0.V_TOP.t39 VDDA.t274 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 bgr_0.NFET_GATE_10uA.t19 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X572 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 bgr_0.NFET_GATE_10uA.t20 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X573 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 VDDA.t356 VDDA.t354 two_stage_opamp_dummy_magic_0.err_amp_out.t10 VDDA.t355 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X575 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VDDA.t37 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t7 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X578 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 bgr_0.V_TOP.t40 VDDA.t273 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 VDDA.t272 bgr_0.V_TOP.t41 bgr_0.Vin+.t2 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X581 VDDA.t353 VDDA.t351 GNDA.t210 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X582 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X584 bgr_0.V_mir1.t3 bgr_0.V_mir1.t2 VDDA.t438 VDDA.t437 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X585 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 two_stage_opamp_dummy_magic_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t21 GNDA.t346 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X587 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.VD4.t8 two_stage_opamp_dummy_magic_0.VD4.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X588 GNDA.t234 GNDA.t233 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X589 bgr_0.V_mir2.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 bgr_0.V_p_2.t4 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X590 bgr_0.PFET_GATE_10uA.t7 VDDA.t348 VDDA.t350 VDDA.t349 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X591 two_stage_opamp_dummy_magic_0.VD1.t3 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.X.t14 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X592 two_stage_opamp_dummy_magic_0.V_source.t2 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X593 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_0.X.t46 VDDA.t13 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X594 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_0.X.t47 VDDA.t178 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X595 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 two_stage_opamp_dummy_magic_0.Y.t46 GNDA.t122 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X596 two_stage_opamp_dummy_magic_0.VD2.t17 VIN+.t7 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X597 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 VOUT-.t15 VDDA.t345 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X599 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 two_stage_opamp_dummy_magic_0.V_err_gate.t1 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X601 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VDDA.t344 VDDA.t342 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X603 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X604 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X605 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 bgr_0.V_TOP.t42 VDDA.t270 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 GNDA.t47 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_0.V_source.t7 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X608 VOUT-.t4 a_5750_2076.t0 GNDA.t72 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X609 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 bgr_0.PFET_GATE_10uA.t26 VDDA.t182 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X610 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 VDDA.t341 VDDA.t339 VOUT+.t15 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X613 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 bgr_0.1st_Vout_2.t6 bgr_0.V_mir2.t21 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X615 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_0.Y.t47 VDDA.t40 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X616 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X617 GNDA.t236 GNDA.t235 bgr_0.Vin-.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X618 two_stage_opamp_dummy_magic_0.VD2.t0 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X619 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 GNDA.t85 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X621 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 VDDA.t42 two_stage_opamp_dummy_magic_0.Y.t48 VOUT-.t2 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X624 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 bgr_0.V_TOP.t43 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X627 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 VDDA.t336 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X629 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.X.t10 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X630 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X631 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t222 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X632 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 VDDA.t61 bgr_0.1st_Vout_2.t32 bgr_0.PFET_GATE_10uA.t1 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X635 VDDA.t335 VDDA.t333 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X636 two_stage_opamp_dummy_magic_0.V_err_p.t1 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X637 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t330 VDDA.t332 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X639 a_5160_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t333 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X640 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_0.X.t48 GNDA.t178 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X642 two_stage_opamp_dummy_magic_0.VD2.t16 VIN+.t8 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA.t316 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X643 GNDA.t232 GNDA.t231 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X644 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X649 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 bgr_0.V_mir1.t13 bgr_0.Vin-.t11 bgr_0.V_p_1.t6 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X651 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 two_stage_opamp_dummy_magic_0.V_source.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X654 two_stage_opamp_dummy_magic_0.VD2.t15 VIN+.t9 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X655 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t163 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X656 two_stage_opamp_dummy_magic_0.VD3.t24 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X657 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 two_stage_opamp_dummy_magic_0.Y.t49 GNDA.t9 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X659 VDDA.t329 VDDA.t327 GNDA.t209 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X660 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 two_stage_opamp_dummy_magic_0.V_err_gate.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X662 a_14710_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA.t152 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X663 GNDA.t120 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X664 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X665 VDDA.t169 two_stage_opamp_dummy_magic_0.X.t50 VOUT+.t3 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X666 GNDA.t49 bgr_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X667 VDDA.t267 bgr_0.V_TOP.t44 bgr_0.START_UP.t2 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X668 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.Y.t12 two_stage_opamp_dummy_magic_0.VD4.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X670 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 VDDA.t27 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X673 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t338 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X674 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 GNDA.t342 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X676 GNDA.t230 GNDA.t229 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X677 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.Y.t16 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X679 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 VDDA.t5 two_stage_opamp_dummy_magic_0.Y.t50 VOUT-.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X681 a_5280_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA.t124 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X682 VDDA.t326 VDDA.t324 VOUT-.t14 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X683 VDDA.t459 bgr_0.V_mir2.t5 bgr_0.V_mir2.t6 VDDA.t458 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X684 VDDA.t203 bgr_0.PFET_GATE_10uA.t27 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X685 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 bgr_0.PFET_GATE_10uA.t28 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X688 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 bgr_0.V_TOP.t45 VDDA.t265 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 two_stage_opamp_dummy_magic_0.V_err_p.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t152 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X691 two_stage_opamp_dummy_magic_0.V_source.t6 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X692 bgr_0.1st_Vout_1.t8 bgr_0.V_mir1.t22 VDDA.t217 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X693 two_stage_opamp_dummy_magic_0.V_err_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X694 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X696 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_0.X.t51 GNDA.t76 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X698 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 bgr_0.1st_Vout_2.t0 bgr_0.V_CUR_REF_REG.t6 bgr_0.V_p_2.t0 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X700 bgr_0.V_TOP.t46 VDDA.t264 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.Y.t18 two_stage_opamp_dummy_magic_0.VD4.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X702 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X703 two_stage_opamp_dummy_magic_0.V_p_mir.t3 VIN-.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X704 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t9 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X705 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 bgr_0.V_p_1.t10 VDDA.t472 GNDA.t208 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X710 GNDA.t131 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 VOUT+.t12 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X711 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 bgr_0.V_mir1.t16 bgr_0.Vin-.t12 bgr_0.V_p_1.t5 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X713 VDDA.t323 VDDA.t321 bgr_0.PFET_GATE_10uA.t6 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X714 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 two_stage_opamp_dummy_magic_0.V_source.t1 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA.t6 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X717 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 two_stage_opamp_dummy_magic_0.VD1.t15 VIN-.t10 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X719 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X720 GNDA.t228 GNDA.t226 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA.t227 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X721 bgr_0.V_TOP.t47 VDDA.t263 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 VDDA.t7 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD4.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X723 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 two_stage_opamp_dummy_magic_0.Y.t51 GNDA.t198 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X724 VDDA.t154 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X725 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 two_stage_opamp_dummy_magic_0.V_err_gate.t12 VDDA.t318 VDDA.t320 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X727 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 bgr_0.V_TOP.t48 VDDA.t262 VDDA.t261 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X729 bgr_0.V_TOP.t11 bgr_0.START_UP.t7 bgr_0.Vin-.t6 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X730 two_stage_opamp_dummy_magic_0.V_err_gate.t0 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X731 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 bgr_0.1st_Vout_2.t1 bgr_0.V_CUR_REF_REG.t7 bgr_0.V_p_2.t1 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X733 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 VDDA.t434 bgr_0.1st_Vout_2.t36 bgr_0.PFET_GATE_10uA.t9 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X735 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X736 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.Y.t10 GNDA.t102 sky130_fd_pr__res_high_po_1p41 l=1.41
X737 GNDA.t331 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 two_stage_opamp_dummy_magic_0.V_source.t36 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X738 a_14590_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t138 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X739 GNDA.t225 GNDA.t223 VOUT+.t17 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X740 VDDA.t15 two_stage_opamp_dummy_magic_0.X.t52 VOUT+.t2 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X741 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 two_stage_opamp_dummy_magic_0.Y.t52 VDDA.t250 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X742 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 VDDA.t428 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t5 VDDA.t427 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X750 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t1 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X751 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.VD4.t33 two_stage_opamp_dummy_magic_0.VD4.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X752 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VDDA.t317 VDDA.t315 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X755 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 bgr_0.PFET_GATE_10uA.t29 VDDA.t462 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X757 two_stage_opamp_dummy_magic_0.VD2.t21 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.Y.t23 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X758 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X759 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X760 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 VDDA.t78 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t5 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X762 VDDA.t129 two_stage_opamp_dummy_magic_0.Y.t53 VOUT-.t5 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X763 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 a_5280_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t143 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X767 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X768 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 two_stage_opamp_dummy_magic_0.V_err_p.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t4 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X770 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t312 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.71 pd=3.95 as=1.42 ps=7.9 w=3.55 l=0.2
X771 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 VDDA.t130 two_stage_opamp_dummy_magic_0.Y.t54 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.4 as=0.8 ps=4.4 w=4 l=0.15
X773 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_0.X.t53 GNDA.t320 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X774 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t329 VDDA.t443 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X778 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 bgr_0.V_TOP.t49 VDDA.t260 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X780 bgr_0.1st_Vout_1.t9 bgr_0.Vin+.t10 bgr_0.V_p_1.t0 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X781 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA.t220 GNDA.t222 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X782 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA.t217 GNDA.t219 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X783 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 two_stage_opamp_dummy_magic_0.VD2.t18 VIN+.t10 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA.t318 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X785 bgr_0.Vin+.t0 bgr_0.Vbe2.t0 GNDA.t101 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X786 VDDA.t229 two_stage_opamp_dummy_magic_0.Vb3.t28 two_stage_opamp_dummy_magic_0.VD3.t27 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X787 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X788 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.V_TOP.n0 bgr_0.V_TOP.t43 369.534
R1 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 339.961
R2 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 339.272
R3 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R4 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R5 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R6 bgr_0.V_TOP.n12 bgr_0.V_TOP.n8 334.772
R7 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R8 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R9 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R10 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R11 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R12 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R13 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R14 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R15 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R16 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R17 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R18 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R19 bgr_0.V_TOP bgr_0.V_TOP.t32 214.222
R20 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R21 bgr_0.V_TOP.n7 bgr_0.V_TOP.t13 176.114
R22 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R23 bgr_0.V_TOP.n27 bgr_0.V_TOP.t31 144.601
R24 bgr_0.V_TOP.n26 bgr_0.V_TOP.t44 144.601
R25 bgr_0.V_TOP.n25 bgr_0.V_TOP.t18 144.601
R26 bgr_0.V_TOP.n24 bgr_0.V_TOP.t26 144.601
R27 bgr_0.V_TOP.n23 bgr_0.V_TOP.t37 144.601
R28 bgr_0.V_TOP.n22 bgr_0.V_TOP.t35 144.601
R29 bgr_0.V_TOP.n21 bgr_0.V_TOP.t48 144.601
R30 bgr_0.V_TOP.n20 bgr_0.V_TOP.t20 144.601
R31 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 144.601
R32 bgr_0.V_TOP.n1 bgr_0.V_TOP.t23 144.601
R33 bgr_0.V_TOP.n2 bgr_0.V_TOP.t14 144.601
R34 bgr_0.V_TOP.n3 bgr_0.V_TOP.t38 144.601
R35 bgr_0.V_TOP.n4 bgr_0.V_TOP.t41 144.601
R36 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R37 bgr_0.V_TOP.n18 bgr_0.V_TOP.t7 95.4466
R38 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R39 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R40 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R41 bgr_0.V_TOP.n6 bgr_0.V_TOP.t0 39.4005
R42 bgr_0.V_TOP.n6 bgr_0.V_TOP.t1 39.4005
R43 bgr_0.V_TOP.n8 bgr_0.V_TOP.t3 39.4005
R44 bgr_0.V_TOP.n8 bgr_0.V_TOP.t4 39.4005
R45 bgr_0.V_TOP.n10 bgr_0.V_TOP.t12 39.4005
R46 bgr_0.V_TOP.n10 bgr_0.V_TOP.t9 39.4005
R47 bgr_0.V_TOP.n9 bgr_0.V_TOP.t8 39.4005
R48 bgr_0.V_TOP.n9 bgr_0.V_TOP.t11 39.4005
R49 bgr_0.V_TOP.n14 bgr_0.V_TOP.t5 39.4005
R50 bgr_0.V_TOP.n14 bgr_0.V_TOP.t6 39.4005
R51 bgr_0.V_TOP.n16 bgr_0.V_TOP.t2 39.4005
R52 bgr_0.V_TOP.n16 bgr_0.V_TOP.t10 39.4005
R53 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 8.313
R54 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R55 bgr_0.V_TOP.n28 bgr_0.V_TOP.t49 4.8295
R56 bgr_0.V_TOP.n29 bgr_0.V_TOP.t25 4.8295
R57 bgr_0.V_TOP.n31 bgr_0.V_TOP.t21 4.8295
R58 bgr_0.V_TOP.n32 bgr_0.V_TOP.t34 4.8295
R59 bgr_0.V_TOP.n34 bgr_0.V_TOP.t30 4.8295
R60 bgr_0.V_TOP.n35 bgr_0.V_TOP.t46 4.8295
R61 bgr_0.V_TOP.n37 bgr_0.V_TOP.t24 4.8295
R62 bgr_0.V_TOP.n28 bgr_0.V_TOP.t39 4.5005
R63 bgr_0.V_TOP.n30 bgr_0.V_TOP.t28 4.5005
R64 bgr_0.V_TOP.n29 bgr_0.V_TOP.t33 4.5005
R65 bgr_0.V_TOP.n31 bgr_0.V_TOP.t15 4.5005
R66 bgr_0.V_TOP.n33 bgr_0.V_TOP.t40 4.5005
R67 bgr_0.V_TOP.n32 bgr_0.V_TOP.t45 4.5005
R68 bgr_0.V_TOP.n34 bgr_0.V_TOP.t22 4.5005
R69 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 4.5005
R70 bgr_0.V_TOP.n35 bgr_0.V_TOP.t19 4.5005
R71 bgr_0.V_TOP.n37 bgr_0.V_TOP.t17 4.5005
R72 bgr_0.V_TOP.n38 bgr_0.V_TOP.t42 4.5005
R73 bgr_0.V_TOP.n39 bgr_0.V_TOP.t47 4.5005
R74 bgr_0.V_TOP.n40 bgr_0.V_TOP.t36 4.5005
R75 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R76 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R77 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R78 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R79 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R80 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R81 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R82 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R83 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R84 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R85 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R86 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R87 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R88 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R89 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R90 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R91 bgr_0.Vin-.n21 bgr_0.Vin-.n20 1850.93
R92 bgr_0.Vin-.n9 bgr_0.Vin-.t10 688.859
R93 bgr_0.Vin-.n11 bgr_0.Vin-.n10 514.134
R94 bgr_0.Vin-.n7 bgr_0.Vin-.n6 345.115
R95 bgr_0.Vin-.n13 bgr_0.Vin-.n12 214.713
R96 bgr_0.Vin-.n9 bgr_0.Vin-.t12 174.726
R97 bgr_0.Vin-.n10 bgr_0.Vin-.t8 174.726
R98 bgr_0.Vin-.n11 bgr_0.Vin-.t11 174.726
R99 bgr_0.Vin-.n12 bgr_0.Vin-.t9 174.726
R100 bgr_0.Vin-.n5 bgr_0.Vin-.n3 173.029
R101 bgr_0.Vin-.n5 bgr_0.Vin-.n4 168.654
R102 bgr_0.Vin-.n7 bgr_0.Vin-.t1 162.921
R103 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R104 bgr_0.Vin-.n12 bgr_0.Vin-.n11 128.534
R105 bgr_0.Vin-.n22 bgr_0.Vin-.n21 84.0884
R106 bgr_0.Vin-.n17 bgr_0.Vin-.n16 83.5719
R107 bgr_0.Vin-.n18 bgr_0.Vin-.n0 83.5719
R108 bgr_0.Vin-.n19 bgr_0.Vin-.n1 83.5719
R109 bgr_0.Vin-.n14 bgr_0.Vin-.t0 65.0299
R110 bgr_0.Vin-.n6 bgr_0.Vin-.t6 39.4005
R111 bgr_0.Vin-.n6 bgr_0.Vin-.t7 39.4005
R112 bgr_0.Vin-.n18 bgr_0.Vin-.n17 26.074
R113 bgr_0.Vin-.n19 bgr_0.Vin-.n18 26.074
R114 bgr_0.Vin-.n21 bgr_0.Vin-.n19 26.074
R115 bgr_0.Vin-.n23 bgr_0.Vin-.n13 17.526
R116 bgr_0.Vin-.n4 bgr_0.Vin-.t3 13.1338
R117 bgr_0.Vin-.n4 bgr_0.Vin-.t2 13.1338
R118 bgr_0.Vin-.n3 bgr_0.Vin-.t5 13.1338
R119 bgr_0.Vin-.n3 bgr_0.Vin-.t4 13.1338
R120 bgr_0.Vin-.n13 bgr_0.Vin-.n8 12.5317
R121 bgr_0.Vin-.n8 bgr_0.Vin-.n7 6.40675
R122 bgr_0.Vin-.n8 bgr_0.Vin-.n5 3.8755
R123 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56363
R124 bgr_0.Vin-.n23 bgr_0.Vin-.n22 1.5505
R125 bgr_0.Vin-.n25 bgr_0.Vin-.n24 1.5505
R126 bgr_0.Vin-.n15 bgr_0.Vin-.n2 1.5505
R127 bgr_0.Vin-.n22 bgr_0.Vin-.n1 1.14402
R128 bgr_0.Vin-.n15 bgr_0.Vin-.n0 0.885803
R129 bgr_0.Vin-.n16 bgr_0.Vin-.n15 0.77514
R130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.756696
R131 bgr_0.Vin-.n25 bgr_0.Vin-.n1 0.701365
R132 bgr_0.Vin-.n14 bgr_0.Vin-.n2 0.537712
R133 bgr_0.Vin-.n17 bgr_0.Vin-.t0 0.290206
R134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n25 0.203382
R135 bgr_0.Vin-.n24 bgr_0.Vin-.n2 0.0183571
R136 bgr_0.Vin-.n24 bgr_0.Vin-.n23 0.0183571
R137 VDDA.n376 VDDA.n343 6600
R138 VDDA.n378 VDDA.n343 6600
R139 VDDA.n378 VDDA.n344 6570
R140 VDDA.n376 VDDA.n344 6570
R141 VDDA.n331 VDDA.n266 4710
R142 VDDA.n331 VDDA.n267 4710
R143 VDDA.n333 VDDA.n266 4710
R144 VDDA.n333 VDDA.n267 4710
R145 VDDA.n289 VDDA.n288 4710
R146 VDDA.n291 VDDA.n288 4710
R147 VDDA.n289 VDDA.n282 4710
R148 VDDA.n291 VDDA.n282 4710
R149 VDDA.n71 VDDA.n55 4605
R150 VDDA.n69 VDDA.n55 4605
R151 VDDA.n143 VDDA.n139 4605
R152 VDDA.n143 VDDA.n140 4605
R153 VDDA.n181 VDDA.n155 4590
R154 VDDA.n179 VDDA.n155 4590
R155 VDDA.n179 VDDA.n156 4590
R156 VDDA.n181 VDDA.n156 4590
R157 VDDA.n69 VDDA.n56 4575
R158 VDDA.n71 VDDA.n56 4575
R159 VDDA.n145 VDDA.n140 4575
R160 VDDA.n145 VDDA.n139 4575
R161 VDDA.n208 VDDA.n199 4020
R162 VDDA.n208 VDDA.n200 4020
R163 VDDA.n206 VDDA.n199 4020
R164 VDDA.n206 VDDA.n200 4020
R165 VDDA.n96 VDDA.n87 4020
R166 VDDA.n96 VDDA.n88 4020
R167 VDDA.n94 VDDA.n87 4020
R168 VDDA.n94 VDDA.n88 4020
R169 VDDA.n442 VDDA.n410 3420
R170 VDDA.n444 VDDA.n410 3420
R171 VDDA.n444 VDDA.n411 3420
R172 VDDA.n442 VDDA.n411 3420
R173 VDDA.n48 VDDA.n41 3390
R174 VDDA.n50 VDDA.n41 3390
R175 VDDA.n48 VDDA.n47 3390
R176 VDDA.n50 VDDA.n47 3390
R177 VDDA.n134 VDDA.n127 3390
R178 VDDA.n136 VDDA.n127 3390
R179 VDDA.n134 VDDA.n133 3390
R180 VDDA.n136 VDDA.n133 3390
R181 VDDA.n21 VDDA.n16 2940
R182 VDDA.n23 VDDA.n16 2940
R183 VDDA.n23 VDDA.n20 2940
R184 VDDA.n21 VDDA.n20 2940
R185 VDDA.n30 VDDA.n12 2940
R186 VDDA.n32 VDDA.n12 2940
R187 VDDA.n32 VDDA.n29 2940
R188 VDDA.n30 VDDA.n29 2940
R189 VDDA.n229 VDDA.n226 2520
R190 VDDA.n232 VDDA.n225 2505
R191 VDDA.n232 VDDA.n226 2475
R192 VDDA.n229 VDDA.n225 2220
R193 VDDA.n458 VDDA.n404 2145
R194 VDDA.n458 VDDA.n405 2100
R195 VDDA.n455 VDDA.n405 2100
R196 VDDA.n423 VDDA.n416 2100
R197 VDDA.n425 VDDA.n416 2100
R198 VDDA.n425 VDDA.n417 2100
R199 VDDA.n423 VDDA.n417 2100
R200 VDDA.n455 VDDA.n404 2055
R201 VDDA.n391 VDDA.n389 1770
R202 VDDA.n393 VDDA.n389 1770
R203 VDDA.n391 VDDA.n386 1770
R204 VDDA.n393 VDDA.n386 1770
R205 VDDA.n352 VDDA.n350 1770
R206 VDDA.n354 VDDA.n350 1770
R207 VDDA.n352 VDDA.n347 1770
R208 VDDA.n354 VDDA.n347 1770
R209 VDDA.n247 VDDA.n243 1566
R210 VDDA.n247 VDDA.n242 1566
R211 VDDA.n246 VDDA.n242 1536
R212 VDDA.n246 VDDA.n243 1536
R213 VDDA.n74 VDDA.t324 1216.42
R214 VDDA.n66 VDDA.t345 1216.42
R215 VDDA.n124 VDDA.t339 1216.42
R216 VDDA.n148 VDDA.t369 1216.42
R217 VDDA.n375 VDDA.n342 704
R218 VDDA.n379 VDDA.n342 704
R219 VDDA.n17 VDDA.t356 689.4
R220 VDDA.n25 VDDA.t380 689.4
R221 VDDA.n13 VDDA.t426 689.4
R222 VDDA.n34 VDDA.t320 689.4
R223 VDDA.n235 VDDA.t312 666.134
R224 VDDA.n223 VDDA.t403 666.134
R225 VDDA.n185 VDDA.t408 663.801
R226 VDDA.n175 VDDA.t402 663.801
R227 VDDA.n203 VDDA.t394 660.109
R228 VDDA.n201 VDDA.t360 660.109
R229 VDDA.n91 VDDA.t415 660.109
R230 VDDA.n89 VDDA.t366 660.109
R231 VDDA.t403 VDDA.n222 658.101
R232 VDDA.n444 VDDA.t413 652.576
R233 VDDA.n239 VDDA.t386 650.668
R234 VDDA.n251 VDDA.t393 650.668
R235 VDDA.n216 VDDA.n215 625.254
R236 VDDA.n174 VDDA.n173 622.268
R237 VDDA.n172 VDDA.n171 622.268
R238 VDDA.n170 VDDA.n169 622.268
R239 VDDA.n168 VDDA.n167 622.268
R240 VDDA.n166 VDDA.n165 622.268
R241 VDDA.n164 VDDA.n163 622.268
R242 VDDA.n162 VDDA.n161 622.268
R243 VDDA.n160 VDDA.n159 622.268
R244 VDDA.n158 VDDA.n157 622.268
R245 VDDA.n152 VDDA.n151 622.268
R246 VDDA.n42 VDDA.t357 573.75
R247 VDDA.n44 VDDA.t327 573.75
R248 VDDA.n128 VDDA.t375 573.75
R249 VDDA.n130 VDDA.t351 573.75
R250 VDDA.n374 VDDA.n341 518.4
R251 VDDA.n380 VDDA.n341 518.4
R252 VDDA.n293 VDDA.n292 496
R253 VDDA.n293 VDDA.n281 496
R254 VDDA.n72 VDDA.n54 491.2
R255 VDDA.n68 VDDA.n54 491.2
R256 VDDA.n142 VDDA.n141 491.2
R257 VDDA.n142 VDDA.n114 491.2
R258 VDDA.n182 VDDA.n154 489.601
R259 VDDA.n178 VDDA.n154 489.601
R260 VDDA.n387 VDDA.t330 419.108
R261 VDDA.n384 VDDA.t333 419.108
R262 VDDA.n209 VDDA.n198 416
R263 VDDA.n209 VDDA.n197 416
R264 VDDA.n97 VDDA.n86 416
R265 VDDA.n97 VDDA.n85 416
R266 VDDA.n348 VDDA.t409 413.084
R267 VDDA.n345 VDDA.t381 413.084
R268 VDDA.n452 VDDA.t397 409.067
R269 VDDA.n461 VDDA.t336 409.067
R270 VDDA.n439 VDDA.t418 409.067
R271 VDDA.n447 VDDA.t412 409.067
R272 VDDA.n420 VDDA.t315 409.067
R273 VDDA.n428 VDDA.t372 390.322
R274 VDDA.t425 VDDA.n29 389.375
R275 VDDA.t319 VDDA.n12 389.375
R276 VDDA.n181 VDDA.t407 389.375
R277 VDDA.t401 VDDA.n179 389.375
R278 VDDA.n387 VDDA.t332 389.185
R279 VDDA.n384 VDDA.t335 389.185
R280 VDDA.n439 VDDA.t420 387.051
R281 VDDA.n447 VDDA.t414 387.051
R282 VDDA.n264 VDDA.t350 384.918
R283 VDDA.n268 VDDA.t323 384.918
R284 VDDA.n283 VDDA.t365 384.918
R285 VDDA.n285 VDDA.t423 384.918
R286 VDDA.n348 VDDA.t411 384.918
R287 VDDA.n345 VDDA.t383 384.918
R288 VDDA.t355 VDDA.n20 384.168
R289 VDDA.t379 VDDA.n16 384.168
R290 VDDA.n270 VDDA.n269 384
R291 VDDA.n269 VDDA.n265 384
R292 VDDA.n287 VDDA.n286 384
R293 VDDA.n287 VDDA.n284 384
R294 VDDA.n183 VDDA.n153 377.601
R295 VDDA.n177 VDDA.n153 377.601
R296 VDDA.n420 VDDA.t317 370.728
R297 VDDA.n428 VDDA.t374 370.728
R298 VDDA.n452 VDDA.t399 370.3
R299 VDDA.n461 VDDA.t338 370.3
R300 VDDA.n441 VDDA.n409 364.8
R301 VDDA.n445 VDDA.n409 364.8
R302 VDDA.n373 VDDA.t342 360.868
R303 VDDA.n381 VDDA.t387 360.868
R304 VDDA.n264 VDDA.t348 358.858
R305 VDDA.n268 VDDA.t321 358.858
R306 VDDA.n283 VDDA.t363 358.858
R307 VDDA.n285 VDDA.t421 358.858
R308 VDDA.n52 VDDA.n51 355.2
R309 VDDA.n52 VDDA.n40 355.2
R310 VDDA.n138 VDDA.n137 355.2
R311 VDDA.n138 VDDA.n126 355.2
R312 VDDA.t322 VDDA.n331 351.591
R313 VDDA.n333 VDDA.t349 351.591
R314 VDDA.t422 VDDA.n289 351.591
R315 VDDA.n291 VDDA.t364 351.591
R316 VDDA.t385 VDDA.n242 349.546
R317 VDDA.t391 VDDA.n243 349.546
R318 VDDA.n413 VDDA.n412 345.127
R319 VDDA.n419 VDDA.n418 345.127
R320 VDDA.n401 VDDA.n400 344.7
R321 VDDA.n450 VDDA.n449 344.7
R322 VDDA.t334 VDDA.n391 344.394
R323 VDDA.n393 VDDA.t331 344.394
R324 VDDA.t382 VDDA.n352 344.394
R325 VDDA.n354 VDDA.t410 344.394
R326 VDDA.t398 VDDA.n455 344.394
R327 VDDA.n458 VDDA.t337 344.394
R328 VDDA.n275 VDDA.n273 342.3
R329 VDDA.n303 VDDA.n302 341.675
R330 VDDA.n301 VDDA.n300 341.675
R331 VDDA.n299 VDDA.n298 341.675
R332 VDDA.n297 VDDA.n296 341.675
R333 VDDA.n279 VDDA.n278 341.675
R334 VDDA.n277 VDDA.n276 341.675
R335 VDDA.n275 VDDA.n274 341.675
R336 VDDA.t419 VDDA.n442 340.635
R337 VDDA.t316 VDDA.n423 340.635
R338 VDDA.n425 VDDA.t373 340.635
R339 VDDA.n407 VDDA.n406 339.272
R340 VDDA.n431 VDDA.n430 339.272
R341 VDDA.n433 VDDA.n432 339.272
R342 VDDA.n435 VDDA.n434 339.272
R343 VDDA.n437 VDDA.n436 339.272
R344 VDDA.n336 VDDA.n260 337.175
R345 VDDA.n262 VDDA.n261 337.175
R346 VDDA.n312 VDDA.n311 337.175
R347 VDDA.n315 VDDA.n309 337.175
R348 VDDA.n307 VDDA.n306 337.175
R349 VDDA.n319 VDDA.n318 337.175
R350 VDDA.n322 VDDA.n305 337.175
R351 VDDA.n325 VDDA.n324 337.175
R352 VDDA.n328 VDDA.n272 337.175
R353 VDDA.n294 VDDA.n280 337.175
R354 VDDA.n397 VDDA.n383 335.022
R355 VDDA.n17 VDDA.t354 332.75
R356 VDDA.n25 VDDA.t378 332.75
R357 VDDA.n13 VDDA.t424 332.75
R358 VDDA.n34 VDDA.t318 332.75
R359 VDDA.n184 VDDA.t406 332.75
R360 VDDA.n176 VDDA.t400 332.75
R361 VDDA.n19 VDDA.n15 313.601
R362 VDDA.n240 VDDA.t384 310.659
R363 VDDA.n250 VDDA.t390 310.659
R364 VDDA.n27 VDDA.n15 307.2
R365 VDDA.n36 VDDA.n11 307.2
R366 VDDA.n28 VDDA.n11 307.2
R367 VDDA.t328 VDDA.n48 285.815
R368 VDDA.n50 VDDA.t358 285.815
R369 VDDA.t352 VDDA.n134 285.815
R370 VDDA.n136 VDDA.t376 285.815
R371 VDDA.t343 VDDA.n376 278.95
R372 VDDA.n378 VDDA.t388 278.95
R373 VDDA.n42 VDDA.t359 277.916
R374 VDDA.n44 VDDA.t329 277.916
R375 VDDA.n128 VDDA.t377 277.916
R376 VDDA.n130 VDDA.t353 277.916
R377 VDDA.n373 VDDA.t344 270.705
R378 VDDA.n381 VDDA.t389 270.705
R379 VDDA.n228 VDDA.n219 268.8
R380 VDDA.n73 VDDA.n72 267.2
R381 VDDA.n68 VDDA.n67 267.2
R382 VDDA.n141 VDDA.n125 267.2
R383 VDDA.n147 VDDA.n114 267.2
R384 VDDA.n440 VDDA.n408 246.4
R385 VDDA.t361 VDDA.n199 239.915
R386 VDDA.t395 VDDA.n200 239.915
R387 VDDA.t367 VDDA.n87 239.915
R388 VDDA.t416 VDDA.n88 239.915
R389 VDDA.n228 VDDA.n227 236.8
R390 VDDA.n459 VDDA.n403 228.8
R391 VDDA.n422 VDDA.n415 224
R392 VDDA.n426 VDDA.n415 224
R393 VDDA.n205 VDDA.n202 220.8
R394 VDDA.n205 VDDA.n204 220.8
R395 VDDA.n93 VDDA.n90 220.8
R396 VDDA.n93 VDDA.n92 220.8
R397 VDDA.n454 VDDA.n403 219.201
R398 VDDA.n227 VDDA.n224 206.4
R399 VDDA.n24 VDDA.n18 201.601
R400 VDDA.n26 VDDA.n24 201.601
R401 VDDA.n35 VDDA.n33 201.601
R402 VDDA.n46 VDDA.n45 201.601
R403 VDDA.n46 VDDA.n43 201.601
R404 VDDA.n132 VDDA.n131 201.601
R405 VDDA.n132 VDDA.n129 201.601
R406 VDDA.n67 VDDA.n53 195.201
R407 VDDA.n73 VDDA.n53 195.201
R408 VDDA.n147 VDDA.n146 195.201
R409 VDDA.n146 VDDA.n125 195.201
R410 VDDA.n33 VDDA.n14 193.371
R411 VDDA.t8 VDDA.t385 191.919
R412 VDDA.t8 VDDA.t391 191.919
R413 VDDA.n234 VDDA.n219 190.4
R414 VDDA.n204 VDDA.n198 188.8
R415 VDDA.n202 VDDA.n197 188.8
R416 VDDA.n92 VDDA.n86 188.8
R417 VDDA.n90 VDDA.n85 188.8
R418 VDDA.n335 VDDA.n334 188.8
R419 VDDA.n330 VDDA.n329 188.8
R420 VDDA.n394 VDDA.n388 188.8
R421 VDDA.n390 VDDA.n388 188.8
R422 VDDA.n355 VDDA.n349 188.8
R423 VDDA.n351 VDDA.n349 188.8
R424 VDDA.n446 VDDA.n445 188.8
R425 VDDA.t99 VDDA.t425 186.607
R426 VDDA.t452 VDDA.t99 186.607
R427 VDDA.t70 VDDA.t452 186.607
R428 VDDA.t218 VDDA.t70 186.607
R429 VDDA.t254 VDDA.t218 186.607
R430 VDDA.t45 VDDA.t82 186.607
R431 VDDA.t82 VDDA.t253 186.607
R432 VDDA.t253 VDDA.t135 186.607
R433 VDDA.t135 VDDA.t225 186.607
R434 VDDA.t225 VDDA.t319 186.607
R435 VDDA.t407 VDDA.t221 186.607
R436 VDDA.t221 VDDA.t210 186.607
R437 VDDA.t210 VDDA.t431 186.607
R438 VDDA.t431 VDDA.t28 186.607
R439 VDDA.t28 VDDA.t151 186.607
R440 VDDA.t151 VDDA.t219 186.607
R441 VDDA.t219 VDDA.t157 186.607
R442 VDDA.t157 VDDA.t86 186.607
R443 VDDA.t86 VDDA.t251 186.607
R444 VDDA.t251 VDDA.t467 186.607
R445 VDDA.t465 VDDA.t223 186.607
R446 VDDA.t223 VDDA.t126 186.607
R447 VDDA.t126 VDDA.t26 186.607
R448 VDDA.t26 VDDA.t212 186.607
R449 VDDA.t212 VDDA.t427 186.607
R450 VDDA.t427 VDDA.t149 186.607
R451 VDDA.t149 VDDA.t79 186.607
R452 VDDA.t79 VDDA.t463 186.607
R453 VDDA.t463 VDDA.t62 186.607
R454 VDDA.t62 VDDA.t401 186.607
R455 VDDA.t175 VDDA.t355 183.333
R456 VDDA.t102 VDDA.t175 183.333
R457 VDDA.t451 VDDA.t102 183.333
R458 VDDA.t144 VDDA.t451 183.333
R459 VDDA.t174 VDDA.t144 183.333
R460 VDDA.t43 VDDA.t98 183.333
R461 VDDA.t98 VDDA.t201 183.333
R462 VDDA.t201 VDDA.t119 183.333
R463 VDDA.t119 VDDA.t447 183.333
R464 VDDA.t447 VDDA.t379 183.333
R465 VDDA.n375 VDDA.n374 182.4
R466 VDDA.n380 VDDA.n379 182.4
R467 VDDA.n75 VDDA.t326 178.124
R468 VDDA.n65 VDDA.t347 178.124
R469 VDDA.n123 VDDA.t341 178.124
R470 VDDA.n149 VDDA.t371 178.124
R471 VDDA.n446 VDDA.n408 176
R472 VDDA.t111 VDDA.t322 172.727
R473 VDDA.t36 VDDA.t111 172.727
R474 VDDA.t208 VDDA.t36 172.727
R475 VDDA.t458 VDDA.t208 172.727
R476 VDDA.t170 VDDA.t458 172.727
R477 VDDA.t60 VDDA.t170 172.727
R478 VDDA.t120 VDDA.t60 172.727
R479 VDDA.t77 VDDA.t120 172.727
R480 VDDA.t34 VDDA.t77 172.727
R481 VDDA.t24 VDDA.t38 172.727
R482 VDDA.t433 VDDA.t24 172.727
R483 VDDA.t199 VDDA.t433 172.727
R484 VDDA.t206 VDDA.t199 172.727
R485 VDDA.t75 VDDA.t206 172.727
R486 VDDA.t124 VDDA.t75 172.727
R487 VDDA.t183 VDDA.t124 172.727
R488 VDDA.t46 VDDA.t183 172.727
R489 VDDA.t349 VDDA.t46 172.727
R490 VDDA.t50 VDDA.t422 172.727
R491 VDDA.t56 VDDA.t50 172.727
R492 VDDA.t54 VDDA.t56 172.727
R493 VDDA.t155 VDDA.t54 172.727
R494 VDDA.t145 VDDA.t155 172.727
R495 VDDA.t66 VDDA.t145 172.727
R496 VDDA.t96 VDDA.t66 172.727
R497 VDDA.t153 VDDA.t96 172.727
R498 VDDA.t58 VDDA.t153 172.727
R499 VDDA.t147 VDDA.t159 172.727
R500 VDDA.t100 VDDA.t147 172.727
R501 VDDA.t108 VDDA.t100 172.727
R502 VDDA.t52 VDDA.t108 172.727
R503 VDDA.t437 VDDA.t52 172.727
R504 VDDA.t161 VDDA.t437 172.727
R505 VDDA.t216 VDDA.t161 172.727
R506 VDDA.t64 VDDA.t216 172.727
R507 VDDA.t364 VDDA.t64 172.727
R508 VDDA.n220 VDDA.n218 170.534
R509 VDDA.n340 VDDA.n339 168.435
R510 VDDA.n359 VDDA.n358 168.435
R511 VDDA.n361 VDDA.n360 168.435
R512 VDDA.n363 VDDA.n362 168.435
R513 VDDA.n365 VDDA.n364 168.435
R514 VDDA.n367 VDDA.n366 168.435
R515 VDDA.n369 VDDA.n368 168.435
R516 VDDA.n371 VDDA.n370 168.435
R517 VDDA.n245 VDDA.n244 163.84
R518 VDDA.n245 VDDA.n217 163.84
R519 VDDA.n71 VDDA.t325 161.817
R520 VDDA.t346 VDDA.n69 161.817
R521 VDDA.t340 VDDA.n139 161.817
R522 VDDA.t370 VDDA.n140 161.817
R523 VDDA.t313 VDDA.n226 161.733
R524 VDDA.t268 VDDA.t343 159.814
R525 VDDA.t289 VDDA.t268 159.814
R526 VDDA.t300 VDDA.t289 159.814
R527 VDDA.t310 VDDA.t300 159.814
R528 VDDA.t275 VDDA.t310 159.814
R529 VDDA.t271 VDDA.t275 159.814
R530 VDDA.t294 VDDA.t271 159.814
R531 VDDA.t302 VDDA.t294 159.814
R532 VDDA.t280 VDDA.t261 159.814
R533 VDDA.t278 VDDA.t280 159.814
R534 VDDA.t296 VDDA.t278 159.814
R535 VDDA.t305 VDDA.t296 159.814
R536 VDDA.t266 VDDA.t305 159.814
R537 VDDA.t286 VDDA.t266 159.814
R538 VDDA.t284 VDDA.t286 159.814
R539 VDDA.t388 VDDA.t284 159.814
R540 VDDA.t404 VDDA.n225 159.147
R541 VDDA.t106 VDDA.t334 158.333
R542 VDDA.t331 VDDA.t445 158.333
R543 VDDA.t429 VDDA.t382 158.333
R544 VDDA.t410 VDDA.t430 158.333
R545 VDDA.t164 VDDA.t398 158.333
R546 VDDA.t115 VDDA.t164 158.333
R547 VDDA.t204 VDDA.t449 158.333
R548 VDDA.t337 VDDA.t204 158.333
R549 VDDA.t73 VDDA.t419 155.97
R550 VDDA.t454 VDDA.t73 155.97
R551 VDDA.t181 VDDA.t454 155.97
R552 VDDA.t48 VDDA.t181 155.97
R553 VDDA.t140 VDDA.t48 155.97
R554 VDDA.t202 VDDA.t140 155.97
R555 VDDA.t16 VDDA.t94 155.97
R556 VDDA.t179 VDDA.t16 155.97
R557 VDDA.t91 VDDA.t179 155.97
R558 VDDA.t413 VDDA.t91 155.97
R559 VDDA.t142 VDDA.t316 155.97
R560 VDDA.t71 VDDA.t142 155.97
R561 VDDA.t113 VDDA.t461 155.97
R562 VDDA.t373 VDDA.t113 155.97
R563 VDDA.n195 VDDA.n193 155.911
R564 VDDA.n192 VDDA.n190 155.911
R565 VDDA.n83 VDDA.n81 155.911
R566 VDDA.n80 VDDA.n78 155.911
R567 VDDA.n195 VDDA.n194 155.536
R568 VDDA.n192 VDDA.n191 155.536
R569 VDDA.n83 VDDA.n82 155.536
R570 VDDA.n80 VDDA.n79 155.536
R571 VDDA.n203 VDDA.t396 155.125
R572 VDDA.n201 VDDA.t362 155.125
R573 VDDA.n91 VDDA.t417 155.125
R574 VDDA.n89 VDDA.t368 155.125
R575 VDDA.n65 VDDA.n64 147.398
R576 VDDA.n123 VDDA.n122 147.398
R577 VDDA.n76 VDDA.n75 147.054
R578 VDDA.n150 VDDA.n149 147.054
R579 VDDA.n211 VDDA.n210 141.736
R580 VDDA.n99 VDDA.n98 141.736
R581 VDDA.n64 VDDA.n63 141.162
R582 VDDA.n62 VDDA.n61 141.162
R583 VDDA.n60 VDDA.n59 141.162
R584 VDDA.n58 VDDA.n57 141.162
R585 VDDA.n39 VDDA.n38 141.162
R586 VDDA.n113 VDDA.n112 141.162
R587 VDDA.n116 VDDA.n115 141.162
R588 VDDA.n118 VDDA.n117 141.162
R589 VDDA.n120 VDDA.n119 141.162
R590 VDDA.n122 VDDA.n121 141.162
R591 VDDA.n51 VDDA.n43 140.8
R592 VDDA.n45 VDDA.n40 140.8
R593 VDDA.n137 VDDA.n129 140.8
R594 VDDA.n131 VDDA.n126 140.8
R595 VDDA.n66 VDDA.n65 135.387
R596 VDDA.n75 VDDA.n74 135.387
R597 VDDA.n149 VDDA.n148 135.387
R598 VDDA.n124 VDDA.n123 135.387
R599 VDDA.t242 VDDA.t328 121.513
R600 VDDA.t249 VDDA.t242 121.513
R601 VDDA.t234 VDDA.t249 121.513
R602 VDDA.t196 VDDA.t234 121.513
R603 VDDA.t257 VDDA.t196 121.513
R604 VDDA.t243 VDDA.t132 121.513
R605 VDDA.t3 VDDA.t243 121.513
R606 VDDA.t241 VDDA.t3 121.513
R607 VDDA.t256 VDDA.t241 121.513
R608 VDDA.t358 VDDA.t256 121.513
R609 VDDA.t93 VDDA.t352 121.513
R610 VDDA.t215 VDDA.t93 121.513
R611 VDDA.t453 VDDA.t215 121.513
R612 VDDA.t83 VDDA.t453 121.513
R613 VDDA.t214 VDDA.t83 121.513
R614 VDDA.t435 VDDA.t443 121.513
R615 VDDA.t436 VDDA.t435 121.513
R616 VDDA.t81 VDDA.t436 121.513
R617 VDDA.t10 VDDA.t81 121.513
R618 VDDA.t376 VDDA.t10 121.513
R619 VDDA.n334 VDDA.n265 118.4
R620 VDDA.n330 VDDA.n270 118.4
R621 VDDA.n292 VDDA.n284 118.4
R622 VDDA.n286 VDDA.n281 118.4
R623 VDDA.n395 VDDA.n394 118.4
R624 VDDA.n390 VDDA.n385 118.4
R625 VDDA.n356 VDDA.n355 118.4
R626 VDDA.n351 VDDA.n346 118.4
R627 VDDA.n454 VDDA.n453 118.4
R628 VDDA.n460 VDDA.n459 118.4
R629 VDDA.n441 VDDA.n440 118.4
R630 VDDA.n422 VDDA.n421 118.4
R631 VDDA.n427 VDDA.n426 118.4
R632 VDDA.n453 VDDA.n402 105.6
R633 VDDA.n460 VDDA.n402 105.6
R634 VDDA.n421 VDDA.n414 105.6
R635 VDDA.n427 VDDA.n414 105.6
R636 VDDA.n237 VDDA.n236 105.534
R637 VDDA.n244 VDDA.n241 99.8405
R638 VDDA.n249 VDDA.n217 99.8405
R639 VDDA.t192 VDDA.t361 98.2764
R640 VDDA.t18 VDDA.t192 98.2764
R641 VDDA.t456 VDDA.t18 98.2764
R642 VDDA.t32 VDDA.t456 98.2764
R643 VDDA.t190 VDDA.t32 98.2764
R644 VDDA.t6 VDDA.t186 98.2764
R645 VDDA.t186 VDDA.t230 98.2764
R646 VDDA.t230 VDDA.t117 98.2764
R647 VDDA.t117 VDDA.t172 98.2764
R648 VDDA.t172 VDDA.t395 98.2764
R649 VDDA.t88 VDDA.t367 98.2764
R650 VDDA.t232 VDDA.t88 98.2764
R651 VDDA.t68 VDDA.t232 98.2764
R652 VDDA.t226 VDDA.t68 98.2764
R653 VDDA.t188 VDDA.t226 98.2764
R654 VDDA.t228 VDDA.t122 98.2764
R655 VDDA.t122 VDDA.t1 98.2764
R656 VDDA.t1 VDDA.t439 98.2764
R657 VDDA.t439 VDDA.t20 98.2764
R658 VDDA.t20 VDDA.t416 98.2764
R659 VDDA.t22 VDDA.t313 96.6107
R660 VDDA.n31 VDDA.t254 93.3041
R661 VDDA.n31 VDDA.t45 93.3041
R662 VDDA.t467 VDDA.n180 93.3041
R663 VDDA.n180 VDDA.t465 93.3041
R664 VDDA.n19 VDDA.n18 92.8005
R665 VDDA.n183 VDDA.n182 92.8005
R666 VDDA.n178 VDDA.n177 92.8005
R667 VDDA.n21 VDDA.n15 92.5005
R668 VDDA.n22 VDDA.n21 92.5005
R669 VDDA.n20 VDDA.n19 92.5005
R670 VDDA.n24 VDDA.n23 92.5005
R671 VDDA.n23 VDDA.n22 92.5005
R672 VDDA.n27 VDDA.n16 92.5005
R673 VDDA.n30 VDDA.n11 92.5005
R674 VDDA.n31 VDDA.n30 92.5005
R675 VDDA.n29 VDDA.n28 92.5005
R676 VDDA.n33 VDDA.n32 92.5005
R677 VDDA.n32 VDDA.n31 92.5005
R678 VDDA.n36 VDDA.n12 92.5005
R679 VDDA.n51 VDDA.n50 92.5005
R680 VDDA.n47 VDDA.n46 92.5005
R681 VDDA.n49 VDDA.n47 92.5005
R682 VDDA.n48 VDDA.n40 92.5005
R683 VDDA.n52 VDDA.n41 92.5005
R684 VDDA.n49 VDDA.n41 92.5005
R685 VDDA.n55 VDDA.n54 92.5005
R686 VDDA.n70 VDDA.n55 92.5005
R687 VDDA.n56 VDDA.n53 92.5005
R688 VDDA.n70 VDDA.n56 92.5005
R689 VDDA.n200 VDDA.n198 92.5005
R690 VDDA.n206 VDDA.n205 92.5005
R691 VDDA.n207 VDDA.n206 92.5005
R692 VDDA.n199 VDDA.n197 92.5005
R693 VDDA.n209 VDDA.n208 92.5005
R694 VDDA.n208 VDDA.n207 92.5005
R695 VDDA.n88 VDDA.n86 92.5005
R696 VDDA.n94 VDDA.n93 92.5005
R697 VDDA.n95 VDDA.n94 92.5005
R698 VDDA.n87 VDDA.n85 92.5005
R699 VDDA.n97 VDDA.n96 92.5005
R700 VDDA.n96 VDDA.n95 92.5005
R701 VDDA.n182 VDDA.n181 92.5005
R702 VDDA.n155 VDDA.n154 92.5005
R703 VDDA.n180 VDDA.n155 92.5005
R704 VDDA.n179 VDDA.n178 92.5005
R705 VDDA.n156 VDDA.n153 92.5005
R706 VDDA.n180 VDDA.n156 92.5005
R707 VDDA.n137 VDDA.n136 92.5005
R708 VDDA.n133 VDDA.n132 92.5005
R709 VDDA.n135 VDDA.n133 92.5005
R710 VDDA.n134 VDDA.n126 92.5005
R711 VDDA.n138 VDDA.n127 92.5005
R712 VDDA.n135 VDDA.n127 92.5005
R713 VDDA.n143 VDDA.n142 92.5005
R714 VDDA.n144 VDDA.n143 92.5005
R715 VDDA.n146 VDDA.n145 92.5005
R716 VDDA.n145 VDDA.n144 92.5005
R717 VDDA.n246 VDDA.n245 92.5005
R718 VDDA.t8 VDDA.n246 92.5005
R719 VDDA.n248 VDDA.n247 92.5005
R720 VDDA.n247 VDDA.t8 92.5005
R721 VDDA.n229 VDDA.n228 92.5005
R722 VDDA.n230 VDDA.n229 92.5005
R723 VDDA.n233 VDDA.n232 92.5005
R724 VDDA.n232 VDDA.n231 92.5005
R725 VDDA.n317 VDDA.n267 92.5005
R726 VDDA.n332 VDDA.n267 92.5005
R727 VDDA.n334 VDDA.n333 92.5005
R728 VDDA.n269 VDDA.n266 92.5005
R729 VDDA.n332 VDDA.n266 92.5005
R730 VDDA.n331 VDDA.n330 92.5005
R731 VDDA.n292 VDDA.n291 92.5005
R732 VDDA.n288 VDDA.n287 92.5005
R733 VDDA.n290 VDDA.n288 92.5005
R734 VDDA.n289 VDDA.n281 92.5005
R735 VDDA.n293 VDDA.n282 92.5005
R736 VDDA.n290 VDDA.n282 92.5005
R737 VDDA.n394 VDDA.n393 92.5005
R738 VDDA.n389 VDDA.n388 92.5005
R739 VDDA.n392 VDDA.n389 92.5005
R740 VDDA.n391 VDDA.n390 92.5005
R741 VDDA.n396 VDDA.n386 92.5005
R742 VDDA.n392 VDDA.n386 92.5005
R743 VDDA.n376 VDDA.n375 92.5005
R744 VDDA.n343 VDDA.n342 92.5005
R745 VDDA.n377 VDDA.n343 92.5005
R746 VDDA.n379 VDDA.n378 92.5005
R747 VDDA.n344 VDDA.n341 92.5005
R748 VDDA.n377 VDDA.n344 92.5005
R749 VDDA.n355 VDDA.n354 92.5005
R750 VDDA.n350 VDDA.n349 92.5005
R751 VDDA.n353 VDDA.n350 92.5005
R752 VDDA.n352 VDDA.n351 92.5005
R753 VDDA.n357 VDDA.n347 92.5005
R754 VDDA.n353 VDDA.n347 92.5005
R755 VDDA.n455 VDDA.n454 92.5005
R756 VDDA.n404 VDDA.n403 92.5005
R757 VDDA.n456 VDDA.n404 92.5005
R758 VDDA.n459 VDDA.n458 92.5005
R759 VDDA.n405 VDDA.n402 92.5005
R760 VDDA.n457 VDDA.n405 92.5005
R761 VDDA.n442 VDDA.n441 92.5005
R762 VDDA.n410 VDDA.n409 92.5005
R763 VDDA.n443 VDDA.n410 92.5005
R764 VDDA.n445 VDDA.n444 92.5005
R765 VDDA.n411 VDDA.n408 92.5005
R766 VDDA.n443 VDDA.n411 92.5005
R767 VDDA.n423 VDDA.n422 92.5005
R768 VDDA.n416 VDDA.n415 92.5005
R769 VDDA.n424 VDDA.n416 92.5005
R770 VDDA.n426 VDDA.n425 92.5005
R771 VDDA.n417 VDDA.n414 92.5005
R772 VDDA.n424 VDDA.n417 92.5005
R773 VDDA.n222 VDDA.n221 91.7338
R774 VDDA.n22 VDDA.t174 91.6672
R775 VDDA.n22 VDDA.t43 91.6672
R776 VDDA.n2 VDDA.n0 91.2452
R777 VDDA.n103 VDDA.n101 91.2452
R778 VDDA.n2 VDDA.n1 90.9014
R779 VDDA.n4 VDDA.n3 90.9014
R780 VDDA.n6 VDDA.n5 90.9014
R781 VDDA.n8 VDDA.n7 90.9014
R782 VDDA.n10 VDDA.n9 90.9014
R783 VDDA.n111 VDDA.n110 90.9014
R784 VDDA.n109 VDDA.n108 90.9014
R785 VDDA.n107 VDDA.n106 90.9014
R786 VDDA.n105 VDDA.n104 90.9014
R787 VDDA.n103 VDDA.n102 90.9014
R788 VDDA.n223 VDDA.n221 87.4672
R789 VDDA.n236 VDDA.n235 87.4672
R790 VDDA.n27 VDDA.n26 86.4005
R791 VDDA.n28 VDDA.n14 86.4005
R792 VDDA.n36 VDDA.n35 86.4005
R793 VDDA.n332 VDDA.t34 86.3641
R794 VDDA.t38 VDDA.n332 86.3641
R795 VDDA.n290 VDDA.t58 86.3641
R796 VDDA.t159 VDDA.n290 86.3641
R797 VDDA.n377 VDDA.t302 79.907
R798 VDDA.t261 VDDA.n377 79.907
R799 VDDA.n392 VDDA.t106 79.1672
R800 VDDA.t445 VDDA.n392 79.1672
R801 VDDA.n353 VDDA.t429 79.1672
R802 VDDA.t430 VDDA.n353 79.1672
R803 VDDA.t449 VDDA.n457 79.1672
R804 VDDA.n173 VDDA.t464 78.8005
R805 VDDA.n173 VDDA.t63 78.8005
R806 VDDA.n171 VDDA.t150 78.8005
R807 VDDA.n171 VDDA.t80 78.8005
R808 VDDA.n169 VDDA.t213 78.8005
R809 VDDA.n169 VDDA.t428 78.8005
R810 VDDA.n167 VDDA.t127 78.8005
R811 VDDA.n167 VDDA.t27 78.8005
R812 VDDA.n165 VDDA.t466 78.8005
R813 VDDA.n165 VDDA.t224 78.8005
R814 VDDA.n163 VDDA.t252 78.8005
R815 VDDA.n163 VDDA.t468 78.8005
R816 VDDA.n161 VDDA.t158 78.8005
R817 VDDA.n161 VDDA.t87 78.8005
R818 VDDA.n159 VDDA.t152 78.8005
R819 VDDA.n159 VDDA.t220 78.8005
R820 VDDA.n157 VDDA.t432 78.8005
R821 VDDA.n157 VDDA.t29 78.8005
R822 VDDA.n151 VDDA.t222 78.8005
R823 VDDA.n151 VDDA.t211 78.8005
R824 VDDA.n443 VDDA.t202 77.9856
R825 VDDA.t94 VDDA.n443 77.9856
R826 VDDA.n424 VDDA.t71 77.9856
R827 VDDA.t461 VDDA.n424 77.9856
R828 VDDA.n230 VDDA.t404 76.4836
R829 VDDA.n236 VDDA.t314 76.0991
R830 VDDA.n221 VDDA.t405 76.0991
R831 VDDA.n215 VDDA.t9 65.6672
R832 VDDA.n215 VDDA.t392 65.6672
R833 VDDA.n329 VDDA.n271 64.0005
R834 VDDA.n321 VDDA.n271 64.0005
R835 VDDA.n321 VDDA.n320 64.0005
R836 VDDA.n320 VDDA.n317 64.0005
R837 VDDA.n317 VDDA.n316 64.0005
R838 VDDA.n316 VDDA.n308 64.0005
R839 VDDA.n308 VDDA.n263 64.0005
R840 VDDA.n335 VDDA.n263 64.0005
R841 VDDA.n357 VDDA.n356 64.0005
R842 VDDA.n357 VDDA.n346 64.0005
R843 VDDA.t325 VDDA.t239 62.9523
R844 VDDA.t239 VDDA.t128 62.9523
R845 VDDA.t128 VDDA.t235 62.9523
R846 VDDA.t235 VDDA.t197 62.9523
R847 VDDA.t197 VDDA.t247 62.9523
R848 VDDA.t41 VDDA.t244 62.9523
R849 VDDA.t244 VDDA.t4 62.9523
R850 VDDA.t4 VDDA.t237 62.9523
R851 VDDA.t237 VDDA.t258 62.9523
R852 VDDA.t258 VDDA.t346 62.9523
R853 VDDA.t104 VDDA.t340 62.9523
R854 VDDA.t168 VDDA.t104 62.9523
R855 VDDA.t30 VDDA.t168 62.9523
R856 VDDA.t14 VDDA.t30 62.9523
R857 VDDA.t166 VDDA.t14 62.9523
R858 VDDA.t136 VDDA.t133 62.9523
R859 VDDA.t133 VDDA.t138 62.9523
R860 VDDA.t138 VDDA.t441 62.9523
R861 VDDA.t441 VDDA.t11 62.9523
R862 VDDA.t11 VDDA.t370 62.9523
R863 VDDA.n396 VDDA.n395 62.7205
R864 VDDA.n396 VDDA.n385 62.7205
R865 VDDA.n72 VDDA.n71 61.6672
R866 VDDA.n69 VDDA.n68 61.6672
R867 VDDA.n141 VDDA.n139 61.6672
R868 VDDA.n140 VDDA.n114 61.6672
R869 VDDA.n244 VDDA.n242 61.6672
R870 VDDA.n243 VDDA.n217 61.6672
R871 VDDA.n49 VDDA.t257 60.7563
R872 VDDA.t132 VDDA.n49 60.7563
R873 VDDA.n135 VDDA.t214 60.7563
R874 VDDA.t443 VDDA.n135 60.7563
R875 VDDA.n256 VDDA.t471 59.5681
R876 VDDA.n255 VDDA.t469 59.5681
R877 VDDA.n456 VDDA.t115 57.5763
R878 VDDA.n234 VDDA.n233 54.4005
R879 VDDA.n255 VDDA.t472 51.8888
R880 VDDA.n207 VDDA.t190 49.1384
R881 VDDA.n207 VDDA.t6 49.1384
R882 VDDA.n95 VDDA.t188 49.1384
R883 VDDA.n95 VDDA.t228 49.1384
R884 VDDA.n257 VDDA.t470 48.9557
R885 VDDA.n248 VDDA.n241 48.0005
R886 VDDA.n249 VDDA.n248 48.0005
R887 VDDA.n233 VDDA.n224 41.6005
R888 VDDA.n252 VDDA.n251 40.2538
R889 VDDA.n260 VDDA.t184 39.4005
R890 VDDA.n260 VDDA.t47 39.4005
R891 VDDA.n261 VDDA.t76 39.4005
R892 VDDA.n261 VDDA.t125 39.4005
R893 VDDA.n311 VDDA.t200 39.4005
R894 VDDA.n311 VDDA.t207 39.4005
R895 VDDA.n309 VDDA.t25 39.4005
R896 VDDA.n309 VDDA.t434 39.4005
R897 VDDA.n306 VDDA.t35 39.4005
R898 VDDA.n306 VDDA.t39 39.4005
R899 VDDA.n318 VDDA.t121 39.4005
R900 VDDA.n318 VDDA.t78 39.4005
R901 VDDA.n305 VDDA.t171 39.4005
R902 VDDA.n305 VDDA.t61 39.4005
R903 VDDA.n324 VDDA.t209 39.4005
R904 VDDA.n324 VDDA.t459 39.4005
R905 VDDA.n272 VDDA.t112 39.4005
R906 VDDA.n272 VDDA.t37 39.4005
R907 VDDA.n302 VDDA.t217 39.4005
R908 VDDA.n302 VDDA.t65 39.4005
R909 VDDA.n300 VDDA.t438 39.4005
R910 VDDA.n300 VDDA.t162 39.4005
R911 VDDA.n298 VDDA.t109 39.4005
R912 VDDA.n298 VDDA.t53 39.4005
R913 VDDA.n296 VDDA.t148 39.4005
R914 VDDA.n296 VDDA.t101 39.4005
R915 VDDA.n280 VDDA.t59 39.4005
R916 VDDA.n280 VDDA.t160 39.4005
R917 VDDA.n278 VDDA.t97 39.4005
R918 VDDA.n278 VDDA.t154 39.4005
R919 VDDA.n276 VDDA.t146 39.4005
R920 VDDA.n276 VDDA.t67 39.4005
R921 VDDA.n274 VDDA.t55 39.4005
R922 VDDA.n274 VDDA.t156 39.4005
R923 VDDA.n273 VDDA.t51 39.4005
R924 VDDA.n273 VDDA.t57 39.4005
R925 VDDA.n383 VDDA.t107 39.4005
R926 VDDA.n383 VDDA.t446 39.4005
R927 VDDA.n400 VDDA.t450 39.4005
R928 VDDA.n400 VDDA.t205 39.4005
R929 VDDA.n449 VDDA.t165 39.4005
R930 VDDA.n449 VDDA.t116 39.4005
R931 VDDA.n406 VDDA.t180 39.4005
R932 VDDA.n406 VDDA.t92 39.4005
R933 VDDA.n430 VDDA.t95 39.4005
R934 VDDA.n430 VDDA.t17 39.4005
R935 VDDA.n432 VDDA.t141 39.4005
R936 VDDA.n432 VDDA.t203 39.4005
R937 VDDA.n434 VDDA.t182 39.4005
R938 VDDA.n434 VDDA.t49 39.4005
R939 VDDA.n436 VDDA.t74 39.4005
R940 VDDA.n436 VDDA.t455 39.4005
R941 VDDA.n412 VDDA.t462 39.4005
R942 VDDA.n412 VDDA.t114 39.4005
R943 VDDA.n418 VDDA.t143 39.4005
R944 VDDA.n418 VDDA.t72 39.4005
R945 VDDA.n175 VDDA.n174 37.6109
R946 VDDA.n186 VDDA.n185 37.2672
R947 VDDA.n239 VDDA.n238 35.7538
R948 VDDA.t247 VDDA.n70 31.4764
R949 VDDA.n70 VDDA.t41 31.4764
R950 VDDA.n144 VDDA.t166 31.4764
R951 VDDA.n144 VDDA.t136 31.4764
R952 VDDA.n28 VDDA.n27 28.1943
R953 VDDA.n251 VDDA.n250 27.7338
R954 VDDA.n240 VDDA.n239 27.7338
R955 VDDA.n176 VDDA.n175 25.6005
R956 VDDA.n185 VDDA.n184 25.6005
R957 VDDA.n258 VDDA.n254 24.7265
R958 VDDA.n250 VDDA.n249 23.4672
R959 VDDA.n241 VDDA.n240 23.4672
R960 VDDA.n224 VDDA.n223 23.4672
R961 VDDA.n235 VDDA.n234 23.4672
R962 VDDA.n457 VDDA.n456 21.5914
R963 VDDA.n18 VDDA.n17 21.3338
R964 VDDA.n26 VDDA.n25 21.3338
R965 VDDA.n14 VDDA.n13 21.3338
R966 VDDA.n35 VDDA.n34 21.3338
R967 VDDA.n43 VDDA.n42 21.3338
R968 VDDA.n45 VDDA.n44 21.3338
R969 VDDA.n67 VDDA.n66 21.3338
R970 VDDA.n74 VDDA.n73 21.3338
R971 VDDA.n204 VDDA.n203 21.3338
R972 VDDA.n202 VDDA.n201 21.3338
R973 VDDA.n92 VDDA.n91 21.3338
R974 VDDA.n90 VDDA.n89 21.3338
R975 VDDA.n177 VDDA.n176 21.3338
R976 VDDA.n184 VDDA.n183 21.3338
R977 VDDA.n129 VDDA.n128 21.3338
R978 VDDA.n131 VDDA.n130 21.3338
R979 VDDA.n148 VDDA.n147 21.3338
R980 VDDA.n125 VDDA.n124 21.3338
R981 VDDA.n265 VDDA.n264 21.3338
R982 VDDA.n270 VDDA.n268 21.3338
R983 VDDA.n284 VDDA.n283 21.3338
R984 VDDA.n286 VDDA.n285 21.3338
R985 VDDA.n395 VDDA.n387 21.3338
R986 VDDA.n385 VDDA.n384 21.3338
R987 VDDA.n356 VDDA.n348 21.3338
R988 VDDA.n346 VDDA.n345 21.3338
R989 VDDA.n381 VDDA.n380 19.2005
R990 VDDA.n374 VDDA.n373 19.2005
R991 VDDA.n461 VDDA.n460 19.2005
R992 VDDA.n453 VDDA.n452 19.2005
R993 VDDA.n447 VDDA.n446 19.2005
R994 VDDA.n440 VDDA.n439 19.2005
R995 VDDA.n428 VDDA.n427 19.2005
R996 VDDA.n421 VDDA.n420 19.2005
R997 VDDA.n53 VDDA.n52 19.1318
R998 VDDA.n146 VDDA.n138 19.1318
R999 VDDA.n37 VDDA.n36 18.988
R1000 VDDA.n226 VDDA.n219 16.8187
R1001 VDDA.n254 VDDA.n253 16.5955
R1002 VDDA.n372 VDDA.n357 16.363
R1003 VDDA.n231 VDDA.t22 16.1022
R1004 VDDA.n211 VDDA.n209 16.0005
R1005 VDDA.n99 VDDA.n97 16.0005
R1006 VDDA.n468 VDDA.t270 15.0181
R1007 VDDA.n420 VDDA.n419 14.363
R1008 VDDA.n227 VDDA.n225 14.2313
R1009 VDDA.n222 VDDA.n218 13.988
R1010 VDDA.n373 VDDA.n372 13.8005
R1011 VDDA.n382 VDDA.n381 13.8005
R1012 VDDA.n452 VDDA.n451 13.8005
R1013 VDDA.n439 VDDA.n438 13.8005
R1014 VDDA.n429 VDDA.n428 13.8005
R1015 VDDA.n448 VDDA.n447 13.8005
R1016 VDDA.n462 VDDA.n461 13.8005
R1017 VDDA.n339 VDDA.t287 13.1338
R1018 VDDA.n339 VDDA.t285 13.1338
R1019 VDDA.n358 VDDA.t306 13.1338
R1020 VDDA.n358 VDDA.t267 13.1338
R1021 VDDA.n360 VDDA.t279 13.1338
R1022 VDDA.n360 VDDA.t297 13.1338
R1023 VDDA.n362 VDDA.t262 13.1338
R1024 VDDA.n362 VDDA.t281 13.1338
R1025 VDDA.n364 VDDA.t295 13.1338
R1026 VDDA.n364 VDDA.t303 13.1338
R1027 VDDA.n366 VDDA.t276 13.1338
R1028 VDDA.n366 VDDA.t272 13.1338
R1029 VDDA.n368 VDDA.t301 13.1338
R1030 VDDA.n368 VDDA.t311 13.1338
R1031 VDDA.n370 VDDA.t269 13.1338
R1032 VDDA.n370 VDDA.t290 13.1338
R1033 VDDA.n210 VDDA.t191 11.2576
R1034 VDDA.n210 VDDA.t7 11.2576
R1035 VDDA.n193 VDDA.t118 11.2576
R1036 VDDA.n193 VDDA.t173 11.2576
R1037 VDDA.n194 VDDA.t187 11.2576
R1038 VDDA.n194 VDDA.t231 11.2576
R1039 VDDA.n191 VDDA.t457 11.2576
R1040 VDDA.n191 VDDA.t33 11.2576
R1041 VDDA.n190 VDDA.t193 11.2576
R1042 VDDA.n190 VDDA.t19 11.2576
R1043 VDDA.n98 VDDA.t189 11.2576
R1044 VDDA.n98 VDDA.t229 11.2576
R1045 VDDA.n81 VDDA.t440 11.2576
R1046 VDDA.n81 VDDA.t21 11.2576
R1047 VDDA.n82 VDDA.t123 11.2576
R1048 VDDA.n82 VDDA.t2 11.2576
R1049 VDDA.n79 VDDA.t69 11.2576
R1050 VDDA.n79 VDDA.t227 11.2576
R1051 VDDA.n78 VDDA.t89 11.2576
R1052 VDDA.n78 VDDA.t233 11.2576
R1053 VDDA.n188 VDDA.n111 11.1255
R1054 VDDA.t405 VDDA.n220 11.0991
R1055 VDDA.n220 VDDA.t23 11.0991
R1056 VDDA.n37 VDDA.n10 9.64112
R1057 VDDA.n212 VDDA.n211 9.3005
R1058 VDDA.n100 VDDA.n99 9.3005
R1059 VDDA.n325 VDDA.n271 9.3005
R1060 VDDA.n322 VDDA.n321 9.3005
R1061 VDDA.n320 VDDA.n319 9.3005
R1062 VDDA.n317 VDDA.n307 9.3005
R1063 VDDA.n316 VDDA.n315 9.3005
R1064 VDDA.n312 VDDA.n308 9.3005
R1065 VDDA.n263 VDDA.n262 9.3005
R1066 VDDA.n336 VDDA.n335 9.3005
R1067 VDDA.n329 VDDA.n328 9.3005
R1068 VDDA.n294 VDDA.n293 9.3005
R1069 VDDA.n397 VDDA.n396 9.3005
R1070 VDDA.n258 VDDA.n257 8.03219
R1071 VDDA.n463 VDDA.n462 7.44175
R1072 VDDA.n189 VDDA.n188 7.07862
R1073 VDDA.n238 VDDA.n237 6.963
R1074 VDDA.n213 VDDA.n189 6.82862
R1075 VDDA.n63 VDDA.t238 6.56717
R1076 VDDA.n63 VDDA.t259 6.56717
R1077 VDDA.n61 VDDA.t245 6.56717
R1078 VDDA.n61 VDDA.t5 6.56717
R1079 VDDA.n59 VDDA.t248 6.56717
R1080 VDDA.n59 VDDA.t42 6.56717
R1081 VDDA.n57 VDDA.t236 6.56717
R1082 VDDA.n57 VDDA.t198 6.56717
R1083 VDDA.n38 VDDA.t240 6.56717
R1084 VDDA.n38 VDDA.t129 6.56717
R1085 VDDA.n112 VDDA.t442 6.56717
R1086 VDDA.n112 VDDA.t12 6.56717
R1087 VDDA.n115 VDDA.t134 6.56717
R1088 VDDA.n115 VDDA.t139 6.56717
R1089 VDDA.n117 VDDA.t167 6.56717
R1090 VDDA.n117 VDDA.t137 6.56717
R1091 VDDA.n119 VDDA.t31 6.56717
R1092 VDDA.n119 VDDA.t15 6.56717
R1093 VDDA.n121 VDDA.t105 6.56717
R1094 VDDA.n121 VDDA.t169 6.56717
R1095 VDDA.n189 VDDA.n100 6.34425
R1096 VDDA.n213 VDDA.n212 6.32862
R1097 VDDA.n399 VDDA.n398 6.13371
R1098 VDDA.n338 VDDA.n337 6.098
R1099 VDDA.n0 VDDA.t250 6.0005
R1100 VDDA.n0 VDDA.t444 6.0005
R1101 VDDA.n1 VDDA.t85 6.0005
R1102 VDDA.n1 VDDA.t195 6.0005
R1103 VDDA.n3 VDDA.t84 6.0005
R1104 VDDA.n3 VDDA.t194 6.0005
R1105 VDDA.n5 VDDA.t40 6.0005
R1106 VDDA.n5 VDDA.t130 6.0005
R1107 VDDA.n7 VDDA.t131 6.0005
R1108 VDDA.n7 VDDA.t246 6.0005
R1109 VDDA.n9 VDDA.t103 6.0005
R1110 VDDA.n9 VDDA.t255 6.0005
R1111 VDDA.n110 VDDA.t163 6.0005
R1112 VDDA.n110 VDDA.t176 6.0005
R1113 VDDA.n108 VDDA.t13 6.0005
R1114 VDDA.n108 VDDA.t185 6.0005
R1115 VDDA.n106 VDDA.t178 6.0005
R1116 VDDA.n106 VDDA.t448 6.0005
R1117 VDDA.n104 VDDA.t0 6.0005
R1118 VDDA.n104 VDDA.t460 6.0005
R1119 VDDA.n102 VDDA.t177 6.0005
R1120 VDDA.n102 VDDA.t90 6.0005
R1121 VDDA.n101 VDDA.t110 6.0005
R1122 VDDA.n101 VDDA.t44 6.0005
R1123 VDDA.n253 VDDA.n252 5.6255
R1124 VDDA.n77 VDDA.n76 5.03175
R1125 VDDA.n238 VDDA.n216 4.8755
R1126 VDDA.n212 VDDA.n196 4.5005
R1127 VDDA.n100 VDDA.n84 4.5005
R1128 VDDA.n188 VDDA.n187 4.5005
R1129 VDDA.n214 VDDA.n213 4.5005
R1130 VDDA.n295 VDDA.n294 4.5005
R1131 VDDA.n328 VDDA.n327 4.5005
R1132 VDDA.n326 VDDA.n325 4.5005
R1133 VDDA.n323 VDDA.n322 4.5005
R1134 VDDA.n319 VDDA.n304 4.5005
R1135 VDDA.n310 VDDA.n307 4.5005
R1136 VDDA.n315 VDDA.n314 4.5005
R1137 VDDA.n313 VDDA.n312 4.5005
R1138 VDDA.n262 VDDA.n259 4.5005
R1139 VDDA.n337 VDDA.n336 4.5005
R1140 VDDA.n398 VDDA.n397 4.5005
R1141 VDDA.n256 VDDA.n255 4.12334
R1142 VDDA.n469 VDDA 4.08025
R1143 VDDA.n231 VDDA.n230 4.02592
R1144 VDDA.n327 VDDA.n303 3.3755
R1145 VDDA.n257 VDDA.n256 2.93377
R1146 VDDA.n214 VDDA.n77 2.57862
R1147 VDDA.n451 VDDA.n448 2.5005
R1148 VDDA.n398 VDDA.n382 2.47371
R1149 VDDA.n438 VDDA.n429 1.813
R1150 VDDA.n187 VDDA.n186 1.51612
R1151 VDDA.n77 VDDA.n37 1.46925
R1152 VDDA VDDA.n469 1.20605
R1153 VDDA VDDA.n468 1.0815
R1154 VDDA.n372 VDDA.n371 1.0005
R1155 VDDA.n371 VDDA.n369 1.0005
R1156 VDDA.n369 VDDA.n367 1.0005
R1157 VDDA.n367 VDDA.n365 1.0005
R1158 VDDA.n365 VDDA.n363 1.0005
R1159 VDDA.n363 VDDA.n361 1.0005
R1160 VDDA.n361 VDDA.n359 1.0005
R1161 VDDA.n359 VDDA.n340 1.0005
R1162 VDDA.n382 VDDA.n340 1.0005
R1163 VDDA.n253 VDDA.n214 0.913
R1164 VDDA.n338 VDDA.n258 0.840625
R1165 VDDA.n469 VDDA.n254 0.8136
R1166 VDDA.n399 VDDA.n338 0.74075
R1167 VDDA.n277 VDDA.n275 0.6255
R1168 VDDA.n279 VDDA.n277 0.6255
R1169 VDDA.n295 VDDA.n279 0.6255
R1170 VDDA.n297 VDDA.n295 0.6255
R1171 VDDA.n299 VDDA.n297 0.6255
R1172 VDDA.n301 VDDA.n299 0.6255
R1173 VDDA.n303 VDDA.n301 0.6255
R1174 VDDA.n327 VDDA.n326 0.6255
R1175 VDDA.n326 VDDA.n323 0.6255
R1176 VDDA.n323 VDDA.n304 0.6255
R1177 VDDA.n310 VDDA.n304 0.6255
R1178 VDDA.n314 VDDA.n310 0.6255
R1179 VDDA.n314 VDDA.n313 0.6255
R1180 VDDA.n313 VDDA.n259 0.6255
R1181 VDDA.n337 VDDA.n259 0.6255
R1182 VDDA.n419 VDDA.n413 0.563
R1183 VDDA.n429 VDDA.n413 0.563
R1184 VDDA.n438 VDDA.n437 0.563
R1185 VDDA.n437 VDDA.n435 0.563
R1186 VDDA.n435 VDDA.n433 0.563
R1187 VDDA.n433 VDDA.n431 0.563
R1188 VDDA.n431 VDDA.n407 0.563
R1189 VDDA.n448 VDDA.n407 0.563
R1190 VDDA.n451 VDDA.n450 0.563
R1191 VDDA.n450 VDDA.n401 0.563
R1192 VDDA.n462 VDDA.n401 0.563
R1193 VDDA.n187 VDDA.n150 0.547375
R1194 VDDA.n463 VDDA.n399 0.546875
R1195 VDDA.n196 VDDA.n192 0.3755
R1196 VDDA.n196 VDDA.n195 0.3755
R1197 VDDA.n84 VDDA.n80 0.3755
R1198 VDDA.n84 VDDA.n83 0.3755
R1199 VDDA.n237 VDDA.n218 0.3755
R1200 VDDA.n468 VDDA.n463 0.370625
R1201 VDDA.n10 VDDA.n8 0.34425
R1202 VDDA.n8 VDDA.n6 0.34425
R1203 VDDA.n6 VDDA.n4 0.34425
R1204 VDDA.n4 VDDA.n2 0.34425
R1205 VDDA.n76 VDDA.n39 0.34425
R1206 VDDA.n58 VDDA.n39 0.34425
R1207 VDDA.n60 VDDA.n58 0.34425
R1208 VDDA.n62 VDDA.n60 0.34425
R1209 VDDA.n64 VDDA.n62 0.34425
R1210 VDDA.n105 VDDA.n103 0.34425
R1211 VDDA.n107 VDDA.n105 0.34425
R1212 VDDA.n109 VDDA.n107 0.34425
R1213 VDDA.n111 VDDA.n109 0.34425
R1214 VDDA.n122 VDDA.n120 0.34425
R1215 VDDA.n120 VDDA.n118 0.34425
R1216 VDDA.n118 VDDA.n116 0.34425
R1217 VDDA.n116 VDDA.n113 0.34425
R1218 VDDA.n150 VDDA.n113 0.34425
R1219 VDDA.n186 VDDA.n152 0.34425
R1220 VDDA.n158 VDDA.n152 0.34425
R1221 VDDA.n160 VDDA.n158 0.34425
R1222 VDDA.n162 VDDA.n160 0.34425
R1223 VDDA.n164 VDDA.n162 0.34425
R1224 VDDA.n166 VDDA.n164 0.34425
R1225 VDDA.n168 VDDA.n166 0.34425
R1226 VDDA.n170 VDDA.n168 0.34425
R1227 VDDA.n172 VDDA.n170 0.34425
R1228 VDDA.n174 VDDA.n172 0.34425
R1229 VDDA.n252 VDDA.n216 0.188
R1230 VDDA.t263 VDDA.t277 0.1603
R1231 VDDA.t307 VDDA.t299 0.1603
R1232 VDDA.t304 VDDA.t264 0.1603
R1233 VDDA.t292 VDDA.t288 0.1603
R1234 VDDA.t265 VDDA.t282 0.1603
R1235 VDDA.t309 VDDA.t293 0.1603
R1236 VDDA.t283 VDDA.t298 0.1603
R1237 VDDA.t274 VDDA.t260 0.1603
R1238 VDDA.n465 VDDA.t291 0.159278
R1239 VDDA.n466 VDDA.t273 0.159278
R1240 VDDA.n467 VDDA.t308 0.159278
R1241 VDDA.n467 VDDA.t263 0.1368
R1242 VDDA.n467 VDDA.t307 0.1368
R1243 VDDA.n466 VDDA.t304 0.1368
R1244 VDDA.n466 VDDA.t292 0.1368
R1245 VDDA.n465 VDDA.t265 0.1368
R1246 VDDA.n465 VDDA.t309 0.1368
R1247 VDDA.n464 VDDA.t283 0.1368
R1248 VDDA.n464 VDDA.t274 0.1368
R1249 VDDA.t291 VDDA.n464 0.00152174
R1250 VDDA.t273 VDDA.n465 0.00152174
R1251 VDDA.t308 VDDA.n466 0.00152174
R1252 VDDA.t270 VDDA.n467 0.00152174
R1253 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t15 354.854
R1254 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t30 346.8
R1255 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n4 339.522
R1256 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 339.522
R1257 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n9 335.022
R1258 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t0 275.909
R1259 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 227.909
R1260 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 222.034
R1261 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t31 184.097
R1262 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t14 184.097
R1263 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t27 184.097
R1264 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t19 184.097
R1265 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 166.05
R1266 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 166.05
R1267 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t1 48.0005
R1268 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t9 48.0005
R1269 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t10 48.0005
R1270 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t2 48.0005
R1271 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t6 39.4005
R1272 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t4 39.4005
R1273 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t7 39.4005
R1274 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t8 39.4005
R1275 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t5 39.4005
R1276 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t3 39.4005
R1277 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n2 33.1711
R1278 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n0 5.6255
R1279 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 5.28175
R1280 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R1281 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t29 4.8295
R1282 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t25 4.8295
R1283 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t35 4.8295
R1284 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t33 4.8295
R1285 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t17 4.8295
R1286 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t28 4.8295
R1287 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n7 4.5005
R1288 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t11 4.5005
R1289 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t32 4.5005
R1290 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t34 4.5005
R1291 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t21 4.5005
R1292 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t12 4.5005
R1293 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t16 4.5005
R1294 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t26 4.5005
R1295 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t22 4.5005
R1296 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.5005
R1297 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.5005
R1298 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t13 4.5005
R1299 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t18 4.5005
R1300 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t36 4.5005
R1301 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.8075
R1302 bgr_0.cap_res1.t20 bgr_0.cap_res1.t17 178.633
R1303 bgr_0.cap_res1.t14 bgr_0.cap_res1.t0 0.1603
R1304 bgr_0.cap_res1.t10 bgr_0.cap_res1.t6 0.1603
R1305 bgr_0.cap_res1.t9 bgr_0.cap_res1.t15 0.1603
R1306 bgr_0.cap_res1.t7 bgr_0.cap_res1.t3 0.1603
R1307 bgr_0.cap_res1.t16 bgr_0.cap_res1.t1 0.1603
R1308 bgr_0.cap_res1.t12 bgr_0.cap_res1.t8 0.1603
R1309 bgr_0.cap_res1.t2 bgr_0.cap_res1.t5 0.1603
R1310 bgr_0.cap_res1.t19 bgr_0.cap_res1.t13 0.1603
R1311 bgr_0.cap_res1.n1 bgr_0.cap_res1.t4 0.159278
R1312 bgr_0.cap_res1.n2 bgr_0.cap_res1.t18 0.159278
R1313 bgr_0.cap_res1.n3 bgr_0.cap_res1.t11 0.159278
R1314 bgr_0.cap_res1.n3 bgr_0.cap_res1.t14 0.1368
R1315 bgr_0.cap_res1.n3 bgr_0.cap_res1.t10 0.1368
R1316 bgr_0.cap_res1.n2 bgr_0.cap_res1.t9 0.1368
R1317 bgr_0.cap_res1.n2 bgr_0.cap_res1.t7 0.1368
R1318 bgr_0.cap_res1.n1 bgr_0.cap_res1.t16 0.1368
R1319 bgr_0.cap_res1.n1 bgr_0.cap_res1.t12 0.1368
R1320 bgr_0.cap_res1.n0 bgr_0.cap_res1.t2 0.1368
R1321 bgr_0.cap_res1.n0 bgr_0.cap_res1.t19 0.1368
R1322 bgr_0.cap_res1.t4 bgr_0.cap_res1.n0 0.00152174
R1323 bgr_0.cap_res1.t18 bgr_0.cap_res1.n1 0.00152174
R1324 bgr_0.cap_res1.t11 bgr_0.cap_res1.n2 0.00152174
R1325 bgr_0.cap_res1.t17 bgr_0.cap_res1.n3 0.00152174
R1326 a_14710_5068.t0 a_14710_5068.t1 169.905
R1327 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t6 327.092
R1328 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R1329 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R1330 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R1331 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 166.488
R1332 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R1333 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R1334 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R1335 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R1336 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R1337 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R1338 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R1339 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R1340 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R1341 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t1 117.591
R1342 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 117.591
R1343 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t2 108.424
R1344 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 108.424
R1345 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 25.9693
R1346 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n0 25.784
R1347 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 9.90675
R1348 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 1.09425
R1349 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 0.688
R1350 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 0.63175
R1351 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n4 0.61925
R1352 GNDA.n341 GNDA.n340 225584
R1353 GNDA.n1677 GNDA.n1676 40282.1
R1354 GNDA.n342 GNDA.n341 35807.6
R1355 GNDA.n2461 GNDA.n2460 30393.4
R1356 GNDA.n344 GNDA.n343 29285.4
R1357 GNDA.n1608 GNDA.n84 28605.1
R1358 GNDA.n2460 GNDA.n59 28430.8
R1359 GNDA.n344 GNDA.n327 28430.8
R1360 GNDA.n1675 GNDA.n1608 26648.4
R1361 GNDA.n327 GNDA.n80 23523.1
R1362 GNDA.n80 GNDA.n59 23523.1
R1363 GNDA.n1676 GNDA.n83 21360.7
R1364 GNDA.n2441 GNDA.n2440 21106.2
R1365 GNDA.n2442 GNDA.n81 20366.8
R1366 GNDA.n1676 GNDA.n84 19892.9
R1367 GNDA.n2443 GNDA.n80 19630.8
R1368 GNDA.n327 GNDA.n81 17609.2
R1369 GNDA.n2445 GNDA.n59 17609.2
R1370 GNDA.n1679 GNDA.n1675 17265.8
R1371 GNDA.n2443 GNDA.n2442 17092.3
R1372 GNDA.n1677 GNDA.n1675 15892.5
R1373 GNDA.n341 GNDA.n59 14416.4
R1374 GNDA.n1681 GNDA.n1610 12361.8
R1375 GNDA.n1685 GNDA.n1610 12312.5
R1376 GNDA.n1681 GNDA.n1611 11918.5
R1377 GNDA.n1685 GNDA.n1611 11869.2
R1378 GNDA.n2444 GNDA.n2443 11513.6
R1379 GNDA.n464 GNDA.n37 11426
R1380 GNDA.n485 GNDA.n81 11060.7
R1381 GNDA.n453 GNDA.n36 10441
R1382 GNDA.n453 GNDA.n37 10441
R1383 GNDA.n1725 GNDA.n1608 10371.4
R1384 GNDA.n464 GNDA.n36 9456
R1385 GNDA.n2487 GNDA.n29 9259
R1386 GNDA.n1688 GNDA.n1637 9062
R1387 GNDA.n2487 GNDA.n30 8865
R1388 GNDA.n107 GNDA.n103 8175.5
R1389 GNDA.n2425 GNDA.n103 8126.25
R1390 GNDA.n1692 GNDA.n1632 7880
R1391 GNDA.n1692 GNDA.n1633 7880
R1392 GNDA.n1731 GNDA.n1605 7880
R1393 GNDA.n1727 GNDA.n1605 7880
R1394 GNDA.n1635 GNDA.n1632 7830.75
R1395 GNDA.n1635 GNDA.n1633 7830.75
R1396 GNDA.n1731 GNDA.n1606 7830.75
R1397 GNDA.n1727 GNDA.n1606 7830.75
R1398 GNDA.n107 GNDA.n101 7732.25
R1399 GNDA.n450 GNDA.n391 7732.25
R1400 GNDA.n446 GNDA.n391 7732.25
R1401 GNDA.n450 GNDA.n392 7732.25
R1402 GNDA.n446 GNDA.n392 7732.25
R1403 GNDA.n475 GNDA.n345 7732.25
R1404 GNDA.n467 GNDA.n345 7732.25
R1405 GNDA.n475 GNDA.n346 7732.25
R1406 GNDA.n467 GNDA.n346 7732.25
R1407 GNDA.n2425 GNDA.n101 7683
R1408 GNDA.n483 GNDA.n318 6944.25
R1409 GNDA.n2172 GNDA.n314 6845.75
R1410 GNDA.n2176 GNDA.n314 6845.75
R1411 GNDA.n2172 GNDA.n313 6796.5
R1412 GNDA.n2176 GNDA.n313 6796.5
R1413 GNDA.n2447 GNDA.n74 6796.5
R1414 GNDA.n354 GNDA.n318 6722.62
R1415 GNDA.n2170 GNDA.n487 6698
R1416 GNDA.n2165 GNDA.n487 6698
R1417 GNDA.n2170 GNDA.n486 6648.75
R1418 GNDA.n2165 GNDA.n486 6648.75
R1419 GNDA.n437 GNDA.n74 6550.25
R1420 GNDA.n437 GNDA.n75 5614.5
R1421 GNDA.n354 GNDA.n319 5589.88
R1422 GNDA.n2462 GNDA.n56 5319
R1423 GNDA.n336 GNDA.n330 5319
R1424 GNDA.n483 GNDA.n319 5269.75
R1425 GNDA.n2447 GNDA.n75 5269.75
R1426 GNDA.n343 GNDA.n342 5240.28
R1427 GNDA.n371 GNDA.n351 5171.25
R1428 GNDA.n2480 GNDA.n29 5171.25
R1429 GNDA.n2482 GNDA.n30 5171.25
R1430 GNDA.n2459 GNDA.n61 5171.25
R1431 GNDA.n2442 GNDA.n2441 5136.31
R1432 GNDA.n353 GNDA.n351 5122
R1433 GNDA.n2455 GNDA.n61 5122
R1434 GNDA.n1690 GNDA.n1637 4974.25
R1435 GNDA.n1709 GNDA.n1623 4974.25
R1436 GNDA.n1713 GNDA.n1623 4974.25
R1437 GNDA.n371 GNDA.n370 4944.7
R1438 GNDA.n2459 GNDA.n62 4944.7
R1439 GNDA.n2473 GNDA.n38 4925
R1440 GNDA.n2473 GNDA.n39 4925
R1441 GNDA.n370 GNDA.n353 4895.45
R1442 GNDA.n2455 GNDA.n62 4895.45
R1443 GNDA.n38 GNDA.n35 4728
R1444 GNDA.n39 GNDA.n35 4728
R1445 GNDA.n2429 GNDA.n96 4678.75
R1446 GNDA.n2429 GNDA.n95 4629.5
R1447 GNDA.n167 GNDA.n96 4629.5
R1448 GNDA.n2439 GNDA.n84 4603.73
R1449 GNDA.n2151 GNDA.n501 4580.25
R1450 GNDA.n2151 GNDA.n502 4580.25
R1451 GNDA.n167 GNDA.n95 4580.25
R1452 GNDA.n2147 GNDA.n500 4580.25
R1453 GNDA.n510 GNDA.n500 4580.25
R1454 GNDA.n1724 GNDA.n1612 4531
R1455 GNDA.n1724 GNDA.n1613 4531
R1456 GNDA.n1612 GNDA.n1609 4531
R1457 GNDA.n1613 GNDA.n1609 4531
R1458 GNDA.n1709 GNDA.n1622 4531
R1459 GNDA.n1713 GNDA.n1622 4531
R1460 GNDA.n2118 GNDA.n501 4481.75
R1461 GNDA.n2118 GNDA.n502 4481.75
R1462 GNDA.n2147 GNDA.n507 4481.75
R1463 GNDA.n510 GNDA.n507 4481.75
R1464 GNDA.n485 GNDA.n484 4289.57
R1465 GNDA.n429 GNDA.n428 4124.69
R1466 GNDA.n1678 GNDA.n1677 4073.68
R1467 GNDA.n2440 GNDA.n2439 3918.75
R1468 GNDA.n342 GNDA.n327 3758.33
R1469 GNDA.n2480 GNDA.n34 3595.25
R1470 GNDA.n457 GNDA.n326 3373.63
R1471 GNDA.n2490 GNDA.n27 3349
R1472 GNDA.n2476 GNDA.n27 3299.75
R1473 GNDA.n2490 GNDA.n28 3250.5
R1474 GNDA.n1680 GNDA.n1679 3209.7
R1475 GNDA.n2482 GNDA.n34 3201.25
R1476 GNDA.n2476 GNDA.n28 3201.25
R1477 GNDA.n459 GNDA.n326 3176.63
R1478 GNDA.n444 GNDA.n429 2425.56
R1479 GNDA.n359 GNDA.n356 2326.02
R1480 GNDA.n367 GNDA.n356 2326.02
R1481 GNDA.n69 GNDA.n66 2326.02
R1482 GNDA.n77 GNDA.n66 2326.02
R1483 GNDA.n1673 GNDA.n1643 2142.38
R1484 GNDA.n1706 GNDA.n1621 2142.38
R1485 GNDA.n1842 GNDA.n597 1852.75
R1486 GNDA.n1643 GNDA.n1642 1846.88
R1487 GNDA.n1717 GNDA.n1621 1846.88
R1488 GNDA.n1678 GNDA.n79 1755.83
R1489 GNDA.n478 GNDA.n326 1636.08
R1490 GNDA.n435 GNDA.n429 1527.38
R1491 GNDA.n1679 GNDA.n1678 1226.55
R1492 GNDA.n2444 GNDA.n79 1126.93
R1493 GNDA.n364 GNDA.n356 1114.8
R1494 GNDA.n2452 GNDA.n66 1114.8
R1495 GNDA.n343 GNDA.n337 1107.91
R1496 GNDA.n1670 GNDA.n1643 991.841
R1497 GNDA.n1701 GNDA.n1621 991.841
R1498 GNDA.n2171 GNDA.n317 989.183
R1499 GNDA.n83 GNDA.n79 954.963
R1500 GNDA.n741 GNDA.n614 942.497
R1501 GNDA.n1439 GNDA.n587 942.497
R1502 GNDA.n2446 GNDA.n2445 938.855
R1503 GNDA.n2445 GNDA.n2444 924.173
R1504 GNDA.n1421 GNDA.n614 922.337
R1505 GNDA.n1866 GNDA.n587 922.337
R1506 GNDA.n456 GNDA.t273 895.083
R1507 GNDA.n323 GNDA.t255 895.083
R1508 GNDA.n441 GNDA.t258 895.083
R1509 GNDA.n430 GNDA.t245 895.083
R1510 GNDA.n1682 GNDA.n1626 803.201
R1511 GNDA.n1684 GNDA.n1626 800
R1512 GNDA.n1683 GNDA.n1682 774.4
R1513 GNDA.n1684 GNDA.n1683 771.201
R1514 GNDA.n463 GNDA.n455 736
R1515 GNDA.n2464 GNDA.n2463 691.201
R1516 GNDA.n335 GNDA.n53 691.201
R1517 GNDA.n455 GNDA.n454 678.4
R1518 GNDA.n2070 GNDA.n543 669.307
R1519 GNDA.n395 GNDA.t248 666.134
R1520 GNDA.n32 GNDA.t287 666.134
R1521 GNDA.n2056 GNDA.n2055 662.155
R1522 GNDA.n2329 GNDA.n145 662.155
R1523 GNDA.n434 GNDA.n431 624
R1524 GNDA.n366 GNDA.n357 617.601
R1525 GNDA.n71 GNDA.n70 617.601
R1526 GNDA.n2486 GNDA.n31 601.601
R1527 GNDA.n2071 GNDA.n544 585
R1528 GNDA.n2073 GNDA.n2072 585
R1529 GNDA.n2074 GNDA.n2073 585
R1530 GNDA.n556 GNDA.n555 585
R1531 GNDA.n2057 GNDA.n556 585
R1532 GNDA.n2060 GNDA.n2059 585
R1533 GNDA.n2059 GNDA.n2058 585
R1534 GNDA.n2061 GNDA.n554 585
R1535 GNDA.n554 GNDA.n553 585
R1536 GNDA.n2063 GNDA.n2062 585
R1537 GNDA.n2064 GNDA.n2063 585
R1538 GNDA.n552 GNDA.n551 585
R1539 GNDA.n2065 GNDA.n552 585
R1540 GNDA.n2068 GNDA.n2067 585
R1541 GNDA.n2067 GNDA.n2066 585
R1542 GNDA.n542 GNDA.n541 585
R1543 GNDA.n2075 GNDA.n542 585
R1544 GNDA.n2078 GNDA.n2077 585
R1545 GNDA.n2077 GNDA.n2076 585
R1546 GNDA.n2079 GNDA.n540 585
R1547 GNDA.n540 GNDA.n539 585
R1548 GNDA.n2082 GNDA.n2081 585
R1549 GNDA.n2083 GNDA.n2082 585
R1550 GNDA.n2080 GNDA.n536 585
R1551 GNDA.n2084 GNDA.n536 585
R1552 GNDA.n2086 GNDA.n538 585
R1553 GNDA.n2086 GNDA.n2085 585
R1554 GNDA.n893 GNDA.n730 585
R1555 GNDA.n730 GNDA.n729 585
R1556 GNDA.n895 GNDA.n894 585
R1557 GNDA.n896 GNDA.n895 585
R1558 GNDA.n728 GNDA.n727 585
R1559 GNDA.n897 GNDA.n728 585
R1560 GNDA.n901 GNDA.n900 585
R1561 GNDA.n900 GNDA.n899 585
R1562 GNDA.n902 GNDA.n726 585
R1563 GNDA.n898 GNDA.n726 585
R1564 GNDA.n904 GNDA.n903 585
R1565 GNDA.n904 GNDA.n610 585
R1566 GNDA.n905 GNDA.n725 585
R1567 GNDA.n905 GNDA.n611 585
R1568 GNDA.n908 GNDA.n907 585
R1569 GNDA.n907 GNDA.n906 585
R1570 GNDA.n909 GNDA.n724 585
R1571 GNDA.n724 GNDA.n723 585
R1572 GNDA.n912 GNDA.n911 585
R1573 GNDA.n913 GNDA.n912 585
R1574 GNDA.n910 GNDA.n720 585
R1575 GNDA.n914 GNDA.n720 585
R1576 GNDA.n916 GNDA.n722 585
R1577 GNDA.n916 GNDA.n915 585
R1578 GNDA.n917 GNDA.n719 585
R1579 GNDA.n917 GNDA.n557 585
R1580 GNDA.n740 GNDA.n739 585
R1581 GNDA.n873 GNDA.n740 585
R1582 GNDA.n876 GNDA.n875 585
R1583 GNDA.n875 GNDA.n874 585
R1584 GNDA.n877 GNDA.n738 585
R1585 GNDA.n738 GNDA.n737 585
R1586 GNDA.n879 GNDA.n878 585
R1587 GNDA.n880 GNDA.n879 585
R1588 GNDA.n736 GNDA.n735 585
R1589 GNDA.n881 GNDA.n736 585
R1590 GNDA.n884 GNDA.n883 585
R1591 GNDA.n883 GNDA.n882 585
R1592 GNDA.n885 GNDA.n734 585
R1593 GNDA.n734 GNDA.n733 585
R1594 GNDA.n887 GNDA.n886 585
R1595 GNDA.n888 GNDA.n887 585
R1596 GNDA.n732 GNDA.n731 585
R1597 GNDA.n889 GNDA.n732 585
R1598 GNDA.n892 GNDA.n891 585
R1599 GNDA.n891 GNDA.n890 585
R1600 GNDA.n1412 GNDA.n1411 585
R1601 GNDA.n1438 GNDA.n1412 585
R1602 GNDA.n1436 GNDA.n1435 585
R1603 GNDA.n1437 GNDA.n1436 585
R1604 GNDA.n1434 GNDA.n1414 585
R1605 GNDA.n1414 GNDA.n1413 585
R1606 GNDA.n1433 GNDA.n1432 585
R1607 GNDA.n1432 GNDA.n1431 585
R1608 GNDA.n1416 GNDA.n1415 585
R1609 GNDA.n1430 GNDA.n1416 585
R1610 GNDA.n1428 GNDA.n1427 585
R1611 GNDA.n1429 GNDA.n1428 585
R1612 GNDA.n1426 GNDA.n1418 585
R1613 GNDA.n1418 GNDA.n1417 585
R1614 GNDA.n1425 GNDA.n1424 585
R1615 GNDA.n1424 GNDA.n1423 585
R1616 GNDA.n1420 GNDA.n1419 585
R1617 GNDA.n1422 GNDA.n1420 585
R1618 GNDA.n622 GNDA.n621 585
R1619 GNDA.n1421 GNDA.n621 585
R1620 GNDA.n1867 GNDA.n585 585
R1621 GNDA.n1867 GNDA.n1866 585
R1622 GNDA.n590 GNDA.n586 585
R1623 GNDA.n1865 GNDA.n586 585
R1624 GNDA.n1863 GNDA.n1862 585
R1625 GNDA.n1864 GNDA.n1863 585
R1626 GNDA.n1861 GNDA.n589 585
R1627 GNDA.n589 GNDA.n588 585
R1628 GNDA.n1860 GNDA.n1859 585
R1629 GNDA.n1859 GNDA.n1858 585
R1630 GNDA.n592 GNDA.n591 585
R1631 GNDA.n1857 GNDA.n592 585
R1632 GNDA.n1855 GNDA.n1854 585
R1633 GNDA.n1856 GNDA.n1855 585
R1634 GNDA.n1853 GNDA.n594 585
R1635 GNDA.n594 GNDA.n593 585
R1636 GNDA.n1852 GNDA.n1851 585
R1637 GNDA.n1851 GNDA.n1850 585
R1638 GNDA.n596 GNDA.n595 585
R1639 GNDA.n1849 GNDA.n596 585
R1640 GNDA.n1848 GNDA.n1847 585
R1641 GNDA.n598 GNDA.n597 585
R1642 GNDA.n1870 GNDA.n1869 585
R1643 GNDA.n1871 GNDA.n584 585
R1644 GNDA.n1873 GNDA.n1872 585
R1645 GNDA.n1875 GNDA.n583 585
R1646 GNDA.n1878 GNDA.n1877 585
R1647 GNDA.n1879 GNDA.n582 585
R1648 GNDA.n1881 GNDA.n1880 585
R1649 GNDA.n1883 GNDA.n581 585
R1650 GNDA.n1886 GNDA.n1885 585
R1651 GNDA.n1887 GNDA.n580 585
R1652 GNDA.n1889 GNDA.n1888 585
R1653 GNDA.n1891 GNDA.n578 585
R1654 GNDA.n1591 GNDA.n1590 585
R1655 GNDA.n1589 GNDA.n620 585
R1656 GNDA.n1588 GNDA.n1587 585
R1657 GNDA.n1586 GNDA.n1585 585
R1658 GNDA.n1584 GNDA.n1583 585
R1659 GNDA.n1582 GNDA.n1581 585
R1660 GNDA.n1580 GNDA.n1579 585
R1661 GNDA.n1578 GNDA.n1577 585
R1662 GNDA.n1576 GNDA.n1575 585
R1663 GNDA.n1574 GNDA.n1573 585
R1664 GNDA.n1572 GNDA.n1571 585
R1665 GNDA.n1570 GNDA.n1569 585
R1666 GNDA.n948 GNDA.n947 585
R1667 GNDA.n936 GNDA.n709 585
R1668 GNDA.n937 GNDA.n712 585
R1669 GNDA.n940 GNDA.n939 585
R1670 GNDA.n935 GNDA.n714 585
R1671 GNDA.n933 GNDA.n932 585
R1672 GNDA.n716 GNDA.n715 585
R1673 GNDA.n926 GNDA.n925 585
R1674 GNDA.n923 GNDA.n718 585
R1675 GNDA.n921 GNDA.n920 585
R1676 GNDA.n1550 GNDA.n644 585
R1677 GNDA.n1551 GNDA.n642 585
R1678 GNDA.n1552 GNDA.n641 585
R1679 GNDA.n639 GNDA.n637 585
R1680 GNDA.n1558 GNDA.n636 585
R1681 GNDA.n1559 GNDA.n634 585
R1682 GNDA.n1560 GNDA.n633 585
R1683 GNDA.n631 GNDA.n629 585
R1684 GNDA.n1565 GNDA.n628 585
R1685 GNDA.n1566 GNDA.n626 585
R1686 GNDA.n562 GNDA.n559 585
R1687 GNDA.n1922 GNDA.n1921 585
R1688 GNDA.n566 GNDA.n565 585
R1689 GNDA.n1912 GNDA.n568 585
R1690 GNDA.n1914 GNDA.n1913 585
R1691 GNDA.n1909 GNDA.n570 585
R1692 GNDA.n1908 GNDA.n1907 585
R1693 GNDA.n1899 GNDA.n572 585
R1694 GNDA.n1901 GNDA.n1900 585
R1695 GNDA.n1897 GNDA.n574 585
R1696 GNDA.n1896 GNDA.n1895 585
R1697 GNDA.n1896 GNDA.n559 585
R1698 GNDA.n920 GNDA.n919 585
R1699 GNDA.n718 GNDA.n717 585
R1700 GNDA.n927 GNDA.n926 585
R1701 GNDA.n929 GNDA.n716 585
R1702 GNDA.n932 GNDA.n931 585
R1703 GNDA.n714 GNDA.n713 585
R1704 GNDA.n941 GNDA.n940 585
R1705 GNDA.n943 GNDA.n712 585
R1706 GNDA.n944 GNDA.n709 585
R1707 GNDA.n947 GNDA.n946 585
R1708 GNDA.n1568 GNDA.n624 585
R1709 GNDA.n1568 GNDA.n577 585
R1710 GNDA.n1567 GNDA.n1566 585
R1711 GNDA.n1565 GNDA.n1564 585
R1712 GNDA.n1563 GNDA.n629 585
R1713 GNDA.n1561 GNDA.n1560 585
R1714 GNDA.n1559 GNDA.n630 585
R1715 GNDA.n1558 GNDA.n1557 585
R1716 GNDA.n1555 GNDA.n637 585
R1717 GNDA.n1553 GNDA.n1552 585
R1718 GNDA.n1551 GNDA.n638 585
R1719 GNDA.n1550 GNDA.n1549 585
R1720 GNDA.n1892 GNDA.n576 585
R1721 GNDA.n1892 GNDA.n577 585
R1722 GNDA.n1895 GNDA.n1894 585
R1723 GNDA.n574 GNDA.n573 585
R1724 GNDA.n1902 GNDA.n1901 585
R1725 GNDA.n1904 GNDA.n572 585
R1726 GNDA.n1907 GNDA.n1906 585
R1727 GNDA.n570 GNDA.n569 585
R1728 GNDA.n1915 GNDA.n1914 585
R1729 GNDA.n1917 GNDA.n568 585
R1730 GNDA.n1918 GNDA.n566 585
R1731 GNDA.n1921 GNDA.n1920 585
R1732 GNDA.n567 GNDA.n558 585
R1733 GNDA.n1809 GNDA.n558 585
R1734 GNDA.n1210 GNDA.n575 585
R1735 GNDA.n1261 GNDA.n1260 585
R1736 GNDA.n1259 GNDA.n1209 585
R1737 GNDA.n1258 GNDA.n1257 585
R1738 GNDA.n1256 GNDA.n1255 585
R1739 GNDA.n1254 GNDA.n1253 585
R1740 GNDA.n1252 GNDA.n1251 585
R1741 GNDA.n1250 GNDA.n1249 585
R1742 GNDA.n1248 GNDA.n1247 585
R1743 GNDA.n1246 GNDA.n1245 585
R1744 GNDA.n1244 GNDA.n1243 585
R1745 GNDA.n1242 GNDA.n1241 585
R1746 GNDA.n678 GNDA.n677 585
R1747 GNDA.n676 GNDA.n655 585
R1748 GNDA.n675 GNDA.n674 585
R1749 GNDA.n673 GNDA.n672 585
R1750 GNDA.n671 GNDA.n670 585
R1751 GNDA.n669 GNDA.n668 585
R1752 GNDA.n667 GNDA.n666 585
R1753 GNDA.n665 GNDA.n664 585
R1754 GNDA.n663 GNDA.n662 585
R1755 GNDA.n661 GNDA.n660 585
R1756 GNDA.n659 GNDA.n658 585
R1757 GNDA.n657 GNDA.n656 585
R1758 GNDA.n2322 GNDA.n146 585
R1759 GNDA.n1221 GNDA.n148 585
R1760 GNDA.n1222 GNDA.n1219 585
R1761 GNDA.n1225 GNDA.n1218 585
R1762 GNDA.n1226 GNDA.n1217 585
R1763 GNDA.n1229 GNDA.n1216 585
R1764 GNDA.n1230 GNDA.n1215 585
R1765 GNDA.n1233 GNDA.n1214 585
R1766 GNDA.n1234 GNDA.n1213 585
R1767 GNDA.n1237 GNDA.n1212 585
R1768 GNDA.n1238 GNDA.n161 585
R1769 GNDA.n2322 GNDA.n161 585
R1770 GNDA.n1240 GNDA.n1211 585
R1771 GNDA.n1240 GNDA.n187 585
R1772 GNDA.n1239 GNDA.n1238 585
R1773 GNDA.n1237 GNDA.n1236 585
R1774 GNDA.n1235 GNDA.n1234 585
R1775 GNDA.n1233 GNDA.n1232 585
R1776 GNDA.n1231 GNDA.n1230 585
R1777 GNDA.n1229 GNDA.n1228 585
R1778 GNDA.n1227 GNDA.n1226 585
R1779 GNDA.n1225 GNDA.n1224 585
R1780 GNDA.n1223 GNDA.n1222 585
R1781 GNDA.n1221 GNDA.n1220 585
R1782 GNDA.n2291 GNDA.n199 585
R1783 GNDA.n2291 GNDA.n205 585
R1784 GNDA.n1194 GNDA.n1070 585
R1785 GNDA.n1068 GNDA.n1065 585
R1786 GNDA.n1064 GNDA.n1063 585
R1787 GNDA.n1062 GNDA.n1059 585
R1788 GNDA.n1058 GNDA.n1057 585
R1789 GNDA.n1056 GNDA.n1053 585
R1790 GNDA.n1052 GNDA.n1051 585
R1791 GNDA.n1050 GNDA.n1047 585
R1792 GNDA.n1046 GNDA.n534 585
R1793 GNDA.n2090 GNDA.n2089 585
R1794 GNDA.n2087 GNDA.n533 585
R1795 GNDA.n2087 GNDA.n535 585
R1796 GNDA.n2089 GNDA.n2088 585
R1797 GNDA.n1048 GNDA.n534 585
R1798 GNDA.n1050 GNDA.n1049 585
R1799 GNDA.n1054 GNDA.n1051 585
R1800 GNDA.n1056 GNDA.n1055 585
R1801 GNDA.n1060 GNDA.n1057 585
R1802 GNDA.n1062 GNDA.n1061 585
R1803 GNDA.n1066 GNDA.n1063 585
R1804 GNDA.n1068 GNDA.n1067 585
R1805 GNDA.n1070 GNDA.n1069 585
R1806 GNDA.n2091 GNDA.n532 585
R1807 GNDA.n2092 GNDA.n2091 585
R1808 GNDA.n2095 GNDA.n2094 585
R1809 GNDA.n2094 GNDA.n2093 585
R1810 GNDA.n2096 GNDA.n531 585
R1811 GNDA.n531 GNDA.n530 585
R1812 GNDA.n2098 GNDA.n2097 585
R1813 GNDA.n2099 GNDA.n2098 585
R1814 GNDA.n529 GNDA.n528 585
R1815 GNDA.n2100 GNDA.n529 585
R1816 GNDA.n2103 GNDA.n2102 585
R1817 GNDA.n2102 GNDA.n2101 585
R1818 GNDA.n2104 GNDA.n527 585
R1819 GNDA.n527 GNDA.n526 585
R1820 GNDA.n2106 GNDA.n2105 585
R1821 GNDA.n2107 GNDA.n2106 585
R1822 GNDA.n525 GNDA.n524 585
R1823 GNDA.n2108 GNDA.n525 585
R1824 GNDA.n2112 GNDA.n2111 585
R1825 GNDA.n2111 GNDA.n2110 585
R1826 GNDA.n2113 GNDA.n523 585
R1827 GNDA.n2109 GNDA.n523 585
R1828 GNDA.n2115 GNDA.n2114 585
R1829 GNDA.n2115 GNDA.n317 585
R1830 GNDA.n1196 GNDA.n1071 585
R1831 GNDA.n1196 GNDA.n1195 585
R1832 GNDA.n1097 GNDA.n1096 585
R1833 GNDA.n1092 GNDA.n1091 585
R1834 GNDA.n1168 GNDA.n1167 585
R1835 GNDA.n1171 GNDA.n1170 585
R1836 GNDA.n1090 GNDA.n1087 585
R1837 GNDA.n1083 GNDA.n1082 585
R1838 GNDA.n1179 GNDA.n1178 585
R1839 GNDA.n1182 GNDA.n1181 585
R1840 GNDA.n1081 GNDA.n1078 585
R1841 GNDA.n1074 GNDA.n1073 585
R1842 GNDA.n1190 GNDA.n1189 585
R1843 GNDA.n1193 GNDA.n1192 585
R1844 GNDA.n951 GNDA.n559 585
R1845 GNDA.n949 GNDA.n559 585
R1846 GNDA.n1201 GNDA.n1200 585
R1847 GNDA.n1043 GNDA.n686 585
R1848 GNDA.n690 GNDA.n689 585
R1849 GNDA.n967 GNDA.n966 585
R1850 GNDA.n969 GNDA.n968 585
R1851 GNDA.n973 GNDA.n972 585
R1852 GNDA.n971 GNDA.n957 585
R1853 GNDA.n980 GNDA.n979 585
R1854 GNDA.n982 GNDA.n981 585
R1855 GNDA.n986 GNDA.n985 585
R1856 GNDA.n984 GNDA.n955 585
R1857 GNDA.n953 GNDA.n952 585
R1858 GNDA.n1199 GNDA.n687 585
R1859 GNDA.n687 GNDA.n187 585
R1860 GNDA.n2291 GNDA.n193 585
R1861 GNDA.n2291 GNDA.n206 585
R1862 GNDA.n869 GNDA.n741 585
R1863 GNDA.n872 GNDA.n871 585
R1864 GNDA.n773 GNDA.n772 585
R1865 GNDA.n764 GNDA.n763 585
R1866 GNDA.n844 GNDA.n843 585
R1867 GNDA.n847 GNDA.n846 585
R1868 GNDA.n762 GNDA.n759 585
R1869 GNDA.n755 GNDA.n754 585
R1870 GNDA.n855 GNDA.n854 585
R1871 GNDA.n858 GNDA.n857 585
R1872 GNDA.n753 GNDA.n750 585
R1873 GNDA.n746 GNDA.n744 585
R1874 GNDA.n866 GNDA.n865 585
R1875 GNDA.n868 GNDA.n743 585
R1876 GNDA.n771 GNDA.n766 585
R1877 GNDA.n771 GNDA.n577 585
R1878 GNDA.n711 GNDA.n558 585
R1879 GNDA.n770 GNDA.n558 585
R1880 GNDA.n2284 GNDA.n281 585
R1881 GNDA.n279 GNDA.n276 585
R1882 GNDA.n275 GNDA.n274 585
R1883 GNDA.n273 GNDA.n270 585
R1884 GNDA.n269 GNDA.n268 585
R1885 GNDA.n267 GNDA.n264 585
R1886 GNDA.n263 GNDA.n262 585
R1887 GNDA.n261 GNDA.n259 585
R1888 GNDA.n258 GNDA.n184 585
R1889 GNDA.n2295 GNDA.n2294 585
R1890 GNDA.n185 GNDA.n183 585
R1891 GNDA.n187 GNDA.n185 585
R1892 GNDA.n2294 GNDA.n2293 585
R1893 GNDA.n186 GNDA.n184 585
R1894 GNDA.n261 GNDA.n260 585
R1895 GNDA.n265 GNDA.n262 585
R1896 GNDA.n267 GNDA.n266 585
R1897 GNDA.n271 GNDA.n268 585
R1898 GNDA.n273 GNDA.n272 585
R1899 GNDA.n277 GNDA.n274 585
R1900 GNDA.n279 GNDA.n278 585
R1901 GNDA.n281 GNDA.n280 585
R1902 GNDA.n2298 GNDA.n2297 585
R1903 GNDA.n2299 GNDA.n181 585
R1904 GNDA.n2301 GNDA.n2300 585
R1905 GNDA.n2303 GNDA.n180 585
R1906 GNDA.n2306 GNDA.n2305 585
R1907 GNDA.n2307 GNDA.n179 585
R1908 GNDA.n2309 GNDA.n2308 585
R1909 GNDA.n2311 GNDA.n178 585
R1910 GNDA.n2314 GNDA.n2313 585
R1911 GNDA.n2315 GNDA.n177 585
R1912 GNDA.n2317 GNDA.n2316 585
R1913 GNDA.n2319 GNDA.n176 585
R1914 GNDA.n2286 GNDA.n282 585
R1915 GNDA.n2286 GNDA.n2285 585
R1916 GNDA.n649 GNDA.n559 585
R1917 GNDA.n646 GNDA.n559 585
R1918 GNDA.n1288 GNDA.n1287 585
R1919 GNDA.n1284 GNDA.n1283 585
R1920 GNDA.n1359 GNDA.n1358 585
R1921 GNDA.n1362 GNDA.n1361 585
R1922 GNDA.n1282 GNDA.n1279 585
R1923 GNDA.n1275 GNDA.n1274 585
R1924 GNDA.n1370 GNDA.n1369 585
R1925 GNDA.n1373 GNDA.n1372 585
R1926 GNDA.n1273 GNDA.n1270 585
R1927 GNDA.n1266 GNDA.n1265 585
R1928 GNDA.n1381 GNDA.n1380 585
R1929 GNDA.n1384 GNDA.n1383 585
R1930 GNDA.n208 GNDA.n207 585
R1931 GNDA.n207 GNDA.n187 585
R1932 GNDA.n2291 GNDA.n188 585
R1933 GNDA.n2291 GNDA.n2290 585
R1934 GNDA.n1439 GNDA.n1410 585
R1935 GNDA.n1441 GNDA.n1440 585
R1936 GNDA.n1542 GNDA.n1388 585
R1937 GNDA.n1540 GNDA.n1539 585
R1938 GNDA.n1461 GNDA.n1389 585
R1939 GNDA.n1459 GNDA.n1458 585
R1940 GNDA.n1468 GNDA.n1467 585
R1941 GNDA.n1471 GNDA.n1470 585
R1942 GNDA.n1456 GNDA.n1453 585
R1943 GNDA.n1449 GNDA.n1448 585
R1944 GNDA.n1479 GNDA.n1478 585
R1945 GNDA.n1482 GNDA.n1481 585
R1946 GNDA.n1447 GNDA.n1408 585
R1947 GNDA.n1445 GNDA.n1444 585
R1948 GNDA.n1544 GNDA.n1543 585
R1949 GNDA.n1543 GNDA.n577 585
R1950 GNDA.n1547 GNDA.n558 585
R1951 GNDA.n1387 GNDA.n558 585
R1952 GNDA.n2187 GNDA.n2186 585
R1953 GNDA.n303 GNDA.n302 585
R1954 GNDA.n2258 GNDA.n2257 585
R1955 GNDA.n2261 GNDA.n2260 585
R1956 GNDA.n301 GNDA.n298 585
R1957 GNDA.n294 GNDA.n293 585
R1958 GNDA.n2269 GNDA.n2268 585
R1959 GNDA.n2272 GNDA.n2271 585
R1960 GNDA.n292 GNDA.n289 585
R1961 GNDA.n285 GNDA.n284 585
R1962 GNDA.n2280 GNDA.n2279 585
R1963 GNDA.n2283 GNDA.n2282 585
R1964 GNDA.n256 GNDA.n255 585
R1965 GNDA.n253 GNDA.n209 585
R1966 GNDA.n252 GNDA.n251 585
R1967 GNDA.n250 GNDA.n249 585
R1968 GNDA.n248 GNDA.n211 585
R1969 GNDA.n246 GNDA.n245 585
R1970 GNDA.n244 GNDA.n212 585
R1971 GNDA.n243 GNDA.n242 585
R1972 GNDA.n240 GNDA.n213 585
R1973 GNDA.n238 GNDA.n237 585
R1974 GNDA.n236 GNDA.n214 585
R1975 GNDA.n235 GNDA.n234 585
R1976 GNDA.n438 GNDA.n437 585
R1977 GNDA.n437 GNDA.n65 585
R1978 GNDA.n354 GNDA.n322 585
R1979 GNDA.n355 GNDA.n354 585
R1980 GNDA.n1094 GNDA.n514 585
R1981 GNDA.n1094 GNDA.n172 585
R1982 GNDA.n2116 GNDA.n522 585
R1983 GNDA.n2117 GNDA.n2116 585
R1984 GNDA.n2122 GNDA.n2121 585
R1985 GNDA.n2121 GNDA.n2120 585
R1986 GNDA.n2123 GNDA.n521 585
R1987 GNDA.n521 GNDA.n520 585
R1988 GNDA.n2125 GNDA.n2124 585
R1989 GNDA.n2126 GNDA.n2125 585
R1990 GNDA.n519 GNDA.n518 585
R1991 GNDA.n2127 GNDA.n519 585
R1992 GNDA.n2131 GNDA.n2130 585
R1993 GNDA.n2130 GNDA.n2129 585
R1994 GNDA.n2132 GNDA.n517 585
R1995 GNDA.n2128 GNDA.n517 585
R1996 GNDA.n2134 GNDA.n2133 585
R1997 GNDA.n2135 GNDA.n2134 585
R1998 GNDA.n516 GNDA.n515 585
R1999 GNDA.n2136 GNDA.n516 585
R2000 GNDA.n2139 GNDA.n2138 585
R2001 GNDA.n2138 GNDA.n2137 585
R2002 GNDA.n2140 GNDA.n512 585
R2003 GNDA.n512 GNDA.n508 585
R2004 GNDA.n2144 GNDA.n2143 585
R2005 GNDA.n513 GNDA.n511 585
R2006 GNDA.n2185 GNDA.n305 585
R2007 GNDA.n2185 GNDA.n169 585
R2008 GNDA.n2320 GNDA.n174 585
R2009 GNDA.n2321 GNDA.n2320 585
R2010 GNDA.n495 GNDA.n175 585
R2011 GNDA.n175 GNDA.n173 585
R2012 GNDA.n496 GNDA.n494 585
R2013 GNDA.n494 GNDA.n493 585
R2014 GNDA.n498 GNDA.n497 585
R2015 GNDA.n499 GNDA.n498 585
R2016 GNDA.n492 GNDA.n491 585
R2017 GNDA.n2153 GNDA.n492 585
R2018 GNDA.n2157 GNDA.n2156 585
R2019 GNDA.n2156 GNDA.n2155 585
R2020 GNDA.n2158 GNDA.n489 585
R2021 GNDA.n2154 GNDA.n489 585
R2022 GNDA.n2162 GNDA.n2161 585
R2023 GNDA.n2163 GNDA.n2162 585
R2024 GNDA.n2160 GNDA.n490 585
R2025 GNDA.n490 GNDA.n312 585
R2026 GNDA.n2159 GNDA.n309 585
R2027 GNDA.n2178 GNDA.n309 585
R2028 GNDA.n2180 GNDA.n311 585
R2029 GNDA.n2180 GNDA.n2179 585
R2030 GNDA.n2182 GNDA.n2181 585
R2031 GNDA.n2184 GNDA.n2183 585
R2032 GNDA.n2433 GNDA.n2432 585
R2033 GNDA.n2432 GNDA.n2431 585
R2034 GNDA.n232 GNDA.n215 585
R2035 GNDA.n232 GNDA.n216 585
R2036 GNDA.n231 GNDA.n218 585
R2037 GNDA.n231 GNDA.n230 585
R2038 GNDA.n221 GNDA.n217 585
R2039 GNDA.n229 GNDA.n217 585
R2040 GNDA.n227 GNDA.n226 585
R2041 GNDA.n228 GNDA.n227 585
R2042 GNDA.n225 GNDA.n220 585
R2043 GNDA.n220 GNDA.n219 585
R2044 GNDA.n224 GNDA.n223 585
R2045 GNDA.n223 GNDA.n222 585
R2046 GNDA.n115 GNDA.n114 585
R2047 GNDA.n117 GNDA.n115 585
R2048 GNDA.n2418 GNDA.n2417 585
R2049 GNDA.n2417 GNDA.n2416 585
R2050 GNDA.n2419 GNDA.n109 585
R2051 GNDA.n109 GNDA.n104 585
R2052 GNDA.n2422 GNDA.n2421 585
R2053 GNDA.n2423 GNDA.n2422 585
R2054 GNDA.n2420 GNDA.n113 585
R2055 GNDA.n113 GNDA.n108 585
R2056 GNDA.n112 GNDA.n111 585
R2057 GNDA.n93 GNDA.n92 585
R2058 GNDA.n2434 GNDA.n88 585
R2059 GNDA.n88 GNDA.n86 585
R2060 GNDA.n2437 GNDA.n2436 585
R2061 GNDA.n2438 GNDA.n2437 585
R2062 GNDA.n2403 GNDA.n87 585
R2063 GNDA.n87 GNDA.n85 585
R2064 GNDA.n2407 GNDA.n2406 585
R2065 GNDA.n2406 GNDA.n2405 585
R2066 GNDA.n124 GNDA.n122 585
R2067 GNDA.n122 GNDA.n120 585
R2068 GNDA.n2414 GNDA.n2413 585
R2069 GNDA.n2415 GNDA.n2414 585
R2070 GNDA.n2333 GNDA.n121 585
R2071 GNDA.n121 GNDA.n119 585
R2072 GNDA.n2340 GNDA.n2339 585
R2073 GNDA.n2341 GNDA.n2340 585
R2074 GNDA.n2331 GNDA.n144 585
R2075 GNDA.n2342 GNDA.n144 585
R2076 GNDA.n2345 GNDA.n2344 585
R2077 GNDA.n2344 GNDA.n2343 585
R2078 GNDA.n143 GNDA.n141 585
R2079 GNDA.n2330 GNDA.n143 585
R2080 GNDA.n2328 GNDA.n2327 585
R2081 GNDA.n2329 GNDA.n2328 585
R2082 GNDA.n2021 GNDA.n1946 585
R2083 GNDA.n1946 GNDA.n1945 585
R2084 GNDA.n2024 GNDA.n2023 585
R2085 GNDA.n2025 GNDA.n2024 585
R2086 GNDA.n1947 GNDA.n1942 585
R2087 GNDA.n2026 GNDA.n1942 585
R2088 GNDA.n2029 GNDA.n2028 585
R2089 GNDA.n2028 GNDA.n2027 585
R2090 GNDA.n1941 GNDA.n1939 585
R2091 GNDA.n1944 GNDA.n1941 585
R2092 GNDA.n1935 GNDA.n1934 585
R2093 GNDA.n1943 GNDA.n1934 585
R2094 GNDA.n2037 GNDA.n2036 585
R2095 GNDA.n2041 GNDA.n2037 585
R2096 GNDA.n2044 GNDA.n2043 585
R2097 GNDA.n2043 GNDA.n2042 585
R2098 GNDA.n1933 GNDA.n1931 585
R2099 GNDA.n2040 GNDA.n1933 585
R2100 GNDA.n2038 GNDA.n1927 585
R2101 GNDA.n2039 GNDA.n2038 585
R2102 GNDA.n2051 GNDA.n563 585
R2103 GNDA.n563 GNDA.n561 585
R2104 GNDA.n2054 GNDA.n2053 585
R2105 GNDA.n2055 GNDA.n2054 585
R2106 GNDA.n2020 GNDA.n2019 585
R2107 GNDA.n2019 GNDA.n2018 585
R2108 GNDA.n1812 GNDA.n1735 585
R2109 GNDA.n1735 GNDA.n1734 585
R2110 GNDA.n1815 GNDA.n1814 585
R2111 GNDA.n1816 GNDA.n1815 585
R2112 GNDA.n1736 GNDA.n1603 585
R2113 GNDA.n1817 GNDA.n1603 585
R2114 GNDA.n1820 GNDA.n1819 585
R2115 GNDA.n1819 GNDA.n1818 585
R2116 GNDA.n1598 GNDA.n1595 585
R2117 GNDA.n1595 GNDA.n1594 585
R2118 GNDA.n1827 GNDA.n1826 585
R2119 GNDA.n1828 GNDA.n1827 585
R2120 GNDA.n1596 GNDA.n609 585
R2121 GNDA.n1829 GNDA.n609 585
R2122 GNDA.n1832 GNDA.n1831 585
R2123 GNDA.n1831 GNDA.n1830 585
R2124 GNDA.n605 GNDA.n602 585
R2125 GNDA.n602 GNDA.n601 585
R2126 GNDA.n1839 GNDA.n1838 585
R2127 GNDA.n1840 GNDA.n1839 585
R2128 GNDA.n603 GNDA.n600 585
R2129 GNDA.n1841 GNDA.n600 585
R2130 GNDA.n1844 GNDA.n1843 585
R2131 GNDA.n1843 GNDA.n1842 585
R2132 GNDA.n1811 GNDA.n1810 585
R2133 GNDA.n1810 GNDA.n560 585
R2134 GNDA.n890 GNDA.n729 574.797
R2135 GNDA.n337 GNDA.t282 553.957
R2136 GNDA.n2461 GNDA.t279 553.957
R2137 GNDA.n1733 GNDA.n1732 540.783
R2138 GNDA.n374 GNDA.t306 535.191
R2139 GNDA.n347 GNDA.t223 535.191
R2140 GNDA.n425 GNDA.t241 535.191
R2141 GNDA.n393 GNDA.t252 535.191
R2142 GNDA.n106 GNDA.n100 531.201
R2143 GNDA.n2426 GNDA.n100 528
R2144 GNDA.n436 GNDA.n434 524
R2145 GNDA.n1693 GNDA.n1630 512
R2146 GNDA.n1693 GNDA.n1631 512
R2147 GNDA.n1728 GNDA.n1607 512
R2148 GNDA.n1730 GNDA.n1607 512
R2149 GNDA.n1634 GNDA.n1630 508.8
R2150 GNDA.n1634 GNDA.n1631 508.8
R2151 GNDA.n1729 GNDA.n1728 508.8
R2152 GNDA.n1730 GNDA.n1729 508.8
R2153 GNDA.n106 GNDA.n105 499.2
R2154 GNDA.t230 GNDA.n118 496.098
R2155 GNDA.n473 GNDA.n468 496
R2156 GNDA.n449 GNDA.n448 496
R2157 GNDA.n54 GNDA.t261 493.418
R2158 GNDA.n57 GNDA.t278 493.418
R2159 GNDA.n331 GNDA.t291 493.418
R2160 GNDA.n333 GNDA.t281 493.418
R2161 GNDA.n379 GNDA.t300 493.418
R2162 GNDA.n380 GNDA.t217 493.418
R2163 GNDA.n381 GNDA.t231 493.418
R2164 GNDA.n385 GNDA.t284 493.418
R2165 GNDA.n387 GNDA.t297 493.418
R2166 GNDA.n389 GNDA.t310 493.418
R2167 GNDA.n474 GNDA.n473 489.601
R2168 GNDA.n448 GNDA.n447 489.601
R2169 GNDA.n2426 GNDA.n99 486.401
R2170 GNDA.n466 GNDA.n465 463.603
R2171 GNDA.n452 GNDA.n451 463.603
R2172 GNDA.n890 GNDA.n889 453.608
R2173 GNDA.n889 GNDA.n888 453.608
R2174 GNDA.n888 GNDA.n733 453.608
R2175 GNDA.n882 GNDA.n733 453.608
R2176 GNDA.n882 GNDA.n881 453.608
R2177 GNDA.n880 GNDA.n737 453.608
R2178 GNDA.n874 GNDA.n737 453.608
R2179 GNDA.n874 GNDA.n873 453.608
R2180 GNDA.n873 GNDA.n872 453.608
R2181 GNDA.n872 GNDA.n741 453.608
R2182 GNDA.n1422 GNDA.n1421 453.608
R2183 GNDA.n1423 GNDA.n1422 453.608
R2184 GNDA.n1423 GNDA.n1417 453.608
R2185 GNDA.n1429 GNDA.n1417 453.608
R2186 GNDA.n1430 GNDA.n1429 453.608
R2187 GNDA.n1431 GNDA.n1413 453.608
R2188 GNDA.n1437 GNDA.n1413 453.608
R2189 GNDA.n1438 GNDA.n1437 453.608
R2190 GNDA.n1440 GNDA.n1438 453.608
R2191 GNDA.n1440 GNDA.n1439 453.608
R2192 GNDA.n1866 GNDA.n1865 453.608
R2193 GNDA.n1865 GNDA.n1864 453.608
R2194 GNDA.n1864 GNDA.n588 453.608
R2195 GNDA.n1858 GNDA.n588 453.608
R2196 GNDA.n1858 GNDA.n1857 453.608
R2197 GNDA.n1856 GNDA.n593 453.608
R2198 GNDA.n1850 GNDA.n593 453.608
R2199 GNDA.n1850 GNDA.n1849 453.608
R2200 GNDA.n1849 GNDA.n1848 453.608
R2201 GNDA.n1848 GNDA.n597 453.608
R2202 GNDA.n2174 GNDA.n2173 444.8
R2203 GNDA.n2175 GNDA.n2174 444.8
R2204 GNDA.n2175 GNDA.n315 441.601
R2205 GNDA.n2173 GNDA.n316 438.401
R2206 GNDA.n322 GNDA.n321 436.8
R2207 GNDA.n2169 GNDA.n2168 435.2
R2208 GNDA.n2056 GNDA.n560 434.906
R2209 GNDA.n2018 GNDA.n145 434.906
R2210 GNDA.n462 GNDA.n325 428.8
R2211 GNDA.n2169 GNDA.n488 425.601
R2212 GNDA.n479 GNDA.n325 425.601
R2213 GNDA.n438 GNDA.n72 425.601
R2214 GNDA.n2167 GNDA.n2166 422.401
R2215 GNDA.n482 GNDA.n320 422.401
R2216 GNDA.n2485 GNDA.n2484 420.8
R2217 GNDA.n2166 GNDA.n488 419.2
R2218 GNDA.n1644 GNDA.t270 413.084
R2219 GNDA.n1645 GNDA.t267 413.084
R2220 GNDA.n1616 GNDA.t264 413.084
R2221 GNDA.n1614 GNDA.t237 413.084
R2222 GNDA.n1618 GNDA.t294 413.084
R2223 GNDA.n1703 GNDA.t303 413.084
R2224 GNDA.n2449 GNDA.n2448 412.8
R2225 GNDA.n58 GNDA.n55 403.2
R2226 GNDA.n334 GNDA.n332 403.2
R2227 GNDA.n384 GNDA.n383 403.2
R2228 GNDA.n390 GNDA.n388 403.2
R2229 GNDA.n1689 GNDA.n1688 383.118
R2230 GNDA.n587 GNDA.n579 370.214
R2231 GNDA.n1593 GNDA.n614 370.214
R2232 GNDA.n612 GNDA.n587 365.957
R2233 GNDA.n614 GNDA.n613 365.957
R2234 GNDA.n1842 GNDA.n1841 352.627
R2235 GNDA.n1841 GNDA.n1840 352.627
R2236 GNDA.n1840 GNDA.n601 352.627
R2237 GNDA.n1830 GNDA.n601 352.627
R2238 GNDA.n1830 GNDA.n1829 352.627
R2239 GNDA.n1828 GNDA.n1594 352.627
R2240 GNDA.n1818 GNDA.n1594 352.627
R2241 GNDA.n1818 GNDA.n1817 352.627
R2242 GNDA.n1817 GNDA.n1816 352.627
R2243 GNDA.n1734 GNDA.n560 352.627
R2244 GNDA.n2055 GNDA.n561 352.627
R2245 GNDA.n2039 GNDA.n561 352.627
R2246 GNDA.n2040 GNDA.n2039 352.627
R2247 GNDA.n2042 GNDA.n2040 352.627
R2248 GNDA.n2042 GNDA.n2041 352.627
R2249 GNDA.n1944 GNDA.n1943 352.627
R2250 GNDA.n2027 GNDA.n1944 352.627
R2251 GNDA.n2027 GNDA.n2026 352.627
R2252 GNDA.n2026 GNDA.n2025 352.627
R2253 GNDA.n2025 GNDA.n1945 352.627
R2254 GNDA.n2018 GNDA.n1945 352.627
R2255 GNDA.n2330 GNDA.n2329 352.627
R2256 GNDA.n2343 GNDA.n2330 352.627
R2257 GNDA.n2343 GNDA.n2342 352.627
R2258 GNDA.n2342 GNDA.n2341 352.627
R2259 GNDA.n2341 GNDA.n119 352.627
R2260 GNDA.n2415 GNDA.n120 352.627
R2261 GNDA.t338 GNDA.t282 348.202
R2262 GNDA.t94 GNDA.t338 348.202
R2263 GNDA.t57 GNDA.t94 348.202
R2264 GNDA.t91 GNDA.t57 348.202
R2265 GNDA.t98 GNDA.t91 348.202
R2266 GNDA.t55 GNDA.t98 348.202
R2267 GNDA.t110 GNDA.t55 348.202
R2268 GNDA.t163 GNDA.t43 348.202
R2269 GNDA.t65 GNDA.t35 348.202
R2270 GNDA.t58 GNDA.t127 348.202
R2271 GNDA.t337 GNDA.t58 348.202
R2272 GNDA.t109 GNDA.t97 348.202
R2273 GNDA.t97 GNDA.t56 348.202
R2274 GNDA.t56 GNDA.t1 348.202
R2275 GNDA.t1 GNDA.t279 348.202
R2276 GNDA.n1708 GNDA.n1604 344.135
R2277 GNDA.n2405 GNDA.n85 343.452
R2278 GNDA.n2438 GNDA.n86 343.452
R2279 GNDA.n482 GNDA.n481 342.401
R2280 GNDA.n2448 GNDA.n73 342.401
R2281 GNDA.n2484 GNDA.n2483 336
R2282 GNDA.n2479 GNDA.n31 336
R2283 GNDA.n352 GNDA.n349 332.8
R2284 GNDA.n2456 GNDA.n64 332.8
R2285 GNDA.n2470 GNDA.t220 332.75
R2286 GNDA.n40 GNDA.t226 332.75
R2287 GNDA.t339 GNDA.n328 332.375
R2288 GNDA.n329 GNDA.t63 332.375
R2289 GNDA.t41 GNDA.n338 332.375
R2290 GNDA.n339 GNDA.t81 332.375
R2291 GNDA.n340 GNDA.t337 332.375
R2292 GNDA.n1687 GNDA.n1686 331.844
R2293 GNDA.t230 GNDA.n166 172.876
R2294 GNDA.t234 GNDA.n612 327.661
R2295 GNDA.t234 GNDA.n613 327.661
R2296 GNDA.n1264 GNDA.t236 172.876
R2297 GNDA.n1203 GNDA.t236 172.876
R2298 GNDA.t230 GNDA.n170 172.876
R2299 GNDA.n439 GNDA.n73 326.401
R2300 GNDA.t230 GNDA.n171 172.615
R2301 GNDA.t234 GNDA.n579 323.404
R2302 GNDA.t234 GNDA.n1593 323.404
R2303 GNDA.n1263 GNDA.t236 172.615
R2304 GNDA.n680 GNDA.t236 172.615
R2305 GNDA.t230 GNDA.n116 172.615
R2306 GNDA.n1711 GNDA.n1710 323.2
R2307 GNDA.n1690 GNDA.n1689 322.861
R2308 GNDA.n372 GNDA.n350 321.281
R2309 GNDA.n2458 GNDA.n2457 321.281
R2310 GNDA.n352 GNDA.n350 318.08
R2311 GNDA.n2457 GNDA.n2456 318.08
R2312 GNDA.n1712 GNDA.n1711 316.8
R2313 GNDA.n1734 GNDA.n1733 309.529
R2314 GNDA.n2428 GNDA.n2427 304
R2315 GNDA.n2405 GNDA.n118 301.474
R2316 GNDA.n2427 GNDA.n98 300.8
R2317 GNDA.n2428 GNDA.n97 300.8
R2318 GNDA.n373 GNDA.n349 300.8
R2319 GNDA.n2469 GNDA.n2468 300.8
R2320 GNDA.n2468 GNDA.n42 300.8
R2321 GNDA.n468 GNDA.n377 300.8
R2322 GNDA.n449 GNDA.n394 300.8
R2323 GNDA.n64 GNDA.n63 300.8
R2324 GNDA.n2150 GNDA.n503 297.601
R2325 GNDA.n2150 GNDA.n2149 297.601
R2326 GNDA.n98 GNDA.n97 297.601
R2327 GNDA.n2148 GNDA.n506 297.601
R2328 GNDA.n509 GNDA.n506 297.601
R2329 GNDA.n366 GNDA.n365 296
R2330 GNDA.n2451 GNDA.n70 296
R2331 GNDA.n1721 GNDA.n1720 294.401
R2332 GNDA.n1720 GNDA.n1719 294.401
R2333 GNDA.n1710 GNDA.n1624 294.401
R2334 GNDA.n474 GNDA.n348 294.401
R2335 GNDA.n447 GNDA.n426 294.401
R2336 GNDA.n2456 GNDA.n2455 292.5
R2337 GNDA.n2455 GNDA.n2454 292.5
R2338 GNDA.n2457 GNDA.n62 292.5
R2339 GNDA.n67 GNDA.n62 292.5
R2340 GNDA.n64 GNDA.n61 292.5
R2341 GNDA.n67 GNDA.n61 292.5
R2342 GNDA.n2448 GNDA.n2447 292.5
R2343 GNDA.n2447 GNDA.n2446 292.5
R2344 GNDA.n75 GNDA.n73 292.5
R2345 GNDA.n76 GNDA.n75 292.5
R2346 GNDA.n74 GNDA.n72 292.5
R2347 GNDA.n76 GNDA.n74 292.5
R2348 GNDA.n2452 GNDA.n2451 292.5
R2349 GNDA.n2453 GNDA.n2452 292.5
R2350 GNDA.n330 GNDA.n53 292.5
R2351 GNDA.n330 GNDA.n329 292.5
R2352 GNDA.n336 GNDA.n335 292.5
R2353 GNDA.n337 GNDA.n336 292.5
R2354 GNDA.n2463 GNDA.n2462 292.5
R2355 GNDA.n2462 GNDA.n2461 292.5
R2356 GNDA.n2464 GNDA.n56 292.5
R2357 GNDA.n338 GNDA.n56 292.5
R2358 GNDA.n2469 GNDA.n39 292.5
R2359 GNDA.n339 GNDA.n39 292.5
R2360 GNDA.n2468 GNDA.n35 292.5
R2361 GNDA.n2474 GNDA.n35 292.5
R2362 GNDA.n42 GNDA.n38 292.5
R2363 GNDA.n328 GNDA.n38 292.5
R2364 GNDA.n2473 GNDA.n2472 292.5
R2365 GNDA.n2474 GNDA.n2473 292.5
R2366 GNDA.n2491 GNDA.n2490 292.5
R2367 GNDA.n2490 GNDA.n2489 292.5
R2368 GNDA.n28 GNDA.n25 292.5
R2369 GNDA.n2474 GNDA.n28 292.5
R2370 GNDA.n2476 GNDA.n2475 292.5
R2371 GNDA.n2477 GNDA.n2476 292.5
R2372 GNDA.n27 GNDA.n26 292.5
R2373 GNDA.n2474 GNDA.n27 292.5
R2374 GNDA.n2487 GNDA.n2486 292.5
R2375 GNDA.n2488 GNDA.n2487 292.5
R2376 GNDA.n2484 GNDA.n30 292.5
R2377 GNDA.n2474 GNDA.n30 292.5
R2378 GNDA.n2483 GNDA.n2482 292.5
R2379 GNDA.n2482 GNDA.n2481 292.5
R2380 GNDA.n2478 GNDA.n34 292.5
R2381 GNDA.n378 GNDA.n34 292.5
R2382 GNDA.n2480 GNDA.n2479 292.5
R2383 GNDA.n2481 GNDA.n2480 292.5
R2384 GNDA.n31 GNDA.n29 292.5
R2385 GNDA.n2474 GNDA.n29 292.5
R2386 GNDA.n468 GNDA.n467 292.5
R2387 GNDA.n467 GNDA.n466 292.5
R2388 GNDA.n473 GNDA.n346 292.5
R2389 GNDA.n458 GNDA.n346 292.5
R2390 GNDA.n475 GNDA.n474 292.5
R2391 GNDA.n476 GNDA.n475 292.5
R2392 GNDA.n376 GNDA.n345 292.5
R2393 GNDA.n458 GNDA.n345 292.5
R2394 GNDA.n2459 GNDA.n2458 292.5
R2395 GNDA.n2460 GNDA.n2459 292.5
R2396 GNDA.n447 GNDA.n446 292.5
R2397 GNDA.n446 GNDA.n445 292.5
R2398 GNDA.n448 GNDA.n392 292.5
R2399 GNDA.n427 GNDA.n392 292.5
R2400 GNDA.n450 GNDA.n449 292.5
R2401 GNDA.n451 GNDA.n450 292.5
R2402 GNDA.n432 GNDA.n391 292.5
R2403 GNDA.n427 GNDA.n391 292.5
R2404 GNDA.n454 GNDA.n453 292.5
R2405 GNDA.n453 GNDA.n452 292.5
R2406 GNDA.n455 GNDA.n37 292.5
R2407 GNDA.n2474 GNDA.n37 292.5
R2408 GNDA.n464 GNDA.n463 292.5
R2409 GNDA.n465 GNDA.n464 292.5
R2410 GNDA.n52 GNDA.n36 292.5
R2411 GNDA.n2474 GNDA.n36 292.5
R2412 GNDA.n457 GNDA.n325 292.5
R2413 GNDA.t130 GNDA.n457 292.5
R2414 GNDA.n479 GNDA.n478 292.5
R2415 GNDA.n478 GNDA.n477 292.5
R2416 GNDA.n460 GNDA.n459 292.5
R2417 GNDA.n459 GNDA.t130 292.5
R2418 GNDA.n436 GNDA.n435 292.5
R2419 GNDA.n435 GNDA.n60 292.5
R2420 GNDA.n434 GNDA.n428 292.5
R2421 GNDA.t31 GNDA.n428 292.5
R2422 GNDA.n444 GNDA.n443 292.5
R2423 GNDA.t31 GNDA.n444 292.5
R2424 GNDA.n372 GNDA.n371 292.5
R2425 GNDA.n371 GNDA.n344 292.5
R2426 GNDA.n370 GNDA.n350 292.5
R2427 GNDA.n370 GNDA.n369 292.5
R2428 GNDA.n353 GNDA.n352 292.5
R2429 GNDA.n362 GNDA.n353 292.5
R2430 GNDA.n351 GNDA.n349 292.5
R2431 GNDA.n369 GNDA.n351 292.5
R2432 GNDA.n481 GNDA.n319 292.5
R2433 GNDA.n361 GNDA.n319 292.5
R2434 GNDA.n483 GNDA.n482 292.5
R2435 GNDA.n484 GNDA.n483 292.5
R2436 GNDA.n321 GNDA.n318 292.5
R2437 GNDA.n361 GNDA.n318 292.5
R2438 GNDA.n365 GNDA.n364 292.5
R2439 GNDA.n364 GNDA.n363 292.5
R2440 GNDA.n2176 GNDA.n2175 292.5
R2441 GNDA.n2177 GNDA.n2176 292.5
R2442 GNDA.n2174 GNDA.n314 292.5
R2443 GNDA.n2145 GNDA.n314 292.5
R2444 GNDA.n2173 GNDA.n2172 292.5
R2445 GNDA.n2172 GNDA.n2171 292.5
R2446 GNDA.n315 GNDA.n313 292.5
R2447 GNDA.n2145 GNDA.n313 292.5
R2448 GNDA.n2166 GNDA.n2165 292.5
R2449 GNDA.n2165 GNDA.n2164 292.5
R2450 GNDA.n2168 GNDA.n487 292.5
R2451 GNDA.n2146 GNDA.n487 292.5
R2452 GNDA.n2170 GNDA.n2169 292.5
R2453 GNDA.n2171 GNDA.n2170 292.5
R2454 GNDA.n488 GNDA.n486 292.5
R2455 GNDA.n2146 GNDA.n486 292.5
R2456 GNDA.n103 GNDA.n100 292.5
R2457 GNDA.n103 GNDA.n102 292.5
R2458 GNDA.n107 GNDA.n106 292.5
R2459 GNDA.n2424 GNDA.n107 292.5
R2460 GNDA.n105 GNDA.n101 292.5
R2461 GNDA.n308 GNDA.n101 292.5
R2462 GNDA.n2426 GNDA.n2425 292.5
R2463 GNDA.n2425 GNDA.n2424 292.5
R2464 GNDA.n506 GNDA.n500 292.5
R2465 GNDA.n2152 GNDA.n500 292.5
R2466 GNDA.n510 GNDA.n509 292.5
R2467 GNDA.n2146 GNDA.n510 292.5
R2468 GNDA.n507 GNDA.n505 292.5
R2469 GNDA.n2119 GNDA.n507 292.5
R2470 GNDA.n2148 GNDA.n2147 292.5
R2471 GNDA.n2147 GNDA.n2146 292.5
R2472 GNDA.n2429 GNDA.n2428 292.5
R2473 GNDA.n2430 GNDA.n2429 292.5
R2474 GNDA.n2427 GNDA.n96 292.5
R2475 GNDA.n2424 GNDA.n96 292.5
R2476 GNDA.n167 GNDA.n98 292.5
R2477 GNDA.n168 GNDA.n167 292.5
R2478 GNDA.n97 GNDA.n95 292.5
R2479 GNDA.n2424 GNDA.n95 292.5
R2480 GNDA.n2151 GNDA.n2150 292.5
R2481 GNDA.n2152 GNDA.n2151 292.5
R2482 GNDA.n2149 GNDA.n502 292.5
R2483 GNDA.n2146 GNDA.n502 292.5
R2484 GNDA.n2118 GNDA.n504 292.5
R2485 GNDA.n2119 GNDA.n2118 292.5
R2486 GNDA.n503 GNDA.n501 292.5
R2487 GNDA.n2146 GNDA.n501 292.5
R2488 GNDA.n1713 GNDA.n1712 292.5
R2489 GNDA.n1714 GNDA.n1713 292.5
R2490 GNDA.n1711 GNDA.n1623 292.5
R2491 GNDA.n1700 GNDA.n1623 292.5
R2492 GNDA.n1710 GNDA.n1709 292.5
R2493 GNDA.n1709 GNDA.n1708 292.5
R2494 GNDA.n1624 GNDA.n1622 292.5
R2495 GNDA.n1700 GNDA.n1622 292.5
R2496 GNDA.n1688 GNDA.n1687 292.5
R2497 GNDA.n1691 GNDA.n1690 292.5
R2498 GNDA.n1637 GNDA.n1625 292.5
R2499 GNDA.n1639 GNDA.n1637 292.5
R2500 GNDA.n1633 GNDA.n1631 292.5
R2501 GNDA.n1680 GNDA.n1633 292.5
R2502 GNDA.n1635 GNDA.n1634 292.5
R2503 GNDA.n1691 GNDA.n1635 292.5
R2504 GNDA.n1632 GNDA.n1630 292.5
R2505 GNDA.n1638 GNDA.n1632 292.5
R2506 GNDA.n1693 GNDA.n1692 292.5
R2507 GNDA.n1692 GNDA.n1691 292.5
R2508 GNDA.n1685 GNDA.n1684 292.5
R2509 GNDA.n1686 GNDA.n1685 292.5
R2510 GNDA.n1626 GNDA.n1610 292.5
R2511 GNDA.n1725 GNDA.n1610 292.5
R2512 GNDA.n1682 GNDA.n1681 292.5
R2513 GNDA.n1681 GNDA.n1604 292.5
R2514 GNDA.n1683 GNDA.n1611 292.5
R2515 GNDA.n1725 GNDA.n1611 292.5
R2516 GNDA.n1718 GNDA.n1717 292.5
R2517 GNDA.n1717 GNDA.n1716 292.5
R2518 GNDA.n1701 GNDA.n1620 292.5
R2519 GNDA.n1702 GNDA.n1701 292.5
R2520 GNDA.n1706 GNDA.n1705 292.5
R2521 GNDA.n1707 GNDA.n1706 292.5
R2522 GNDA.n1721 GNDA.n1613 292.5
R2523 GNDA.n1640 GNDA.n1613 292.5
R2524 GNDA.n1720 GNDA.n1609 292.5
R2525 GNDA.n1725 GNDA.n1609 292.5
R2526 GNDA.n1719 GNDA.n1612 292.5
R2527 GNDA.n1715 GNDA.n1612 292.5
R2528 GNDA.n1724 GNDA.n1723 292.5
R2529 GNDA.n1725 GNDA.n1724 292.5
R2530 GNDA.n1673 GNDA.n1672 292.5
R2531 GNDA.n1674 GNDA.n1673 292.5
R2532 GNDA.n1671 GNDA.n1670 292.5
R2533 GNDA.n1670 GNDA.n1636 292.5
R2534 GNDA.n1642 GNDA.n1617 292.5
R2535 GNDA.n1642 GNDA.n1641 292.5
R2536 GNDA.n1728 GNDA.n1727 292.5
R2537 GNDA.n1727 GNDA.n1726 292.5
R2538 GNDA.n1729 GNDA.n1606 292.5
R2539 GNDA.n1700 GNDA.n1606 292.5
R2540 GNDA.n1731 GNDA.n1730 292.5
R2541 GNDA.n1732 GNDA.n1731 292.5
R2542 GNDA.n1607 GNDA.n1605 292.5
R2543 GNDA.n1700 GNDA.n1605 292.5
R2544 GNDA.n504 GNDA.n503 291.2
R2545 GNDA.n2149 GNDA.n504 291.2
R2546 GNDA.n2148 GNDA.n505 291.2
R2547 GNDA.n509 GNDA.n505 291.2
R2548 GNDA.n1712 GNDA.n1624 288
R2549 GNDA.n1647 GNDA.n1646 281.601
R2550 GNDA.n1704 GNDA.n1619 281.601
R2551 GNDA.n1672 GNDA.n1671 278.401
R2552 GNDA.n1705 GNDA.n1620 278.401
R2553 GNDA.n2282 GNDA.n282 259.416
R2554 GNDA.n2328 GNDA.n146 259.416
R2555 GNDA.n2054 GNDA.n562 259.416
R2556 GNDA.n1383 GNDA.n649 259.416
R2557 GNDA.n1843 GNDA.n598 259.416
R2558 GNDA.n1445 GNDA.n1410 259.416
R2559 GNDA.n869 GNDA.n868 259.416
R2560 GNDA.n952 GNDA.n951 259.416
R2561 GNDA.n1192 GNDA.n1071 259.416
R2562 GNDA.n2470 GNDA.t222 258.601
R2563 GNDA.n40 GNDA.t228 258.601
R2564 GNDA.n1686 GNDA.n1680 258.101
R2565 GNDA.n1846 GNDA.n1845 254.494
R2566 GNDA.n870 GNDA.n742 254.392
R2567 GNDA.n1443 GNDA.n1442 254.392
R2568 GNDA.n1868 GNDA.n579 254.34
R2569 GNDA.n1874 GNDA.n579 254.34
R2570 GNDA.n1876 GNDA.n579 254.34
R2571 GNDA.n1882 GNDA.n579 254.34
R2572 GNDA.n1884 GNDA.n579 254.34
R2573 GNDA.n1890 GNDA.n579 254.34
R2574 GNDA.n1593 GNDA.n1592 254.34
R2575 GNDA.n1593 GNDA.n619 254.34
R2576 GNDA.n1593 GNDA.n618 254.34
R2577 GNDA.n1593 GNDA.n617 254.34
R2578 GNDA.n1593 GNDA.n616 254.34
R2579 GNDA.n1593 GNDA.n615 254.34
R2580 GNDA.n708 GNDA.n559 254.34
R2581 GNDA.n938 GNDA.n559 254.34
R2582 GNDA.n934 GNDA.n559 254.34
R2583 GNDA.n924 GNDA.n559 254.34
R2584 GNDA.n922 GNDA.n559 254.34
R2585 GNDA.n643 GNDA.n559 254.34
R2586 GNDA.n640 GNDA.n559 254.34
R2587 GNDA.n635 GNDA.n559 254.34
R2588 GNDA.n632 GNDA.n559 254.34
R2589 GNDA.n627 GNDA.n559 254.34
R2590 GNDA.n1925 GNDA.n1924 254.34
R2591 GNDA.n1923 GNDA.n559 254.34
R2592 GNDA.n1911 GNDA.n559 254.34
R2593 GNDA.n1910 GNDA.n559 254.34
R2594 GNDA.n571 GNDA.n559 254.34
R2595 GNDA.n1898 GNDA.n559 254.34
R2596 GNDA.n918 GNDA.n558 254.34
R2597 GNDA.n928 GNDA.n558 254.34
R2598 GNDA.n930 GNDA.n558 254.34
R2599 GNDA.n942 GNDA.n558 254.34
R2600 GNDA.n945 GNDA.n558 254.34
R2601 GNDA.n625 GNDA.n558 254.34
R2602 GNDA.n1562 GNDA.n558 254.34
R2603 GNDA.n1556 GNDA.n558 254.34
R2604 GNDA.n1554 GNDA.n558 254.34
R2605 GNDA.n1548 GNDA.n558 254.34
R2606 GNDA.n1893 GNDA.n558 254.34
R2607 GNDA.n1903 GNDA.n558 254.34
R2608 GNDA.n1905 GNDA.n558 254.34
R2609 GNDA.n1916 GNDA.n558 254.34
R2610 GNDA.n1919 GNDA.n558 254.34
R2611 GNDA.n1808 GNDA.n1807 254.34
R2612 GNDA.n1263 GNDA.n1262 254.34
R2613 GNDA.n1263 GNDA.n1208 254.34
R2614 GNDA.n1263 GNDA.n1207 254.34
R2615 GNDA.n1263 GNDA.n1206 254.34
R2616 GNDA.n1263 GNDA.n1205 254.34
R2617 GNDA.n1263 GNDA.n1204 254.34
R2618 GNDA.n680 GNDA.n679 254.34
R2619 GNDA.n680 GNDA.n654 254.34
R2620 GNDA.n680 GNDA.n653 254.34
R2621 GNDA.n680 GNDA.n652 254.34
R2622 GNDA.n680 GNDA.n651 254.34
R2623 GNDA.n680 GNDA.n650 254.34
R2624 GNDA.n2325 GNDA.n2324 254.34
R2625 GNDA.n2323 GNDA.n2322 254.34
R2626 GNDA.n2322 GNDA.n165 254.34
R2627 GNDA.n2322 GNDA.n164 254.34
R2628 GNDA.n2322 GNDA.n163 254.34
R2629 GNDA.n2322 GNDA.n162 254.34
R2630 GNDA.n2291 GNDA.n204 254.34
R2631 GNDA.n2291 GNDA.n203 254.34
R2632 GNDA.n2291 GNDA.n202 254.34
R2633 GNDA.n2291 GNDA.n201 254.34
R2634 GNDA.n2291 GNDA.n200 254.34
R2635 GNDA.n2017 GNDA.n2016 254.34
R2636 GNDA.n2322 GNDA.n160 254.34
R2637 GNDA.n2322 GNDA.n159 254.34
R2638 GNDA.n2322 GNDA.n158 254.34
R2639 GNDA.n2322 GNDA.n157 254.34
R2640 GNDA.n2322 GNDA.n156 254.34
R2641 GNDA.n2291 GNDA.n198 254.34
R2642 GNDA.n2291 GNDA.n197 254.34
R2643 GNDA.n2291 GNDA.n196 254.34
R2644 GNDA.n2291 GNDA.n195 254.34
R2645 GNDA.n2291 GNDA.n194 254.34
R2646 GNDA.n2322 GNDA.n155 254.34
R2647 GNDA.n1095 GNDA.n166 254.34
R2648 GNDA.n1169 GNDA.n166 254.34
R2649 GNDA.n1089 GNDA.n166 254.34
R2650 GNDA.n1180 GNDA.n166 254.34
R2651 GNDA.n1080 GNDA.n166 254.34
R2652 GNDA.n1191 GNDA.n166 254.34
R2653 GNDA.n950 GNDA.n707 254.34
R2654 GNDA.n1203 GNDA.n1202 254.34
R2655 GNDA.n1203 GNDA.n685 254.34
R2656 GNDA.n1203 GNDA.n684 254.34
R2657 GNDA.n1203 GNDA.n683 254.34
R2658 GNDA.n1203 GNDA.n682 254.34
R2659 GNDA.n1203 GNDA.n681 254.34
R2660 GNDA.n1198 GNDA.n1045 254.34
R2661 GNDA.n767 GNDA.n613 254.34
R2662 GNDA.n845 GNDA.n613 254.34
R2663 GNDA.n761 GNDA.n613 254.34
R2664 GNDA.n856 GNDA.n613 254.34
R2665 GNDA.n752 GNDA.n613 254.34
R2666 GNDA.n867 GNDA.n613 254.34
R2667 GNDA.n769 GNDA.n768 254.34
R2668 GNDA.n2322 GNDA.n154 254.34
R2669 GNDA.n2322 GNDA.n153 254.34
R2670 GNDA.n2322 GNDA.n152 254.34
R2671 GNDA.n2322 GNDA.n151 254.34
R2672 GNDA.n2322 GNDA.n150 254.34
R2673 GNDA.n2292 GNDA.n2291 254.34
R2674 GNDA.n2291 GNDA.n192 254.34
R2675 GNDA.n2291 GNDA.n191 254.34
R2676 GNDA.n2291 GNDA.n190 254.34
R2677 GNDA.n2291 GNDA.n189 254.34
R2678 GNDA.n2296 GNDA.n171 254.34
R2679 GNDA.n2302 GNDA.n171 254.34
R2680 GNDA.n2304 GNDA.n171 254.34
R2681 GNDA.n2310 GNDA.n171 254.34
R2682 GNDA.n2312 GNDA.n171 254.34
R2683 GNDA.n2318 GNDA.n171 254.34
R2684 GNDA.n2322 GNDA.n149 254.34
R2685 GNDA.n1385 GNDA.n647 254.34
R2686 GNDA.n1286 GNDA.n1264 254.34
R2687 GNDA.n1360 GNDA.n1264 254.34
R2688 GNDA.n1281 GNDA.n1264 254.34
R2689 GNDA.n1371 GNDA.n1264 254.34
R2690 GNDA.n1272 GNDA.n1264 254.34
R2691 GNDA.n1382 GNDA.n1264 254.34
R2692 GNDA.n2289 GNDA.n2288 254.34
R2693 GNDA.n1541 GNDA.n612 254.34
R2694 GNDA.n1457 GNDA.n612 254.34
R2695 GNDA.n1469 GNDA.n612 254.34
R2696 GNDA.n1455 GNDA.n612 254.34
R2697 GNDA.n1480 GNDA.n612 254.34
R2698 GNDA.n1446 GNDA.n612 254.34
R2699 GNDA.n1546 GNDA.n1545 254.34
R2700 GNDA.n306 GNDA.n170 254.34
R2701 GNDA.n2259 GNDA.n170 254.34
R2702 GNDA.n300 GNDA.n170 254.34
R2703 GNDA.n2270 GNDA.n170 254.34
R2704 GNDA.n291 GNDA.n170 254.34
R2705 GNDA.n2281 GNDA.n170 254.34
R2706 GNDA.n254 GNDA.n116 254.34
R2707 GNDA.n210 GNDA.n116 254.34
R2708 GNDA.n247 GNDA.n116 254.34
R2709 GNDA.n241 GNDA.n116 254.34
R2710 GNDA.n239 GNDA.n116 254.34
R2711 GNDA.n233 GNDA.n116 254.34
R2712 GNDA.n2142 GNDA.n2141 254.34
R2713 GNDA.n310 GNDA.n307 254.34
R2714 GNDA.n110 GNDA.n91 254.34
R2715 GNDA.n2074 GNDA.n543 250.349
R2716 GNDA.n2297 GNDA.n2295 249.663
R2717 GNDA.n255 GNDA.n161 249.663
R2718 GNDA.n1896 GNDA.n575 249.663
R2719 GNDA.n678 GNDA.n626 249.663
R2720 GNDA.n1869 GNDA.n1867 249.663
R2721 GNDA.n1591 GNDA.n621 249.663
R2722 GNDA.n891 GNDA.n730 249.663
R2723 GNDA.n921 GNDA.n556 249.663
R2724 GNDA.n2091 GNDA.n2090 249.663
R2725 GNDA.n2439 GNDA.n2438 248.049
R2726 GNDA.n1732 GNDA.n1604 245.81
R2727 GNDA.n2440 GNDA.n83 243.252
R2728 GNDA.n1671 GNDA.n1617 240
R2729 GNDA.n1718 GNDA.n1620 240
R2730 GNDA.n1829 GNDA.t234 239.004
R2731 GNDA.n2041 GNDA.t236 239.004
R2732 GNDA.t230 GNDA.n119 239.004
R2733 GNDA.n881 GNDA.t234 236.885
R2734 GNDA.t234 GNDA.n1430 236.885
R2735 GNDA.n1857 GNDA.t234 236.885
R2736 GNDA.n2479 GNDA.n2478 233.601
R2737 GNDA.n358 GNDA.n357 228.8
R2738 GNDA.n2450 GNDA.n71 228.8
R2739 GNDA.n481 GNDA.n480 227.201
R2740 GNDA.n374 GNDA.t308 224.525
R2741 GNDA.n347 GNDA.t225 224.525
R2742 GNDA.n425 GNDA.t243 224.525
R2743 GNDA.n393 GNDA.t254 224.525
R2744 GNDA.n48 GNDA.n46 222.611
R2745 GNDA.n45 GNDA.n43 222.611
R2746 GNDA.n48 GNDA.n47 222.268
R2747 GNDA.n45 GNDA.n44 222.268
R2748 GNDA.n1522 GNDA.n1397 221.667
R2749 GNDA.n1339 GNDA.n1338 221.667
R2750 GNDA.n2238 GNDA.n2237 221.667
R2751 GNDA.n824 GNDA.n823 221.667
R2752 GNDA.n1024 GNDA.n1023 221.667
R2753 GNDA.n1148 GNDA.n1147 221.667
R2754 GNDA.n1791 GNDA.n1745 221.667
R2755 GNDA.n2000 GNDA.n1956 221.667
R2756 GNDA.n2383 GNDA.n2382 221.667
R2757 GNDA.t227 GNDA.t339 221.583
R2758 GNDA.t67 GNDA.t80 221.583
R2759 GNDA.t39 GNDA.t106 221.583
R2760 GNDA.t63 GNDA.t292 221.583
R2761 GNDA.t262 GNDA.t41 221.583
R2762 GNDA.t105 GNDA.t77 221.583
R2763 GNDA.t18 GNDA.t37 221.583
R2764 GNDA.t81 GNDA.t221 221.583
R2765 GNDA.n51 GNDA.n50 217.768
R2766 GNDA.n2491 GNDA.n26 217.601
R2767 GNDA.t234 GNDA.n880 216.725
R2768 GNDA.n1431 GNDA.t234 216.725
R2769 GNDA.t234 GNDA.n1856 216.725
R2770 GNDA.n2475 GNDA.n26 214.4
R2771 GNDA.n2475 GNDA.n25 203.201
R2772 GNDA.n2492 GNDA.n2491 201.601
R2773 GNDA.n2472 GNDA.n41 201.601
R2774 GNDA.n2472 GNDA.n2471 201.601
R2775 GNDA.n460 GNDA.n324 201.601
R2776 GNDA.n461 GNDA.n460 201.601
R2777 GNDA.n443 GNDA.n431 201.601
R2778 GNDA.n443 GNDA.n442 201.601
R2779 GNDA.n15 GNDA.n13 201.566
R2780 GNDA.n4 GNDA.n2 201.566
R2781 GNDA.n23 GNDA.n22 201.222
R2782 GNDA.n21 GNDA.n20 201.222
R2783 GNDA.n19 GNDA.n18 201.222
R2784 GNDA.n17 GNDA.n16 201.222
R2785 GNDA.n15 GNDA.n14 201.222
R2786 GNDA.n4 GNDA.n3 201.222
R2787 GNDA.n6 GNDA.n5 201.222
R2788 GNDA.n8 GNDA.n7 201.222
R2789 GNDA.n10 GNDA.n9 201.222
R2790 GNDA.n12 GNDA.n11 201.222
R2791 GNDA.n2431 GNDA.n2430 199.727
R2792 GNDA.n2185 GNDA.n2184 197
R2793 GNDA.n2432 GNDA.n92 197
R2794 GNDA.n2019 GNDA.n205 197
R2795 GNDA.n2290 GNDA.n207 197
R2796 GNDA.n1810 GNDA.n1809 197
R2797 GNDA.n1543 GNDA.n1387 197
R2798 GNDA.n771 GNDA.n770 197
R2799 GNDA.n687 GNDA.n206 197
R2800 GNDA.n2073 GNDA.n544 197
R2801 GNDA.n1094 GNDA.n513 197
R2802 GNDA.n77 GNDA.n71 195
R2803 GNDA.n78 GNDA.n77 195
R2804 GNDA.n70 GNDA.n69 195
R2805 GNDA.n69 GNDA.n68 195
R2806 GNDA.n367 GNDA.n366 195
R2807 GNDA.n368 GNDA.n367 195
R2808 GNDA.n359 GNDA.n357 195
R2809 GNDA.n360 GNDA.n359 195
R2810 GNDA.n2320 GNDA.n175 187.249
R2811 GNDA.n232 GNDA.n231 187.249
R2812 GNDA.n1240 GNDA.n1239 187.249
R2813 GNDA.n2293 GNDA.n185 187.249
R2814 GNDA.n1894 GNDA.n1892 187.249
R2815 GNDA.n1568 GNDA.n1567 187.249
R2816 GNDA.n919 GNDA.n917 187.249
R2817 GNDA.n2088 GNDA.n2087 187.249
R2818 GNDA.n2121 GNDA.n2116 187.249
R2819 GNDA.n479 GNDA.n324 185.601
R2820 GNDA.n1487 GNDA.n1486 185
R2821 GNDA.n1488 GNDA.n1405 185
R2822 GNDA.n1405 GNDA.t233 185
R2823 GNDA.n1490 GNDA.n1489 185
R2824 GNDA.n1492 GNDA.n1404 185
R2825 GNDA.n1495 GNDA.n1494 185
R2826 GNDA.n1496 GNDA.n1403 185
R2827 GNDA.n1498 GNDA.n1497 185
R2828 GNDA.n1500 GNDA.n1402 185
R2829 GNDA.n1503 GNDA.n1502 185
R2830 GNDA.n1504 GNDA.n1401 185
R2831 GNDA.n1506 GNDA.n1505 185
R2832 GNDA.n1508 GNDA.n1400 185
R2833 GNDA.n1511 GNDA.n1510 185
R2834 GNDA.n1512 GNDA.n1399 185
R2835 GNDA.n1514 GNDA.n1513 185
R2836 GNDA.n1516 GNDA.n1398 185
R2837 GNDA.n1519 GNDA.n1518 185
R2838 GNDA.n1520 GNDA.n1397 185
R2839 GNDA.n1537 GNDA.n1536 185
R2840 GNDA.n1534 GNDA.n1391 185
R2841 GNDA.n1533 GNDA.n1393 185
R2842 GNDA.n1531 GNDA.n1530 185
R2843 GNDA.n1529 GNDA.n1394 185
R2844 GNDA.n1528 GNDA.n1527 185
R2845 GNDA.n1525 GNDA.n1395 185
R2846 GNDA.n1525 GNDA.t233 185
R2847 GNDA.n1524 GNDA.n1396 185
R2848 GNDA.n1522 GNDA.n1521 185
R2849 GNDA.n1305 GNDA.n1304 185
R2850 GNDA.n1306 GNDA.n1303 185
R2851 GNDA.n1306 GNDA.t235 185
R2852 GNDA.n1309 GNDA.n1308 185
R2853 GNDA.n1310 GNDA.n1302 185
R2854 GNDA.n1312 GNDA.n1311 185
R2855 GNDA.n1314 GNDA.n1301 185
R2856 GNDA.n1317 GNDA.n1316 185
R2857 GNDA.n1318 GNDA.n1300 185
R2858 GNDA.n1320 GNDA.n1319 185
R2859 GNDA.n1322 GNDA.n1299 185
R2860 GNDA.n1325 GNDA.n1324 185
R2861 GNDA.n1326 GNDA.n1298 185
R2862 GNDA.n1328 GNDA.n1327 185
R2863 GNDA.n1330 GNDA.n1297 185
R2864 GNDA.n1333 GNDA.n1332 185
R2865 GNDA.n1334 GNDA.n1296 185
R2866 GNDA.n1336 GNDA.n1335 185
R2867 GNDA.n1338 GNDA.n1295 185
R2868 GNDA.n1355 GNDA.n1290 185
R2869 GNDA.n1353 GNDA.n1352 185
R2870 GNDA.n1351 GNDA.n1291 185
R2871 GNDA.n1350 GNDA.n1349 185
R2872 GNDA.n1347 GNDA.n1292 185
R2873 GNDA.n1345 GNDA.n1344 185
R2874 GNDA.n1343 GNDA.n1293 185
R2875 GNDA.n1293 GNDA.t235 185
R2876 GNDA.n1342 GNDA.n1341 185
R2877 GNDA.n1339 GNDA.n1294 185
R2878 GNDA.n2204 GNDA.n2203 185
R2879 GNDA.n2205 GNDA.n2202 185
R2880 GNDA.n2205 GNDA.t309 185
R2881 GNDA.n2208 GNDA.n2207 185
R2882 GNDA.n2209 GNDA.n2201 185
R2883 GNDA.n2211 GNDA.n2210 185
R2884 GNDA.n2213 GNDA.n2200 185
R2885 GNDA.n2216 GNDA.n2215 185
R2886 GNDA.n2217 GNDA.n2199 185
R2887 GNDA.n2219 GNDA.n2218 185
R2888 GNDA.n2221 GNDA.n2198 185
R2889 GNDA.n2224 GNDA.n2223 185
R2890 GNDA.n2225 GNDA.n2197 185
R2891 GNDA.n2227 GNDA.n2226 185
R2892 GNDA.n2229 GNDA.n2196 185
R2893 GNDA.n2232 GNDA.n2231 185
R2894 GNDA.n2233 GNDA.n2195 185
R2895 GNDA.n2235 GNDA.n2234 185
R2896 GNDA.n2237 GNDA.n2194 185
R2897 GNDA.n2254 GNDA.n2189 185
R2898 GNDA.n2252 GNDA.n2251 185
R2899 GNDA.n2250 GNDA.n2190 185
R2900 GNDA.n2249 GNDA.n2248 185
R2901 GNDA.n2246 GNDA.n2191 185
R2902 GNDA.n2244 GNDA.n2243 185
R2903 GNDA.n2242 GNDA.n2192 185
R2904 GNDA.n2192 GNDA.t309 185
R2905 GNDA.n2241 GNDA.n2240 185
R2906 GNDA.n2238 GNDA.n2193 185
R2907 GNDA.n790 GNDA.n789 185
R2908 GNDA.n791 GNDA.n788 185
R2909 GNDA.n791 GNDA.t277 185
R2910 GNDA.n794 GNDA.n793 185
R2911 GNDA.n795 GNDA.n787 185
R2912 GNDA.n797 GNDA.n796 185
R2913 GNDA.n799 GNDA.n786 185
R2914 GNDA.n802 GNDA.n801 185
R2915 GNDA.n803 GNDA.n785 185
R2916 GNDA.n805 GNDA.n804 185
R2917 GNDA.n807 GNDA.n784 185
R2918 GNDA.n810 GNDA.n809 185
R2919 GNDA.n811 GNDA.n783 185
R2920 GNDA.n813 GNDA.n812 185
R2921 GNDA.n815 GNDA.n782 185
R2922 GNDA.n818 GNDA.n817 185
R2923 GNDA.n819 GNDA.n781 185
R2924 GNDA.n821 GNDA.n820 185
R2925 GNDA.n823 GNDA.n780 185
R2926 GNDA.n840 GNDA.n775 185
R2927 GNDA.n838 GNDA.n837 185
R2928 GNDA.n836 GNDA.n776 185
R2929 GNDA.n835 GNDA.n834 185
R2930 GNDA.n832 GNDA.n777 185
R2931 GNDA.n830 GNDA.n829 185
R2932 GNDA.n828 GNDA.n778 185
R2933 GNDA.n778 GNDA.t277 185
R2934 GNDA.n827 GNDA.n826 185
R2935 GNDA.n824 GNDA.n779 185
R2936 GNDA.n990 GNDA.n705 185
R2937 GNDA.n991 GNDA.n704 185
R2938 GNDA.n991 GNDA.t276 185
R2939 GNDA.n994 GNDA.n993 185
R2940 GNDA.n995 GNDA.n703 185
R2941 GNDA.n997 GNDA.n996 185
R2942 GNDA.n999 GNDA.n702 185
R2943 GNDA.n1002 GNDA.n1001 185
R2944 GNDA.n1003 GNDA.n701 185
R2945 GNDA.n1005 GNDA.n1004 185
R2946 GNDA.n1007 GNDA.n700 185
R2947 GNDA.n1010 GNDA.n1009 185
R2948 GNDA.n1011 GNDA.n699 185
R2949 GNDA.n1013 GNDA.n1012 185
R2950 GNDA.n1015 GNDA.n698 185
R2951 GNDA.n1018 GNDA.n1017 185
R2952 GNDA.n1019 GNDA.n697 185
R2953 GNDA.n1021 GNDA.n1020 185
R2954 GNDA.n1023 GNDA.n696 185
R2955 GNDA.n1040 GNDA.n688 185
R2956 GNDA.n1038 GNDA.n1037 185
R2957 GNDA.n1036 GNDA.n692 185
R2958 GNDA.n1035 GNDA.n1034 185
R2959 GNDA.n1032 GNDA.n693 185
R2960 GNDA.n1030 GNDA.n1029 185
R2961 GNDA.n1028 GNDA.n694 185
R2962 GNDA.n694 GNDA.t276 185
R2963 GNDA.n1027 GNDA.n1026 185
R2964 GNDA.n1024 GNDA.n695 185
R2965 GNDA.n1114 GNDA.n1113 185
R2966 GNDA.n1115 GNDA.n1112 185
R2967 GNDA.n1115 GNDA.t251 185
R2968 GNDA.n1118 GNDA.n1117 185
R2969 GNDA.n1119 GNDA.n1111 185
R2970 GNDA.n1121 GNDA.n1120 185
R2971 GNDA.n1123 GNDA.n1110 185
R2972 GNDA.n1126 GNDA.n1125 185
R2973 GNDA.n1127 GNDA.n1109 185
R2974 GNDA.n1129 GNDA.n1128 185
R2975 GNDA.n1131 GNDA.n1108 185
R2976 GNDA.n1134 GNDA.n1133 185
R2977 GNDA.n1135 GNDA.n1107 185
R2978 GNDA.n1137 GNDA.n1136 185
R2979 GNDA.n1139 GNDA.n1106 185
R2980 GNDA.n1142 GNDA.n1141 185
R2981 GNDA.n1143 GNDA.n1105 185
R2982 GNDA.n1145 GNDA.n1144 185
R2983 GNDA.n1147 GNDA.n1104 185
R2984 GNDA.n1164 GNDA.n1099 185
R2985 GNDA.n1162 GNDA.n1161 185
R2986 GNDA.n1160 GNDA.n1100 185
R2987 GNDA.n1159 GNDA.n1158 185
R2988 GNDA.n1156 GNDA.n1101 185
R2989 GNDA.n1154 GNDA.n1153 185
R2990 GNDA.n1152 GNDA.n1102 185
R2991 GNDA.n1102 GNDA.t251 185
R2992 GNDA.n1151 GNDA.n1150 185
R2993 GNDA.n1148 GNDA.n1103 185
R2994 GNDA.n1756 GNDA.n1755 185
R2995 GNDA.n1757 GNDA.n1753 185
R2996 GNDA.n1753 GNDA.t244 185
R2997 GNDA.n1759 GNDA.n1758 185
R2998 GNDA.n1761 GNDA.n1752 185
R2999 GNDA.n1764 GNDA.n1763 185
R3000 GNDA.n1765 GNDA.n1751 185
R3001 GNDA.n1767 GNDA.n1766 185
R3002 GNDA.n1769 GNDA.n1750 185
R3003 GNDA.n1772 GNDA.n1771 185
R3004 GNDA.n1773 GNDA.n1749 185
R3005 GNDA.n1775 GNDA.n1774 185
R3006 GNDA.n1777 GNDA.n1748 185
R3007 GNDA.n1780 GNDA.n1779 185
R3008 GNDA.n1781 GNDA.n1747 185
R3009 GNDA.n1783 GNDA.n1782 185
R3010 GNDA.n1785 GNDA.n1746 185
R3011 GNDA.n1788 GNDA.n1787 185
R3012 GNDA.n1789 GNDA.n1745 185
R3013 GNDA.n1806 GNDA.n1805 185
R3014 GNDA.n1803 GNDA.n1738 185
R3015 GNDA.n1802 GNDA.n1741 185
R3016 GNDA.n1800 GNDA.n1799 185
R3017 GNDA.n1798 GNDA.n1742 185
R3018 GNDA.n1797 GNDA.n1796 185
R3019 GNDA.n1794 GNDA.n1743 185
R3020 GNDA.n1794 GNDA.t244 185
R3021 GNDA.n1793 GNDA.n1744 185
R3022 GNDA.n1791 GNDA.n1790 185
R3023 GNDA.n1964 GNDA.n1926 185
R3024 GNDA.n1966 GNDA.n1965 185
R3025 GNDA.n1965 GNDA.t240 185
R3026 GNDA.n1968 GNDA.n1967 185
R3027 GNDA.n1970 GNDA.n1963 185
R3028 GNDA.n1973 GNDA.n1972 185
R3029 GNDA.n1974 GNDA.n1962 185
R3030 GNDA.n1976 GNDA.n1975 185
R3031 GNDA.n1978 GNDA.n1961 185
R3032 GNDA.n1981 GNDA.n1980 185
R3033 GNDA.n1982 GNDA.n1960 185
R3034 GNDA.n1984 GNDA.n1983 185
R3035 GNDA.n1986 GNDA.n1959 185
R3036 GNDA.n1989 GNDA.n1988 185
R3037 GNDA.n1990 GNDA.n1958 185
R3038 GNDA.n1992 GNDA.n1991 185
R3039 GNDA.n1994 GNDA.n1957 185
R3040 GNDA.n1997 GNDA.n1996 185
R3041 GNDA.n1998 GNDA.n1956 185
R3042 GNDA.n2015 GNDA.n2014 185
R3043 GNDA.n2012 GNDA.n1949 185
R3044 GNDA.n2011 GNDA.n1952 185
R3045 GNDA.n2009 GNDA.n2008 185
R3046 GNDA.n2007 GNDA.n1953 185
R3047 GNDA.n2006 GNDA.n2005 185
R3048 GNDA.n2003 GNDA.n1954 185
R3049 GNDA.n2003 GNDA.t240 185
R3050 GNDA.n2002 GNDA.n1955 185
R3051 GNDA.n2000 GNDA.n1999 185
R3052 GNDA.n2349 GNDA.n139 185
R3053 GNDA.n2350 GNDA.n138 185
R3054 GNDA.n2350 GNDA.t229 185
R3055 GNDA.n2353 GNDA.n2352 185
R3056 GNDA.n2354 GNDA.n137 185
R3057 GNDA.n2356 GNDA.n2355 185
R3058 GNDA.n2358 GNDA.n136 185
R3059 GNDA.n2361 GNDA.n2360 185
R3060 GNDA.n2362 GNDA.n135 185
R3061 GNDA.n2364 GNDA.n2363 185
R3062 GNDA.n2366 GNDA.n134 185
R3063 GNDA.n2369 GNDA.n2368 185
R3064 GNDA.n2370 GNDA.n133 185
R3065 GNDA.n2372 GNDA.n2371 185
R3066 GNDA.n2374 GNDA.n132 185
R3067 GNDA.n2377 GNDA.n2376 185
R3068 GNDA.n2378 GNDA.n131 185
R3069 GNDA.n2380 GNDA.n2379 185
R3070 GNDA.n2382 GNDA.n130 185
R3071 GNDA.n2399 GNDA.n90 185
R3072 GNDA.n2397 GNDA.n2396 185
R3073 GNDA.n2395 GNDA.n126 185
R3074 GNDA.n2394 GNDA.n2393 185
R3075 GNDA.n2391 GNDA.n127 185
R3076 GNDA.n2389 GNDA.n2388 185
R3077 GNDA.n2387 GNDA.n128 185
R3078 GNDA.n128 GNDA.t229 185
R3079 GNDA.n2386 GNDA.n2385 185
R3080 GNDA.n2383 GNDA.n129 185
R3081 GNDA.n2400 GNDA.n89 185
R3082 GNDA.n2404 GNDA.n2402 185
R3083 GNDA.n2409 GNDA.n2408 185
R3084 GNDA.n2412 GNDA.n2411 185
R3085 GNDA.n125 GNDA.n123 185
R3086 GNDA.n2338 GNDA.n2337 185
R3087 GNDA.n2335 GNDA.n2332 185
R3088 GNDA.n142 GNDA.n140 185
R3089 GNDA.n2347 GNDA.n2346 185
R3090 GNDA.n1951 GNDA.n1948 185
R3091 GNDA.n1940 GNDA.n1938 185
R3092 GNDA.n2031 GNDA.n2030 185
R3093 GNDA.n2033 GNDA.n1937 185
R3094 GNDA.n2035 GNDA.n2034 185
R3095 GNDA.n1932 GNDA.n1930 185
R3096 GNDA.n2046 GNDA.n2045 185
R3097 GNDA.n2048 GNDA.n1929 185
R3098 GNDA.n2050 GNDA.n2049 185
R3099 GNDA.n1740 GNDA.n1737 185
R3100 GNDA.n1602 GNDA.n1601 185
R3101 GNDA.n1822 GNDA.n1821 185
R3102 GNDA.n1825 GNDA.n1824 185
R3103 GNDA.n1600 GNDA.n1597 185
R3104 GNDA.n608 GNDA.n607 185
R3105 GNDA.n1834 GNDA.n1833 185
R3106 GNDA.n1837 GNDA.n1836 185
R3107 GNDA.n606 GNDA.n604 185
R3108 GNDA.n1166 GNDA.n1165 185
R3109 GNDA.n1088 GNDA.n1086 185
R3110 GNDA.n1173 GNDA.n1172 185
R3111 GNDA.n1175 GNDA.n1085 185
R3112 GNDA.n1177 GNDA.n1176 185
R3113 GNDA.n1079 GNDA.n1077 185
R3114 GNDA.n1184 GNDA.n1183 185
R3115 GNDA.n1186 GNDA.n1076 185
R3116 GNDA.n1188 GNDA.n1187 185
R3117 GNDA.n1042 GNDA.n1041 185
R3118 GNDA.n965 GNDA.n964 185
R3119 GNDA.n963 GNDA.n961 185
R3120 GNDA.n970 GNDA.n960 185
R3121 GNDA.n975 GNDA.n974 185
R3122 GNDA.n978 GNDA.n977 185
R3123 GNDA.n959 GNDA.n956 185
R3124 GNDA.n983 GNDA.n706 185
R3125 GNDA.n988 GNDA.n987 185
R3126 GNDA.n842 GNDA.n841 185
R3127 GNDA.n760 GNDA.n758 185
R3128 GNDA.n849 GNDA.n848 185
R3129 GNDA.n851 GNDA.n757 185
R3130 GNDA.n853 GNDA.n852 185
R3131 GNDA.n751 GNDA.n749 185
R3132 GNDA.n860 GNDA.n859 185
R3133 GNDA.n862 GNDA.n748 185
R3134 GNDA.n864 GNDA.n863 185
R3135 GNDA.n2256 GNDA.n2255 185
R3136 GNDA.n299 GNDA.n297 185
R3137 GNDA.n2263 GNDA.n2262 185
R3138 GNDA.n2265 GNDA.n296 185
R3139 GNDA.n2267 GNDA.n2266 185
R3140 GNDA.n290 GNDA.n288 185
R3141 GNDA.n2274 GNDA.n2273 185
R3142 GNDA.n2276 GNDA.n287 185
R3143 GNDA.n2278 GNDA.n2277 185
R3144 GNDA.n1357 GNDA.n1356 185
R3145 GNDA.n1280 GNDA.n1278 185
R3146 GNDA.n1364 GNDA.n1363 185
R3147 GNDA.n1366 GNDA.n1277 185
R3148 GNDA.n1368 GNDA.n1367 185
R3149 GNDA.n1271 GNDA.n1269 185
R3150 GNDA.n1375 GNDA.n1374 185
R3151 GNDA.n1377 GNDA.n1268 185
R3152 GNDA.n1379 GNDA.n1378 185
R3153 GNDA.n1392 GNDA.n1390 185
R3154 GNDA.n1464 GNDA.n1462 185
R3155 GNDA.n1466 GNDA.n1465 185
R3156 GNDA.n1454 GNDA.n1452 185
R3157 GNDA.n1473 GNDA.n1472 185
R3158 GNDA.n1475 GNDA.n1451 185
R3159 GNDA.n1477 GNDA.n1476 185
R3160 GNDA.n1409 GNDA.n1407 185
R3161 GNDA.n1484 GNDA.n1483 185
R3162 GNDA.n462 GNDA.n461 182.4
R3163 GNDA.n377 GNDA.n376 182.4
R3164 GNDA.n432 GNDA.n394 182.4
R3165 GNDA.n2057 GNDA.n2056 181.233
R3166 GNDA.n2092 GNDA.n145 181.233
R3167 GNDA.n466 GNDA.t274 181.226
R3168 GNDA.n451 GNDA.t246 181.226
R3169 GNDA.n1689 GNDA.n1625 179.917
R3170 GNDA.n1723 GNDA.n1615 176
R3171 GNDA.n1723 GNDA.n1722 176
R3172 GNDA.n2280 GNDA.n284 175.546
R3173 GNDA.n2271 GNDA.n292 175.546
R3174 GNDA.n2269 GNDA.n293 175.546
R3175 GNDA.n2260 GNDA.n301 175.546
R3176 GNDA.n2258 GNDA.n302 175.546
R3177 GNDA.n494 GNDA.n175 175.546
R3178 GNDA.n498 GNDA.n494 175.546
R3179 GNDA.n498 GNDA.n492 175.546
R3180 GNDA.n2156 GNDA.n492 175.546
R3181 GNDA.n2156 GNDA.n489 175.546
R3182 GNDA.n2162 GNDA.n489 175.546
R3183 GNDA.n2162 GNDA.n490 175.546
R3184 GNDA.n490 GNDA.n309 175.546
R3185 GNDA.n2180 GNDA.n309 175.546
R3186 GNDA.n2181 GNDA.n2180 175.546
R3187 GNDA.n2301 GNDA.n181 175.546
R3188 GNDA.n2305 GNDA.n2303 175.546
R3189 GNDA.n2309 GNDA.n179 175.546
R3190 GNDA.n2313 GNDA.n2311 175.546
R3191 GNDA.n2317 GNDA.n177 175.546
R3192 GNDA.n259 GNDA.n258 175.546
R3193 GNDA.n264 GNDA.n263 175.546
R3194 GNDA.n270 GNDA.n269 175.546
R3195 GNDA.n276 GNDA.n275 175.546
R3196 GNDA.n2285 GNDA.n2284 175.546
R3197 GNDA.n2328 GNDA.n143 175.546
R3198 GNDA.n2344 GNDA.n143 175.546
R3199 GNDA.n2344 GNDA.n144 175.546
R3200 GNDA.n2340 GNDA.n144 175.546
R3201 GNDA.n2340 GNDA.n121 175.546
R3202 GNDA.n2414 GNDA.n121 175.546
R3203 GNDA.n2414 GNDA.n122 175.546
R3204 GNDA.n2406 GNDA.n122 175.546
R3205 GNDA.n2406 GNDA.n87 175.546
R3206 GNDA.n2437 GNDA.n87 175.546
R3207 GNDA.n2437 GNDA.n88 175.546
R3208 GNDA.n231 GNDA.n217 175.546
R3209 GNDA.n227 GNDA.n217 175.546
R3210 GNDA.n227 GNDA.n220 175.546
R3211 GNDA.n223 GNDA.n220 175.546
R3212 GNDA.n223 GNDA.n115 175.546
R3213 GNDA.n2417 GNDA.n115 175.546
R3214 GNDA.n2417 GNDA.n109 175.546
R3215 GNDA.n2422 GNDA.n109 175.546
R3216 GNDA.n2422 GNDA.n113 175.546
R3217 GNDA.n113 GNDA.n112 175.546
R3218 GNDA.n253 GNDA.n252 175.546
R3219 GNDA.n249 GNDA.n248 175.546
R3220 GNDA.n246 GNDA.n212 175.546
R3221 GNDA.n242 GNDA.n240 175.546
R3222 GNDA.n238 GNDA.n214 175.546
R3223 GNDA.n1212 GNDA.n161 175.546
R3224 GNDA.n1214 GNDA.n1213 175.546
R3225 GNDA.n1216 GNDA.n1215 175.546
R3226 GNDA.n1218 GNDA.n1217 175.546
R3227 GNDA.n1219 GNDA.n148 175.546
R3228 GNDA.n2054 GNDA.n563 175.546
R3229 GNDA.n2038 GNDA.n563 175.546
R3230 GNDA.n2038 GNDA.n1933 175.546
R3231 GNDA.n2043 GNDA.n1933 175.546
R3232 GNDA.n2043 GNDA.n2037 175.546
R3233 GNDA.n2037 GNDA.n1934 175.546
R3234 GNDA.n1941 GNDA.n1934 175.546
R3235 GNDA.n2028 GNDA.n1941 175.546
R3236 GNDA.n2028 GNDA.n1942 175.546
R3237 GNDA.n2024 GNDA.n1942 175.546
R3238 GNDA.n2024 GNDA.n1946 175.546
R3239 GNDA.n1236 GNDA.n1235 175.546
R3240 GNDA.n1232 GNDA.n1231 175.546
R3241 GNDA.n1228 GNDA.n1227 175.546
R3242 GNDA.n1224 GNDA.n1223 175.546
R3243 GNDA.n1220 GNDA.n199 175.546
R3244 GNDA.n1261 GNDA.n1209 175.546
R3245 GNDA.n1257 GNDA.n1256 175.546
R3246 GNDA.n1253 GNDA.n1252 175.546
R3247 GNDA.n1249 GNDA.n1248 175.546
R3248 GNDA.n1245 GNDA.n1244 175.546
R3249 GNDA.n1897 GNDA.n1896 175.546
R3250 GNDA.n1900 GNDA.n1899 175.546
R3251 GNDA.n1909 GNDA.n1908 175.546
R3252 GNDA.n1913 GNDA.n1912 175.546
R3253 GNDA.n1922 GNDA.n565 175.546
R3254 GNDA.n1381 GNDA.n1265 175.546
R3255 GNDA.n1372 GNDA.n1273 175.546
R3256 GNDA.n1370 GNDA.n1274 175.546
R3257 GNDA.n1361 GNDA.n1282 175.546
R3258 GNDA.n1359 GNDA.n1283 175.546
R3259 GNDA.n260 GNDA.n186 175.546
R3260 GNDA.n266 GNDA.n265 175.546
R3261 GNDA.n272 GNDA.n271 175.546
R3262 GNDA.n278 GNDA.n277 175.546
R3263 GNDA.n280 GNDA.n188 175.546
R3264 GNDA.n674 GNDA.n655 175.546
R3265 GNDA.n672 GNDA.n671 175.546
R3266 GNDA.n668 GNDA.n667 175.546
R3267 GNDA.n664 GNDA.n663 175.546
R3268 GNDA.n660 GNDA.n659 175.546
R3269 GNDA.n631 GNDA.n628 175.546
R3270 GNDA.n634 GNDA.n633 175.546
R3271 GNDA.n639 GNDA.n636 175.546
R3272 GNDA.n642 GNDA.n641 175.546
R3273 GNDA.n646 GNDA.n644 175.546
R3274 GNDA.n1843 GNDA.n600 175.546
R3275 GNDA.n1839 GNDA.n600 175.546
R3276 GNDA.n1839 GNDA.n602 175.546
R3277 GNDA.n1831 GNDA.n602 175.546
R3278 GNDA.n1831 GNDA.n609 175.546
R3279 GNDA.n1827 GNDA.n609 175.546
R3280 GNDA.n1827 GNDA.n1595 175.546
R3281 GNDA.n1819 GNDA.n1595 175.546
R3282 GNDA.n1819 GNDA.n1603 175.546
R3283 GNDA.n1815 GNDA.n1603 175.546
R3284 GNDA.n1815 GNDA.n1735 175.546
R3285 GNDA.n1902 GNDA.n573 175.546
R3286 GNDA.n1906 GNDA.n1904 175.546
R3287 GNDA.n1915 GNDA.n569 175.546
R3288 GNDA.n1918 GNDA.n1917 175.546
R3289 GNDA.n1920 GNDA.n567 175.546
R3290 GNDA.n1873 GNDA.n584 175.546
R3291 GNDA.n1877 GNDA.n1875 175.546
R3292 GNDA.n1881 GNDA.n582 175.546
R3293 GNDA.n1885 GNDA.n1883 175.546
R3294 GNDA.n1889 GNDA.n580 175.546
R3295 GNDA.n1867 GNDA.n586 175.546
R3296 GNDA.n1863 GNDA.n586 175.546
R3297 GNDA.n1863 GNDA.n589 175.546
R3298 GNDA.n1859 GNDA.n589 175.546
R3299 GNDA.n1859 GNDA.n592 175.546
R3300 GNDA.n1855 GNDA.n592 175.546
R3301 GNDA.n1855 GNDA.n594 175.546
R3302 GNDA.n1851 GNDA.n594 175.546
R3303 GNDA.n1851 GNDA.n596 175.546
R3304 GNDA.n1847 GNDA.n596 175.546
R3305 GNDA.n1481 GNDA.n1447 175.546
R3306 GNDA.n1479 GNDA.n1448 175.546
R3307 GNDA.n1470 GNDA.n1456 175.546
R3308 GNDA.n1468 GNDA.n1458 175.546
R3309 GNDA.n1540 GNDA.n1389 175.546
R3310 GNDA.n1564 GNDA.n1563 175.546
R3311 GNDA.n1561 GNDA.n630 175.546
R3312 GNDA.n1557 GNDA.n1555 175.546
R3313 GNDA.n1553 GNDA.n638 175.546
R3314 GNDA.n1549 GNDA.n1547 175.546
R3315 GNDA.n1587 GNDA.n620 175.546
R3316 GNDA.n1585 GNDA.n1584 175.546
R3317 GNDA.n1581 GNDA.n1580 175.546
R3318 GNDA.n1577 GNDA.n1576 175.546
R3319 GNDA.n1573 GNDA.n1572 175.546
R3320 GNDA.n1420 GNDA.n621 175.546
R3321 GNDA.n1424 GNDA.n1420 175.546
R3322 GNDA.n1424 GNDA.n1418 175.546
R3323 GNDA.n1428 GNDA.n1418 175.546
R3324 GNDA.n1428 GNDA.n1416 175.546
R3325 GNDA.n1432 GNDA.n1416 175.546
R3326 GNDA.n1432 GNDA.n1414 175.546
R3327 GNDA.n1436 GNDA.n1414 175.546
R3328 GNDA.n1436 GNDA.n1412 175.546
R3329 GNDA.n1441 GNDA.n1412 175.546
R3330 GNDA.n866 GNDA.n744 175.546
R3331 GNDA.n857 GNDA.n753 175.546
R3332 GNDA.n855 GNDA.n754 175.546
R3333 GNDA.n846 GNDA.n762 175.546
R3334 GNDA.n844 GNDA.n763 175.546
R3335 GNDA.n891 GNDA.n732 175.546
R3336 GNDA.n887 GNDA.n732 175.546
R3337 GNDA.n887 GNDA.n734 175.546
R3338 GNDA.n883 GNDA.n734 175.546
R3339 GNDA.n883 GNDA.n736 175.546
R3340 GNDA.n879 GNDA.n736 175.546
R3341 GNDA.n879 GNDA.n738 175.546
R3342 GNDA.n875 GNDA.n738 175.546
R3343 GNDA.n875 GNDA.n740 175.546
R3344 GNDA.n871 GNDA.n740 175.546
R3345 GNDA.n927 GNDA.n717 175.546
R3346 GNDA.n931 GNDA.n929 175.546
R3347 GNDA.n941 GNDA.n713 175.546
R3348 GNDA.n944 GNDA.n943 175.546
R3349 GNDA.n946 GNDA.n711 175.546
R3350 GNDA.n895 GNDA.n730 175.546
R3351 GNDA.n895 GNDA.n728 175.546
R3352 GNDA.n900 GNDA.n728 175.546
R3353 GNDA.n900 GNDA.n726 175.546
R3354 GNDA.n904 GNDA.n726 175.546
R3355 GNDA.n905 GNDA.n904 175.546
R3356 GNDA.n907 GNDA.n905 175.546
R3357 GNDA.n907 GNDA.n724 175.546
R3358 GNDA.n912 GNDA.n724 175.546
R3359 GNDA.n912 GNDA.n720 175.546
R3360 GNDA.n916 GNDA.n720 175.546
R3361 GNDA.n985 GNDA.n984 175.546
R3362 GNDA.n981 GNDA.n980 175.546
R3363 GNDA.n972 GNDA.n971 175.546
R3364 GNDA.n968 GNDA.n967 175.546
R3365 GNDA.n689 GNDA.n686 175.546
R3366 GNDA.n925 GNDA.n923 175.546
R3367 GNDA.n933 GNDA.n715 175.546
R3368 GNDA.n939 GNDA.n935 175.546
R3369 GNDA.n937 GNDA.n936 175.546
R3370 GNDA.n949 GNDA.n948 175.546
R3371 GNDA.n1049 GNDA.n1048 175.546
R3372 GNDA.n1055 GNDA.n1054 175.546
R3373 GNDA.n1061 GNDA.n1060 175.546
R3374 GNDA.n1067 GNDA.n1066 175.546
R3375 GNDA.n1069 GNDA.n193 175.546
R3376 GNDA.n2059 GNDA.n556 175.546
R3377 GNDA.n2059 GNDA.n554 175.546
R3378 GNDA.n2063 GNDA.n554 175.546
R3379 GNDA.n2063 GNDA.n552 175.546
R3380 GNDA.n2067 GNDA.n552 175.546
R3381 GNDA.n2067 GNDA.n542 175.546
R3382 GNDA.n2077 GNDA.n542 175.546
R3383 GNDA.n2077 GNDA.n540 175.546
R3384 GNDA.n2082 GNDA.n540 175.546
R3385 GNDA.n2082 GNDA.n536 175.546
R3386 GNDA.n2086 GNDA.n536 175.546
R3387 GNDA.n1190 GNDA.n1073 175.546
R3388 GNDA.n1181 GNDA.n1081 175.546
R3389 GNDA.n1179 GNDA.n1082 175.546
R3390 GNDA.n1170 GNDA.n1090 175.546
R3391 GNDA.n1168 GNDA.n1091 175.546
R3392 GNDA.n2121 GNDA.n521 175.546
R3393 GNDA.n2125 GNDA.n521 175.546
R3394 GNDA.n2125 GNDA.n519 175.546
R3395 GNDA.n2130 GNDA.n519 175.546
R3396 GNDA.n2130 GNDA.n517 175.546
R3397 GNDA.n2134 GNDA.n517 175.546
R3398 GNDA.n2134 GNDA.n516 175.546
R3399 GNDA.n2138 GNDA.n516 175.546
R3400 GNDA.n2138 GNDA.n512 175.546
R3401 GNDA.n2143 GNDA.n512 175.546
R3402 GNDA.n2094 GNDA.n2091 175.546
R3403 GNDA.n2094 GNDA.n531 175.546
R3404 GNDA.n2098 GNDA.n531 175.546
R3405 GNDA.n2098 GNDA.n529 175.546
R3406 GNDA.n2102 GNDA.n529 175.546
R3407 GNDA.n2102 GNDA.n527 175.546
R3408 GNDA.n2106 GNDA.n527 175.546
R3409 GNDA.n2106 GNDA.n525 175.546
R3410 GNDA.n2111 GNDA.n525 175.546
R3411 GNDA.n2111 GNDA.n523 175.546
R3412 GNDA.n2115 GNDA.n523 175.546
R3413 GNDA.n1047 GNDA.n1046 175.546
R3414 GNDA.n1053 GNDA.n1052 175.546
R3415 GNDA.n1059 GNDA.n1058 175.546
R3416 GNDA.n1065 GNDA.n1064 175.546
R3417 GNDA.n1195 GNDA.n1194 175.546
R3418 GNDA.n2474 GNDA.t43 174.101
R3419 GNDA.n2474 GNDA.t35 174.101
R3420 GNDA.n456 GNDA.t275 169.566
R3421 GNDA.n323 GNDA.t257 169.566
R3422 GNDA.n441 GNDA.t260 169.566
R3423 GNDA.n430 GNDA.t247 169.566
R3424 GNDA.n1536 GNDA.n1392 163.333
R3425 GNDA.n1356 GNDA.n1355 163.333
R3426 GNDA.n2255 GNDA.n2254 163.333
R3427 GNDA.n841 GNDA.n840 163.333
R3428 GNDA.n1041 GNDA.n1040 163.333
R3429 GNDA.n1165 GNDA.n1164 163.333
R3430 GNDA.n1805 GNDA.n1740 163.333
R3431 GNDA.n2014 GNDA.n1951 163.333
R3432 GNDA.n2400 GNDA.n2399 163.333
R3433 GNDA.n1644 GNDA.t272 160.725
R3434 GNDA.n1645 GNDA.t269 160.725
R3435 GNDA.n1616 GNDA.t266 160.725
R3436 GNDA.n1614 GNDA.t239 160.725
R3437 GNDA.n1618 GNDA.t296 160.725
R3438 GNDA.n1703 GNDA.t305 160.725
R3439 GNDA.n1715 GNDA.n1714 159.778
R3440 GNDA.n1640 GNDA.n1639 159.778
R3441 GNDA.n548 GNDA.t139 157.555
R3442 GNDA.n547 GNDA.t334 157.555
R3443 GNDA.n1648 GNDA.t126 153.294
R3444 GNDA.n2324 GNDA.n2323 152.643
R3445 GNDA.n1924 GNDA.n1923 152.643
R3446 GNDA.n102 GNDA.n94 150.614
R3447 GNDA.n1484 GNDA.n1407 150
R3448 GNDA.n1476 GNDA.n1475 150
R3449 GNDA.n1473 GNDA.n1452 150
R3450 GNDA.n1465 GNDA.n1464 150
R3451 GNDA.n1525 GNDA.n1524 150
R3452 GNDA.n1527 GNDA.n1525 150
R3453 GNDA.n1531 GNDA.n1394 150
R3454 GNDA.n1534 GNDA.n1533 150
R3455 GNDA.n1506 GNDA.n1401 150
R3456 GNDA.n1510 GNDA.n1508 150
R3457 GNDA.n1514 GNDA.n1399 150
R3458 GNDA.n1518 GNDA.n1516 150
R3459 GNDA.n1502 GNDA.n1500 150
R3460 GNDA.n1498 GNDA.n1403 150
R3461 GNDA.n1494 GNDA.n1492 150
R3462 GNDA.n1490 GNDA.n1405 150
R3463 GNDA.n1486 GNDA.n1405 150
R3464 GNDA.n1378 GNDA.n1377 150
R3465 GNDA.n1375 GNDA.n1269 150
R3466 GNDA.n1367 GNDA.n1366 150
R3467 GNDA.n1364 GNDA.n1278 150
R3468 GNDA.n1341 GNDA.n1293 150
R3469 GNDA.n1345 GNDA.n1293 150
R3470 GNDA.n1349 GNDA.n1347 150
R3471 GNDA.n1353 GNDA.n1291 150
R3472 GNDA.n1324 GNDA.n1322 150
R3473 GNDA.n1328 GNDA.n1298 150
R3474 GNDA.n1332 GNDA.n1330 150
R3475 GNDA.n1336 GNDA.n1296 150
R3476 GNDA.n1320 GNDA.n1300 150
R3477 GNDA.n1316 GNDA.n1314 150
R3478 GNDA.n1312 GNDA.n1302 150
R3479 GNDA.n1308 GNDA.n1306 150
R3480 GNDA.n1306 GNDA.n1305 150
R3481 GNDA.n2277 GNDA.n2276 150
R3482 GNDA.n2274 GNDA.n288 150
R3483 GNDA.n2266 GNDA.n2265 150
R3484 GNDA.n2263 GNDA.n297 150
R3485 GNDA.n2240 GNDA.n2192 150
R3486 GNDA.n2244 GNDA.n2192 150
R3487 GNDA.n2248 GNDA.n2246 150
R3488 GNDA.n2252 GNDA.n2190 150
R3489 GNDA.n2223 GNDA.n2221 150
R3490 GNDA.n2227 GNDA.n2197 150
R3491 GNDA.n2231 GNDA.n2229 150
R3492 GNDA.n2235 GNDA.n2195 150
R3493 GNDA.n2219 GNDA.n2199 150
R3494 GNDA.n2215 GNDA.n2213 150
R3495 GNDA.n2211 GNDA.n2201 150
R3496 GNDA.n2207 GNDA.n2205 150
R3497 GNDA.n2205 GNDA.n2204 150
R3498 GNDA.n863 GNDA.n862 150
R3499 GNDA.n860 GNDA.n749 150
R3500 GNDA.n852 GNDA.n851 150
R3501 GNDA.n849 GNDA.n758 150
R3502 GNDA.n826 GNDA.n778 150
R3503 GNDA.n830 GNDA.n778 150
R3504 GNDA.n834 GNDA.n832 150
R3505 GNDA.n838 GNDA.n776 150
R3506 GNDA.n809 GNDA.n807 150
R3507 GNDA.n813 GNDA.n783 150
R3508 GNDA.n817 GNDA.n815 150
R3509 GNDA.n821 GNDA.n781 150
R3510 GNDA.n805 GNDA.n785 150
R3511 GNDA.n801 GNDA.n799 150
R3512 GNDA.n797 GNDA.n787 150
R3513 GNDA.n793 GNDA.n791 150
R3514 GNDA.n791 GNDA.n790 150
R3515 GNDA.n988 GNDA.n706 150
R3516 GNDA.n977 GNDA.n959 150
R3517 GNDA.n975 GNDA.n960 150
R3518 GNDA.n964 GNDA.n963 150
R3519 GNDA.n1026 GNDA.n694 150
R3520 GNDA.n1030 GNDA.n694 150
R3521 GNDA.n1034 GNDA.n1032 150
R3522 GNDA.n1038 GNDA.n692 150
R3523 GNDA.n1009 GNDA.n1007 150
R3524 GNDA.n1013 GNDA.n699 150
R3525 GNDA.n1017 GNDA.n1015 150
R3526 GNDA.n1021 GNDA.n697 150
R3527 GNDA.n1005 GNDA.n701 150
R3528 GNDA.n1001 GNDA.n999 150
R3529 GNDA.n997 GNDA.n703 150
R3530 GNDA.n993 GNDA.n991 150
R3531 GNDA.n991 GNDA.n990 150
R3532 GNDA.n1187 GNDA.n1186 150
R3533 GNDA.n1184 GNDA.n1077 150
R3534 GNDA.n1176 GNDA.n1175 150
R3535 GNDA.n1173 GNDA.n1086 150
R3536 GNDA.n1150 GNDA.n1102 150
R3537 GNDA.n1154 GNDA.n1102 150
R3538 GNDA.n1158 GNDA.n1156 150
R3539 GNDA.n1162 GNDA.n1100 150
R3540 GNDA.n1133 GNDA.n1131 150
R3541 GNDA.n1137 GNDA.n1107 150
R3542 GNDA.n1141 GNDA.n1139 150
R3543 GNDA.n1145 GNDA.n1105 150
R3544 GNDA.n1129 GNDA.n1109 150
R3545 GNDA.n1125 GNDA.n1123 150
R3546 GNDA.n1121 GNDA.n1111 150
R3547 GNDA.n1117 GNDA.n1115 150
R3548 GNDA.n1115 GNDA.n1114 150
R3549 GNDA.n1836 GNDA.n606 150
R3550 GNDA.n1834 GNDA.n607 150
R3551 GNDA.n1824 GNDA.n1600 150
R3552 GNDA.n1822 GNDA.n1601 150
R3553 GNDA.n1794 GNDA.n1793 150
R3554 GNDA.n1796 GNDA.n1794 150
R3555 GNDA.n1800 GNDA.n1742 150
R3556 GNDA.n1803 GNDA.n1802 150
R3557 GNDA.n1775 GNDA.n1749 150
R3558 GNDA.n1779 GNDA.n1777 150
R3559 GNDA.n1783 GNDA.n1747 150
R3560 GNDA.n1787 GNDA.n1785 150
R3561 GNDA.n1771 GNDA.n1769 150
R3562 GNDA.n1767 GNDA.n1751 150
R3563 GNDA.n1763 GNDA.n1761 150
R3564 GNDA.n1759 GNDA.n1753 150
R3565 GNDA.n1755 GNDA.n1753 150
R3566 GNDA.n2049 GNDA.n2048 150
R3567 GNDA.n2046 GNDA.n1930 150
R3568 GNDA.n2034 GNDA.n2033 150
R3569 GNDA.n2031 GNDA.n1938 150
R3570 GNDA.n2003 GNDA.n2002 150
R3571 GNDA.n2005 GNDA.n2003 150
R3572 GNDA.n2009 GNDA.n1953 150
R3573 GNDA.n2012 GNDA.n2011 150
R3574 GNDA.n1984 GNDA.n1960 150
R3575 GNDA.n1988 GNDA.n1986 150
R3576 GNDA.n1992 GNDA.n1958 150
R3577 GNDA.n1996 GNDA.n1994 150
R3578 GNDA.n1980 GNDA.n1978 150
R3579 GNDA.n1976 GNDA.n1962 150
R3580 GNDA.n1972 GNDA.n1970 150
R3581 GNDA.n1968 GNDA.n1965 150
R3582 GNDA.n1965 GNDA.n1964 150
R3583 GNDA.n2347 GNDA.n140 150
R3584 GNDA.n2337 GNDA.n2335 150
R3585 GNDA.n2411 GNDA.n125 150
R3586 GNDA.n2409 GNDA.n2402 150
R3587 GNDA.n2385 GNDA.n128 150
R3588 GNDA.n2389 GNDA.n128 150
R3589 GNDA.n2393 GNDA.n2391 150
R3590 GNDA.n2397 GNDA.n126 150
R3591 GNDA.n2368 GNDA.n2366 150
R3592 GNDA.n2372 GNDA.n133 150
R3593 GNDA.n2376 GNDA.n2374 150
R3594 GNDA.n2380 GNDA.n131 150
R3595 GNDA.n2364 GNDA.n135 150
R3596 GNDA.n2360 GNDA.n2358 150
R3597 GNDA.n2356 GNDA.n137 150
R3598 GNDA.n2352 GNDA.n2350 150
R3599 GNDA.n2350 GNDA.n2349 150
R3600 GNDA.n545 GNDA.t22 148.906
R3601 GNDA.n2478 GNDA.n33 148.8
R3602 GNDA.n545 GNDA.t321 148.653
R3603 GNDA.n465 GNDA.t301 147.511
R3604 GNDA.n452 GNDA.t311 147.511
R3605 GNDA.n2486 GNDA.n2485 145.601
R3606 GNDA.n94 GNDA.n86 145.013
R3607 GNDA.n375 GNDA.n348 144
R3608 GNDA.n433 GNDA.n426 144
R3609 GNDA.t295 GNDA.t34 141.341
R3610 GNDA.t99 GNDA.t268 141.341
R3611 GNDA.n1651 GNDA.n1649 139.638
R3612 GNDA.n1667 GNDA.n1666 139.077
R3613 GNDA.n1665 GNDA.n1664 139.077
R3614 GNDA.n1663 GNDA.n1662 139.077
R3615 GNDA.n1661 GNDA.n1660 139.077
R3616 GNDA.n1659 GNDA.n1658 139.077
R3617 GNDA.n1657 GNDA.n1656 139.077
R3618 GNDA.n1655 GNDA.n1654 139.077
R3619 GNDA.n1653 GNDA.n1652 139.077
R3620 GNDA.n1651 GNDA.n1650 139.077
R3621 GNDA.t238 GNDA.t324 135.196
R3622 GNDA.t324 GNDA.t132 135.196
R3623 GNDA.t132 GNDA.t141 135.196
R3624 GNDA.t116 GNDA.t84 135.196
R3625 GNDA.t196 GNDA.t116 135.196
R3626 GNDA.t265 GNDA.t196 135.196
R3627 GNDA.n477 GNDA.n476 134.867
R3628 GNDA.n445 GNDA.n60 134.867
R3629 GNDA.n1726 GNDA.t141 129.05
R3630 GNDA.t84 GNDA.n1638 129.05
R3631 GNDA.t80 GNDA.t227 126.62
R3632 GNDA.t106 GNDA.t67 126.62
R3633 GNDA.t292 GNDA.t39 126.62
R3634 GNDA.t77 GNDA.t262 126.62
R3635 GNDA.t37 GNDA.t105 126.62
R3636 GNDA.t221 GNDA.t18 126.62
R3637 GNDA.n2186 GNDA.n2185 124.832
R3638 GNDA.n2320 GNDA.n2319 124.832
R3639 GNDA.n2432 GNDA.n88 124.832
R3640 GNDA.n234 GNDA.n232 124.832
R3641 GNDA.n2019 GNDA.n1946 124.832
R3642 GNDA.n1241 GNDA.n1240 124.832
R3643 GNDA.n1287 GNDA.n207 124.832
R3644 GNDA.n656 GNDA.n185 124.832
R3645 GNDA.n1810 GNDA.n1735 124.832
R3646 GNDA.n1892 GNDA.n1891 124.832
R3647 GNDA.n1543 GNDA.n1542 124.832
R3648 GNDA.n1569 GNDA.n1568 124.832
R3649 GNDA.n772 GNDA.n771 124.832
R3650 GNDA.n917 GNDA.n916 124.832
R3651 GNDA.n1201 GNDA.n687 124.832
R3652 GNDA.n2087 GNDA.n2086 124.832
R3653 GNDA.n1096 GNDA.n1094 124.832
R3654 GNDA.n2116 GNDA.n2115 124.832
R3655 GNDA.n2464 GNDA.n55 124.8
R3656 GNDA.n2463 GNDA.n58 124.8
R3657 GNDA.n332 GNDA.n53 124.8
R3658 GNDA.n335 GNDA.n334 124.8
R3659 GNDA.n454 GNDA.n390 124.8
R3660 GNDA.n480 GNDA.n322 123.201
R3661 GNDA.n1707 GNDA.t17 122.906
R3662 GNDA.n1674 GNDA.t159 122.906
R3663 GNDA.n2056 GNDA.n557 119.035
R3664 GNDA.n535 GNDA.n145 119.035
R3665 GNDA.n1646 GNDA.n1617 118.4
R3666 GNDA.n1672 GNDA.n1647 118.4
R3667 GNDA.n1719 GNDA.n1615 118.4
R3668 GNDA.n1722 GNDA.n1721 118.4
R3669 GNDA.n1705 GNDA.n1704 118.4
R3670 GNDA.n1718 GNDA.n1619 118.4
R3671 GNDA.t128 GNDA.t203 116.76
R3672 GNDA.t4 GNDA.t167 116.76
R3673 GNDA.n54 GNDA.t263 113.974
R3674 GNDA.n57 GNDA.t280 113.974
R3675 GNDA.n331 GNDA.t293 113.974
R3676 GNDA.n333 GNDA.t283 113.974
R3677 GNDA.n379 GNDA.t302 113.974
R3678 GNDA.n380 GNDA.t219 113.974
R3679 GNDA.n381 GNDA.t232 113.974
R3680 GNDA.n385 GNDA.t286 113.974
R3681 GNDA.n387 GNDA.t299 113.974
R3682 GNDA.n389 GNDA.t312 113.974
R3683 GNDA.t234 GNDA.n1828 113.624
R3684 GNDA.n1943 GNDA.t236 113.624
R3685 GNDA.t230 GNDA.n2415 113.624
R3686 GNDA.n2056 GNDA.n558 103.144
R3687 GNDA.n2291 GNDA.n145 103.144
R3688 GNDA.n2056 GNDA.n559 99.6276
R3689 GNDA.n2322 GNDA.n145 99.6276
R3690 GNDA.n2471 GNDA.n2469 99.2005
R3691 GNDA.n42 GNDA.n41 99.2005
R3692 GNDA.n1708 GNDA.n1707 98.3245
R3693 GNDA.t313 GNDA.t343 98.3245
R3694 GNDA.t71 GNDA.t125 98.3245
R3695 GNDA.n1687 GNDA.n1674 98.3245
R3696 GNDA.n2439 GNDA.n82 98.227
R3697 GNDA.n896 GNDA.n729 96.5152
R3698 GNDA.n897 GNDA.n896 96.5152
R3699 GNDA.n899 GNDA.n897 96.5152
R3700 GNDA.n899 GNDA.n898 96.5152
R3701 GNDA.n898 GNDA.n610 96.5152
R3702 GNDA.n906 GNDA.n611 96.5152
R3703 GNDA.n906 GNDA.n723 96.5152
R3704 GNDA.n913 GNDA.n723 96.5152
R3705 GNDA.n914 GNDA.n913 96.5152
R3706 GNDA.n915 GNDA.n914 96.5152
R3707 GNDA.n915 GNDA.n557 96.5152
R3708 GNDA.n2058 GNDA.n2057 96.5152
R3709 GNDA.n2058 GNDA.n553 96.5152
R3710 GNDA.n2064 GNDA.n553 96.5152
R3711 GNDA.n2065 GNDA.n2064 96.5152
R3712 GNDA.n2066 GNDA.n2065 96.5152
R3713 GNDA.n2076 GNDA.n2075 96.5152
R3714 GNDA.n2076 GNDA.n539 96.5152
R3715 GNDA.n2083 GNDA.n539 96.5152
R3716 GNDA.n2084 GNDA.n2083 96.5152
R3717 GNDA.n2085 GNDA.n2084 96.5152
R3718 GNDA.n2085 GNDA.n535 96.5152
R3719 GNDA.n2093 GNDA.n2092 96.5152
R3720 GNDA.n2093 GNDA.n530 96.5152
R3721 GNDA.n2099 GNDA.n530 96.5152
R3722 GNDA.n2100 GNDA.n2099 96.5152
R3723 GNDA.n2101 GNDA.n2100 96.5152
R3724 GNDA.n2107 GNDA.n526 96.5152
R3725 GNDA.n2108 GNDA.n2107 96.5152
R3726 GNDA.n2110 GNDA.n2108 96.5152
R3727 GNDA.n2110 GNDA.n2109 96.5152
R3728 GNDA.n2109 GNDA.n317 96.5152
R3729 GNDA.n2171 GNDA.n485 95.4985
R3730 GNDA.n2439 GNDA.n85 95.4038
R3731 GNDA.n418 GNDA.n417 94.8175
R3732 GNDA.n416 GNDA.n415 94.8175
R3733 GNDA.n414 GNDA.n413 94.8175
R3734 GNDA.n412 GNDA.n411 94.8175
R3735 GNDA.n410 GNDA.n409 94.8175
R3736 GNDA.n408 GNDA.n407 94.8175
R3737 GNDA.n406 GNDA.n405 94.8175
R3738 GNDA.n404 GNDA.n403 94.8175
R3739 GNDA.n402 GNDA.n401 94.8175
R3740 GNDA.n400 GNDA.n399 94.8175
R3741 GNDA.n398 GNDA.n397 94.8175
R3742 GNDA.t45 GNDA.t256 92.7208
R3743 GNDA.t89 GNDA.t146 92.7208
R3744 GNDA.t347 GNDA.t0 92.7208
R3745 GNDA.t20 GNDA.t151 92.7208
R3746 GNDA.t301 GNDA.t182 92.7208
R3747 GNDA.t182 GNDA.t108 92.7208
R3748 GNDA.t318 GNDA.t154 92.7208
R3749 GNDA.t340 GNDA.t119 92.7208
R3750 GNDA.t119 GNDA.t15 92.7208
R3751 GNDA.t15 GNDA.t100 92.7208
R3752 GNDA.t73 GNDA.t285 92.7208
R3753 GNDA.t285 GNDA.t61 92.7208
R3754 GNDA.t61 GNDA.t92 92.7208
R3755 GNDA.t160 GNDA.t181 92.7208
R3756 GNDA.t311 GNDA.t314 92.7208
R3757 GNDA.t192 GNDA.t121 92.7208
R3758 GNDA.t157 GNDA.t86 92.7208
R3759 GNDA.t158 GNDA.t87 92.7208
R3760 GNDA.t259 GNDA.t199 92.7208
R3761 GNDA.t17 GNDA.t304 92.1793
R3762 GNDA.t345 GNDA.t185 92.1793
R3763 GNDA.t194 GNDA.t107 92.1793
R3764 GNDA.t159 GNDA.t271 92.1793
R3765 GNDA.t236 GNDA.n559 91.423
R3766 GNDA.n2322 GNDA.t230 91.423
R3767 GNDA.n424 GNDA.n423 90.6469
R3768 GNDA.n472 GNDA.n469 90.6469
R3769 GNDA.n395 GNDA.t250 90.6175
R3770 GNDA.n32 GNDA.t290 90.6175
R3771 GNDA.n422 GNDA.n421 90.3344
R3772 GNDA.n471 GNDA.n470 90.3344
R3773 GNDA.t140 GNDA.t307 88.5063
R3774 GNDA.t200 GNDA.t253 88.5063
R3775 GNDA.n442 GNDA.n440 85.6005
R3776 GNDA.n1695 GNDA.n1694 85.2845
R3777 GNDA.n1628 GNDA.n1627 85.2845
R3778 GNDA.n544 GNDA.n543 84.306
R3779 GNDA.t224 GNDA.t45 80.0771
R3780 GNDA.t69 GNDA.t140 80.0771
R3781 GNDA.n2488 GNDA.t314 80.0771
R3782 GNDA.t155 GNDA.t200 80.0771
R3783 GNDA.t199 GNDA.t242 80.0771
R3784 GNDA.t206 GNDA.t114 79.8888
R3785 GNDA.t136 GNDA.t23 79.8888
R3786 GNDA.t112 GNDA.t54 79.8888
R3787 GNDA.t95 GNDA.t27 79.8888
R3788 GNDA.n2281 GNDA.n2280 76.3222
R3789 GNDA.n292 GNDA.n291 76.3222
R3790 GNDA.n2270 GNDA.n2269 76.3222
R3791 GNDA.n301 GNDA.n300 76.3222
R3792 GNDA.n2259 GNDA.n2258 76.3222
R3793 GNDA.n2186 GNDA.n306 76.3222
R3794 GNDA.n2181 GNDA.n307 76.3222
R3795 GNDA.n2297 GNDA.n2296 76.3222
R3796 GNDA.n2302 GNDA.n2301 76.3222
R3797 GNDA.n2305 GNDA.n2304 76.3222
R3798 GNDA.n2310 GNDA.n2309 76.3222
R3799 GNDA.n2313 GNDA.n2312 76.3222
R3800 GNDA.n2318 GNDA.n2317 76.3222
R3801 GNDA.n2295 GNDA.n150 76.3222
R3802 GNDA.n259 GNDA.n151 76.3222
R3803 GNDA.n264 GNDA.n152 76.3222
R3804 GNDA.n270 GNDA.n153 76.3222
R3805 GNDA.n2284 GNDA.n154 76.3222
R3806 GNDA.n2285 GNDA.n149 76.3222
R3807 GNDA.n112 GNDA.n110 76.3222
R3808 GNDA.n255 GNDA.n254 76.3222
R3809 GNDA.n252 GNDA.n210 76.3222
R3810 GNDA.n248 GNDA.n247 76.3222
R3811 GNDA.n241 GNDA.n212 76.3222
R3812 GNDA.n240 GNDA.n239 76.3222
R3813 GNDA.n233 GNDA.n214 76.3222
R3814 GNDA.n1213 GNDA.n162 76.3222
R3815 GNDA.n1215 GNDA.n163 76.3222
R3816 GNDA.n1217 GNDA.n164 76.3222
R3817 GNDA.n1219 GNDA.n165 76.3222
R3818 GNDA.n2324 GNDA.n146 76.3222
R3819 GNDA.n1239 GNDA.n204 76.3222
R3820 GNDA.n1235 GNDA.n203 76.3222
R3821 GNDA.n1231 GNDA.n202 76.3222
R3822 GNDA.n1227 GNDA.n201 76.3222
R3823 GNDA.n1223 GNDA.n200 76.3222
R3824 GNDA.n2016 GNDA.n199 76.3222
R3825 GNDA.n1262 GNDA.n575 76.3222
R3826 GNDA.n1209 GNDA.n1208 76.3222
R3827 GNDA.n1256 GNDA.n1207 76.3222
R3828 GNDA.n1252 GNDA.n1206 76.3222
R3829 GNDA.n1248 GNDA.n1205 76.3222
R3830 GNDA.n1244 GNDA.n1204 76.3222
R3831 GNDA.n1900 GNDA.n1898 76.3222
R3832 GNDA.n1908 GNDA.n571 76.3222
R3833 GNDA.n1913 GNDA.n1910 76.3222
R3834 GNDA.n1911 GNDA.n565 76.3222
R3835 GNDA.n1924 GNDA.n562 76.3222
R3836 GNDA.n1382 GNDA.n1381 76.3222
R3837 GNDA.n1273 GNDA.n1272 76.3222
R3838 GNDA.n1371 GNDA.n1370 76.3222
R3839 GNDA.n1282 GNDA.n1281 76.3222
R3840 GNDA.n1360 GNDA.n1359 76.3222
R3841 GNDA.n1287 GNDA.n1286 76.3222
R3842 GNDA.n2293 GNDA.n2292 76.3222
R3843 GNDA.n260 GNDA.n192 76.3222
R3844 GNDA.n266 GNDA.n191 76.3222
R3845 GNDA.n272 GNDA.n190 76.3222
R3846 GNDA.n278 GNDA.n189 76.3222
R3847 GNDA.n2289 GNDA.n188 76.3222
R3848 GNDA.n679 GNDA.n678 76.3222
R3849 GNDA.n674 GNDA.n654 76.3222
R3850 GNDA.n671 GNDA.n653 76.3222
R3851 GNDA.n667 GNDA.n652 76.3222
R3852 GNDA.n663 GNDA.n651 76.3222
R3853 GNDA.n659 GNDA.n650 76.3222
R3854 GNDA.n628 GNDA.n627 76.3222
R3855 GNDA.n633 GNDA.n632 76.3222
R3856 GNDA.n636 GNDA.n635 76.3222
R3857 GNDA.n641 GNDA.n640 76.3222
R3858 GNDA.n644 GNDA.n643 76.3222
R3859 GNDA.n649 GNDA.n647 76.3222
R3860 GNDA.n1894 GNDA.n1893 76.3222
R3861 GNDA.n1903 GNDA.n1902 76.3222
R3862 GNDA.n1906 GNDA.n1905 76.3222
R3863 GNDA.n1916 GNDA.n1915 76.3222
R3864 GNDA.n1919 GNDA.n1918 76.3222
R3865 GNDA.n1808 GNDA.n567 76.3222
R3866 GNDA.n1869 GNDA.n1868 76.3222
R3867 GNDA.n1874 GNDA.n1873 76.3222
R3868 GNDA.n1877 GNDA.n1876 76.3222
R3869 GNDA.n1882 GNDA.n1881 76.3222
R3870 GNDA.n1885 GNDA.n1884 76.3222
R3871 GNDA.n1890 GNDA.n1889 76.3222
R3872 GNDA.n1847 GNDA.n1846 76.3222
R3873 GNDA.n1447 GNDA.n1446 76.3222
R3874 GNDA.n1480 GNDA.n1479 76.3222
R3875 GNDA.n1456 GNDA.n1455 76.3222
R3876 GNDA.n1469 GNDA.n1468 76.3222
R3877 GNDA.n1457 GNDA.n1389 76.3222
R3878 GNDA.n1542 GNDA.n1541 76.3222
R3879 GNDA.n1567 GNDA.n625 76.3222
R3880 GNDA.n1563 GNDA.n1562 76.3222
R3881 GNDA.n1556 GNDA.n630 76.3222
R3882 GNDA.n1555 GNDA.n1554 76.3222
R3883 GNDA.n1548 GNDA.n638 76.3222
R3884 GNDA.n1547 GNDA.n1546 76.3222
R3885 GNDA.n1592 GNDA.n1591 76.3222
R3886 GNDA.n1587 GNDA.n619 76.3222
R3887 GNDA.n1584 GNDA.n618 76.3222
R3888 GNDA.n1580 GNDA.n617 76.3222
R3889 GNDA.n1576 GNDA.n616 76.3222
R3890 GNDA.n1572 GNDA.n615 76.3222
R3891 GNDA.n1442 GNDA.n1410 76.3222
R3892 GNDA.n867 GNDA.n866 76.3222
R3893 GNDA.n753 GNDA.n752 76.3222
R3894 GNDA.n856 GNDA.n855 76.3222
R3895 GNDA.n762 GNDA.n761 76.3222
R3896 GNDA.n845 GNDA.n844 76.3222
R3897 GNDA.n772 GNDA.n767 76.3222
R3898 GNDA.n870 GNDA.n869 76.3222
R3899 GNDA.n919 GNDA.n918 76.3222
R3900 GNDA.n928 GNDA.n927 76.3222
R3901 GNDA.n931 GNDA.n930 76.3222
R3902 GNDA.n942 GNDA.n941 76.3222
R3903 GNDA.n945 GNDA.n944 76.3222
R3904 GNDA.n769 GNDA.n711 76.3222
R3905 GNDA.n984 GNDA.n681 76.3222
R3906 GNDA.n981 GNDA.n682 76.3222
R3907 GNDA.n971 GNDA.n683 76.3222
R3908 GNDA.n968 GNDA.n684 76.3222
R3909 GNDA.n689 GNDA.n685 76.3222
R3910 GNDA.n1202 GNDA.n1201 76.3222
R3911 GNDA.n923 GNDA.n922 76.3222
R3912 GNDA.n924 GNDA.n715 76.3222
R3913 GNDA.n935 GNDA.n934 76.3222
R3914 GNDA.n938 GNDA.n937 76.3222
R3915 GNDA.n948 GNDA.n708 76.3222
R3916 GNDA.n951 GNDA.n950 76.3222
R3917 GNDA.n2088 GNDA.n198 76.3222
R3918 GNDA.n1049 GNDA.n197 76.3222
R3919 GNDA.n1055 GNDA.n196 76.3222
R3920 GNDA.n1061 GNDA.n195 76.3222
R3921 GNDA.n1067 GNDA.n194 76.3222
R3922 GNDA.n1045 GNDA.n193 76.3222
R3923 GNDA.n1846 GNDA.n598 76.3222
R3924 GNDA.n1868 GNDA.n584 76.3222
R3925 GNDA.n1875 GNDA.n1874 76.3222
R3926 GNDA.n1876 GNDA.n582 76.3222
R3927 GNDA.n1883 GNDA.n1882 76.3222
R3928 GNDA.n1884 GNDA.n580 76.3222
R3929 GNDA.n1891 GNDA.n1890 76.3222
R3930 GNDA.n1592 GNDA.n620 76.3222
R3931 GNDA.n1585 GNDA.n619 76.3222
R3932 GNDA.n1581 GNDA.n618 76.3222
R3933 GNDA.n1577 GNDA.n617 76.3222
R3934 GNDA.n1573 GNDA.n616 76.3222
R3935 GNDA.n1569 GNDA.n615 76.3222
R3936 GNDA.n936 GNDA.n708 76.3222
R3937 GNDA.n939 GNDA.n938 76.3222
R3938 GNDA.n934 GNDA.n933 76.3222
R3939 GNDA.n925 GNDA.n924 76.3222
R3940 GNDA.n922 GNDA.n921 76.3222
R3941 GNDA.n643 GNDA.n642 76.3222
R3942 GNDA.n640 GNDA.n639 76.3222
R3943 GNDA.n635 GNDA.n634 76.3222
R3944 GNDA.n632 GNDA.n631 76.3222
R3945 GNDA.n627 GNDA.n626 76.3222
R3946 GNDA.n1923 GNDA.n1922 76.3222
R3947 GNDA.n1912 GNDA.n1911 76.3222
R3948 GNDA.n1910 GNDA.n1909 76.3222
R3949 GNDA.n1899 GNDA.n571 76.3222
R3950 GNDA.n1898 GNDA.n1897 76.3222
R3951 GNDA.n918 GNDA.n717 76.3222
R3952 GNDA.n929 GNDA.n928 76.3222
R3953 GNDA.n930 GNDA.n713 76.3222
R3954 GNDA.n943 GNDA.n942 76.3222
R3955 GNDA.n946 GNDA.n945 76.3222
R3956 GNDA.n1564 GNDA.n625 76.3222
R3957 GNDA.n1562 GNDA.n1561 76.3222
R3958 GNDA.n1557 GNDA.n1556 76.3222
R3959 GNDA.n1554 GNDA.n1553 76.3222
R3960 GNDA.n1549 GNDA.n1548 76.3222
R3961 GNDA.n1893 GNDA.n573 76.3222
R3962 GNDA.n1904 GNDA.n1903 76.3222
R3963 GNDA.n1905 GNDA.n569 76.3222
R3964 GNDA.n1917 GNDA.n1916 76.3222
R3965 GNDA.n1920 GNDA.n1919 76.3222
R3966 GNDA.n1809 GNDA.n1808 76.3222
R3967 GNDA.n1262 GNDA.n1261 76.3222
R3968 GNDA.n1257 GNDA.n1208 76.3222
R3969 GNDA.n1253 GNDA.n1207 76.3222
R3970 GNDA.n1249 GNDA.n1206 76.3222
R3971 GNDA.n1245 GNDA.n1205 76.3222
R3972 GNDA.n1241 GNDA.n1204 76.3222
R3973 GNDA.n679 GNDA.n655 76.3222
R3974 GNDA.n672 GNDA.n654 76.3222
R3975 GNDA.n668 GNDA.n653 76.3222
R3976 GNDA.n664 GNDA.n652 76.3222
R3977 GNDA.n660 GNDA.n651 76.3222
R3978 GNDA.n656 GNDA.n650 76.3222
R3979 GNDA.n2323 GNDA.n148 76.3222
R3980 GNDA.n1218 GNDA.n165 76.3222
R3981 GNDA.n1216 GNDA.n164 76.3222
R3982 GNDA.n1214 GNDA.n163 76.3222
R3983 GNDA.n1212 GNDA.n162 76.3222
R3984 GNDA.n1236 GNDA.n204 76.3222
R3985 GNDA.n1232 GNDA.n203 76.3222
R3986 GNDA.n1228 GNDA.n202 76.3222
R3987 GNDA.n1224 GNDA.n201 76.3222
R3988 GNDA.n1220 GNDA.n200 76.3222
R3989 GNDA.n2016 GNDA.n205 76.3222
R3990 GNDA.n1192 GNDA.n1191 76.3222
R3991 GNDA.n1080 GNDA.n1073 76.3222
R3992 GNDA.n1181 GNDA.n1180 76.3222
R3993 GNDA.n1089 GNDA.n1082 76.3222
R3994 GNDA.n1170 GNDA.n1169 76.3222
R3995 GNDA.n1095 GNDA.n1091 76.3222
R3996 GNDA.n2143 GNDA.n2142 76.3222
R3997 GNDA.n2090 GNDA.n156 76.3222
R3998 GNDA.n1047 GNDA.n157 76.3222
R3999 GNDA.n1053 GNDA.n158 76.3222
R4000 GNDA.n1059 GNDA.n159 76.3222
R4001 GNDA.n1065 GNDA.n160 76.3222
R4002 GNDA.n1195 GNDA.n155 76.3222
R4003 GNDA.n1194 GNDA.n160 76.3222
R4004 GNDA.n1064 GNDA.n159 76.3222
R4005 GNDA.n1058 GNDA.n158 76.3222
R4006 GNDA.n1052 GNDA.n157 76.3222
R4007 GNDA.n1046 GNDA.n156 76.3222
R4008 GNDA.n1048 GNDA.n198 76.3222
R4009 GNDA.n1054 GNDA.n197 76.3222
R4010 GNDA.n1060 GNDA.n196 76.3222
R4011 GNDA.n1066 GNDA.n195 76.3222
R4012 GNDA.n1069 GNDA.n194 76.3222
R4013 GNDA.n1071 GNDA.n155 76.3222
R4014 GNDA.n1096 GNDA.n1095 76.3222
R4015 GNDA.n1169 GNDA.n1168 76.3222
R4016 GNDA.n1090 GNDA.n1089 76.3222
R4017 GNDA.n1180 GNDA.n1179 76.3222
R4018 GNDA.n1081 GNDA.n1080 76.3222
R4019 GNDA.n1191 GNDA.n1190 76.3222
R4020 GNDA.n950 GNDA.n949 76.3222
R4021 GNDA.n1202 GNDA.n686 76.3222
R4022 GNDA.n967 GNDA.n685 76.3222
R4023 GNDA.n972 GNDA.n684 76.3222
R4024 GNDA.n980 GNDA.n683 76.3222
R4025 GNDA.n985 GNDA.n682 76.3222
R4026 GNDA.n952 GNDA.n681 76.3222
R4027 GNDA.n1045 GNDA.n206 76.3222
R4028 GNDA.n871 GNDA.n870 76.3222
R4029 GNDA.n767 GNDA.n763 76.3222
R4030 GNDA.n846 GNDA.n845 76.3222
R4031 GNDA.n761 GNDA.n754 76.3222
R4032 GNDA.n857 GNDA.n856 76.3222
R4033 GNDA.n752 GNDA.n744 76.3222
R4034 GNDA.n868 GNDA.n867 76.3222
R4035 GNDA.n770 GNDA.n769 76.3222
R4036 GNDA.n276 GNDA.n154 76.3222
R4037 GNDA.n275 GNDA.n153 76.3222
R4038 GNDA.n269 GNDA.n152 76.3222
R4039 GNDA.n263 GNDA.n151 76.3222
R4040 GNDA.n258 GNDA.n150 76.3222
R4041 GNDA.n2292 GNDA.n186 76.3222
R4042 GNDA.n265 GNDA.n192 76.3222
R4043 GNDA.n271 GNDA.n191 76.3222
R4044 GNDA.n277 GNDA.n190 76.3222
R4045 GNDA.n280 GNDA.n189 76.3222
R4046 GNDA.n2296 GNDA.n181 76.3222
R4047 GNDA.n2303 GNDA.n2302 76.3222
R4048 GNDA.n2304 GNDA.n179 76.3222
R4049 GNDA.n2311 GNDA.n2310 76.3222
R4050 GNDA.n2312 GNDA.n177 76.3222
R4051 GNDA.n2319 GNDA.n2318 76.3222
R4052 GNDA.n282 GNDA.n149 76.3222
R4053 GNDA.n647 GNDA.n646 76.3222
R4054 GNDA.n1286 GNDA.n1283 76.3222
R4055 GNDA.n1361 GNDA.n1360 76.3222
R4056 GNDA.n1281 GNDA.n1274 76.3222
R4057 GNDA.n1372 GNDA.n1371 76.3222
R4058 GNDA.n1272 GNDA.n1265 76.3222
R4059 GNDA.n1383 GNDA.n1382 76.3222
R4060 GNDA.n2290 GNDA.n2289 76.3222
R4061 GNDA.n1442 GNDA.n1441 76.3222
R4062 GNDA.n1541 GNDA.n1540 76.3222
R4063 GNDA.n1458 GNDA.n1457 76.3222
R4064 GNDA.n1470 GNDA.n1469 76.3222
R4065 GNDA.n1455 GNDA.n1448 76.3222
R4066 GNDA.n1481 GNDA.n1480 76.3222
R4067 GNDA.n1446 GNDA.n1445 76.3222
R4068 GNDA.n1546 GNDA.n1387 76.3222
R4069 GNDA.n306 GNDA.n302 76.3222
R4070 GNDA.n2260 GNDA.n2259 76.3222
R4071 GNDA.n300 GNDA.n293 76.3222
R4072 GNDA.n2271 GNDA.n2270 76.3222
R4073 GNDA.n291 GNDA.n284 76.3222
R4074 GNDA.n2282 GNDA.n2281 76.3222
R4075 GNDA.n254 GNDA.n253 76.3222
R4076 GNDA.n249 GNDA.n210 76.3222
R4077 GNDA.n247 GNDA.n246 76.3222
R4078 GNDA.n242 GNDA.n241 76.3222
R4079 GNDA.n239 GNDA.n238 76.3222
R4080 GNDA.n234 GNDA.n233 76.3222
R4081 GNDA.n2142 GNDA.n513 76.3222
R4082 GNDA.n2184 GNDA.n307 76.3222
R4083 GNDA.n110 GNDA.n92 76.3222
R4084 GNDA.n1501 GNDA.n1401 76.062
R4085 GNDA.n1502 GNDA.n1501 76.062
R4086 GNDA.n1322 GNDA.n1321 76.062
R4087 GNDA.n1321 GNDA.n1320 76.062
R4088 GNDA.n2221 GNDA.n2220 76.062
R4089 GNDA.n2220 GNDA.n2219 76.062
R4090 GNDA.n807 GNDA.n806 76.062
R4091 GNDA.n806 GNDA.n805 76.062
R4092 GNDA.n1007 GNDA.n1006 76.062
R4093 GNDA.n1006 GNDA.n1005 76.062
R4094 GNDA.n1131 GNDA.n1130 76.062
R4095 GNDA.n1130 GNDA.n1129 76.062
R4096 GNDA.n1770 GNDA.n1749 76.062
R4097 GNDA.n1771 GNDA.n1770 76.062
R4098 GNDA.n1979 GNDA.n1960 76.062
R4099 GNDA.n1980 GNDA.n1979 76.062
R4100 GNDA.n2366 GNDA.n2365 76.062
R4101 GNDA.n2365 GNDA.n2364 76.062
R4102 GNDA.n1485 GNDA.n1484 74.5978
R4103 GNDA.n1486 GNDA.n1485 74.5978
R4104 GNDA.n1378 GNDA.n1267 74.5978
R4105 GNDA.n1305 GNDA.n1267 74.5978
R4106 GNDA.n2277 GNDA.n286 74.5978
R4107 GNDA.n2204 GNDA.n286 74.5978
R4108 GNDA.n863 GNDA.n747 74.5978
R4109 GNDA.n790 GNDA.n747 74.5978
R4110 GNDA.n989 GNDA.n988 74.5978
R4111 GNDA.n990 GNDA.n989 74.5978
R4112 GNDA.n1187 GNDA.n1075 74.5978
R4113 GNDA.n1114 GNDA.n1075 74.5978
R4114 GNDA.n1754 GNDA.n606 74.5978
R4115 GNDA.n1755 GNDA.n1754 74.5978
R4116 GNDA.n2049 GNDA.n1928 74.5978
R4117 GNDA.n1964 GNDA.n1928 74.5978
R4118 GNDA.n2348 GNDA.n2347 74.5978
R4119 GNDA.n2349 GNDA.n2348 74.5978
R4120 GNDA.n1700 GNDA.t207 73.7435
R4121 GNDA.n1716 GNDA.t34 73.7435
R4122 GNDA.n1716 GNDA.t205 73.7435
R4123 GNDA.n1641 GNDA.t212 73.7435
R4124 GNDA.n1641 GNDA.t99 73.7435
R4125 GNDA.n1691 GNDA.t166 73.7435
R4126 GNDA.n2430 GNDA.n94 73.1246
R4127 GNDA.n2460 GNDA.t72 72.3996
R4128 GNDA.n2446 GNDA.t333 72.3996
R4129 GNDA.n484 GNDA.t344 72.3996
R4130 GNDA.t150 GNDA.n344 72.3996
R4131 GNDA.t108 GNDA.n378 71.648
R4132 GNDA.t114 GNDA.t204 67.5983
R4133 GNDA.t204 GNDA.t136 67.5983
R4134 GNDA.t175 GNDA.n1725 67.5983
R4135 GNDA.n1725 GNDA.t173 67.5983
R4136 GNDA.t79 GNDA.t112 67.5983
R4137 GNDA.t27 GNDA.t79 67.5983
R4138 GNDA.n1491 GNDA.t233 65.8183
R4139 GNDA.n1493 GNDA.t233 65.8183
R4140 GNDA.n1499 GNDA.t233 65.8183
R4141 GNDA.n1507 GNDA.t233 65.8183
R4142 GNDA.n1509 GNDA.t233 65.8183
R4143 GNDA.n1515 GNDA.t233 65.8183
R4144 GNDA.n1517 GNDA.t233 65.8183
R4145 GNDA.n1535 GNDA.t233 65.8183
R4146 GNDA.n1532 GNDA.t233 65.8183
R4147 GNDA.n1526 GNDA.t233 65.8183
R4148 GNDA.n1523 GNDA.t233 65.8183
R4149 GNDA.n1307 GNDA.t235 65.8183
R4150 GNDA.n1313 GNDA.t235 65.8183
R4151 GNDA.n1315 GNDA.t235 65.8183
R4152 GNDA.n1323 GNDA.t235 65.8183
R4153 GNDA.n1329 GNDA.t235 65.8183
R4154 GNDA.n1331 GNDA.t235 65.8183
R4155 GNDA.n1337 GNDA.t235 65.8183
R4156 GNDA.n1354 GNDA.t235 65.8183
R4157 GNDA.n1348 GNDA.t235 65.8183
R4158 GNDA.n1346 GNDA.t235 65.8183
R4159 GNDA.n1340 GNDA.t235 65.8183
R4160 GNDA.n2206 GNDA.t309 65.8183
R4161 GNDA.n2212 GNDA.t309 65.8183
R4162 GNDA.n2214 GNDA.t309 65.8183
R4163 GNDA.n2222 GNDA.t309 65.8183
R4164 GNDA.n2228 GNDA.t309 65.8183
R4165 GNDA.n2230 GNDA.t309 65.8183
R4166 GNDA.n2236 GNDA.t309 65.8183
R4167 GNDA.n2253 GNDA.t309 65.8183
R4168 GNDA.n2247 GNDA.t309 65.8183
R4169 GNDA.n2245 GNDA.t309 65.8183
R4170 GNDA.n2239 GNDA.t309 65.8183
R4171 GNDA.n792 GNDA.t277 65.8183
R4172 GNDA.n798 GNDA.t277 65.8183
R4173 GNDA.n800 GNDA.t277 65.8183
R4174 GNDA.n808 GNDA.t277 65.8183
R4175 GNDA.n814 GNDA.t277 65.8183
R4176 GNDA.n816 GNDA.t277 65.8183
R4177 GNDA.n822 GNDA.t277 65.8183
R4178 GNDA.n839 GNDA.t277 65.8183
R4179 GNDA.n833 GNDA.t277 65.8183
R4180 GNDA.n831 GNDA.t277 65.8183
R4181 GNDA.n825 GNDA.t277 65.8183
R4182 GNDA.n992 GNDA.t276 65.8183
R4183 GNDA.n998 GNDA.t276 65.8183
R4184 GNDA.n1000 GNDA.t276 65.8183
R4185 GNDA.n1008 GNDA.t276 65.8183
R4186 GNDA.n1014 GNDA.t276 65.8183
R4187 GNDA.n1016 GNDA.t276 65.8183
R4188 GNDA.n1022 GNDA.t276 65.8183
R4189 GNDA.n1039 GNDA.t276 65.8183
R4190 GNDA.n1033 GNDA.t276 65.8183
R4191 GNDA.n1031 GNDA.t276 65.8183
R4192 GNDA.n1025 GNDA.t276 65.8183
R4193 GNDA.n1116 GNDA.t251 65.8183
R4194 GNDA.n1122 GNDA.t251 65.8183
R4195 GNDA.n1124 GNDA.t251 65.8183
R4196 GNDA.n1132 GNDA.t251 65.8183
R4197 GNDA.n1138 GNDA.t251 65.8183
R4198 GNDA.n1140 GNDA.t251 65.8183
R4199 GNDA.n1146 GNDA.t251 65.8183
R4200 GNDA.n1163 GNDA.t251 65.8183
R4201 GNDA.n1157 GNDA.t251 65.8183
R4202 GNDA.n1155 GNDA.t251 65.8183
R4203 GNDA.n1149 GNDA.t251 65.8183
R4204 GNDA.n1760 GNDA.t244 65.8183
R4205 GNDA.n1762 GNDA.t244 65.8183
R4206 GNDA.n1768 GNDA.t244 65.8183
R4207 GNDA.n1776 GNDA.t244 65.8183
R4208 GNDA.n1778 GNDA.t244 65.8183
R4209 GNDA.n1784 GNDA.t244 65.8183
R4210 GNDA.n1786 GNDA.t244 65.8183
R4211 GNDA.n1804 GNDA.t244 65.8183
R4212 GNDA.n1801 GNDA.t244 65.8183
R4213 GNDA.n1795 GNDA.t244 65.8183
R4214 GNDA.n1792 GNDA.t244 65.8183
R4215 GNDA.n1969 GNDA.t240 65.8183
R4216 GNDA.n1971 GNDA.t240 65.8183
R4217 GNDA.n1977 GNDA.t240 65.8183
R4218 GNDA.n1985 GNDA.t240 65.8183
R4219 GNDA.n1987 GNDA.t240 65.8183
R4220 GNDA.n1993 GNDA.t240 65.8183
R4221 GNDA.n1995 GNDA.t240 65.8183
R4222 GNDA.n2013 GNDA.t240 65.8183
R4223 GNDA.n2010 GNDA.t240 65.8183
R4224 GNDA.n2004 GNDA.t240 65.8183
R4225 GNDA.n2001 GNDA.t240 65.8183
R4226 GNDA.n2351 GNDA.t229 65.8183
R4227 GNDA.n2357 GNDA.t229 65.8183
R4228 GNDA.n2359 GNDA.t229 65.8183
R4229 GNDA.n2367 GNDA.t229 65.8183
R4230 GNDA.n2373 GNDA.t229 65.8183
R4231 GNDA.n2375 GNDA.t229 65.8183
R4232 GNDA.n2381 GNDA.t229 65.8183
R4233 GNDA.n2398 GNDA.t229 65.8183
R4234 GNDA.n2392 GNDA.t229 65.8183
R4235 GNDA.n2390 GNDA.t229 65.8183
R4236 GNDA.n2384 GNDA.t229 65.8183
R4237 GNDA.n2401 GNDA.t229 65.8183
R4238 GNDA.n2410 GNDA.t229 65.8183
R4239 GNDA.n2336 GNDA.t229 65.8183
R4240 GNDA.n2334 GNDA.t229 65.8183
R4241 GNDA.n1950 GNDA.t240 65.8183
R4242 GNDA.n2032 GNDA.t240 65.8183
R4243 GNDA.n1936 GNDA.t240 65.8183
R4244 GNDA.n2047 GNDA.t240 65.8183
R4245 GNDA.n1739 GNDA.t244 65.8183
R4246 GNDA.n1823 GNDA.t244 65.8183
R4247 GNDA.n1599 GNDA.t244 65.8183
R4248 GNDA.n1835 GNDA.t244 65.8183
R4249 GNDA.n1093 GNDA.t251 65.8183
R4250 GNDA.n1174 GNDA.t251 65.8183
R4251 GNDA.n1084 GNDA.t251 65.8183
R4252 GNDA.n1185 GNDA.t251 65.8183
R4253 GNDA.t276 GNDA.n691 65.8183
R4254 GNDA.n962 GNDA.t276 65.8183
R4255 GNDA.n976 GNDA.t276 65.8183
R4256 GNDA.n958 GNDA.t276 65.8183
R4257 GNDA.n765 GNDA.t277 65.8183
R4258 GNDA.n850 GNDA.t277 65.8183
R4259 GNDA.n756 GNDA.t277 65.8183
R4260 GNDA.n861 GNDA.t277 65.8183
R4261 GNDA.n304 GNDA.t309 65.8183
R4262 GNDA.n2264 GNDA.t309 65.8183
R4263 GNDA.n295 GNDA.t309 65.8183
R4264 GNDA.n2275 GNDA.t309 65.8183
R4265 GNDA.n1285 GNDA.t235 65.8183
R4266 GNDA.n1365 GNDA.t235 65.8183
R4267 GNDA.n1276 GNDA.t235 65.8183
R4268 GNDA.n1376 GNDA.t235 65.8183
R4269 GNDA.n1463 GNDA.t233 65.8183
R4270 GNDA.n1460 GNDA.t233 65.8183
R4271 GNDA.n1474 GNDA.t233 65.8183
R4272 GNDA.n1450 GNDA.t233 65.8183
R4273 GNDA.n102 GNDA.n82 65.4848
R4274 GNDA.t234 GNDA.n610 65.4161
R4275 GNDA.n2066 GNDA.t236 65.4161
R4276 GNDA.n2101 GNDA.t230 65.4161
R4277 GNDA.t134 GNDA.t89 63.2189
R4278 GNDA.t52 GNDA.t20 63.2189
R4279 GNDA.t50 GNDA.t192 63.2189
R4280 GNDA.t87 GNDA.t326 63.2189
R4281 GNDA.t205 GNDA.n1715 61.453
R4282 GNDA.t212 GNDA.n1640 61.453
R4283 GNDA.n2441 GNDA.n82 61.1116
R4284 GNDA.t234 GNDA.n577 60.9488
R4285 GNDA.t236 GNDA.n187 60.9488
R4286 GNDA.t304 GNDA.t206 55.3078
R4287 GNDA.t23 GNDA.t345 55.3078
R4288 GNDA.n1714 GNDA.t238 55.3078
R4289 GNDA.n1639 GNDA.t265 55.3078
R4290 GNDA.t54 GNDA.t194 55.3078
R4291 GNDA.t271 GNDA.t95 55.3078
R4292 GNDA.n2348 GNDA.t229 55.2026
R4293 GNDA.t240 GNDA.n1928 55.2026
R4294 GNDA.n1754 GNDA.t244 55.2026
R4295 GNDA.t251 GNDA.n1075 55.2026
R4296 GNDA.n989 GNDA.t276 55.2026
R4297 GNDA.t277 GNDA.n747 55.2026
R4298 GNDA.t309 GNDA.n286 55.2026
R4299 GNDA.t235 GNDA.n1267 55.2026
R4300 GNDA.n1485 GNDA.t233 55.2026
R4301 GNDA.n511 GNDA.n172 55.1165
R4302 GNDA.n2183 GNDA.n169 55.1165
R4303 GNDA.n2431 GNDA.n93 55.1165
R4304 GNDA.n458 GNDA.t330 54.7898
R4305 GNDA.n427 GNDA.t33 54.7898
R4306 GNDA.n1501 GNDA.t233 54.4705
R4307 GNDA.n1321 GNDA.t235 54.4705
R4308 GNDA.n2220 GNDA.t309 54.4705
R4309 GNDA.n806 GNDA.t277 54.4705
R4310 GNDA.n1006 GNDA.t276 54.4705
R4311 GNDA.n1130 GNDA.t251 54.4705
R4312 GNDA.n1770 GNDA.t244 54.4705
R4313 GNDA.n1979 GNDA.t240 54.4705
R4314 GNDA.n2365 GNDA.t229 54.4705
R4315 GNDA.n365 GNDA.n358 54.4005
R4316 GNDA.n463 GNDA.n384 54.4005
R4317 GNDA.n382 GNDA.n52 54.4005
R4318 GNDA.n386 GNDA.n52 54.4005
R4319 GNDA.n2451 GNDA.n2450 54.4005
R4320 GNDA.n1476 GNDA.n1450 53.3664
R4321 GNDA.n1474 GNDA.n1473 53.3664
R4322 GNDA.n1465 GNDA.n1460 53.3664
R4323 GNDA.n1463 GNDA.n1392 53.3664
R4324 GNDA.n1523 GNDA.n1522 53.3664
R4325 GNDA.n1527 GNDA.n1526 53.3664
R4326 GNDA.n1532 GNDA.n1531 53.3664
R4327 GNDA.n1535 GNDA.n1534 53.3664
R4328 GNDA.n1507 GNDA.n1506 53.3664
R4329 GNDA.n1510 GNDA.n1509 53.3664
R4330 GNDA.n1515 GNDA.n1514 53.3664
R4331 GNDA.n1518 GNDA.n1517 53.3664
R4332 GNDA.n1500 GNDA.n1499 53.3664
R4333 GNDA.n1493 GNDA.n1403 53.3664
R4334 GNDA.n1492 GNDA.n1491 53.3664
R4335 GNDA.n1491 GNDA.n1490 53.3664
R4336 GNDA.n1494 GNDA.n1493 53.3664
R4337 GNDA.n1499 GNDA.n1498 53.3664
R4338 GNDA.n1508 GNDA.n1507 53.3664
R4339 GNDA.n1509 GNDA.n1399 53.3664
R4340 GNDA.n1516 GNDA.n1515 53.3664
R4341 GNDA.n1517 GNDA.n1397 53.3664
R4342 GNDA.n1536 GNDA.n1535 53.3664
R4343 GNDA.n1533 GNDA.n1532 53.3664
R4344 GNDA.n1526 GNDA.n1394 53.3664
R4345 GNDA.n1524 GNDA.n1523 53.3664
R4346 GNDA.n1376 GNDA.n1375 53.3664
R4347 GNDA.n1367 GNDA.n1276 53.3664
R4348 GNDA.n1365 GNDA.n1364 53.3664
R4349 GNDA.n1356 GNDA.n1285 53.3664
R4350 GNDA.n1340 GNDA.n1339 53.3664
R4351 GNDA.n1346 GNDA.n1345 53.3664
R4352 GNDA.n1349 GNDA.n1348 53.3664
R4353 GNDA.n1354 GNDA.n1353 53.3664
R4354 GNDA.n1324 GNDA.n1323 53.3664
R4355 GNDA.n1329 GNDA.n1328 53.3664
R4356 GNDA.n1332 GNDA.n1331 53.3664
R4357 GNDA.n1337 GNDA.n1336 53.3664
R4358 GNDA.n1315 GNDA.n1300 53.3664
R4359 GNDA.n1314 GNDA.n1313 53.3664
R4360 GNDA.n1307 GNDA.n1302 53.3664
R4361 GNDA.n1308 GNDA.n1307 53.3664
R4362 GNDA.n1313 GNDA.n1312 53.3664
R4363 GNDA.n1316 GNDA.n1315 53.3664
R4364 GNDA.n1323 GNDA.n1298 53.3664
R4365 GNDA.n1330 GNDA.n1329 53.3664
R4366 GNDA.n1331 GNDA.n1296 53.3664
R4367 GNDA.n1338 GNDA.n1337 53.3664
R4368 GNDA.n1355 GNDA.n1354 53.3664
R4369 GNDA.n1348 GNDA.n1291 53.3664
R4370 GNDA.n1347 GNDA.n1346 53.3664
R4371 GNDA.n1341 GNDA.n1340 53.3664
R4372 GNDA.n2275 GNDA.n2274 53.3664
R4373 GNDA.n2266 GNDA.n295 53.3664
R4374 GNDA.n2264 GNDA.n2263 53.3664
R4375 GNDA.n2255 GNDA.n304 53.3664
R4376 GNDA.n2239 GNDA.n2238 53.3664
R4377 GNDA.n2245 GNDA.n2244 53.3664
R4378 GNDA.n2248 GNDA.n2247 53.3664
R4379 GNDA.n2253 GNDA.n2252 53.3664
R4380 GNDA.n2223 GNDA.n2222 53.3664
R4381 GNDA.n2228 GNDA.n2227 53.3664
R4382 GNDA.n2231 GNDA.n2230 53.3664
R4383 GNDA.n2236 GNDA.n2235 53.3664
R4384 GNDA.n2214 GNDA.n2199 53.3664
R4385 GNDA.n2213 GNDA.n2212 53.3664
R4386 GNDA.n2206 GNDA.n2201 53.3664
R4387 GNDA.n2207 GNDA.n2206 53.3664
R4388 GNDA.n2212 GNDA.n2211 53.3664
R4389 GNDA.n2215 GNDA.n2214 53.3664
R4390 GNDA.n2222 GNDA.n2197 53.3664
R4391 GNDA.n2229 GNDA.n2228 53.3664
R4392 GNDA.n2230 GNDA.n2195 53.3664
R4393 GNDA.n2237 GNDA.n2236 53.3664
R4394 GNDA.n2254 GNDA.n2253 53.3664
R4395 GNDA.n2247 GNDA.n2190 53.3664
R4396 GNDA.n2246 GNDA.n2245 53.3664
R4397 GNDA.n2240 GNDA.n2239 53.3664
R4398 GNDA.n861 GNDA.n860 53.3664
R4399 GNDA.n852 GNDA.n756 53.3664
R4400 GNDA.n850 GNDA.n849 53.3664
R4401 GNDA.n841 GNDA.n765 53.3664
R4402 GNDA.n825 GNDA.n824 53.3664
R4403 GNDA.n831 GNDA.n830 53.3664
R4404 GNDA.n834 GNDA.n833 53.3664
R4405 GNDA.n839 GNDA.n838 53.3664
R4406 GNDA.n809 GNDA.n808 53.3664
R4407 GNDA.n814 GNDA.n813 53.3664
R4408 GNDA.n817 GNDA.n816 53.3664
R4409 GNDA.n822 GNDA.n821 53.3664
R4410 GNDA.n800 GNDA.n785 53.3664
R4411 GNDA.n799 GNDA.n798 53.3664
R4412 GNDA.n792 GNDA.n787 53.3664
R4413 GNDA.n793 GNDA.n792 53.3664
R4414 GNDA.n798 GNDA.n797 53.3664
R4415 GNDA.n801 GNDA.n800 53.3664
R4416 GNDA.n808 GNDA.n783 53.3664
R4417 GNDA.n815 GNDA.n814 53.3664
R4418 GNDA.n816 GNDA.n781 53.3664
R4419 GNDA.n823 GNDA.n822 53.3664
R4420 GNDA.n840 GNDA.n839 53.3664
R4421 GNDA.n833 GNDA.n776 53.3664
R4422 GNDA.n832 GNDA.n831 53.3664
R4423 GNDA.n826 GNDA.n825 53.3664
R4424 GNDA.n959 GNDA.n958 53.3664
R4425 GNDA.n976 GNDA.n975 53.3664
R4426 GNDA.n963 GNDA.n962 53.3664
R4427 GNDA.n1041 GNDA.n691 53.3664
R4428 GNDA.n1025 GNDA.n1024 53.3664
R4429 GNDA.n1031 GNDA.n1030 53.3664
R4430 GNDA.n1034 GNDA.n1033 53.3664
R4431 GNDA.n1039 GNDA.n1038 53.3664
R4432 GNDA.n1009 GNDA.n1008 53.3664
R4433 GNDA.n1014 GNDA.n1013 53.3664
R4434 GNDA.n1017 GNDA.n1016 53.3664
R4435 GNDA.n1022 GNDA.n1021 53.3664
R4436 GNDA.n1000 GNDA.n701 53.3664
R4437 GNDA.n999 GNDA.n998 53.3664
R4438 GNDA.n992 GNDA.n703 53.3664
R4439 GNDA.n993 GNDA.n992 53.3664
R4440 GNDA.n998 GNDA.n997 53.3664
R4441 GNDA.n1001 GNDA.n1000 53.3664
R4442 GNDA.n1008 GNDA.n699 53.3664
R4443 GNDA.n1015 GNDA.n1014 53.3664
R4444 GNDA.n1016 GNDA.n697 53.3664
R4445 GNDA.n1023 GNDA.n1022 53.3664
R4446 GNDA.n1040 GNDA.n1039 53.3664
R4447 GNDA.n1033 GNDA.n692 53.3664
R4448 GNDA.n1032 GNDA.n1031 53.3664
R4449 GNDA.n1026 GNDA.n1025 53.3664
R4450 GNDA.n1185 GNDA.n1184 53.3664
R4451 GNDA.n1176 GNDA.n1084 53.3664
R4452 GNDA.n1174 GNDA.n1173 53.3664
R4453 GNDA.n1165 GNDA.n1093 53.3664
R4454 GNDA.n1149 GNDA.n1148 53.3664
R4455 GNDA.n1155 GNDA.n1154 53.3664
R4456 GNDA.n1158 GNDA.n1157 53.3664
R4457 GNDA.n1163 GNDA.n1162 53.3664
R4458 GNDA.n1133 GNDA.n1132 53.3664
R4459 GNDA.n1138 GNDA.n1137 53.3664
R4460 GNDA.n1141 GNDA.n1140 53.3664
R4461 GNDA.n1146 GNDA.n1145 53.3664
R4462 GNDA.n1124 GNDA.n1109 53.3664
R4463 GNDA.n1123 GNDA.n1122 53.3664
R4464 GNDA.n1116 GNDA.n1111 53.3664
R4465 GNDA.n1117 GNDA.n1116 53.3664
R4466 GNDA.n1122 GNDA.n1121 53.3664
R4467 GNDA.n1125 GNDA.n1124 53.3664
R4468 GNDA.n1132 GNDA.n1107 53.3664
R4469 GNDA.n1139 GNDA.n1138 53.3664
R4470 GNDA.n1140 GNDA.n1105 53.3664
R4471 GNDA.n1147 GNDA.n1146 53.3664
R4472 GNDA.n1164 GNDA.n1163 53.3664
R4473 GNDA.n1157 GNDA.n1100 53.3664
R4474 GNDA.n1156 GNDA.n1155 53.3664
R4475 GNDA.n1150 GNDA.n1149 53.3664
R4476 GNDA.n1835 GNDA.n1834 53.3664
R4477 GNDA.n1600 GNDA.n1599 53.3664
R4478 GNDA.n1823 GNDA.n1822 53.3664
R4479 GNDA.n1740 GNDA.n1739 53.3664
R4480 GNDA.n1792 GNDA.n1791 53.3664
R4481 GNDA.n1796 GNDA.n1795 53.3664
R4482 GNDA.n1801 GNDA.n1800 53.3664
R4483 GNDA.n1804 GNDA.n1803 53.3664
R4484 GNDA.n1776 GNDA.n1775 53.3664
R4485 GNDA.n1779 GNDA.n1778 53.3664
R4486 GNDA.n1784 GNDA.n1783 53.3664
R4487 GNDA.n1787 GNDA.n1786 53.3664
R4488 GNDA.n1769 GNDA.n1768 53.3664
R4489 GNDA.n1762 GNDA.n1751 53.3664
R4490 GNDA.n1761 GNDA.n1760 53.3664
R4491 GNDA.n1760 GNDA.n1759 53.3664
R4492 GNDA.n1763 GNDA.n1762 53.3664
R4493 GNDA.n1768 GNDA.n1767 53.3664
R4494 GNDA.n1777 GNDA.n1776 53.3664
R4495 GNDA.n1778 GNDA.n1747 53.3664
R4496 GNDA.n1785 GNDA.n1784 53.3664
R4497 GNDA.n1786 GNDA.n1745 53.3664
R4498 GNDA.n1805 GNDA.n1804 53.3664
R4499 GNDA.n1802 GNDA.n1801 53.3664
R4500 GNDA.n1795 GNDA.n1742 53.3664
R4501 GNDA.n1793 GNDA.n1792 53.3664
R4502 GNDA.n2047 GNDA.n2046 53.3664
R4503 GNDA.n2034 GNDA.n1936 53.3664
R4504 GNDA.n2032 GNDA.n2031 53.3664
R4505 GNDA.n1951 GNDA.n1950 53.3664
R4506 GNDA.n2001 GNDA.n2000 53.3664
R4507 GNDA.n2005 GNDA.n2004 53.3664
R4508 GNDA.n2010 GNDA.n2009 53.3664
R4509 GNDA.n2013 GNDA.n2012 53.3664
R4510 GNDA.n1985 GNDA.n1984 53.3664
R4511 GNDA.n1988 GNDA.n1987 53.3664
R4512 GNDA.n1993 GNDA.n1992 53.3664
R4513 GNDA.n1996 GNDA.n1995 53.3664
R4514 GNDA.n1978 GNDA.n1977 53.3664
R4515 GNDA.n1971 GNDA.n1962 53.3664
R4516 GNDA.n1970 GNDA.n1969 53.3664
R4517 GNDA.n1969 GNDA.n1968 53.3664
R4518 GNDA.n1972 GNDA.n1971 53.3664
R4519 GNDA.n1977 GNDA.n1976 53.3664
R4520 GNDA.n1986 GNDA.n1985 53.3664
R4521 GNDA.n1987 GNDA.n1958 53.3664
R4522 GNDA.n1994 GNDA.n1993 53.3664
R4523 GNDA.n1995 GNDA.n1956 53.3664
R4524 GNDA.n2014 GNDA.n2013 53.3664
R4525 GNDA.n2011 GNDA.n2010 53.3664
R4526 GNDA.n2004 GNDA.n1953 53.3664
R4527 GNDA.n2002 GNDA.n2001 53.3664
R4528 GNDA.n2335 GNDA.n2334 53.3664
R4529 GNDA.n2336 GNDA.n125 53.3664
R4530 GNDA.n2410 GNDA.n2409 53.3664
R4531 GNDA.n2401 GNDA.n2400 53.3664
R4532 GNDA.n2384 GNDA.n2383 53.3664
R4533 GNDA.n2390 GNDA.n2389 53.3664
R4534 GNDA.n2393 GNDA.n2392 53.3664
R4535 GNDA.n2398 GNDA.n2397 53.3664
R4536 GNDA.n2368 GNDA.n2367 53.3664
R4537 GNDA.n2373 GNDA.n2372 53.3664
R4538 GNDA.n2376 GNDA.n2375 53.3664
R4539 GNDA.n2381 GNDA.n2380 53.3664
R4540 GNDA.n2359 GNDA.n135 53.3664
R4541 GNDA.n2358 GNDA.n2357 53.3664
R4542 GNDA.n2351 GNDA.n137 53.3664
R4543 GNDA.n2352 GNDA.n2351 53.3664
R4544 GNDA.n2357 GNDA.n2356 53.3664
R4545 GNDA.n2360 GNDA.n2359 53.3664
R4546 GNDA.n2367 GNDA.n133 53.3664
R4547 GNDA.n2374 GNDA.n2373 53.3664
R4548 GNDA.n2375 GNDA.n131 53.3664
R4549 GNDA.n2382 GNDA.n2381 53.3664
R4550 GNDA.n2399 GNDA.n2398 53.3664
R4551 GNDA.n2392 GNDA.n126 53.3664
R4552 GNDA.n2391 GNDA.n2390 53.3664
R4553 GNDA.n2385 GNDA.n2384 53.3664
R4554 GNDA.n2402 GNDA.n2401 53.3664
R4555 GNDA.n2411 GNDA.n2410 53.3664
R4556 GNDA.n2337 GNDA.n2336 53.3664
R4557 GNDA.n2334 GNDA.n140 53.3664
R4558 GNDA.n1950 GNDA.n1938 53.3664
R4559 GNDA.n2033 GNDA.n2032 53.3664
R4560 GNDA.n1936 GNDA.n1930 53.3664
R4561 GNDA.n2048 GNDA.n2047 53.3664
R4562 GNDA.n1739 GNDA.n1601 53.3664
R4563 GNDA.n1824 GNDA.n1823 53.3664
R4564 GNDA.n1599 GNDA.n607 53.3664
R4565 GNDA.n1836 GNDA.n1835 53.3664
R4566 GNDA.n1093 GNDA.n1086 53.3664
R4567 GNDA.n1175 GNDA.n1174 53.3664
R4568 GNDA.n1084 GNDA.n1077 53.3664
R4569 GNDA.n1186 GNDA.n1185 53.3664
R4570 GNDA.n964 GNDA.n691 53.3664
R4571 GNDA.n962 GNDA.n960 53.3664
R4572 GNDA.n977 GNDA.n976 53.3664
R4573 GNDA.n958 GNDA.n706 53.3664
R4574 GNDA.n765 GNDA.n758 53.3664
R4575 GNDA.n851 GNDA.n850 53.3664
R4576 GNDA.n756 GNDA.n749 53.3664
R4577 GNDA.n862 GNDA.n861 53.3664
R4578 GNDA.n304 GNDA.n297 53.3664
R4579 GNDA.n2265 GNDA.n2264 53.3664
R4580 GNDA.n295 GNDA.n288 53.3664
R4581 GNDA.n2276 GNDA.n2275 53.3664
R4582 GNDA.n1285 GNDA.n1278 53.3664
R4583 GNDA.n1366 GNDA.n1365 53.3664
R4584 GNDA.n1276 GNDA.n1269 53.3664
R4585 GNDA.n1377 GNDA.n1376 53.3664
R4586 GNDA.n1464 GNDA.n1463 53.3664
R4587 GNDA.n1460 GNDA.n1452 53.3664
R4588 GNDA.n1475 GNDA.n1474 53.3664
R4589 GNDA.n1450 GNDA.n1407 53.3664
R4590 GNDA.n2120 GNDA.n2117 52.3879
R4591 GNDA.n2321 GNDA.n173 52.3879
R4592 GNDA.n230 GNDA.n216 52.3879
R4593 GNDA.n477 GNDA.n344 50.5752
R4594 GNDA.t249 GNDA.t328 50.5752
R4595 GNDA.t186 GNDA.t193 50.5752
R4596 GNDA.t183 GNDA.t316 50.5752
R4597 GNDA.t29 GNDA.t323 50.5752
R4598 GNDA.t144 GNDA.t24 50.5752
R4599 GNDA.t2 GNDA.t123 50.5752
R4600 GNDA.t111 GNDA.t13 50.5752
R4601 GNDA.t332 GNDA.t103 50.5752
R4602 GNDA.t317 GNDA.t11 50.5752
R4603 GNDA.t161 GNDA.t5 50.5752
R4604 GNDA.t322 GNDA.t59 50.5752
R4605 GNDA.t335 GNDA.t25 50.5752
R4606 GNDA.t315 GNDA.t288 50.5752
R4607 GNDA.n2460 GNDA.n60 50.5752
R4608 GNDA.n2483 GNDA.n33 49.6005
R4609 GNDA.n2126 GNDA.n520 49.1137
R4610 GNDA.n2127 GNDA.n2126 49.1137
R4611 GNDA.n2129 GNDA.n2127 49.1137
R4612 GNDA.n2129 GNDA.n2128 49.1137
R4613 GNDA.n2136 GNDA.n2135 49.1137
R4614 GNDA.n2137 GNDA.n2136 49.1137
R4615 GNDA.n2137 GNDA.n508 49.1137
R4616 GNDA.n2144 GNDA.n511 49.1137
R4617 GNDA.n493 GNDA.n173 49.1137
R4618 GNDA.n499 GNDA.n493 49.1137
R4619 GNDA.n2155 GNDA.n2153 49.1137
R4620 GNDA.n2155 GNDA.n2154 49.1137
R4621 GNDA.n2179 GNDA.n2178 49.1137
R4622 GNDA.n2183 GNDA.n2182 49.1137
R4623 GNDA.n230 GNDA.n229 49.1137
R4624 GNDA.n229 GNDA.n228 49.1137
R4625 GNDA.n228 GNDA.n219 49.1137
R4626 GNDA.n222 GNDA.n219 49.1137
R4627 GNDA.n222 GNDA.n117 49.1137
R4628 GNDA.n2416 GNDA.n104 49.1137
R4629 GNDA.n2423 GNDA.n108 49.1137
R4630 GNDA.n111 GNDA.n108 49.1137
R4631 GNDA.n111 GNDA.n93 49.1137
R4632 GNDA.n50 GNDA.t44 48.0005
R4633 GNDA.n50 GNDA.t36 48.0005
R4634 GNDA.n46 GNDA.t78 48.0005
R4635 GNDA.n46 GNDA.t38 48.0005
R4636 GNDA.n47 GNDA.t66 48.0005
R4637 GNDA.n47 GNDA.t42 48.0005
R4638 GNDA.n44 GNDA.t64 48.0005
R4639 GNDA.n44 GNDA.t164 48.0005
R4640 GNDA.n43 GNDA.t68 48.0005
R4641 GNDA.n43 GNDA.t40 48.0005
R4642 GNDA.t230 GNDA.n2321 47.4766
R4643 GNDA.n2164 GNDA.n2163 47.4766
R4644 GNDA.t230 GNDA.n172 46.9309
R4645 GNDA.t230 GNDA.n169 46.9309
R4646 GNDA.t130 GNDA.t347 46.3607
R4647 GNDA.t130 GNDA.t147 46.3607
R4648 GNDA.t100 GNDA.n2474 46.3607
R4649 GNDA.t31 GNDA.t118 46.3607
R4650 GNDA.t86 GNDA.t31 46.3607
R4651 GNDA.n1816 GNDA.n1733 43.0993
R4652 GNDA.n120 GNDA.n118 43.0993
R4653 GNDA.t185 GNDA.t169 43.0173
R4654 GNDA.t107 GNDA.t82 43.0173
R4655 GNDA.t154 GNDA.t249 42.1461
R4656 GNDA.t193 GNDA.t183 42.1461
R4657 GNDA.t316 GNDA.t29 42.1461
R4658 GNDA.t323 GNDA.t144 42.1461
R4659 GNDA.t24 GNDA.t2 42.1461
R4660 GNDA.t123 GNDA.t46 42.1461
R4661 GNDA.t218 GNDA.t340 42.1461
R4662 GNDA.t92 GNDA.t298 42.1461
R4663 GNDA.t7 GNDA.t111 42.1461
R4664 GNDA.t13 GNDA.t332 42.1461
R4665 GNDA.t103 GNDA.t317 42.1461
R4666 GNDA.t11 GNDA.t161 42.1461
R4667 GNDA.t5 GNDA.t322 42.1461
R4668 GNDA.t59 GNDA.t335 42.1461
R4669 GNDA.t25 GNDA.t315 42.1461
R4670 GNDA.t288 GNDA.t160 42.1461
R4671 GNDA.n2152 GNDA.n499 42.0196
R4672 GNDA.n78 GNDA.t143 39.7033
R4673 GNDA.t165 GNDA.n360 39.7033
R4674 GNDA.t147 GNDA.n458 37.9315
R4675 GNDA.n2481 GNDA.t328 37.9315
R4676 GNDA.t46 GNDA.n2477 37.9315
R4677 GNDA.t10 GNDA.t73 37.9315
R4678 GNDA.t118 GNDA.n427 37.9315
R4679 GNDA.n2454 GNDA.n65 37.3678
R4680 GNDA.n362 GNDA.n355 37.3678
R4681 GNDA.n2179 GNDA.n308 36.5626
R4682 GNDA.n2454 GNDA.t180 35.0323
R4683 GNDA.t138 GNDA.n362 35.0323
R4684 GNDA.n2117 GNDA.n485 33.8341
R4685 GNDA.n383 GNDA.n382 32.0005
R4686 GNDA.n388 GNDA.n386 32.0005
R4687 GNDA.n2120 GNDA.n2119 31.1055
R4688 GNDA.n2177 GNDA.n312 31.1055
R4689 GNDA.n216 GNDA.n168 31.1055
R4690 GNDA.t234 GNDA.n611 31.0997
R4691 GNDA.n526 GNDA.t230 31.0997
R4692 GNDA.t207 GNDA.t128 30.7268
R4693 GNDA.t48 GNDA.t313 30.7268
R4694 GNDA.t125 GNDA.t171 30.7268
R4695 GNDA.t167 GNDA.t166 30.7268
R4696 GNDA.n67 GNDA.t72 30.3614
R4697 GNDA.t180 GNDA.n2453 30.3614
R4698 GNDA.n76 GNDA.t124 30.3614
R4699 GNDA.t152 GNDA.n361 30.3614
R4700 GNDA.n363 GNDA.t138 30.3614
R4701 GNDA.n369 GNDA.t150 30.3614
R4702 GNDA.t0 GNDA.t134 29.5024
R4703 GNDA.t330 GNDA.t52 29.5024
R4704 GNDA.n2489 GNDA.t7 29.5024
R4705 GNDA.t33 GNDA.t50 29.5024
R4706 GNDA.t326 GNDA.t157 29.5024
R4707 GNDA.n463 GNDA.n462 28.5224
R4708 GNDA.n440 GNDA.n439 28.1864
R4709 GNDA.n480 GNDA.n479 28.1786
R4710 GNDA.n2166 GNDA.n99 28.1318
R4711 GNDA.n474 GNDA.n373 27.8818
R4712 GNDA.n447 GNDA.n63 27.8818
R4713 GNDA.n1721 GNDA.n1617 27.8193
R4714 GNDA.n1719 GNDA.n1718 27.8193
R4715 GNDA.n1504 GNDA.n1503 27.5561
R4716 GNDA.n1319 GNDA.n1299 27.5561
R4717 GNDA.n2218 GNDA.n2198 27.5561
R4718 GNDA.n804 GNDA.n784 27.5561
R4719 GNDA.n1004 GNDA.n700 27.5561
R4720 GNDA.n1128 GNDA.n1108 27.5561
R4721 GNDA.n1773 GNDA.n1772 27.5561
R4722 GNDA.n1982 GNDA.n1981 27.5561
R4723 GNDA.n2363 GNDA.n134 27.5561
R4724 GNDA.n577 GNDA.n558 26.9584
R4725 GNDA.n2291 GNDA.n187 26.9584
R4726 GNDA.t149 GNDA.n67 25.6905
R4727 GNDA.t143 GNDA.n76 25.6905
R4728 GNDA.n361 GNDA.t165 25.6905
R4729 GNDA.n369 GNDA.t179 25.6905
R4730 GNDA.n2128 GNDA.t230 25.6485
R4731 GNDA.n2154 GNDA.t230 25.6485
R4732 GNDA.t230 GNDA.n117 25.6485
R4733 GNDA.n376 GNDA.n375 25.6005
R4734 GNDA.n439 GNDA.n438 25.6005
R4735 GNDA.n433 GNDA.n432 25.6005
R4736 GNDA.t124 GNDA.t102 25.2234
R4737 GNDA.t153 GNDA.t152 25.2234
R4738 GNDA.n1702 GNDA.n1700 24.5815
R4739 GNDA.n1691 GNDA.n1636 24.5815
R4740 GNDA.n1666 GNDA.t113 24.0005
R4741 GNDA.n1666 GNDA.t28 24.0005
R4742 GNDA.n1664 GNDA.t83 24.0005
R4743 GNDA.n1664 GNDA.t195 24.0005
R4744 GNDA.n1662 GNDA.t172 24.0005
R4745 GNDA.n1662 GNDA.t168 24.0005
R4746 GNDA.n1660 GNDA.t117 24.0005
R4747 GNDA.n1660 GNDA.t197 24.0005
R4748 GNDA.n1658 GNDA.t174 24.0005
R4749 GNDA.n1658 GNDA.t85 24.0005
R4750 GNDA.n1656 GNDA.t142 24.0005
R4751 GNDA.n1656 GNDA.t176 24.0005
R4752 GNDA.n1654 GNDA.t325 24.0005
R4753 GNDA.n1654 GNDA.t133 24.0005
R4754 GNDA.n1652 GNDA.t129 24.0005
R4755 GNDA.n1652 GNDA.t49 24.0005
R4756 GNDA.n1650 GNDA.t346 24.0005
R4757 GNDA.n1650 GNDA.t170 24.0005
R4758 GNDA.n1649 GNDA.t115 24.0005
R4759 GNDA.n1649 GNDA.t137 24.0005
R4760 GNDA.n1521 GNDA.n1520 23.6449
R4761 GNDA.n1295 GNDA.n1294 23.6449
R4762 GNDA.n2194 GNDA.n2193 23.6449
R4763 GNDA.n780 GNDA.n779 23.6449
R4764 GNDA.n696 GNDA.n695 23.6449
R4765 GNDA.n1104 GNDA.n1103 23.6449
R4766 GNDA.n1790 GNDA.n1789 23.6449
R4767 GNDA.n1999 GNDA.n1998 23.6449
R4768 GNDA.n130 GNDA.n129 23.6449
R4769 GNDA.n2135 GNDA.t230 23.4657
R4770 GNDA.n2163 GNDA.t230 23.4657
R4771 GNDA.n2416 GNDA.t230 23.4657
R4772 GNDA.n2494 GNDA.n12 22.688
R4773 GNDA.n24 GNDA.n23 22.5943
R4774 GNDA.n373 GNDA.n372 22.4005
R4775 GNDA.n2458 GNDA.n63 22.4005
R4776 GNDA.t101 GNDA.t21 21.8286
R4777 GNDA.n549 GNDA.n488 21.4917
R4778 GNDA.n2074 GNDA.t236 21.4482
R4779 GNDA.n55 GNDA.n54 21.3338
R4780 GNDA.n58 GNDA.n57 21.3338
R4781 GNDA.n332 GNDA.n331 21.3338
R4782 GNDA.n334 GNDA.n333 21.3338
R4783 GNDA.n2471 GNDA.n2470 21.3338
R4784 GNDA.n41 GNDA.n40 21.3338
R4785 GNDA.n384 GNDA.n379 21.3338
R4786 GNDA.n383 GNDA.n380 21.3338
R4787 GNDA.n382 GNDA.n381 21.3338
R4788 GNDA.n386 GNDA.n385 21.3338
R4789 GNDA.n388 GNDA.n387 21.3338
R4790 GNDA.n390 GNDA.n389 21.3338
R4791 GNDA.n461 GNDA.n456 21.3338
R4792 GNDA.n324 GNDA.n323 21.3338
R4793 GNDA.n377 GNDA.n374 21.3338
R4794 GNDA.n348 GNDA.n347 21.3338
R4795 GNDA.n442 GNDA.n441 21.3338
R4796 GNDA.n431 GNDA.n430 21.3338
R4797 GNDA.n426 GNDA.n425 21.3338
R4798 GNDA.n394 GNDA.n393 21.3338
R4799 GNDA.n1647 GNDA.n1644 21.3338
R4800 GNDA.n1646 GNDA.n1645 21.3338
R4801 GNDA.n1722 GNDA.n1616 21.3338
R4802 GNDA.n1615 GNDA.n1614 21.3338
R4803 GNDA.n1619 GNDA.n1618 21.3338
R4804 GNDA.n1704 GNDA.n1703 21.3338
R4805 GNDA.n1672 GNDA.n1669 21.1792
R4806 GNDA.n378 GNDA.t318 21.0733
R4807 GNDA.n2489 GNDA.t298 21.0733
R4808 GNDA.n2496 GNDA.n0 20.0005
R4809 GNDA.n22 GNDA.t201 19.7005
R4810 GNDA.n22 GNDA.t211 19.7005
R4811 GNDA.n20 GNDA.t9 19.7005
R4812 GNDA.n20 GNDA.t189 19.7005
R4813 GNDA.n18 GNDA.t122 19.7005
R4814 GNDA.n18 GNDA.t191 19.7005
R4815 GNDA.n16 GNDA.t162 19.7005
R4816 GNDA.n16 GNDA.t202 19.7005
R4817 GNDA.n14 GNDA.t198 19.7005
R4818 GNDA.n14 GNDA.t188 19.7005
R4819 GNDA.n13 GNDA.t209 19.7005
R4820 GNDA.n13 GNDA.t190 19.7005
R4821 GNDA.n2 GNDA.t19 19.7005
R4822 GNDA.n2 GNDA.t215 19.7005
R4823 GNDA.n3 GNDA.t320 19.7005
R4824 GNDA.n3 GNDA.t75 19.7005
R4825 GNDA.n5 GNDA.t329 19.7005
R4826 GNDA.n5 GNDA.t319 19.7005
R4827 GNDA.n7 GNDA.t76 19.7005
R4828 GNDA.n7 GNDA.t177 19.7005
R4829 GNDA.n9 GNDA.t178 19.7005
R4830 GNDA.n9 GNDA.t336 19.7005
R4831 GNDA.n11 GNDA.t210 19.7005
R4832 GNDA.n11 GNDA.t96 19.7005
R4833 GNDA.n546 GNDA.n545 19.4279
R4834 GNDA.n1695 GNDA.n1693 19.2005
R4835 GNDA.n2149 GNDA.n2148 19.2005
R4836 GNDA.n2427 GNDA.n2426 19.2005
R4837 GNDA.n509 GNDA.n488 19.2005
R4838 GNDA.n2167 GNDA.n316 19.2005
R4839 GNDA.n1628 GNDA.n1607 19.2005
R4840 GNDA.n2450 GNDA.n2449 19.1943
R4841 GNDA.n358 GNDA.n320 19.1474
R4842 GNDA.n375 GNDA.n325 18.913
R4843 GNDA.n434 GNDA.n433 18.913
R4844 GNDA.n68 GNDA.n65 18.6842
R4845 GNDA.n368 GNDA.n355 18.6842
R4846 GNDA.t203 GNDA.t48 18.4363
R4847 GNDA.t171 GNDA.t4 18.4363
R4848 GNDA.n2119 GNDA.n520 18.0087
R4849 GNDA.n2178 GNDA.n2177 18.0087
R4850 GNDA.n1697 GNDA.n1628 17.613
R4851 GNDA.n2072 GNDA.n550 17.4917
R4852 GNDA.n2070 GNDA.n2069 16.9605
R4853 GNDA.n1870 GNDA.n585 16.9379
R4854 GNDA.n1590 GNDA.n622 16.9379
R4855 GNDA.n893 GNDA.n892 16.9379
R4856 GNDA.t230 GNDA.n168 16.3716
R4857 GNDA.n68 GNDA.t149 16.3487
R4858 GNDA.t333 GNDA.n78 16.3487
R4859 GNDA.n360 GNDA.t344 16.3487
R4860 GNDA.t179 GNDA.n368 16.3487
R4861 GNDA.n1503 GNDA.n1402 16.0005
R4862 GNDA.n1497 GNDA.n1402 16.0005
R4863 GNDA.n1497 GNDA.n1496 16.0005
R4864 GNDA.n1496 GNDA.n1495 16.0005
R4865 GNDA.n1495 GNDA.n1404 16.0005
R4866 GNDA.n1489 GNDA.n1404 16.0005
R4867 GNDA.n1489 GNDA.n1488 16.0005
R4868 GNDA.n1488 GNDA.n1487 16.0005
R4869 GNDA.n1505 GNDA.n1504 16.0005
R4870 GNDA.n1505 GNDA.n1400 16.0005
R4871 GNDA.n1511 GNDA.n1400 16.0005
R4872 GNDA.n1512 GNDA.n1511 16.0005
R4873 GNDA.n1513 GNDA.n1512 16.0005
R4874 GNDA.n1513 GNDA.n1398 16.0005
R4875 GNDA.n1519 GNDA.n1398 16.0005
R4876 GNDA.n1520 GNDA.n1519 16.0005
R4877 GNDA.n1521 GNDA.n1396 16.0005
R4878 GNDA.n1396 GNDA.n1395 16.0005
R4879 GNDA.n1528 GNDA.n1395 16.0005
R4880 GNDA.n1529 GNDA.n1528 16.0005
R4881 GNDA.n1530 GNDA.n1393 16.0005
R4882 GNDA.n1393 GNDA.n1391 16.0005
R4883 GNDA.n1537 GNDA.n1391 16.0005
R4884 GNDA.n1319 GNDA.n1318 16.0005
R4885 GNDA.n1318 GNDA.n1317 16.0005
R4886 GNDA.n1317 GNDA.n1301 16.0005
R4887 GNDA.n1311 GNDA.n1301 16.0005
R4888 GNDA.n1311 GNDA.n1310 16.0005
R4889 GNDA.n1310 GNDA.n1309 16.0005
R4890 GNDA.n1309 GNDA.n1303 16.0005
R4891 GNDA.n1304 GNDA.n1303 16.0005
R4892 GNDA.n1325 GNDA.n1299 16.0005
R4893 GNDA.n1326 GNDA.n1325 16.0005
R4894 GNDA.n1327 GNDA.n1326 16.0005
R4895 GNDA.n1327 GNDA.n1297 16.0005
R4896 GNDA.n1333 GNDA.n1297 16.0005
R4897 GNDA.n1334 GNDA.n1333 16.0005
R4898 GNDA.n1335 GNDA.n1334 16.0005
R4899 GNDA.n1335 GNDA.n1295 16.0005
R4900 GNDA.n1342 GNDA.n1294 16.0005
R4901 GNDA.n1343 GNDA.n1342 16.0005
R4902 GNDA.n1344 GNDA.n1343 16.0005
R4903 GNDA.n1344 GNDA.n1292 16.0005
R4904 GNDA.n1351 GNDA.n1350 16.0005
R4905 GNDA.n1352 GNDA.n1351 16.0005
R4906 GNDA.n1352 GNDA.n1290 16.0005
R4907 GNDA.n2218 GNDA.n2217 16.0005
R4908 GNDA.n2217 GNDA.n2216 16.0005
R4909 GNDA.n2216 GNDA.n2200 16.0005
R4910 GNDA.n2210 GNDA.n2200 16.0005
R4911 GNDA.n2210 GNDA.n2209 16.0005
R4912 GNDA.n2209 GNDA.n2208 16.0005
R4913 GNDA.n2208 GNDA.n2202 16.0005
R4914 GNDA.n2203 GNDA.n2202 16.0005
R4915 GNDA.n2224 GNDA.n2198 16.0005
R4916 GNDA.n2225 GNDA.n2224 16.0005
R4917 GNDA.n2226 GNDA.n2225 16.0005
R4918 GNDA.n2226 GNDA.n2196 16.0005
R4919 GNDA.n2232 GNDA.n2196 16.0005
R4920 GNDA.n2233 GNDA.n2232 16.0005
R4921 GNDA.n2234 GNDA.n2233 16.0005
R4922 GNDA.n2234 GNDA.n2194 16.0005
R4923 GNDA.n2241 GNDA.n2193 16.0005
R4924 GNDA.n2242 GNDA.n2241 16.0005
R4925 GNDA.n2243 GNDA.n2242 16.0005
R4926 GNDA.n2243 GNDA.n2191 16.0005
R4927 GNDA.n2250 GNDA.n2249 16.0005
R4928 GNDA.n2251 GNDA.n2250 16.0005
R4929 GNDA.n2251 GNDA.n2189 16.0005
R4930 GNDA.n804 GNDA.n803 16.0005
R4931 GNDA.n803 GNDA.n802 16.0005
R4932 GNDA.n802 GNDA.n786 16.0005
R4933 GNDA.n796 GNDA.n786 16.0005
R4934 GNDA.n796 GNDA.n795 16.0005
R4935 GNDA.n795 GNDA.n794 16.0005
R4936 GNDA.n794 GNDA.n788 16.0005
R4937 GNDA.n789 GNDA.n788 16.0005
R4938 GNDA.n810 GNDA.n784 16.0005
R4939 GNDA.n811 GNDA.n810 16.0005
R4940 GNDA.n812 GNDA.n811 16.0005
R4941 GNDA.n812 GNDA.n782 16.0005
R4942 GNDA.n818 GNDA.n782 16.0005
R4943 GNDA.n819 GNDA.n818 16.0005
R4944 GNDA.n820 GNDA.n819 16.0005
R4945 GNDA.n820 GNDA.n780 16.0005
R4946 GNDA.n827 GNDA.n779 16.0005
R4947 GNDA.n828 GNDA.n827 16.0005
R4948 GNDA.n829 GNDA.n828 16.0005
R4949 GNDA.n829 GNDA.n777 16.0005
R4950 GNDA.n836 GNDA.n835 16.0005
R4951 GNDA.n837 GNDA.n836 16.0005
R4952 GNDA.n837 GNDA.n775 16.0005
R4953 GNDA.n1004 GNDA.n1003 16.0005
R4954 GNDA.n1003 GNDA.n1002 16.0005
R4955 GNDA.n1002 GNDA.n702 16.0005
R4956 GNDA.n996 GNDA.n702 16.0005
R4957 GNDA.n996 GNDA.n995 16.0005
R4958 GNDA.n995 GNDA.n994 16.0005
R4959 GNDA.n994 GNDA.n704 16.0005
R4960 GNDA.n705 GNDA.n704 16.0005
R4961 GNDA.n1010 GNDA.n700 16.0005
R4962 GNDA.n1011 GNDA.n1010 16.0005
R4963 GNDA.n1012 GNDA.n1011 16.0005
R4964 GNDA.n1012 GNDA.n698 16.0005
R4965 GNDA.n1018 GNDA.n698 16.0005
R4966 GNDA.n1019 GNDA.n1018 16.0005
R4967 GNDA.n1020 GNDA.n1019 16.0005
R4968 GNDA.n1020 GNDA.n696 16.0005
R4969 GNDA.n1027 GNDA.n695 16.0005
R4970 GNDA.n1028 GNDA.n1027 16.0005
R4971 GNDA.n1029 GNDA.n1028 16.0005
R4972 GNDA.n1029 GNDA.n693 16.0005
R4973 GNDA.n1036 GNDA.n1035 16.0005
R4974 GNDA.n1037 GNDA.n1036 16.0005
R4975 GNDA.n1037 GNDA.n688 16.0005
R4976 GNDA.n1128 GNDA.n1127 16.0005
R4977 GNDA.n1127 GNDA.n1126 16.0005
R4978 GNDA.n1126 GNDA.n1110 16.0005
R4979 GNDA.n1120 GNDA.n1110 16.0005
R4980 GNDA.n1120 GNDA.n1119 16.0005
R4981 GNDA.n1119 GNDA.n1118 16.0005
R4982 GNDA.n1118 GNDA.n1112 16.0005
R4983 GNDA.n1113 GNDA.n1112 16.0005
R4984 GNDA.n1134 GNDA.n1108 16.0005
R4985 GNDA.n1135 GNDA.n1134 16.0005
R4986 GNDA.n1136 GNDA.n1135 16.0005
R4987 GNDA.n1136 GNDA.n1106 16.0005
R4988 GNDA.n1142 GNDA.n1106 16.0005
R4989 GNDA.n1143 GNDA.n1142 16.0005
R4990 GNDA.n1144 GNDA.n1143 16.0005
R4991 GNDA.n1144 GNDA.n1104 16.0005
R4992 GNDA.n1151 GNDA.n1103 16.0005
R4993 GNDA.n1152 GNDA.n1151 16.0005
R4994 GNDA.n1153 GNDA.n1152 16.0005
R4995 GNDA.n1153 GNDA.n1101 16.0005
R4996 GNDA.n1160 GNDA.n1159 16.0005
R4997 GNDA.n1161 GNDA.n1160 16.0005
R4998 GNDA.n1161 GNDA.n1099 16.0005
R4999 GNDA.n1772 GNDA.n1750 16.0005
R5000 GNDA.n1766 GNDA.n1750 16.0005
R5001 GNDA.n1766 GNDA.n1765 16.0005
R5002 GNDA.n1765 GNDA.n1764 16.0005
R5003 GNDA.n1764 GNDA.n1752 16.0005
R5004 GNDA.n1758 GNDA.n1752 16.0005
R5005 GNDA.n1758 GNDA.n1757 16.0005
R5006 GNDA.n1757 GNDA.n1756 16.0005
R5007 GNDA.n1774 GNDA.n1773 16.0005
R5008 GNDA.n1774 GNDA.n1748 16.0005
R5009 GNDA.n1780 GNDA.n1748 16.0005
R5010 GNDA.n1781 GNDA.n1780 16.0005
R5011 GNDA.n1782 GNDA.n1781 16.0005
R5012 GNDA.n1782 GNDA.n1746 16.0005
R5013 GNDA.n1788 GNDA.n1746 16.0005
R5014 GNDA.n1789 GNDA.n1788 16.0005
R5015 GNDA.n1790 GNDA.n1744 16.0005
R5016 GNDA.n1744 GNDA.n1743 16.0005
R5017 GNDA.n1797 GNDA.n1743 16.0005
R5018 GNDA.n1798 GNDA.n1797 16.0005
R5019 GNDA.n1799 GNDA.n1741 16.0005
R5020 GNDA.n1741 GNDA.n1738 16.0005
R5021 GNDA.n1806 GNDA.n1738 16.0005
R5022 GNDA.n1981 GNDA.n1961 16.0005
R5023 GNDA.n1975 GNDA.n1961 16.0005
R5024 GNDA.n1975 GNDA.n1974 16.0005
R5025 GNDA.n1974 GNDA.n1973 16.0005
R5026 GNDA.n1973 GNDA.n1963 16.0005
R5027 GNDA.n1967 GNDA.n1963 16.0005
R5028 GNDA.n1967 GNDA.n1966 16.0005
R5029 GNDA.n1966 GNDA.n1926 16.0005
R5030 GNDA.n1983 GNDA.n1982 16.0005
R5031 GNDA.n1983 GNDA.n1959 16.0005
R5032 GNDA.n1989 GNDA.n1959 16.0005
R5033 GNDA.n1990 GNDA.n1989 16.0005
R5034 GNDA.n1991 GNDA.n1990 16.0005
R5035 GNDA.n1991 GNDA.n1957 16.0005
R5036 GNDA.n1997 GNDA.n1957 16.0005
R5037 GNDA.n1998 GNDA.n1997 16.0005
R5038 GNDA.n1999 GNDA.n1955 16.0005
R5039 GNDA.n1955 GNDA.n1954 16.0005
R5040 GNDA.n2006 GNDA.n1954 16.0005
R5041 GNDA.n2007 GNDA.n2006 16.0005
R5042 GNDA.n2008 GNDA.n1952 16.0005
R5043 GNDA.n1952 GNDA.n1949 16.0005
R5044 GNDA.n2015 GNDA.n1949 16.0005
R5045 GNDA.n2363 GNDA.n2362 16.0005
R5046 GNDA.n2362 GNDA.n2361 16.0005
R5047 GNDA.n2361 GNDA.n136 16.0005
R5048 GNDA.n2355 GNDA.n136 16.0005
R5049 GNDA.n2355 GNDA.n2354 16.0005
R5050 GNDA.n2354 GNDA.n2353 16.0005
R5051 GNDA.n2353 GNDA.n138 16.0005
R5052 GNDA.n139 GNDA.n138 16.0005
R5053 GNDA.n2369 GNDA.n134 16.0005
R5054 GNDA.n2370 GNDA.n2369 16.0005
R5055 GNDA.n2371 GNDA.n2370 16.0005
R5056 GNDA.n2371 GNDA.n132 16.0005
R5057 GNDA.n2377 GNDA.n132 16.0005
R5058 GNDA.n2378 GNDA.n2377 16.0005
R5059 GNDA.n2379 GNDA.n2378 16.0005
R5060 GNDA.n2379 GNDA.n130 16.0005
R5061 GNDA.n2386 GNDA.n129 16.0005
R5062 GNDA.n2387 GNDA.n2386 16.0005
R5063 GNDA.n2388 GNDA.n2387 16.0005
R5064 GNDA.n2388 GNDA.n127 16.0005
R5065 GNDA.n2395 GNDA.n2394 16.0005
R5066 GNDA.n2396 GNDA.n2395 16.0005
R5067 GNDA.n2396 GNDA.n90 16.0005
R5068 GNDA.n2072 GNDA.n2071 16.0005
R5069 GNDA.n2071 GNDA.n2070 16.0005
R5070 GNDA.n321 GNDA.n320 16.0005
R5071 GNDA.n2449 GNDA.n72 16.0005
R5072 GNDA.n328 GNDA.t110 15.8278
R5073 GNDA.n329 GNDA.t163 15.8278
R5074 GNDA.n338 GNDA.t65 15.8278
R5075 GNDA.t127 GNDA.n339 15.8278
R5076 GNDA.n340 GNDA.t109 15.8278
R5077 GNDA.n1699 GNDA.n1625 15.363
R5078 GNDA.n1712 GNDA.n1699 15.363
R5079 GNDA.t90 GNDA.n2144 14.7345
R5080 GNDA.t21 GNDA.n2423 14.7345
R5081 GNDA.n2493 GNDA.n2492 14.238
R5082 GNDA.n2496 GNDA.n2495 14.133
R5083 GNDA.n2465 GNDA.n2464 14.0661
R5084 GNDA.n2465 GNDA.n53 14.0661
R5085 GNDA.n1530 GNDA 14.0449
R5086 GNDA.n1350 GNDA 14.0449
R5087 GNDA.n2249 GNDA 14.0449
R5088 GNDA.n835 GNDA 14.0449
R5089 GNDA.n1035 GNDA 14.0449
R5090 GNDA.n1159 GNDA 14.0449
R5091 GNDA.n1799 GNDA 14.0449
R5092 GNDA.n2008 GNDA 14.0449
R5093 GNDA.n2394 GNDA 14.0449
R5094 GNDA.n473 GNDA.n472 13.988
R5095 GNDA.n448 GNDA.n424 13.988
R5096 GNDA.n396 GNDA.n395 13.8005
R5097 GNDA.n419 GNDA.n32 13.8005
R5098 GNDA.n1696 GNDA.n1695 13.8005
R5099 GNDA.n1669 GNDA.n550 13.7706
R5100 GNDA.n2287 GNDA.n257 12.9309
R5101 GNDA.n1386 GNDA.n645 12.9309
R5102 GNDA.n710 GNDA.n623 12.9309
R5103 GNDA.n1197 GNDA.n182 12.9309
R5104 GNDA.n476 GNDA.t256 12.6442
R5105 GNDA.t146 GNDA.t224 12.6442
R5106 GNDA.t151 GNDA.t69 12.6442
R5107 GNDA.n2477 GNDA.t218 12.6442
R5108 GNDA.t181 GNDA.n2488 12.6442
R5109 GNDA.t121 GNDA.t155 12.6442
R5110 GNDA.t242 GNDA.t158 12.6442
R5111 GNDA.n445 GNDA.t259 12.6442
R5112 GNDA.n2182 GNDA.n308 12.5517
R5113 GNDA.n218 GNDA.n215 12.4126
R5114 GNDA.n2122 GNDA.n522 12.4126
R5115 GNDA.n495 GNDA.n174 12.4126
R5116 GNDA.n1260 GNDA.n1210 11.6369
R5117 GNDA.n1260 GNDA.n1259 11.6369
R5118 GNDA.n1259 GNDA.n1258 11.6369
R5119 GNDA.n1258 GNDA.n1255 11.6369
R5120 GNDA.n1255 GNDA.n1254 11.6369
R5121 GNDA.n1254 GNDA.n1251 11.6369
R5122 GNDA.n1251 GNDA.n1250 11.6369
R5123 GNDA.n1250 GNDA.n1247 11.6369
R5124 GNDA.n1247 GNDA.n1246 11.6369
R5125 GNDA.n1246 GNDA.n1243 11.6369
R5126 GNDA.n1243 GNDA.n1242 11.6369
R5127 GNDA.n256 GNDA.n209 11.6369
R5128 GNDA.n251 GNDA.n209 11.6369
R5129 GNDA.n251 GNDA.n250 11.6369
R5130 GNDA.n250 GNDA.n211 11.6369
R5131 GNDA.n245 GNDA.n211 11.6369
R5132 GNDA.n245 GNDA.n244 11.6369
R5133 GNDA.n244 GNDA.n243 11.6369
R5134 GNDA.n243 GNDA.n213 11.6369
R5135 GNDA.n237 GNDA.n213 11.6369
R5136 GNDA.n237 GNDA.n236 11.6369
R5137 GNDA.n236 GNDA.n235 11.6369
R5138 GNDA.n221 GNDA.n218 11.6369
R5139 GNDA.n226 GNDA.n221 11.6369
R5140 GNDA.n226 GNDA.n225 11.6369
R5141 GNDA.n225 GNDA.n224 11.6369
R5142 GNDA.n224 GNDA.n114 11.6369
R5143 GNDA.n2418 GNDA.n114 11.6369
R5144 GNDA.n2421 GNDA.n2419 11.6369
R5145 GNDA.n2421 GNDA.n2420 11.6369
R5146 GNDA.n1871 GNDA.n1870 11.6369
R5147 GNDA.n1872 GNDA.n1871 11.6369
R5148 GNDA.n1872 GNDA.n583 11.6369
R5149 GNDA.n1878 GNDA.n583 11.6369
R5150 GNDA.n1879 GNDA.n1878 11.6369
R5151 GNDA.n1880 GNDA.n1879 11.6369
R5152 GNDA.n1880 GNDA.n581 11.6369
R5153 GNDA.n1886 GNDA.n581 11.6369
R5154 GNDA.n1887 GNDA.n1886 11.6369
R5155 GNDA.n1888 GNDA.n1887 11.6369
R5156 GNDA.n1888 GNDA.n578 11.6369
R5157 GNDA.n590 GNDA.n585 11.6369
R5158 GNDA.n1862 GNDA.n590 11.6369
R5159 GNDA.n1862 GNDA.n1861 11.6369
R5160 GNDA.n1861 GNDA.n1860 11.6369
R5161 GNDA.n1860 GNDA.n591 11.6369
R5162 GNDA.n1854 GNDA.n591 11.6369
R5163 GNDA.n1854 GNDA.n1853 11.6369
R5164 GNDA.n1853 GNDA.n1852 11.6369
R5165 GNDA.n1852 GNDA.n595 11.6369
R5166 GNDA.n677 GNDA.n676 11.6369
R5167 GNDA.n676 GNDA.n675 11.6369
R5168 GNDA.n675 GNDA.n673 11.6369
R5169 GNDA.n673 GNDA.n670 11.6369
R5170 GNDA.n670 GNDA.n669 11.6369
R5171 GNDA.n669 GNDA.n666 11.6369
R5172 GNDA.n666 GNDA.n665 11.6369
R5173 GNDA.n665 GNDA.n662 11.6369
R5174 GNDA.n662 GNDA.n661 11.6369
R5175 GNDA.n661 GNDA.n658 11.6369
R5176 GNDA.n658 GNDA.n657 11.6369
R5177 GNDA.n1590 GNDA.n1589 11.6369
R5178 GNDA.n1589 GNDA.n1588 11.6369
R5179 GNDA.n1588 GNDA.n1586 11.6369
R5180 GNDA.n1586 GNDA.n1583 11.6369
R5181 GNDA.n1583 GNDA.n1582 11.6369
R5182 GNDA.n1582 GNDA.n1579 11.6369
R5183 GNDA.n1579 GNDA.n1578 11.6369
R5184 GNDA.n1578 GNDA.n1575 11.6369
R5185 GNDA.n1575 GNDA.n1574 11.6369
R5186 GNDA.n1574 GNDA.n1571 11.6369
R5187 GNDA.n1571 GNDA.n1570 11.6369
R5188 GNDA.n1419 GNDA.n622 11.6369
R5189 GNDA.n1425 GNDA.n1419 11.6369
R5190 GNDA.n1426 GNDA.n1425 11.6369
R5191 GNDA.n1427 GNDA.n1426 11.6369
R5192 GNDA.n1427 GNDA.n1415 11.6369
R5193 GNDA.n1433 GNDA.n1415 11.6369
R5194 GNDA.n1434 GNDA.n1433 11.6369
R5195 GNDA.n1435 GNDA.n1434 11.6369
R5196 GNDA.n1435 GNDA.n1411 11.6369
R5197 GNDA.n892 GNDA.n731 11.6369
R5198 GNDA.n886 GNDA.n731 11.6369
R5199 GNDA.n886 GNDA.n885 11.6369
R5200 GNDA.n885 GNDA.n884 11.6369
R5201 GNDA.n884 GNDA.n735 11.6369
R5202 GNDA.n878 GNDA.n735 11.6369
R5203 GNDA.n878 GNDA.n877 11.6369
R5204 GNDA.n877 GNDA.n876 11.6369
R5205 GNDA.n876 GNDA.n739 11.6369
R5206 GNDA.n894 GNDA.n893 11.6369
R5207 GNDA.n894 GNDA.n727 11.6369
R5208 GNDA.n901 GNDA.n727 11.6369
R5209 GNDA.n902 GNDA.n901 11.6369
R5210 GNDA.n903 GNDA.n902 11.6369
R5211 GNDA.n903 GNDA.n725 11.6369
R5212 GNDA.n908 GNDA.n725 11.6369
R5213 GNDA.n909 GNDA.n908 11.6369
R5214 GNDA.n911 GNDA.n909 11.6369
R5215 GNDA.n911 GNDA.n910 11.6369
R5216 GNDA.n910 GNDA.n722 11.6369
R5217 GNDA.n2060 GNDA.n555 11.6369
R5218 GNDA.n2061 GNDA.n2060 11.6369
R5219 GNDA.n2062 GNDA.n2061 11.6369
R5220 GNDA.n2062 GNDA.n551 11.6369
R5221 GNDA.n2068 GNDA.n551 11.6369
R5222 GNDA.n2078 GNDA.n541 11.6369
R5223 GNDA.n2079 GNDA.n2078 11.6369
R5224 GNDA.n2081 GNDA.n2079 11.6369
R5225 GNDA.n2081 GNDA.n2080 11.6369
R5226 GNDA.n2080 GNDA.n538 11.6369
R5227 GNDA.n2095 GNDA.n532 11.6369
R5228 GNDA.n2096 GNDA.n2095 11.6369
R5229 GNDA.n2097 GNDA.n2096 11.6369
R5230 GNDA.n2097 GNDA.n528 11.6369
R5231 GNDA.n2103 GNDA.n528 11.6369
R5232 GNDA.n2104 GNDA.n2103 11.6369
R5233 GNDA.n2105 GNDA.n2104 11.6369
R5234 GNDA.n2105 GNDA.n524 11.6369
R5235 GNDA.n2112 GNDA.n524 11.6369
R5236 GNDA.n2113 GNDA.n2112 11.6369
R5237 GNDA.n2114 GNDA.n2113 11.6369
R5238 GNDA.n2123 GNDA.n2122 11.6369
R5239 GNDA.n2124 GNDA.n2123 11.6369
R5240 GNDA.n2124 GNDA.n518 11.6369
R5241 GNDA.n2131 GNDA.n518 11.6369
R5242 GNDA.n2132 GNDA.n2131 11.6369
R5243 GNDA.n2133 GNDA.n2132 11.6369
R5244 GNDA.n2139 GNDA.n515 11.6369
R5245 GNDA.n2140 GNDA.n2139 11.6369
R5246 GNDA.n2299 GNDA.n2298 11.6369
R5247 GNDA.n2300 GNDA.n2299 11.6369
R5248 GNDA.n2300 GNDA.n180 11.6369
R5249 GNDA.n2306 GNDA.n180 11.6369
R5250 GNDA.n2307 GNDA.n2306 11.6369
R5251 GNDA.n2308 GNDA.n2307 11.6369
R5252 GNDA.n2308 GNDA.n178 11.6369
R5253 GNDA.n2314 GNDA.n178 11.6369
R5254 GNDA.n2315 GNDA.n2314 11.6369
R5255 GNDA.n2316 GNDA.n2315 11.6369
R5256 GNDA.n2316 GNDA.n176 11.6369
R5257 GNDA.n496 GNDA.n495 11.6369
R5258 GNDA.n497 GNDA.n496 11.6369
R5259 GNDA.n497 GNDA.n491 11.6369
R5260 GNDA.n2157 GNDA.n491 11.6369
R5261 GNDA.n2158 GNDA.n2157 11.6369
R5262 GNDA.n2161 GNDA.n2158 11.6369
R5263 GNDA.n2160 GNDA.n2159 11.6369
R5264 GNDA.n2159 GNDA.n311 11.6369
R5265 GNDA.n2419 GNDA 11.5076
R5266 GNDA GNDA.n515 11.5076
R5267 GNDA GNDA.n2160 11.5076
R5268 GNDA.n2420 GNDA.n91 11.4026
R5269 GNDA.n2141 GNDA.n2140 11.4026
R5270 GNDA.n311 GNDA.n310 11.4026
R5271 GNDA.n1845 GNDA.n595 11.249
R5272 GNDA.n1443 GNDA.n1411 11.249
R5273 GNDA.n742 GNDA.n739 11.249
R5274 GNDA.n2069 GNDA.n2068 10.4732
R5275 GNDA.n2466 GNDA.n52 10.3161
R5276 GNDA.n1698 GNDA.n1626 9.78488
R5277 GNDA GNDA.n0 9.67325
R5278 GNDA.n2075 GNDA.n2074 9.65197
R5279 GNDA.n1694 GNDA.t213 9.6005
R5280 GNDA.n1694 GNDA.t214 9.6005
R5281 GNDA.n417 GNDA.t26 9.6005
R5282 GNDA.n417 GNDA.t289 9.6005
R5283 GNDA.n415 GNDA.t6 9.6005
R5284 GNDA.n415 GNDA.t60 9.6005
R5285 GNDA.n413 GNDA.t104 9.6005
R5286 GNDA.n413 GNDA.t12 9.6005
R5287 GNDA.n411 GNDA.t8 9.6005
R5288 GNDA.n411 GNDA.t14 9.6005
R5289 GNDA.n409 GNDA.t62 9.6005
R5290 GNDA.n409 GNDA.t93 9.6005
R5291 GNDA.n407 GNDA.t74 9.6005
R5292 GNDA.n407 GNDA.t342 9.6005
R5293 GNDA.n405 GNDA.t16 9.6005
R5294 GNDA.n405 GNDA.t331 9.6005
R5295 GNDA.n403 GNDA.t341 9.6005
R5296 GNDA.n403 GNDA.t120 9.6005
R5297 GNDA.n401 GNDA.t3 9.6005
R5298 GNDA.n401 GNDA.t47 9.6005
R5299 GNDA.n399 GNDA.t30 9.6005
R5300 GNDA.n399 GNDA.t145 9.6005
R5301 GNDA.n397 GNDA.t187 9.6005
R5302 GNDA.n397 GNDA.t184 9.6005
R5303 GNDA.n1627 GNDA.t208 9.6005
R5304 GNDA.n1627 GNDA.t216 9.6005
R5305 GNDA.n1696 GNDA.n1629 9.37925
R5306 GNDA.n2468 GNDA.n2467 9.3005
R5307 GNDA.n2146 GNDA.n508 9.27744
R5308 GNDA.n2424 GNDA.n104 9.27744
R5309 GNDA.n2145 GNDA.t90 8.73174
R5310 GNDA.n235 GNDA.n215 8.66313
R5311 GNDA.n2114 GNDA.n522 8.66313
R5312 GNDA.n176 GNDA.n174 8.66313
R5313 GNDA.n1242 GNDA.n257 8.53383
R5314 GNDA.n645 GNDA.n578 8.53383
R5315 GNDA.n657 GNDA.n182 8.53383
R5316 GNDA.n1570 GNDA.n623 8.53383
R5317 GNDA.n722 GNDA.n721 8.53383
R5318 GNDA.n538 GNDA.n537 8.53383
R5319 GNDA.n1668 GNDA.n1667 8.44175
R5320 GNDA.n2474 GNDA.t10 8.42962
R5321 GNDA.n1487 GNDA.n1406 8.35606
R5322 GNDA.n1304 GNDA.n648 8.35606
R5323 GNDA.n2203 GNDA.n283 8.35606
R5324 GNDA.n789 GNDA.n745 8.35606
R5325 GNDA.n954 GNDA.n705 8.35606
R5326 GNDA.n1113 GNDA.n1072 8.35606
R5327 GNDA.n1756 GNDA.n599 8.35606
R5328 GNDA.n2052 GNDA.n1926 8.35606
R5329 GNDA.n2326 GNDA.n139 8.35606
R5330 GNDA.n1699 GNDA.n1698 7.71925
R5331 GNDA.t88 GNDA.n2145 7.64034
R5332 GNDA.n396 GNDA.n1 7.28175
R5333 GNDA.n420 GNDA.n419 7.20362
R5334 GNDA.n2153 GNDA.n2152 7.09463
R5335 GNDA.n2168 GNDA.n2167 6.4005
R5336 GNDA.n2485 GNDA.n32 6.4005
R5337 GNDA.n395 GNDA.n33 6.4005
R5338 GNDA.t169 GNDA.n1702 6.14575
R5339 GNDA.t343 GNDA.t295 6.14575
R5340 GNDA.n1726 GNDA.t175 6.14575
R5341 GNDA.n1638 GNDA.t173 6.14575
R5342 GNDA.t268 GNDA.t71 6.14575
R5343 GNDA.t82 GNDA.n1636 6.14575
R5344 GNDA.n471 GNDA.n1 5.65675
R5345 GNDA.n422 GNDA.n420 5.563
R5346 GNDA.n546 GNDA.n0 5.02613
R5347 GNDA.n2146 GNDA.t148 4.91182
R5348 GNDA.n420 GNDA.n24 4.85988
R5349 GNDA GNDA.n2496 4.8133
R5350 GNDA.n1812 GNDA.n1811 4.6085
R5351 GNDA.n2021 GNDA.n2020 4.6085
R5352 GNDA.n2434 GNDA.n2433 4.6085
R5353 GNDA.n773 GNDA.n766 4.6085
R5354 GNDA.n1200 GNDA.n1199 4.6085
R5355 GNDA.n1097 GNDA.n514 4.6085
R5356 GNDA.n1544 GNDA.n1388 4.6085
R5357 GNDA.n1288 GNDA.n208 4.6085
R5358 GNDA.n2187 GNDA.n305 4.6085
R5359 GNDA.n1238 GNDA.n1211 4.55161
R5360 GNDA.n1895 GNDA.n576 4.55161
R5361 GNDA.n1566 GNDA.n624 4.55161
R5362 GNDA.n920 GNDA.n719 4.55161
R5363 GNDA.n2089 GNDA.n533 4.55161
R5364 GNDA.n2294 GNDA.n183 4.55161
R5365 GNDA.n1807 GNDA.n564 4.5061
R5366 GNDA.n2017 GNDA.n147 4.5061
R5367 GNDA.n768 GNDA.n710 4.5061
R5368 GNDA.n1198 GNDA.n1197 4.5061
R5369 GNDA.n1545 GNDA.n1386 4.5061
R5370 GNDA.n2288 GNDA.n2287 4.5061
R5371 GNDA.n2466 GNDA.n2465 4.5005
R5372 GNDA.n51 GNDA.n49 4.5005
R5373 GNDA.n2495 GNDA.n2494 4.5005
R5374 GNDA.n1698 GNDA.n1697 4.5005
R5375 GNDA.n1210 GNDA.n645 4.39646
R5376 GNDA.n257 GNDA.n256 4.39646
R5377 GNDA.n677 GNDA.n623 4.39646
R5378 GNDA.n721 GNDA.n555 4.39646
R5379 GNDA.n537 GNDA.n532 4.39646
R5380 GNDA.n2298 GNDA.n182 4.39646
R5381 GNDA.n1925 GNDA.n564 4.3525
R5382 GNDA.n2325 GNDA.n147 4.3525
R5383 GNDA.n710 GNDA.n707 4.3525
R5384 GNDA.n1197 GNDA.n1196 4.3525
R5385 GNDA.n1386 GNDA.n1385 4.3525
R5386 GNDA.n2287 GNDA.n2286 4.3525
R5387 GNDA.n2053 GNDA.n1925 4.3013
R5388 GNDA.n2327 GNDA.n2325 4.3013
R5389 GNDA.n953 GNDA.n707 4.3013
R5390 GNDA.n1196 GNDA.n1193 4.3013
R5391 GNDA.n1385 GNDA.n1384 4.3013
R5392 GNDA.n2286 GNDA.n2283 4.3013
R5393 GNDA.n1238 GNDA.n1237 4.26717
R5394 GNDA.n1237 GNDA.n1234 4.26717
R5395 GNDA.n1234 GNDA.n1233 4.26717
R5396 GNDA.n1233 GNDA.n1230 4.26717
R5397 GNDA.n1230 GNDA.n1229 4.26717
R5398 GNDA.n1229 GNDA.n1226 4.26717
R5399 GNDA.n1225 GNDA.n1222 4.26717
R5400 GNDA.n1222 GNDA.n1221 4.26717
R5401 GNDA.n1895 GNDA.n574 4.26717
R5402 GNDA.n1901 GNDA.n574 4.26717
R5403 GNDA.n1901 GNDA.n572 4.26717
R5404 GNDA.n1907 GNDA.n572 4.26717
R5405 GNDA.n1907 GNDA.n570 4.26717
R5406 GNDA.n1914 GNDA.n570 4.26717
R5407 GNDA.n568 GNDA.n566 4.26717
R5408 GNDA.n1921 GNDA.n566 4.26717
R5409 GNDA.n1566 GNDA.n1565 4.26717
R5410 GNDA.n1565 GNDA.n629 4.26717
R5411 GNDA.n1560 GNDA.n629 4.26717
R5412 GNDA.n1560 GNDA.n1559 4.26717
R5413 GNDA.n1559 GNDA.n1558 4.26717
R5414 GNDA.n1558 GNDA.n637 4.26717
R5415 GNDA.n1552 GNDA.n1551 4.26717
R5416 GNDA.n1551 GNDA.n1550 4.26717
R5417 GNDA.n920 GNDA.n718 4.26717
R5418 GNDA.n926 GNDA.n718 4.26717
R5419 GNDA.n926 GNDA.n716 4.26717
R5420 GNDA.n932 GNDA.n716 4.26717
R5421 GNDA.n932 GNDA.n714 4.26717
R5422 GNDA.n940 GNDA.n714 4.26717
R5423 GNDA.n712 GNDA.n709 4.26717
R5424 GNDA.n947 GNDA.n709 4.26717
R5425 GNDA.n2089 GNDA.n534 4.26717
R5426 GNDA.n1050 GNDA.n534 4.26717
R5427 GNDA.n1051 GNDA.n1050 4.26717
R5428 GNDA.n1056 GNDA.n1051 4.26717
R5429 GNDA.n1057 GNDA.n1056 4.26717
R5430 GNDA.n1062 GNDA.n1057 4.26717
R5431 GNDA.n1068 GNDA.n1063 4.26717
R5432 GNDA.n1070 GNDA.n1068 4.26717
R5433 GNDA.n2294 GNDA.n184 4.26717
R5434 GNDA.n261 GNDA.n184 4.26717
R5435 GNDA.n262 GNDA.n261 4.26717
R5436 GNDA.n267 GNDA.n262 4.26717
R5437 GNDA.n268 GNDA.n267 4.26717
R5438 GNDA.n273 GNDA.n268 4.26717
R5439 GNDA.n279 GNDA.n274 4.26717
R5440 GNDA.n281 GNDA.n279 4.26717
R5441 GNDA.n743 GNDA.n742 4.2501
R5442 GNDA.n1444 GNDA.n1443 4.2501
R5443 GNDA GNDA.n1225 4.21976
R5444 GNDA GNDA.n568 4.21976
R5445 GNDA.n1552 GNDA 4.21976
R5446 GNDA GNDA.n712 4.21976
R5447 GNDA.n1063 GNDA 4.21976
R5448 GNDA.n274 GNDA 4.21976
R5449 GNDA.t307 GNDA.t274 4.21506
R5450 GNDA.n2481 GNDA.t186 4.21506
R5451 GNDA.t253 GNDA.t246 4.21506
R5452 GNDA.n1845 GNDA.n1844 4.1477
R5453 GNDA.n1221 GNDA.n147 4.12494
R5454 GNDA.n1921 GNDA.n564 4.12494
R5455 GNDA.n1550 GNDA.n1386 4.12494
R5456 GNDA.n947 GNDA.n710 4.12494
R5457 GNDA.n1197 GNDA.n1070 4.12494
R5458 GNDA.n2287 GNDA.n281 4.12494
R5459 GNDA.t148 GNDA.t88 3.82042
R5460 GNDA.n1697 GNDA.n1696 3.813
R5461 GNDA.n1629 GNDA 3.68412
R5462 GNDA.n604 GNDA.n603 3.5845
R5463 GNDA.n1838 GNDA.n1837 3.5845
R5464 GNDA.n1833 GNDA.n605 3.5845
R5465 GNDA.n1832 GNDA.n608 3.5845
R5466 GNDA.n1597 GNDA.n1596 3.5845
R5467 GNDA.n1826 GNDA.n1825 3.5845
R5468 GNDA.n1821 GNDA.n1598 3.5845
R5469 GNDA.n1820 GNDA.n1602 3.5845
R5470 GNDA.n1737 GNDA.n1736 3.5845
R5471 GNDA.n2051 GNDA.n2050 3.5845
R5472 GNDA.n1929 GNDA.n1927 3.5845
R5473 GNDA.n2045 GNDA.n1931 3.5845
R5474 GNDA.n2044 GNDA.n1932 3.5845
R5475 GNDA.n2036 GNDA.n2035 3.5845
R5476 GNDA.n1937 GNDA.n1935 3.5845
R5477 GNDA.n2030 GNDA.n1939 3.5845
R5478 GNDA.n2029 GNDA.n1940 3.5845
R5479 GNDA.n1948 GNDA.n1947 3.5845
R5480 GNDA.n2346 GNDA.n141 3.5845
R5481 GNDA.n2345 GNDA.n142 3.5845
R5482 GNDA.n2332 GNDA.n2331 3.5845
R5483 GNDA.n2339 GNDA.n2338 3.5845
R5484 GNDA.n2333 GNDA.n123 3.5845
R5485 GNDA.n2413 GNDA.n2412 3.5845
R5486 GNDA.n2408 GNDA.n124 3.5845
R5487 GNDA.n2407 GNDA.n2404 3.5845
R5488 GNDA.n2403 GNDA.n89 3.5845
R5489 GNDA.n865 GNDA.n864 3.5845
R5490 GNDA.n748 GNDA.n746 3.5845
R5491 GNDA.n859 GNDA.n750 3.5845
R5492 GNDA.n858 GNDA.n751 3.5845
R5493 GNDA.n854 GNDA.n853 3.5845
R5494 GNDA.n757 GNDA.n755 3.5845
R5495 GNDA.n848 GNDA.n759 3.5845
R5496 GNDA.n847 GNDA.n760 3.5845
R5497 GNDA.n843 GNDA.n842 3.5845
R5498 GNDA.n987 GNDA.n955 3.5845
R5499 GNDA.n986 GNDA.n983 3.5845
R5500 GNDA.n982 GNDA.n956 3.5845
R5501 GNDA.n979 GNDA.n978 3.5845
R5502 GNDA.n974 GNDA.n957 3.5845
R5503 GNDA.n973 GNDA.n970 3.5845
R5504 GNDA.n969 GNDA.n961 3.5845
R5505 GNDA.n966 GNDA.n965 3.5845
R5506 GNDA.n1042 GNDA.n690 3.5845
R5507 GNDA.n1189 GNDA.n1188 3.5845
R5508 GNDA.n1076 GNDA.n1074 3.5845
R5509 GNDA.n1183 GNDA.n1078 3.5845
R5510 GNDA.n1182 GNDA.n1079 3.5845
R5511 GNDA.n1178 GNDA.n1177 3.5845
R5512 GNDA.n1085 GNDA.n1083 3.5845
R5513 GNDA.n1172 GNDA.n1087 3.5845
R5514 GNDA.n1171 GNDA.n1088 3.5845
R5515 GNDA.n1167 GNDA.n1166 3.5845
R5516 GNDA.n1483 GNDA.n1408 3.5845
R5517 GNDA.n1482 GNDA.n1409 3.5845
R5518 GNDA.n1478 GNDA.n1477 3.5845
R5519 GNDA.n1451 GNDA.n1449 3.5845
R5520 GNDA.n1472 GNDA.n1453 3.5845
R5521 GNDA.n1471 GNDA.n1454 3.5845
R5522 GNDA.n1467 GNDA.n1466 3.5845
R5523 GNDA.n1462 GNDA.n1459 3.5845
R5524 GNDA.n1461 GNDA.n1390 3.5845
R5525 GNDA.n1380 GNDA.n1379 3.5845
R5526 GNDA.n1268 GNDA.n1266 3.5845
R5527 GNDA.n1374 GNDA.n1270 3.5845
R5528 GNDA.n1373 GNDA.n1271 3.5845
R5529 GNDA.n1369 GNDA.n1368 3.5845
R5530 GNDA.n1277 GNDA.n1275 3.5845
R5531 GNDA.n1363 GNDA.n1279 3.5845
R5532 GNDA.n1362 GNDA.n1280 3.5845
R5533 GNDA.n1358 GNDA.n1357 3.5845
R5534 GNDA.n2279 GNDA.n2278 3.5845
R5535 GNDA.n287 GNDA.n285 3.5845
R5536 GNDA.n2273 GNDA.n289 3.5845
R5537 GNDA.n2272 GNDA.n290 3.5845
R5538 GNDA.n2268 GNDA.n2267 3.5845
R5539 GNDA.n296 GNDA.n294 3.5845
R5540 GNDA.n2262 GNDA.n298 3.5845
R5541 GNDA.n2261 GNDA.n299 3.5845
R5542 GNDA.n2257 GNDA.n2256 3.5845
R5543 GNDA.n2493 GNDA.n24 3.438
R5544 GNDA.n423 GNDA.t32 3.42907
R5545 GNDA.n423 GNDA.t327 3.42907
R5546 GNDA.n421 GNDA.t156 3.42907
R5547 GNDA.n421 GNDA.t51 3.42907
R5548 GNDA.n470 GNDA.t53 3.42907
R5549 GNDA.n470 GNDA.t70 3.42907
R5550 GNDA.n469 GNDA.t135 3.42907
R5551 GNDA.n469 GNDA.t131 3.42907
R5552 GNDA.n1844 GNDA.n599 3.3797
R5553 GNDA.n2053 GNDA.n2052 3.3797
R5554 GNDA.n2327 GNDA.n2326 3.3797
R5555 GNDA.n745 GNDA.n743 3.3797
R5556 GNDA.n954 GNDA.n953 3.3797
R5557 GNDA.n1193 GNDA.n1072 3.3797
R5558 GNDA.n1444 GNDA.n1406 3.3797
R5559 GNDA.n1384 GNDA.n648 3.3797
R5560 GNDA.n2283 GNDA.n283 3.3797
R5561 GNDA.n2494 GNDA.n2493 3.3755
R5562 GNDA.n2424 GNDA.t101 3.27472
R5563 GNDA.n105 GNDA.n99 3.2005
R5564 GNDA.n316 GNDA.n315 3.2005
R5565 GNDA.n1814 GNDA.n1813 2.8677
R5566 GNDA.n2023 GNDA.n2022 2.8677
R5567 GNDA.n2436 GNDA.n2435 2.8677
R5568 GNDA.n774 GNDA.n764 2.8677
R5569 GNDA.n1044 GNDA.n1043 2.8677
R5570 GNDA.n1098 GNDA.n1092 2.8677
R5571 GNDA.n1539 GNDA.n1538 2.8677
R5572 GNDA.n1289 GNDA.n1284 2.8677
R5573 GNDA.n2188 GNDA.n303 2.8677
R5574 GNDA.n1655 GNDA.n1653 2.34425
R5575 GNDA.n1663 GNDA.n1661 2.34425
R5576 GNDA.n1538 GNDA.n1537 2.31161
R5577 GNDA.n1290 GNDA.n1289 2.31161
R5578 GNDA.n2189 GNDA.n2188 2.31161
R5579 GNDA.n775 GNDA.n774 2.31161
R5580 GNDA.n1044 GNDA.n688 2.31161
R5581 GNDA.n1099 GNDA.n1098 2.31161
R5582 GNDA.n1813 GNDA.n1806 2.31161
R5583 GNDA.n2022 GNDA.n2015 2.31161
R5584 GNDA.n2435 GNDA.n90 2.31161
R5585 GNDA GNDA.n1529 1.95606
R5586 GNDA.n1292 GNDA 1.95606
R5587 GNDA.n2191 GNDA 1.95606
R5588 GNDA.n777 GNDA 1.95606
R5589 GNDA.n693 GNDA 1.95606
R5590 GNDA.n1101 GNDA 1.95606
R5591 GNDA GNDA.n1798 1.95606
R5592 GNDA GNDA.n2007 1.95606
R5593 GNDA.n127 GNDA 1.95606
R5594 GNDA.n1813 GNDA.n1812 1.7413
R5595 GNDA.n2022 GNDA.n2021 1.7413
R5596 GNDA.n2435 GNDA.n2434 1.7413
R5597 GNDA.n774 GNDA.n773 1.7413
R5598 GNDA.n1200 GNDA.n1044 1.7413
R5599 GNDA.n1098 GNDA.n1097 1.7413
R5600 GNDA.n1538 GNDA.n1388 1.7413
R5601 GNDA.n1289 GNDA.n1288 1.7413
R5602 GNDA.n2188 GNDA.n2187 1.7413
R5603 GNDA.n550 GNDA.n549 1.73362
R5604 GNDA.n2164 GNDA.n312 1.63761
R5605 GNDA.n2492 GNDA.n25 1.6005
R5606 GNDA.n440 GNDA.n436 1.6005
R5607 GNDA.n603 GNDA.n599 1.2293
R5608 GNDA.n2052 GNDA.n2051 1.2293
R5609 GNDA.n2326 GNDA.n141 1.2293
R5610 GNDA.n865 GNDA.n745 1.2293
R5611 GNDA.n955 GNDA.n954 1.2293
R5612 GNDA.n1189 GNDA.n1072 1.2293
R5613 GNDA.n1408 GNDA.n1406 1.2293
R5614 GNDA.n1380 GNDA.n648 1.2293
R5615 GNDA.n2279 GNDA.n283 1.2293
R5616 GNDA.n1811 GNDA.n1807 1.1781
R5617 GNDA.n2020 GNDA.n2017 1.1781
R5618 GNDA.n2433 GNDA.n91 1.1781
R5619 GNDA.n768 GNDA.n766 1.1781
R5620 GNDA.n1199 GNDA.n1198 1.1781
R5621 GNDA.n2141 GNDA.n514 1.1781
R5622 GNDA.n1545 GNDA.n1544 1.1781
R5623 GNDA.n2288 GNDA.n208 1.1781
R5624 GNDA.n310 GNDA.n305 1.1781
R5625 GNDA.n2069 GNDA.n541 1.16414
R5626 GNDA.n1838 GNDA.n604 1.0245
R5627 GNDA.n1837 GNDA.n605 1.0245
R5628 GNDA.n1833 GNDA.n1832 1.0245
R5629 GNDA.n1596 GNDA.n608 1.0245
R5630 GNDA.n1826 GNDA.n1597 1.0245
R5631 GNDA.n1825 GNDA.n1598 1.0245
R5632 GNDA.n1821 GNDA.n1820 1.0245
R5633 GNDA.n1736 GNDA.n1602 1.0245
R5634 GNDA.n1814 GNDA.n1737 1.0245
R5635 GNDA.n2050 GNDA.n1927 1.0245
R5636 GNDA.n1931 GNDA.n1929 1.0245
R5637 GNDA.n2045 GNDA.n2044 1.0245
R5638 GNDA.n2036 GNDA.n1932 1.0245
R5639 GNDA.n2035 GNDA.n1935 1.0245
R5640 GNDA.n1939 GNDA.n1937 1.0245
R5641 GNDA.n2030 GNDA.n2029 1.0245
R5642 GNDA.n1947 GNDA.n1940 1.0245
R5643 GNDA.n2023 GNDA.n1948 1.0245
R5644 GNDA.n2346 GNDA.n2345 1.0245
R5645 GNDA.n2331 GNDA.n142 1.0245
R5646 GNDA.n2339 GNDA.n2332 1.0245
R5647 GNDA.n2338 GNDA.n2333 1.0245
R5648 GNDA.n2413 GNDA.n123 1.0245
R5649 GNDA.n2412 GNDA.n124 1.0245
R5650 GNDA.n2408 GNDA.n2407 1.0245
R5651 GNDA.n2404 GNDA.n2403 1.0245
R5652 GNDA.n2436 GNDA.n89 1.0245
R5653 GNDA.n864 GNDA.n746 1.0245
R5654 GNDA.n750 GNDA.n748 1.0245
R5655 GNDA.n859 GNDA.n858 1.0245
R5656 GNDA.n854 GNDA.n751 1.0245
R5657 GNDA.n853 GNDA.n755 1.0245
R5658 GNDA.n759 GNDA.n757 1.0245
R5659 GNDA.n848 GNDA.n847 1.0245
R5660 GNDA.n843 GNDA.n760 1.0245
R5661 GNDA.n842 GNDA.n764 1.0245
R5662 GNDA.n987 GNDA.n986 1.0245
R5663 GNDA.n983 GNDA.n982 1.0245
R5664 GNDA.n979 GNDA.n956 1.0245
R5665 GNDA.n978 GNDA.n957 1.0245
R5666 GNDA.n974 GNDA.n973 1.0245
R5667 GNDA.n970 GNDA.n969 1.0245
R5668 GNDA.n966 GNDA.n961 1.0245
R5669 GNDA.n965 GNDA.n690 1.0245
R5670 GNDA.n1043 GNDA.n1042 1.0245
R5671 GNDA.n1188 GNDA.n1074 1.0245
R5672 GNDA.n1078 GNDA.n1076 1.0245
R5673 GNDA.n1183 GNDA.n1182 1.0245
R5674 GNDA.n1178 GNDA.n1079 1.0245
R5675 GNDA.n1177 GNDA.n1083 1.0245
R5676 GNDA.n1087 GNDA.n1085 1.0245
R5677 GNDA.n1172 GNDA.n1171 1.0245
R5678 GNDA.n1167 GNDA.n1088 1.0245
R5679 GNDA.n1166 GNDA.n1092 1.0245
R5680 GNDA.n1483 GNDA.n1482 1.0245
R5681 GNDA.n1478 GNDA.n1409 1.0245
R5682 GNDA.n1477 GNDA.n1449 1.0245
R5683 GNDA.n1453 GNDA.n1451 1.0245
R5684 GNDA.n1472 GNDA.n1471 1.0245
R5685 GNDA.n1467 GNDA.n1454 1.0245
R5686 GNDA.n1466 GNDA.n1459 1.0245
R5687 GNDA.n1462 GNDA.n1461 1.0245
R5688 GNDA.n1539 GNDA.n1390 1.0245
R5689 GNDA.n1379 GNDA.n1266 1.0245
R5690 GNDA.n1270 GNDA.n1268 1.0245
R5691 GNDA.n1374 GNDA.n1373 1.0245
R5692 GNDA.n1369 GNDA.n1271 1.0245
R5693 GNDA.n1368 GNDA.n1275 1.0245
R5694 GNDA.n1279 GNDA.n1277 1.0245
R5695 GNDA.n1363 GNDA.n1362 1.0245
R5696 GNDA.n1358 GNDA.n1280 1.0245
R5697 GNDA.n1357 GNDA.n1284 1.0245
R5698 GNDA.n2278 GNDA.n285 1.0245
R5699 GNDA.n289 GNDA.n287 1.0245
R5700 GNDA.n2273 GNDA.n2272 1.0245
R5701 GNDA.n2268 GNDA.n290 1.0245
R5702 GNDA.n2267 GNDA.n294 1.0245
R5703 GNDA.n298 GNDA.n296 1.0245
R5704 GNDA.n2262 GNDA.n2261 1.0245
R5705 GNDA.n2257 GNDA.n299 1.0245
R5706 GNDA.n2256 GNDA.n303 1.0245
R5707 GNDA.n2467 GNDA.n2466 0.65675
R5708 GNDA.n1653 GNDA.n1651 0.563
R5709 GNDA.n1657 GNDA.n1655 0.563
R5710 GNDA.n1659 GNDA.n1657 0.563
R5711 GNDA.n1661 GNDA.n1659 0.563
R5712 GNDA.n1665 GNDA.n1663 0.563
R5713 GNDA.n1667 GNDA.n1665 0.563
R5714 GNDA.n2453 GNDA.t102 0.467591
R5715 GNDA.n363 GNDA.t153 0.467591
R5716 GNDA.n547 GNDA.n546 0.41175
R5717 GNDA.n2495 GNDA.n1 0.359875
R5718 GNDA.n398 GNDA.n396 0.359875
R5719 GNDA.n17 GNDA.n15 0.34425
R5720 GNDA.n19 GNDA.n17 0.34425
R5721 GNDA.n21 GNDA.n19 0.34425
R5722 GNDA.n23 GNDA.n21 0.34425
R5723 GNDA.n12 GNDA.n10 0.34425
R5724 GNDA.n10 GNDA.n8 0.34425
R5725 GNDA.n8 GNDA.n6 0.34425
R5726 GNDA.n6 GNDA.n4 0.34425
R5727 GNDA.n49 GNDA.n45 0.34425
R5728 GNDA.n49 GNDA.n48 0.34425
R5729 GNDA.n400 GNDA.n398 0.34425
R5730 GNDA.n402 GNDA.n400 0.34425
R5731 GNDA.n404 GNDA.n402 0.34425
R5732 GNDA.n406 GNDA.n404 0.34425
R5733 GNDA.n408 GNDA.n406 0.34425
R5734 GNDA.n410 GNDA.n408 0.34425
R5735 GNDA.n412 GNDA.n410 0.34425
R5736 GNDA.n414 GNDA.n412 0.34425
R5737 GNDA.n416 GNDA.n414 0.34425
R5738 GNDA.n418 GNDA.n416 0.34425
R5739 GNDA.n472 GNDA.n471 0.313
R5740 GNDA.n424 GNDA.n422 0.313
R5741 GNDA.n548 GNDA.n547 0.311875
R5742 GNDA.n1648 GNDA.n1629 0.276625
R5743 GNDA.n1668 GNDA.n1648 0.22375
R5744 GNDA.n2467 GNDA.n51 0.188
R5745 GNDA.n419 GNDA.n418 0.188
R5746 GNDA GNDA.n2418 0.129793
R5747 GNDA.n2133 GNDA 0.129793
R5748 GNDA.n2161 GNDA 0.129793
R5749 GNDA.n1669 GNDA.n1668 0.100375
R5750 GNDA.n549 GNDA.n548 0.076875
R5751 GNDA.n1211 GNDA.n257 0.0479074
R5752 GNDA.n1226 GNDA 0.0479074
R5753 GNDA.n645 GNDA.n576 0.0479074
R5754 GNDA.n1914 GNDA 0.0479074
R5755 GNDA.n624 GNDA.n623 0.0479074
R5756 GNDA GNDA.n637 0.0479074
R5757 GNDA.n721 GNDA.n719 0.0479074
R5758 GNDA.n940 GNDA 0.0479074
R5759 GNDA.n537 GNDA.n533 0.0479074
R5760 GNDA GNDA.n1062 0.0479074
R5761 GNDA.n183 GNDA.n182 0.0479074
R5762 GNDA GNDA.n273 0.0479074
R5763 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.n3 110.171
R5764 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.n2 110.171
R5765 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.n4 109.828
R5766 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.n5 109.828
R5767 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 108.966
R5768 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n14 108.965
R5769 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 107.716
R5770 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 107.716
R5771 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 107.716
R5772 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.n1 105.314
R5773 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n8 103.216
R5774 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5775 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5776 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5777 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5778 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5779 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5780 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5781 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5782 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5783 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5784 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5785 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5786 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5787 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5788 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5789 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5790 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5791 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5792 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5793 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5794 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5795 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5796 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.n6 4.5005
R5797 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 4.5005
R5798 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.n13 3.6255
R5799 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n11 1.2505
R5800 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5801 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.n0 0.688
R5802 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n7 0.51925
R5803 VOUT-.n14 VOUT-.n6 141.722
R5804 VOUT-.n9 VOUT-.n7 141.722
R5805 VOUT-.n13 VOUT-.n12 141.161
R5806 VOUT-.n11 VOUT-.n10 141.161
R5807 VOUT-.n9 VOUT-.n8 141.161
R5808 VOUT-.n16 VOUT-.n15 136.661
R5809 VOUT-.n5 VOUT-.t4 113.129
R5810 VOUT-.n2 VOUT-.n0 90.9636
R5811 VOUT-.n4 VOUT-.n3 90.3386
R5812 VOUT-.n2 VOUT-.n1 90.3386
R5813 VOUT-.n96 VOUT-.n16 15.0943
R5814 VOUT-.n96 VOUT-.n95 11.6871
R5815 VOUT-.n15 VOUT-.t5 6.56717
R5816 VOUT-.n15 VOUT-.t8 6.56717
R5817 VOUT-.n12 VOUT-.t7 6.56717
R5818 VOUT-.n12 VOUT-.t12 6.56717
R5819 VOUT-.n10 VOUT-.t2 6.56717
R5820 VOUT-.n10 VOUT-.t11 6.56717
R5821 VOUT-.n8 VOUT-.t0 6.56717
R5822 VOUT-.n8 VOUT-.t9 6.56717
R5823 VOUT-.n7 VOUT-.t13 6.56717
R5824 VOUT-.n7 VOUT-.t15 6.56717
R5825 VOUT-.n6 VOUT-.t14 6.56717
R5826 VOUT-.n6 VOUT-.t10 6.56717
R5827 VOUT- VOUT-.n96 6.48488
R5828 VOUT-.n43 VOUT-.t85 4.8295
R5829 VOUT-.n45 VOUT-.t131 4.8295
R5830 VOUT-.n47 VOUT-.t31 4.8295
R5831 VOUT-.n49 VOUT-.t62 4.8295
R5832 VOUT-.n51 VOUT-.t114 4.8295
R5833 VOUT-.n63 VOUT-.t40 4.8295
R5834 VOUT-.n65 VOUT-.t34 4.8295
R5835 VOUT-.n66 VOUT-.t136 4.8295
R5836 VOUT-.n68 VOUT-.t70 4.8295
R5837 VOUT-.n69 VOUT-.t36 4.8295
R5838 VOUT-.n71 VOUT-.t95 4.8295
R5839 VOUT-.n72 VOUT-.t66 4.8295
R5840 VOUT-.n74 VOUT-.t55 4.8295
R5841 VOUT-.n75 VOUT-.t29 4.8295
R5842 VOUT-.n77 VOUT-.t91 4.8295
R5843 VOUT-.n78 VOUT-.t58 4.8295
R5844 VOUT-.n80 VOUT-.t49 4.8295
R5845 VOUT-.n81 VOUT-.t20 4.8295
R5846 VOUT-.n83 VOUT-.t148 4.8295
R5847 VOUT-.n84 VOUT-.t122 4.8295
R5848 VOUT-.n86 VOUT-.t44 4.8295
R5849 VOUT-.n87 VOUT-.t152 4.8295
R5850 VOUT-.n89 VOUT-.t142 4.8295
R5851 VOUT-.n90 VOUT-.t116 4.8295
R5852 VOUT-.n17 VOUT-.t108 4.8295
R5853 VOUT-.n29 VOUT-.t28 4.8295
R5854 VOUT-.n31 VOUT-.t24 4.8295
R5855 VOUT-.n32 VOUT-.t129 4.8295
R5856 VOUT-.n34 VOUT-.t61 4.8295
R5857 VOUT-.n35 VOUT-.t32 4.8295
R5858 VOUT-.n37 VOUT-.t100 4.8295
R5859 VOUT-.n38 VOUT-.t71 4.8295
R5860 VOUT-.n40 VOUT-.t69 4.8295
R5861 VOUT-.n41 VOUT-.t35 4.8295
R5862 VOUT-.n92 VOUT-.t77 4.8295
R5863 VOUT-.n56 VOUT-.t26 4.8154
R5864 VOUT-.n55 VOUT-.t59 4.8154
R5865 VOUT-.n54 VOUT-.t37 4.8154
R5866 VOUT-.n53 VOUT-.t81 4.8154
R5867 VOUT-.n62 VOUT-.t132 4.806
R5868 VOUT-.n61 VOUT-.t115 4.806
R5869 VOUT-.n60 VOUT-.t146 4.806
R5870 VOUT-.n59 VOUT-.t46 4.806
R5871 VOUT-.n58 VOUT-.t87 4.806
R5872 VOUT-.n57 VOUT-.t65 4.806
R5873 VOUT-.n56 VOUT-.t102 4.806
R5874 VOUT-.n55 VOUT-.t134 4.806
R5875 VOUT-.n54 VOUT-.t120 4.806
R5876 VOUT-.n53 VOUT-.t155 4.806
R5877 VOUT-.n28 VOUT-.t48 4.806
R5878 VOUT-.n27 VOUT-.t92 4.806
R5879 VOUT-.n26 VOUT-.t42 4.806
R5880 VOUT-.n25 VOUT-.t130 4.806
R5881 VOUT-.n24 VOUT-.t84 4.806
R5882 VOUT-.n23 VOUT-.t125 4.806
R5883 VOUT-.n22 VOUT-.t74 4.806
R5884 VOUT-.n21 VOUT-.t23 4.806
R5885 VOUT-.n20 VOUT-.t64 4.806
R5886 VOUT-.n19 VOUT-.t150 4.806
R5887 VOUT-.n44 VOUT-.t96 4.5005
R5888 VOUT-.n43 VOUT-.t57 4.5005
R5889 VOUT-.n45 VOUT-.t104 4.5005
R5890 VOUT-.n46 VOUT-.t73 4.5005
R5891 VOUT-.n47 VOUT-.t138 4.5005
R5892 VOUT-.n48 VOUT-.t107 4.5005
R5893 VOUT-.n49 VOUT-.t41 4.5005
R5894 VOUT-.n50 VOUT-.t143 4.5005
R5895 VOUT-.n51 VOUT-.t21 4.5005
R5896 VOUT-.n52 VOUT-.t126 4.5005
R5897 VOUT-.n53 VOUT-.t119 4.5005
R5898 VOUT-.n54 VOUT-.t82 4.5005
R5899 VOUT-.n55 VOUT-.t97 4.5005
R5900 VOUT-.n56 VOUT-.t63 4.5005
R5901 VOUT-.n57 VOUT-.t27 4.5005
R5902 VOUT-.n58 VOUT-.t45 4.5005
R5903 VOUT-.n59 VOUT-.t144 4.5005
R5904 VOUT-.n60 VOUT-.t112 4.5005
R5905 VOUT-.n61 VOUT-.t76 4.5005
R5906 VOUT-.n62 VOUT-.t93 4.5005
R5907 VOUT-.n64 VOUT-.t56 4.5005
R5908 VOUT-.n63 VOUT-.t19 4.5005
R5909 VOUT-.n65 VOUT-.t52 4.5005
R5910 VOUT-.n67 VOUT-.t156 4.5005
R5911 VOUT-.n66 VOUT-.t121 4.5005
R5912 VOUT-.n68 VOUT-.t89 4.5005
R5913 VOUT-.n70 VOUT-.t50 4.5005
R5914 VOUT-.n69 VOUT-.t151 4.5005
R5915 VOUT-.n71 VOUT-.t43 4.5005
R5916 VOUT-.n73 VOUT-.t145 4.5005
R5917 VOUT-.n72 VOUT-.t118 4.5005
R5918 VOUT-.n74 VOUT-.t141 4.5005
R5919 VOUT-.n76 VOUT-.t111 4.5005
R5920 VOUT-.n75 VOUT-.t80 4.5005
R5921 VOUT-.n77 VOUT-.t39 4.5005
R5922 VOUT-.n79 VOUT-.t139 4.5005
R5923 VOUT-.n78 VOUT-.t109 4.5005
R5924 VOUT-.n80 VOUT-.t135 4.5005
R5925 VOUT-.n82 VOUT-.t103 4.5005
R5926 VOUT-.n81 VOUT-.t72 4.5005
R5927 VOUT-.n83 VOUT-.t99 4.5005
R5928 VOUT-.n85 VOUT-.t68 4.5005
R5929 VOUT-.n84 VOUT-.t33 4.5005
R5930 VOUT-.n86 VOUT-.t133 4.5005
R5931 VOUT-.n88 VOUT-.t98 4.5005
R5932 VOUT-.n87 VOUT-.t67 4.5005
R5933 VOUT-.n89 VOUT-.t94 4.5005
R5934 VOUT-.n91 VOUT-.t60 4.5005
R5935 VOUT-.n90 VOUT-.t30 4.5005
R5936 VOUT-.n18 VOUT-.t101 4.5005
R5937 VOUT-.n17 VOUT-.t149 4.5005
R5938 VOUT-.n19 VOUT-.t88 4.5005
R5939 VOUT-.n20 VOUT-.t51 4.5005
R5940 VOUT-.n21 VOUT-.t137 4.5005
R5941 VOUT-.n22 VOUT-.t106 4.5005
R5942 VOUT-.n23 VOUT-.t75 4.5005
R5943 VOUT-.n24 VOUT-.t25 4.5005
R5944 VOUT-.n25 VOUT-.t128 4.5005
R5945 VOUT-.n26 VOUT-.t90 4.5005
R5946 VOUT-.n27 VOUT-.t54 4.5005
R5947 VOUT-.n28 VOUT-.t140 4.5005
R5948 VOUT-.n30 VOUT-.t110 4.5005
R5949 VOUT-.n29 VOUT-.t79 4.5005
R5950 VOUT-.n31 VOUT-.t113 4.5005
R5951 VOUT-.n33 VOUT-.t78 4.5005
R5952 VOUT-.n32 VOUT-.t38 4.5005
R5953 VOUT-.n34 VOUT-.t147 4.5005
R5954 VOUT-.n36 VOUT-.t117 4.5005
R5955 VOUT-.n35 VOUT-.t83 4.5005
R5956 VOUT-.n37 VOUT-.t47 4.5005
R5957 VOUT-.n39 VOUT-.t153 4.5005
R5958 VOUT-.n38 VOUT-.t123 4.5005
R5959 VOUT-.n40 VOUT-.t154 4.5005
R5960 VOUT-.n42 VOUT-.t124 4.5005
R5961 VOUT-.n41 VOUT-.t86 4.5005
R5962 VOUT-.n95 VOUT-.t105 4.5005
R5963 VOUT-.n94 VOUT-.t53 4.5005
R5964 VOUT-.n93 VOUT-.t22 4.5005
R5965 VOUT-.n92 VOUT-.t127 4.5005
R5966 VOUT-.n16 VOUT-.n14 4.5005
R5967 VOUT-.n3 VOUT-.t18 3.42907
R5968 VOUT-.n3 VOUT-.t16 3.42907
R5969 VOUT-.n1 VOUT-.t3 3.42907
R5970 VOUT-.n1 VOUT-.t1 3.42907
R5971 VOUT-.n0 VOUT-.t17 3.42907
R5972 VOUT-.n0 VOUT-.t6 3.42907
R5973 VOUT- VOUT-.n5 1.54738
R5974 VOUT-.n5 VOUT-.n4 1.07862
R5975 VOUT-.n4 VOUT-.n2 0.6255
R5976 VOUT-.n11 VOUT-.n9 0.563
R5977 VOUT-.n13 VOUT-.n11 0.563
R5978 VOUT-.n14 VOUT-.n13 0.563
R5979 VOUT-.n44 VOUT-.n43 0.3295
R5980 VOUT-.n46 VOUT-.n45 0.3295
R5981 VOUT-.n48 VOUT-.n47 0.3295
R5982 VOUT-.n50 VOUT-.n49 0.3295
R5983 VOUT-.n52 VOUT-.n51 0.3295
R5984 VOUT-.n54 VOUT-.n53 0.3295
R5985 VOUT-.n55 VOUT-.n54 0.3295
R5986 VOUT-.n56 VOUT-.n55 0.3295
R5987 VOUT-.n57 VOUT-.n56 0.3295
R5988 VOUT-.n58 VOUT-.n57 0.3295
R5989 VOUT-.n59 VOUT-.n58 0.3295
R5990 VOUT-.n60 VOUT-.n59 0.3295
R5991 VOUT-.n61 VOUT-.n60 0.3295
R5992 VOUT-.n62 VOUT-.n61 0.3295
R5993 VOUT-.n64 VOUT-.n62 0.3295
R5994 VOUT-.n64 VOUT-.n63 0.3295
R5995 VOUT-.n67 VOUT-.n65 0.3295
R5996 VOUT-.n67 VOUT-.n66 0.3295
R5997 VOUT-.n70 VOUT-.n68 0.3295
R5998 VOUT-.n70 VOUT-.n69 0.3295
R5999 VOUT-.n73 VOUT-.n71 0.3295
R6000 VOUT-.n73 VOUT-.n72 0.3295
R6001 VOUT-.n76 VOUT-.n74 0.3295
R6002 VOUT-.n76 VOUT-.n75 0.3295
R6003 VOUT-.n79 VOUT-.n77 0.3295
R6004 VOUT-.n79 VOUT-.n78 0.3295
R6005 VOUT-.n82 VOUT-.n80 0.3295
R6006 VOUT-.n82 VOUT-.n81 0.3295
R6007 VOUT-.n85 VOUT-.n83 0.3295
R6008 VOUT-.n85 VOUT-.n84 0.3295
R6009 VOUT-.n88 VOUT-.n86 0.3295
R6010 VOUT-.n88 VOUT-.n87 0.3295
R6011 VOUT-.n91 VOUT-.n89 0.3295
R6012 VOUT-.n91 VOUT-.n90 0.3295
R6013 VOUT-.n18 VOUT-.n17 0.3295
R6014 VOUT-.n20 VOUT-.n19 0.3295
R6015 VOUT-.n21 VOUT-.n20 0.3295
R6016 VOUT-.n22 VOUT-.n21 0.3295
R6017 VOUT-.n23 VOUT-.n22 0.3295
R6018 VOUT-.n24 VOUT-.n23 0.3295
R6019 VOUT-.n25 VOUT-.n24 0.3295
R6020 VOUT-.n26 VOUT-.n25 0.3295
R6021 VOUT-.n27 VOUT-.n26 0.3295
R6022 VOUT-.n28 VOUT-.n27 0.3295
R6023 VOUT-.n30 VOUT-.n28 0.3295
R6024 VOUT-.n30 VOUT-.n29 0.3295
R6025 VOUT-.n33 VOUT-.n31 0.3295
R6026 VOUT-.n33 VOUT-.n32 0.3295
R6027 VOUT-.n36 VOUT-.n34 0.3295
R6028 VOUT-.n36 VOUT-.n35 0.3295
R6029 VOUT-.n39 VOUT-.n37 0.3295
R6030 VOUT-.n39 VOUT-.n38 0.3295
R6031 VOUT-.n42 VOUT-.n40 0.3295
R6032 VOUT-.n42 VOUT-.n41 0.3295
R6033 VOUT-.n95 VOUT-.n94 0.3295
R6034 VOUT-.n94 VOUT-.n93 0.3295
R6035 VOUT-.n93 VOUT-.n92 0.3295
R6036 VOUT-.n60 VOUT-.n46 0.306
R6037 VOUT-.n59 VOUT-.n48 0.306
R6038 VOUT-.n58 VOUT-.n50 0.306
R6039 VOUT-.n57 VOUT-.n52 0.306
R6040 VOUT-.n64 VOUT-.n44 0.2825
R6041 VOUT-.n67 VOUT-.n64 0.2825
R6042 VOUT-.n70 VOUT-.n67 0.2825
R6043 VOUT-.n73 VOUT-.n70 0.2825
R6044 VOUT-.n76 VOUT-.n73 0.2825
R6045 VOUT-.n79 VOUT-.n76 0.2825
R6046 VOUT-.n82 VOUT-.n79 0.2825
R6047 VOUT-.n85 VOUT-.n82 0.2825
R6048 VOUT-.n88 VOUT-.n85 0.2825
R6049 VOUT-.n91 VOUT-.n88 0.2825
R6050 VOUT-.n30 VOUT-.n18 0.2825
R6051 VOUT-.n33 VOUT-.n30 0.2825
R6052 VOUT-.n36 VOUT-.n33 0.2825
R6053 VOUT-.n39 VOUT-.n36 0.2825
R6054 VOUT-.n42 VOUT-.n39 0.2825
R6055 VOUT-.n93 VOUT-.n42 0.2825
R6056 VOUT-.n93 VOUT-.n91 0.2825
R6057 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t138 48.958
R6058 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.922875
R6059 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1603
R6060 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1603
R6061 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1603
R6062 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1603
R6063 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R6064 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1603
R6065 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R6066 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.1603
R6067 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1603
R6068 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R6069 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1603
R6070 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1603
R6071 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R6072 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.1603
R6073 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1603
R6074 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1603
R6075 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1603
R6076 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.1603
R6077 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R6078 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R6079 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.1603
R6080 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1603
R6081 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R6082 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R6083 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1603
R6084 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1603
R6085 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1603
R6086 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R6087 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1603
R6088 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.1603
R6089 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R6090 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1603
R6091 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R6092 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1603
R6093 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.1603
R6094 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1603
R6095 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1603
R6096 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1603
R6097 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1603
R6098 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.1603
R6099 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1603
R6100 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R6101 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.1603
R6102 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R6103 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R6104 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1603
R6105 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1603
R6106 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R6107 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.1603
R6108 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1603
R6109 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R6110 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1603
R6111 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.1603
R6112 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R6113 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R6114 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R6115 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R6116 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.1603
R6117 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.159278
R6118 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R6119 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R6120 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R6121 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R6122 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R6123 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R6124 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R6125 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R6126 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R6127 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R6128 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.159278
R6129 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.159278
R6130 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.159278
R6131 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.159278
R6132 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.159278
R6133 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.159278
R6134 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.159278
R6135 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.159278
R6136 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.159278
R6137 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.159278
R6138 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.159278
R6139 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.159278
R6140 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.159278
R6141 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.159278
R6142 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.159278
R6143 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.159278
R6144 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.137822
R6145 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1368
R6146 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1368
R6147 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1368
R6148 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1368
R6149 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.1368
R6150 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.1368
R6151 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1368
R6152 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1368
R6153 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R6154 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1368
R6155 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R6156 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1368
R6157 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1368
R6158 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1368
R6159 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R6160 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1368
R6161 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.1368
R6162 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1368
R6163 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1368
R6164 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.1368
R6165 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.1368
R6166 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.1368
R6167 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.1368
R6168 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.1368
R6169 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1368
R6170 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1368
R6171 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1368
R6172 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R6173 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1368
R6174 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1368
R6175 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.1368
R6176 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.114322
R6177 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R6178 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R6179 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R6180 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.1133
R6181 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.1133
R6182 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.1133
R6183 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.1133
R6184 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.1133
R6185 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.1133
R6186 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R6187 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R6188 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R6189 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R6190 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R6191 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R6192 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R6193 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R6194 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R6195 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R6196 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.00152174
R6197 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R6198 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.00152174
R6199 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.00152174
R6200 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.00152174
R6201 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.00152174
R6202 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.00152174
R6203 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.00152174
R6204 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.00152174
R6205 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.00152174
R6206 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R6207 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.00152174
R6208 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.00152174
R6209 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.00152174
R6210 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.00152174
R6211 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.00152174
R6212 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.00152174
R6213 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.00152174
R6214 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.00152174
R6215 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.00152174
R6216 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.00152174
R6217 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.00152174
R6218 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.00152174
R6219 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R6220 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 0.00152174
R6221 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.00152174
R6222 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.00152174
R6223 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.00152174
R6224 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R6225 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R6226 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.00152174
R6227 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.00152174
R6228 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.00152174
R6229 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.00152174
R6230 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.00152174
R6231 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R6232 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 627.971
R6233 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 626.721
R6234 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 622.221
R6235 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 289.2
R6236 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 289.2
R6237 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 222.751
R6238 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 208.468
R6239 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 208.468
R6240 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 176.733
R6241 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 176.733
R6242 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 176.733
R6243 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 176.733
R6244 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 176.733
R6245 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 152
R6246 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 152
R6247 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 112.468
R6248 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 112.468
R6249 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R6250 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R6251 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 112.468
R6252 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R6253 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R6254 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 112.468
R6255 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 78.8005
R6256 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 78.8005
R6257 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R6258 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R6259 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R6260 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R6261 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R6262 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 48.0005
R6263 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 48.0005
R6264 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 48.0005
R6265 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 48.0005
R6266 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R6267 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 45.5227
R6268 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 45.5227
R6269 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 45.5227
R6270 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 45.5227
R6271 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 14.7693
R6272 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 14.0818
R6273 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 5.7505
R6274 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 5.5005
R6275 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t12 662.393
R6276 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 631.188
R6277 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n3 626.894
R6278 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 626.894
R6279 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 222.268
R6280 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 222.268
R6281 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n4 217.768
R6282 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t4 78.8005
R6283 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R6284 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R6285 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R6286 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t10 78.8005
R6287 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R6288 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R6289 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t11 48.0005
R6290 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R6291 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t5 48.0005
R6292 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R6293 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R6294 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 6.8755
R6295 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 5.188
R6296 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n2 0.7505
R6297 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 0.688
R6298 bgr_0.Vbe2.n125 bgr_0.Vbe2.t0 162.458
R6299 bgr_0.Vbe2.n142 bgr_0.Vbe2.n1 83.5719
R6300 bgr_0.Vbe2.n134 bgr_0.Vbe2.n2 83.5719
R6301 bgr_0.Vbe2.n136 bgr_0.Vbe2.n135 83.5719
R6302 bgr_0.Vbe2.n128 bgr_0.Vbe2.n7 83.5719
R6303 bgr_0.Vbe2.n120 bgr_0.Vbe2.n8 83.5719
R6304 bgr_0.Vbe2.n122 bgr_0.Vbe2.n121 83.5719
R6305 bgr_0.Vbe2.n114 bgr_0.Vbe2.n12 83.5719
R6306 bgr_0.Vbe2.n109 bgr_0.Vbe2.n13 83.5719
R6307 bgr_0.Vbe2.n51 bgr_0.Vbe2.n50 83.5719
R6308 bgr_0.Vbe2.n49 bgr_0.Vbe2.n48 83.5719
R6309 bgr_0.Vbe2.n47 bgr_0.Vbe2.n46 83.5719
R6310 bgr_0.Vbe2.n65 bgr_0.Vbe2.n64 83.5719
R6311 bgr_0.Vbe2.n63 bgr_0.Vbe2.n62 83.5719
R6312 bgr_0.Vbe2.n33 bgr_0.Vbe2.n32 83.5719
R6313 bgr_0.Vbe2.n73 bgr_0.Vbe2.n72 83.5719
R6314 bgr_0.Vbe2.n28 bgr_0.Vbe2.n26 83.5719
R6315 bgr_0.Vbe2.n78 bgr_0.Vbe2.n25 83.5719
R6316 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 83.5719
R6317 bgr_0.Vbe2.n23 bgr_0.Vbe2.n22 83.5719
R6318 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 83.5719
R6319 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 83.5719
R6320 bgr_0.Vbe2.n97 bgr_0.Vbe2.n96 83.5719
R6321 bgr_0.Vbe2.n59 bgr_0.Vbe2.n32 73.8495
R6322 bgr_0.Vbe2.n144 bgr_0.Vbe2.n1 73.3165
R6323 bgr_0.Vbe2.n130 bgr_0.Vbe2.n7 73.3165
R6324 bgr_0.Vbe2.n116 bgr_0.Vbe2.n12 73.3165
R6325 bgr_0.Vbe2.n50 bgr_0.Vbe2.n42 73.3165
R6326 bgr_0.Vbe2.n72 bgr_0.Vbe2.n71 73.3165
R6327 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 73.3165
R6328 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 73.3165
R6329 bgr_0.Vbe2.n135 bgr_0.Vbe2.n133 73.19
R6330 bgr_0.Vbe2.n121 bgr_0.Vbe2.n119 73.19
R6331 bgr_0.Vbe2.n47 bgr_0.Vbe2.n45 73.19
R6332 bgr_0.Vbe2.n64 bgr_0.Vbe2.n29 73.19
R6333 bgr_0.Vbe2.n80 bgr_0.Vbe2.n25 73.19
R6334 bgr_0.Vbe2.n97 bgr_0.Vbe2.n19 73.19
R6335 bgr_0.Vbe2.n110 bgr_0.Vbe2.t5 65.0299
R6336 bgr_0.Vbe2.t7 bgr_0.Vbe2.n20 65.0299
R6337 bgr_0.Vbe2.n134 bgr_0.Vbe2.n1 26.074
R6338 bgr_0.Vbe2.n120 bgr_0.Vbe2.n7 26.074
R6339 bgr_0.Vbe2.n109 bgr_0.Vbe2.n12 26.074
R6340 bgr_0.Vbe2.n50 bgr_0.Vbe2.n49 26.074
R6341 bgr_0.Vbe2.n63 bgr_0.Vbe2.n32 26.074
R6342 bgr_0.Vbe2.n72 bgr_0.Vbe2.n28 26.074
R6343 bgr_0.Vbe2.n85 bgr_0.Vbe2.n23 26.074
R6344 bgr_0.Vbe2.n101 bgr_0.Vbe2.n99 26.074
R6345 bgr_0.Vbe2.n135 bgr_0.Vbe2.t1 25.7843
R6346 bgr_0.Vbe2.n121 bgr_0.Vbe2.t8 25.7843
R6347 bgr_0.Vbe2.t3 bgr_0.Vbe2.n47 25.7843
R6348 bgr_0.Vbe2.n64 bgr_0.Vbe2.t4 25.7843
R6349 bgr_0.Vbe2.t2 bgr_0.Vbe2.n25 25.7843
R6350 bgr_0.Vbe2.t6 bgr_0.Vbe2.n97 25.7843
R6351 bgr_0.Vbe2.n103 bgr_0.Vbe2.n91 9.3005
R6352 bgr_0.Vbe2.n91 bgr_0.Vbe2.n17 9.3005
R6353 bgr_0.Vbe2.n91 bgr_0.Vbe2.n18 9.3005
R6354 bgr_0.Vbe2.n107 bgr_0.Vbe2.n91 9.3005
R6355 bgr_0.Vbe2.n93 bgr_0.Vbe2.n17 9.3005
R6356 bgr_0.Vbe2.n93 bgr_0.Vbe2.n18 9.3005
R6357 bgr_0.Vbe2.n93 bgr_0.Vbe2.n15 9.3005
R6358 bgr_0.Vbe2.n107 bgr_0.Vbe2.n93 9.3005
R6359 bgr_0.Vbe2.n108 bgr_0.Vbe2.n17 9.3005
R6360 bgr_0.Vbe2.n108 bgr_0.Vbe2.n16 9.3005
R6361 bgr_0.Vbe2.n108 bgr_0.Vbe2.n18 9.3005
R6362 bgr_0.Vbe2.n108 bgr_0.Vbe2.n15 9.3005
R6363 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 9.3005
R6364 bgr_0.Vbe2.n107 bgr_0.Vbe2.n95 9.3005
R6365 bgr_0.Vbe2.n95 bgr_0.Vbe2.n15 9.3005
R6366 bgr_0.Vbe2.n95 bgr_0.Vbe2.n18 9.3005
R6367 bgr_0.Vbe2.n95 bgr_0.Vbe2.n16 9.3005
R6368 bgr_0.Vbe2.n107 bgr_0.Vbe2.n90 9.3005
R6369 bgr_0.Vbe2.n90 bgr_0.Vbe2.n15 9.3005
R6370 bgr_0.Vbe2.n90 bgr_0.Vbe2.n18 9.3005
R6371 bgr_0.Vbe2.n90 bgr_0.Vbe2.n16 9.3005
R6372 bgr_0.Vbe2.n103 bgr_0.Vbe2.n90 9.3005
R6373 bgr_0.Vbe2.n106 bgr_0.Vbe2.n17 9.3005
R6374 bgr_0.Vbe2.n106 bgr_0.Vbe2.n16 9.3005
R6375 bgr_0.Vbe2.n106 bgr_0.Vbe2.n18 9.3005
R6376 bgr_0.Vbe2.n107 bgr_0.Vbe2.n106 9.3005
R6377 bgr_0.Vbe2.n56 bgr_0.Vbe2.n55 9.3005
R6378 bgr_0.Vbe2.n55 bgr_0.Vbe2.n54 9.3005
R6379 bgr_0.Vbe2.n55 bgr_0.Vbe2.n35 9.3005
R6380 bgr_0.Vbe2.n55 bgr_0.Vbe2.n36 9.3005
R6381 bgr_0.Vbe2.n54 bgr_0.Vbe2.n52 9.3005
R6382 bgr_0.Vbe2.n52 bgr_0.Vbe2.n35 9.3005
R6383 bgr_0.Vbe2.n52 bgr_0.Vbe2.n37 9.3005
R6384 bgr_0.Vbe2.n52 bgr_0.Vbe2.n36 9.3005
R6385 bgr_0.Vbe2.n54 bgr_0.Vbe2.n3 9.3005
R6386 bgr_0.Vbe2.n38 bgr_0.Vbe2.n3 9.3005
R6387 bgr_0.Vbe2.n35 bgr_0.Vbe2.n3 9.3005
R6388 bgr_0.Vbe2.n37 bgr_0.Vbe2.n3 9.3005
R6389 bgr_0.Vbe2.n36 bgr_0.Vbe2.n3 9.3005
R6390 bgr_0.Vbe2.n39 bgr_0.Vbe2.n36 9.3005
R6391 bgr_0.Vbe2.n39 bgr_0.Vbe2.n37 9.3005
R6392 bgr_0.Vbe2.n39 bgr_0.Vbe2.n35 9.3005
R6393 bgr_0.Vbe2.n39 bgr_0.Vbe2.n38 9.3005
R6394 bgr_0.Vbe2.n57 bgr_0.Vbe2.n36 9.3005
R6395 bgr_0.Vbe2.n57 bgr_0.Vbe2.n37 9.3005
R6396 bgr_0.Vbe2.n57 bgr_0.Vbe2.n35 9.3005
R6397 bgr_0.Vbe2.n57 bgr_0.Vbe2.n38 9.3005
R6398 bgr_0.Vbe2.n57 bgr_0.Vbe2.n56 9.3005
R6399 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 9.3005
R6400 bgr_0.Vbe2.n53 bgr_0.Vbe2.n38 9.3005
R6401 bgr_0.Vbe2.n53 bgr_0.Vbe2.n35 9.3005
R6402 bgr_0.Vbe2.n53 bgr_0.Vbe2.n36 9.3005
R6403 bgr_0.Vbe2.n105 bgr_0.Vbe2.n15 4.64654
R6404 bgr_0.Vbe2.n92 bgr_0.Vbe2.n16 4.64654
R6405 bgr_0.Vbe2.n103 bgr_0.Vbe2.n14 4.64654
R6406 bgr_0.Vbe2.n94 bgr_0.Vbe2.n17 4.64654
R6407 bgr_0.Vbe2.n104 bgr_0.Vbe2.n103 4.64654
R6408 bgr_0.Vbe2.n43 bgr_0.Vbe2.n37 4.64654
R6409 bgr_0.Vbe2.n44 bgr_0.Vbe2.n38 4.64654
R6410 bgr_0.Vbe2.n56 bgr_0.Vbe2.n41 4.64654
R6411 bgr_0.Vbe2.n54 bgr_0.Vbe2.n34 4.64654
R6412 bgr_0.Vbe2.n56 bgr_0.Vbe2.n40 4.64654
R6413 bgr_0.Vbe2.n133 bgr_0.Vbe2.n132 2.36206
R6414 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 2.36206
R6415 bgr_0.Vbe2.n68 bgr_0.Vbe2.n29 2.36206
R6416 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 2.36206
R6417 bgr_0.Vbe2.n145 bgr_0.Vbe2.n144 2.19742
R6418 bgr_0.Vbe2.n131 bgr_0.Vbe2.n130 2.19742
R6419 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 2.19742
R6420 bgr_0.Vbe2.n71 bgr_0.Vbe2.n69 2.19742
R6421 bgr_0.Vbe2.n84 bgr_0.Vbe2.n82 2.19742
R6422 bgr_0.Vbe2.n110 bgr_0.Vbe2.n13 1.56363
R6423 bgr_0.Vbe2.n22 bgr_0.Vbe2.n20 1.56363
R6424 bgr_0.Vbe2.n83 bgr_0.Vbe2.n21 1.5505
R6425 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 1.5505
R6426 bgr_0.Vbe2.n70 bgr_0.Vbe2.n27 1.5505
R6427 bgr_0.Vbe2.n75 bgr_0.Vbe2.n74 1.5505
R6428 bgr_0.Vbe2.n77 bgr_0.Vbe2.n76 1.5505
R6429 bgr_0.Vbe2.n79 bgr_0.Vbe2.n24 1.5505
R6430 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 1.5505
R6431 bgr_0.Vbe2.n67 bgr_0.Vbe2.n66 1.5505
R6432 bgr_0.Vbe2.n31 bgr_0.Vbe2.n30 1.5505
R6433 bgr_0.Vbe2.n115 bgr_0.Vbe2.n11 1.5505
R6434 bgr_0.Vbe2.n113 bgr_0.Vbe2.n112 1.5505
R6435 bgr_0.Vbe2.n129 bgr_0.Vbe2.n6 1.5505
R6436 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 1.5505
R6437 bgr_0.Vbe2.n124 bgr_0.Vbe2.n123 1.5505
R6438 bgr_0.Vbe2.n10 bgr_0.Vbe2.n9 1.5505
R6439 bgr_0.Vbe2.n143 bgr_0.Vbe2.n0 1.5505
R6440 bgr_0.Vbe2.n141 bgr_0.Vbe2.n140 1.5505
R6441 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 1.5505
R6442 bgr_0.Vbe2.n5 bgr_0.Vbe2.n4 1.5505
R6443 bgr_0.Vbe2.n136 bgr_0.Vbe2.n5 1.25468
R6444 bgr_0.Vbe2.n122 bgr_0.Vbe2.n10 1.25468
R6445 bgr_0.Vbe2.n46 bgr_0.Vbe2.n37 1.25468
R6446 bgr_0.Vbe2.n66 bgr_0.Vbe2.n65 1.25468
R6447 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 1.25468
R6448 bgr_0.Vbe2.n96 bgr_0.Vbe2.n15 1.25468
R6449 bgr_0.Vbe2.n144 bgr_0.Vbe2.n143 1.19225
R6450 bgr_0.Vbe2.n130 bgr_0.Vbe2.n129 1.19225
R6451 bgr_0.Vbe2.n116 bgr_0.Vbe2.n115 1.19225
R6452 bgr_0.Vbe2.n54 bgr_0.Vbe2.n42 1.19225
R6453 bgr_0.Vbe2.n71 bgr_0.Vbe2.n70 1.19225
R6454 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 1.19225
R6455 bgr_0.Vbe2.n102 bgr_0.Vbe2.n17 1.19225
R6456 bgr_0.Vbe2.n137 bgr_0.Vbe2.n2 1.07024
R6457 bgr_0.Vbe2.n123 bgr_0.Vbe2.n8 1.07024
R6458 bgr_0.Vbe2.n48 bgr_0.Vbe2.n35 1.07024
R6459 bgr_0.Vbe2.n62 bgr_0.Vbe2.n31 1.07024
R6460 bgr_0.Vbe2.n77 bgr_0.Vbe2.n26 1.07024
R6461 bgr_0.Vbe2.n98 bgr_0.Vbe2.n18 1.07024
R6462 bgr_0.Vbe2.n133 bgr_0.Vbe2.n5 1.0237
R6463 bgr_0.Vbe2.n119 bgr_0.Vbe2.n10 1.0237
R6464 bgr_0.Vbe2.n45 bgr_0.Vbe2.n37 1.0237
R6465 bgr_0.Vbe2.n66 bgr_0.Vbe2.n29 1.0237
R6466 bgr_0.Vbe2.n80 bgr_0.Vbe2.n79 1.0237
R6467 bgr_0.Vbe2.n19 bgr_0.Vbe2.n15 1.0237
R6468 bgr_0.Vbe2.n142 bgr_0.Vbe2.n141 0.885803
R6469 bgr_0.Vbe2.n128 bgr_0.Vbe2.n127 0.885803
R6470 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 0.885803
R6471 bgr_0.Vbe2.n51 bgr_0.Vbe2.n38 0.885803
R6472 bgr_0.Vbe2.n61 bgr_0.Vbe2.n33 0.885803
R6473 bgr_0.Vbe2.n74 bgr_0.Vbe2.n73 0.885803
R6474 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 0.885803
R6475 bgr_0.Vbe2.n100 bgr_0.Vbe2.n16 0.885803
R6476 bgr_0.Vbe2.n45 bgr_0.Vbe2.n36 0.812055
R6477 bgr_0.Vbe2.n107 bgr_0.Vbe2.n19 0.812055
R6478 bgr_0.Vbe2.n141 bgr_0.Vbe2.n2 0.77514
R6479 bgr_0.Vbe2.n127 bgr_0.Vbe2.n8 0.77514
R6480 bgr_0.Vbe2.n113 bgr_0.Vbe2.n13 0.77514
R6481 bgr_0.Vbe2.n48 bgr_0.Vbe2.n38 0.77514
R6482 bgr_0.Vbe2.n62 bgr_0.Vbe2.n61 0.77514
R6483 bgr_0.Vbe2.n74 bgr_0.Vbe2.n26 0.77514
R6484 bgr_0.Vbe2.n87 bgr_0.Vbe2.n22 0.77514
R6485 bgr_0.Vbe2.n98 bgr_0.Vbe2.n16 0.77514
R6486 bgr_0.Vbe2 bgr_0.Vbe2.n142 0.756696
R6487 bgr_0.Vbe2 bgr_0.Vbe2.n128 0.756696
R6488 bgr_0.Vbe2 bgr_0.Vbe2.n114 0.756696
R6489 bgr_0.Vbe2 bgr_0.Vbe2.n51 0.756696
R6490 bgr_0.Vbe2 bgr_0.Vbe2.n33 0.756696
R6491 bgr_0.Vbe2.n73 bgr_0.Vbe2 0.756696
R6492 bgr_0.Vbe2.n86 bgr_0.Vbe2 0.756696
R6493 bgr_0.Vbe2.n100 bgr_0.Vbe2 0.756696
R6494 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 0.711459
R6495 bgr_0.Vbe2.n56 bgr_0.Vbe2.n42 0.647417
R6496 bgr_0.Vbe2.n103 bgr_0.Vbe2.n102 0.647417
R6497 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 0.590702
R6498 bgr_0.Vbe2.n123 bgr_0.Vbe2.n122 0.590702
R6499 bgr_0.Vbe2.n46 bgr_0.Vbe2.n35 0.590702
R6500 bgr_0.Vbe2.n65 bgr_0.Vbe2.n31 0.590702
R6501 bgr_0.Vbe2.n78 bgr_0.Vbe2.n77 0.590702
R6502 bgr_0.Vbe2.n96 bgr_0.Vbe2.n18 0.590702
R6503 bgr_0.Vbe2.n59 bgr_0.Vbe2 0.576566
R6504 bgr_0.Vbe2.n89 bgr_0.Vbe2.n20 0.530034
R6505 bgr_0.Vbe2.n111 bgr_0.Vbe2.n110 0.530034
R6506 bgr_0.Vbe2.t1 bgr_0.Vbe2.n134 0.290206
R6507 bgr_0.Vbe2.t8 bgr_0.Vbe2.n120 0.290206
R6508 bgr_0.Vbe2.t5 bgr_0.Vbe2.n109 0.290206
R6509 bgr_0.Vbe2.n49 bgr_0.Vbe2.t3 0.290206
R6510 bgr_0.Vbe2.t4 bgr_0.Vbe2.n63 0.290206
R6511 bgr_0.Vbe2.n28 bgr_0.Vbe2.t2 0.290206
R6512 bgr_0.Vbe2.n23 bgr_0.Vbe2.t7 0.290206
R6513 bgr_0.Vbe2.n99 bgr_0.Vbe2.t6 0.290206
R6514 bgr_0.Vbe2.n143 bgr_0.Vbe2 0.203382
R6515 bgr_0.Vbe2.n129 bgr_0.Vbe2 0.203382
R6516 bgr_0.Vbe2.n115 bgr_0.Vbe2 0.203382
R6517 bgr_0.Vbe2.n54 bgr_0.Vbe2 0.203382
R6518 bgr_0.Vbe2.n70 bgr_0.Vbe2 0.203382
R6519 bgr_0.Vbe2.n83 bgr_0.Vbe2 0.203382
R6520 bgr_0.Vbe2 bgr_0.Vbe2.n17 0.203382
R6521 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 0.154071
R6522 bgr_0.Vbe2.n69 bgr_0.Vbe2.n68 0.154071
R6523 bgr_0.Vbe2.n118 bgr_0.Vbe2.n117 0.154071
R6524 bgr_0.Vbe2.n132 bgr_0.Vbe2.n131 0.154071
R6525 bgr_0.Vbe2.n111 bgr_0.Vbe2.n108 0.137464
R6526 bgr_0.Vbe2.n139 bgr_0.Vbe2.n3 0.137464
R6527 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 0.134964
R6528 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 0.134964
R6529 bgr_0.Vbe2 bgr_0.Vbe2.n145 0.0196071
R6530 bgr_0.Vbe2.n88 bgr_0.Vbe2.n21 0.0183571
R6531 bgr_0.Vbe2.n82 bgr_0.Vbe2.n21 0.0183571
R6532 bgr_0.Vbe2.n81 bgr_0.Vbe2.n24 0.0183571
R6533 bgr_0.Vbe2.n76 bgr_0.Vbe2.n24 0.0183571
R6534 bgr_0.Vbe2.n76 bgr_0.Vbe2.n75 0.0183571
R6535 bgr_0.Vbe2.n75 bgr_0.Vbe2.n27 0.0183571
R6536 bgr_0.Vbe2.n69 bgr_0.Vbe2.n27 0.0183571
R6537 bgr_0.Vbe2.n68 bgr_0.Vbe2.n67 0.0183571
R6538 bgr_0.Vbe2.n67 bgr_0.Vbe2.n30 0.0183571
R6539 bgr_0.Vbe2.n112 bgr_0.Vbe2.n11 0.0183571
R6540 bgr_0.Vbe2.n117 bgr_0.Vbe2.n11 0.0183571
R6541 bgr_0.Vbe2.n118 bgr_0.Vbe2.n9 0.0183571
R6542 bgr_0.Vbe2.n124 bgr_0.Vbe2.n9 0.0183571
R6543 bgr_0.Vbe2.n126 bgr_0.Vbe2.n6 0.0183571
R6544 bgr_0.Vbe2.n131 bgr_0.Vbe2.n6 0.0183571
R6545 bgr_0.Vbe2.n132 bgr_0.Vbe2.n4 0.0183571
R6546 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 0.0183571
R6547 bgr_0.Vbe2.n140 bgr_0.Vbe2.n0 0.0183571
R6548 bgr_0.Vbe2.n145 bgr_0.Vbe2.n0 0.0183571
R6549 bgr_0.Vbe2.n58 bgr_0.Vbe2.n30 0.0106786
R6550 bgr_0.Vbe2.n139 bgr_0.Vbe2.n138 0.0106786
R6551 bgr_0.Vbe2.n126 bgr_0.Vbe2.n125 0.00996429
R6552 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.00992001
R6553 bgr_0.Vbe2.n106 bgr_0.Vbe2.n104 0.00992001
R6554 bgr_0.Vbe2.n105 bgr_0.Vbe2.n91 0.00992001
R6555 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 0.00992001
R6556 bgr_0.Vbe2.n108 bgr_0.Vbe2.n14 0.00992001
R6557 bgr_0.Vbe2.n92 bgr_0.Vbe2.n91 0.00992001
R6558 bgr_0.Vbe2.n93 bgr_0.Vbe2.n14 0.00992001
R6559 bgr_0.Vbe2.n104 bgr_0.Vbe2.n95 0.00992001
R6560 bgr_0.Vbe2.n94 bgr_0.Vbe2.n90 0.00992001
R6561 bgr_0.Vbe2.n106 bgr_0.Vbe2.n105 0.00992001
R6562 bgr_0.Vbe2.n39 bgr_0.Vbe2.n34 0.00992001
R6563 bgr_0.Vbe2.n53 bgr_0.Vbe2.n40 0.00992001
R6564 bgr_0.Vbe2.n55 bgr_0.Vbe2.n43 0.00992001
R6565 bgr_0.Vbe2.n52 bgr_0.Vbe2.n44 0.00992001
R6566 bgr_0.Vbe2.n41 bgr_0.Vbe2.n3 0.00992001
R6567 bgr_0.Vbe2.n55 bgr_0.Vbe2.n44 0.00992001
R6568 bgr_0.Vbe2.n52 bgr_0.Vbe2.n41 0.00992001
R6569 bgr_0.Vbe2.n40 bgr_0.Vbe2.n39 0.00992001
R6570 bgr_0.Vbe2.n57 bgr_0.Vbe2.n34 0.00992001
R6571 bgr_0.Vbe2.n53 bgr_0.Vbe2.n43 0.00992001
R6572 bgr_0.Vbe2.n125 bgr_0.Vbe2.n124 0.00889286
R6573 bgr_0.Vbe2.n89 bgr_0.Vbe2.n88 0.00817857
R6574 bgr_0.Vbe2.n60 bgr_0.Vbe2.n58 0.00817857
R6575 bgr_0.Vbe2.n112 bgr_0.Vbe2.n111 0.00817857
R6576 bgr_0.Vbe2.n140 bgr_0.Vbe2.n139 0.00817857
R6577 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t32 1172.87
R6578 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t40 1172.87
R6579 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t50 996.134
R6580 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t39 996.134
R6581 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t53 996.134
R6582 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t42 996.134
R6583 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t26 996.134
R6584 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t34 996.134
R6585 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R6586 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t36 996.134
R6587 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t52 851.534
R6588 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t29 851.534
R6589 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t28 674.801
R6590 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t44 674.801
R6591 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t27 674.801
R6592 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t43 674.801
R6593 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t54 674.801
R6594 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t47 674.801
R6595 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t33 674.801
R6596 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 674.801
R6597 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t30 530.201
R6598 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t38 530.201
R6599 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R6600 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t25 353.467
R6601 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t31 353.467
R6602 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t46 353.467
R6603 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t35 353.467
R6604 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t49 353.467
R6605 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t37 353.467
R6606 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t51 353.467
R6607 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n28 176.733
R6608 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R6609 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R6610 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6611 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6612 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6613 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 176.733
R6614 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R6615 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R6616 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R6617 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R6618 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R6619 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 176.733
R6620 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R6621 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R6622 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R6623 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R6624 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R6625 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n51 166.175
R6626 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.639
R6627 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.577
R6628 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n11 155.91
R6629 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 155.535
R6630 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 155.535
R6631 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 155.535
R6632 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n12 155.535
R6633 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 151.035
R6634 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n8 110.156
R6635 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n1 110.156
R6636 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n6 109.812
R6637 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n4 109.812
R6638 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n2 109.812
R6639 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n0 105.312
R6640 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R6641 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n22 51.9494
R6642 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R6643 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n31 51.9494
R6644 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 51.9494
R6645 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R6646 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.Y.n52 47.4599
R6647 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R6648 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R6649 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t0 16.0005
R6650 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t21 16.0005
R6651 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t23 16.0005
R6652 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R6653 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t16 16.0005
R6654 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t7 16.0005
R6655 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R6656 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t8 16.0005
R6657 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t20 16.0005
R6658 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t13 16.0005
R6659 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n21 13.4224
R6660 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 11.5786
R6661 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t12 11.2576
R6662 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t17 11.2576
R6663 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t2 11.2576
R6664 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t4 11.2576
R6665 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t24 11.2576
R6666 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t14 11.2576
R6667 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t18 11.2576
R6668 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t3 11.2576
R6669 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t22 11.2576
R6670 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t19 11.2576
R6671 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t5 11.2576
R6672 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t11 11.2576
R6673 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n10 6.96925
R6674 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n19 4.8755
R6675 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 4.5005
R6676 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 4.5005
R6677 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n42 1.73488
R6678 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n13 0.3755
R6679 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n15 0.3755
R6680 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n17 0.3755
R6681 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n3 0.34425
R6682 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n5 0.34425
R6683 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n7 0.34425
R6684 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.045
R6685 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 344.7
R6686 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R6687 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 201.565
R6688 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 201.222
R6689 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 201.222
R6690 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 201.222
R6691 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 201.222
R6692 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 120.16
R6693 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 39.4005
R6694 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R6695 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 39.4005
R6696 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 39.4005
R6697 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R6698 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 39.4005
R6699 two_stage_opamp_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 35.3599
R6700 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R6701 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R6702 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R6703 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 19.7005
R6704 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R6705 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 19.7005
R6706 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 19.7005
R6707 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R6708 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R6709 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 19.7005
R6710 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 5.46925
R6711 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 3.15675
R6712 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 0.34425
R6713 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 0.34425
R6714 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 0.34425
R6715 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.34425
R6716 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3 0.188
R6717 two_stage_opamp_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 0.063
R6718 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t1 384.967
R6719 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t5 369.534
R6720 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t20 369.534
R6721 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t23 369.534
R6722 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t15 369.534
R6723 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t17 369.534
R6724 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.n18 369.534
R6725 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 365.491
R6726 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t12 192.8
R6727 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t11 192.8
R6728 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t19 192.8
R6729 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t6 192.8
R6730 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t14 192.8
R6731 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t13 192.8
R6732 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t21 192.8
R6733 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t7 192.8
R6734 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t16 192.8
R6735 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t22 192.8
R6736 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t9 192.8
R6737 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t10 192.8
R6738 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t18 192.8
R6739 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t8 192.8
R6740 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R6741 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R6742 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R6743 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R6744 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R6745 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R6746 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R6747 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R6748 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R6749 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R6750 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R6751 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R6752 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R6753 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R6754 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R6755 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R6756 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R6757 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R6758 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t3 39.4005
R6759 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t0 39.4005
R6760 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 28.6755
R6761 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t4 24.0005
R6762 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t2 24.0005
R6763 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6764 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 514.134
R6765 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 323.142
R6766 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 322.692
R6767 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6768 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6769 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 270.591
R6770 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 270.591
R6771 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 233.374
R6772 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 233.374
R6773 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 233.374
R6774 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 233.374
R6775 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 208.838
R6776 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 197.964
R6777 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 174.726
R6778 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 174.726
R6779 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 174.726
R6780 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6781 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 169.216
R6782 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 169.216
R6783 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 169.216
R6784 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 129.24
R6785 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 129.24
R6786 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6787 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6788 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 128.534
R6789 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 128.534
R6790 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 16.8443
R6791 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6792 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6793 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6794 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6795 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6796 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6797 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 4.3755
R6798 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 4.3755
R6799 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 1.89425
R6800 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 1.59425
R6801 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 1.0255
R6802 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 0.688
R6803 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 0.688
R6804 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 0.4505
R6805 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 632.186
R6806 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 625.9
R6807 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 625.9
R6808 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 625.9
R6809 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 623.126
R6810 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 623.126
R6811 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 622.439
R6812 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 622.439
R6813 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 621.38
R6814 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 617.914
R6815 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6816 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6817 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6818 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6819 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6820 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6821 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6822 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6823 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6824 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6825 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6826 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6827 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6828 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6829 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6830 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6831 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6832 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6833 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 78.8005
R6834 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6835 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 6.3775
R6836 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 6.188
R6837 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 630.221
R6838 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n3 626.742
R6839 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n2 622.986
R6840 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 622.455
R6841 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 622.455
R6842 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.n24 585
R6843 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6844 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6845 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.n21 176.733
R6846 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R6847 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6848 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6849 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6850 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6851 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6852 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6853 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6854 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6855 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6856 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6857 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6858 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6859 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6860 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6861 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n23 161.808
R6862 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 135.232
R6863 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6864 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6865 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6866 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6867 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6868 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6869 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6870 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6871 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6872 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6873 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6874 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6875 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6876 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6877 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6878 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6879 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6880 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6881 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n1 82.5474
R6882 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6883 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6884 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6885 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6886 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6887 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6888 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6889 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6890 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6891 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R6892 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6893 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6894 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 49.8072
R6895 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n20 49.8072
R6896 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n25 41.7422
R6897 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate 35.4265
R6898 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t6 24.0005
R6899 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t5 24.0005
R6900 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 2.313
R6901 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R6902 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R6903 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R6904 bgr_0.V_mir2.n16 bgr_0.V_mir2.t22 310.488
R6905 bgr_0.V_mir2.n9 bgr_0.V_mir2.t17 310.488
R6906 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R6907 bgr_0.V_mir2.n2 bgr_0.V_mir2.t4 278.312
R6908 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R6909 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R6910 bgr_0.V_mir2.n18 bgr_0.V_mir2.t11 184.097
R6911 bgr_0.V_mir2.n11 bgr_0.V_mir2.t7 184.097
R6912 bgr_0.V_mir2.n6 bgr_0.V_mir2.t9 184.097
R6913 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R6914 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R6915 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R6916 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R6917 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R6918 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R6919 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R6920 bgr_0.V_mir2.n17 bgr_0.V_mir2.t13 120.501
R6921 bgr_0.V_mir2.n9 bgr_0.V_mir2.t21 120.501
R6922 bgr_0.V_mir2.n10 bgr_0.V_mir2.t15 120.501
R6923 bgr_0.V_mir2.n4 bgr_0.V_mir2.t18 120.501
R6924 bgr_0.V_mir2.n5 bgr_0.V_mir2.t5 120.501
R6925 bgr_0.V_mir2.n1 bgr_0.V_mir2.t3 48.0005
R6926 bgr_0.V_mir2.n1 bgr_0.V_mir2.t2 48.0005
R6927 bgr_0.V_mir2.n0 bgr_0.V_mir2.t1 48.0005
R6928 bgr_0.V_mir2.n0 bgr_0.V_mir2.t0 48.0005
R6929 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R6930 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R6931 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R6932 bgr_0.V_mir2.n12 bgr_0.V_mir2.t16 39.4005
R6933 bgr_0.V_mir2.n12 bgr_0.V_mir2.t8 39.4005
R6934 bgr_0.V_mir2.n7 bgr_0.V_mir2.t6 39.4005
R6935 bgr_0.V_mir2.n7 bgr_0.V_mir2.t10 39.4005
R6936 bgr_0.V_mir2.t14 bgr_0.V_mir2.n20 39.4005
R6937 bgr_0.V_mir2.n20 bgr_0.V_mir2.t12 39.4005
R6938 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R6939 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R6940 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R6941 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R6942 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R6943 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R6944 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t13 672.831
R6945 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 613.801
R6946 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t28 611.739
R6947 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t17 611.739
R6948 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R6949 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t31 611.739
R6950 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R6951 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R6952 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t16 421.75
R6953 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R6954 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R6955 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t12 421.75
R6956 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R6957 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t24 421.75
R6958 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t27 421.75
R6959 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R6960 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R6961 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t18 421.75
R6962 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R6963 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R6964 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R6965 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R6966 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t0 284.55
R6967 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n10 167.675
R6968 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 167.488
R6969 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R6970 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R6971 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R6972 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R6973 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R6974 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R6975 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R6976 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R6977 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R6978 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R6979 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.n3 167.094
R6980 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R6981 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n24 139.639
R6982 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n25 139.638
R6983 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n26 139.077
R6984 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n23 134.577
R6985 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t8 65.6672
R6986 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t1 65.6672
R6987 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n22 64.7974
R6988 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n18 40.7027
R6989 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n14 40.7027
R6990 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 40.7027
R6991 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n5 40.7027
R6992 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R6993 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R6994 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R6995 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R6996 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t10 24.0005
R6997 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R6998 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R6999 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R7000 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n1 16.0505
R7001 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 11.0786
R7002 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 4.5005
R7003 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 2.23488
R7004 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 0.766125
R7005 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 0.563
R7006 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n4 4020
R7007 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n4 4020
R7008 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 4020
R7009 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n10 4020
R7010 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t31 660.109
R7011 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t34 660.109
R7012 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n14 422.401
R7013 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n3 422.401
R7014 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.VD4.n11 239.915
R7015 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t32 239.915
R7016 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n8 220.8
R7017 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n6 220.8
R7018 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n6 188.8
R7019 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n3 188.8
R7020 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n0 155.911
R7021 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n23 155.91
R7022 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 155.537
R7023 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n19 155.536
R7024 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n1 155.536
R7025 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 155.535
R7026 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 155.535
R7027 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n28 155.535
R7028 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 155.535
R7029 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 155.535
R7030 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t33 155.125
R7031 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t36 155.125
R7032 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 151.036
R7033 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.VD4.t35 98.2764
R7034 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.VD4.t11 98.2764
R7035 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t15 98.2764
R7036 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.VD4.t19 98.2764
R7037 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.VD4.t3 98.2764
R7038 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.t9 98.2764
R7039 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t13 98.2764
R7040 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.VD4.t17 98.2764
R7041 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.VD4.t21 98.2764
R7042 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.VD4.t5 98.2764
R7043 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n13 92.5005
R7044 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n9 92.5005
R7045 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R7046 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 92.5005
R7047 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n4 92.5005
R7048 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n4 92.5005
R7049 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.t7 49.1384
R7050 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.VD4.n12 49.1384
R7051 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 21.3338
R7052 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 21.3338
R7053 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R7054 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R7055 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t14 11.2576
R7056 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t18 11.2576
R7057 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t20 11.2576
R7058 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t4 11.2576
R7059 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t12 11.2576
R7060 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t16 11.2576
R7061 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t24 11.2576
R7062 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t30 11.2576
R7063 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t28 11.2576
R7064 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R7065 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R7066 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R7067 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t2 11.2576
R7068 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t26 11.2576
R7069 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R7070 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t37 11.2576
R7071 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R7072 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R7073 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.t22 11.2576
R7074 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R7075 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 9.488
R7076 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n33 6.53175
R7077 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n22 5.3755
R7078 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n17 4.5005
R7079 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n31 0.3755
R7080 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n29 0.3755
R7081 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n27 0.3755
R7082 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.3755
R7083 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n2 0.3755
R7084 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n18 0.3755
R7085 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n20 0.3755
R7086 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t29 1172.87
R7087 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t35 1172.87
R7088 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t52 996.134
R7089 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.t39 996.134
R7090 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t26 996.134
R7091 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.t43 996.134
R7092 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t25 996.134
R7093 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t42 996.134
R7094 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t50 996.134
R7095 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t37 996.134
R7096 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t49 851.534
R7097 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.t27 851.534
R7098 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t33 674.801
R7099 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t46 674.801
R7100 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t34 674.801
R7101 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t47 674.801
R7102 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t31 674.801
R7103 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t45 674.801
R7104 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.t30 674.801
R7105 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.t44 674.801
R7106 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t28 530.201
R7107 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t32 530.201
R7108 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t40 353.467
R7109 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t48 353.467
R7110 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t36 353.467
R7111 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t51 353.467
R7112 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t38 353.467
R7113 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t54 353.467
R7114 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t41 353.467
R7115 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 353.467
R7116 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 176.733
R7117 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R7118 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R7119 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R7120 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R7121 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R7122 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 176.733
R7123 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.n42 176.733
R7124 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R7125 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R7126 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R7127 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R7128 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n17 176.733
R7129 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 176.733
R7130 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.n15 176.733
R7131 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 176.733
R7132 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n13 176.733
R7133 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.n11 176.733
R7134 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 166.175
R7135 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n40 161.637
R7136 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 161.577
R7137 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n21 155.91
R7138 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 155.535
R7139 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 155.535
R7140 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 155.535
R7141 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 155.535
R7142 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 151.035
R7143 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 110.374
R7144 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n1 110.374
R7145 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 109.812
R7146 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 109.812
R7147 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 109.812
R7148 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n0 105.312
R7149 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R7150 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n38 51.9494
R7151 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R7152 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n47 51.9494
R7153 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 51.9494
R7154 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n12 51.9494
R7155 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t20 47.46
R7156 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R7157 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t2 16.0005
R7158 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R7159 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t16 16.0005
R7160 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t1 16.0005
R7161 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t18 16.0005
R7162 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t24 16.0005
R7163 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R7164 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R7165 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t22 16.0005
R7166 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R7167 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t23 16.0005
R7168 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n31 13.4067
R7169 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 11.5943
R7170 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t19 11.2576
R7171 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R7172 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t12 11.2576
R7173 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R7174 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t9 11.2576
R7175 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R7176 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R7177 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t4 11.2576
R7178 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t8 11.2576
R7179 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t13 11.2576
R7180 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t10 11.2576
R7181 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t11 11.2576
R7182 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.X.n52 6.07862
R7183 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n29 4.8755
R7184 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 4.5005
R7185 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 4.5005
R7186 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n20 1.7505
R7187 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.X.n10 0.8755
R7188 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.563
R7189 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.563
R7190 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n8 0.563
R7191 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n27 0.3755
R7192 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n25 0.3755
R7193 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n23 0.3755
R7194 VOUT+.n2 VOUT+.n0 141.504
R7195 VOUT+.n8 VOUT+.n7 141.504
R7196 VOUT+.n6 VOUT+.n5 141.161
R7197 VOUT+.n4 VOUT+.n3 141.161
R7198 VOUT+.n2 VOUT+.n1 141.161
R7199 VOUT+.n10 VOUT+.n9 136.661
R7200 VOUT+.n96 VOUT+.t14 113.129
R7201 VOUT+.n93 VOUT+.n91 90.9636
R7202 VOUT+.n93 VOUT+.n92 90.3386
R7203 VOUT+.n95 VOUT+.n94 90.3386
R7204 VOUT+.n90 VOUT+.n10 15.0943
R7205 VOUT+.n90 VOUT+.n89 11.6871
R7206 VOUT+.n9 VOUT+.t11 6.56717
R7207 VOUT+.n9 VOUT+.t5 6.56717
R7208 VOUT+.n7 VOUT+.t9 6.56717
R7209 VOUT+.n7 VOUT+.t16 6.56717
R7210 VOUT+.n5 VOUT+.t10 6.56717
R7211 VOUT+.n5 VOUT+.t4 6.56717
R7212 VOUT+.n3 VOUT+.t2 6.56717
R7213 VOUT+.n3 VOUT+.t6 6.56717
R7214 VOUT+.n1 VOUT+.t3 6.56717
R7215 VOUT+.n1 VOUT+.t7 6.56717
R7216 VOUT+.n0 VOUT+.t15 6.56717
R7217 VOUT+.n0 VOUT+.t8 6.56717
R7218 VOUT+ VOUT+.n90 6.48488
R7219 VOUT+.n37 VOUT+.t108 4.8295
R7220 VOUT+.n46 VOUT+.t65 4.8295
R7221 VOUT+.n44 VOUT+.t118 4.8295
R7222 VOUT+.n42 VOUT+.t151 4.8295
R7223 VOUT+.n40 VOUT+.t44 4.8295
R7224 VOUT+.n39 VOUT+.t67 4.8295
R7225 VOUT+.n59 VOUT+.t27 4.8295
R7226 VOUT+.n60 VOUT+.t76 4.8295
R7227 VOUT+.n62 VOUT+.t62 4.8295
R7228 VOUT+.n63 VOUT+.t112 4.8295
R7229 VOUT+.n65 VOUT+.t114 4.8295
R7230 VOUT+.n66 VOUT+.t99 4.8295
R7231 VOUT+.n68 VOUT+.t74 4.8295
R7232 VOUT+.n69 VOUT+.t55 4.8295
R7233 VOUT+.n71 VOUT+.t109 4.8295
R7234 VOUT+.n72 VOUT+.t91 4.8295
R7235 VOUT+.n74 VOUT+.t68 4.8295
R7236 VOUT+.n75 VOUT+.t52 4.8295
R7237 VOUT+.n77 VOUT+.t29 4.8295
R7238 VOUT+.n78 VOUT+.t153 4.8295
R7239 VOUT+.n80 VOUT+.t63 4.8295
R7240 VOUT+.n81 VOUT+.t46 4.8295
R7241 VOUT+.n83 VOUT+.t22 4.8295
R7242 VOUT+.n84 VOUT+.t146 4.8295
R7243 VOUT+.n11 VOUT+.t117 4.8295
R7244 VOUT+.n13 VOUT+.t72 4.8295
R7245 VOUT+.n25 VOUT+.t37 4.8295
R7246 VOUT+.n26 VOUT+.t20 4.8295
R7247 VOUT+.n28 VOUT+.t79 4.8295
R7248 VOUT+.n29 VOUT+.t60 4.8295
R7249 VOUT+.n31 VOUT+.t121 4.8295
R7250 VOUT+.n32 VOUT+.t104 4.8295
R7251 VOUT+.n34 VOUT+.t84 4.8295
R7252 VOUT+.n35 VOUT+.t66 4.8295
R7253 VOUT+.n86 VOUT+.t123 4.8295
R7254 VOUT+.n48 VOUT+.t95 4.8154
R7255 VOUT+.n49 VOUT+.t70 4.8154
R7256 VOUT+.n50 VOUT+.t110 4.8154
R7257 VOUT+.n51 VOUT+.t145 4.8154
R7258 VOUT+.n48 VOUT+.t32 4.806
R7259 VOUT+.n49 VOUT+.t150 4.806
R7260 VOUT+.n50 VOUT+.t50 4.806
R7261 VOUT+.n51 VOUT+.t87 4.806
R7262 VOUT+.n52 VOUT+.t125 4.806
R7263 VOUT+.n53 VOUT+.t105 4.806
R7264 VOUT+.n54 VOUT+.t140 4.806
R7265 VOUT+.n55 VOUT+.t36 4.806
R7266 VOUT+.n56 VOUT+.t156 4.806
R7267 VOUT+.n57 VOUT+.t53 4.806
R7268 VOUT+.n14 VOUT+.t73 4.806
R7269 VOUT+.n15 VOUT+.t116 4.806
R7270 VOUT+.n16 VOUT+.t64 4.806
R7271 VOUT+.n17 VOUT+.t154 4.806
R7272 VOUT+.n18 VOUT+.t106 4.806
R7273 VOUT+.n19 VOUT+.t143 4.806
R7274 VOUT+.n20 VOUT+.t96 4.806
R7275 VOUT+.n21 VOUT+.t42 4.806
R7276 VOUT+.n22 VOUT+.t86 4.806
R7277 VOUT+.n23 VOUT+.t34 4.806
R7278 VOUT+.n37 VOUT+.t69 4.5005
R7279 VOUT+.n38 VOUT+.t90 4.5005
R7280 VOUT+.n46 VOUT+.t80 4.5005
R7281 VOUT+.n47 VOUT+.t43 4.5005
R7282 VOUT+.n44 VOUT+.t56 4.5005
R7283 VOUT+.n45 VOUT+.t21 4.5005
R7284 VOUT+.n42 VOUT+.t98 4.5005
R7285 VOUT+.n43 VOUT+.t59 4.5005
R7286 VOUT+.n40 VOUT+.t136 4.5005
R7287 VOUT+.n41 VOUT+.t101 4.5005
R7288 VOUT+.n39 VOUT+.t30 4.5005
R7289 VOUT+.n58 VOUT+.t51 4.5005
R7290 VOUT+.n57 VOUT+.t155 4.5005
R7291 VOUT+.n56 VOUT+.t119 4.5005
R7292 VOUT+.n55 VOUT+.t139 4.5005
R7293 VOUT+.n54 VOUT+.t102 4.5005
R7294 VOUT+.n53 VOUT+.t61 4.5005
R7295 VOUT+.n52 VOUT+.t85 4.5005
R7296 VOUT+.n51 VOUT+.t45 4.5005
R7297 VOUT+.n50 VOUT+.t147 4.5005
R7298 VOUT+.n49 VOUT+.t111 4.5005
R7299 VOUT+.n48 VOUT+.t134 4.5005
R7300 VOUT+.n59 VOUT+.t130 4.5005
R7301 VOUT+.n61 VOUT+.t152 4.5005
R7302 VOUT+.n60 VOUT+.t115 4.5005
R7303 VOUT+.n62 VOUT+.t23 4.5005
R7304 VOUT+.n64 VOUT+.t47 4.5005
R7305 VOUT+.n63 VOUT+.t148 4.5005
R7306 VOUT+.n65 VOUT+.t78 4.5005
R7307 VOUT+.n67 VOUT+.t26 4.5005
R7308 VOUT+.n66 VOUT+.t132 4.5005
R7309 VOUT+.n68 VOUT+.t39 4.5005
R7310 VOUT+.n70 VOUT+.t128 4.5005
R7311 VOUT+.n69 VOUT+.t92 4.5005
R7312 VOUT+.n71 VOUT+.t71 4.5005
R7313 VOUT+.n73 VOUT+.t19 4.5005
R7314 VOUT+.n72 VOUT+.t126 4.5005
R7315 VOUT+.n74 VOUT+.t33 4.5005
R7316 VOUT+.n76 VOUT+.t122 4.5005
R7317 VOUT+.n75 VOUT+.t88 4.5005
R7318 VOUT+.n77 VOUT+.t135 4.5005
R7319 VOUT+.n79 VOUT+.t82 4.5005
R7320 VOUT+.n78 VOUT+.t48 4.5005
R7321 VOUT+.n80 VOUT+.t28 4.5005
R7322 VOUT+.n82 VOUT+.t120 4.5005
R7323 VOUT+.n81 VOUT+.t81 4.5005
R7324 VOUT+.n83 VOUT+.t129 4.5005
R7325 VOUT+.n85 VOUT+.t77 4.5005
R7326 VOUT+.n84 VOUT+.t40 4.5005
R7327 VOUT+.n11 VOUT+.t25 4.5005
R7328 VOUT+.n12 VOUT+.t124 4.5005
R7329 VOUT+.n13 VOUT+.t38 4.5005
R7330 VOUT+.n24 VOUT+.t127 4.5005
R7331 VOUT+.n23 VOUT+.t94 4.5005
R7332 VOUT+.n22 VOUT+.t54 4.5005
R7333 VOUT+.n21 VOUT+.t144 4.5005
R7334 VOUT+.n20 VOUT+.t113 4.5005
R7335 VOUT+.n19 VOUT+.t75 4.5005
R7336 VOUT+.n18 VOUT+.t24 4.5005
R7337 VOUT+.n17 VOUT+.t131 4.5005
R7338 VOUT+.n16 VOUT+.t97 4.5005
R7339 VOUT+.n15 VOUT+.t58 4.5005
R7340 VOUT+.n14 VOUT+.t149 4.5005
R7341 VOUT+.n25 VOUT+.t142 4.5005
R7342 VOUT+.n27 VOUT+.t93 4.5005
R7343 VOUT+.n26 VOUT+.t57 4.5005
R7344 VOUT+.n28 VOUT+.t41 4.5005
R7345 VOUT+.n30 VOUT+.t133 4.5005
R7346 VOUT+.n29 VOUT+.t100 4.5005
R7347 VOUT+.n31 VOUT+.t83 4.5005
R7348 VOUT+.n33 VOUT+.t31 4.5005
R7349 VOUT+.n32 VOUT+.t137 4.5005
R7350 VOUT+.n34 VOUT+.t49 4.5005
R7351 VOUT+.n36 VOUT+.t138 4.5005
R7352 VOUT+.n35 VOUT+.t103 4.5005
R7353 VOUT+.n86 VOUT+.t89 4.5005
R7354 VOUT+.n87 VOUT+.t35 4.5005
R7355 VOUT+.n88 VOUT+.t141 4.5005
R7356 VOUT+.n89 VOUT+.t107 4.5005
R7357 VOUT+.n10 VOUT+.n8 4.5005
R7358 VOUT+.n91 VOUT+.t1 3.42907
R7359 VOUT+.n91 VOUT+.t18 3.42907
R7360 VOUT+.n92 VOUT+.t12 3.42907
R7361 VOUT+.n92 VOUT+.t0 3.42907
R7362 VOUT+.n94 VOUT+.t17 3.42907
R7363 VOUT+.n94 VOUT+.t13 3.42907
R7364 VOUT+ VOUT+.n96 1.54738
R7365 VOUT+.n96 VOUT+.n95 1.07862
R7366 VOUT+.n95 VOUT+.n93 0.6255
R7367 VOUT+.n4 VOUT+.n2 0.34425
R7368 VOUT+.n6 VOUT+.n4 0.34425
R7369 VOUT+.n8 VOUT+.n6 0.34425
R7370 VOUT+.n38 VOUT+.n37 0.3295
R7371 VOUT+.n47 VOUT+.n46 0.3295
R7372 VOUT+.n45 VOUT+.n44 0.3295
R7373 VOUT+.n43 VOUT+.n42 0.3295
R7374 VOUT+.n41 VOUT+.n40 0.3295
R7375 VOUT+.n58 VOUT+.n39 0.3295
R7376 VOUT+.n58 VOUT+.n57 0.3295
R7377 VOUT+.n57 VOUT+.n56 0.3295
R7378 VOUT+.n56 VOUT+.n55 0.3295
R7379 VOUT+.n55 VOUT+.n54 0.3295
R7380 VOUT+.n54 VOUT+.n53 0.3295
R7381 VOUT+.n53 VOUT+.n52 0.3295
R7382 VOUT+.n52 VOUT+.n51 0.3295
R7383 VOUT+.n51 VOUT+.n50 0.3295
R7384 VOUT+.n50 VOUT+.n49 0.3295
R7385 VOUT+.n49 VOUT+.n48 0.3295
R7386 VOUT+.n61 VOUT+.n59 0.3295
R7387 VOUT+.n61 VOUT+.n60 0.3295
R7388 VOUT+.n64 VOUT+.n62 0.3295
R7389 VOUT+.n64 VOUT+.n63 0.3295
R7390 VOUT+.n67 VOUT+.n65 0.3295
R7391 VOUT+.n67 VOUT+.n66 0.3295
R7392 VOUT+.n70 VOUT+.n68 0.3295
R7393 VOUT+.n70 VOUT+.n69 0.3295
R7394 VOUT+.n73 VOUT+.n71 0.3295
R7395 VOUT+.n73 VOUT+.n72 0.3295
R7396 VOUT+.n76 VOUT+.n74 0.3295
R7397 VOUT+.n76 VOUT+.n75 0.3295
R7398 VOUT+.n79 VOUT+.n77 0.3295
R7399 VOUT+.n79 VOUT+.n78 0.3295
R7400 VOUT+.n82 VOUT+.n80 0.3295
R7401 VOUT+.n82 VOUT+.n81 0.3295
R7402 VOUT+.n85 VOUT+.n83 0.3295
R7403 VOUT+.n85 VOUT+.n84 0.3295
R7404 VOUT+.n12 VOUT+.n11 0.3295
R7405 VOUT+.n24 VOUT+.n13 0.3295
R7406 VOUT+.n24 VOUT+.n23 0.3295
R7407 VOUT+.n23 VOUT+.n22 0.3295
R7408 VOUT+.n22 VOUT+.n21 0.3295
R7409 VOUT+.n21 VOUT+.n20 0.3295
R7410 VOUT+.n20 VOUT+.n19 0.3295
R7411 VOUT+.n19 VOUT+.n18 0.3295
R7412 VOUT+.n18 VOUT+.n17 0.3295
R7413 VOUT+.n17 VOUT+.n16 0.3295
R7414 VOUT+.n16 VOUT+.n15 0.3295
R7415 VOUT+.n15 VOUT+.n14 0.3295
R7416 VOUT+.n27 VOUT+.n25 0.3295
R7417 VOUT+.n27 VOUT+.n26 0.3295
R7418 VOUT+.n30 VOUT+.n28 0.3295
R7419 VOUT+.n30 VOUT+.n29 0.3295
R7420 VOUT+.n33 VOUT+.n31 0.3295
R7421 VOUT+.n33 VOUT+.n32 0.3295
R7422 VOUT+.n36 VOUT+.n34 0.3295
R7423 VOUT+.n36 VOUT+.n35 0.3295
R7424 VOUT+.n87 VOUT+.n86 0.3295
R7425 VOUT+.n88 VOUT+.n87 0.3295
R7426 VOUT+.n89 VOUT+.n88 0.3295
R7427 VOUT+.n52 VOUT+.n47 0.306
R7428 VOUT+.n53 VOUT+.n45 0.306
R7429 VOUT+.n54 VOUT+.n43 0.306
R7430 VOUT+.n55 VOUT+.n41 0.306
R7431 VOUT+.n58 VOUT+.n38 0.2825
R7432 VOUT+.n61 VOUT+.n58 0.2825
R7433 VOUT+.n64 VOUT+.n61 0.2825
R7434 VOUT+.n67 VOUT+.n64 0.2825
R7435 VOUT+.n70 VOUT+.n67 0.2825
R7436 VOUT+.n73 VOUT+.n70 0.2825
R7437 VOUT+.n76 VOUT+.n73 0.2825
R7438 VOUT+.n79 VOUT+.n76 0.2825
R7439 VOUT+.n82 VOUT+.n79 0.2825
R7440 VOUT+.n85 VOUT+.n82 0.2825
R7441 VOUT+.n24 VOUT+.n12 0.2825
R7442 VOUT+.n27 VOUT+.n24 0.2825
R7443 VOUT+.n30 VOUT+.n27 0.2825
R7444 VOUT+.n33 VOUT+.n30 0.2825
R7445 VOUT+.n36 VOUT+.n33 0.2825
R7446 VOUT+.n87 VOUT+.n36 0.2825
R7447 VOUT+.n87 VOUT+.n85 0.2825
R7448 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t25 369.534
R7449 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t24 369.534
R7450 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t15 369.534
R7451 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t11 369.534
R7452 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t17 369.534
R7453 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t16 369.534
R7454 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7455 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7456 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7457 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7458 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t21 238.322
R7459 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t13 238.322
R7460 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t4 194.895
R7461 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t18 192.8
R7462 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t10 192.8
R7463 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t14 192.8
R7464 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t22 192.8
R7465 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t28 192.8
R7466 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t19 192.8
R7467 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t26 192.8
R7468 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t12 192.8
R7469 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t20 192.8
R7470 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t27 192.8
R7471 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t29 192.8
R7472 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t23 192.8
R7473 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7474 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7475 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7476 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7477 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7478 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7479 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7480 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 169.394
R7481 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7482 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7483 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t8 100.635
R7484 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7485 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7486 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7487 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7488 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7489 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7490 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t6 39.4005
R7491 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t2 39.4005
R7492 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t1 39.4005
R7493 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t3 39.4005
R7494 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t9 39.4005
R7495 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t5 39.4005
R7496 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t0 39.4005
R7497 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t7 39.4005
R7498 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 26.9067
R7499 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 5.15675
R7500 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7501 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n14 4.188
R7502 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 3.03175
R7503 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7504 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7505 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t20 449.868
R7506 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t25 449.868
R7507 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7508 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t21 449.868
R7509 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R7510 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R7511 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7512 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t18 273.134
R7513 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7514 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7515 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t13 273.134
R7516 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7517 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7518 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7519 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7520 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t16 273.134
R7521 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7522 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t14 273.134
R7523 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7524 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7525 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7526 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7527 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R7528 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R7529 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R7530 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 176.733
R7531 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R7532 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7533 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R7534 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R7535 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R7536 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R7537 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R7538 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7539 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t3 175.566
R7540 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n11 168.769
R7541 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 165.8
R7542 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t2 61.057
R7543 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 56.563
R7544 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 56.2338
R7545 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n15 56.2338
R7546 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 56.2338
R7547 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n6 56.2338
R7548 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7549 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7550 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7551 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t1 39.4005
R7552 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 11.5673
R7553 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n21 11.0786
R7554 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 2.26612
R7555 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 112.338
R7556 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.62
R7557 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.62
R7558 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 110.306
R7559 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 110.306
R7560 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 110.171
R7561 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 110.171
R7562 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n7 109.828
R7563 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 109.828
R7564 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.12
R7565 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 105.309
R7566 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7567 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7568 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7569 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7570 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7571 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7572 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7573 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7574 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7575 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7576 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7577 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7578 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7579 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7580 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7581 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7582 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7583 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7584 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7585 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7586 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7587 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7588 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7589 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7590 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 1.84425
R7591 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 0.71925
R7592 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 0.688
R7593 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 0.688
R7594 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n6 0.34425
R7595 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n8 0.34425
R7596 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.170955
R7597 a_5160_5068.t0 a_5160_5068.t1 422.339
R7598 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 144.827
R7599 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 134.577
R7600 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 119.198
R7601 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 91.2435
R7602 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 90.8997
R7603 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 90.8997
R7604 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 90.8997
R7605 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 90.8997
R7606 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 24.0005
R7607 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R7608 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R7609 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 24.0005
R7610 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 6.0005
R7611 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 6.0005
R7612 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 6.0005
R7613 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 6.0005
R7614 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 6.0005
R7615 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 6.0005
R7616 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 6.0005
R7617 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 6.0005
R7618 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 6.0005
R7619 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 6.0005
R7620 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 5.29738
R7621 two_stage_opamp_dummy_magic_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 0.766125
R7622 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 0.34425
R7623 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 0.34425
R7624 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.34425
R7625 two_stage_opamp_dummy_magic_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 0.063
R7626 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7627 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7628 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7629 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 310.488
R7630 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7631 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7632 bgr_0.V_mir1.n7 bgr_0.V_mir1.t15 278.312
R7633 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7634 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7635 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R7636 bgr_0.V_mir1.n11 bgr_0.V_mir1.t0 184.097
R7637 bgr_0.V_mir1.n2 bgr_0.V_mir1.t8 184.097
R7638 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7639 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7640 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7641 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7642 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7643 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7644 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 120.501
R7645 bgr_0.V_mir1.n17 bgr_0.V_mir1.t2 120.501
R7646 bgr_0.V_mir1.n9 bgr_0.V_mir1.t18 120.501
R7647 bgr_0.V_mir1.n10 bgr_0.V_mir1.t4 120.501
R7648 bgr_0.V_mir1.n0 bgr_0.V_mir1.t17 120.501
R7649 bgr_0.V_mir1.n1 bgr_0.V_mir1.t6 120.501
R7650 bgr_0.V_mir1.n6 bgr_0.V_mir1.t14 48.0005
R7651 bgr_0.V_mir1.n6 bgr_0.V_mir1.t16 48.0005
R7652 bgr_0.V_mir1.n5 bgr_0.V_mir1.t12 48.0005
R7653 bgr_0.V_mir1.n5 bgr_0.V_mir1.t13 48.0005
R7654 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7655 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7656 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7657 bgr_0.V_mir1.n12 bgr_0.V_mir1.t1 39.4005
R7658 bgr_0.V_mir1.n12 bgr_0.V_mir1.t5 39.4005
R7659 bgr_0.V_mir1.n3 bgr_0.V_mir1.t9 39.4005
R7660 bgr_0.V_mir1.n3 bgr_0.V_mir1.t7 39.4005
R7661 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7662 bgr_0.V_mir1.n20 bgr_0.V_mir1.t3 39.4005
R7663 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7664 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7665 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7666 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7667 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7668 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7669 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t5 49.8805
R7670 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.1603
R7671 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R7672 two_stage_opamp_dummy_magic_0.cap_res_X.t9 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.1603
R7673 two_stage_opamp_dummy_magic_0.cap_res_X.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.1603
R7674 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R7675 two_stage_opamp_dummy_magic_0.cap_res_X.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1603
R7676 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R7677 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.1603
R7678 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1603
R7679 two_stage_opamp_dummy_magic_0.cap_res_X.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.1603
R7680 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R7681 two_stage_opamp_dummy_magic_0.cap_res_X.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1603
R7682 two_stage_opamp_dummy_magic_0.cap_res_X.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.1603
R7683 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R7684 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1603
R7685 two_stage_opamp_dummy_magic_0.cap_res_X.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.1603
R7686 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1603
R7687 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1603
R7688 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.1603
R7689 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.1603
R7690 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1603
R7691 two_stage_opamp_dummy_magic_0.cap_res_X.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.1603
R7692 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.1603
R7693 two_stage_opamp_dummy_magic_0.cap_res_X.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R7694 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1603
R7695 two_stage_opamp_dummy_magic_0.cap_res_X.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1603
R7696 two_stage_opamp_dummy_magic_0.cap_res_X.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1603
R7697 two_stage_opamp_dummy_magic_0.cap_res_X.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R7698 two_stage_opamp_dummy_magic_0.cap_res_X.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1603
R7699 two_stage_opamp_dummy_magic_0.cap_res_X.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R7700 two_stage_opamp_dummy_magic_0.cap_res_X.t15 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1603
R7701 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.1603
R7702 two_stage_opamp_dummy_magic_0.cap_res_X.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R7703 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.1603
R7704 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.1603
R7705 two_stage_opamp_dummy_magic_0.cap_res_X.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1603
R7706 two_stage_opamp_dummy_magic_0.cap_res_X.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.1603
R7707 two_stage_opamp_dummy_magic_0.cap_res_X.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1603
R7708 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R7709 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1603
R7710 two_stage_opamp_dummy_magic_0.cap_res_X.t7 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R7711 two_stage_opamp_dummy_magic_0.cap_res_X.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1603
R7712 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1603
R7713 two_stage_opamp_dummy_magic_0.cap_res_X.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.1603
R7714 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R7715 two_stage_opamp_dummy_magic_0.cap_res_X.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R7716 two_stage_opamp_dummy_magic_0.cap_res_X.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.1603
R7717 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R7718 two_stage_opamp_dummy_magic_0.cap_res_X.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.1603
R7719 two_stage_opamp_dummy_magic_0.cap_res_X.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R7720 two_stage_opamp_dummy_magic_0.cap_res_X.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1603
R7721 two_stage_opamp_dummy_magic_0.cap_res_X.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1603
R7722 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.1603
R7723 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.1603
R7724 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.1603
R7725 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1603
R7726 two_stage_opamp_dummy_magic_0.cap_res_X.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R7727 two_stage_opamp_dummy_magic_0.cap_res_X.t5 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R7728 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.159278
R7729 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.159278
R7730 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.159278
R7731 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.159278
R7732 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.159278
R7733 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.159278
R7734 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.159278
R7735 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.159278
R7736 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.159278
R7737 two_stage_opamp_dummy_magic_0.cap_res_X.t23 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.159278
R7738 two_stage_opamp_dummy_magic_0.cap_res_X.t125 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.159278
R7739 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.159278
R7740 two_stage_opamp_dummy_magic_0.cap_res_X.t121 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.159278
R7741 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R7742 two_stage_opamp_dummy_magic_0.cap_res_X.t36 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R7743 two_stage_opamp_dummy_magic_0.cap_res_X.t74 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R7744 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R7745 two_stage_opamp_dummy_magic_0.cap_res_X.t137 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R7746 two_stage_opamp_dummy_magic_0.cap_res_X.t28 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R7747 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R7748 two_stage_opamp_dummy_magic_0.cap_res_X.t109 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R7749 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R7750 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R7751 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.159278
R7752 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t0 0.159278
R7753 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.159278
R7754 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.159278
R7755 two_stage_opamp_dummy_magic_0.cap_res_X.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.137822
R7756 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.1368
R7757 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.1368
R7758 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1368
R7759 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R7760 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1368
R7761 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R7762 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R7763 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.1368
R7764 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1368
R7765 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.1368
R7766 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1368
R7767 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R7768 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1368
R7769 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1368
R7770 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1368
R7771 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.1368
R7772 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1368
R7773 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1368
R7774 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1368
R7775 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1368
R7776 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.1368
R7777 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1368
R7778 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.1368
R7779 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1368
R7780 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1368
R7781 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.1368
R7782 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1368
R7783 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.1368
R7784 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1368
R7785 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1368
R7786 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1368
R7787 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.114322
R7788 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.1133
R7789 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.1133
R7790 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R7791 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R7792 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R7793 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R7794 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R7795 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R7796 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R7797 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R7798 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R7799 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R7800 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R7801 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R7802 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.1133
R7803 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.1133
R7804 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.1133
R7805 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.1133
R7806 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R7807 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.00152174
R7808 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.00152174
R7809 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.00152174
R7810 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.00152174
R7811 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.00152174
R7812 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.00152174
R7813 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.00152174
R7814 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.00152174
R7815 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.00152174
R7816 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R7817 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.00152174
R7818 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.00152174
R7819 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R7820 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.00152174
R7821 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.00152174
R7822 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.00152174
R7823 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R7824 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.00152174
R7825 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.00152174
R7826 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.00152174
R7827 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R7828 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.00152174
R7829 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.00152174
R7830 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.00152174
R7831 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.00152174
R7832 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.00152174
R7833 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.00152174
R7834 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.00152174
R7835 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R7836 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.00152174
R7837 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R7838 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.00152174
R7839 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R7840 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.00152174
R7841 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R7842 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R7843 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R7844 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 145.046
R7845 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 134.797
R7846 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 118.885
R7847 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 91.2435
R7848 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 90.8997
R7849 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 90.8997
R7850 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 90.8997
R7851 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 90.8997
R7852 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 24.0005
R7853 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R7854 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 24.0005
R7855 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 24.0005
R7856 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 6.0005
R7857 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 6.0005
R7858 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 6.0005
R7859 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 6.0005
R7860 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 6.0005
R7861 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 6.0005
R7862 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 6.0005
R7863 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 6.0005
R7864 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 6.0005
R7865 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 6.0005
R7866 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 5.29738
R7867 two_stage_opamp_dummy_magic_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 0.59425
R7868 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.34425
R7869 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 0.34425
R7870 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 0.34425
R7871 two_stage_opamp_dummy_magic_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 0.063
R7872 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 525.38
R7873 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 525.38
R7874 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 366.856
R7875 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 360.43
R7876 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7877 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 281.168
R7878 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 281.168
R7879 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 281.168
R7880 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7881 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7882 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 165.972
R7883 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 165.972
R7884 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 115.52
R7885 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 115.52
R7886 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7887 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 79.2627
R7888 two_stage_opamp_dummy_magic_0.V_b_2nd_stage two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 18.4432
R7889 two_stage_opamp_dummy_magic_0.V_b_2nd_stage two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 11.6047
R7890 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 229.562
R7891 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7892 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7893 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7894 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7895 bgr_0.V_p_2.n1 bgr_0.V_p_2.t10 98.2279
R7896 bgr_0.V_p_2.n5 bgr_0.V_p_2.t0 48.0005
R7897 bgr_0.V_p_2.n5 bgr_0.V_p_2.t7 48.0005
R7898 bgr_0.V_p_2.n4 bgr_0.V_p_2.t4 48.0005
R7899 bgr_0.V_p_2.n4 bgr_0.V_p_2.t3 48.0005
R7900 bgr_0.V_p_2.n3 bgr_0.V_p_2.t1 48.0005
R7901 bgr_0.V_p_2.n3 bgr_0.V_p_2.t6 48.0005
R7902 bgr_0.V_p_2.n2 bgr_0.V_p_2.t5 48.0005
R7903 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R7904 bgr_0.V_p_2.t8 bgr_0.V_p_2.n6 48.0005
R7905 bgr_0.V_p_2.n6 bgr_0.V_p_2.t9 48.0005
R7906 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7907 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7908 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7909 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7910 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7911 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7912 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 622.955
R7913 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 622.955
R7914 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 622.268
R7915 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 622.268
R7916 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 622.268
R7917 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 617.768
R7918 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7919 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7920 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7921 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7922 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7923 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7924 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7925 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7926 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7927 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7928 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7929 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7930 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7931 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7932 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7933 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7934 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7935 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7936 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7937 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7938 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7939 two_stage_opamp_dummy_magic_0.V_err_p.t14 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7940 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7941 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7942 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 0.764705
R7943 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 0.688
R7944 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 0.688
R7945 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 0.688
R7946 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7947 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7948 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R7949 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R7950 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R7951 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 201.565
R7952 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 201.222
R7953 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 201.222
R7954 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 201.222
R7955 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 201.222
R7956 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 120.16
R7957 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 71.2813
R7958 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R7959 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 47.2974
R7960 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 39.4005
R7961 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R7962 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R7963 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R7964 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R7965 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 39.4005
R7966 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R7967 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 19.7005
R7968 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R7969 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R7970 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R7971 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R7972 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R7973 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R7974 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R7975 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R7976 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 5.46925
R7977 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1 1.15675
R7978 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 0.34425
R7979 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 0.34425
R7980 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 0.34425
R7981 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 0.063
R7982 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7983 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7984 bgr_0.Vin+.n0 bgr_0.Vin+.t6 303.259
R7985 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R7986 bgr_0.Vin+.n0 bgr_0.Vin+.t8 174.726
R7987 bgr_0.Vin+.n1 bgr_0.Vin+.t10 174.726
R7988 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R7989 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R7990 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R7991 bgr_0.Vin+.t0 bgr_0.Vin+.n8 158.796
R7992 bgr_0.Vin+.n8 bgr_0.Vin+.t1 147.981
R7993 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7994 bgr_0.Vin+.n3 bgr_0.Vin+.t9 96.4005
R7995 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R7996 bgr_0.Vin+.n5 bgr_0.Vin+.t2 13.1338
R7997 bgr_0.Vin+.n5 bgr_0.Vin+.t5 13.1338
R7998 bgr_0.Vin+.n4 bgr_0.Vin+.t4 13.1338
R7999 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R8000 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R8001 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 229.562
R8002 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R8003 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R8004 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R8005 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R8006 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.2279
R8007 bgr_0.V_p_1.n5 bgr_0.V_p_1.t5 48.0005
R8008 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R8009 bgr_0.V_p_1.n4 bgr_0.V_p_1.t0 48.0005
R8010 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8011 bgr_0.V_p_1.n3 bgr_0.V_p_1.t6 48.0005
R8012 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R8013 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R8014 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R8015 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8016 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R8017 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R8018 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t13 355.293
R8019 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.t14 346.8
R8020 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.n20 339.522
R8021 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 339.522
R8022 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n14 335.022
R8023 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t4 275.909
R8024 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 227.909
R8025 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 222.034
R8026 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t26 184.097
R8027 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t36 184.097
R8028 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t19 184.097
R8029 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t32 184.097
R8030 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n17 166.05
R8031 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n8 166.05
R8032 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n4 57.7228
R8033 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t3 48.0005
R8034 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t0 48.0005
R8035 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t2 48.0005
R8036 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t1 48.0005
R8037 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t5 39.4005
R8038 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t8 39.4005
R8039 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t7 39.4005
R8040 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t9 39.4005
R8041 bgr_0.1st_Vout_2.t10 bgr_0.1st_Vout_2.n21 39.4005
R8042 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.t6 39.4005
R8043 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t17 4.8295
R8044 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t16 4.8295
R8045 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t27 4.8295
R8046 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t23 4.8295
R8047 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t35 4.8295
R8048 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t34 4.8295
R8049 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t28 4.8295
R8050 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R8051 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t15 4.5005
R8052 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t12 4.5005
R8053 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t30 4.5005
R8054 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t22 4.5005
R8055 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t18 4.5005
R8056 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t11 4.5005
R8057 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R8058 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t29 4.5005
R8059 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.5005
R8060 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t24 4.5005
R8061 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R8062 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.5005
R8063 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n11 4.5005
R8064 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n15 4.5005
R8065 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n7 1.3755
R8066 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n16 1.3755
R8067 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 1.188
R8068 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 0.9405
R8069 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n0 0.8935
R8070 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n13 0.78175
R8071 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 0.6585
R8072 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n3 0.6585
R8073 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n1 0.6585
R8074 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n9 0.6255
R8075 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n18 0.6255
R8076 bgr_0.cap_res2 bgr_0.cap_res2.t20 188.315
R8077 bgr_0.cap_res2 bgr_0.cap_res2.t9 0.259
R8078 bgr_0.cap_res2.t13 bgr_0.cap_res2.t8 0.1603
R8079 bgr_0.cap_res2.t2 bgr_0.cap_res2.t6 0.1603
R8080 bgr_0.cap_res2.t5 bgr_0.cap_res2.t1 0.1603
R8081 bgr_0.cap_res2.t19 bgr_0.cap_res2.t0 0.1603
R8082 bgr_0.cap_res2.t14 bgr_0.cap_res2.t10 0.1603
R8083 bgr_0.cap_res2.t4 bgr_0.cap_res2.t7 0.1603
R8084 bgr_0.cap_res2.t18 bgr_0.cap_res2.t16 0.1603
R8085 bgr_0.cap_res2.t12 bgr_0.cap_res2.t15 0.1603
R8086 bgr_0.cap_res2.n1 bgr_0.cap_res2.t17 0.159278
R8087 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.159278
R8088 bgr_0.cap_res2.n3 bgr_0.cap_res2.t3 0.159278
R8089 bgr_0.cap_res2.n3 bgr_0.cap_res2.t13 0.1368
R8090 bgr_0.cap_res2.n3 bgr_0.cap_res2.t2 0.1368
R8091 bgr_0.cap_res2.n2 bgr_0.cap_res2.t5 0.1368
R8092 bgr_0.cap_res2.n2 bgr_0.cap_res2.t19 0.1368
R8093 bgr_0.cap_res2.n1 bgr_0.cap_res2.t14 0.1368
R8094 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R8095 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R8096 bgr_0.cap_res2.n0 bgr_0.cap_res2.t12 0.1368
R8097 bgr_0.cap_res2.t17 bgr_0.cap_res2.n0 0.00152174
R8098 bgr_0.cap_res2.t11 bgr_0.cap_res2.n1 0.00152174
R8099 bgr_0.cap_res2.t3 bgr_0.cap_res2.n2 0.00152174
R8100 bgr_0.cap_res2.t9 bgr_0.cap_res2.n3 0.00152174
R8101 VIN-.n4 VIN-.t8 485.021
R8102 VIN-.n1 VIN-.t6 483.925
R8103 VIN-.n5 VIN-.t7 483.358
R8104 VIN-.n8 VIN-.t10 431.536
R8105 VIN-.n2 VIN-.t9 431.536
R8106 VIN-.n6 VIN-.t1 431.257
R8107 VIN-.n0 VIN-.t0 431.257
R8108 VIN-.n6 VIN-.t2 289.908
R8109 VIN-.n0 VIN-.t5 289.908
R8110 VIN-.n8 VIN-.t4 279.183
R8111 VIN-.n2 VIN-.t3 279.183
R8112 VIN-.n7 VIN-.n6 233.374
R8113 VIN-.n1 VIN-.n0 233.374
R8114 VIN-.n9 VIN-.n8 188.989
R8115 VIN-.n3 VIN-.n2 188.989
R8116 VIN-.n4 VIN-.n3 1.6755
R8117 VIN- VIN-.n9 1.20467
R8118 VIN-.n5 VIN-.n4 1.0755
R8119 VIN-.n3 VIN-.n1 0.883833
R8120 VIN-.n9 VIN-.n7 0.883833
R8121 VIN-.n7 VIN-.n5 0.567167
R8122 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.t8 198.992
R8123 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n8 116.8
R8124 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.n0 113.108
R8125 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.n1 112.564
R8126 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n6 112.002
R8127 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n15 112.002
R8128 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n13 112.002
R8129 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n11 112.002
R8130 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n9 112.002
R8131 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.n2 112.002
R8132 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n4 112.001
R8133 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n19 99.7407
R8134 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.n22 95.3803
R8135 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n34 94.8178
R8136 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.n32 94.8178
R8137 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.n30 94.8178
R8138 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.n28 94.8178
R8139 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.n23 94.8178
R8140 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n20 94.8178
R8141 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.n37 90.3178
R8142 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.n25 90.3178
R8143 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t33 16.0005
R8144 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t21 16.0005
R8145 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t16 16.0005
R8146 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t25 16.0005
R8147 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t17 16.0005
R8148 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t37 16.0005
R8149 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t34 16.0005
R8150 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t22 16.0005
R8151 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t23 16.0005
R8152 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t38 16.0005
R8153 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.t32 16.0005
R8154 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.t20 16.0005
R8155 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t15 16.0005
R8156 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t31 16.0005
R8157 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.t35 16.0005
R8158 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.t19 16.0005
R8159 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t18 16.0005
R8160 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t13 16.0005
R8161 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t24 16.0005
R8162 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t29 16.0005
R8163 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.t26 9.6005
R8164 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.t0 9.6005
R8165 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.t7 9.6005
R8166 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.t39 9.6005
R8167 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.t14 9.6005
R8168 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.t5 9.6005
R8169 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.t36 9.6005
R8170 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.t10 9.6005
R8171 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.t40 9.6005
R8172 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.t9 9.6005
R8173 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.t11 9.6005
R8174 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.t2 9.6005
R8175 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.t4 9.6005
R8176 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.t12 9.6005
R8177 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t3 9.6005
R8178 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t1 9.6005
R8179 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t28 9.6005
R8180 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t6 9.6005
R8181 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.t30 9.6005
R8182 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.t27 9.6005
R8183 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.n26 4.5005
R8184 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.n36 4.5005
R8185 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.n17 4.5005
R8186 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.n16 3.65675
R8187 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.n24 0.563
R8188 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.n27 0.563
R8189 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.n29 0.563
R8190 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.n31 0.563
R8191 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n33 0.563
R8192 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n35 0.563
R8193 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n21 0.563
R8194 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n10 0.563
R8195 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n12 0.563
R8196 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n14 0.563
R8197 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n5 0.563
R8198 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n3 0.563
R8199 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.n7 0.53175
R8200 two_stage_opamp_dummy_magic_0.V_source two_stage_opamp_dummy_magic_0.V_source.n38 0.422375
R8201 two_stage_opamp_dummy_magic_0.V_source two_stage_opamp_dummy_magic_0.V_source.n18 0.328625
R8202 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 610.534
R8203 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 610.534
R8204 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R8205 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R8206 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R8207 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R8208 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 433.8
R8209 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 433.8
R8210 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 433.8
R8211 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R8212 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R8213 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R8214 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 433.8
R8215 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R8216 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R8217 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R8218 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R8219 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R8220 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R8221 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R8222 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.836
R8223 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 339.834
R8224 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R8225 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 334.772
R8226 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 218.266
R8227 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 176.733
R8228 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R8229 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R8230 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R8231 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R8232 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R8233 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R8234 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R8235 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R8236 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R8237 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R8238 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R8239 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R8240 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R8241 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R8242 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 176.733
R8243 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 118.117
R8244 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 65.8738
R8245 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 64.5042
R8246 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n29 57.2661
R8247 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 53.2453
R8248 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 46.5938
R8249 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R8250 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R8251 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R8252 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 39.4005
R8253 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R8254 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R8255 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R8256 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R8257 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n6 18.3911
R8258 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 16.0005
R8259 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R8260 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R8261 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R8262 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 4.5005
R8263 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R8264 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n4 4020
R8265 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n4 4020
R8266 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n10 4020
R8267 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n10 4020
R8268 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t32 660.109
R8269 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t35 660.109
R8270 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n14 422.401
R8271 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n3 422.401
R8272 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.n11 239.915
R8273 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.t33 239.915
R8274 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n8 220.8
R8275 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n6 220.8
R8276 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.n6 188.8
R8277 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n3 188.8
R8278 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 155.911
R8279 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n23 155.91
R8280 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 155.536
R8281 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.n19 155.536
R8282 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n21 155.536
R8283 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 155.535
R8284 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 155.535
R8285 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n28 155.535
R8286 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n26 155.535
R8287 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 155.535
R8288 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t34 155.125
R8289 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t37 155.125
R8290 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n16 151.037
R8291 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.t36 98.2764
R8292 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t4 98.2764
R8293 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.t10 98.2764
R8294 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.t18 98.2764
R8295 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.VD3.t14 98.2764
R8296 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.VD3.t22 98.2764
R8297 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t6 98.2764
R8298 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t12 98.2764
R8299 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t8 98.2764
R8300 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.VD3.t16 98.2764
R8301 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.n13 92.5005
R8302 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 92.5005
R8303 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n10 92.5005
R8304 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n3 92.5005
R8305 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n4 92.5005
R8306 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n4 92.5005
R8307 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t20 49.1384
R8308 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.VD3.n12 49.1384
R8309 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 21.3338
R8310 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 21.3338
R8311 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R8312 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R8313 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R8314 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R8315 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.t19 11.2576
R8316 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R8317 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R8318 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R8319 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R8320 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R8321 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t0 11.2576
R8322 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R8323 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R8324 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R8325 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t26 11.2576
R8326 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R8327 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t28 11.2576
R8328 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t2 11.2576
R8329 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.t29 11.2576
R8330 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R8331 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R8332 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R8333 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 9.488
R8334 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n33 6.51612
R8335 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n22 5.39112
R8336 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.n17 4.5005
R8337 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n25 0.3755
R8338 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.n27 0.3755
R8339 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n29 0.3755
R8340 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n31 0.3755
R8341 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.n20 0.3755
R8342 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.n18 0.3755
R8343 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.n2 0.3755
R8344 a_14240_2076.t0 a_14240_2076.t1 169.905
R8345 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8346 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2595
R8347 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 2280
R8348 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 2250
R8349 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 672.159
R8350 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 672.159
R8351 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 276.8
R8352 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 240
R8353 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 196.8
R8354 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 195.201
R8355 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 174.417
R8356 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 166.034
R8357 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 160.517
R8358 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 160.517
R8359 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 105.909
R8360 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 105.722
R8361 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 95.7988
R8362 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 92.5005
R8363 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 92.5005
R8364 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 92.5005
R8365 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 92.5005
R8366 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8367 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8368 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 75.9449
R8369 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 75.9449
R8370 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 67.2005
R8371 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 47.8997
R8372 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 47.8997
R8373 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 28.8005
R8374 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 23.4672
R8375 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 23.4672
R8376 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 16.8187
R8377 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 16.8187
R8378 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 11.0991
R8379 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 11.0991
R8380 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 10.9449
R8381 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 10.9449
R8382 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 5.60988
R8383 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8384 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t8 661.375
R8385 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t13 611.739
R8386 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t25 611.739
R8387 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.t12 611.739
R8388 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t21 611.739
R8389 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R8390 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R8391 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R8392 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R8393 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R8394 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t20 421.75
R8395 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R8396 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R8397 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R8398 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R8399 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t26 421.75
R8400 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R8401 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R8402 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t11 421.75
R8403 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R8404 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R8405 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 172.667
R8406 two_stage_opamp_dummy_magic_0.Vb3 two_stage_opamp_dummy_magic_0.Vb3.n17 171.84
R8407 two_stage_opamp_dummy_magic_0.Vb3 two_stage_opamp_dummy_magic_0.Vb3.n8 171.376
R8408 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n13 167.094
R8409 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R8410 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R8411 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R8412 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R8413 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R8414 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.n4 167.094
R8415 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R8416 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R8417 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.n0 167.094
R8418 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n1 167.094
R8419 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 167.094
R8420 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n22 139.639
R8421 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 139.638
R8422 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n21 134.577
R8423 two_stage_opamp_dummy_magic_0.Vb3 two_stage_opamp_dummy_magic_0.Vb3.n20 65.6099
R8424 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 40.7027
R8425 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n12 40.7027
R8426 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 40.7027
R8427 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n3 40.7027
R8428 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R8429 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R8430 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R8431 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R8432 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R8433 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R8434 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t0 10.9449
R8435 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t1 10.9449
R8436 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3 7.313
R8437 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n18 6.70362
R8438 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n24 4.5005
R8439 two_stage_opamp_dummy_magic_0.Vb3 two_stage_opamp_dummy_magic_0.Vb3.n25 0.65675
R8440 a_11220_17410.t0 a_11220_17410.t1 258.591
R8441 a_14590_5068.t0 a_14590_5068.t1 433.31
R8442 VIN+.n9 VIN+.t5 485.127
R8443 VIN+.n3 VIN+.t4 485.127
R8444 VIN+.n4 VIN+.t3 485.125
R8445 VIN+.n7 VIN+.t9 318.656
R8446 VIN+.n7 VIN+.t2 318.656
R8447 VIN+.n5 VIN+.t7 318.656
R8448 VIN+.n5 VIN+.t1 318.656
R8449 VIN+.n1 VIN+.t8 318.656
R8450 VIN+.n1 VIN+.t6 318.656
R8451 VIN+.n0 VIN+.t10 318.656
R8452 VIN+.n0 VIN+.t0 318.656
R8453 VIN+.n2 VIN+.n0 166.488
R8454 VIN+.n8 VIN+.n7 165.8
R8455 VIN+.n6 VIN+.n5 165.8
R8456 VIN+.n2 VIN+.n1 165.8
R8457 VIN+.n6 VIN+.n4 1.22862
R8458 VIN+.n4 VIN+.n3 0.7005
R8459 VIN+.n8 VIN+.n6 0.688
R8460 VIN+.n3 VIN+.n2 0.634875
R8461 VIN+.n9 VIN+.n8 0.634875
R8462 VIN+ VIN+.n9 0.50675
R8463 a_13730_17020.t0 a_13730_17020.t1 258.591
R8464 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R8465 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R8466 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t3 303.259
R8467 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R8468 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R8469 bgr_0.V_CUR_REF_REG.t1 bgr_0.V_CUR_REF_REG.n5 245.284
R8470 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t7 174.726
R8471 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 174.726
R8472 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R8473 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R8474 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 96.4005
R8475 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t0 39.4005
R8476 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t2 39.4005
R8477 a_12828_17530.t0 a_12828_17530.t1 376.99
R8478 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8479 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8480 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8481 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8482 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8483 bgr_0.START_UP.n0 bgr_0.START_UP.t1 130.001
R8484 bgr_0.START_UP.n0 bgr_0.START_UP.t0 81.7074
R8485 bgr_0.START_UP bgr_0.START_UP.n0 38.2614
R8486 bgr_0.START_UP bgr_0.START_UP.n5 14.7817
R8487 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8488 bgr_0.START_UP.n1 bgr_0.START_UP.t3 13.1338
R8489 bgr_0.START_UP.n2 bgr_0.START_UP.t4 13.1338
R8490 bgr_0.START_UP.n2 bgr_0.START_UP.t5 13.1338
R8491 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8492 a_11220_17290.t0 a_11220_17290.t1 376.99
R8493 a_12828_17650.t0 a_12828_17650.t1 258.591
R8494 two_stage_opamp_dummy_magic_0.V_p_mir two_stage_opamp_dummy_magic_0.V_p_mir.n0 112.165
R8495 two_stage_opamp_dummy_magic_0.V_p_mir two_stage_opamp_dummy_magic_0.V_p_mir.n1 102.007
R8496 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R8497 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t3 16.0005
R8498 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t2 9.6005
R8499 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t1 9.6005
R8500 a_5750_2076.t0 a_5750_2076.t1 169.905
R8501 a_13790_17550.t0 a_13790_17550.t1 258.591
R8502 a_5280_5068.t0 a_5280_5068.t1 169.905
C0 VOUT- VOUT+ 0.305434f
C1 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.V_err_gate 0.651421f
C2 two_stage_opamp_dummy_magic_0.V_CMFB_S2 VOUT+ 0.228059f
C3 bgr_0.V_TOP VDDA 16.1451f
C4 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.err_amp_out 0.719451f
C5 bgr_0.NFET_GATE_10uA bgr_0.START_UP 0.518703f
C6 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.V_err_gate 0.0135f
C7 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_source 0.318635f
C8 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.V_err_gate 0.080391f
C9 bgr_0.cap_res2 bgr_0.PFET_GATE_10uA 0.018633f
C10 bgr_0.1st_Vout_1 VDDA 2.06087f
C11 two_stage_opamp_dummy_magic_0.cap_res_Y VDDA 1.14388f
C12 two_stage_opamp_dummy_magic_0.Vb3 VOUT+ 0.10139f
C13 two_stage_opamp_dummy_magic_0.X VDDA 6.1633f
C14 bgr_0.Vbe2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.014154f
C15 bgr_0.cap_res2 VDDA 0.586627f
C16 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.050552f
C17 two_stage_opamp_dummy_magic_0.Vb3 bgr_0.Vbe2 0.180547f
C18 two_stage_opamp_dummy_magic_0.V_CMFB_S1 VOUT- 0.019638f
C19 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.01385f
C20 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S2 6.24062f
C21 two_stage_opamp_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S4 9.52539f
C22 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_b_2nd_stage 0.339961f
C23 bgr_0.NFET_GATE_10uA VDDA 1.08124f
C24 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.13839f
C25 two_stage_opamp_dummy_magic_0.VD3 VDDA 4.51742f
C26 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.Vb3 0.058654f
C27 two_stage_opamp_dummy_magic_0.VD4 VDDA 4.77525f
C28 two_stage_opamp_dummy_magic_0.cap_res_Y VOUT- 50.843f
C29 two_stage_opamp_dummy_magic_0.V_CMFB_S1 VOUT+ 0.268674f
C30 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.1st_Vout_1 0.477103f
C31 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.00548f
C32 two_stage_opamp_dummy_magic_0.V_b_2nd_stage VDDA 0.233238f
C33 two_stage_opamp_dummy_magic_0.Vb2_Vb3 VDDA 0.955772f
C34 two_stage_opamp_dummy_magic_0.V_CMFB_S4 VDDA 3.82305f
C35 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_gate 0.33956f
C36 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.V_CMFB_S2 0.964122f
C37 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.551434f
C38 bgr_0.START_UP bgr_0.PFET_GATE_10uA 0.166283f
C39 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.Vb3 0.05378f
C40 two_stage_opamp_dummy_magic_0.V_err_gate VDDA 5.35733f
C41 two_stage_opamp_dummy_magic_0.cap_res_Y VOUT+ 0.028842f
C42 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.Vb3 0.289615f
C43 VIN- VIN+ 0.597231f
C44 two_stage_opamp_dummy_magic_0.X VOUT+ 2.44233f
C45 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.Vb3 0.12531f
C46 bgr_0.START_UP VDDA 1.37621f
C47 bgr_0.Vbe2 bgr_0.V_TOP 0.285619f
C48 bgr_0.PFET_GATE_10uA m2_7180_19780# 0.012f
C49 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.559544f
C50 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_CMFB_S2 0.090225f
C51 two_stage_opamp_dummy_magic_0.V_CMFB_S3 bgr_0.PFET_GATE_10uA 0.345554f
C52 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.V_CMFB_S2 0.024757f
C53 two_stage_opamp_dummy_magic_0.V_p_mir VIN- 0.055745f
C54 bgr_0.V_TOP m2_8540_19780# 0.012f
C55 m2_7180_19780# VDDA 0.010446f
C56 two_stage_opamp_dummy_magic_0.V_b_2nd_stage VOUT- 2.57317f
C57 two_stage_opamp_dummy_magic_0.V_source VIN- 0.416969f
C58 two_stage_opamp_dummy_magic_0.V_CMFB_S1 bgr_0.V_TOP 0.211793f
C59 two_stage_opamp_dummy_magic_0.V_CMFB_S4 VOUT- 0.223667f
C60 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.Vb3 0.489974f
C61 two_stage_opamp_dummy_magic_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.501436f
C62 two_stage_opamp_dummy_magic_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S4 0.572712f
C63 two_stage_opamp_dummy_magic_0.V_CMFB_S3 VDDA 1.91443f
C64 two_stage_opamp_dummy_magic_0.VD1 VIN- 0.948002f
C65 bgr_0.1st_Vout_1 m2_8540_19780# 0.075543f
C66 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.Vb3 1.44805f
C67 bgr_0.PFET_GATE_10uA VDDA 10.4821f
C68 two_stage_opamp_dummy_magic_0.err_amp_out VDDA 1.77275f
C69 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.V_CMFB_S1 0.097112f
C70 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.318695f
C71 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.Vb3 1.24376f
C72 two_stage_opamp_dummy_magic_0.V_p_mir VIN+ 0.14435f
C73 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.V_CMFB_S1 0.794783f
C74 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.61857f
C75 two_stage_opamp_dummy_magic_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.Vb3 0.038649f
C76 two_stage_opamp_dummy_magic_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_err_gate 1.90164f
C77 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb3 0.904138f
C78 two_stage_opamp_dummy_magic_0.V_b_2nd_stage VOUT+ 2.57386f
C79 two_stage_opamp_dummy_magic_0.V_source VIN+ 2.73629f
C80 bgr_0.V_TOP bgr_0.1st_Vout_1 0.925484f
C81 two_stage_opamp_dummy_magic_0.Vb2_Vb3 VOUT+ 0.043377f
C82 two_stage_opamp_dummy_magic_0.V_CMFB_S1 bgr_0.cap_res2 0.092994f
C83 two_stage_opamp_dummy_magic_0.VD1 VIN+ 0.065465f
C84 two_stage_opamp_dummy_magic_0.V_CMFB_S4 bgr_0.START_UP_NFET1 0.011716f
C85 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.09763f
C86 bgr_0.NFET_GATE_10uA bgr_0.Vbe2 0.021455f
C87 two_stage_opamp_dummy_magic_0.Vb3 two_stage_opamp_dummy_magic_0.V_err_gate 14.9057f
C88 two_stage_opamp_dummy_magic_0.V_err_gate VOUT+ 0.095951f
C89 two_stage_opamp_dummy_magic_0.V_source two_stage_opamp_dummy_magic_0.V_p_mir 0.859683f
C90 two_stage_opamp_dummy_magic_0.Vb3 bgr_0.START_UP 0.023308f
C91 bgr_0.cap_res2 bgr_0.1st_Vout_1 0.822981f
C92 two_stage_opamp_dummy_magic_0.cap_res_Y bgr_0.cap_res2 0.048779f
C93 two_stage_opamp_dummy_magic_0.V_CMFB_S1 bgr_0.NFET_GATE_10uA 0.067783f
C94 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.VD1 1.05762f
C95 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C96 two_stage_opamp_dummy_magic_0.V_CMFB_S3 VOUT- 0.26403f
C97 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.V_source 0.979041f
C98 two_stage_opamp_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.505117f
C99 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.577673f
C100 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.4652f
C101 bgr_0.NFET_GATE_10uA bgr_0.V_TOP 0.080353f
C102 two_stage_opamp_dummy_magic_0.V_b_2nd_stage VIN+ 0.107903f
C103 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S4 1.85524f
C104 bgr_0.NFET_GATE_10uA bgr_0.1st_Vout_1 1.02268f
C105 bgr_0.START_UP bgr_0.Vbe2 0.193132f
C106 VDDA VOUT- 6.81753f
C107 two_stage_opamp_dummy_magic_0.V_err_amp_ref VDDA 5.17627f
C108 two_stage_opamp_dummy_magic_0.V_CMFB_S2 VDDA 3.86448f
C109 two_stage_opamp_dummy_magic_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_err_gate 0.529958f
C110 two_stage_opamp_dummy_magic_0.err_amp_out VOUT+ 0.01087f
C111 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.VD3 3.51341f
C112 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.VD4 0.035948f
C113 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.V_b_2nd_stage 0.066774f
C114 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.V_CMFB_S4 0.563927f
C115 two_stage_opamp_dummy_magic_0.V_p_mir two_stage_opamp_dummy_magic_0.V_b_2nd_stage 0.165253f
C116 two_stage_opamp_dummy_magic_0.Vb3 VDDA 5.84291f
C117 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.V_b_2nd_stage 0.017284f
C118 two_stage_opamp_dummy_magic_0.V_source two_stage_opamp_dummy_magic_0.V_b_2nd_stage 2.55867f
C119 VDDA VOUT+ 6.753f
C120 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage 0.010152f
C121 bgr_0.START_UP_NFET1 VDDA 0.150493f
C122 bgr_0.Vbe2 bgr_0.PFET_GATE_10uA 0.242909f
C123 bgr_0.START_UP bgr_0.V_TOP 0.815644f
C124 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.V_err_gate 0.218048f
C125 bgr_0.START_UP bgr_0.1st_Vout_1 0.030647f
C126 bgr_0.Vbe2 VDDA 0.02318f
C127 two_stage_opamp_dummy_magic_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S1 0.128019f
C128 two_stage_opamp_dummy_magic_0.V_CMFB_S1 bgr_0.PFET_GATE_10uA 1.72424f
C129 two_stage_opamp_dummy_magic_0.V_err_amp_ref VOUT- 0.11443f
C130 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_CMFB_S4 0.053993f
C131 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD3 0.107225f
C132 two_stage_opamp_dummy_magic_0.V_CMFB_S3 bgr_0.V_TOP 0.032614f
C133 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.VD3 0.079359f
C134 m2_8540_19780# VDDA 0.010446f
C135 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 2.47366f
C136 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.V_CMFB_S4 0.024757f
C137 two_stage_opamp_dummy_magic_0.V_CMFB_S1 VDDA 3.31408f
C138 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.V_CMFB_S3 0.660179f
C139 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 0.145581f
C140 two_stage_opamp_dummy_magic_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.Vb3 0.272073f
C141 bgr_0.PFET_GATE_10uA bgr_0.1st_Vout_1 0.035393f
C142 VIN+ GNDA 2.10937f
C143 VIN- GNDA 2.159328f
C144 VOUT+ GNDA 17.91994f
C145 VOUT- GNDA 17.84433f
C146 VDDA GNDA 0.152182p
C147 two_stage_opamp_dummy_magic_0.V_b_2nd_stage GNDA 7.5997f
C148 two_stage_opamp_dummy_magic_0.V_p_mir GNDA 0.810478f
C149 two_stage_opamp_dummy_magic_0.V_source GNDA 8.309299f
C150 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.62122f
C151 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.895637f
C152 two_stage_opamp_dummy_magic_0.cap_res_Y GNDA 32.792385f
C153 two_stage_opamp_dummy_magic_0.X GNDA 5.64241f
C154 bgr_0.cap_res2 GNDA 7.923826f
C155 two_stage_opamp_dummy_magic_0.V_CMFB_S1 GNDA 13.349511f
C156 two_stage_opamp_dummy_magic_0.V_CMFB_S3 GNDA 9.152886f
C157 bgr_0.1st_Vout_1 GNDA 4.985791f
C158 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 18.89328f
C159 bgr_0.V_TOP GNDA 6.831777f
C160 bgr_0.PFET_GATE_10uA GNDA 5.08629f
C161 bgr_0.Vbe2 GNDA 17.0692f
C162 bgr_0.START_UP GNDA 7.196543f
C163 bgr_0.START_UP_NFET1 GNDA 5.28327f
C164 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 18.889242f
C165 two_stage_opamp_dummy_magic_0.Vb3 GNDA 19.293179f
C166 two_stage_opamp_dummy_magic_0.V_CMFB_S4 GNDA 16.472971f
C167 two_stage_opamp_dummy_magic_0.V_CMFB_S2 GNDA 23.537739f
C168 bgr_0.NFET_GATE_10uA GNDA 7.33111f
C169 two_stage_opamp_dummy_magic_0.VD3 GNDA 6.465442f
C170 two_stage_opamp_dummy_magic_0.VD4 GNDA 6.52597f
C171 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.66568f
C172 bgr_0.START_UP.t0 GNDA 1.6623f
C173 bgr_0.START_UP.t1 GNDA 0.043697f
C174 bgr_0.START_UP.n0 GNDA 1.12862f
C175 bgr_0.START_UP.t2 GNDA 0.041701f
C176 bgr_0.START_UP.t3 GNDA 0.041701f
C177 bgr_0.START_UP.n1 GNDA 0.151283f
C178 bgr_0.START_UP.t4 GNDA 0.041701f
C179 bgr_0.START_UP.t5 GNDA 0.041701f
C180 bgr_0.START_UP.n2 GNDA 0.139173f
C181 bgr_0.START_UP.n3 GNDA 0.720787f
C182 bgr_0.START_UP.t7 GNDA 0.01567f
C183 bgr_0.START_UP.t6 GNDA 0.01567f
C184 bgr_0.START_UP.n4 GNDA 0.044238f
C185 bgr_0.START_UP.n5 GNDA 0.445182f
C186 bgr_0.V_CUR_REF_REG.t3 GNDA 0.014208f
C187 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C188 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C189 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C190 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C191 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C192 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C193 bgr_0.V_CUR_REF_REG.t1 GNDA 0.42777f
C194 VIN+.t0 GNDA 0.036562f
C195 VIN+.t10 GNDA 0.036562f
C196 VIN+.n0 GNDA 0.075254f
C197 VIN+.t6 GNDA 0.036562f
C198 VIN+.t8 GNDA 0.036562f
C199 VIN+.n1 GNDA 0.074514f
C200 VIN+.n2 GNDA 0.428602f
C201 VIN+.t4 GNDA 0.051438f
C202 VIN+.n3 GNDA 0.267734f
C203 VIN+.t3 GNDA 0.051438f
C204 VIN+.n4 GNDA 0.350523f
C205 VIN+.t1 GNDA 0.036562f
C206 VIN+.t7 GNDA 0.036562f
C207 VIN+.n5 GNDA 0.074514f
C208 VIN+.n6 GNDA 0.332972f
C209 VIN+.t2 GNDA 0.036562f
C210 VIN+.t9 GNDA 0.036562f
C211 VIN+.n7 GNDA 0.074514f
C212 VIN+.n8 GNDA 0.250183f
C213 VIN+.t5 GNDA 0.051438f
C214 VIN+.n9 GNDA 0.240718f
C215 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.163549f
C216 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.130451f
C217 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.130451f
C218 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.130451f
C219 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.130451f
C220 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.150539f
C221 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.122221f
C222 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.075108f
C223 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.075108f
C224 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.071883f
C225 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.130451f
C226 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.130451f
C227 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.130451f
C228 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.130451f
C229 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.150539f
C230 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.122221f
C231 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.075108f
C232 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.075108f
C233 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.071883f
C234 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.072871f
C235 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.130451f
C236 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.130451f
C237 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.130451f
C238 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.130451f
C239 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.150539f
C240 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.122221f
C241 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.075108f
C242 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.075108f
C243 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.071883f
C244 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.130451f
C245 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.130451f
C246 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.130451f
C247 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.130451f
C248 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.150539f
C249 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.122221f
C250 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.075108f
C251 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.075108f
C252 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.071883f
C253 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.077166f
C254 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.97833f
C255 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.094873f
C256 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.094873f
C257 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.340545f
C258 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 7.854681f
C259 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.026354f
C260 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.026354f
C261 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.079599f
C262 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.026354f
C263 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.026354f
C264 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.084888f
C265 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.026354f
C266 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.026354f
C267 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 0.084888f
C268 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.467983f
C269 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.228738f
C270 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.025546f
C271 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.025546f
C272 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.087918f
C273 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.025546f
C274 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.025546f
C275 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.087704f
C276 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.189325f
C277 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.070868f
C278 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.098895f
C279 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.126025f
C280 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.044485f
C281 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.08331f
C282 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.055614f
C283 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.126025f
C284 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.044485f
C285 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.08331f
C286 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.055614f
C287 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.050363f
C288 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.098895f
C289 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.294724f
C290 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.439919f
C291 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.254003f
C292 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.254003f
C293 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.254003f
C294 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.254003f
C295 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.190502f
C296 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.127002f
C297 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.190502f
C298 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.254003f
C299 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.254003f
C300 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.254003f
C301 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.254003f
C302 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.439919f
C303 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.294724f
C304 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.070868f
C305 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.106202f
C306 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.025546f
C307 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.025546f
C308 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.08575f
C309 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.073309f
C310 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.035035f
C311 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.025546f
C312 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.025546f
C313 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.087704f
C314 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.100609f
C315 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.025546f
C316 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.025546f
C317 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.087704f
C318 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.150083f
C319 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.025546f
C320 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.025546f
C321 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.087918f
C322 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.025546f
C323 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.025546f
C324 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.087704f
C325 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.189325f
C326 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.025546f
C327 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.025546f
C328 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.087704f
C329 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.100608f
C330 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.025546f
C331 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.025546f
C332 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.087704f
C333 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.100608f
C334 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.025546f
C335 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.025546f
C336 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.087704f
C337 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.100608f
C338 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.025546f
C339 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.025546f
C340 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.087704f
C341 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.175735f
C342 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.024321f
C343 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.024321f
C344 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.058658f
C345 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.024321f
C346 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.024321f
C347 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.060884f
C348 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.024321f
C349 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.024321f
C350 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.060557f
C351 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.411197f
C352 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.024321f
C353 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.024321f
C354 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.060884f
C355 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.269887f
C356 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.626981f
C357 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.036482f
C358 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.036482f
C359 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.132506f
C360 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.064756f
C361 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.064756f
C362 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.064756f
C363 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.064756f
C364 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.064756f
C365 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.064756f
C366 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.064756f
C367 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.064756f
C368 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.064756f
C369 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.07558f
C370 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.07126f
C371 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.04469f
C372 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.04469f
C373 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.04469f
C374 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.04469f
C375 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.04469f
C376 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.04469f
C377 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.04469f
C378 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.040177f
C379 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.064756f
C380 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.064756f
C381 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.064756f
C382 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.064756f
C383 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.064756f
C384 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.064756f
C385 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.064756f
C386 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.064756f
C387 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.064756f
C388 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.07558f
C389 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.07126f
C390 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.04469f
C391 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.04469f
C392 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.04469f
C393 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.04469f
C394 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.04469f
C395 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.04469f
C396 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.04469f
C397 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.039819f
C398 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.11518f
C399 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.036482f
C400 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.036482f
C401 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.072964f
C402 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.338266f
C403 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 5.42356f
C404 bgr_0.TAIL_CUR_MIR_BIAS GNDA 5.36303f
C405 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA 0.014411f
C406 two_stage_opamp_dummy_magic_0.V_source.t25 GNDA 0.014411f
C407 two_stage_opamp_dummy_magic_0.V_source.n0 GNDA 0.048951f
C408 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA 0.014411f
C409 two_stage_opamp_dummy_magic_0.V_source.t13 GNDA 0.014411f
C410 two_stage_opamp_dummy_magic_0.V_source.n1 GNDA 0.051603f
C411 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA 0.014411f
C412 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA 0.014411f
C413 two_stage_opamp_dummy_magic_0.V_source.n2 GNDA 0.051153f
C414 two_stage_opamp_dummy_magic_0.V_source.n3 GNDA 0.186431f
C415 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA 0.014411f
C416 two_stage_opamp_dummy_magic_0.V_source.t29 GNDA 0.014411f
C417 two_stage_opamp_dummy_magic_0.V_source.n4 GNDA 0.051153f
C418 two_stage_opamp_dummy_magic_0.V_source.n5 GNDA 0.096803f
C419 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA 0.014411f
C420 two_stage_opamp_dummy_magic_0.V_source.t21 GNDA 0.014411f
C421 two_stage_opamp_dummy_magic_0.V_source.n6 GNDA 0.051153f
C422 two_stage_opamp_dummy_magic_0.V_source.n7 GNDA 0.096323f
C423 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA 0.014411f
C424 two_stage_opamp_dummy_magic_0.V_source.t31 GNDA 0.014411f
C425 two_stage_opamp_dummy_magic_0.V_source.n8 GNDA 0.051839f
C426 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA 0.014411f
C427 two_stage_opamp_dummy_magic_0.V_source.t20 GNDA 0.014411f
C428 two_stage_opamp_dummy_magic_0.V_source.n9 GNDA 0.051153f
C429 two_stage_opamp_dummy_magic_0.V_source.n10 GNDA 0.183313f
C430 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA 0.014411f
C431 two_stage_opamp_dummy_magic_0.V_source.t38 GNDA 0.014411f
C432 two_stage_opamp_dummy_magic_0.V_source.n11 GNDA 0.051153f
C433 two_stage_opamp_dummy_magic_0.V_source.n12 GNDA 0.096803f
C434 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA 0.014411f
C435 two_stage_opamp_dummy_magic_0.V_source.t22 GNDA 0.014411f
C436 two_stage_opamp_dummy_magic_0.V_source.n13 GNDA 0.051153f
C437 two_stage_opamp_dummy_magic_0.V_source.n14 GNDA 0.096803f
C438 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA 0.014411f
C439 two_stage_opamp_dummy_magic_0.V_source.t37 GNDA 0.014411f
C440 two_stage_opamp_dummy_magic_0.V_source.n15 GNDA 0.051153f
C441 two_stage_opamp_dummy_magic_0.V_source.n16 GNDA 0.144361f
C442 two_stage_opamp_dummy_magic_0.V_source.n17 GNDA 0.0759f
C443 two_stage_opamp_dummy_magic_0.V_source.n18 GNDA 0.076908f
C444 two_stage_opamp_dummy_magic_0.V_source.t30 GNDA 0.024019f
C445 two_stage_opamp_dummy_magic_0.V_source.t27 GNDA 0.024019f
C446 two_stage_opamp_dummy_magic_0.V_source.n19 GNDA 0.095892f
C447 two_stage_opamp_dummy_magic_0.V_source.t28 GNDA 0.024019f
C448 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA 0.024019f
C449 two_stage_opamp_dummy_magic_0.V_source.n20 GNDA 0.094792f
C450 two_stage_opamp_dummy_magic_0.V_source.n21 GNDA 0.168638f
C451 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA 0.024019f
C452 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA 0.024019f
C453 two_stage_opamp_dummy_magic_0.V_source.n22 GNDA 0.09527f
C454 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA 0.024019f
C455 two_stage_opamp_dummy_magic_0.V_source.t12 GNDA 0.024019f
C456 two_stage_opamp_dummy_magic_0.V_source.n23 GNDA 0.094792f
C457 two_stage_opamp_dummy_magic_0.V_source.n24 GNDA 0.1683f
C458 two_stage_opamp_dummy_magic_0.V_source.t8 GNDA 0.120338f
C459 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA 0.024019f
C460 two_stage_opamp_dummy_magic_0.V_source.t2 GNDA 0.024019f
C461 two_stage_opamp_dummy_magic_0.V_source.n25 GNDA 0.091856f
C462 two_stage_opamp_dummy_magic_0.V_source.n26 GNDA 1.02382f
C463 two_stage_opamp_dummy_magic_0.V_source.n27 GNDA 0.028823f
C464 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA 0.024019f
C465 two_stage_opamp_dummy_magic_0.V_source.t9 GNDA 0.024019f
C466 two_stage_opamp_dummy_magic_0.V_source.n28 GNDA 0.094792f
C467 two_stage_opamp_dummy_magic_0.V_source.n29 GNDA 0.087751f
C468 two_stage_opamp_dummy_magic_0.V_source.t36 GNDA 0.024019f
C469 two_stage_opamp_dummy_magic_0.V_source.t10 GNDA 0.024019f
C470 two_stage_opamp_dummy_magic_0.V_source.n30 GNDA 0.094792f
C471 two_stage_opamp_dummy_magic_0.V_source.n31 GNDA 0.087751f
C472 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA 0.024019f
C473 two_stage_opamp_dummy_magic_0.V_source.t5 GNDA 0.024019f
C474 two_stage_opamp_dummy_magic_0.V_source.n32 GNDA 0.094792f
C475 two_stage_opamp_dummy_magic_0.V_source.n33 GNDA 0.087751f
C476 two_stage_opamp_dummy_magic_0.V_source.t7 GNDA 0.024019f
C477 two_stage_opamp_dummy_magic_0.V_source.t39 GNDA 0.024019f
C478 two_stage_opamp_dummy_magic_0.V_source.n34 GNDA 0.094792f
C479 two_stage_opamp_dummy_magic_0.V_source.n35 GNDA 0.087751f
C480 two_stage_opamp_dummy_magic_0.V_source.n36 GNDA 0.028823f
C481 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA 0.024019f
C482 two_stage_opamp_dummy_magic_0.V_source.t0 GNDA 0.024019f
C483 two_stage_opamp_dummy_magic_0.V_source.n37 GNDA 0.091856f
C484 two_stage_opamp_dummy_magic_0.V_source.n38 GNDA 0.086382f
C485 VIN-.t6 GNDA 0.046059f
C486 VIN-.t5 GNDA 0.030419f
C487 VIN-.t0 GNDA 0.037555f
C488 VIN-.n0 GNDA 0.053964f
C489 VIN-.n1 GNDA 0.293957f
C490 VIN-.t3 GNDA 0.029919f
C491 VIN-.t9 GNDA 0.037568f
C492 VIN-.n2 GNDA 0.059078f
C493 VIN-.n3 GNDA 0.237445f
C494 VIN-.t8 GNDA 0.045592f
C495 VIN-.n4 GNDA 0.274074f
C496 VIN-.t7 GNDA 0.045908f
C497 VIN-.n5 GNDA 0.197794f
C498 VIN-.t2 GNDA 0.030419f
C499 VIN-.t1 GNDA 0.037555f
C500 VIN-.n6 GNDA 0.053964f
C501 VIN-.n7 GNDA 0.165144f
C502 VIN-.t4 GNDA 0.029919f
C503 VIN-.t10 GNDA 0.037568f
C504 VIN-.n8 GNDA 0.059078f
C505 VIN-.n9 GNDA 0.204653f
C506 bgr_0.cap_res2.t6 GNDA 0.406156f
C507 bgr_0.cap_res2.t2 GNDA 0.407628f
C508 bgr_0.cap_res2.t8 GNDA 0.406156f
C509 bgr_0.cap_res2.t13 GNDA 0.407628f
C510 bgr_0.cap_res2.t0 GNDA 0.406156f
C511 bgr_0.cap_res2.t19 GNDA 0.407628f
C512 bgr_0.cap_res2.t1 GNDA 0.406156f
C513 bgr_0.cap_res2.t5 GNDA 0.407628f
C514 bgr_0.cap_res2.t7 GNDA 0.406156f
C515 bgr_0.cap_res2.t4 GNDA 0.407628f
C516 bgr_0.cap_res2.t10 GNDA 0.406156f
C517 bgr_0.cap_res2.t14 GNDA 0.407628f
C518 bgr_0.cap_res2.t15 GNDA 0.406156f
C519 bgr_0.cap_res2.t12 GNDA 0.407628f
C520 bgr_0.cap_res2.t16 GNDA 0.406156f
C521 bgr_0.cap_res2.t18 GNDA 0.407628f
C522 bgr_0.cap_res2.n0 GNDA 0.272247f
C523 bgr_0.cap_res2.t17 GNDA 0.216805f
C524 bgr_0.cap_res2.n1 GNDA 0.295394f
C525 bgr_0.cap_res2.t11 GNDA 0.216805f
C526 bgr_0.cap_res2.n2 GNDA 0.295394f
C527 bgr_0.cap_res2.t3 GNDA 0.216805f
C528 bgr_0.cap_res2.n3 GNDA 0.295394f
C529 bgr_0.cap_res2.t9 GNDA 0.214043f
C530 bgr_0.cap_res2.t20 GNDA 0.133038f
C531 bgr_0.1st_Vout_2.n0 GNDA 0.995956f
C532 bgr_0.1st_Vout_2.n1 GNDA 0.240335f
C533 bgr_0.1st_Vout_2.n2 GNDA 0.995956f
C534 bgr_0.1st_Vout_2.n3 GNDA 0.240335f
C535 bgr_0.1st_Vout_2.n4 GNDA 0.805677f
C536 bgr_0.1st_Vout_2.n5 GNDA 0.240335f
C537 bgr_0.1st_Vout_2.t13 GNDA 0.021508f
C538 bgr_0.1st_Vout_2.n6 GNDA 0.02259f
C539 bgr_0.1st_Vout_2.n7 GNDA 0.171874f
C540 bgr_0.1st_Vout_2.t32 GNDA 0.013652f
C541 bgr_0.1st_Vout_2.t19 GNDA 0.013652f
C542 bgr_0.1st_Vout_2.n8 GNDA 0.03037f
C543 bgr_0.1st_Vout_2.n9 GNDA 0.083918f
C544 bgr_0.1st_Vout_2.n10 GNDA 0.012945f
C545 bgr_0.1st_Vout_2.t4 GNDA 0.018875f
C546 bgr_0.1st_Vout_2.n11 GNDA 0.195802f
C547 bgr_0.1st_Vout_2.n12 GNDA 0.011712f
C548 bgr_0.1st_Vout_2.n13 GNDA 0.049674f
C549 bgr_0.1st_Vout_2.n14 GNDA 0.021654f
C550 bgr_0.1st_Vout_2.n15 GNDA 0.080059f
C551 bgr_0.1st_Vout_2.n16 GNDA 0.03943f
C552 bgr_0.1st_Vout_2.t36 GNDA 0.013652f
C553 bgr_0.1st_Vout_2.t26 GNDA 0.013652f
C554 bgr_0.1st_Vout_2.n17 GNDA 0.03037f
C555 bgr_0.1st_Vout_2.n18 GNDA 0.083918f
C556 bgr_0.1st_Vout_2.t17 GNDA 0.364565f
C557 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C558 bgr_0.1st_Vout_2.t15 GNDA 0.358459f
C559 bgr_0.1st_Vout_2.t16 GNDA 0.364565f
C560 bgr_0.1st_Vout_2.t12 GNDA 0.358459f
C561 bgr_0.1st_Vout_2.t27 GNDA 0.364565f
C562 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C563 bgr_0.1st_Vout_2.t22 GNDA 0.358459f
C564 bgr_0.1st_Vout_2.t23 GNDA 0.364565f
C565 bgr_0.1st_Vout_2.t18 GNDA 0.358459f
C566 bgr_0.1st_Vout_2.t35 GNDA 0.364565f
C567 bgr_0.1st_Vout_2.t11 GNDA 0.358459f
C568 bgr_0.1st_Vout_2.t31 GNDA 0.358459f
C569 bgr_0.1st_Vout_2.t34 GNDA 0.364565f
C570 bgr_0.1st_Vout_2.t29 GNDA 0.358459f
C571 bgr_0.1st_Vout_2.t28 GNDA 0.364565f
C572 bgr_0.1st_Vout_2.t33 GNDA 0.358459f
C573 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C574 bgr_0.1st_Vout_2.t20 GNDA 0.358459f
C575 bgr_0.1st_Vout_2.t25 GNDA 0.358459f
C576 bgr_0.1st_Vout_2.t14 GNDA 0.023417f
C577 bgr_0.1st_Vout_2.n19 GNDA 0.516024f
C578 bgr_0.1st_Vout_2.n20 GNDA 0.106455f
C579 bgr_0.1st_Vout_2.n21 GNDA 0.02259f
C580 bgr_0.Vin+.t6 GNDA 0.020459f
C581 bgr_0.Vin+.t8 GNDA 0.013299f
C582 bgr_0.Vin+.n0 GNDA 0.04388f
C583 bgr_0.Vin+.t10 GNDA 0.013299f
C584 bgr_0.Vin+.n1 GNDA 0.034146f
C585 bgr_0.Vin+.t7 GNDA 0.013299f
C586 bgr_0.Vin+.n2 GNDA 0.034607f
C587 bgr_0.Vin+.n3 GNDA 0.074523f
C588 bgr_0.Vin+.t4 GNDA 0.043132f
C589 bgr_0.Vin+.t3 GNDA 0.043132f
C590 bgr_0.Vin+.n4 GNDA 0.144858f
C591 bgr_0.Vin+.t2 GNDA 0.043132f
C592 bgr_0.Vin+.t5 GNDA 0.043132f
C593 bgr_0.Vin+.n5 GNDA 0.142495f
C594 bgr_0.Vin+.n6 GNDA 0.656763f
C595 bgr_0.Vin+.n7 GNDA 0.71769f
C596 bgr_0.Vin+.t1 GNDA 0.125873f
C597 bgr_0.Vin+.n8 GNDA 0.446219f
C598 bgr_0.Vin+.t0 GNDA 0.137433f
C599 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.013337f
C600 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.013337f
C601 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.033433f
C602 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.013337f
C603 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.013337f
C604 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.033256f
C605 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.295581f
C606 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.013337f
C607 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.013337f
C608 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.026675f
C609 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.149082f
C610 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 3.24594f
C611 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.170331f
C612 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.026675f
C613 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.026675f
C614 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.077329f
C615 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.026675f
C616 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.026675f
C617 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.077085f
C618 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.304398f
C619 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.026675f
C620 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.026675f
C621 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.077085f
C622 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.161657f
C623 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.026675f
C624 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.026675f
C625 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.077085f
C626 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.161657f
C627 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.026675f
C628 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.026675f
C629 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.077085f
C630 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 0.291832f
C631 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 0.574104f
C632 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.018562f
C633 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.017814f
C634 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.017897f
C635 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.018631f
C636 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.018518f
C637 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.263092f
C638 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.018518f
C639 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.137234f
C640 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.018518f
C641 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.167483f
C642 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.173327f
C643 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.155565f
C644 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.30324f
C645 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.018562f
C646 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.018383f
C647 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.381398f
C648 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.018383f
C649 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.21975f
C650 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.21975f
C651 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.018383f
C652 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.233772f
C653 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.588067f
C654 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.588067f
C655 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.697944f
C656 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.368648f
C657 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.233458f
C658 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.638139f
C659 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.222663f
C660 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 1.15528f
C661 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.233772f
C662 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.641216f
C663 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.588067f
C664 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.588067f
C665 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.697944f
C666 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.368648f
C667 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.23331f
C668 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.215887f
C669 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 1.41875f
C670 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.02014f
C671 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.02014f
C672 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.061008f
C673 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.02014f
C674 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.02014f
C675 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.076053f
C676 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.471161f
C677 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.265651f
C678 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.080559f
C679 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.080559f
C680 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.347776f
C681 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.080559f
C682 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.080559f
C683 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.347073f
C684 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.400756f
C685 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.080559f
C686 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.080559f
C687 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.347073f
C688 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.214827f
C689 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.080559f
C690 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.080559f
C691 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.347073f
C692 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.214827f
C693 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.080559f
C694 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.080559f
C695 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.347073f
C696 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.374181f
C697 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.956082f
C698 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.344611f
C699 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.34586f
C700 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.344611f
C701 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.347313f
C702 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.377753f
C703 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.344611f
C704 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.34586f
C705 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.344611f
C706 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.34586f
C707 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344611f
C708 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.34586f
C709 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.344611f
C710 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.34586f
C711 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.344611f
C712 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.34586f
C713 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.344611f
C714 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.34586f
C715 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.344611f
C716 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.34586f
C717 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.344611f
C718 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.34586f
C719 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.344611f
C720 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.34586f
C721 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.344611f
C722 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.34586f
C723 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.344611f
C724 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.34586f
C725 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.344611f
C726 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.34586f
C727 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.344611f
C728 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.34586f
C729 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.344611f
C730 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.34586f
C731 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.344611f
C732 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.34586f
C733 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.344611f
C734 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.34586f
C735 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.344611f
C736 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.34586f
C737 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.344611f
C738 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.34586f
C739 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.344611f
C740 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.34586f
C741 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.344611f
C742 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.34586f
C743 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344611f
C744 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.34586f
C745 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.344611f
C746 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.34586f
C747 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.344611f
C748 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.34586f
C749 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.344611f
C750 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.34586f
C751 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.344611f
C752 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.34586f
C753 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.344611f
C754 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.34586f
C755 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.344611f
C756 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.34586f
C757 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.344611f
C758 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.34586f
C759 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.344611f
C760 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.34586f
C761 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.344611f
C762 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.361508f
C763 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.344611f
C764 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.185098f
C765 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.1981f
C766 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.344611f
C767 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.185098f
C768 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.196502f
C769 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.344611f
C770 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.185098f
C771 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.196502f
C772 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.344611f
C773 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185098f
C774 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.196502f
C775 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.344611f
C776 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.185098f
C777 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.196502f
C778 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.344611f
C779 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.185098f
C780 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.196502f
C781 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.344611f
C782 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.185098f
C783 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.196502f
C784 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.344611f
C785 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.185098f
C786 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.196502f
C787 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.344611f
C788 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.185098f
C789 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.196502f
C790 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.344611f
C791 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.34586f
C792 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.166603f
C793 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.214893f
C794 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.183952f
C795 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.233388f
C796 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.183952f
C797 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.250633f
C798 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.183952f
C799 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.250633f
C800 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.183952f
C801 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.250633f
C802 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.183952f
C803 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.250633f
C804 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.183952f
C805 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.250633f
C806 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.183952f
C807 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.250633f
C808 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.183952f
C809 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.250633f
C810 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.183952f
C811 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.250633f
C812 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.183952f
C813 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.250633f
C814 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.183952f
C815 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.250633f
C816 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.183952f
C817 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.250633f
C818 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.183952f
C819 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.250633f
C820 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.183952f
C821 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.250633f
C822 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.183952f
C823 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.250633f
C824 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.183952f
C825 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.233388f
C826 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.343466f
C827 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.166603f
C828 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.216142f
C829 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.343466f
C830 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.166603f
C831 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.216142f
C832 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.343466f
C833 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.344611f
C834 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.363106f
C835 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.363106f
C836 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185098f
C837 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.216142f
C838 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.343466f
C839 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.344611f
C840 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.185098f
C841 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.197648f
C842 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.343466f
C843 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.344611f
C844 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.185098f
C845 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.216142f
C846 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.343466f
C847 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.344611f
C848 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.185098f
C849 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.216142f
C850 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.343466f
C851 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344611f
C852 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.185098f
C853 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216142f
C854 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.343466f
C855 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.344611f
C856 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.363106f
C857 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.363106f
C858 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.185098f
C859 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216142f
C860 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.343466f
C861 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.344611f
C862 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.363106f
C863 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.363106f
C864 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.185098f
C865 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216142f
C866 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.343466f
C867 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216142f
C868 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.185098f
C869 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.363106f
C870 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.363106f
C871 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.769243f
C872 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.303799f
C873 bgr_0.V_mir1.t8 GNDA 0.053881f
C874 bgr_0.V_mir1.t6 GNDA 0.042444f
C875 bgr_0.V_mir1.t17 GNDA 0.042444f
C876 bgr_0.V_mir1.t20 GNDA 0.06851f
C877 bgr_0.V_mir1.n0 GNDA 0.076506f
C878 bgr_0.V_mir1.n1 GNDA 0.052264f
C879 bgr_0.V_mir1.n2 GNDA 0.081315f
C880 bgr_0.V_mir1.t9 GNDA 0.03537f
C881 bgr_0.V_mir1.t7 GNDA 0.03537f
C882 bgr_0.V_mir1.n3 GNDA 0.08097f
C883 bgr_0.V_mir1.n4 GNDA 0.203577f
C884 bgr_0.V_mir1.t12 GNDA 0.017685f
C885 bgr_0.V_mir1.t13 GNDA 0.017685f
C886 bgr_0.V_mir1.n5 GNDA 0.046242f
C887 bgr_0.V_mir1.t15 GNDA 0.075466f
C888 bgr_0.V_mir1.t14 GNDA 0.017685f
C889 bgr_0.V_mir1.t16 GNDA 0.017685f
C890 bgr_0.V_mir1.n6 GNDA 0.050199f
C891 bgr_0.V_mir1.n7 GNDA 0.827814f
C892 bgr_0.V_mir1.n8 GNDA 0.268286f
C893 bgr_0.V_mir1.t0 GNDA 0.053881f
C894 bgr_0.V_mir1.t4 GNDA 0.042444f
C895 bgr_0.V_mir1.t18 GNDA 0.042444f
C896 bgr_0.V_mir1.t21 GNDA 0.06851f
C897 bgr_0.V_mir1.n9 GNDA 0.076506f
C898 bgr_0.V_mir1.n10 GNDA 0.052264f
C899 bgr_0.V_mir1.n11 GNDA 0.081315f
C900 bgr_0.V_mir1.t1 GNDA 0.03537f
C901 bgr_0.V_mir1.t5 GNDA 0.03537f
C902 bgr_0.V_mir1.n12 GNDA 0.08097f
C903 bgr_0.V_mir1.n13 GNDA 0.156007f
C904 bgr_0.V_mir1.n14 GNDA 0.09373f
C905 bgr_0.V_mir1.n15 GNDA 0.699157f
C906 bgr_0.V_mir1.t10 GNDA 0.053881f
C907 bgr_0.V_mir1.t2 GNDA 0.042444f
C908 bgr_0.V_mir1.t19 GNDA 0.042444f
C909 bgr_0.V_mir1.t22 GNDA 0.06851f
C910 bgr_0.V_mir1.n16 GNDA 0.076506f
C911 bgr_0.V_mir1.n17 GNDA 0.052264f
C912 bgr_0.V_mir1.n18 GNDA 0.081315f
C913 bgr_0.V_mir1.n19 GNDA 0.201563f
C914 bgr_0.V_mir1.t3 GNDA 0.03537f
C915 bgr_0.V_mir1.n20 GNDA 0.08097f
C916 bgr_0.V_mir1.t11 GNDA 0.03537f
C917 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.018232f
C918 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.018232f
C919 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.066269f
C920 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.018232f
C921 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.018232f
C922 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.055069f
C923 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.380049f
C924 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.227039f
C925 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.072929f
C926 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.072929f
C927 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.314837f
C928 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.072929f
C929 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.072929f
C930 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.3142f
C931 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.362799f
C932 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.072929f
C933 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.072929f
C934 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.3142f
C935 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.19448f
C936 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.072929f
C937 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.072929f
C938 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.3142f
C939 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.19448f
C940 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.072929f
C941 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.072929f
C942 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.3142f
C943 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.338741f
C944 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.587263f
C945 two_stage_opamp_dummy_magic_0.Vb1.n2 GNDA 0.084204f
C946 two_stage_opamp_dummy_magic_0.Vb1.n21 GNDA 0.216598f
C947 two_stage_opamp_dummy_magic_0.Vb1.t3 GNDA 0.012763f
C948 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA 0.080271f
C949 two_stage_opamp_dummy_magic_0.Vb1.n22 GNDA 0.113928f
C950 two_stage_opamp_dummy_magic_0.Vb1.n23 GNDA 0.949496f
C951 bgr_0.VB1_CUR_BIAS GNDA 0.847546f
C952 bgr_0.PFET_GATE_10uA.t23 GNDA 0.039433f
C953 bgr_0.PFET_GATE_10uA.t16 GNDA 0.058292f
C954 bgr_0.PFET_GATE_10uA.n0 GNDA 0.064232f
C955 bgr_0.PFET_GATE_10uA.t29 GNDA 0.039433f
C956 bgr_0.PFET_GATE_10uA.t17 GNDA 0.058292f
C957 bgr_0.PFET_GATE_10uA.n1 GNDA 0.064232f
C958 bgr_0.PFET_GATE_10uA.n2 GNDA 0.077289f
C959 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039433f
C960 bgr_0.PFET_GATE_10uA.t24 GNDA 0.058292f
C961 bgr_0.PFET_GATE_10uA.n3 GNDA 0.064232f
C962 bgr_0.PFET_GATE_10uA.t18 GNDA 0.039433f
C963 bgr_0.PFET_GATE_10uA.t25 GNDA 0.058292f
C964 bgr_0.PFET_GATE_10uA.n4 GNDA 0.064232f
C965 bgr_0.PFET_GATE_10uA.n5 GNDA 0.064438f
C966 bgr_0.PFET_GATE_10uA.t4 GNDA 0.786496f
C967 bgr_0.PFET_GATE_10uA.t8 GNDA 0.590788f
C968 bgr_0.PFET_GATE_10uA.t0 GNDA 0.040444f
C969 bgr_0.PFET_GATE_10uA.t7 GNDA 0.040444f
C970 bgr_0.PFET_GATE_10uA.n6 GNDA 0.103372f
C971 bgr_0.PFET_GATE_10uA.t9 GNDA 0.040444f
C972 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040444f
C973 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100701f
C974 bgr_0.PFET_GATE_10uA.n8 GNDA 0.984984f
C975 bgr_0.PFET_GATE_10uA.t1 GNDA 0.040444f
C976 bgr_0.PFET_GATE_10uA.t3 GNDA 0.040444f
C977 bgr_0.PFET_GATE_10uA.n9 GNDA 0.100701f
C978 bgr_0.PFET_GATE_10uA.n10 GNDA 0.558538f
C979 bgr_0.PFET_GATE_10uA.n11 GNDA 1.14022f
C980 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040444f
C981 bgr_0.PFET_GATE_10uA.t2 GNDA 0.040444f
C982 bgr_0.PFET_GATE_10uA.n12 GNDA 0.097542f
C983 bgr_0.PFET_GATE_10uA.n13 GNDA 0.358998f
C984 bgr_0.PFET_GATE_10uA.n14 GNDA 3.87496f
C985 bgr_0.PFET_GATE_10uA.t13 GNDA 0.045593f
C986 bgr_0.PFET_GATE_10uA.t21 GNDA 0.045593f
C987 bgr_0.PFET_GATE_10uA.n15 GNDA 0.138029f
C988 bgr_0.PFET_GATE_10uA.n16 GNDA 1.80019f
C989 bgr_0.PFET_GATE_10uA.n17 GNDA 1.42645f
C990 bgr_0.PFET_GATE_10uA.t27 GNDA 0.039433f
C991 bgr_0.PFET_GATE_10uA.t20 GNDA 0.039433f
C992 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039433f
C993 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039433f
C994 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039433f
C995 bgr_0.PFET_GATE_10uA.t11 GNDA 0.058292f
C996 bgr_0.PFET_GATE_10uA.n18 GNDA 0.07214f
C997 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051566f
C998 bgr_0.PFET_GATE_10uA.n20 GNDA 0.051566f
C999 bgr_0.PFET_GATE_10uA.n21 GNDA 0.051566f
C1000 bgr_0.PFET_GATE_10uA.n22 GNDA 0.043658f
C1001 bgr_0.PFET_GATE_10uA.t14 GNDA 0.039433f
C1002 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039433f
C1003 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039433f
C1004 bgr_0.PFET_GATE_10uA.t15 GNDA 0.058292f
C1005 bgr_0.PFET_GATE_10uA.n23 GNDA 0.07214f
C1006 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051566f
C1007 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043658f
C1008 bgr_0.PFET_GATE_10uA.n26 GNDA 0.059927f
C1009 VOUT+.t15 GNDA 0.043783f
C1010 VOUT+.t8 GNDA 0.043783f
C1011 VOUT+.n0 GNDA 0.174842f
C1012 VOUT+.t3 GNDA 0.043783f
C1013 VOUT+.t7 GNDA 0.043783f
C1014 VOUT+.n1 GNDA 0.17462f
C1015 VOUT+.n2 GNDA 0.193447f
C1016 VOUT+.t2 GNDA 0.043783f
C1017 VOUT+.t6 GNDA 0.043783f
C1018 VOUT+.n3 GNDA 0.17462f
C1019 VOUT+.n4 GNDA 0.101943f
C1020 VOUT+.t10 GNDA 0.043783f
C1021 VOUT+.t4 GNDA 0.043783f
C1022 VOUT+.n5 GNDA 0.17462f
C1023 VOUT+.n6 GNDA 0.101943f
C1024 VOUT+.t9 GNDA 0.043783f
C1025 VOUT+.t16 GNDA 0.043783f
C1026 VOUT+.n7 GNDA 0.174842f
C1027 VOUT+.n8 GNDA 0.123612f
C1028 VOUT+.t11 GNDA 0.043783f
C1029 VOUT+.t5 GNDA 0.043783f
C1030 VOUT+.n9 GNDA 0.17232f
C1031 VOUT+.n10 GNDA 0.32492f
C1032 VOUT+.t117 GNDA 0.296858f
C1033 VOUT+.t25 GNDA 0.291887f
C1034 VOUT+.n11 GNDA 0.1957f
C1035 VOUT+.t124 GNDA 0.291887f
C1036 VOUT+.n12 GNDA 0.1277f
C1037 VOUT+.t72 GNDA 0.296858f
C1038 VOUT+.t38 GNDA 0.291887f
C1039 VOUT+.n13 GNDA 0.1957f
C1040 VOUT+.t127 GNDA 0.291887f
C1041 VOUT+.t34 GNDA 0.296236f
C1042 VOUT+.t86 GNDA 0.296236f
C1043 VOUT+.t42 GNDA 0.296236f
C1044 VOUT+.t96 GNDA 0.296236f
C1045 VOUT+.t143 GNDA 0.296236f
C1046 VOUT+.t106 GNDA 0.296236f
C1047 VOUT+.t154 GNDA 0.296236f
C1048 VOUT+.t64 GNDA 0.296236f
C1049 VOUT+.t116 GNDA 0.296236f
C1050 VOUT+.t73 GNDA 0.296236f
C1051 VOUT+.t149 GNDA 0.291887f
C1052 VOUT+.n14 GNDA 0.196323f
C1053 VOUT+.t58 GNDA 0.291887f
C1054 VOUT+.n15 GNDA 0.251052f
C1055 VOUT+.t97 GNDA 0.291887f
C1056 VOUT+.n16 GNDA 0.251052f
C1057 VOUT+.t131 GNDA 0.291887f
C1058 VOUT+.n17 GNDA 0.251052f
C1059 VOUT+.t24 GNDA 0.291887f
C1060 VOUT+.n18 GNDA 0.251052f
C1061 VOUT+.t75 GNDA 0.291887f
C1062 VOUT+.n19 GNDA 0.251052f
C1063 VOUT+.t113 GNDA 0.291887f
C1064 VOUT+.n20 GNDA 0.251052f
C1065 VOUT+.t144 GNDA 0.291887f
C1066 VOUT+.n21 GNDA 0.251052f
C1067 VOUT+.t54 GNDA 0.291887f
C1068 VOUT+.n22 GNDA 0.251052f
C1069 VOUT+.t94 GNDA 0.291887f
C1070 VOUT+.n23 GNDA 0.251052f
C1071 VOUT+.n24 GNDA 0.237158f
C1072 VOUT+.t37 GNDA 0.296858f
C1073 VOUT+.t142 GNDA 0.291887f
C1074 VOUT+.n25 GNDA 0.1957f
C1075 VOUT+.t93 GNDA 0.291887f
C1076 VOUT+.t20 GNDA 0.296858f
C1077 VOUT+.t57 GNDA 0.291887f
C1078 VOUT+.n26 GNDA 0.1957f
C1079 VOUT+.n27 GNDA 0.237158f
C1080 VOUT+.t79 GNDA 0.296858f
C1081 VOUT+.t41 GNDA 0.291887f
C1082 VOUT+.n28 GNDA 0.1957f
C1083 VOUT+.t133 GNDA 0.291887f
C1084 VOUT+.t60 GNDA 0.296858f
C1085 VOUT+.t100 GNDA 0.291887f
C1086 VOUT+.n29 GNDA 0.1957f
C1087 VOUT+.n30 GNDA 0.237158f
C1088 VOUT+.t121 GNDA 0.296858f
C1089 VOUT+.t83 GNDA 0.291887f
C1090 VOUT+.n31 GNDA 0.1957f
C1091 VOUT+.t31 GNDA 0.291887f
C1092 VOUT+.t104 GNDA 0.296858f
C1093 VOUT+.t137 GNDA 0.291887f
C1094 VOUT+.n32 GNDA 0.1957f
C1095 VOUT+.n33 GNDA 0.237158f
C1096 VOUT+.t84 GNDA 0.296858f
C1097 VOUT+.t49 GNDA 0.291887f
C1098 VOUT+.n34 GNDA 0.1957f
C1099 VOUT+.t138 GNDA 0.291887f
C1100 VOUT+.t66 GNDA 0.296858f
C1101 VOUT+.t103 GNDA 0.291887f
C1102 VOUT+.n35 GNDA 0.1957f
C1103 VOUT+.n36 GNDA 0.237158f
C1104 VOUT+.t108 GNDA 0.296858f
C1105 VOUT+.t69 GNDA 0.291887f
C1106 VOUT+.n37 GNDA 0.1957f
C1107 VOUT+.t90 GNDA 0.291887f
C1108 VOUT+.n38 GNDA 0.1277f
C1109 VOUT+.t67 GNDA 0.296858f
C1110 VOUT+.t30 GNDA 0.291887f
C1111 VOUT+.n39 GNDA 0.1957f
C1112 VOUT+.t51 GNDA 0.291887f
C1113 VOUT+.t53 GNDA 0.296236f
C1114 VOUT+.t156 GNDA 0.296236f
C1115 VOUT+.t44 GNDA 0.296858f
C1116 VOUT+.t136 GNDA 0.291887f
C1117 VOUT+.n40 GNDA 0.1957f
C1118 VOUT+.t101 GNDA 0.291887f
C1119 VOUT+.n41 GNDA 0.12314f
C1120 VOUT+.t36 GNDA 0.296236f
C1121 VOUT+.t151 GNDA 0.296858f
C1122 VOUT+.t98 GNDA 0.291887f
C1123 VOUT+.n42 GNDA 0.1957f
C1124 VOUT+.t59 GNDA 0.291887f
C1125 VOUT+.n43 GNDA 0.12314f
C1126 VOUT+.t140 GNDA 0.296236f
C1127 VOUT+.t118 GNDA 0.296858f
C1128 VOUT+.t56 GNDA 0.291887f
C1129 VOUT+.n44 GNDA 0.1957f
C1130 VOUT+.t21 GNDA 0.291887f
C1131 VOUT+.n45 GNDA 0.12314f
C1132 VOUT+.t105 GNDA 0.296236f
C1133 VOUT+.t65 GNDA 0.296858f
C1134 VOUT+.t80 GNDA 0.291887f
C1135 VOUT+.n46 GNDA 0.1957f
C1136 VOUT+.t43 GNDA 0.291887f
C1137 VOUT+.n47 GNDA 0.12314f
C1138 VOUT+.t125 GNDA 0.296236f
C1139 VOUT+.t145 GNDA 0.29648f
C1140 VOUT+.t87 GNDA 0.296236f
C1141 VOUT+.t110 GNDA 0.29648f
C1142 VOUT+.t50 GNDA 0.296236f
C1143 VOUT+.t70 GNDA 0.29648f
C1144 VOUT+.t150 GNDA 0.296236f
C1145 VOUT+.t95 GNDA 0.29648f
C1146 VOUT+.t32 GNDA 0.296236f
C1147 VOUT+.t134 GNDA 0.291887f
C1148 VOUT+.n48 GNDA 0.323078f
C1149 VOUT+.t111 GNDA 0.291887f
C1150 VOUT+.n49 GNDA 0.377807f
C1151 VOUT+.t147 GNDA 0.291887f
C1152 VOUT+.n50 GNDA 0.377807f
C1153 VOUT+.t45 GNDA 0.291887f
C1154 VOUT+.n51 GNDA 0.377807f
C1155 VOUT+.t85 GNDA 0.291887f
C1156 VOUT+.n52 GNDA 0.310341f
C1157 VOUT+.t61 GNDA 0.291887f
C1158 VOUT+.n53 GNDA 0.310341f
C1159 VOUT+.t102 GNDA 0.291887f
C1160 VOUT+.n54 GNDA 0.310341f
C1161 VOUT+.t139 GNDA 0.291887f
C1162 VOUT+.n55 GNDA 0.310341f
C1163 VOUT+.t119 GNDA 0.291887f
C1164 VOUT+.n56 GNDA 0.251052f
C1165 VOUT+.t155 GNDA 0.291887f
C1166 VOUT+.n57 GNDA 0.251052f
C1167 VOUT+.n58 GNDA 0.237158f
C1168 VOUT+.t27 GNDA 0.296858f
C1169 VOUT+.t130 GNDA 0.291887f
C1170 VOUT+.n59 GNDA 0.1957f
C1171 VOUT+.t152 GNDA 0.291887f
C1172 VOUT+.t76 GNDA 0.296858f
C1173 VOUT+.t115 GNDA 0.291887f
C1174 VOUT+.n60 GNDA 0.1957f
C1175 VOUT+.n61 GNDA 0.237158f
C1176 VOUT+.t62 GNDA 0.296858f
C1177 VOUT+.t23 GNDA 0.291887f
C1178 VOUT+.n62 GNDA 0.1957f
C1179 VOUT+.t47 GNDA 0.291887f
C1180 VOUT+.t112 GNDA 0.296858f
C1181 VOUT+.t148 GNDA 0.291887f
C1182 VOUT+.n63 GNDA 0.1957f
C1183 VOUT+.n64 GNDA 0.237158f
C1184 VOUT+.t114 GNDA 0.296858f
C1185 VOUT+.t78 GNDA 0.291887f
C1186 VOUT+.n65 GNDA 0.1957f
C1187 VOUT+.t26 GNDA 0.291887f
C1188 VOUT+.t99 GNDA 0.296858f
C1189 VOUT+.t132 GNDA 0.291887f
C1190 VOUT+.n66 GNDA 0.1957f
C1191 VOUT+.n67 GNDA 0.237158f
C1192 VOUT+.t74 GNDA 0.296858f
C1193 VOUT+.t39 GNDA 0.291887f
C1194 VOUT+.n68 GNDA 0.1957f
C1195 VOUT+.t128 GNDA 0.291887f
C1196 VOUT+.t55 GNDA 0.296858f
C1197 VOUT+.t92 GNDA 0.291887f
C1198 VOUT+.n69 GNDA 0.1957f
C1199 VOUT+.n70 GNDA 0.237158f
C1200 VOUT+.t109 GNDA 0.296858f
C1201 VOUT+.t71 GNDA 0.291887f
C1202 VOUT+.n71 GNDA 0.1957f
C1203 VOUT+.t19 GNDA 0.291887f
C1204 VOUT+.t91 GNDA 0.296858f
C1205 VOUT+.t126 GNDA 0.291887f
C1206 VOUT+.n72 GNDA 0.1957f
C1207 VOUT+.n73 GNDA 0.237158f
C1208 VOUT+.t68 GNDA 0.296858f
C1209 VOUT+.t33 GNDA 0.291887f
C1210 VOUT+.n74 GNDA 0.1957f
C1211 VOUT+.t122 GNDA 0.291887f
C1212 VOUT+.t52 GNDA 0.296858f
C1213 VOUT+.t88 GNDA 0.291887f
C1214 VOUT+.n75 GNDA 0.1957f
C1215 VOUT+.n76 GNDA 0.237158f
C1216 VOUT+.t29 GNDA 0.296858f
C1217 VOUT+.t135 GNDA 0.291887f
C1218 VOUT+.n77 GNDA 0.1957f
C1219 VOUT+.t82 GNDA 0.291887f
C1220 VOUT+.t153 GNDA 0.296858f
C1221 VOUT+.t48 GNDA 0.291887f
C1222 VOUT+.n78 GNDA 0.1957f
C1223 VOUT+.n79 GNDA 0.237158f
C1224 VOUT+.t63 GNDA 0.296858f
C1225 VOUT+.t28 GNDA 0.291887f
C1226 VOUT+.n80 GNDA 0.1957f
C1227 VOUT+.t120 GNDA 0.291887f
C1228 VOUT+.t46 GNDA 0.296858f
C1229 VOUT+.t81 GNDA 0.291887f
C1230 VOUT+.n81 GNDA 0.1957f
C1231 VOUT+.n82 GNDA 0.237158f
C1232 VOUT+.t22 GNDA 0.296858f
C1233 VOUT+.t129 GNDA 0.291887f
C1234 VOUT+.n83 GNDA 0.1957f
C1235 VOUT+.t77 GNDA 0.291887f
C1236 VOUT+.t146 GNDA 0.296858f
C1237 VOUT+.t40 GNDA 0.291887f
C1238 VOUT+.n84 GNDA 0.1957f
C1239 VOUT+.n85 GNDA 0.237158f
C1240 VOUT+.t123 GNDA 0.296858f
C1241 VOUT+.t89 GNDA 0.291887f
C1242 VOUT+.n86 GNDA 0.1957f
C1243 VOUT+.t35 GNDA 0.291887f
C1244 VOUT+.n87 GNDA 0.237158f
C1245 VOUT+.t141 GNDA 0.291887f
C1246 VOUT+.n88 GNDA 0.1277f
C1247 VOUT+.t107 GNDA 0.291887f
C1248 VOUT+.n89 GNDA 0.232121f
C1249 VOUT+.n90 GNDA 0.521129f
C1250 VOUT+.t1 GNDA 0.05108f
C1251 VOUT+.t18 GNDA 0.05108f
C1252 VOUT+.n91 GNDA 0.235555f
C1253 VOUT+.t12 GNDA 0.05108f
C1254 VOUT+.t0 GNDA 0.05108f
C1255 VOUT+.n92 GNDA 0.234998f
C1256 VOUT+.n93 GNDA 0.184732f
C1257 VOUT+.t17 GNDA 0.05108f
C1258 VOUT+.t13 GNDA 0.05108f
C1259 VOUT+.n94 GNDA 0.234998f
C1260 VOUT+.n95 GNDA 0.125481f
C1261 VOUT+.t14 GNDA 0.084549f
C1262 VOUT+.n96 GNDA 0.179426f
C1263 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.023034f
C1264 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.023034f
C1265 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.076867f
C1266 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.023034f
C1267 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.023034f
C1268 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.082819f
C1269 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.023034f
C1270 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.023034f
C1271 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.082819f
C1272 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.023034f
C1273 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.023034f
C1274 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.082024f
C1275 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.321952f
C1276 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.023034f
C1277 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.023034f
C1278 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.082024f
C1279 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.166748f
C1280 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.023034f
C1281 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.023034f
C1282 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.082024f
C1283 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.166748f
C1284 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.201273f
C1285 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.199546f
C1286 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.734081f
C1287 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.101352f
C1288 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.101352f
C1289 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.107946f
C1290 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.085543f
C1291 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.04573f
C1292 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.101352f
C1293 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.101352f
C1294 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.101352f
C1295 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.101352f
C1296 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.101352f
C1297 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.101352f
C1298 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.107946f
C1299 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.085543f
C1300 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.048372f
C1301 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.048372f
C1302 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.048372f
C1303 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.048372f
C1304 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.04573f
C1305 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.025502f
C1306 two_stage_opamp_dummy_magic_0.X.n20 GNDA 1.2196f
C1307 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.053747f
C1308 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.053747f
C1309 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.184971f
C1310 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.053747f
C1311 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.053747f
C1312 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.184521f
C1313 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.398323f
C1314 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.053747f
C1315 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.053747f
C1316 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.184521f
C1317 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.211671f
C1318 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.053747f
C1319 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.053747f
C1320 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.184521f
C1321 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.211671f
C1322 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.053747f
C1323 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.053747f
C1324 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.184521f
C1325 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.257031f
C1326 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.053747f
C1327 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.053747f
C1328 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.180411f
C1329 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.513007f
C1330 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.032248f
C1331 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.032248f
C1332 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.032248f
C1333 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.032248f
C1334 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.032248f
C1335 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.032248f
C1336 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.032248f
C1337 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.039159f
C1338 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.039159f
C1339 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.025338f
C1340 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.025338f
C1341 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.025338f
C1342 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.025338f
C1343 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.025338f
C1344 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.022696f
C1345 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.032248f
C1346 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.039159f
C1347 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.036516f
C1348 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.022278f
C1349 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.0668f
C1350 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.0668f
C1351 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.0668f
C1352 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.0668f
C1353 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.0668f
C1354 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.0668f
C1355 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.0668f
C1356 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.073493f
C1357 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.06241f
C1358 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.036855f
C1359 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.036855f
C1360 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.036855f
C1361 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.036855f
C1362 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.036855f
C1363 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.034213f
C1364 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.0668f
C1365 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.073493f
C1366 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.059768f
C1367 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.022245f
C1368 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.314383f
C1369 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.941608f
C1370 two_stage_opamp_dummy_magic_0.X.n52 GNDA 0.451014f
C1371 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.026504f
C1372 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.026504f
C1373 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.091215f
C1374 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.026504f
C1375 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.026504f
C1376 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.090993f
C1377 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.196425f
C1378 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.073525f
C1379 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.102604f
C1380 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.130751f
C1381 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.046153f
C1382 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.086435f
C1383 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.0577f
C1384 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.130751f
C1385 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.046153f
C1386 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.086435f
C1387 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.0577f
C1388 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.052251f
C1389 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.102604f
C1390 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.305777f
C1391 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.456416f
C1392 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.263528f
C1393 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.263528f
C1394 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.263528f
C1395 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.263528f
C1396 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.197646f
C1397 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.131764f
C1398 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.197646f
C1399 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.263528f
C1400 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.263528f
C1401 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.263528f
C1402 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.263528f
C1403 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.456416f
C1404 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.305777f
C1405 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.073525f
C1406 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.110185f
C1407 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.026504f
C1408 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.026504f
C1409 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.088966f
C1410 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.076058f
C1411 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.036349f
C1412 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.026504f
C1413 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.026504f
C1414 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.090993f
C1415 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.104381f
C1416 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.026504f
C1417 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.026504f
C1418 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.090993f
C1419 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.158094f
C1420 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.026504f
C1421 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.026504f
C1422 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.091215f
C1423 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.026504f
C1424 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.026504f
C1425 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.090993f
C1426 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.196424f
C1427 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.026504f
C1428 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.026504f
C1429 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.090993f
C1430 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.104381f
C1431 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.026504f
C1432 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.026504f
C1433 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.090993f
C1434 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.104381f
C1435 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.026504f
C1436 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.026504f
C1437 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.090993f
C1438 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.104381f
C1439 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.026504f
C1440 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.026504f
C1441 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.090993f
C1442 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.180564f
C1443 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.016652f
C1444 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.016652f
C1445 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.035974f
C1446 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.053205f
C1447 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.261863f
C1448 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.137379f
C1449 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.137379f
C1450 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.137379f
C1451 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.137379f
C1452 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.158535f
C1453 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.128713f
C1454 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.079097f
C1455 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.079097f
C1456 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.075701f
C1457 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.137379f
C1458 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.137379f
C1459 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.137379f
C1460 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.137379f
C1461 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.158535f
C1462 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.128713f
C1463 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.079097f
C1464 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.079097f
C1465 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.075701f
C1466 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.051501f
C1467 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.137379f
C1468 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.137379f
C1469 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.137379f
C1470 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.137379f
C1471 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.158535f
C1472 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.128713f
C1473 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.079097f
C1474 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.079097f
C1475 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.075701f
C1476 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.137379f
C1477 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.137379f
C1478 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.137379f
C1479 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.137379f
C1480 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.158535f
C1481 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.128713f
C1482 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.079097f
C1483 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.079097f
C1484 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.075701f
C1485 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.050681f
C1486 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 1.85691f
C1487 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 1.54451f
C1488 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.166013f
C1489 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 7.99036f
C1490 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.027753f
C1491 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.027753f
C1492 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.083827f
C1493 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.027753f
C1494 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.027753f
C1495 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.089396f
C1496 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.027753f
C1497 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.027753f
C1498 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.089396f
C1499 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.027753f
C1500 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.027753f
C1501 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.088568f
C1502 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.429835f
C1503 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.28805f
C1504 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.260315f
C1505 bgr_0.VB2_CUR_BIAS GNDA 8.02162f
C1506 bgr_0.V_mir2.t1 GNDA 0.017685f
C1507 bgr_0.V_mir2.t0 GNDA 0.017685f
C1508 bgr_0.V_mir2.n0 GNDA 0.046242f
C1509 bgr_0.V_mir2.t4 GNDA 0.075466f
C1510 bgr_0.V_mir2.t3 GNDA 0.017685f
C1511 bgr_0.V_mir2.t2 GNDA 0.017685f
C1512 bgr_0.V_mir2.n1 GNDA 0.050199f
C1513 bgr_0.V_mir2.n2 GNDA 0.827814f
C1514 bgr_0.V_mir2.n3 GNDA 0.268286f
C1515 bgr_0.V_mir2.t5 GNDA 0.042444f
C1516 bgr_0.V_mir2.t18 GNDA 0.042444f
C1517 bgr_0.V_mir2.t20 GNDA 0.06851f
C1518 bgr_0.V_mir2.n4 GNDA 0.076506f
C1519 bgr_0.V_mir2.n5 GNDA 0.052264f
C1520 bgr_0.V_mir2.t9 GNDA 0.053881f
C1521 bgr_0.V_mir2.n6 GNDA 0.081315f
C1522 bgr_0.V_mir2.t6 GNDA 0.03537f
C1523 bgr_0.V_mir2.t10 GNDA 0.03537f
C1524 bgr_0.V_mir2.n7 GNDA 0.08097f
C1525 bgr_0.V_mir2.n8 GNDA 0.201563f
C1526 bgr_0.V_mir2.t15 GNDA 0.042444f
C1527 bgr_0.V_mir2.t21 GNDA 0.042444f
C1528 bgr_0.V_mir2.t17 GNDA 0.06851f
C1529 bgr_0.V_mir2.n9 GNDA 0.076506f
C1530 bgr_0.V_mir2.n10 GNDA 0.052264f
C1531 bgr_0.V_mir2.t7 GNDA 0.053881f
C1532 bgr_0.V_mir2.n11 GNDA 0.081315f
C1533 bgr_0.V_mir2.t16 GNDA 0.03537f
C1534 bgr_0.V_mir2.t8 GNDA 0.03537f
C1535 bgr_0.V_mir2.n12 GNDA 0.08097f
C1536 bgr_0.V_mir2.n13 GNDA 0.203577f
C1537 bgr_0.V_mir2.n14 GNDA 0.699157f
C1538 bgr_0.V_mir2.n15 GNDA 0.09373f
C1539 bgr_0.V_mir2.t13 GNDA 0.042444f
C1540 bgr_0.V_mir2.t19 GNDA 0.042444f
C1541 bgr_0.V_mir2.t22 GNDA 0.06851f
C1542 bgr_0.V_mir2.n16 GNDA 0.076506f
C1543 bgr_0.V_mir2.n17 GNDA 0.052264f
C1544 bgr_0.V_mir2.t11 GNDA 0.053881f
C1545 bgr_0.V_mir2.n18 GNDA 0.081315f
C1546 bgr_0.V_mir2.n19 GNDA 0.156007f
C1547 bgr_0.V_mir2.t12 GNDA 0.03537f
C1548 bgr_0.V_mir2.n20 GNDA 0.08097f
C1549 bgr_0.V_mir2.t14 GNDA 0.03537f
C1550 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.36379f
C1551 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 11.624901f
C1552 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.018358f
C1553 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.018358f
C1554 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.042939f
C1555 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.018358f
C1556 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.018358f
C1557 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.042615f
C1558 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.018358f
C1559 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.018358f
C1560 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.042642f
C1561 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.015145f
C1562 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.015145f
C1563 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.015145f
C1564 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.015145f
C1565 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.015145f
C1566 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.015145f
C1567 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.015145f
C1568 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.015145f
C1569 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.015145f
C1570 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.015145f
C1571 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.015145f
C1572 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.015145f
C1573 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.015145f
C1574 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.015145f
C1575 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.015145f
C1576 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.015145f
C1577 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.032814f
C1578 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.051172f
C1579 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.039928f
C1580 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.039928f
C1581 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.039928f
C1582 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.039928f
C1583 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.039928f
C1584 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.039928f
C1585 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.039928f
C1586 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.039928f
C1587 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.039928f
C1588 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.039928f
C1589 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.039928f
C1590 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.039928f
C1591 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.039928f
C1592 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.039928f
C1593 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.034167f
C1594 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.015145f
C1595 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.015145f
C1596 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.032814f
C1597 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.051172f
C1598 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.034167f
C1599 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.054821f
C1600 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.018358f
C1601 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.018358f
C1602 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.036715f
C1603 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.116293f
C1604 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.018358f
C1605 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.018358f
C1606 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.042642f
C1607 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.018358f
C1608 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.018358f
C1609 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.042301f
C1610 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.036715f
C1611 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.036715f
C1612 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.112441f
C1613 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.065343f
C1614 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.024434f
C1615 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.076638f
C1616 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.024434f
C1617 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.062736f
C1618 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.024434f
C1619 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.062736f
C1620 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.024434f
C1621 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.096248f
C1622 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.623974f
C1623 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.079245f
C1624 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.079245f
C1625 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.265552f
C1626 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 2.99217f
C1627 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.079245f
C1628 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.079245f
C1629 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.265552f
C1630 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.717088f
C1631 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.079245f
C1632 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.079245f
C1633 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.265552f
C1634 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 1.0252f
C1635 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 1.01347f
C1636 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.038072f
C1637 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.011995f
C1638 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.022383f
C1639 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.053439f
C1640 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.44626f
C1641 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.011995f
C1642 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.022383f
C1643 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.053439f
C1644 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.509955f
C1645 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.037821f
C1646 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.481763f
C1647 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.011995f
C1648 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.022383f
C1649 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.053439f
C1650 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.26588f
C1651 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.011995f
C1652 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.022383f
C1653 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.053439f
C1654 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.363087f
C1655 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.02389f
C1656 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.02389f
C1657 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.059804f
C1658 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.02389f
C1659 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.02389f
C1660 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.059594f
C1661 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.453962f
C1662 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.02389f
C1663 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.02389f
C1664 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.059594f
C1665 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.673829f
C1666 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 3.27646f
C1667 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.305094f
C1668 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.04778f
C1669 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.04778f
C1670 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.13851f
C1671 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.04778f
C1672 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.04778f
C1673 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.138073f
C1674 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.545233f
C1675 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.04778f
C1676 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.04778f
C1677 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.138073f
C1678 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.289558f
C1679 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.04778f
C1680 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.04778f
C1681 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.138073f
C1682 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.289558f
C1683 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.04778f
C1684 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.04778f
C1685 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.138073f
C1686 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 0.522724f
C1687 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 GNDA 1.02833f
C1688 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.022266f
C1689 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.022266f
C1690 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.074304f
C1691 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.022266f
C1692 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.022266f
C1693 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.079792f
C1694 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.022266f
C1695 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.022266f
C1696 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.079289f
C1697 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.342655f
C1698 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.022266f
C1699 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.022266f
C1700 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.079289f
C1701 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.18197f
C1702 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.022266f
C1703 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.022266f
C1704 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.079289f
C1705 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.18197f
C1706 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.022266f
C1707 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.022266f
C1708 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.079792f
C1709 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.226f
C1710 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.313311f
C1711 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.051955f
C1712 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.051955f
C1713 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.178804f
C1714 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.051955f
C1715 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.051955f
C1716 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.178369f
C1717 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.385041f
C1718 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.051955f
C1719 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.051955f
C1720 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.178369f
C1721 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.204613f
C1722 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.051955f
C1723 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.051955f
C1724 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.178369f
C1725 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.204613f
C1726 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.051955f
C1727 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.051955f
C1728 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.178369f
C1729 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.248461f
C1730 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.051955f
C1731 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.051955f
C1732 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.174395f
C1733 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.497474f
C1734 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.031173f
C1735 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.037853f
C1736 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.035299f
C1737 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.031173f
C1738 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.031173f
C1739 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.031173f
C1740 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.031173f
C1741 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.031173f
C1742 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.031173f
C1743 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.031173f
C1744 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.037853f
C1745 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.037853f
C1746 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.024493f
C1747 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.024493f
C1748 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.024493f
C1749 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.024493f
C1750 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.024493f
C1751 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.021939f
C1752 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.021535f
C1753 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.064573f
C1754 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.071042f
C1755 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.057775f
C1756 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.064573f
C1757 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.064573f
C1758 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.064573f
C1759 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.064573f
C1760 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.064573f
C1761 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.064573f
C1762 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.064573f
C1763 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.071042f
C1764 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.060329f
C1765 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.035626f
C1766 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.035626f
C1767 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.035626f
C1768 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.035626f
C1769 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.035626f
C1770 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.033072f
C1771 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.021503f
C1772 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.301806f
C1773 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.910287f
C1774 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.454055f
C1775 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.097972f
C1776 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.097972f
C1777 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.097972f
C1778 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.097972f
C1779 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.097972f
C1780 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.097972f
C1781 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.104347f
C1782 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.082691f
C1783 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.046759f
C1784 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.046759f
C1785 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.046759f
C1786 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.046759f
C1787 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.044205f
C1788 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.097972f
C1789 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.097972f
C1790 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.104347f
C1791 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.082691f
C1792 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 0.044205f
C1793 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.024652f
C1794 two_stage_opamp_dummy_magic_0.Y.n52 GNDA 1.17745f
C1795 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.709602f
C1796 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.015165f
C1797 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.015129f
C1798 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.404283f
C1799 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.015129f
C1800 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.01672f
C1801 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.06287f
C1802 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 0.017939f
C1803 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 1.57415f
C1804 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.017939f
C1805 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.229687f
C1806 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.205215f
C1807 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.360369f
C1808 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.361571f
C1809 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.194207f
C1810 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.207375f
C1811 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.360369f
C1812 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.361571f
C1813 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.194207f
C1814 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.226779f
C1815 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.360369f
C1816 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.361571f
C1817 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.194207f
C1818 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.226779f
C1819 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.360369f
C1820 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.361571f
C1821 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.194207f
C1822 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.226779f
C1823 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.360369f
C1824 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.361571f
C1825 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.380975f
C1826 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.380975f
C1827 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.194207f
C1828 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.226779f
C1829 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.360369f
C1830 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.361571f
C1831 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.380975f
C1832 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.380975f
C1833 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.194207f
C1834 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.226779f
C1835 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.361571f
C1836 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.362881f
C1837 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.361571f
C1838 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.364405f
C1839 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.396343f
C1840 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.361571f
C1841 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.362881f
C1842 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.361571f
C1843 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.362881f
C1844 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.361571f
C1845 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.362881f
C1846 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.361571f
C1847 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.362881f
C1848 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.361571f
C1849 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.362881f
C1850 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.361571f
C1851 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.362881f
C1852 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.361571f
C1853 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.362881f
C1854 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.361571f
C1855 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.362881f
C1856 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.361571f
C1857 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.362881f
C1858 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.361571f
C1859 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.362881f
C1860 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.361571f
C1861 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.362881f
C1862 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.361571f
C1863 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.362881f
C1864 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.361571f
C1865 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.362881f
C1866 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.361571f
C1867 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.362881f
C1868 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.361571f
C1869 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.362881f
C1870 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.361571f
C1871 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.362881f
C1872 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.361571f
C1873 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.362881f
C1874 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.361571f
C1875 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.362881f
C1876 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.361571f
C1877 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.362881f
C1878 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.361571f
C1879 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.362881f
C1880 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.361571f
C1881 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.362881f
C1882 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.361571f
C1883 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.362881f
C1884 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.361571f
C1885 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.362881f
C1886 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.361571f
C1887 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.362881f
C1888 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.361571f
C1889 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.362881f
C1890 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.361571f
C1891 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.362881f
C1892 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.361571f
C1893 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.362881f
C1894 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.361571f
C1895 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.362881f
C1896 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.361571f
C1897 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.379298f
C1898 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.361571f
C1899 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.194207f
C1900 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.207849f
C1901 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.361571f
C1902 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.194207f
C1903 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.206173f
C1904 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.361571f
C1905 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.194207f
C1906 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.206173f
C1907 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.361571f
C1908 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.194207f
C1909 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.206173f
C1910 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.361571f
C1911 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.194207f
C1912 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.206173f
C1913 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.361571f
C1914 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.194207f
C1915 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.206173f
C1916 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.361571f
C1917 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.194207f
C1918 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.206173f
C1919 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.361571f
C1920 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.194207f
C1921 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.206173f
C1922 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.361571f
C1923 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.194207f
C1924 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.206173f
C1925 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.361571f
C1926 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.362881f
C1927 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.361571f
C1928 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.362881f
C1929 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.174802f
C1930 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.225469f
C1931 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.193005f
C1932 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.244873f
C1933 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.193005f
C1934 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.262967f
C1935 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.193005f
C1936 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.262967f
C1937 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.193005f
C1938 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.262967f
C1939 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.193005f
C1940 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.262967f
C1941 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.193005f
C1942 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.262967f
C1943 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.193005f
C1944 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.262967f
C1945 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.193005f
C1946 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.262967f
C1947 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.193005f
C1948 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.262967f
C1949 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.193005f
C1950 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.262967f
C1951 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.193005f
C1952 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.262967f
C1953 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.193005f
C1954 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.262967f
C1955 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.193005f
C1956 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.262967f
C1957 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.193005f
C1958 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.262967f
C1959 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.193005f
C1960 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.262967f
C1961 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.193005f
C1962 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.244873f
C1963 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.360369f
C1964 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.174802f
C1965 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.226779f
C1966 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.360369f
C1967 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.174802f
C1968 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.226779f
C1969 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.360369f
C1970 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.361571f
C1971 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.380975f
C1972 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.380975f
C1973 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.194207f
C1974 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.226779f
C1975 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.360369f
C1976 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.226779f
C1977 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.194207f
C1978 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.380975f
C1979 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.380975f
C1980 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.455833f
C1981 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.312131f
C1982 VOUT-.t17 GNDA 0.051122f
C1983 VOUT-.t6 GNDA 0.051122f
C1984 VOUT-.n0 GNDA 0.235747f
C1985 VOUT-.t3 GNDA 0.051122f
C1986 VOUT-.t1 GNDA 0.051122f
C1987 VOUT-.n1 GNDA 0.23519f
C1988 VOUT-.n2 GNDA 0.184883f
C1989 VOUT-.t18 GNDA 0.051122f
C1990 VOUT-.t16 GNDA 0.051122f
C1991 VOUT-.n3 GNDA 0.23519f
C1992 VOUT-.n4 GNDA 0.125584f
C1993 VOUT-.t4 GNDA 0.084618f
C1994 VOUT-.n5 GNDA 0.179572f
C1995 VOUT-.t14 GNDA 0.043819f
C1996 VOUT-.t10 GNDA 0.043819f
C1997 VOUT-.n6 GNDA 0.175106f
C1998 VOUT-.t13 GNDA 0.043819f
C1999 VOUT-.t15 GNDA 0.043819f
C2000 VOUT-.n7 GNDA 0.175106f
C2001 VOUT-.t0 GNDA 0.043819f
C2002 VOUT-.t9 GNDA 0.043819f
C2003 VOUT-.n8 GNDA 0.174762f
C2004 VOUT-.n9 GNDA 0.178148f
C2005 VOUT-.t2 GNDA 0.043819f
C2006 VOUT-.t11 GNDA 0.043819f
C2007 VOUT-.n10 GNDA 0.174762f
C2008 VOUT-.n11 GNDA 0.091802f
C2009 VOUT-.t7 GNDA 0.043819f
C2010 VOUT-.t12 GNDA 0.043819f
C2011 VOUT-.n12 GNDA 0.174762f
C2012 VOUT-.n13 GNDA 0.091802f
C2013 VOUT-.n14 GNDA 0.108255f
C2014 VOUT-.t5 GNDA 0.043819f
C2015 VOUT-.t8 GNDA 0.043819f
C2016 VOUT-.n15 GNDA 0.172461f
C2017 VOUT-.n16 GNDA 0.325185f
C2018 VOUT-.t101 GNDA 0.292125f
C2019 VOUT-.t108 GNDA 0.297101f
C2020 VOUT-.t149 GNDA 0.292125f
C2021 VOUT-.n17 GNDA 0.19586f
C2022 VOUT-.n18 GNDA 0.127805f
C2023 VOUT-.t48 GNDA 0.296478f
C2024 VOUT-.t92 GNDA 0.296478f
C2025 VOUT-.t42 GNDA 0.296478f
C2026 VOUT-.t130 GNDA 0.296478f
C2027 VOUT-.t84 GNDA 0.296478f
C2028 VOUT-.t125 GNDA 0.296478f
C2029 VOUT-.t74 GNDA 0.296478f
C2030 VOUT-.t23 GNDA 0.296478f
C2031 VOUT-.t64 GNDA 0.296478f
C2032 VOUT-.t150 GNDA 0.296478f
C2033 VOUT-.t88 GNDA 0.292125f
C2034 VOUT-.n19 GNDA 0.196483f
C2035 VOUT-.t51 GNDA 0.292125f
C2036 VOUT-.n20 GNDA 0.251257f
C2037 VOUT-.t137 GNDA 0.292125f
C2038 VOUT-.n21 GNDA 0.251257f
C2039 VOUT-.t106 GNDA 0.292125f
C2040 VOUT-.n22 GNDA 0.251257f
C2041 VOUT-.t75 GNDA 0.292125f
C2042 VOUT-.n23 GNDA 0.251257f
C2043 VOUT-.t25 GNDA 0.292125f
C2044 VOUT-.n24 GNDA 0.251257f
C2045 VOUT-.t128 GNDA 0.292125f
C2046 VOUT-.n25 GNDA 0.251257f
C2047 VOUT-.t90 GNDA 0.292125f
C2048 VOUT-.n26 GNDA 0.251257f
C2049 VOUT-.t54 GNDA 0.292125f
C2050 VOUT-.n27 GNDA 0.251257f
C2051 VOUT-.t140 GNDA 0.292125f
C2052 VOUT-.n28 GNDA 0.251257f
C2053 VOUT-.t110 GNDA 0.292125f
C2054 VOUT-.t28 GNDA 0.297101f
C2055 VOUT-.t79 GNDA 0.292125f
C2056 VOUT-.n29 GNDA 0.19586f
C2057 VOUT-.n30 GNDA 0.237352f
C2058 VOUT-.t24 GNDA 0.297101f
C2059 VOUT-.t113 GNDA 0.292125f
C2060 VOUT-.n31 GNDA 0.19586f
C2061 VOUT-.t78 GNDA 0.292125f
C2062 VOUT-.t129 GNDA 0.297101f
C2063 VOUT-.t38 GNDA 0.292125f
C2064 VOUT-.n32 GNDA 0.19586f
C2065 VOUT-.n33 GNDA 0.237352f
C2066 VOUT-.t61 GNDA 0.297101f
C2067 VOUT-.t147 GNDA 0.292125f
C2068 VOUT-.n34 GNDA 0.19586f
C2069 VOUT-.t117 GNDA 0.292125f
C2070 VOUT-.t32 GNDA 0.297101f
C2071 VOUT-.t83 GNDA 0.292125f
C2072 VOUT-.n35 GNDA 0.19586f
C2073 VOUT-.n36 GNDA 0.237352f
C2074 VOUT-.t100 GNDA 0.297101f
C2075 VOUT-.t47 GNDA 0.292125f
C2076 VOUT-.n37 GNDA 0.19586f
C2077 VOUT-.t153 GNDA 0.292125f
C2078 VOUT-.t71 GNDA 0.297101f
C2079 VOUT-.t123 GNDA 0.292125f
C2080 VOUT-.n38 GNDA 0.19586f
C2081 VOUT-.n39 GNDA 0.237352f
C2082 VOUT-.t69 GNDA 0.297101f
C2083 VOUT-.t154 GNDA 0.292125f
C2084 VOUT-.n40 GNDA 0.19586f
C2085 VOUT-.t124 GNDA 0.292125f
C2086 VOUT-.t35 GNDA 0.297101f
C2087 VOUT-.t86 GNDA 0.292125f
C2088 VOUT-.n41 GNDA 0.19586f
C2089 VOUT-.n42 GNDA 0.237352f
C2090 VOUT-.t96 GNDA 0.292125f
C2091 VOUT-.t85 GNDA 0.297101f
C2092 VOUT-.t57 GNDA 0.292125f
C2093 VOUT-.n43 GNDA 0.19586f
C2094 VOUT-.n44 GNDA 0.127805f
C2095 VOUT-.t132 GNDA 0.296478f
C2096 VOUT-.t115 GNDA 0.296478f
C2097 VOUT-.t131 GNDA 0.297101f
C2098 VOUT-.t104 GNDA 0.292125f
C2099 VOUT-.n45 GNDA 0.19586f
C2100 VOUT-.t73 GNDA 0.292125f
C2101 VOUT-.n46 GNDA 0.12324f
C2102 VOUT-.t146 GNDA 0.296478f
C2103 VOUT-.t31 GNDA 0.297101f
C2104 VOUT-.t138 GNDA 0.292125f
C2105 VOUT-.n47 GNDA 0.19586f
C2106 VOUT-.t107 GNDA 0.292125f
C2107 VOUT-.n48 GNDA 0.12324f
C2108 VOUT-.t46 GNDA 0.296478f
C2109 VOUT-.t62 GNDA 0.297101f
C2110 VOUT-.t41 GNDA 0.292125f
C2111 VOUT-.n49 GNDA 0.19586f
C2112 VOUT-.t143 GNDA 0.292125f
C2113 VOUT-.n50 GNDA 0.12324f
C2114 VOUT-.t87 GNDA 0.296478f
C2115 VOUT-.t114 GNDA 0.297101f
C2116 VOUT-.t21 GNDA 0.292125f
C2117 VOUT-.n51 GNDA 0.19586f
C2118 VOUT-.t126 GNDA 0.292125f
C2119 VOUT-.n52 GNDA 0.12324f
C2120 VOUT-.t65 GNDA 0.296478f
C2121 VOUT-.t26 GNDA 0.296722f
C2122 VOUT-.t102 GNDA 0.296478f
C2123 VOUT-.t59 GNDA 0.296722f
C2124 VOUT-.t134 GNDA 0.296478f
C2125 VOUT-.t37 GNDA 0.296722f
C2126 VOUT-.t120 GNDA 0.296478f
C2127 VOUT-.t81 GNDA 0.296722f
C2128 VOUT-.t155 GNDA 0.296478f
C2129 VOUT-.t119 GNDA 0.292125f
C2130 VOUT-.n53 GNDA 0.323342f
C2131 VOUT-.t82 GNDA 0.292125f
C2132 VOUT-.n54 GNDA 0.378116f
C2133 VOUT-.t97 GNDA 0.292125f
C2134 VOUT-.n55 GNDA 0.378116f
C2135 VOUT-.t63 GNDA 0.292125f
C2136 VOUT-.n56 GNDA 0.378116f
C2137 VOUT-.t27 GNDA 0.292125f
C2138 VOUT-.n57 GNDA 0.310595f
C2139 VOUT-.t45 GNDA 0.292125f
C2140 VOUT-.n58 GNDA 0.310595f
C2141 VOUT-.t144 GNDA 0.292125f
C2142 VOUT-.n59 GNDA 0.310595f
C2143 VOUT-.t112 GNDA 0.292125f
C2144 VOUT-.n60 GNDA 0.310595f
C2145 VOUT-.t76 GNDA 0.292125f
C2146 VOUT-.n61 GNDA 0.251257f
C2147 VOUT-.t93 GNDA 0.292125f
C2148 VOUT-.n62 GNDA 0.251257f
C2149 VOUT-.t56 GNDA 0.292125f
C2150 VOUT-.t40 GNDA 0.297101f
C2151 VOUT-.t19 GNDA 0.292125f
C2152 VOUT-.n63 GNDA 0.19586f
C2153 VOUT-.n64 GNDA 0.237352f
C2154 VOUT-.t34 GNDA 0.297101f
C2155 VOUT-.t52 GNDA 0.292125f
C2156 VOUT-.n65 GNDA 0.19586f
C2157 VOUT-.t156 GNDA 0.292125f
C2158 VOUT-.t136 GNDA 0.297101f
C2159 VOUT-.t121 GNDA 0.292125f
C2160 VOUT-.n66 GNDA 0.19586f
C2161 VOUT-.n67 GNDA 0.237352f
C2162 VOUT-.t70 GNDA 0.297101f
C2163 VOUT-.t89 GNDA 0.292125f
C2164 VOUT-.n68 GNDA 0.19586f
C2165 VOUT-.t50 GNDA 0.292125f
C2166 VOUT-.t36 GNDA 0.297101f
C2167 VOUT-.t151 GNDA 0.292125f
C2168 VOUT-.n69 GNDA 0.19586f
C2169 VOUT-.n70 GNDA 0.237352f
C2170 VOUT-.t95 GNDA 0.297101f
C2171 VOUT-.t43 GNDA 0.292125f
C2172 VOUT-.n71 GNDA 0.19586f
C2173 VOUT-.t145 GNDA 0.292125f
C2174 VOUT-.t66 GNDA 0.297101f
C2175 VOUT-.t118 GNDA 0.292125f
C2176 VOUT-.n72 GNDA 0.19586f
C2177 VOUT-.n73 GNDA 0.237352f
C2178 VOUT-.t55 GNDA 0.297101f
C2179 VOUT-.t141 GNDA 0.292125f
C2180 VOUT-.n74 GNDA 0.19586f
C2181 VOUT-.t111 GNDA 0.292125f
C2182 VOUT-.t29 GNDA 0.297101f
C2183 VOUT-.t80 GNDA 0.292125f
C2184 VOUT-.n75 GNDA 0.19586f
C2185 VOUT-.n76 GNDA 0.237352f
C2186 VOUT-.t91 GNDA 0.297101f
C2187 VOUT-.t39 GNDA 0.292125f
C2188 VOUT-.n77 GNDA 0.19586f
C2189 VOUT-.t139 GNDA 0.292125f
C2190 VOUT-.t58 GNDA 0.297101f
C2191 VOUT-.t109 GNDA 0.292125f
C2192 VOUT-.n78 GNDA 0.19586f
C2193 VOUT-.n79 GNDA 0.237352f
C2194 VOUT-.t49 GNDA 0.297101f
C2195 VOUT-.t135 GNDA 0.292125f
C2196 VOUT-.n80 GNDA 0.19586f
C2197 VOUT-.t103 GNDA 0.292125f
C2198 VOUT-.t20 GNDA 0.297101f
C2199 VOUT-.t72 GNDA 0.292125f
C2200 VOUT-.n81 GNDA 0.19586f
C2201 VOUT-.n82 GNDA 0.237352f
C2202 VOUT-.t148 GNDA 0.297101f
C2203 VOUT-.t99 GNDA 0.292125f
C2204 VOUT-.n83 GNDA 0.19586f
C2205 VOUT-.t68 GNDA 0.292125f
C2206 VOUT-.t122 GNDA 0.297101f
C2207 VOUT-.t33 GNDA 0.292125f
C2208 VOUT-.n84 GNDA 0.19586f
C2209 VOUT-.n85 GNDA 0.237352f
C2210 VOUT-.t44 GNDA 0.297101f
C2211 VOUT-.t133 GNDA 0.292125f
C2212 VOUT-.n86 GNDA 0.19586f
C2213 VOUT-.t98 GNDA 0.292125f
C2214 VOUT-.t152 GNDA 0.297101f
C2215 VOUT-.t67 GNDA 0.292125f
C2216 VOUT-.n87 GNDA 0.19586f
C2217 VOUT-.n88 GNDA 0.237352f
C2218 VOUT-.t142 GNDA 0.297101f
C2219 VOUT-.t94 GNDA 0.292125f
C2220 VOUT-.n89 GNDA 0.19586f
C2221 VOUT-.t60 GNDA 0.292125f
C2222 VOUT-.t116 GNDA 0.297101f
C2223 VOUT-.t30 GNDA 0.292125f
C2224 VOUT-.n90 GNDA 0.19586f
C2225 VOUT-.n91 GNDA 0.237352f
C2226 VOUT-.t77 GNDA 0.297101f
C2227 VOUT-.t127 GNDA 0.292125f
C2228 VOUT-.n92 GNDA 0.19586f
C2229 VOUT-.t22 GNDA 0.292125f
C2230 VOUT-.n93 GNDA 0.237352f
C2231 VOUT-.t53 GNDA 0.292125f
C2232 VOUT-.n94 GNDA 0.127805f
C2233 VOUT-.t105 GNDA 0.292125f
C2234 VOUT-.n95 GNDA 0.23231f
C2235 VOUT-.n96 GNDA 0.521555f
C2236 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.325502f
C2237 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013595f
C2238 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013595f
C2239 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.045371f
C2240 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013595f
C2241 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013595f
C2242 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.048807f
C2243 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013595f
C2244 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013595f
C2245 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.048807f
C2246 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013595f
C2247 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013595f
C2248 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.048495f
C2249 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013595f
C2250 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013595f
C2251 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.048495f
C2252 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.139712f
C2253 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.103838f
C2254 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013595f
C2255 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013595f
C2256 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.044102f
C2257 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013595f
C2258 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013595f
C2259 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.047844f
C2260 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013595f
C2261 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013595f
C2262 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.046785f
C2263 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.199933f
C2264 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013595f
C2265 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013595f
C2266 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.046785f
C2267 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.143094f
C2268 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013595f
C2269 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013595f
C2270 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.047844f
C2271 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013595f
C2272 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013595f
C2273 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.046785f
C2274 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.199933f
C2275 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.081571f
C2276 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.087203f
C2277 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.19992f
C2278 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.212963f
C2279 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.19992f
C2280 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 1.62043f
C2281 two_stage_opamp_dummy_magic_0.V_tot.t11 GNDA 0.010451f
C2282 two_stage_opamp_dummy_magic_0.V_tot.t5 GNDA 0.010451f
C2283 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.046799f
C2284 two_stage_opamp_dummy_magic_0.V_tot.t12 GNDA 0.010451f
C2285 two_stage_opamp_dummy_magic_0.V_tot.t8 GNDA 0.010451f
C2286 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.046195f
C2287 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.349166f
C2288 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.023984f
C2289 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.19579f
C2290 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.024032f
C2291 two_stage_opamp_dummy_magic_0.V_tot.t9 GNDA 0.010835f
C2292 two_stage_opamp_dummy_magic_0.V_tot.t10 GNDA 0.010835f
C2293 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.039314f
C2294 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.324506f
C2295 two_stage_opamp_dummy_magic_0.V_tot.t7 GNDA 0.010451f
C2296 two_stage_opamp_dummy_magic_0.V_tot.t13 GNDA 0.010451f
C2297 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.046195f
C2298 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.256256f
C2299 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.311983f
C2300 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 3.27399f
C2301 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 1.6312f
C2302 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.212987f
C2303 bgr_0.cap_res1.t6 GNDA 0.417173f
C2304 bgr_0.cap_res1.t10 GNDA 0.418684f
C2305 bgr_0.cap_res1.t0 GNDA 0.417173f
C2306 bgr_0.cap_res1.t14 GNDA 0.418684f
C2307 bgr_0.cap_res1.t3 GNDA 0.417173f
C2308 bgr_0.cap_res1.t7 GNDA 0.418684f
C2309 bgr_0.cap_res1.t15 GNDA 0.417173f
C2310 bgr_0.cap_res1.t9 GNDA 0.418684f
C2311 bgr_0.cap_res1.t8 GNDA 0.417173f
C2312 bgr_0.cap_res1.t12 GNDA 0.418684f
C2313 bgr_0.cap_res1.t1 GNDA 0.417173f
C2314 bgr_0.cap_res1.t16 GNDA 0.418684f
C2315 bgr_0.cap_res1.t13 GNDA 0.417173f
C2316 bgr_0.cap_res1.t19 GNDA 0.418684f
C2317 bgr_0.cap_res1.t5 GNDA 0.417173f
C2318 bgr_0.cap_res1.t2 GNDA 0.418684f
C2319 bgr_0.cap_res1.n0 GNDA 0.279631f
C2320 bgr_0.cap_res1.t4 GNDA 0.222685f
C2321 bgr_0.cap_res1.n1 GNDA 0.303406f
C2322 bgr_0.cap_res1.t18 GNDA 0.222685f
C2323 bgr_0.cap_res1.n2 GNDA 0.303406f
C2324 bgr_0.cap_res1.t11 GNDA 0.222685f
C2325 bgr_0.cap_res1.n3 GNDA 0.303406f
C2326 bgr_0.cap_res1.t17 GNDA 0.649059f
C2327 bgr_0.cap_res1.t20 GNDA 0.10618f
C2328 bgr_0.1st_Vout_1.n0 GNDA 0.573726f
C2329 bgr_0.1st_Vout_1.n1 GNDA 1.42916f
C2330 bgr_0.1st_Vout_1.n2 GNDA 1.78489f
C2331 bgr_0.1st_Vout_1.n3 GNDA 0.125562f
C2332 bgr_0.1st_Vout_1.t20 GNDA 0.352846f
C2333 bgr_0.1st_Vout_1.t11 GNDA 0.346937f
C2334 bgr_0.1st_Vout_1.t32 GNDA 0.346937f
C2335 bgr_0.1st_Vout_1.t29 GNDA 0.352846f
C2336 bgr_0.1st_Vout_1.t34 GNDA 0.346937f
C2337 bgr_0.1st_Vout_1.t25 GNDA 0.352846f
C2338 bgr_0.1st_Vout_1.t21 GNDA 0.346937f
C2339 bgr_0.1st_Vout_1.t12 GNDA 0.346937f
C2340 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C2341 bgr_0.1st_Vout_1.t16 GNDA 0.346937f
C2342 bgr_0.1st_Vout_1.t33 GNDA 0.352846f
C2343 bgr_0.1st_Vout_1.t26 GNDA 0.346937f
C2344 bgr_0.1st_Vout_1.t22 GNDA 0.346937f
C2345 bgr_0.1st_Vout_1.t17 GNDA 0.352846f
C2346 bgr_0.1st_Vout_1.t24 GNDA 0.346937f
C2347 bgr_0.1st_Vout_1.t28 GNDA 0.352846f
C2348 bgr_0.1st_Vout_1.t23 GNDA 0.346937f
C2349 bgr_0.1st_Vout_1.t13 GNDA 0.346937f
C2350 bgr_0.1st_Vout_1.t18 GNDA 0.346937f
C2351 bgr_0.1st_Vout_1.t36 GNDA 0.346937f
C2352 bgr_0.1st_Vout_1.t30 GNDA 0.022665f
C2353 bgr_0.1st_Vout_1.n4 GNDA 0.021864f
C2354 bgr_0.1st_Vout_1.t14 GNDA 0.013213f
C2355 bgr_0.1st_Vout_1.t31 GNDA 0.013213f
C2356 bgr_0.1st_Vout_1.n5 GNDA 0.029393f
C2357 bgr_0.1st_Vout_1.t0 GNDA 0.018268f
C2358 bgr_0.1st_Vout_1.n6 GNDA 0.012529f
C2359 bgr_0.1st_Vout_1.n7 GNDA 0.189508f
C2360 bgr_0.1st_Vout_1.n8 GNDA 0.011336f
C2361 bgr_0.1st_Vout_1.n9 GNDA 0.020958f
C2362 bgr_0.1st_Vout_1.t19 GNDA 0.013213f
C2363 bgr_0.1st_Vout_1.t27 GNDA 0.013213f
C2364 bgr_0.1st_Vout_1.n10 GNDA 0.029393f
C2365 bgr_0.1st_Vout_1.n11 GNDA 0.021864f
C2366 bgr_0.1st_Vout_1.t15 GNDA 0.020738f
C2367 VDDA.t250 GNDA 0.027842f
C2368 VDDA.t444 GNDA 0.027842f
C2369 VDDA.n0 GNDA 0.120197f
C2370 VDDA.t85 GNDA 0.027842f
C2371 VDDA.t195 GNDA 0.027842f
C2372 VDDA.n1 GNDA 0.119954f
C2373 VDDA.n2 GNDA 0.138502f
C2374 VDDA.t84 GNDA 0.027842f
C2375 VDDA.t194 GNDA 0.027842f
C2376 VDDA.n3 GNDA 0.119954f
C2377 VDDA.n4 GNDA 0.074245f
C2378 VDDA.t40 GNDA 0.027842f
C2379 VDDA.t130 GNDA 0.027842f
C2380 VDDA.n5 GNDA 0.119954f
C2381 VDDA.n6 GNDA 0.074245f
C2382 VDDA.t131 GNDA 0.027842f
C2383 VDDA.t246 GNDA 0.027842f
C2384 VDDA.n7 GNDA 0.119954f
C2385 VDDA.n8 GNDA 0.074245f
C2386 VDDA.t103 GNDA 0.027842f
C2387 VDDA.t255 GNDA 0.027842f
C2388 VDDA.n9 GNDA 0.119954f
C2389 VDDA.n10 GNDA 0.218007f
C2390 VDDA.n11 GNDA 0.06743f
C2391 VDDA.n12 GNDA 0.180018f
C2392 VDDA.t426 GNDA 0.013115f
C2393 VDDA.n13 GNDA 0.028951f
C2394 VDDA.n14 GNDA 0.043275f
C2395 VDDA.n15 GNDA 0.068106f
C2396 VDDA.n16 GNDA 0.181504f
C2397 VDDA.t356 GNDA 0.013115f
C2398 VDDA.n17 GNDA 0.028951f
C2399 VDDA.n18 GNDA 0.040287f
C2400 VDDA.n19 GNDA 0.045739f
C2401 VDDA.n20 GNDA 0.181504f
C2402 VDDA.t355 GNDA 0.176569f
C2403 VDDA.t175 GNDA 0.109106f
C2404 VDDA.t102 GNDA 0.109106f
C2405 VDDA.t451 GNDA 0.109106f
C2406 VDDA.t144 GNDA 0.109106f
C2407 VDDA.t174 GNDA 0.08183f
C2408 VDDA.t379 GNDA 0.176569f
C2409 VDDA.t447 GNDA 0.109106f
C2410 VDDA.t119 GNDA 0.109106f
C2411 VDDA.t201 GNDA 0.109106f
C2412 VDDA.t98 GNDA 0.109106f
C2413 VDDA.t43 GNDA 0.08183f
C2414 VDDA.n21 GNDA 0.068781f
C2415 VDDA.n22 GNDA 0.054553f
C2416 VDDA.n23 GNDA 0.068781f
C2417 VDDA.n24 GNDA 0.043851f
C2418 VDDA.t380 GNDA 0.013115f
C2419 VDDA.n25 GNDA 0.028951f
C2420 VDDA.n26 GNDA 0.039714f
C2421 VDDA.n27 GNDA 0.095712f
C2422 VDDA.n28 GNDA 0.095712f
C2423 VDDA.n29 GNDA 0.180018f
C2424 VDDA.t425 GNDA 0.173008f
C2425 VDDA.t99 GNDA 0.107192f
C2426 VDDA.t452 GNDA 0.107192f
C2427 VDDA.t70 GNDA 0.107192f
C2428 VDDA.t218 GNDA 0.107192f
C2429 VDDA.t254 GNDA 0.080394f
C2430 VDDA.t319 GNDA 0.173008f
C2431 VDDA.t225 GNDA 0.107192f
C2432 VDDA.t135 GNDA 0.107192f
C2433 VDDA.t253 GNDA 0.107192f
C2434 VDDA.t82 GNDA 0.107192f
C2435 VDDA.t45 GNDA 0.080394f
C2436 VDDA.n30 GNDA 0.068781f
C2437 VDDA.n31 GNDA 0.053596f
C2438 VDDA.n32 GNDA 0.068781f
C2439 VDDA.n33 GNDA 0.043422f
C2440 VDDA.t320 GNDA 0.013115f
C2441 VDDA.n34 GNDA 0.028951f
C2442 VDDA.n35 GNDA 0.039714f
C2443 VDDA.n36 GNDA 0.076706f
C2444 VDDA.n37 GNDA 0.43487f
C2445 VDDA.t240 GNDA 0.041763f
C2446 VDDA.t129 GNDA 0.041763f
C2447 VDDA.n38 GNDA 0.166563f
C2448 VDDA.n39 GNDA 0.097241f
C2449 VDDA.t326 GNDA 0.041603f
C2450 VDDA.n40 GNDA 0.05522f
C2451 VDDA.n41 GNDA 0.079516f
C2452 VDDA.t359 GNDA 0.046205f
C2453 VDDA.t357 GNDA 0.020234f
C2454 VDDA.n42 GNDA 0.074338f
C2455 VDDA.n43 GNDA 0.045655f
C2456 VDDA.t329 GNDA 0.046205f
C2457 VDDA.t327 GNDA 0.020234f
C2458 VDDA.n44 GNDA 0.074338f
C2459 VDDA.n45 GNDA 0.045655f
C2460 VDDA.n46 GNDA 0.043851f
C2461 VDDA.n47 GNDA 0.079516f
C2462 VDDA.n48 GNDA 0.229873f
C2463 VDDA.t328 GNDA 0.284691f
C2464 VDDA.t242 GNDA 0.164616f
C2465 VDDA.t249 GNDA 0.164616f
C2466 VDDA.t234 GNDA 0.164616f
C2467 VDDA.t196 GNDA 0.164616f
C2468 VDDA.t257 GNDA 0.123462f
C2469 VDDA.n49 GNDA 0.082308f
C2470 VDDA.t132 GNDA 0.123462f
C2471 VDDA.t243 GNDA 0.164616f
C2472 VDDA.t3 GNDA 0.164616f
C2473 VDDA.t241 GNDA 0.164616f
C2474 VDDA.t256 GNDA 0.164616f
C2475 VDDA.t358 GNDA 0.284691f
C2476 VDDA.n50 GNDA 0.229873f
C2477 VDDA.n51 GNDA 0.05522f
C2478 VDDA.n52 GNDA 0.115651f
C2479 VDDA.n53 GNDA 0.079909f
C2480 VDDA.n54 GNDA 0.108214f
C2481 VDDA.n55 GNDA 0.108214f
C2482 VDDA.n56 GNDA 0.107508f
C2483 VDDA.t347 GNDA 0.041603f
C2484 VDDA.t236 GNDA 0.041763f
C2485 VDDA.t198 GNDA 0.041763f
C2486 VDDA.n57 GNDA 0.166563f
C2487 VDDA.n58 GNDA 0.097241f
C2488 VDDA.t248 GNDA 0.041763f
C2489 VDDA.t42 GNDA 0.041763f
C2490 VDDA.n59 GNDA 0.166563f
C2491 VDDA.n60 GNDA 0.097241f
C2492 VDDA.t245 GNDA 0.041763f
C2493 VDDA.t5 GNDA 0.041763f
C2494 VDDA.n61 GNDA 0.166563f
C2495 VDDA.n62 GNDA 0.097241f
C2496 VDDA.t238 GNDA 0.041763f
C2497 VDDA.t259 GNDA 0.041763f
C2498 VDDA.n63 GNDA 0.166563f
C2499 VDDA.n64 GNDA 0.19871f
C2500 VDDA.n65 GNDA 0.133588f
C2501 VDDA.t345 GNDA 0.050479f
C2502 VDDA.n66 GNDA 0.097627f
C2503 VDDA.n67 GNDA 0.058909f
C2504 VDDA.n68 GNDA 0.08334f
C2505 VDDA.n69 GNDA 0.371616f
C2506 VDDA.t346 GNDA 0.573999f
C2507 VDDA.t258 GNDA 0.317748f
C2508 VDDA.t237 GNDA 0.317748f
C2509 VDDA.t4 GNDA 0.317748f
C2510 VDDA.t244 GNDA 0.317748f
C2511 VDDA.t41 GNDA 0.238311f
C2512 VDDA.n70 GNDA 0.158874f
C2513 VDDA.t247 GNDA 0.238311f
C2514 VDDA.t197 GNDA 0.317748f
C2515 VDDA.t235 GNDA 0.317748f
C2516 VDDA.t128 GNDA 0.317748f
C2517 VDDA.t239 GNDA 0.317748f
C2518 VDDA.t325 GNDA 0.573999f
C2519 VDDA.n71 GNDA 0.371616f
C2520 VDDA.n72 GNDA 0.08334f
C2521 VDDA.n73 GNDA 0.058909f
C2522 VDDA.t324 GNDA 0.050479f
C2523 VDDA.n74 GNDA 0.097627f
C2524 VDDA.n75 GNDA 0.13335f
C2525 VDDA.n76 GNDA 0.145951f
C2526 VDDA.n77 GNDA 0.183365f
C2527 VDDA.t89 GNDA 0.024362f
C2528 VDDA.t233 GNDA 0.024362f
C2529 VDDA.n78 GNDA 0.083842f
C2530 VDDA.t69 GNDA 0.024362f
C2531 VDDA.t227 GNDA 0.024362f
C2532 VDDA.n79 GNDA 0.083638f
C2533 VDDA.n80 GNDA 0.180547f
C2534 VDDA.t440 GNDA 0.024362f
C2535 VDDA.t21 GNDA 0.024362f
C2536 VDDA.n81 GNDA 0.083842f
C2537 VDDA.t123 GNDA 0.024362f
C2538 VDDA.t2 GNDA 0.024362f
C2539 VDDA.n82 GNDA 0.083638f
C2540 VDDA.n83 GNDA 0.180547f
C2541 VDDA.n84 GNDA 0.033411f
C2542 VDDA.n85 GNDA 0.066846f
C2543 VDDA.n86 GNDA 0.066846f
C2544 VDDA.n87 GNDA 0.28106f
C2545 VDDA.n88 GNDA 0.28106f
C2546 VDDA.t367 GNDA 0.419522f
C2547 VDDA.t88 GNDA 0.242226f
C2548 VDDA.t232 GNDA 0.242226f
C2549 VDDA.t68 GNDA 0.242226f
C2550 VDDA.t226 GNDA 0.242226f
C2551 VDDA.t188 GNDA 0.18167f
C2552 VDDA.t368 GNDA 0.120182f
C2553 VDDA.t366 GNDA 0.042422f
C2554 VDDA.n89 GNDA 0.079448f
C2555 VDDA.n90 GNDA 0.053036f
C2556 VDDA.t417 GNDA 0.120182f
C2557 VDDA.t415 GNDA 0.042422f
C2558 VDDA.n91 GNDA 0.079448f
C2559 VDDA.n92 GNDA 0.053036f
C2560 VDDA.n93 GNDA 0.048028f
C2561 VDDA.n94 GNDA 0.09431f
C2562 VDDA.t416 GNDA 0.419522f
C2563 VDDA.t20 GNDA 0.242226f
C2564 VDDA.t439 GNDA 0.242226f
C2565 VDDA.t1 GNDA 0.242226f
C2566 VDDA.t122 GNDA 0.242226f
C2567 VDDA.t228 GNDA 0.18167f
C2568 VDDA.n95 GNDA 0.121113f
C2569 VDDA.n96 GNDA 0.09431f
C2570 VDDA.n97 GNDA 0.101302f
C2571 VDDA.t189 GNDA 0.024362f
C2572 VDDA.t229 GNDA 0.024362f
C2573 VDDA.n98 GNDA 0.07828f
C2574 VDDA.n99 GNDA 0.058147f
C2575 VDDA.n100 GNDA 0.058709f
C2576 VDDA.t110 GNDA 0.027842f
C2577 VDDA.t44 GNDA 0.027842f
C2578 VDDA.n101 GNDA 0.120197f
C2579 VDDA.t177 GNDA 0.027842f
C2580 VDDA.t90 GNDA 0.027842f
C2581 VDDA.n102 GNDA 0.119954f
C2582 VDDA.n103 GNDA 0.138502f
C2583 VDDA.t0 GNDA 0.027842f
C2584 VDDA.t460 GNDA 0.027842f
C2585 VDDA.n104 GNDA 0.119954f
C2586 VDDA.n105 GNDA 0.074245f
C2587 VDDA.t178 GNDA 0.027842f
C2588 VDDA.t448 GNDA 0.027842f
C2589 VDDA.n106 GNDA 0.119954f
C2590 VDDA.n107 GNDA 0.074245f
C2591 VDDA.t13 GNDA 0.027842f
C2592 VDDA.t185 GNDA 0.027842f
C2593 VDDA.n108 GNDA 0.119954f
C2594 VDDA.n109 GNDA 0.074245f
C2595 VDDA.t163 GNDA 0.027842f
C2596 VDDA.t176 GNDA 0.027842f
C2597 VDDA.n110 GNDA 0.119954f
C2598 VDDA.n111 GNDA 0.268748f
C2599 VDDA.t442 GNDA 0.041763f
C2600 VDDA.t12 GNDA 0.041763f
C2601 VDDA.n112 GNDA 0.166563f
C2602 VDDA.n113 GNDA 0.097241f
C2603 VDDA.t371 GNDA 0.041603f
C2604 VDDA.n114 GNDA 0.08334f
C2605 VDDA.t341 GNDA 0.041603f
C2606 VDDA.t134 GNDA 0.041763f
C2607 VDDA.t139 GNDA 0.041763f
C2608 VDDA.n115 GNDA 0.166563f
C2609 VDDA.n116 GNDA 0.097241f
C2610 VDDA.t167 GNDA 0.041763f
C2611 VDDA.t137 GNDA 0.041763f
C2612 VDDA.n117 GNDA 0.166563f
C2613 VDDA.n118 GNDA 0.097241f
C2614 VDDA.t31 GNDA 0.041763f
C2615 VDDA.t15 GNDA 0.041763f
C2616 VDDA.n119 GNDA 0.166563f
C2617 VDDA.n120 GNDA 0.097241f
C2618 VDDA.t105 GNDA 0.041763f
C2619 VDDA.t169 GNDA 0.041763f
C2620 VDDA.n121 GNDA 0.166563f
C2621 VDDA.n122 GNDA 0.19871f
C2622 VDDA.n123 GNDA 0.133588f
C2623 VDDA.t339 GNDA 0.050479f
C2624 VDDA.n124 GNDA 0.097627f
C2625 VDDA.n125 GNDA 0.058909f
C2626 VDDA.n126 GNDA 0.05522f
C2627 VDDA.n127 GNDA 0.079516f
C2628 VDDA.t377 GNDA 0.046205f
C2629 VDDA.t375 GNDA 0.020234f
C2630 VDDA.n128 GNDA 0.074338f
C2631 VDDA.n129 GNDA 0.045655f
C2632 VDDA.t353 GNDA 0.046205f
C2633 VDDA.t351 GNDA 0.020234f
C2634 VDDA.n130 GNDA 0.074338f
C2635 VDDA.n131 GNDA 0.045655f
C2636 VDDA.n132 GNDA 0.043851f
C2637 VDDA.n133 GNDA 0.079516f
C2638 VDDA.n134 GNDA 0.229873f
C2639 VDDA.t352 GNDA 0.284691f
C2640 VDDA.t93 GNDA 0.164616f
C2641 VDDA.t215 GNDA 0.164616f
C2642 VDDA.t453 GNDA 0.164616f
C2643 VDDA.t83 GNDA 0.164616f
C2644 VDDA.t214 GNDA 0.123462f
C2645 VDDA.n135 GNDA 0.082308f
C2646 VDDA.t443 GNDA 0.123462f
C2647 VDDA.t435 GNDA 0.164616f
C2648 VDDA.t436 GNDA 0.164616f
C2649 VDDA.t81 GNDA 0.164616f
C2650 VDDA.t10 GNDA 0.164616f
C2651 VDDA.t376 GNDA 0.284691f
C2652 VDDA.n136 GNDA 0.229873f
C2653 VDDA.n137 GNDA 0.05522f
C2654 VDDA.n138 GNDA 0.115651f
C2655 VDDA.n139 GNDA 0.371616f
C2656 VDDA.n140 GNDA 0.371616f
C2657 VDDA.t340 GNDA 0.573999f
C2658 VDDA.t104 GNDA 0.317748f
C2659 VDDA.t168 GNDA 0.317748f
C2660 VDDA.t30 GNDA 0.317748f
C2661 VDDA.t14 GNDA 0.317748f
C2662 VDDA.t166 GNDA 0.238311f
C2663 VDDA.t370 GNDA 0.573999f
C2664 VDDA.t11 GNDA 0.317748f
C2665 VDDA.t441 GNDA 0.317748f
C2666 VDDA.t138 GNDA 0.317748f
C2667 VDDA.t133 GNDA 0.317748f
C2668 VDDA.t136 GNDA 0.238311f
C2669 VDDA.n141 GNDA 0.08334f
C2670 VDDA.n142 GNDA 0.108214f
C2671 VDDA.n143 GNDA 0.108214f
C2672 VDDA.n144 GNDA 0.158874f
C2673 VDDA.n145 GNDA 0.107508f
C2674 VDDA.n146 GNDA 0.079909f
C2675 VDDA.n147 GNDA 0.058909f
C2676 VDDA.t369 GNDA 0.050479f
C2677 VDDA.n148 GNDA 0.097627f
C2678 VDDA.n149 GNDA 0.13335f
C2679 VDDA.n150 GNDA 0.1205f
C2680 VDDA.n152 GNDA 0.064437f
C2681 VDDA.n153 GNDA 0.082134f
C2682 VDDA.n154 GNDA 0.10686f
C2683 VDDA.n155 GNDA 0.10686f
C2684 VDDA.n156 GNDA 0.10686f
C2685 VDDA.n158 GNDA 0.064437f
C2686 VDDA.n160 GNDA 0.064437f
C2687 VDDA.n162 GNDA 0.064437f
C2688 VDDA.n164 GNDA 0.064437f
C2689 VDDA.n166 GNDA 0.064437f
C2690 VDDA.n168 GNDA 0.064437f
C2691 VDDA.n170 GNDA 0.064437f
C2692 VDDA.n172 GNDA 0.064437f
C2693 VDDA.n174 GNDA 0.1032f
C2694 VDDA.t402 GNDA 0.012682f
C2695 VDDA.n175 GNDA 0.020249f
C2696 VDDA.n176 GNDA 0.017705f
C2697 VDDA.n177 GNDA 0.059428f
C2698 VDDA.n178 GNDA 0.064983f
C2699 VDDA.n179 GNDA 0.218506f
C2700 VDDA.t401 GNDA 0.173008f
C2701 VDDA.t62 GNDA 0.107192f
C2702 VDDA.t463 GNDA 0.107192f
C2703 VDDA.t79 GNDA 0.107192f
C2704 VDDA.t149 GNDA 0.107192f
C2705 VDDA.t427 GNDA 0.107192f
C2706 VDDA.t212 GNDA 0.107192f
C2707 VDDA.t26 GNDA 0.107192f
C2708 VDDA.t126 GNDA 0.107192f
C2709 VDDA.t223 GNDA 0.107192f
C2710 VDDA.t465 GNDA 0.080394f
C2711 VDDA.n180 GNDA 0.053596f
C2712 VDDA.t467 GNDA 0.080394f
C2713 VDDA.t251 GNDA 0.107192f
C2714 VDDA.t86 GNDA 0.107192f
C2715 VDDA.t157 GNDA 0.107192f
C2716 VDDA.t219 GNDA 0.107192f
C2717 VDDA.t151 GNDA 0.107192f
C2718 VDDA.t28 GNDA 0.107192f
C2719 VDDA.t431 GNDA 0.107192f
C2720 VDDA.t210 GNDA 0.107192f
C2721 VDDA.t221 GNDA 0.107192f
C2722 VDDA.t407 GNDA 0.173008f
C2723 VDDA.n181 GNDA 0.218506f
C2724 VDDA.n182 GNDA 0.064983f
C2725 VDDA.n183 GNDA 0.059428f
C2726 VDDA.n184 GNDA 0.017705f
C2727 VDDA.t408 GNDA 0.012682f
C2728 VDDA.n185 GNDA 0.019891f
C2729 VDDA.n186 GNDA 0.10107f
C2730 VDDA.n187 GNDA 0.091879f
C2731 VDDA.n188 GNDA 0.582978f
C2732 VDDA.n189 GNDA 0.470301f
C2733 VDDA.t193 GNDA 0.024362f
C2734 VDDA.t19 GNDA 0.024362f
C2735 VDDA.n190 GNDA 0.083842f
C2736 VDDA.t457 GNDA 0.024362f
C2737 VDDA.t33 GNDA 0.024362f
C2738 VDDA.n191 GNDA 0.083638f
C2739 VDDA.n192 GNDA 0.180547f
C2740 VDDA.t118 GNDA 0.024362f
C2741 VDDA.t173 GNDA 0.024362f
C2742 VDDA.n193 GNDA 0.083842f
C2743 VDDA.t187 GNDA 0.024362f
C2744 VDDA.t231 GNDA 0.024362f
C2745 VDDA.n194 GNDA 0.083638f
C2746 VDDA.n195 GNDA 0.180547f
C2747 VDDA.n196 GNDA 0.033411f
C2748 VDDA.n197 GNDA 0.066846f
C2749 VDDA.n198 GNDA 0.066846f
C2750 VDDA.n199 GNDA 0.28106f
C2751 VDDA.n200 GNDA 0.28106f
C2752 VDDA.t361 GNDA 0.419522f
C2753 VDDA.t192 GNDA 0.242226f
C2754 VDDA.t18 GNDA 0.242226f
C2755 VDDA.t456 GNDA 0.242226f
C2756 VDDA.t32 GNDA 0.242226f
C2757 VDDA.t190 GNDA 0.18167f
C2758 VDDA.t362 GNDA 0.120182f
C2759 VDDA.t360 GNDA 0.042422f
C2760 VDDA.n201 GNDA 0.079448f
C2761 VDDA.n202 GNDA 0.053036f
C2762 VDDA.t396 GNDA 0.120182f
C2763 VDDA.t394 GNDA 0.042422f
C2764 VDDA.n203 GNDA 0.079448f
C2765 VDDA.n204 GNDA 0.053036f
C2766 VDDA.n205 GNDA 0.048028f
C2767 VDDA.n206 GNDA 0.09431f
C2768 VDDA.t395 GNDA 0.419522f
C2769 VDDA.t172 GNDA 0.242226f
C2770 VDDA.t117 GNDA 0.242226f
C2771 VDDA.t230 GNDA 0.242226f
C2772 VDDA.t186 GNDA 0.242226f
C2773 VDDA.t6 GNDA 0.18167f
C2774 VDDA.n207 GNDA 0.121113f
C2775 VDDA.n208 GNDA 0.09431f
C2776 VDDA.n209 GNDA 0.101302f
C2777 VDDA.t191 GNDA 0.024362f
C2778 VDDA.t7 GNDA 0.024362f
C2779 VDDA.n210 GNDA 0.07828f
C2780 VDDA.n211 GNDA 0.058147f
C2781 VDDA.n212 GNDA 0.058408f
C2782 VDDA.n213 GNDA 0.425348f
C2783 VDDA.n214 GNDA 0.155498f
C2784 VDDA.n216 GNDA 0.081762f
C2785 VDDA.n217 GNDA 0.029895f
C2786 VDDA.n218 GNDA 0.106671f
C2787 VDDA.n219 GNDA 0.050691f
C2788 VDDA.t23 GNDA 0.02471f
C2789 VDDA.n220 GNDA 0.087437f
C2790 VDDA.t405 GNDA 0.112738f
C2791 VDDA.n221 GNDA 0.054748f
C2792 VDDA.n222 GNDA 0.053709f
C2793 VDDA.t403 GNDA 0.040912f
C2794 VDDA.n223 GNDA 0.044942f
C2795 VDDA.n224 GNDA 0.036f
C2796 VDDA.n225 GNDA 0.33626f
C2797 VDDA.n226 GNDA 0.335f
C2798 VDDA.t404 GNDA 0.309878f
C2799 VDDA.n227 GNDA 0.048913f
C2800 VDDA.n228 GNDA 0.056716f
C2801 VDDA.n229 GNDA 0.056716f
C2802 VDDA.n230 GNDA 0.102668f
C2803 VDDA.t313 GNDA 0.340032f
C2804 VDDA.t22 GNDA 0.143735f
C2805 VDDA.n231 GNDA 0.025667f
C2806 VDDA.n232 GNDA 0.05955f
C2807 VDDA.n233 GNDA 0.010441f
C2808 VDDA.n234 GNDA 0.035636f
C2809 VDDA.t312 GNDA 0.042935f
C2810 VDDA.n235 GNDA 0.044942f
C2811 VDDA.t314 GNDA 0.088028f
C2812 VDDA.n236 GNDA 0.059194f
C2813 VDDA.n237 GNDA 0.1867f
C2814 VDDA.n238 GNDA 0.115372f
C2815 VDDA.t386 GNDA 0.015441f
C2816 VDDA.n239 GNDA 0.018508f
C2817 VDDA.t384 GNDA 0.013363f
C2818 VDDA.n240 GNDA 0.01883f
C2819 VDDA.n241 GNDA 0.0249f
C2820 VDDA.n242 GNDA 0.165294f
C2821 VDDA.n243 GNDA 0.165294f
C2822 VDDA.t385 GNDA 0.182399f
C2823 VDDA.t391 GNDA 0.182399f
C2824 VDDA.n244 GNDA 0.029895f
C2825 VDDA.n245 GNDA 0.036791f
C2826 VDDA.n246 GNDA 0.036791f
C2827 VDDA.t8 GNDA 0.124037f
C2828 VDDA.n247 GNDA 0.037518f
C2829 VDDA.n248 GNDA 0.010441f
C2830 VDDA.n249 GNDA 0.0249f
C2831 VDDA.t390 GNDA 0.013363f
C2832 VDDA.n250 GNDA 0.01883f
C2833 VDDA.t393 GNDA 0.015441f
C2834 VDDA.n251 GNDA 0.020926f
C2835 VDDA.n252 GNDA 0.122228f
C2836 VDDA.n253 GNDA 0.470112f
C2837 VDDA.n254 GNDA 4.61119f
C2838 VDDA.t470 GNDA 0.769516f
C2839 VDDA.t471 GNDA 0.820156f
C2840 VDDA.t469 GNDA 0.820156f
C2841 VDDA.t472 GNDA 0.786455f
C2842 VDDA.n255 GNDA 0.549754f
C2843 VDDA.n256 GNDA 0.266904f
C2844 VDDA.n257 GNDA 0.342188f
C2845 VDDA.n258 GNDA 2.44178f
C2846 VDDA.n259 GNDA 0.022274f
C2847 VDDA.n260 GNDA 0.016858f
C2848 VDDA.n261 GNDA 0.016858f
C2849 VDDA.n262 GNDA 0.049267f
C2850 VDDA.n263 GNDA 0.022274f
C2851 VDDA.t350 GNDA 0.026148f
C2852 VDDA.t348 GNDA 0.01723f
C2853 VDDA.n264 GNDA 0.041019f
C2854 VDDA.n265 GNDA 0.058365f
C2855 VDDA.n266 GNDA 0.109724f
C2856 VDDA.n267 GNDA 0.109724f
C2857 VDDA.t323 GNDA 0.026148f
C2858 VDDA.t321 GNDA 0.01723f
C2859 VDDA.n268 GNDA 0.041019f
C2860 VDDA.n269 GNDA 0.083526f
C2861 VDDA.n270 GNDA 0.058365f
C2862 VDDA.n271 GNDA 0.022274f
C2863 VDDA.n272 GNDA 0.016858f
C2864 VDDA.n273 GNDA 0.017626f
C2865 VDDA.n274 GNDA 0.017507f
C2866 VDDA.n275 GNDA 0.136095f
C2867 VDDA.n276 GNDA 0.017507f
C2868 VDDA.n277 GNDA 0.070891f
C2869 VDDA.n278 GNDA 0.017507f
C2870 VDDA.n279 GNDA 0.070891f
C2871 VDDA.n280 GNDA 0.016858f
C2872 VDDA.n281 GNDA 0.068467f
C2873 VDDA.n282 GNDA 0.109724f
C2874 VDDA.t365 GNDA 0.026148f
C2875 VDDA.t363 GNDA 0.01723f
C2876 VDDA.n283 GNDA 0.041019f
C2877 VDDA.n284 GNDA 0.058365f
C2878 VDDA.t423 GNDA 0.026148f
C2879 VDDA.t421 GNDA 0.01723f
C2880 VDDA.n285 GNDA 0.041019f
C2881 VDDA.n286 GNDA 0.058365f
C2882 VDDA.n287 GNDA 0.083526f
C2883 VDDA.n288 GNDA 0.109724f
C2884 VDDA.n289 GNDA 0.238571f
C2885 VDDA.t422 GNDA 0.217596f
C2886 VDDA.t50 GNDA 0.137818f
C2887 VDDA.t56 GNDA 0.137818f
C2888 VDDA.t54 GNDA 0.137818f
C2889 VDDA.t155 GNDA 0.137818f
C2890 VDDA.t145 GNDA 0.137818f
C2891 VDDA.t66 GNDA 0.137818f
C2892 VDDA.t96 GNDA 0.137818f
C2893 VDDA.t153 GNDA 0.137818f
C2894 VDDA.t58 GNDA 0.103364f
C2895 VDDA.n290 GNDA 0.068909f
C2896 VDDA.t159 GNDA 0.103364f
C2897 VDDA.t147 GNDA 0.137818f
C2898 VDDA.t100 GNDA 0.137818f
C2899 VDDA.t108 GNDA 0.137818f
C2900 VDDA.t52 GNDA 0.137818f
C2901 VDDA.t437 GNDA 0.137818f
C2902 VDDA.t161 GNDA 0.137818f
C2903 VDDA.t216 GNDA 0.137818f
C2904 VDDA.t64 GNDA 0.137818f
C2905 VDDA.t364 GNDA 0.217596f
C2906 VDDA.n291 GNDA 0.238571f
C2907 VDDA.n292 GNDA 0.068467f
C2908 VDDA.n293 GNDA 0.116636f
C2909 VDDA.n294 GNDA 0.049267f
C2910 VDDA.n295 GNDA 0.022274f
C2911 VDDA.n296 GNDA 0.017507f
C2912 VDDA.n297 GNDA 0.070891f
C2913 VDDA.n298 GNDA 0.017507f
C2914 VDDA.n299 GNDA 0.070891f
C2915 VDDA.n300 GNDA 0.017507f
C2916 VDDA.n301 GNDA 0.070891f
C2917 VDDA.n302 GNDA 0.017507f
C2918 VDDA.n303 GNDA 0.101518f
C2919 VDDA.n304 GNDA 0.022274f
C2920 VDDA.n305 GNDA 0.016858f
C2921 VDDA.n306 GNDA 0.016858f
C2922 VDDA.n307 GNDA 0.049267f
C2923 VDDA.n308 GNDA 0.022274f
C2924 VDDA.n309 GNDA 0.016858f
C2925 VDDA.n310 GNDA 0.022274f
C2926 VDDA.n311 GNDA 0.016858f
C2927 VDDA.n312 GNDA 0.049267f
C2928 VDDA.n313 GNDA 0.022274f
C2929 VDDA.n314 GNDA 0.022274f
C2930 VDDA.n315 GNDA 0.049267f
C2931 VDDA.n316 GNDA 0.022274f
C2932 VDDA.n317 GNDA 0.022274f
C2933 VDDA.n318 GNDA 0.016858f
C2934 VDDA.n319 GNDA 0.049267f
C2935 VDDA.n320 GNDA 0.022274f
C2936 VDDA.n321 GNDA 0.022274f
C2937 VDDA.n322 GNDA 0.049267f
C2938 VDDA.n323 GNDA 0.022274f
C2939 VDDA.n324 GNDA 0.016858f
C2940 VDDA.n325 GNDA 0.049267f
C2941 VDDA.n326 GNDA 0.022274f
C2942 VDDA.n327 GNDA 0.0529f
C2943 VDDA.n328 GNDA 0.049267f
C2944 VDDA.n329 GNDA 0.036366f
C2945 VDDA.n330 GNDA 0.034735f
C2946 VDDA.n331 GNDA 0.238571f
C2947 VDDA.t322 GNDA 0.217596f
C2948 VDDA.t111 GNDA 0.137818f
C2949 VDDA.t36 GNDA 0.137818f
C2950 VDDA.t208 GNDA 0.137818f
C2951 VDDA.t458 GNDA 0.137818f
C2952 VDDA.t170 GNDA 0.137818f
C2953 VDDA.t60 GNDA 0.137818f
C2954 VDDA.t120 GNDA 0.137818f
C2955 VDDA.t77 GNDA 0.137818f
C2956 VDDA.t34 GNDA 0.103364f
C2957 VDDA.n332 GNDA 0.068909f
C2958 VDDA.t38 GNDA 0.103364f
C2959 VDDA.t24 GNDA 0.137818f
C2960 VDDA.t433 GNDA 0.137818f
C2961 VDDA.t199 GNDA 0.137818f
C2962 VDDA.t206 GNDA 0.137818f
C2963 VDDA.t75 GNDA 0.137818f
C2964 VDDA.t124 GNDA 0.137818f
C2965 VDDA.t183 GNDA 0.137818f
C2966 VDDA.t46 GNDA 0.137818f
C2967 VDDA.t349 GNDA 0.217596f
C2968 VDDA.n333 GNDA 0.238571f
C2969 VDDA.n334 GNDA 0.034735f
C2970 VDDA.n335 GNDA 0.036366f
C2971 VDDA.n336 GNDA 0.049267f
C2972 VDDA.n337 GNDA 0.067432f
C2973 VDDA.n338 GNDA 0.204725f
C2974 VDDA.t287 GNDA 0.020882f
C2975 VDDA.t285 GNDA 0.020882f
C2976 VDDA.n339 GNDA 0.068986f
C2977 VDDA.n340 GNDA 0.089018f
C2978 VDDA.t389 GNDA 0.063993f
C2979 VDDA.n341 GNDA 0.112761f
C2980 VDDA.n342 GNDA 0.153714f
C2981 VDDA.n343 GNDA 0.153714f
C2982 VDDA.n344 GNDA 0.153008f
C2983 VDDA.t344 GNDA 0.063993f
C2984 VDDA.t342 GNDA 0.099572f
C2985 VDDA.t383 GNDA 0.026148f
C2986 VDDA.t381 GNDA 0.013196f
C2987 VDDA.n345 GNDA 0.041225f
C2988 VDDA.n346 GNDA 0.023771f
C2989 VDDA.n347 GNDA 0.042247f
C2990 VDDA.t411 GNDA 0.026148f
C2991 VDDA.t409 GNDA 0.013196f
C2992 VDDA.n348 GNDA 0.041225f
C2993 VDDA.n349 GNDA 0.042247f
C2994 VDDA.n350 GNDA 0.042247f
C2995 VDDA.n351 GNDA 0.034664f
C2996 VDDA.n352 GNDA 0.166574f
C2997 VDDA.t382 GNDA 0.209159f
C2998 VDDA.t429 GNDA 0.09475f
C2999 VDDA.n353 GNDA 0.063167f
C3000 VDDA.t430 GNDA 0.09475f
C3001 VDDA.t410 GNDA 0.212243f
C3002 VDDA.n354 GNDA 0.174974f
C3003 VDDA.n355 GNDA 0.034664f
C3004 VDDA.n356 GNDA 0.023771f
C3005 VDDA.n357 GNDA 0.033396f
C3006 VDDA.t306 GNDA 0.020882f
C3007 VDDA.t267 GNDA 0.020882f
C3008 VDDA.n358 GNDA 0.068986f
C3009 VDDA.n359 GNDA 0.089018f
C3010 VDDA.t279 GNDA 0.020882f
C3011 VDDA.t297 GNDA 0.020882f
C3012 VDDA.n360 GNDA 0.068986f
C3013 VDDA.n361 GNDA 0.089018f
C3014 VDDA.t262 GNDA 0.020882f
C3015 VDDA.t281 GNDA 0.020882f
C3016 VDDA.n362 GNDA 0.068986f
C3017 VDDA.n363 GNDA 0.089018f
C3018 VDDA.t295 GNDA 0.020882f
C3019 VDDA.t303 GNDA 0.020882f
C3020 VDDA.n364 GNDA 0.068986f
C3021 VDDA.n365 GNDA 0.089018f
C3022 VDDA.t276 GNDA 0.020882f
C3023 VDDA.t272 GNDA 0.020882f
C3024 VDDA.n366 GNDA 0.068986f
C3025 VDDA.n367 GNDA 0.089018f
C3026 VDDA.t301 GNDA 0.020882f
C3027 VDDA.t311 GNDA 0.020882f
C3028 VDDA.n368 GNDA 0.068986f
C3029 VDDA.n369 GNDA 0.089018f
C3030 VDDA.t269 GNDA 0.020882f
C3031 VDDA.t290 GNDA 0.020882f
C3032 VDDA.n370 GNDA 0.068986f
C3033 VDDA.n371 GNDA 0.089018f
C3034 VDDA.n372 GNDA 0.098286f
C3035 VDDA.n373 GNDA 0.118836f
C3036 VDDA.n374 GNDA 0.080101f
C3037 VDDA.n375 GNDA 0.097797f
C3038 VDDA.n376 GNDA 0.360336f
C3039 VDDA.t343 GNDA 0.464953f
C3040 VDDA.t268 GNDA 0.335149f
C3041 VDDA.t289 GNDA 0.335149f
C3042 VDDA.t300 GNDA 0.335149f
C3043 VDDA.t310 GNDA 0.335149f
C3044 VDDA.t275 GNDA 0.335149f
C3045 VDDA.t271 GNDA 0.335149f
C3046 VDDA.t294 GNDA 0.335149f
C3047 VDDA.t302 GNDA 0.251362f
C3048 VDDA.n377 GNDA 0.167575f
C3049 VDDA.t261 GNDA 0.251362f
C3050 VDDA.t280 GNDA 0.335149f
C3051 VDDA.t278 GNDA 0.335149f
C3052 VDDA.t296 GNDA 0.335149f
C3053 VDDA.t305 GNDA 0.335149f
C3054 VDDA.t266 GNDA 0.335149f
C3055 VDDA.t286 GNDA 0.335149f
C3056 VDDA.t284 GNDA 0.335149f
C3057 VDDA.t388 GNDA 0.464953f
C3058 VDDA.n378 GNDA 0.360336f
C3059 VDDA.n379 GNDA 0.097797f
C3060 VDDA.n380 GNDA 0.080101f
C3061 VDDA.t387 GNDA 0.099572f
C3062 VDDA.n381 GNDA 0.118836f
C3063 VDDA.n382 GNDA 0.05455f
C3064 VDDA.n383 GNDA 0.016811f
C3065 VDDA.t335 GNDA 0.026342f
C3066 VDDA.t333 GNDA 0.012854f
C3067 VDDA.n384 GNDA 0.039458f
C3068 VDDA.n385 GNDA 0.023662f
C3069 VDDA.n386 GNDA 0.042247f
C3070 VDDA.t332 GNDA 0.026342f
C3071 VDDA.t330 GNDA 0.012854f
C3072 VDDA.n387 GNDA 0.039458f
C3073 VDDA.n388 GNDA 0.042247f
C3074 VDDA.n389 GNDA 0.042247f
C3075 VDDA.n390 GNDA 0.034664f
C3076 VDDA.n391 GNDA 0.166574f
C3077 VDDA.t334 GNDA 0.209159f
C3078 VDDA.t106 GNDA 0.09475f
C3079 VDDA.n392 GNDA 0.063167f
C3080 VDDA.t445 GNDA 0.09475f
C3081 VDDA.t331 GNDA 0.209159f
C3082 VDDA.n393 GNDA 0.166574f
C3083 VDDA.n394 GNDA 0.034664f
C3084 VDDA.n395 GNDA 0.023662f
C3085 VDDA.n396 GNDA 0.024859f
C3086 VDDA.n397 GNDA 0.04653f
C3087 VDDA.n398 GNDA 0.098034f
C3088 VDDA.n399 GNDA 0.170233f
C3089 VDDA.n400 GNDA 0.017363f
C3090 VDDA.n401 GNDA 0.061291f
C3091 VDDA.t338 GNDA 0.02747f
C3092 VDDA.n402 GNDA 0.02297f
C3093 VDDA.n403 GNDA 0.049718f
C3094 VDDA.n404 GNDA 0.049718f
C3095 VDDA.n405 GNDA 0.049718f
C3096 VDDA.t399 GNDA 0.02747f
C3097 VDDA.t397 GNDA 0.013708f
C3098 VDDA.n406 GNDA 0.017331f
C3099 VDDA.n407 GNDA 0.061323f
C3100 VDDA.t414 GNDA 0.026215f
C3101 VDDA.n408 GNDA 0.04594f
C3102 VDDA.n409 GNDA 0.079961f
C3103 VDDA.n410 GNDA 0.079961f
C3104 VDDA.n411 GNDA 0.079961f
C3105 VDDA.t420 GNDA 0.026215f
C3106 VDDA.t418 GNDA 0.013708f
C3107 VDDA.n412 GNDA 0.01737f
C3108 VDDA.n413 GNDA 0.061284f
C3109 VDDA.t374 GNDA 0.027481f
C3110 VDDA.n414 GNDA 0.02297f
C3111 VDDA.n415 GNDA 0.049718f
C3112 VDDA.n416 GNDA 0.049718f
C3113 VDDA.n417 GNDA 0.049718f
C3114 VDDA.t317 GNDA 0.027481f
C3115 VDDA.t315 GNDA 0.013708f
C3116 VDDA.n418 GNDA 0.01737f
C3117 VDDA.n419 GNDA 0.083877f
C3118 VDDA.n420 GNDA 0.047064f
C3119 VDDA.n421 GNDA 0.028087f
C3120 VDDA.n422 GNDA 0.038585f
C3121 VDDA.n423 GNDA 0.175784f
C3122 VDDA.t316 GNDA 0.212838f
C3123 VDDA.t142 GNDA 0.128248f
C3124 VDDA.t71 GNDA 0.096186f
C3125 VDDA.n424 GNDA 0.064124f
C3126 VDDA.t461 GNDA 0.096186f
C3127 VDDA.t113 GNDA 0.128248f
C3128 VDDA.t373 GNDA 0.212838f
C3129 VDDA.n425 GNDA 0.175784f
C3130 VDDA.n426 GNDA 0.038585f
C3131 VDDA.n427 GNDA 0.028087f
C3132 VDDA.t372 GNDA 0.014143f
C3133 VDDA.n428 GNDA 0.046578f
C3134 VDDA.n429 GNDA 0.042308f
C3135 VDDA.n430 GNDA 0.017331f
C3136 VDDA.n431 GNDA 0.061323f
C3137 VDDA.n432 GNDA 0.017331f
C3138 VDDA.n433 GNDA 0.061323f
C3139 VDDA.n434 GNDA 0.017331f
C3140 VDDA.n435 GNDA 0.061323f
C3141 VDDA.n436 GNDA 0.017331f
C3142 VDDA.n437 GNDA 0.061323f
C3143 VDDA.n438 GNDA 0.042308f
C3144 VDDA.n439 GNDA 0.04741f
C3145 VDDA.n440 GNDA 0.0434f
C3146 VDDA.n441 GNDA 0.05409f
C3147 VDDA.n442 GNDA 0.206794f
C3148 VDDA.t419 GNDA 0.212838f
C3149 VDDA.t73 GNDA 0.128248f
C3150 VDDA.t454 GNDA 0.128248f
C3151 VDDA.t181 GNDA 0.128248f
C3152 VDDA.t48 GNDA 0.128248f
C3153 VDDA.t140 GNDA 0.128248f
C3154 VDDA.t202 GNDA 0.096186f
C3155 VDDA.n443 GNDA 0.064124f
C3156 VDDA.t94 GNDA 0.096186f
C3157 VDDA.t16 GNDA 0.128248f
C3158 VDDA.t179 GNDA 0.128248f
C3159 VDDA.t91 GNDA 0.128248f
C3160 VDDA.t413 GNDA 0.336941f
C3161 VDDA.n444 GNDA 0.339185f
C3162 VDDA.n445 GNDA 0.062098f
C3163 VDDA.n446 GNDA 0.043049f
C3164 VDDA.t412 GNDA 0.013708f
C3165 VDDA.n447 GNDA 0.04741f
C3166 VDDA.n448 GNDA 0.049965f
C3167 VDDA.n449 GNDA 0.017363f
C3168 VDDA.n450 GNDA 0.061291f
C3169 VDDA.n451 GNDA 0.049965f
C3170 VDDA.n452 GNDA 0.046154f
C3171 VDDA.n453 GNDA 0.028087f
C3172 VDDA.n454 GNDA 0.038052f
C3173 VDDA.n455 GNDA 0.173883f
C3174 VDDA.t398 GNDA 0.209159f
C3175 VDDA.t164 GNDA 0.126334f
C3176 VDDA.t115 GNDA 0.086136f
C3177 VDDA.n456 GNDA 0.031583f
C3178 VDDA.n457 GNDA 0.040197f
C3179 VDDA.t449 GNDA 0.09475f
C3180 VDDA.t204 GNDA 0.126334f
C3181 VDDA.t337 GNDA 0.209159f
C3182 VDDA.n458 GNDA 0.174949f
C3183 VDDA.n459 GNDA 0.039118f
C3184 VDDA.n460 GNDA 0.028087f
C3185 VDDA.t336 GNDA 0.013708f
C3186 VDDA.n461 GNDA 0.046154f
C3187 VDDA.n462 GNDA 0.092057f
C3188 VDDA.n463 GNDA 0.138185f
C3189 VDDA.t299 GNDA 0.389094f
C3190 VDDA.t307 GNDA 0.390504f
C3191 VDDA.t277 GNDA 0.389094f
C3192 VDDA.t263 GNDA 0.390504f
C3193 VDDA.t288 GNDA 0.389094f
C3194 VDDA.t292 GNDA 0.390504f
C3195 VDDA.t264 GNDA 0.389094f
C3196 VDDA.t304 GNDA 0.390504f
C3197 VDDA.t293 GNDA 0.389094f
C3198 VDDA.t309 GNDA 0.390504f
C3199 VDDA.t282 GNDA 0.389094f
C3200 VDDA.t265 GNDA 0.390504f
C3201 VDDA.t260 GNDA 0.389094f
C3202 VDDA.t274 GNDA 0.390504f
C3203 VDDA.t298 GNDA 0.389094f
C3204 VDDA.t283 GNDA 0.390504f
C3205 VDDA.n464 GNDA 0.26081f
C3206 VDDA.t291 GNDA 0.207697f
C3207 VDDA.n465 GNDA 0.282985f
C3208 VDDA.t273 GNDA 0.207697f
C3209 VDDA.n466 GNDA 0.282985f
C3210 VDDA.t308 GNDA 0.207697f
C3211 VDDA.n467 GNDA 0.282985f
C3212 VDDA.t270 GNDA 0.309925f
C3213 VDDA.n468 GNDA 0.270061f
C3214 VDDA.n469 GNDA 0.853205f
C3215 bgr_0.Vin-.n0 GNDA 0.073641f
C3216 bgr_0.Vin-.n1 GNDA 0.082742f
C3217 bgr_0.Vin-.n2 GNDA 0.998979f
C3218 bgr_0.Vin-.t5 GNDA 0.028614f
C3219 bgr_0.Vin-.t4 GNDA 0.028614f
C3220 bgr_0.Vin-.n3 GNDA 0.099613f
C3221 bgr_0.Vin-.t3 GNDA 0.028614f
C3222 bgr_0.Vin-.t2 GNDA 0.028614f
C3223 bgr_0.Vin-.n4 GNDA 0.095121f
C3224 bgr_0.Vin-.n5 GNDA 0.408067f
C3225 bgr_0.Vin-.t1 GNDA 0.098662f
C3226 bgr_0.Vin-.n6 GNDA 0.025702f
C3227 bgr_0.Vin-.n7 GNDA 0.469862f
C3228 bgr_0.Vin-.n8 GNDA 0.222852f
C3229 bgr_0.Vin-.t10 GNDA 0.023594f
C3230 bgr_0.Vin-.n9 GNDA 0.027673f
C3231 bgr_0.Vin-.n10 GNDA 0.022653f
C3232 bgr_0.Vin-.n11 GNDA 0.022653f
C3233 bgr_0.Vin-.n12 GNDA 0.040466f
C3234 bgr_0.Vin-.n13 GNDA 0.524007f
C3235 bgr_0.Vin-.t0 GNDA 0.276208f
C3236 bgr_0.Vin-.n14 GNDA 0.510829f
C3237 bgr_0.Vin-.n15 GNDA 0.074468f
C3238 bgr_0.Vin-.n16 GNDA 0.126176f
C3239 bgr_0.Vin-.n17 GNDA 0.073776f
C3240 bgr_0.Vin-.n18 GNDA 0.145931f
C3241 bgr_0.Vin-.n19 GNDA 0.145931f
C3242 bgr_0.Vin-.n20 GNDA -5.06787f
C3243 bgr_0.Vin-.n21 GNDA 5.25363f
C3244 bgr_0.Vin-.n22 GNDA 0.222489f
C3245 bgr_0.Vin-.n23 GNDA 0.382836f
C3246 bgr_0.Vin-.n24 GNDA 0.166915f
C3247 bgr_0.Vin-.n25 GNDA 0.040544f
C3248 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.043026f
C3249 bgr_0.V_TOP.t31 GNDA 0.115045f
C3250 bgr_0.V_TOP.t44 GNDA 0.115045f
C3251 bgr_0.V_TOP.t18 GNDA 0.115045f
C3252 bgr_0.V_TOP.t26 GNDA 0.115045f
C3253 bgr_0.V_TOP.t37 GNDA 0.115045f
C3254 bgr_0.V_TOP.t35 GNDA 0.115045f
C3255 bgr_0.V_TOP.t48 GNDA 0.115045f
C3256 bgr_0.V_TOP.t20 GNDA 0.115045f
C3257 bgr_0.V_TOP.t27 GNDA 0.115045f
C3258 bgr_0.V_TOP.t41 GNDA 0.115045f
C3259 bgr_0.V_TOP.t38 GNDA 0.115045f
C3260 bgr_0.V_TOP.t14 GNDA 0.115045f
C3261 bgr_0.V_TOP.t23 GNDA 0.115045f
C3262 bgr_0.V_TOP.t29 GNDA 0.115045f
C3263 bgr_0.V_TOP.t43 GNDA 0.150392f
C3264 bgr_0.V_TOP.n0 GNDA 0.084081f
C3265 bgr_0.V_TOP.n1 GNDA 0.061357f
C3266 bgr_0.V_TOP.n2 GNDA 0.061357f
C3267 bgr_0.V_TOP.n3 GNDA 0.061357f
C3268 bgr_0.V_TOP.n4 GNDA 0.061357f
C3269 bgr_0.V_TOP.n5 GNDA 0.057217f
C3270 bgr_0.V_TOP.t7 GNDA 0.147947f
C3271 bgr_0.V_TOP.t13 GNDA 0.155772f
C3272 bgr_0.V_TOP.t0 GNDA 0.010957f
C3273 bgr_0.V_TOP.t1 GNDA 0.010957f
C3274 bgr_0.V_TOP.n6 GNDA 0.027281f
C3275 bgr_0.V_TOP.n7 GNDA 0.726844f
C3276 bgr_0.V_TOP.t3 GNDA 0.010957f
C3277 bgr_0.V_TOP.t4 GNDA 0.010957f
C3278 bgr_0.V_TOP.n8 GNDA 0.026425f
C3279 bgr_0.V_TOP.t8 GNDA 0.010957f
C3280 bgr_0.V_TOP.t11 GNDA 0.010957f
C3281 bgr_0.V_TOP.n9 GNDA 0.027465f
C3282 bgr_0.V_TOP.t12 GNDA 0.010957f
C3283 bgr_0.V_TOP.t9 GNDA 0.010957f
C3284 bgr_0.V_TOP.n10 GNDA 0.027281f
C3285 bgr_0.V_TOP.n11 GNDA 0.252824f
C3286 bgr_0.V_TOP.n12 GNDA 0.153577f
C3287 bgr_0.V_TOP.n13 GNDA 0.087653f
C3288 bgr_0.V_TOP.t5 GNDA 0.010957f
C3289 bgr_0.V_TOP.t6 GNDA 0.010957f
C3290 bgr_0.V_TOP.n14 GNDA 0.027281f
C3291 bgr_0.V_TOP.n15 GNDA 0.151313f
C3292 bgr_0.V_TOP.t2 GNDA 0.010957f
C3293 bgr_0.V_TOP.t10 GNDA 0.010957f
C3294 bgr_0.V_TOP.n16 GNDA 0.027281f
C3295 bgr_0.V_TOP.n17 GNDA 0.149874f
C3296 bgr_0.V_TOP.n18 GNDA 0.329448f
C3297 bgr_0.V_TOP.n19 GNDA 0.023183f
C3298 bgr_0.V_TOP.n20 GNDA 0.057217f
C3299 bgr_0.V_TOP.n21 GNDA 0.061357f
C3300 bgr_0.V_TOP.n22 GNDA 0.061357f
C3301 bgr_0.V_TOP.n23 GNDA 0.061357f
C3302 bgr_0.V_TOP.n24 GNDA 0.061357f
C3303 bgr_0.V_TOP.n25 GNDA 0.061357f
C3304 bgr_0.V_TOP.n26 GNDA 0.061357f
C3305 bgr_0.V_TOP.n27 GNDA 0.057217f
C3306 bgr_0.V_TOP.t32 GNDA 0.132572f
C3307 bgr_0.V_TOP.t49 GNDA 0.445732f
C3308 bgr_0.V_TOP.t39 GNDA 0.438267f
C3309 bgr_0.V_TOP.n28 GNDA 0.293844f
C3310 bgr_0.V_TOP.t28 GNDA 0.438267f
C3311 bgr_0.V_TOP.t25 GNDA 0.445732f
C3312 bgr_0.V_TOP.t33 GNDA 0.438267f
C3313 bgr_0.V_TOP.n29 GNDA 0.293844f
C3314 bgr_0.V_TOP.n30 GNDA 0.273917f
C3315 bgr_0.V_TOP.t21 GNDA 0.445732f
C3316 bgr_0.V_TOP.t15 GNDA 0.438267f
C3317 bgr_0.V_TOP.n31 GNDA 0.293844f
C3318 bgr_0.V_TOP.t40 GNDA 0.438267f
C3319 bgr_0.V_TOP.t34 GNDA 0.445732f
C3320 bgr_0.V_TOP.t45 GNDA 0.438267f
C3321 bgr_0.V_TOP.n32 GNDA 0.293844f
C3322 bgr_0.V_TOP.n33 GNDA 0.356092f
C3323 bgr_0.V_TOP.t30 GNDA 0.445732f
C3324 bgr_0.V_TOP.t22 GNDA 0.438267f
C3325 bgr_0.V_TOP.n34 GNDA 0.293844f
C3326 bgr_0.V_TOP.t16 GNDA 0.438267f
C3327 bgr_0.V_TOP.t46 GNDA 0.445732f
C3328 bgr_0.V_TOP.t19 GNDA 0.438267f
C3329 bgr_0.V_TOP.n35 GNDA 0.293844f
C3330 bgr_0.V_TOP.n36 GNDA 0.356092f
C3331 bgr_0.V_TOP.t24 GNDA 0.445732f
C3332 bgr_0.V_TOP.t17 GNDA 0.438267f
C3333 bgr_0.V_TOP.n37 GNDA 0.293844f
C3334 bgr_0.V_TOP.t42 GNDA 0.438267f
C3335 bgr_0.V_TOP.n38 GNDA 0.273917f
C3336 bgr_0.V_TOP.t47 GNDA 0.438267f
C3337 bgr_0.V_TOP.n39 GNDA 0.191742f
C3338 bgr_0.V_TOP.t36 GNDA 0.438267f
C3339 bgr_0.V_TOP.n40 GNDA 0.893239f
.ends

