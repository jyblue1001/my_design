* NGSPICE file created from B.ext - technology: sky130A

**.subckt B
X0 a_4510_n8350# p_right a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X1 w_5530_n8860# p_bias v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X2 p_left a_4510_n7380# v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X3 a_4510_n8350# n_right w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 n_right VOUT v_common_n a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X5 v_common_p p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X6 a_5700_n9470# p_right a_4510_n8350# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X7 p_right p_left a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X8 p_bias n_bias a_5700_n9470# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X9 v_common_p p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X10 w_5530_n8860# n_right a_4510_n8350# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X11 v_common_n VOUT n_right a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X12 w_5530_n8860# p_bias p_bias w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X13 a_5700_n9470# p_left p_right a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X14 a_4510_n8350# a_8196_n10872# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X15 n_right n_left w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X16 p_left p_left a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X17 n_left a_4510_n7380# v_common_n a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X18 w_5530_n8860# p_bias p_bias w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 a_4510_n8350# n_right w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X20 v_common_n n_bias a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X21 w_5530_n8860# n_left n_right w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X22 a_5700_n9470# n_bias n_bias a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X23 v_common_p a_4510_n7380# p_left w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X24 w_5530_n8860# n_right a_4510_n8350# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X25 a_5700_n9470# p_left p_left a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X26 a_4510_n8350# a_5270_n10872# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X27 p_bias p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X28 a_4510_n8350# p_right a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X29 n_right a_8196_n10872# a_5700_n9470# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X30 n_left n_left w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X31 p_right VOUT v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X32 p_bias p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X33 a_5270_n10872# p_right a_5700_n9470# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X34 w_5530_n8860# p_bias v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X35 v_common_p VOUT p_right w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X36 w_5530_n8860# n_left n_left w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X37 a_5700_n9470# p_right a_4510_n8350# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X38 n_bias n_bias a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X39 a_5700_n9470# n_bias v_common_n a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X40 v_common_n a_4510_n7380# n_left a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
**.ends

