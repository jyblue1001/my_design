** sch_path: /foss/designs/my_design/projects/montecarlo/xschem_ngspice/inverter/inverter_monte_carlo.sch
**.subckt inverter_monte_carlo
XM1 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdd VDD GND 1.8
Vin Vin GND 0.5
**** begin user architecture code



.option wnflag=1

.control

  let runs=10
  let run=1

  dowhile run <= runs
    save all
    dc vin 0 1.8 0.01
    write inverter_monte_carlo_mc.raw
    set appendwrite
    reset
    let run = run + 1
  end

.endc




.param mc_mm_switch=0
.param mc_pr_switch=1
.include /foss/pdks/sky130A/libs.tech/ngspice/parameters/critical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/parameters/montecarlo.spice

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
