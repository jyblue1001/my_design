magic
tech sky130A
timestamp 1756186613
<< nwell >>
rect 16915 520 17735 660
rect 17865 520 18685 660
rect 16375 120 16760 260
rect 16910 20 18690 360
rect 16360 -560 17725 -420
rect 17875 -560 19240 -420
<< pwell >>
rect 17780 -4275 17820 -4120
<< nmos >>
rect 17000 -1055 17020 -805
rect 17060 -1055 17080 -805
rect 18520 -1055 18540 -805
rect 18580 -1055 18600 -805
rect 16570 -1565 17070 -1315
rect 17190 -1565 17690 -1315
rect 17910 -1565 18410 -1315
rect 18530 -1565 19030 -1315
rect 16780 -1870 17780 -1770
rect 17820 -1870 18820 -1770
<< pmos >>
rect 17015 540 17030 640
rect 17070 540 17085 640
rect 17125 540 17140 640
rect 17180 540 17195 640
rect 17235 540 17250 640
rect 17290 540 17305 640
rect 17345 540 17360 640
rect 17400 540 17415 640
rect 17455 540 17470 640
rect 17510 540 17525 640
rect 17565 540 17580 640
rect 17620 540 17635 640
rect 17965 540 17980 640
rect 18020 540 18035 640
rect 18075 540 18090 640
rect 18130 540 18145 640
rect 18185 540 18200 640
rect 18240 540 18255 640
rect 18295 540 18310 640
rect 18350 540 18365 640
rect 18405 540 18420 640
rect 18460 540 18475 640
rect 18515 540 18530 640
rect 18570 540 18585 640
rect 16475 140 16490 240
rect 16530 140 16545 240
rect 16585 140 16600 240
rect 16640 140 16655 240
rect 17010 40 17060 340
rect 17100 40 17150 340
rect 17190 40 17240 340
rect 17280 40 17330 340
rect 17370 40 17420 340
rect 17460 40 17510 340
rect 17550 40 17600 340
rect 17640 40 17690 340
rect 17730 40 17780 340
rect 17820 40 17870 340
rect 17910 40 17960 340
rect 18000 40 18050 340
rect 18090 40 18140 340
rect 18180 40 18230 340
rect 18270 40 18320 340
rect 18360 40 18410 340
rect 18450 40 18500 340
rect 18540 40 18590 340
rect 16460 -540 16480 -440
rect 16520 -540 16540 -440
rect 16580 -540 16600 -440
rect 16640 -540 16660 -440
rect 16700 -540 16720 -440
rect 16760 -540 16780 -440
rect 16820 -540 16840 -440
rect 16880 -540 16900 -440
rect 16940 -540 16960 -440
rect 17000 -540 17020 -440
rect 17060 -540 17080 -440
rect 17120 -540 17140 -440
rect 17180 -540 17200 -440
rect 17240 -540 17260 -440
rect 17300 -540 17320 -440
rect 17360 -540 17380 -440
rect 17420 -540 17440 -440
rect 17480 -540 17500 -440
rect 17540 -540 17560 -440
rect 17600 -540 17620 -440
rect 17980 -540 18000 -440
rect 18040 -540 18060 -440
rect 18100 -540 18120 -440
rect 18160 -540 18180 -440
rect 18220 -540 18240 -440
rect 18280 -540 18300 -440
rect 18340 -540 18360 -440
rect 18400 -540 18420 -440
rect 18460 -540 18480 -440
rect 18520 -540 18540 -440
rect 18580 -540 18600 -440
rect 18640 -540 18660 -440
rect 18700 -540 18720 -440
rect 18760 -540 18780 -440
rect 18820 -540 18840 -440
rect 18880 -540 18900 -440
rect 18940 -540 18960 -440
rect 19000 -540 19020 -440
rect 19060 -540 19080 -440
rect 19120 -540 19140 -440
<< ndiff >>
rect 16960 -820 17000 -805
rect 16960 -840 16970 -820
rect 16990 -840 17000 -820
rect 16960 -870 17000 -840
rect 16960 -890 16970 -870
rect 16990 -890 17000 -870
rect 16960 -920 17000 -890
rect 16960 -940 16970 -920
rect 16990 -940 17000 -920
rect 16960 -970 17000 -940
rect 16960 -990 16970 -970
rect 16990 -990 17000 -970
rect 16960 -1020 17000 -990
rect 16960 -1040 16970 -1020
rect 16990 -1040 17000 -1020
rect 16960 -1055 17000 -1040
rect 17020 -820 17060 -805
rect 17020 -840 17030 -820
rect 17050 -840 17060 -820
rect 17020 -870 17060 -840
rect 17020 -890 17030 -870
rect 17050 -890 17060 -870
rect 17020 -920 17060 -890
rect 17020 -940 17030 -920
rect 17050 -940 17060 -920
rect 17020 -970 17060 -940
rect 17020 -990 17030 -970
rect 17050 -990 17060 -970
rect 17020 -1020 17060 -990
rect 17020 -1040 17030 -1020
rect 17050 -1040 17060 -1020
rect 17020 -1055 17060 -1040
rect 17080 -820 17120 -805
rect 17080 -840 17090 -820
rect 17110 -840 17120 -820
rect 17080 -870 17120 -840
rect 17080 -890 17090 -870
rect 17110 -890 17120 -870
rect 17080 -920 17120 -890
rect 17080 -940 17090 -920
rect 17110 -940 17120 -920
rect 18480 -820 18520 -805
rect 18480 -840 18490 -820
rect 18510 -840 18520 -820
rect 18480 -870 18520 -840
rect 18480 -890 18490 -870
rect 18510 -890 18520 -870
rect 18480 -920 18520 -890
rect 17080 -970 17120 -940
rect 17080 -990 17090 -970
rect 17110 -990 17120 -970
rect 17080 -1020 17120 -990
rect 17080 -1040 17090 -1020
rect 17110 -1040 17120 -1020
rect 17080 -1055 17120 -1040
rect 18480 -940 18490 -920
rect 18510 -940 18520 -920
rect 18480 -970 18520 -940
rect 18480 -990 18490 -970
rect 18510 -990 18520 -970
rect 18480 -1020 18520 -990
rect 18480 -1040 18490 -1020
rect 18510 -1040 18520 -1020
rect 18480 -1055 18520 -1040
rect 18540 -820 18580 -805
rect 18540 -840 18550 -820
rect 18570 -840 18580 -820
rect 18540 -870 18580 -840
rect 18540 -890 18550 -870
rect 18570 -890 18580 -870
rect 18540 -920 18580 -890
rect 18540 -940 18550 -920
rect 18570 -940 18580 -920
rect 18540 -970 18580 -940
rect 18540 -990 18550 -970
rect 18570 -990 18580 -970
rect 18540 -1020 18580 -990
rect 18540 -1040 18550 -1020
rect 18570 -1040 18580 -1020
rect 18540 -1055 18580 -1040
rect 18600 -820 18640 -805
rect 18600 -840 18610 -820
rect 18630 -840 18640 -820
rect 18600 -870 18640 -840
rect 18600 -890 18610 -870
rect 18630 -890 18640 -870
rect 18600 -920 18640 -890
rect 18600 -940 18610 -920
rect 18630 -940 18640 -920
rect 18600 -970 18640 -940
rect 18600 -990 18610 -970
rect 18630 -990 18640 -970
rect 18600 -1020 18640 -990
rect 18600 -1040 18610 -1020
rect 18630 -1040 18640 -1020
rect 18600 -1055 18640 -1040
rect 16530 -1330 16570 -1315
rect 16530 -1350 16540 -1330
rect 16560 -1350 16570 -1330
rect 16530 -1380 16570 -1350
rect 16530 -1400 16540 -1380
rect 16560 -1400 16570 -1380
rect 16530 -1430 16570 -1400
rect 16530 -1450 16540 -1430
rect 16560 -1450 16570 -1430
rect 16530 -1480 16570 -1450
rect 16530 -1500 16540 -1480
rect 16560 -1500 16570 -1480
rect 16530 -1530 16570 -1500
rect 16530 -1550 16540 -1530
rect 16560 -1550 16570 -1530
rect 16530 -1565 16570 -1550
rect 17070 -1330 17110 -1315
rect 17150 -1330 17190 -1315
rect 17070 -1350 17080 -1330
rect 17100 -1350 17110 -1330
rect 17150 -1350 17160 -1330
rect 17180 -1350 17190 -1330
rect 17070 -1380 17110 -1350
rect 17150 -1380 17190 -1350
rect 17070 -1400 17080 -1380
rect 17100 -1400 17110 -1380
rect 17150 -1400 17160 -1380
rect 17180 -1400 17190 -1380
rect 17070 -1430 17110 -1400
rect 17150 -1430 17190 -1400
rect 17070 -1450 17080 -1430
rect 17100 -1450 17110 -1430
rect 17150 -1450 17160 -1430
rect 17180 -1450 17190 -1430
rect 17070 -1480 17110 -1450
rect 17150 -1480 17190 -1450
rect 17070 -1500 17080 -1480
rect 17100 -1500 17110 -1480
rect 17150 -1500 17160 -1480
rect 17180 -1500 17190 -1480
rect 17070 -1530 17110 -1500
rect 17150 -1530 17190 -1500
rect 17070 -1550 17080 -1530
rect 17100 -1550 17110 -1530
rect 17150 -1550 17160 -1530
rect 17180 -1550 17190 -1530
rect 17070 -1560 17110 -1550
rect 17150 -1560 17190 -1550
rect 17070 -1565 17190 -1560
rect 17690 -1330 17730 -1315
rect 17690 -1350 17700 -1330
rect 17720 -1350 17730 -1330
rect 17690 -1380 17730 -1350
rect 17690 -1400 17700 -1380
rect 17720 -1400 17730 -1380
rect 17690 -1430 17730 -1400
rect 17690 -1450 17700 -1430
rect 17720 -1450 17730 -1430
rect 17690 -1480 17730 -1450
rect 17690 -1500 17700 -1480
rect 17720 -1500 17730 -1480
rect 17690 -1530 17730 -1500
rect 17690 -1550 17700 -1530
rect 17720 -1550 17730 -1530
rect 17690 -1565 17730 -1550
rect 17870 -1330 17910 -1315
rect 17870 -1350 17880 -1330
rect 17900 -1350 17910 -1330
rect 17870 -1380 17910 -1350
rect 17870 -1400 17880 -1380
rect 17900 -1400 17910 -1380
rect 17870 -1430 17910 -1400
rect 17870 -1450 17880 -1430
rect 17900 -1450 17910 -1430
rect 17870 -1480 17910 -1450
rect 17870 -1500 17880 -1480
rect 17900 -1500 17910 -1480
rect 17870 -1530 17910 -1500
rect 17870 -1550 17880 -1530
rect 17900 -1550 17910 -1530
rect 17870 -1565 17910 -1550
rect 18410 -1330 18450 -1315
rect 18490 -1330 18530 -1315
rect 18410 -1350 18420 -1330
rect 18440 -1350 18450 -1330
rect 18490 -1350 18500 -1330
rect 18520 -1350 18530 -1330
rect 18410 -1380 18450 -1350
rect 18490 -1380 18530 -1350
rect 18410 -1400 18420 -1380
rect 18440 -1400 18450 -1380
rect 18490 -1400 18500 -1380
rect 18520 -1400 18530 -1380
rect 18410 -1430 18450 -1400
rect 18490 -1430 18530 -1400
rect 18410 -1450 18420 -1430
rect 18440 -1450 18450 -1430
rect 18490 -1450 18500 -1430
rect 18520 -1450 18530 -1430
rect 18410 -1480 18450 -1450
rect 18490 -1480 18530 -1450
rect 18410 -1500 18420 -1480
rect 18440 -1500 18450 -1480
rect 18490 -1500 18500 -1480
rect 18520 -1500 18530 -1480
rect 18410 -1530 18450 -1500
rect 18490 -1530 18530 -1500
rect 18410 -1550 18420 -1530
rect 18440 -1550 18450 -1530
rect 18490 -1550 18500 -1530
rect 18520 -1550 18530 -1530
rect 18410 -1565 18450 -1550
rect 18490 -1565 18530 -1550
rect 19030 -1330 19070 -1315
rect 19030 -1350 19040 -1330
rect 19060 -1350 19070 -1330
rect 19030 -1380 19070 -1350
rect 19030 -1400 19040 -1380
rect 19060 -1400 19070 -1380
rect 19030 -1430 19070 -1400
rect 19030 -1450 19040 -1430
rect 19060 -1450 19070 -1430
rect 19030 -1480 19070 -1450
rect 19030 -1500 19040 -1480
rect 19060 -1500 19070 -1480
rect 19030 -1530 19070 -1500
rect 19030 -1550 19040 -1530
rect 19060 -1550 19070 -1530
rect 19030 -1565 19070 -1550
rect 16740 -1785 16780 -1770
rect 16740 -1805 16750 -1785
rect 16770 -1805 16780 -1785
rect 16740 -1835 16780 -1805
rect 16740 -1855 16750 -1835
rect 16770 -1855 16780 -1835
rect 16740 -1870 16780 -1855
rect 17780 -1785 17820 -1770
rect 17780 -1805 17790 -1785
rect 17810 -1805 17820 -1785
rect 17780 -1835 17820 -1805
rect 17780 -1855 17790 -1835
rect 17810 -1855 17820 -1835
rect 17780 -1870 17820 -1855
rect 18820 -1785 18860 -1770
rect 18820 -1805 18830 -1785
rect 18850 -1805 18860 -1785
rect 18820 -1835 18860 -1805
rect 18820 -1855 18830 -1835
rect 18850 -1855 18860 -1835
rect 18820 -1870 18860 -1855
<< pdiff >>
rect 16975 625 17015 640
rect 16975 605 16985 625
rect 17005 605 17015 625
rect 16975 575 17015 605
rect 16975 555 16985 575
rect 17005 555 17015 575
rect 16975 540 17015 555
rect 17030 625 17070 640
rect 17030 605 17040 625
rect 17060 605 17070 625
rect 17030 575 17070 605
rect 17030 555 17040 575
rect 17060 555 17070 575
rect 17030 540 17070 555
rect 17085 625 17125 640
rect 17085 605 17095 625
rect 17115 605 17125 625
rect 17085 575 17125 605
rect 17085 555 17095 575
rect 17115 555 17125 575
rect 17085 540 17125 555
rect 17140 625 17180 640
rect 17140 605 17150 625
rect 17170 605 17180 625
rect 17140 575 17180 605
rect 17140 555 17150 575
rect 17170 555 17180 575
rect 17140 540 17180 555
rect 17195 625 17235 640
rect 17195 605 17205 625
rect 17225 605 17235 625
rect 17195 575 17235 605
rect 17195 555 17205 575
rect 17225 555 17235 575
rect 17195 540 17235 555
rect 17250 625 17290 640
rect 17250 605 17260 625
rect 17280 605 17290 625
rect 17250 575 17290 605
rect 17250 555 17260 575
rect 17280 555 17290 575
rect 17250 540 17290 555
rect 17305 625 17345 640
rect 17305 605 17315 625
rect 17335 605 17345 625
rect 17305 575 17345 605
rect 17305 555 17315 575
rect 17335 555 17345 575
rect 17305 540 17345 555
rect 17360 625 17400 640
rect 17360 605 17370 625
rect 17390 605 17400 625
rect 17360 575 17400 605
rect 17360 555 17370 575
rect 17390 555 17400 575
rect 17360 540 17400 555
rect 17415 625 17455 640
rect 17415 605 17425 625
rect 17445 605 17455 625
rect 17415 575 17455 605
rect 17415 555 17425 575
rect 17445 555 17455 575
rect 17415 540 17455 555
rect 17470 625 17510 640
rect 17470 605 17480 625
rect 17500 605 17510 625
rect 17470 575 17510 605
rect 17470 555 17480 575
rect 17500 555 17510 575
rect 17470 540 17510 555
rect 17525 625 17565 640
rect 17525 605 17535 625
rect 17555 605 17565 625
rect 17525 575 17565 605
rect 17525 555 17535 575
rect 17555 555 17565 575
rect 17525 540 17565 555
rect 17580 625 17620 640
rect 17580 605 17590 625
rect 17610 605 17620 625
rect 17580 575 17620 605
rect 17580 555 17590 575
rect 17610 555 17620 575
rect 17580 540 17620 555
rect 17635 625 17675 640
rect 17635 605 17645 625
rect 17665 605 17675 625
rect 17635 575 17675 605
rect 17635 555 17645 575
rect 17665 555 17675 575
rect 17635 540 17675 555
rect 17925 625 17965 640
rect 17925 605 17935 625
rect 17955 605 17965 625
rect 17925 575 17965 605
rect 17925 555 17935 575
rect 17955 555 17965 575
rect 17925 540 17965 555
rect 17980 625 18020 640
rect 17980 605 17990 625
rect 18010 605 18020 625
rect 17980 575 18020 605
rect 17980 555 17990 575
rect 18010 555 18020 575
rect 17980 540 18020 555
rect 18035 625 18075 640
rect 18035 605 18045 625
rect 18065 605 18075 625
rect 18035 575 18075 605
rect 18035 555 18045 575
rect 18065 555 18075 575
rect 18035 540 18075 555
rect 18090 625 18130 640
rect 18090 605 18100 625
rect 18120 605 18130 625
rect 18090 575 18130 605
rect 18090 555 18100 575
rect 18120 555 18130 575
rect 18090 540 18130 555
rect 18145 625 18185 640
rect 18145 605 18155 625
rect 18175 605 18185 625
rect 18145 575 18185 605
rect 18145 555 18155 575
rect 18175 555 18185 575
rect 18145 540 18185 555
rect 18200 625 18240 640
rect 18200 605 18210 625
rect 18230 605 18240 625
rect 18200 575 18240 605
rect 18200 555 18210 575
rect 18230 555 18240 575
rect 18200 540 18240 555
rect 18255 625 18295 640
rect 18255 605 18265 625
rect 18285 605 18295 625
rect 18255 575 18295 605
rect 18255 555 18265 575
rect 18285 555 18295 575
rect 18255 540 18295 555
rect 18310 625 18350 640
rect 18310 605 18320 625
rect 18340 605 18350 625
rect 18310 575 18350 605
rect 18310 555 18320 575
rect 18340 555 18350 575
rect 18310 540 18350 555
rect 18365 625 18405 640
rect 18365 605 18375 625
rect 18395 605 18405 625
rect 18365 575 18405 605
rect 18365 555 18375 575
rect 18395 555 18405 575
rect 18365 540 18405 555
rect 18420 625 18460 640
rect 18420 605 18430 625
rect 18450 605 18460 625
rect 18420 575 18460 605
rect 18420 555 18430 575
rect 18450 555 18460 575
rect 18420 540 18460 555
rect 18475 625 18515 640
rect 18475 605 18485 625
rect 18505 605 18515 625
rect 18475 575 18515 605
rect 18475 555 18485 575
rect 18505 555 18515 575
rect 18475 540 18515 555
rect 18530 625 18570 640
rect 18530 605 18540 625
rect 18560 605 18570 625
rect 18530 575 18570 605
rect 18530 555 18540 575
rect 18560 555 18570 575
rect 18530 540 18570 555
rect 18585 625 18625 640
rect 18585 605 18595 625
rect 18615 605 18625 625
rect 18585 575 18625 605
rect 18585 555 18595 575
rect 18615 555 18625 575
rect 18585 540 18625 555
rect 16970 325 17010 340
rect 16970 305 16980 325
rect 17000 305 17010 325
rect 16970 275 17010 305
rect 16970 255 16980 275
rect 17000 255 17010 275
rect 16435 225 16475 240
rect 16435 205 16445 225
rect 16465 205 16475 225
rect 16435 175 16475 205
rect 16435 155 16445 175
rect 16465 155 16475 175
rect 16435 140 16475 155
rect 16490 225 16530 240
rect 16490 205 16500 225
rect 16520 205 16530 225
rect 16490 175 16530 205
rect 16490 155 16500 175
rect 16520 155 16530 175
rect 16490 140 16530 155
rect 16545 225 16585 240
rect 16545 205 16555 225
rect 16575 205 16585 225
rect 16545 175 16585 205
rect 16545 155 16555 175
rect 16575 155 16585 175
rect 16545 140 16585 155
rect 16600 225 16640 240
rect 16600 205 16610 225
rect 16630 205 16640 225
rect 16600 175 16640 205
rect 16600 155 16610 175
rect 16630 155 16640 175
rect 16600 140 16640 155
rect 16655 225 16700 240
rect 16655 205 16665 225
rect 16685 205 16700 225
rect 16655 175 16700 205
rect 16655 155 16665 175
rect 16685 155 16700 175
rect 16655 140 16700 155
rect 16970 225 17010 255
rect 16970 205 16980 225
rect 17000 205 17010 225
rect 16970 175 17010 205
rect 16970 155 16980 175
rect 17000 155 17010 175
rect 16970 125 17010 155
rect 16970 105 16980 125
rect 17000 105 17010 125
rect 16970 75 17010 105
rect 16970 55 16980 75
rect 17000 55 17010 75
rect 16970 40 17010 55
rect 17060 325 17100 340
rect 17060 305 17070 325
rect 17090 305 17100 325
rect 17060 275 17100 305
rect 17060 255 17070 275
rect 17090 255 17100 275
rect 17060 225 17100 255
rect 17060 205 17070 225
rect 17090 205 17100 225
rect 17060 175 17100 205
rect 17060 155 17070 175
rect 17090 155 17100 175
rect 17060 125 17100 155
rect 17060 105 17070 125
rect 17090 105 17100 125
rect 17060 75 17100 105
rect 17060 55 17070 75
rect 17090 55 17100 75
rect 17060 40 17100 55
rect 17150 325 17190 340
rect 17150 305 17160 325
rect 17180 305 17190 325
rect 17150 275 17190 305
rect 17150 255 17160 275
rect 17180 255 17190 275
rect 17150 225 17190 255
rect 17150 205 17160 225
rect 17180 205 17190 225
rect 17150 175 17190 205
rect 17150 155 17160 175
rect 17180 155 17190 175
rect 17150 125 17190 155
rect 17150 105 17160 125
rect 17180 105 17190 125
rect 17150 75 17190 105
rect 17150 55 17160 75
rect 17180 55 17190 75
rect 17150 40 17190 55
rect 17240 325 17280 340
rect 17240 305 17250 325
rect 17270 305 17280 325
rect 17240 275 17280 305
rect 17240 255 17250 275
rect 17270 255 17280 275
rect 17240 225 17280 255
rect 17240 205 17250 225
rect 17270 205 17280 225
rect 17240 175 17280 205
rect 17240 155 17250 175
rect 17270 155 17280 175
rect 17240 125 17280 155
rect 17240 105 17250 125
rect 17270 105 17280 125
rect 17240 75 17280 105
rect 17240 55 17250 75
rect 17270 55 17280 75
rect 17240 40 17280 55
rect 17330 325 17370 340
rect 17330 305 17340 325
rect 17360 305 17370 325
rect 17330 275 17370 305
rect 17330 255 17340 275
rect 17360 255 17370 275
rect 17330 225 17370 255
rect 17330 205 17340 225
rect 17360 205 17370 225
rect 17330 175 17370 205
rect 17330 155 17340 175
rect 17360 155 17370 175
rect 17330 125 17370 155
rect 17330 105 17340 125
rect 17360 105 17370 125
rect 17330 75 17370 105
rect 17330 55 17340 75
rect 17360 55 17370 75
rect 17330 40 17370 55
rect 17420 325 17460 340
rect 17420 305 17430 325
rect 17450 305 17460 325
rect 17420 275 17460 305
rect 17420 255 17430 275
rect 17450 255 17460 275
rect 17420 225 17460 255
rect 17420 205 17430 225
rect 17450 205 17460 225
rect 17420 175 17460 205
rect 17420 155 17430 175
rect 17450 155 17460 175
rect 17420 125 17460 155
rect 17420 105 17430 125
rect 17450 105 17460 125
rect 17420 75 17460 105
rect 17420 55 17430 75
rect 17450 55 17460 75
rect 17420 40 17460 55
rect 17510 325 17550 340
rect 17510 305 17520 325
rect 17540 305 17550 325
rect 17510 275 17550 305
rect 17510 255 17520 275
rect 17540 255 17550 275
rect 17510 225 17550 255
rect 17510 205 17520 225
rect 17540 205 17550 225
rect 17510 175 17550 205
rect 17510 155 17520 175
rect 17540 155 17550 175
rect 17510 125 17550 155
rect 17510 105 17520 125
rect 17540 105 17550 125
rect 17510 75 17550 105
rect 17510 55 17520 75
rect 17540 55 17550 75
rect 17510 40 17550 55
rect 17600 325 17640 340
rect 17600 305 17610 325
rect 17630 305 17640 325
rect 17600 275 17640 305
rect 17600 255 17610 275
rect 17630 255 17640 275
rect 17600 225 17640 255
rect 17600 205 17610 225
rect 17630 205 17640 225
rect 17600 175 17640 205
rect 17600 155 17610 175
rect 17630 155 17640 175
rect 17600 125 17640 155
rect 17600 105 17610 125
rect 17630 105 17640 125
rect 17600 75 17640 105
rect 17600 55 17610 75
rect 17630 55 17640 75
rect 17600 40 17640 55
rect 17690 325 17730 340
rect 17690 305 17700 325
rect 17720 305 17730 325
rect 17690 275 17730 305
rect 17690 255 17700 275
rect 17720 255 17730 275
rect 17690 225 17730 255
rect 17690 205 17700 225
rect 17720 205 17730 225
rect 17690 175 17730 205
rect 17690 155 17700 175
rect 17720 155 17730 175
rect 17690 125 17730 155
rect 17690 105 17700 125
rect 17720 105 17730 125
rect 17690 75 17730 105
rect 17690 55 17700 75
rect 17720 55 17730 75
rect 17690 40 17730 55
rect 17780 325 17820 340
rect 17780 305 17790 325
rect 17810 305 17820 325
rect 17780 275 17820 305
rect 17780 255 17790 275
rect 17810 255 17820 275
rect 17780 225 17820 255
rect 17780 205 17790 225
rect 17810 205 17820 225
rect 17780 175 17820 205
rect 17780 155 17790 175
rect 17810 155 17820 175
rect 17780 125 17820 155
rect 17780 105 17790 125
rect 17810 105 17820 125
rect 17780 75 17820 105
rect 17780 55 17790 75
rect 17810 55 17820 75
rect 17780 40 17820 55
rect 17870 325 17910 340
rect 17870 305 17880 325
rect 17900 305 17910 325
rect 17870 275 17910 305
rect 17870 255 17880 275
rect 17900 255 17910 275
rect 17870 225 17910 255
rect 17870 205 17880 225
rect 17900 205 17910 225
rect 17870 175 17910 205
rect 17870 155 17880 175
rect 17900 155 17910 175
rect 17870 125 17910 155
rect 17870 105 17880 125
rect 17900 105 17910 125
rect 17870 75 17910 105
rect 17870 55 17880 75
rect 17900 55 17910 75
rect 17870 40 17910 55
rect 17960 325 18000 340
rect 17960 305 17970 325
rect 17990 305 18000 325
rect 17960 275 18000 305
rect 17960 255 17970 275
rect 17990 255 18000 275
rect 17960 225 18000 255
rect 17960 205 17970 225
rect 17990 205 18000 225
rect 17960 175 18000 205
rect 17960 155 17970 175
rect 17990 155 18000 175
rect 17960 125 18000 155
rect 17960 105 17970 125
rect 17990 105 18000 125
rect 17960 75 18000 105
rect 17960 55 17970 75
rect 17990 55 18000 75
rect 17960 40 18000 55
rect 18050 325 18090 340
rect 18050 305 18060 325
rect 18080 305 18090 325
rect 18050 275 18090 305
rect 18050 255 18060 275
rect 18080 255 18090 275
rect 18050 225 18090 255
rect 18050 205 18060 225
rect 18080 205 18090 225
rect 18050 175 18090 205
rect 18050 155 18060 175
rect 18080 155 18090 175
rect 18050 125 18090 155
rect 18050 105 18060 125
rect 18080 105 18090 125
rect 18050 75 18090 105
rect 18050 55 18060 75
rect 18080 55 18090 75
rect 18050 40 18090 55
rect 18140 325 18180 340
rect 18140 305 18150 325
rect 18170 305 18180 325
rect 18140 275 18180 305
rect 18140 255 18150 275
rect 18170 255 18180 275
rect 18140 225 18180 255
rect 18140 205 18150 225
rect 18170 205 18180 225
rect 18140 175 18180 205
rect 18140 155 18150 175
rect 18170 155 18180 175
rect 18140 125 18180 155
rect 18140 105 18150 125
rect 18170 105 18180 125
rect 18140 75 18180 105
rect 18140 55 18150 75
rect 18170 55 18180 75
rect 18140 40 18180 55
rect 18230 325 18270 340
rect 18230 305 18240 325
rect 18260 305 18270 325
rect 18230 275 18270 305
rect 18230 255 18240 275
rect 18260 255 18270 275
rect 18230 225 18270 255
rect 18230 205 18240 225
rect 18260 205 18270 225
rect 18230 175 18270 205
rect 18230 155 18240 175
rect 18260 155 18270 175
rect 18230 125 18270 155
rect 18230 105 18240 125
rect 18260 105 18270 125
rect 18230 75 18270 105
rect 18230 55 18240 75
rect 18260 55 18270 75
rect 18230 40 18270 55
rect 18320 325 18360 340
rect 18320 305 18330 325
rect 18350 305 18360 325
rect 18320 275 18360 305
rect 18320 255 18330 275
rect 18350 255 18360 275
rect 18320 225 18360 255
rect 18320 205 18330 225
rect 18350 205 18360 225
rect 18320 175 18360 205
rect 18320 155 18330 175
rect 18350 155 18360 175
rect 18320 125 18360 155
rect 18320 105 18330 125
rect 18350 105 18360 125
rect 18320 75 18360 105
rect 18320 55 18330 75
rect 18350 55 18360 75
rect 18320 40 18360 55
rect 18410 325 18450 340
rect 18410 305 18420 325
rect 18440 305 18450 325
rect 18410 275 18450 305
rect 18410 255 18420 275
rect 18440 255 18450 275
rect 18410 225 18450 255
rect 18410 205 18420 225
rect 18440 205 18450 225
rect 18410 175 18450 205
rect 18410 155 18420 175
rect 18440 155 18450 175
rect 18410 125 18450 155
rect 18410 105 18420 125
rect 18440 105 18450 125
rect 18410 75 18450 105
rect 18410 55 18420 75
rect 18440 55 18450 75
rect 18410 40 18450 55
rect 18500 325 18540 340
rect 18500 305 18510 325
rect 18530 305 18540 325
rect 18500 275 18540 305
rect 18500 255 18510 275
rect 18530 255 18540 275
rect 18500 225 18540 255
rect 18500 205 18510 225
rect 18530 205 18540 225
rect 18500 175 18540 205
rect 18500 155 18510 175
rect 18530 155 18540 175
rect 18500 125 18540 155
rect 18500 105 18510 125
rect 18530 105 18540 125
rect 18500 75 18540 105
rect 18500 55 18510 75
rect 18530 55 18540 75
rect 18500 40 18540 55
rect 18590 325 18630 340
rect 18590 305 18600 325
rect 18620 305 18630 325
rect 18590 275 18630 305
rect 18590 255 18600 275
rect 18620 255 18630 275
rect 18590 225 18630 255
rect 18590 205 18600 225
rect 18620 205 18630 225
rect 18590 175 18630 205
rect 18590 155 18600 175
rect 18620 155 18630 175
rect 18590 125 18630 155
rect 18590 105 18600 125
rect 18620 105 18630 125
rect 18590 75 18630 105
rect 18590 55 18600 75
rect 18620 55 18630 75
rect 18590 40 18630 55
rect 16420 -455 16460 -440
rect 16420 -475 16430 -455
rect 16450 -475 16460 -455
rect 16420 -505 16460 -475
rect 16420 -525 16430 -505
rect 16450 -525 16460 -505
rect 16420 -540 16460 -525
rect 16480 -455 16520 -440
rect 16480 -475 16490 -455
rect 16510 -475 16520 -455
rect 16480 -505 16520 -475
rect 16480 -525 16490 -505
rect 16510 -525 16520 -505
rect 16480 -540 16520 -525
rect 16540 -455 16580 -440
rect 16540 -475 16550 -455
rect 16570 -475 16580 -455
rect 16540 -505 16580 -475
rect 16540 -525 16550 -505
rect 16570 -525 16580 -505
rect 16540 -540 16580 -525
rect 16600 -455 16640 -440
rect 16600 -475 16610 -455
rect 16630 -475 16640 -455
rect 16600 -505 16640 -475
rect 16600 -525 16610 -505
rect 16630 -525 16640 -505
rect 16600 -540 16640 -525
rect 16660 -455 16700 -440
rect 16660 -475 16670 -455
rect 16690 -475 16700 -455
rect 16660 -505 16700 -475
rect 16660 -525 16670 -505
rect 16690 -525 16700 -505
rect 16660 -540 16700 -525
rect 16720 -455 16760 -440
rect 16720 -475 16730 -455
rect 16750 -475 16760 -455
rect 16720 -505 16760 -475
rect 16720 -525 16730 -505
rect 16750 -525 16760 -505
rect 16720 -540 16760 -525
rect 16780 -455 16820 -440
rect 16780 -475 16790 -455
rect 16810 -475 16820 -455
rect 16780 -505 16820 -475
rect 16780 -525 16790 -505
rect 16810 -525 16820 -505
rect 16780 -540 16820 -525
rect 16840 -455 16880 -440
rect 16840 -475 16850 -455
rect 16870 -475 16880 -455
rect 16840 -505 16880 -475
rect 16840 -525 16850 -505
rect 16870 -525 16880 -505
rect 16840 -540 16880 -525
rect 16900 -455 16940 -440
rect 16900 -475 16910 -455
rect 16930 -475 16940 -455
rect 16900 -505 16940 -475
rect 16900 -525 16910 -505
rect 16930 -525 16940 -505
rect 16900 -540 16940 -525
rect 16960 -455 17000 -440
rect 16960 -475 16970 -455
rect 16990 -475 17000 -455
rect 16960 -505 17000 -475
rect 16960 -525 16970 -505
rect 16990 -525 17000 -505
rect 16960 -540 17000 -525
rect 17020 -455 17060 -440
rect 17020 -475 17030 -455
rect 17050 -475 17060 -455
rect 17020 -505 17060 -475
rect 17020 -525 17030 -505
rect 17050 -525 17060 -505
rect 17020 -540 17060 -525
rect 17080 -455 17120 -440
rect 17080 -475 17090 -455
rect 17110 -475 17120 -455
rect 17080 -505 17120 -475
rect 17080 -525 17090 -505
rect 17110 -525 17120 -505
rect 17080 -540 17120 -525
rect 17140 -455 17180 -440
rect 17140 -475 17150 -455
rect 17170 -475 17180 -455
rect 17140 -505 17180 -475
rect 17140 -525 17150 -505
rect 17170 -525 17180 -505
rect 17140 -540 17180 -525
rect 17200 -455 17240 -440
rect 17200 -475 17210 -455
rect 17230 -475 17240 -455
rect 17200 -505 17240 -475
rect 17200 -525 17210 -505
rect 17230 -525 17240 -505
rect 17200 -540 17240 -525
rect 17260 -455 17300 -440
rect 17260 -475 17270 -455
rect 17290 -475 17300 -455
rect 17260 -505 17300 -475
rect 17260 -525 17270 -505
rect 17290 -525 17300 -505
rect 17260 -540 17300 -525
rect 17320 -455 17360 -440
rect 17320 -475 17330 -455
rect 17350 -475 17360 -455
rect 17320 -505 17360 -475
rect 17320 -525 17330 -505
rect 17350 -525 17360 -505
rect 17320 -540 17360 -525
rect 17380 -455 17420 -440
rect 17380 -475 17390 -455
rect 17410 -475 17420 -455
rect 17380 -505 17420 -475
rect 17380 -525 17390 -505
rect 17410 -525 17420 -505
rect 17380 -540 17420 -525
rect 17440 -455 17480 -440
rect 17440 -475 17450 -455
rect 17470 -475 17480 -455
rect 17440 -505 17480 -475
rect 17440 -525 17450 -505
rect 17470 -525 17480 -505
rect 17440 -540 17480 -525
rect 17500 -455 17540 -440
rect 17500 -475 17510 -455
rect 17530 -475 17540 -455
rect 17500 -505 17540 -475
rect 17500 -525 17510 -505
rect 17530 -525 17540 -505
rect 17500 -540 17540 -525
rect 17560 -455 17600 -440
rect 17560 -475 17570 -455
rect 17590 -475 17600 -455
rect 17560 -505 17600 -475
rect 17560 -525 17570 -505
rect 17590 -525 17600 -505
rect 17560 -540 17600 -525
rect 17620 -455 17660 -440
rect 17620 -475 17630 -455
rect 17650 -475 17660 -455
rect 17620 -505 17660 -475
rect 17620 -525 17630 -505
rect 17650 -525 17660 -505
rect 17620 -540 17660 -525
rect 17940 -455 17980 -440
rect 17940 -475 17950 -455
rect 17970 -475 17980 -455
rect 17940 -505 17980 -475
rect 17940 -525 17950 -505
rect 17970 -525 17980 -505
rect 17940 -540 17980 -525
rect 18000 -455 18040 -440
rect 18000 -475 18010 -455
rect 18030 -475 18040 -455
rect 18000 -505 18040 -475
rect 18000 -525 18010 -505
rect 18030 -525 18040 -505
rect 18000 -540 18040 -525
rect 18060 -455 18100 -440
rect 18060 -475 18070 -455
rect 18090 -475 18100 -455
rect 18060 -505 18100 -475
rect 18060 -525 18070 -505
rect 18090 -525 18100 -505
rect 18060 -540 18100 -525
rect 18120 -455 18160 -440
rect 18120 -475 18130 -455
rect 18150 -475 18160 -455
rect 18120 -505 18160 -475
rect 18120 -525 18130 -505
rect 18150 -525 18160 -505
rect 18120 -540 18160 -525
rect 18180 -455 18220 -440
rect 18180 -475 18190 -455
rect 18210 -475 18220 -455
rect 18180 -505 18220 -475
rect 18180 -525 18190 -505
rect 18210 -525 18220 -505
rect 18180 -540 18220 -525
rect 18240 -455 18280 -440
rect 18240 -475 18250 -455
rect 18270 -475 18280 -455
rect 18240 -505 18280 -475
rect 18240 -525 18250 -505
rect 18270 -525 18280 -505
rect 18240 -540 18280 -525
rect 18300 -455 18340 -440
rect 18300 -475 18310 -455
rect 18330 -475 18340 -455
rect 18300 -505 18340 -475
rect 18300 -525 18310 -505
rect 18330 -525 18340 -505
rect 18300 -540 18340 -525
rect 18360 -455 18400 -440
rect 18360 -475 18370 -455
rect 18390 -475 18400 -455
rect 18360 -505 18400 -475
rect 18360 -525 18370 -505
rect 18390 -525 18400 -505
rect 18360 -540 18400 -525
rect 18420 -455 18460 -440
rect 18420 -475 18430 -455
rect 18450 -475 18460 -455
rect 18420 -505 18460 -475
rect 18420 -525 18430 -505
rect 18450 -525 18460 -505
rect 18420 -540 18460 -525
rect 18480 -455 18520 -440
rect 18480 -475 18490 -455
rect 18510 -475 18520 -455
rect 18480 -505 18520 -475
rect 18480 -525 18490 -505
rect 18510 -525 18520 -505
rect 18480 -540 18520 -525
rect 18540 -455 18580 -440
rect 18540 -475 18550 -455
rect 18570 -475 18580 -455
rect 18540 -505 18580 -475
rect 18540 -525 18550 -505
rect 18570 -525 18580 -505
rect 18540 -540 18580 -525
rect 18600 -455 18640 -440
rect 18600 -475 18610 -455
rect 18630 -475 18640 -455
rect 18600 -505 18640 -475
rect 18600 -525 18610 -505
rect 18630 -525 18640 -505
rect 18600 -540 18640 -525
rect 18660 -455 18700 -440
rect 18660 -475 18670 -455
rect 18690 -475 18700 -455
rect 18660 -505 18700 -475
rect 18660 -525 18670 -505
rect 18690 -525 18700 -505
rect 18660 -540 18700 -525
rect 18720 -455 18760 -440
rect 18720 -475 18730 -455
rect 18750 -475 18760 -455
rect 18720 -505 18760 -475
rect 18720 -525 18730 -505
rect 18750 -525 18760 -505
rect 18720 -540 18760 -525
rect 18780 -455 18820 -440
rect 18780 -475 18790 -455
rect 18810 -475 18820 -455
rect 18780 -505 18820 -475
rect 18780 -525 18790 -505
rect 18810 -525 18820 -505
rect 18780 -540 18820 -525
rect 18840 -455 18880 -440
rect 18840 -475 18850 -455
rect 18870 -475 18880 -455
rect 18840 -505 18880 -475
rect 18840 -525 18850 -505
rect 18870 -525 18880 -505
rect 18840 -540 18880 -525
rect 18900 -455 18940 -440
rect 18900 -475 18910 -455
rect 18930 -475 18940 -455
rect 18900 -505 18940 -475
rect 18900 -525 18910 -505
rect 18930 -525 18940 -505
rect 18900 -540 18940 -525
rect 18960 -455 19000 -440
rect 18960 -475 18970 -455
rect 18990 -475 19000 -455
rect 18960 -505 19000 -475
rect 18960 -525 18970 -505
rect 18990 -525 19000 -505
rect 18960 -540 19000 -525
rect 19020 -455 19060 -440
rect 19020 -475 19030 -455
rect 19050 -475 19060 -455
rect 19020 -505 19060 -475
rect 19020 -525 19030 -505
rect 19050 -525 19060 -505
rect 19020 -540 19060 -525
rect 19080 -455 19120 -440
rect 19080 -475 19090 -455
rect 19110 -475 19120 -455
rect 19080 -505 19120 -475
rect 19080 -525 19090 -505
rect 19110 -525 19120 -505
rect 19080 -540 19120 -525
rect 19140 -455 19180 -440
rect 19140 -475 19150 -455
rect 19170 -475 19180 -455
rect 19140 -505 19180 -475
rect 19140 -525 19150 -505
rect 19170 -525 19180 -505
rect 19140 -540 19180 -525
<< ndiffc >>
rect 16970 -840 16990 -820
rect 16970 -890 16990 -870
rect 16970 -940 16990 -920
rect 16970 -990 16990 -970
rect 16970 -1040 16990 -1020
rect 17030 -840 17050 -820
rect 17030 -890 17050 -870
rect 17030 -940 17050 -920
rect 17030 -990 17050 -970
rect 17030 -1040 17050 -1020
rect 17090 -840 17110 -820
rect 17090 -890 17110 -870
rect 17090 -940 17110 -920
rect 18490 -840 18510 -820
rect 18490 -890 18510 -870
rect 17090 -990 17110 -970
rect 17090 -1040 17110 -1020
rect 18490 -940 18510 -920
rect 18490 -990 18510 -970
rect 18490 -1040 18510 -1020
rect 18550 -840 18570 -820
rect 18550 -890 18570 -870
rect 18550 -940 18570 -920
rect 18550 -990 18570 -970
rect 18550 -1040 18570 -1020
rect 18610 -840 18630 -820
rect 18610 -890 18630 -870
rect 18610 -940 18630 -920
rect 18610 -990 18630 -970
rect 18610 -1040 18630 -1020
rect 16540 -1350 16560 -1330
rect 16540 -1400 16560 -1380
rect 16540 -1450 16560 -1430
rect 16540 -1500 16560 -1480
rect 16540 -1550 16560 -1530
rect 17080 -1350 17100 -1330
rect 17160 -1350 17180 -1330
rect 17080 -1400 17100 -1380
rect 17160 -1400 17180 -1380
rect 17080 -1450 17100 -1430
rect 17160 -1450 17180 -1430
rect 17080 -1500 17100 -1480
rect 17160 -1500 17180 -1480
rect 17080 -1550 17100 -1530
rect 17160 -1550 17180 -1530
rect 17700 -1350 17720 -1330
rect 17700 -1400 17720 -1380
rect 17700 -1450 17720 -1430
rect 17700 -1500 17720 -1480
rect 17700 -1550 17720 -1530
rect 17880 -1350 17900 -1330
rect 17880 -1400 17900 -1380
rect 17880 -1450 17900 -1430
rect 17880 -1500 17900 -1480
rect 17880 -1550 17900 -1530
rect 18420 -1350 18440 -1330
rect 18500 -1350 18520 -1330
rect 18420 -1400 18440 -1380
rect 18500 -1400 18520 -1380
rect 18420 -1450 18440 -1430
rect 18500 -1450 18520 -1430
rect 18420 -1500 18440 -1480
rect 18500 -1500 18520 -1480
rect 18420 -1550 18440 -1530
rect 18500 -1550 18520 -1530
rect 19040 -1350 19060 -1330
rect 19040 -1400 19060 -1380
rect 19040 -1450 19060 -1430
rect 19040 -1500 19060 -1480
rect 19040 -1550 19060 -1530
rect 16750 -1805 16770 -1785
rect 16750 -1855 16770 -1835
rect 17790 -1805 17810 -1785
rect 17790 -1855 17810 -1835
rect 18830 -1805 18850 -1785
rect 18830 -1855 18850 -1835
<< pdiffc >>
rect 16985 605 17005 625
rect 16985 555 17005 575
rect 17040 605 17060 625
rect 17040 555 17060 575
rect 17095 605 17115 625
rect 17095 555 17115 575
rect 17150 605 17170 625
rect 17150 555 17170 575
rect 17205 605 17225 625
rect 17205 555 17225 575
rect 17260 605 17280 625
rect 17260 555 17280 575
rect 17315 605 17335 625
rect 17315 555 17335 575
rect 17370 605 17390 625
rect 17370 555 17390 575
rect 17425 605 17445 625
rect 17425 555 17445 575
rect 17480 605 17500 625
rect 17480 555 17500 575
rect 17535 605 17555 625
rect 17535 555 17555 575
rect 17590 605 17610 625
rect 17590 555 17610 575
rect 17645 605 17665 625
rect 17645 555 17665 575
rect 17935 605 17955 625
rect 17935 555 17955 575
rect 17990 605 18010 625
rect 17990 555 18010 575
rect 18045 605 18065 625
rect 18045 555 18065 575
rect 18100 605 18120 625
rect 18100 555 18120 575
rect 18155 605 18175 625
rect 18155 555 18175 575
rect 18210 605 18230 625
rect 18210 555 18230 575
rect 18265 605 18285 625
rect 18265 555 18285 575
rect 18320 605 18340 625
rect 18320 555 18340 575
rect 18375 605 18395 625
rect 18375 555 18395 575
rect 18430 605 18450 625
rect 18430 555 18450 575
rect 18485 605 18505 625
rect 18485 555 18505 575
rect 18540 605 18560 625
rect 18540 555 18560 575
rect 18595 605 18615 625
rect 18595 555 18615 575
rect 16980 305 17000 325
rect 16980 255 17000 275
rect 16445 205 16465 225
rect 16445 155 16465 175
rect 16500 205 16520 225
rect 16500 155 16520 175
rect 16555 205 16575 225
rect 16555 155 16575 175
rect 16610 205 16630 225
rect 16610 155 16630 175
rect 16665 205 16685 225
rect 16665 155 16685 175
rect 16980 205 17000 225
rect 16980 155 17000 175
rect 16980 105 17000 125
rect 16980 55 17000 75
rect 17070 305 17090 325
rect 17070 255 17090 275
rect 17070 205 17090 225
rect 17070 155 17090 175
rect 17070 105 17090 125
rect 17070 55 17090 75
rect 17160 305 17180 325
rect 17160 255 17180 275
rect 17160 205 17180 225
rect 17160 155 17180 175
rect 17160 105 17180 125
rect 17160 55 17180 75
rect 17250 305 17270 325
rect 17250 255 17270 275
rect 17250 205 17270 225
rect 17250 155 17270 175
rect 17250 105 17270 125
rect 17250 55 17270 75
rect 17340 305 17360 325
rect 17340 255 17360 275
rect 17340 205 17360 225
rect 17340 155 17360 175
rect 17340 105 17360 125
rect 17340 55 17360 75
rect 17430 305 17450 325
rect 17430 255 17450 275
rect 17430 205 17450 225
rect 17430 155 17450 175
rect 17430 105 17450 125
rect 17430 55 17450 75
rect 17520 305 17540 325
rect 17520 255 17540 275
rect 17520 205 17540 225
rect 17520 155 17540 175
rect 17520 105 17540 125
rect 17520 55 17540 75
rect 17610 305 17630 325
rect 17610 255 17630 275
rect 17610 205 17630 225
rect 17610 155 17630 175
rect 17610 105 17630 125
rect 17610 55 17630 75
rect 17700 305 17720 325
rect 17700 255 17720 275
rect 17700 205 17720 225
rect 17700 155 17720 175
rect 17700 105 17720 125
rect 17700 55 17720 75
rect 17790 305 17810 325
rect 17790 255 17810 275
rect 17790 205 17810 225
rect 17790 155 17810 175
rect 17790 105 17810 125
rect 17790 55 17810 75
rect 17880 305 17900 325
rect 17880 255 17900 275
rect 17880 205 17900 225
rect 17880 155 17900 175
rect 17880 105 17900 125
rect 17880 55 17900 75
rect 17970 305 17990 325
rect 17970 255 17990 275
rect 17970 205 17990 225
rect 17970 155 17990 175
rect 17970 105 17990 125
rect 17970 55 17990 75
rect 18060 305 18080 325
rect 18060 255 18080 275
rect 18060 205 18080 225
rect 18060 155 18080 175
rect 18060 105 18080 125
rect 18060 55 18080 75
rect 18150 305 18170 325
rect 18150 255 18170 275
rect 18150 205 18170 225
rect 18150 155 18170 175
rect 18150 105 18170 125
rect 18150 55 18170 75
rect 18240 305 18260 325
rect 18240 255 18260 275
rect 18240 205 18260 225
rect 18240 155 18260 175
rect 18240 105 18260 125
rect 18240 55 18260 75
rect 18330 305 18350 325
rect 18330 255 18350 275
rect 18330 205 18350 225
rect 18330 155 18350 175
rect 18330 105 18350 125
rect 18330 55 18350 75
rect 18420 305 18440 325
rect 18420 255 18440 275
rect 18420 205 18440 225
rect 18420 155 18440 175
rect 18420 105 18440 125
rect 18420 55 18440 75
rect 18510 305 18530 325
rect 18510 255 18530 275
rect 18510 205 18530 225
rect 18510 155 18530 175
rect 18510 105 18530 125
rect 18510 55 18530 75
rect 18600 305 18620 325
rect 18600 255 18620 275
rect 18600 205 18620 225
rect 18600 155 18620 175
rect 18600 105 18620 125
rect 18600 55 18620 75
rect 16430 -475 16450 -455
rect 16430 -525 16450 -505
rect 16490 -475 16510 -455
rect 16490 -525 16510 -505
rect 16550 -475 16570 -455
rect 16550 -525 16570 -505
rect 16610 -475 16630 -455
rect 16610 -525 16630 -505
rect 16670 -475 16690 -455
rect 16670 -525 16690 -505
rect 16730 -475 16750 -455
rect 16730 -525 16750 -505
rect 16790 -475 16810 -455
rect 16790 -525 16810 -505
rect 16850 -475 16870 -455
rect 16850 -525 16870 -505
rect 16910 -475 16930 -455
rect 16910 -525 16930 -505
rect 16970 -475 16990 -455
rect 16970 -525 16990 -505
rect 17030 -475 17050 -455
rect 17030 -525 17050 -505
rect 17090 -475 17110 -455
rect 17090 -525 17110 -505
rect 17150 -475 17170 -455
rect 17150 -525 17170 -505
rect 17210 -475 17230 -455
rect 17210 -525 17230 -505
rect 17270 -475 17290 -455
rect 17270 -525 17290 -505
rect 17330 -475 17350 -455
rect 17330 -525 17350 -505
rect 17390 -475 17410 -455
rect 17390 -525 17410 -505
rect 17450 -475 17470 -455
rect 17450 -525 17470 -505
rect 17510 -475 17530 -455
rect 17510 -525 17530 -505
rect 17570 -475 17590 -455
rect 17570 -525 17590 -505
rect 17630 -475 17650 -455
rect 17630 -525 17650 -505
rect 17950 -475 17970 -455
rect 17950 -525 17970 -505
rect 18010 -475 18030 -455
rect 18010 -525 18030 -505
rect 18070 -475 18090 -455
rect 18070 -525 18090 -505
rect 18130 -475 18150 -455
rect 18130 -525 18150 -505
rect 18190 -475 18210 -455
rect 18190 -525 18210 -505
rect 18250 -475 18270 -455
rect 18250 -525 18270 -505
rect 18310 -475 18330 -455
rect 18310 -525 18330 -505
rect 18370 -475 18390 -455
rect 18370 -525 18390 -505
rect 18430 -475 18450 -455
rect 18430 -525 18450 -505
rect 18490 -475 18510 -455
rect 18490 -525 18510 -505
rect 18550 -475 18570 -455
rect 18550 -525 18570 -505
rect 18610 -475 18630 -455
rect 18610 -525 18630 -505
rect 18670 -475 18690 -455
rect 18670 -525 18690 -505
rect 18730 -475 18750 -455
rect 18730 -525 18750 -505
rect 18790 -475 18810 -455
rect 18790 -525 18810 -505
rect 18850 -475 18870 -455
rect 18850 -525 18870 -505
rect 18910 -475 18930 -455
rect 18910 -525 18930 -505
rect 18970 -475 18990 -455
rect 18970 -525 18990 -505
rect 19030 -475 19050 -455
rect 19030 -525 19050 -505
rect 19090 -475 19110 -455
rect 19090 -525 19110 -505
rect 19150 -475 19170 -455
rect 19150 -525 19170 -505
<< psubdiff >>
rect 17560 -820 17600 -805
rect 17560 -840 17570 -820
rect 17590 -840 17600 -820
rect 17560 -860 17600 -840
rect 17560 -880 17570 -860
rect 17590 -880 17600 -860
rect 17560 -900 17600 -880
rect 17560 -920 17570 -900
rect 17590 -920 17600 -900
rect 17560 -935 17600 -920
rect 18000 -820 18040 -805
rect 18000 -840 18010 -820
rect 18030 -840 18040 -820
rect 18000 -860 18040 -840
rect 18000 -880 18010 -860
rect 18030 -880 18040 -860
rect 18000 -900 18040 -880
rect 18000 -920 18010 -900
rect 18030 -920 18040 -900
rect 18000 -935 18040 -920
rect 17110 -1330 17150 -1315
rect 17110 -1350 17120 -1330
rect 17140 -1350 17150 -1330
rect 17110 -1380 17150 -1350
rect 17110 -1400 17120 -1380
rect 17140 -1400 17150 -1380
rect 17110 -1430 17150 -1400
rect 17110 -1450 17120 -1430
rect 17140 -1450 17150 -1430
rect 17110 -1480 17150 -1450
rect 17110 -1500 17120 -1480
rect 17140 -1500 17150 -1480
rect 17110 -1530 17150 -1500
rect 17110 -1550 17120 -1530
rect 17140 -1550 17150 -1530
rect 17110 -1560 17150 -1550
rect 18450 -1330 18490 -1315
rect 18450 -1350 18460 -1330
rect 18480 -1350 18490 -1330
rect 18450 -1380 18490 -1350
rect 18450 -1400 18460 -1380
rect 18480 -1400 18490 -1380
rect 18450 -1430 18490 -1400
rect 18450 -1450 18460 -1430
rect 18480 -1450 18490 -1430
rect 18450 -1480 18490 -1450
rect 18450 -1500 18460 -1480
rect 18480 -1500 18490 -1480
rect 18450 -1530 18490 -1500
rect 18450 -1550 18460 -1530
rect 18480 -1550 18490 -1530
rect 18450 -1565 18490 -1550
rect 18860 -1785 18900 -1770
rect 18860 -1805 18870 -1785
rect 18890 -1805 18900 -1785
rect 18860 -1835 18900 -1805
rect 18860 -1855 18870 -1835
rect 18890 -1855 18900 -1835
rect 18860 -1870 18900 -1855
rect 17775 -4165 17825 -4150
rect 17775 -4185 17790 -4165
rect 17810 -4185 17825 -4165
rect 17775 -4205 17825 -4185
rect 17775 -4225 17790 -4205
rect 17810 -4225 17825 -4205
rect 17775 -4245 17825 -4225
rect 17775 -4265 17790 -4245
rect 17810 -4265 17825 -4245
rect 17775 -4280 17825 -4265
<< nsubdiff >>
rect 16935 625 16975 640
rect 16935 605 16945 625
rect 16965 605 16975 625
rect 16935 575 16975 605
rect 16935 555 16945 575
rect 16965 555 16975 575
rect 16935 540 16975 555
rect 17675 625 17715 640
rect 17675 605 17685 625
rect 17705 605 17715 625
rect 17675 575 17715 605
rect 17675 555 17685 575
rect 17705 555 17715 575
rect 17675 540 17715 555
rect 17885 625 17925 640
rect 17885 605 17895 625
rect 17915 605 17925 625
rect 17885 575 17925 605
rect 17885 555 17895 575
rect 17915 555 17925 575
rect 17885 540 17925 555
rect 18625 625 18665 640
rect 18625 605 18635 625
rect 18655 605 18665 625
rect 18625 575 18665 605
rect 18625 555 18635 575
rect 18655 555 18665 575
rect 18625 540 18665 555
rect 16930 325 16970 340
rect 16930 305 16940 325
rect 16960 305 16970 325
rect 16930 275 16970 305
rect 16930 255 16940 275
rect 16960 255 16970 275
rect 16395 225 16435 240
rect 16395 205 16405 225
rect 16425 205 16435 225
rect 16395 175 16435 205
rect 16395 155 16405 175
rect 16425 155 16435 175
rect 16395 140 16435 155
rect 16700 225 16740 240
rect 16700 205 16710 225
rect 16730 205 16740 225
rect 16700 175 16740 205
rect 16700 155 16710 175
rect 16730 155 16740 175
rect 16700 140 16740 155
rect 16930 225 16970 255
rect 16930 205 16940 225
rect 16960 205 16970 225
rect 16930 175 16970 205
rect 16930 155 16940 175
rect 16960 155 16970 175
rect 16930 125 16970 155
rect 16930 105 16940 125
rect 16960 105 16970 125
rect 16930 75 16970 105
rect 16930 55 16940 75
rect 16960 55 16970 75
rect 16930 40 16970 55
rect 18630 325 18670 340
rect 18630 305 18640 325
rect 18660 305 18670 325
rect 18630 275 18670 305
rect 18630 255 18640 275
rect 18660 255 18670 275
rect 18630 225 18670 255
rect 18630 205 18640 225
rect 18660 205 18670 225
rect 18630 175 18670 205
rect 18630 155 18640 175
rect 18660 155 18670 175
rect 18630 125 18670 155
rect 18630 105 18640 125
rect 18660 105 18670 125
rect 18630 75 18670 105
rect 18630 55 18640 75
rect 18660 55 18670 75
rect 18630 40 18670 55
rect 16380 -455 16420 -440
rect 16380 -475 16390 -455
rect 16410 -475 16420 -455
rect 16380 -505 16420 -475
rect 16380 -525 16390 -505
rect 16410 -525 16420 -505
rect 16380 -540 16420 -525
rect 17660 -455 17700 -440
rect 17660 -475 17670 -455
rect 17690 -475 17700 -455
rect 17660 -505 17700 -475
rect 17660 -525 17670 -505
rect 17690 -525 17700 -505
rect 17660 -540 17700 -525
rect 17900 -455 17940 -440
rect 17900 -475 17910 -455
rect 17930 -475 17940 -455
rect 17900 -505 17940 -475
rect 17900 -525 17910 -505
rect 17930 -525 17940 -505
rect 17900 -540 17940 -525
rect 19180 -455 19220 -440
rect 19180 -475 19190 -455
rect 19210 -475 19220 -455
rect 19180 -505 19220 -475
rect 19180 -525 19190 -505
rect 19210 -525 19220 -505
rect 19180 -540 19220 -525
<< psubdiffcont >>
rect 17570 -840 17590 -820
rect 17570 -880 17590 -860
rect 17570 -920 17590 -900
rect 18010 -840 18030 -820
rect 18010 -880 18030 -860
rect 18010 -920 18030 -900
rect 17120 -1350 17140 -1330
rect 17120 -1400 17140 -1380
rect 17120 -1450 17140 -1430
rect 17120 -1500 17140 -1480
rect 17120 -1550 17140 -1530
rect 18460 -1350 18480 -1330
rect 18460 -1400 18480 -1380
rect 18460 -1450 18480 -1430
rect 18460 -1500 18480 -1480
rect 18460 -1550 18480 -1530
rect 18870 -1805 18890 -1785
rect 18870 -1855 18890 -1835
rect 17790 -4185 17810 -4165
rect 17790 -4225 17810 -4205
rect 17790 -4265 17810 -4245
<< nsubdiffcont >>
rect 16945 605 16965 625
rect 16945 555 16965 575
rect 17685 605 17705 625
rect 17685 555 17705 575
rect 17895 605 17915 625
rect 17895 555 17915 575
rect 18635 605 18655 625
rect 18635 555 18655 575
rect 16940 305 16960 325
rect 16940 255 16960 275
rect 16405 205 16425 225
rect 16405 155 16425 175
rect 16710 205 16730 225
rect 16710 155 16730 175
rect 16940 205 16960 225
rect 16940 155 16960 175
rect 16940 105 16960 125
rect 16940 55 16960 75
rect 18640 305 18660 325
rect 18640 255 18660 275
rect 18640 205 18660 225
rect 18640 155 18660 175
rect 18640 105 18660 125
rect 18640 55 18660 75
rect 16390 -475 16410 -455
rect 16390 -525 16410 -505
rect 17670 -475 17690 -455
rect 17670 -525 17690 -505
rect 17910 -475 17930 -455
rect 17910 -525 17930 -505
rect 19190 -475 19210 -455
rect 19190 -525 19210 -505
<< poly >>
rect 16975 685 17015 695
rect 16975 665 16985 685
rect 17005 670 17015 685
rect 17635 685 17675 695
rect 17635 670 17645 685
rect 17005 665 17030 670
rect 16975 655 17030 665
rect 17620 665 17645 670
rect 17665 665 17675 685
rect 17620 655 17675 665
rect 17925 685 17965 695
rect 17925 665 17935 685
rect 17955 670 17965 685
rect 18585 685 18625 695
rect 18585 670 18595 685
rect 17955 665 17980 670
rect 17925 655 17980 665
rect 18570 665 18595 670
rect 18615 665 18625 685
rect 18570 655 18625 665
rect 17015 640 17030 655
rect 17070 640 17085 655
rect 17125 640 17140 655
rect 17180 640 17195 655
rect 17235 640 17250 655
rect 17290 640 17305 655
rect 17345 640 17360 655
rect 17400 640 17415 655
rect 17455 640 17470 655
rect 17510 640 17525 655
rect 17565 640 17580 655
rect 17620 640 17635 655
rect 17965 640 17980 655
rect 18020 640 18035 655
rect 18075 640 18090 655
rect 18130 640 18145 655
rect 18185 640 18200 655
rect 18240 640 18255 655
rect 18295 640 18310 655
rect 18350 640 18365 655
rect 18405 640 18420 655
rect 18460 640 18475 655
rect 18515 640 18530 655
rect 18570 640 18585 655
rect 17015 525 17030 540
rect 17070 525 17085 540
rect 17125 525 17140 540
rect 17180 525 17195 540
rect 17235 525 17250 540
rect 17290 525 17305 540
rect 17345 525 17360 540
rect 17400 525 17415 540
rect 17455 525 17470 540
rect 17510 525 17525 540
rect 17565 525 17580 540
rect 17620 525 17635 540
rect 17965 525 17980 540
rect 18020 525 18035 540
rect 18075 525 18090 540
rect 18130 525 18145 540
rect 18185 525 18200 540
rect 18240 525 18255 540
rect 18295 525 18310 540
rect 18350 525 18365 540
rect 18405 525 18420 540
rect 18460 525 18475 540
rect 18515 525 18530 540
rect 18570 525 18585 540
rect 17063 516 17092 525
rect 17063 499 17069 516
rect 17086 499 17092 516
rect 17063 490 17092 499
rect 17118 516 17147 525
rect 17118 499 17124 516
rect 17141 499 17147 516
rect 17118 490 17147 499
rect 17173 516 17202 525
rect 17173 499 17179 516
rect 17196 499 17202 516
rect 17173 490 17202 499
rect 17228 516 17257 525
rect 17228 499 17234 516
rect 17251 499 17257 516
rect 17228 490 17257 499
rect 17283 516 17312 525
rect 17283 499 17289 516
rect 17306 499 17312 516
rect 17283 490 17312 499
rect 17338 516 17367 525
rect 17338 499 17344 516
rect 17361 499 17367 516
rect 17338 490 17367 499
rect 17393 516 17422 525
rect 17393 499 17399 516
rect 17416 499 17422 516
rect 17393 490 17422 499
rect 17448 516 17477 525
rect 17448 499 17454 516
rect 17471 499 17477 516
rect 17448 490 17477 499
rect 17503 516 17532 525
rect 17503 499 17509 516
rect 17526 499 17532 516
rect 17503 490 17532 499
rect 17558 516 17587 525
rect 17558 499 17564 516
rect 17581 499 17587 516
rect 17558 490 17587 499
rect 18013 516 18042 525
rect 18013 499 18019 516
rect 18036 499 18042 516
rect 18013 490 18042 499
rect 18068 516 18097 525
rect 18068 499 18074 516
rect 18091 499 18097 516
rect 18068 490 18097 499
rect 18123 516 18152 525
rect 18123 499 18129 516
rect 18146 499 18152 516
rect 18123 490 18152 499
rect 18178 516 18207 525
rect 18178 499 18184 516
rect 18201 499 18207 516
rect 18178 490 18207 499
rect 18233 516 18262 525
rect 18233 499 18239 516
rect 18256 499 18262 516
rect 18233 490 18262 499
rect 18288 516 18317 525
rect 18288 499 18294 516
rect 18311 499 18317 516
rect 18288 490 18317 499
rect 18343 516 18372 525
rect 18343 499 18349 516
rect 18366 499 18372 516
rect 18343 490 18372 499
rect 18398 516 18427 525
rect 18398 499 18404 516
rect 18421 499 18427 516
rect 18398 490 18427 499
rect 18453 516 18482 525
rect 18453 499 18459 516
rect 18476 499 18482 516
rect 18453 490 18482 499
rect 18508 516 18537 525
rect 18508 499 18514 516
rect 18531 499 18537 516
rect 18508 490 18537 499
rect 16970 385 17010 395
rect 16970 365 16980 385
rect 17000 370 17010 385
rect 18590 385 18630 395
rect 18590 370 18600 385
rect 17000 365 17060 370
rect 16970 355 17060 365
rect 18540 365 18600 370
rect 18620 365 18630 385
rect 18540 355 18630 365
rect 17010 340 17060 355
rect 17100 340 17150 355
rect 17190 340 17240 355
rect 17280 340 17330 355
rect 17370 340 17420 355
rect 17460 340 17510 355
rect 17550 340 17600 355
rect 17640 340 17690 355
rect 17730 340 17780 355
rect 17820 340 17870 355
rect 17910 340 17960 355
rect 18000 340 18050 355
rect 18090 340 18140 355
rect 18180 340 18230 355
rect 18270 340 18320 355
rect 18360 340 18410 355
rect 18450 340 18500 355
rect 18540 340 18590 355
rect 16440 285 16470 295
rect 16440 265 16445 285
rect 16465 265 16470 285
rect 16660 285 16690 295
rect 16660 265 16665 285
rect 16685 265 16690 285
rect 16440 250 16490 265
rect 16475 240 16490 250
rect 16530 240 16545 255
rect 16585 240 16600 255
rect 16640 250 16690 265
rect 16640 240 16655 250
rect 16475 125 16490 140
rect 16530 130 16545 140
rect 16585 130 16600 140
rect 16530 115 16600 130
rect 16640 125 16655 140
rect 16545 95 16555 115
rect 16575 95 16585 115
rect 16545 85 16585 95
rect 17010 25 17060 40
rect 17100 20 17150 40
rect 17190 25 17240 40
rect 17280 25 17330 40
rect 17370 25 17420 40
rect 17460 25 17510 40
rect 17550 25 17600 40
rect 17640 25 17690 40
rect 17730 25 17780 40
rect 17820 25 17870 40
rect 17910 25 17960 40
rect 18000 25 18050 40
rect 18090 25 18140 40
rect 18180 25 18230 40
rect 18270 25 18320 40
rect 18360 25 18410 40
rect 18450 25 18500 40
rect 18540 25 18590 40
rect 17110 15 17145 20
rect 17110 -5 17115 15
rect 17135 -5 17145 15
rect 17110 -15 17145 -5
rect 17195 15 17235 25
rect 17195 -5 17205 15
rect 17225 -5 17235 15
rect 17195 -15 17235 -5
rect 17285 15 17325 25
rect 17285 -5 17295 15
rect 17315 -5 17325 15
rect 17285 -15 17325 -5
rect 17375 15 17415 25
rect 17375 -5 17385 15
rect 17405 -5 17415 15
rect 17375 -15 17415 -5
rect 17465 15 17505 25
rect 17465 -5 17475 15
rect 17495 -5 17505 15
rect 17465 -15 17505 -5
rect 17555 15 17595 25
rect 17555 -5 17565 15
rect 17585 -5 17595 15
rect 17555 -15 17595 -5
rect 17645 15 17685 25
rect 17645 -5 17655 15
rect 17675 -5 17685 15
rect 17645 -15 17685 -5
rect 17735 15 17770 25
rect 17735 -5 17745 15
rect 17765 -5 17770 15
rect 17735 -15 17770 -5
rect 17830 15 17865 25
rect 17830 -5 17835 15
rect 17855 -5 17865 15
rect 17830 -15 17865 -5
rect 17915 15 17955 25
rect 17915 -5 17925 15
rect 17945 -5 17955 15
rect 17915 -15 17955 -5
rect 18005 15 18045 25
rect 18005 -5 18015 15
rect 18035 -5 18045 15
rect 18005 -15 18045 -5
rect 18095 15 18135 25
rect 18095 -5 18105 15
rect 18125 -5 18135 15
rect 18095 -15 18135 -5
rect 18185 15 18225 25
rect 18185 -5 18195 15
rect 18215 -5 18225 15
rect 18185 -15 18225 -5
rect 18275 15 18315 25
rect 18275 -5 18285 15
rect 18305 -5 18315 15
rect 18275 -15 18315 -5
rect 18365 15 18405 25
rect 18365 -5 18375 15
rect 18395 -5 18405 15
rect 18365 -15 18405 -5
rect 18455 15 18490 25
rect 18455 -5 18465 15
rect 18485 -5 18490 15
rect 18455 -15 18490 -5
rect 16425 -395 16455 -385
rect 16425 -415 16430 -395
rect 16450 -410 16455 -395
rect 17625 -395 17655 -385
rect 17625 -410 17630 -395
rect 16450 -415 16480 -410
rect 16425 -425 16480 -415
rect 17600 -415 17630 -410
rect 17650 -415 17655 -395
rect 17600 -425 17655 -415
rect 17945 -395 17975 -385
rect 17945 -415 17950 -395
rect 17970 -410 17975 -395
rect 19145 -395 19175 -385
rect 19145 -410 19150 -395
rect 17970 -415 18000 -410
rect 17945 -425 18000 -415
rect 19120 -415 19150 -410
rect 19170 -415 19175 -395
rect 19120 -425 19175 -415
rect 16460 -440 16480 -425
rect 16520 -440 16540 -425
rect 16580 -440 16600 -425
rect 16640 -440 16660 -425
rect 16700 -440 16720 -425
rect 16760 -440 16780 -425
rect 16820 -440 16840 -425
rect 16880 -440 16900 -425
rect 16940 -440 16960 -425
rect 17000 -440 17020 -425
rect 17060 -440 17080 -425
rect 17120 -440 17140 -425
rect 17180 -440 17200 -425
rect 17240 -440 17260 -425
rect 17300 -440 17320 -425
rect 17360 -440 17380 -425
rect 17420 -440 17440 -425
rect 17480 -440 17500 -425
rect 17540 -440 17560 -425
rect 17600 -440 17620 -425
rect 17980 -440 18000 -425
rect 18040 -440 18060 -425
rect 18100 -440 18120 -425
rect 18160 -440 18180 -425
rect 18220 -440 18240 -425
rect 18280 -440 18300 -425
rect 18340 -440 18360 -425
rect 18400 -440 18420 -425
rect 18460 -440 18480 -425
rect 18520 -440 18540 -425
rect 18580 -440 18600 -425
rect 18640 -440 18660 -425
rect 18700 -440 18720 -425
rect 18760 -440 18780 -425
rect 18820 -440 18840 -425
rect 18880 -440 18900 -425
rect 18940 -440 18960 -425
rect 19000 -440 19020 -425
rect 19060 -440 19080 -425
rect 19120 -440 19140 -425
rect 16460 -555 16480 -540
rect 16520 -560 16540 -540
rect 16580 -550 16600 -540
rect 16640 -550 16660 -540
rect 16700 -550 16720 -540
rect 16760 -550 16780 -540
rect 16515 -570 16545 -560
rect 16580 -565 16780 -550
rect 16820 -550 16840 -540
rect 16880 -550 16900 -540
rect 16820 -565 16900 -550
rect 16940 -550 16960 -540
rect 17000 -550 17020 -540
rect 17060 -550 17080 -540
rect 17120 -550 17140 -540
rect 16940 -565 17140 -550
rect 17180 -550 17200 -540
rect 17240 -550 17260 -540
rect 17180 -565 17260 -550
rect 17300 -550 17320 -540
rect 17360 -550 17380 -540
rect 17420 -550 17440 -540
rect 17480 -550 17500 -540
rect 17300 -565 17500 -550
rect 17540 -555 17560 -540
rect 17600 -555 17620 -540
rect 17980 -555 18000 -540
rect 18040 -555 18060 -540
rect 18100 -550 18120 -540
rect 18160 -550 18180 -540
rect 18220 -550 18240 -540
rect 18280 -550 18300 -540
rect 17535 -565 17565 -555
rect 16515 -590 16520 -570
rect 16540 -590 16545 -570
rect 16515 -600 16545 -590
rect 16600 -585 16610 -565
rect 16630 -585 16640 -565
rect 16600 -595 16640 -585
rect 16845 -585 16850 -565
rect 16870 -585 16875 -565
rect 16845 -595 16875 -585
rect 16960 -585 16970 -565
rect 16990 -585 17000 -565
rect 16960 -595 17000 -585
rect 17205 -585 17210 -565
rect 17230 -585 17235 -565
rect 17205 -595 17235 -585
rect 17320 -585 17330 -565
rect 17350 -585 17360 -565
rect 17320 -595 17360 -585
rect 17535 -585 17540 -565
rect 17560 -585 17565 -565
rect 17535 -595 17565 -585
rect 18035 -565 18065 -555
rect 18100 -565 18300 -550
rect 18340 -550 18360 -540
rect 18400 -550 18420 -540
rect 18340 -565 18420 -550
rect 18460 -550 18480 -540
rect 18520 -550 18540 -540
rect 18580 -550 18600 -540
rect 18640 -550 18660 -540
rect 18460 -565 18660 -550
rect 18700 -550 18720 -540
rect 18760 -550 18780 -540
rect 18700 -565 18780 -550
rect 18820 -550 18840 -540
rect 18880 -550 18900 -540
rect 18940 -550 18960 -540
rect 19000 -550 19020 -540
rect 18820 -565 19020 -550
rect 19060 -560 19080 -540
rect 19120 -555 19140 -540
rect 18035 -585 18040 -565
rect 18060 -585 18065 -565
rect 18035 -595 18065 -585
rect 18240 -585 18250 -565
rect 18270 -585 18280 -565
rect 18240 -595 18280 -585
rect 18365 -585 18370 -565
rect 18390 -585 18395 -565
rect 18365 -595 18395 -585
rect 18600 -585 18610 -565
rect 18630 -585 18640 -565
rect 18600 -595 18640 -585
rect 18725 -585 18730 -565
rect 18750 -585 18755 -565
rect 18725 -595 18755 -585
rect 18960 -585 18970 -565
rect 18990 -585 19000 -565
rect 18960 -595 19000 -585
rect 19055 -570 19085 -560
rect 19055 -590 19060 -570
rect 19080 -590 19085 -570
rect 19055 -600 19085 -590
rect 17007 -760 17037 -750
rect 17007 -775 17012 -760
rect 17000 -780 17012 -775
rect 17032 -780 17037 -760
rect 17000 -790 17037 -780
rect 18563 -760 18593 -750
rect 18563 -780 18568 -760
rect 18588 -775 18593 -760
rect 18588 -780 18600 -775
rect 18563 -790 18600 -780
rect 17000 -805 17020 -790
rect 17060 -805 17080 -790
rect 18520 -805 18540 -790
rect 18580 -805 18600 -790
rect 17000 -1070 17020 -1055
rect 17060 -1070 17080 -1055
rect 18520 -1070 18540 -1055
rect 18580 -1070 18600 -1055
rect 17060 -1080 17105 -1070
rect 17060 -1100 17080 -1080
rect 17100 -1100 17105 -1080
rect 17060 -1110 17105 -1100
rect 18440 -1080 18540 -1070
rect 18440 -1100 18445 -1080
rect 18465 -1085 18540 -1080
rect 18465 -1100 18470 -1085
rect 18440 -1110 18470 -1100
rect 16620 -1270 16660 -1260
rect 16620 -1290 16630 -1270
rect 16650 -1290 16660 -1270
rect 16620 -1300 16660 -1290
rect 16740 -1270 16780 -1260
rect 16740 -1290 16750 -1270
rect 16770 -1290 16780 -1270
rect 16740 -1300 16780 -1290
rect 16860 -1270 16900 -1260
rect 16860 -1290 16870 -1270
rect 16890 -1290 16900 -1270
rect 16860 -1300 16900 -1290
rect 16980 -1270 17020 -1260
rect 16980 -1290 16990 -1270
rect 17010 -1290 17020 -1270
rect 16980 -1300 17020 -1290
rect 17300 -1270 17340 -1260
rect 17300 -1290 17310 -1270
rect 17330 -1290 17340 -1270
rect 17300 -1300 17340 -1290
rect 17420 -1270 17460 -1260
rect 17420 -1290 17430 -1270
rect 17450 -1290 17460 -1270
rect 17420 -1300 17460 -1290
rect 17540 -1270 17580 -1260
rect 17540 -1290 17550 -1270
rect 17570 -1290 17580 -1270
rect 17540 -1300 17580 -1290
rect 18020 -1270 18060 -1260
rect 18020 -1290 18030 -1270
rect 18050 -1290 18060 -1270
rect 18020 -1300 18060 -1290
rect 18140 -1270 18180 -1260
rect 18140 -1290 18150 -1270
rect 18170 -1290 18180 -1270
rect 18140 -1300 18180 -1290
rect 18260 -1270 18300 -1260
rect 18260 -1290 18270 -1270
rect 18290 -1290 18300 -1270
rect 18260 -1300 18300 -1290
rect 18580 -1270 18620 -1260
rect 18580 -1290 18590 -1270
rect 18610 -1290 18620 -1270
rect 18580 -1300 18620 -1290
rect 18700 -1270 18740 -1260
rect 18700 -1290 18710 -1270
rect 18730 -1290 18740 -1270
rect 18700 -1300 18740 -1290
rect 18820 -1270 18860 -1260
rect 18820 -1290 18830 -1270
rect 18850 -1290 18860 -1270
rect 18820 -1300 18860 -1290
rect 18940 -1270 18980 -1260
rect 18940 -1290 18950 -1270
rect 18970 -1290 18980 -1270
rect 18940 -1300 18980 -1290
rect 16570 -1315 17070 -1300
rect 17190 -1315 17690 -1300
rect 17910 -1315 18410 -1300
rect 18530 -1315 19030 -1300
rect 16570 -1580 17070 -1565
rect 17190 -1580 17690 -1565
rect 17910 -1580 18410 -1565
rect 18530 -1580 19030 -1565
rect 16820 -1725 16860 -1715
rect 16820 -1745 16830 -1725
rect 16850 -1745 16860 -1725
rect 16820 -1755 16860 -1745
rect 16900 -1725 16940 -1715
rect 16900 -1745 16910 -1725
rect 16930 -1745 16940 -1725
rect 16900 -1755 16940 -1745
rect 16980 -1725 17020 -1715
rect 16980 -1745 16990 -1725
rect 17010 -1745 17020 -1725
rect 16980 -1755 17020 -1745
rect 17060 -1725 17100 -1715
rect 17060 -1745 17070 -1725
rect 17090 -1745 17100 -1725
rect 17060 -1755 17100 -1745
rect 17140 -1725 17180 -1715
rect 17140 -1745 17150 -1725
rect 17170 -1745 17180 -1725
rect 17140 -1755 17180 -1745
rect 17220 -1725 17260 -1715
rect 17220 -1745 17230 -1725
rect 17250 -1745 17260 -1725
rect 17220 -1755 17260 -1745
rect 17300 -1725 17340 -1715
rect 17300 -1745 17310 -1725
rect 17330 -1745 17340 -1725
rect 17300 -1755 17340 -1745
rect 17380 -1725 17420 -1715
rect 17380 -1745 17390 -1725
rect 17410 -1745 17420 -1725
rect 17380 -1755 17420 -1745
rect 17460 -1725 17500 -1715
rect 17460 -1745 17470 -1725
rect 17490 -1745 17500 -1725
rect 17460 -1755 17500 -1745
rect 17540 -1725 17580 -1715
rect 17540 -1745 17550 -1725
rect 17570 -1745 17580 -1725
rect 17540 -1755 17580 -1745
rect 17620 -1725 17660 -1715
rect 17620 -1745 17630 -1725
rect 17650 -1745 17660 -1725
rect 17620 -1755 17660 -1745
rect 17700 -1725 17740 -1715
rect 17700 -1745 17710 -1725
rect 17730 -1745 17740 -1725
rect 17700 -1755 17740 -1745
rect 17860 -1725 17900 -1715
rect 17860 -1745 17870 -1725
rect 17890 -1745 17900 -1725
rect 17860 -1755 17900 -1745
rect 17940 -1725 17980 -1715
rect 17940 -1745 17950 -1725
rect 17970 -1745 17980 -1725
rect 17940 -1755 17980 -1745
rect 18020 -1725 18060 -1715
rect 18020 -1745 18030 -1725
rect 18050 -1745 18060 -1725
rect 18020 -1755 18060 -1745
rect 18100 -1725 18140 -1715
rect 18100 -1745 18110 -1725
rect 18130 -1745 18140 -1725
rect 18100 -1755 18140 -1745
rect 18180 -1725 18220 -1715
rect 18180 -1745 18190 -1725
rect 18210 -1745 18220 -1725
rect 18180 -1755 18220 -1745
rect 18260 -1725 18300 -1715
rect 18260 -1745 18270 -1725
rect 18290 -1745 18300 -1725
rect 18260 -1755 18300 -1745
rect 18340 -1725 18380 -1715
rect 18340 -1745 18350 -1725
rect 18370 -1745 18380 -1725
rect 18340 -1755 18380 -1745
rect 18420 -1725 18460 -1715
rect 18420 -1745 18430 -1725
rect 18450 -1745 18460 -1725
rect 18420 -1755 18460 -1745
rect 18500 -1725 18540 -1715
rect 18500 -1745 18510 -1725
rect 18530 -1745 18540 -1725
rect 18500 -1755 18540 -1745
rect 18580 -1725 18620 -1715
rect 18580 -1745 18590 -1725
rect 18610 -1745 18620 -1725
rect 18580 -1755 18620 -1745
rect 18660 -1725 18700 -1715
rect 18660 -1745 18670 -1725
rect 18690 -1745 18700 -1725
rect 18660 -1755 18700 -1745
rect 18740 -1725 18780 -1715
rect 18740 -1745 18750 -1725
rect 18770 -1745 18780 -1725
rect 18740 -1755 18780 -1745
rect 16780 -1770 17780 -1755
rect 17820 -1770 18820 -1755
rect 16780 -1885 17780 -1870
rect 17820 -1885 18820 -1870
<< polycont >>
rect 16985 665 17005 685
rect 17645 665 17665 685
rect 17935 665 17955 685
rect 18595 665 18615 685
rect 17069 499 17086 516
rect 17124 499 17141 516
rect 17179 499 17196 516
rect 17234 499 17251 516
rect 17289 499 17306 516
rect 17344 499 17361 516
rect 17399 499 17416 516
rect 17454 499 17471 516
rect 17509 499 17526 516
rect 17564 499 17581 516
rect 18019 499 18036 516
rect 18074 499 18091 516
rect 18129 499 18146 516
rect 18184 499 18201 516
rect 18239 499 18256 516
rect 18294 499 18311 516
rect 18349 499 18366 516
rect 18404 499 18421 516
rect 18459 499 18476 516
rect 18514 499 18531 516
rect 16980 365 17000 385
rect 18600 365 18620 385
rect 16445 265 16465 285
rect 16665 265 16685 285
rect 16555 95 16575 115
rect 17115 -5 17135 15
rect 17205 -5 17225 15
rect 17295 -5 17315 15
rect 17385 -5 17405 15
rect 17475 -5 17495 15
rect 17565 -5 17585 15
rect 17655 -5 17675 15
rect 17745 -5 17765 15
rect 17835 -5 17855 15
rect 17925 -5 17945 15
rect 18015 -5 18035 15
rect 18105 -5 18125 15
rect 18195 -5 18215 15
rect 18285 -5 18305 15
rect 18375 -5 18395 15
rect 18465 -5 18485 15
rect 16430 -415 16450 -395
rect 17630 -415 17650 -395
rect 17950 -415 17970 -395
rect 19150 -415 19170 -395
rect 16520 -590 16540 -570
rect 16610 -585 16630 -565
rect 16850 -585 16870 -565
rect 16970 -585 16990 -565
rect 17210 -585 17230 -565
rect 17330 -585 17350 -565
rect 17540 -585 17560 -565
rect 18040 -585 18060 -565
rect 18250 -585 18270 -565
rect 18370 -585 18390 -565
rect 18610 -585 18630 -565
rect 18730 -585 18750 -565
rect 18970 -585 18990 -565
rect 19060 -590 19080 -570
rect 17012 -780 17032 -760
rect 18568 -780 18588 -760
rect 17080 -1100 17100 -1080
rect 18445 -1100 18465 -1080
rect 16630 -1290 16650 -1270
rect 16750 -1290 16770 -1270
rect 16870 -1290 16890 -1270
rect 16990 -1290 17010 -1270
rect 17310 -1290 17330 -1270
rect 17430 -1290 17450 -1270
rect 17550 -1290 17570 -1270
rect 18030 -1290 18050 -1270
rect 18150 -1290 18170 -1270
rect 18270 -1290 18290 -1270
rect 18590 -1290 18610 -1270
rect 18710 -1290 18730 -1270
rect 18830 -1290 18850 -1270
rect 18950 -1290 18970 -1270
rect 16830 -1745 16850 -1725
rect 16910 -1745 16930 -1725
rect 16990 -1745 17010 -1725
rect 17070 -1745 17090 -1725
rect 17150 -1745 17170 -1725
rect 17230 -1745 17250 -1725
rect 17310 -1745 17330 -1725
rect 17390 -1745 17410 -1725
rect 17470 -1745 17490 -1725
rect 17550 -1745 17570 -1725
rect 17630 -1745 17650 -1725
rect 17710 -1745 17730 -1725
rect 17870 -1745 17890 -1725
rect 17950 -1745 17970 -1725
rect 18030 -1745 18050 -1725
rect 18110 -1745 18130 -1725
rect 18190 -1745 18210 -1725
rect 18270 -1745 18290 -1725
rect 18350 -1745 18370 -1725
rect 18430 -1745 18450 -1725
rect 18510 -1745 18530 -1725
rect 18590 -1745 18610 -1725
rect 18670 -1745 18690 -1725
rect 18750 -1745 18770 -1725
<< xpolycontact >>
rect 17470 -2035 17690 -2000
rect 17904 -2035 18124 -2000
rect 16485 -3160 16520 -2940
rect 16100 -3481 16135 -3261
rect 16100 -3889 16135 -3670
rect 16210 -3585 16245 -3365
rect 16210 -3889 16245 -3669
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19185 -3350 19220 -3130
rect 19185 -3889 19220 -3669
rect 19245 -3350 19280 -3130
rect 19245 -3889 19280 -3669
rect 19305 -3350 19340 -3130
rect 19305 -3889 19340 -3669
rect 19465 -3376 19500 -3156
rect 19465 -3784 19500 -3565
<< ppolyres >>
rect 16100 -3670 16135 -3481
rect 19465 -3565 19500 -3376
<< xpolyres >>
rect 17690 -2035 17904 -2000
rect 16210 -3669 16245 -3585
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19185 -3669 19220 -3350
rect 19245 -3669 19280 -3350
rect 19305 -3669 19340 -3350
<< locali >>
rect 16975 685 17015 695
rect 16975 665 16985 685
rect 17005 665 17015 685
rect 16975 655 17015 665
rect 17635 685 17675 695
rect 17635 665 17645 685
rect 17665 665 17675 685
rect 17635 655 17675 665
rect 17925 685 17965 695
rect 17925 665 17935 685
rect 17955 665 17965 685
rect 17925 655 17965 665
rect 18585 685 18625 695
rect 18585 665 18595 685
rect 18615 665 18625 685
rect 18585 655 18625 665
rect 16940 625 17010 635
rect 16940 605 16945 625
rect 16965 605 16985 625
rect 17005 605 17010 625
rect 16940 575 17010 605
rect 16940 555 16945 575
rect 16965 555 16985 575
rect 17005 555 17010 575
rect 16940 545 17010 555
rect 17035 625 17065 635
rect 17035 605 17040 625
rect 17060 605 17065 625
rect 17035 575 17065 605
rect 17035 555 17040 575
rect 17060 555 17065 575
rect 17035 545 17065 555
rect 17090 625 17120 635
rect 17090 605 17095 625
rect 17115 605 17120 625
rect 17090 575 17120 605
rect 17090 555 17095 575
rect 17115 555 17120 575
rect 17090 545 17120 555
rect 17145 625 17175 635
rect 17145 605 17150 625
rect 17170 605 17175 625
rect 17145 575 17175 605
rect 17145 555 17150 575
rect 17170 555 17175 575
rect 17145 545 17175 555
rect 17200 625 17230 635
rect 17200 605 17205 625
rect 17225 605 17230 625
rect 17200 575 17230 605
rect 17200 555 17205 575
rect 17225 555 17230 575
rect 17200 545 17230 555
rect 17255 625 17285 635
rect 17255 605 17260 625
rect 17280 605 17285 625
rect 17255 575 17285 605
rect 17255 555 17260 575
rect 17280 555 17285 575
rect 17255 545 17285 555
rect 17310 625 17340 635
rect 17310 605 17315 625
rect 17335 605 17340 625
rect 17310 575 17340 605
rect 17310 555 17315 575
rect 17335 555 17340 575
rect 17310 545 17340 555
rect 17365 625 17395 635
rect 17365 605 17370 625
rect 17390 605 17395 625
rect 17365 575 17395 605
rect 17365 555 17370 575
rect 17390 555 17395 575
rect 17365 545 17395 555
rect 17420 625 17450 635
rect 17420 605 17425 625
rect 17445 605 17450 625
rect 17420 575 17450 605
rect 17420 555 17425 575
rect 17445 555 17450 575
rect 17420 545 17450 555
rect 17475 625 17505 635
rect 17475 605 17480 625
rect 17500 605 17505 625
rect 17475 575 17505 605
rect 17475 555 17480 575
rect 17500 555 17505 575
rect 17475 545 17505 555
rect 17530 625 17560 635
rect 17530 605 17535 625
rect 17555 605 17560 625
rect 17530 575 17560 605
rect 17530 555 17535 575
rect 17555 555 17560 575
rect 17530 545 17560 555
rect 17585 625 17615 635
rect 17585 605 17590 625
rect 17610 605 17615 625
rect 17585 575 17615 605
rect 17585 555 17590 575
rect 17610 555 17615 575
rect 17585 545 17615 555
rect 17640 625 17710 635
rect 17640 605 17645 625
rect 17665 605 17685 625
rect 17705 605 17710 625
rect 17640 575 17710 605
rect 17640 555 17645 575
rect 17665 555 17685 575
rect 17705 555 17710 575
rect 17640 545 17710 555
rect 17890 625 17960 635
rect 17890 605 17895 625
rect 17915 605 17935 625
rect 17955 605 17960 625
rect 17890 575 17960 605
rect 17890 555 17895 575
rect 17915 555 17935 575
rect 17955 555 17960 575
rect 17890 545 17960 555
rect 17985 625 18015 635
rect 17985 605 17990 625
rect 18010 605 18015 625
rect 17985 575 18015 605
rect 17985 555 17990 575
rect 18010 555 18015 575
rect 17985 545 18015 555
rect 18040 625 18070 635
rect 18040 605 18045 625
rect 18065 605 18070 625
rect 18040 575 18070 605
rect 18040 555 18045 575
rect 18065 555 18070 575
rect 18040 545 18070 555
rect 18095 625 18125 635
rect 18095 605 18100 625
rect 18120 605 18125 625
rect 18095 575 18125 605
rect 18095 555 18100 575
rect 18120 555 18125 575
rect 18095 545 18125 555
rect 18150 625 18180 635
rect 18150 605 18155 625
rect 18175 605 18180 625
rect 18150 575 18180 605
rect 18150 555 18155 575
rect 18175 555 18180 575
rect 18150 545 18180 555
rect 18205 625 18235 635
rect 18205 605 18210 625
rect 18230 605 18235 625
rect 18205 575 18235 605
rect 18205 555 18210 575
rect 18230 555 18235 575
rect 18205 545 18235 555
rect 18260 625 18290 635
rect 18260 605 18265 625
rect 18285 605 18290 625
rect 18260 575 18290 605
rect 18260 555 18265 575
rect 18285 555 18290 575
rect 18260 545 18290 555
rect 18315 625 18345 635
rect 18315 605 18320 625
rect 18340 605 18345 625
rect 18315 575 18345 605
rect 18315 555 18320 575
rect 18340 555 18345 575
rect 18315 545 18345 555
rect 18370 625 18400 635
rect 18370 605 18375 625
rect 18395 605 18400 625
rect 18370 575 18400 605
rect 18370 555 18375 575
rect 18395 555 18400 575
rect 18370 545 18400 555
rect 18425 625 18455 635
rect 18425 605 18430 625
rect 18450 605 18455 625
rect 18425 575 18455 605
rect 18425 555 18430 575
rect 18450 555 18455 575
rect 18425 545 18455 555
rect 18480 625 18510 635
rect 18480 605 18485 625
rect 18505 605 18510 625
rect 18480 575 18510 605
rect 18480 555 18485 575
rect 18505 555 18510 575
rect 18480 545 18510 555
rect 18535 625 18565 635
rect 18535 605 18540 625
rect 18560 605 18565 625
rect 18535 575 18565 605
rect 18535 555 18540 575
rect 18560 555 18565 575
rect 18535 545 18565 555
rect 18590 625 18660 635
rect 18590 605 18595 625
rect 18615 605 18635 625
rect 18655 605 18660 625
rect 18590 575 18660 605
rect 18590 555 18595 575
rect 18615 555 18635 575
rect 18655 555 18660 575
rect 18590 545 18660 555
rect 17063 516 17092 525
rect 17063 499 17069 516
rect 17086 499 17092 516
rect 17063 490 17092 499
rect 17118 516 17147 525
rect 17118 499 17124 516
rect 17141 499 17147 516
rect 17118 490 17147 499
rect 17173 516 17202 525
rect 17173 499 17179 516
rect 17196 499 17202 516
rect 17173 490 17202 499
rect 17228 516 17257 525
rect 17228 499 17234 516
rect 17251 499 17257 516
rect 17228 490 17257 499
rect 17283 516 17312 525
rect 17283 499 17289 516
rect 17306 499 17312 516
rect 17283 490 17312 499
rect 17338 516 17367 525
rect 17338 499 17344 516
rect 17361 499 17367 516
rect 17338 490 17367 499
rect 17393 516 17422 525
rect 17393 499 17399 516
rect 17416 499 17422 516
rect 17393 490 17422 499
rect 17448 516 17477 525
rect 17448 499 17454 516
rect 17471 499 17477 516
rect 17448 490 17477 499
rect 17503 516 17532 525
rect 17503 499 17509 516
rect 17526 499 17532 516
rect 17503 490 17532 499
rect 17558 516 17587 525
rect 17558 499 17564 516
rect 17581 499 17587 516
rect 17558 490 17587 499
rect 18013 516 18042 525
rect 18013 499 18019 516
rect 18036 499 18042 516
rect 18013 490 18042 499
rect 18068 516 18097 525
rect 18068 499 18074 516
rect 18091 499 18097 516
rect 18068 490 18097 499
rect 18123 516 18152 525
rect 18123 499 18129 516
rect 18146 499 18152 516
rect 18123 490 18152 499
rect 18178 516 18207 525
rect 18178 499 18184 516
rect 18201 499 18207 516
rect 18178 490 18207 499
rect 18233 516 18262 525
rect 18233 499 18239 516
rect 18256 499 18262 516
rect 18233 490 18262 499
rect 18288 516 18317 525
rect 18288 499 18294 516
rect 18311 499 18317 516
rect 18288 490 18317 499
rect 18343 516 18372 525
rect 18343 499 18349 516
rect 18366 499 18372 516
rect 18343 490 18372 499
rect 18398 516 18427 525
rect 18398 499 18404 516
rect 18421 499 18427 516
rect 18398 490 18427 499
rect 18453 516 18482 525
rect 18453 499 18459 516
rect 18476 499 18482 516
rect 18453 490 18482 499
rect 18508 516 18537 525
rect 18508 499 18514 516
rect 18531 499 18537 516
rect 18508 490 18537 499
rect 16970 385 17010 395
rect 16970 365 16980 385
rect 17000 365 17010 385
rect 16970 355 17010 365
rect 17150 385 17190 395
rect 17150 365 17160 385
rect 17180 365 17190 385
rect 17150 355 17190 365
rect 17330 385 17370 395
rect 17330 365 17340 385
rect 17360 365 17370 385
rect 17330 355 17370 365
rect 17510 385 17550 395
rect 17510 365 17520 385
rect 17540 365 17550 385
rect 17510 355 17550 365
rect 17690 385 17730 395
rect 17690 365 17700 385
rect 17720 365 17730 385
rect 17690 355 17730 365
rect 17870 385 17910 395
rect 17870 365 17880 385
rect 17900 365 17910 385
rect 17870 355 17910 365
rect 18050 385 18090 395
rect 18050 365 18060 385
rect 18080 365 18090 385
rect 18050 355 18090 365
rect 18230 385 18270 395
rect 18230 365 18240 385
rect 18260 365 18270 385
rect 18230 355 18270 365
rect 18410 385 18450 395
rect 18410 365 18420 385
rect 18440 365 18450 385
rect 18410 355 18450 365
rect 18590 385 18630 395
rect 18590 365 18600 385
rect 18620 365 18630 385
rect 18590 355 18630 365
rect 16980 335 17000 355
rect 17160 335 17180 355
rect 17340 335 17360 355
rect 17520 335 17540 355
rect 17700 335 17720 355
rect 17880 335 17900 355
rect 18060 335 18080 355
rect 18240 335 18260 355
rect 18420 335 18440 355
rect 18600 335 18620 355
rect 16935 325 17005 335
rect 16935 305 16940 325
rect 16960 305 16980 325
rect 17000 305 17005 325
rect 16440 285 16470 295
rect 16440 265 16445 285
rect 16465 265 16470 285
rect 16440 255 16470 265
rect 16545 285 16585 295
rect 16545 265 16555 285
rect 16575 265 16585 285
rect 16545 255 16585 265
rect 16655 285 16695 295
rect 16655 265 16665 285
rect 16685 265 16695 285
rect 16655 255 16695 265
rect 16935 275 17005 305
rect 16935 255 16940 275
rect 16960 255 16980 275
rect 17000 255 17005 275
rect 16400 225 16470 235
rect 16400 205 16405 225
rect 16425 205 16445 225
rect 16465 205 16470 225
rect 16400 175 16470 205
rect 16400 155 16405 175
rect 16425 155 16445 175
rect 16465 155 16470 175
rect 16400 145 16470 155
rect 16495 225 16525 235
rect 16495 205 16500 225
rect 16520 205 16525 225
rect 16495 175 16525 205
rect 16495 155 16500 175
rect 16520 155 16525 175
rect 16495 145 16525 155
rect 16550 225 16580 235
rect 16550 205 16555 225
rect 16575 205 16580 225
rect 16550 175 16580 205
rect 16550 155 16555 175
rect 16575 155 16580 175
rect 16550 145 16580 155
rect 16605 225 16635 235
rect 16605 205 16610 225
rect 16630 205 16635 225
rect 16605 175 16635 205
rect 16605 155 16610 175
rect 16630 155 16635 175
rect 16605 145 16635 155
rect 16660 225 16735 235
rect 16660 205 16665 225
rect 16685 205 16710 225
rect 16730 205 16735 225
rect 16660 175 16735 205
rect 16660 155 16665 175
rect 16685 155 16710 175
rect 16730 155 16735 175
rect 16660 145 16735 155
rect 16935 225 17005 255
rect 16935 205 16940 225
rect 16960 205 16980 225
rect 17000 205 17005 225
rect 16935 175 17005 205
rect 16935 155 16940 175
rect 16960 155 16980 175
rect 17000 155 17005 175
rect 16935 125 17005 155
rect 16485 115 16525 125
rect 16485 95 16495 115
rect 16515 95 16525 115
rect 16485 85 16525 95
rect 16545 115 16585 125
rect 16545 95 16555 115
rect 16575 95 16585 115
rect 16545 85 16585 95
rect 16605 115 16645 125
rect 16605 95 16615 115
rect 16635 95 16645 115
rect 16605 85 16645 95
rect 16935 105 16940 125
rect 16960 105 16980 125
rect 17000 105 17005 125
rect 16935 75 17005 105
rect 16935 55 16940 75
rect 16960 55 16980 75
rect 17000 55 17005 75
rect 16935 45 17005 55
rect 17065 325 17095 335
rect 17065 305 17070 325
rect 17090 305 17095 325
rect 17065 275 17095 305
rect 17065 255 17070 275
rect 17090 255 17095 275
rect 17065 225 17095 255
rect 17065 205 17070 225
rect 17090 205 17095 225
rect 17065 175 17095 205
rect 17065 155 17070 175
rect 17090 155 17095 175
rect 17065 125 17095 155
rect 17065 105 17070 125
rect 17090 105 17095 125
rect 17065 75 17095 105
rect 17065 55 17070 75
rect 17090 55 17095 75
rect 17065 45 17095 55
rect 17155 325 17185 335
rect 17155 305 17160 325
rect 17180 305 17185 325
rect 17155 275 17185 305
rect 17155 255 17160 275
rect 17180 255 17185 275
rect 17155 225 17185 255
rect 17155 205 17160 225
rect 17180 205 17185 225
rect 17155 175 17185 205
rect 17155 155 17160 175
rect 17180 155 17185 175
rect 17155 125 17185 155
rect 17155 105 17160 125
rect 17180 105 17185 125
rect 17155 75 17185 105
rect 17155 55 17160 75
rect 17180 55 17185 75
rect 17155 45 17185 55
rect 17245 325 17275 335
rect 17245 305 17250 325
rect 17270 305 17275 325
rect 17245 275 17275 305
rect 17245 255 17250 275
rect 17270 255 17275 275
rect 17245 225 17275 255
rect 17245 205 17250 225
rect 17270 205 17275 225
rect 17245 175 17275 205
rect 17245 155 17250 175
rect 17270 155 17275 175
rect 17245 125 17275 155
rect 17245 105 17250 125
rect 17270 105 17275 125
rect 17245 75 17275 105
rect 17245 55 17250 75
rect 17270 55 17275 75
rect 17245 45 17275 55
rect 17335 325 17365 335
rect 17335 305 17340 325
rect 17360 305 17365 325
rect 17335 275 17365 305
rect 17335 255 17340 275
rect 17360 255 17365 275
rect 17335 225 17365 255
rect 17335 205 17340 225
rect 17360 205 17365 225
rect 17335 175 17365 205
rect 17335 155 17340 175
rect 17360 155 17365 175
rect 17335 125 17365 155
rect 17335 105 17340 125
rect 17360 105 17365 125
rect 17335 75 17365 105
rect 17335 55 17340 75
rect 17360 55 17365 75
rect 17335 45 17365 55
rect 17425 325 17455 335
rect 17425 305 17430 325
rect 17450 305 17455 325
rect 17425 275 17455 305
rect 17425 255 17430 275
rect 17450 255 17455 275
rect 17425 225 17455 255
rect 17425 205 17430 225
rect 17450 205 17455 225
rect 17425 175 17455 205
rect 17425 155 17430 175
rect 17450 155 17455 175
rect 17425 125 17455 155
rect 17425 105 17430 125
rect 17450 105 17455 125
rect 17425 75 17455 105
rect 17425 55 17430 75
rect 17450 55 17455 75
rect 17425 45 17455 55
rect 17515 325 17545 335
rect 17515 305 17520 325
rect 17540 305 17545 325
rect 17515 275 17545 305
rect 17515 255 17520 275
rect 17540 255 17545 275
rect 17515 225 17545 255
rect 17515 205 17520 225
rect 17540 205 17545 225
rect 17515 175 17545 205
rect 17515 155 17520 175
rect 17540 155 17545 175
rect 17515 125 17545 155
rect 17515 105 17520 125
rect 17540 105 17545 125
rect 17515 75 17545 105
rect 17515 55 17520 75
rect 17540 55 17545 75
rect 17515 45 17545 55
rect 17605 325 17635 335
rect 17605 305 17610 325
rect 17630 305 17635 325
rect 17605 275 17635 305
rect 17605 255 17610 275
rect 17630 255 17635 275
rect 17605 225 17635 255
rect 17605 205 17610 225
rect 17630 205 17635 225
rect 17605 175 17635 205
rect 17605 155 17610 175
rect 17630 155 17635 175
rect 17605 125 17635 155
rect 17605 105 17610 125
rect 17630 105 17635 125
rect 17605 75 17635 105
rect 17605 55 17610 75
rect 17630 55 17635 75
rect 17605 45 17635 55
rect 17695 325 17725 335
rect 17695 305 17700 325
rect 17720 305 17725 325
rect 17695 275 17725 305
rect 17695 255 17700 275
rect 17720 255 17725 275
rect 17695 225 17725 255
rect 17695 205 17700 225
rect 17720 205 17725 225
rect 17695 175 17725 205
rect 17695 155 17700 175
rect 17720 155 17725 175
rect 17695 125 17725 155
rect 17695 105 17700 125
rect 17720 105 17725 125
rect 17695 75 17725 105
rect 17695 55 17700 75
rect 17720 55 17725 75
rect 17695 45 17725 55
rect 17785 325 17815 335
rect 17785 305 17790 325
rect 17810 305 17815 325
rect 17785 275 17815 305
rect 17785 255 17790 275
rect 17810 255 17815 275
rect 17785 225 17815 255
rect 17785 205 17790 225
rect 17810 205 17815 225
rect 17785 175 17815 205
rect 17785 155 17790 175
rect 17810 155 17815 175
rect 17785 125 17815 155
rect 17785 105 17790 125
rect 17810 105 17815 125
rect 17785 75 17815 105
rect 17785 55 17790 75
rect 17810 55 17815 75
rect 17785 45 17815 55
rect 17875 325 17905 335
rect 17875 305 17880 325
rect 17900 305 17905 325
rect 17875 275 17905 305
rect 17875 255 17880 275
rect 17900 255 17905 275
rect 17875 225 17905 255
rect 17875 205 17880 225
rect 17900 205 17905 225
rect 17875 175 17905 205
rect 17875 155 17880 175
rect 17900 155 17905 175
rect 17875 125 17905 155
rect 17875 105 17880 125
rect 17900 105 17905 125
rect 17875 75 17905 105
rect 17875 55 17880 75
rect 17900 55 17905 75
rect 17875 45 17905 55
rect 17965 325 17995 335
rect 17965 305 17970 325
rect 17990 305 17995 325
rect 17965 275 17995 305
rect 17965 255 17970 275
rect 17990 255 17995 275
rect 17965 225 17995 255
rect 17965 205 17970 225
rect 17990 205 17995 225
rect 17965 175 17995 205
rect 17965 155 17970 175
rect 17990 155 17995 175
rect 17965 125 17995 155
rect 17965 105 17970 125
rect 17990 105 17995 125
rect 17965 75 17995 105
rect 17965 55 17970 75
rect 17990 55 17995 75
rect 17965 45 17995 55
rect 18055 325 18085 335
rect 18055 305 18060 325
rect 18080 305 18085 325
rect 18055 275 18085 305
rect 18055 255 18060 275
rect 18080 255 18085 275
rect 18055 225 18085 255
rect 18055 205 18060 225
rect 18080 205 18085 225
rect 18055 175 18085 205
rect 18055 155 18060 175
rect 18080 155 18085 175
rect 18055 125 18085 155
rect 18055 105 18060 125
rect 18080 105 18085 125
rect 18055 75 18085 105
rect 18055 55 18060 75
rect 18080 55 18085 75
rect 18055 45 18085 55
rect 18145 325 18175 335
rect 18145 305 18150 325
rect 18170 305 18175 325
rect 18145 275 18175 305
rect 18145 255 18150 275
rect 18170 255 18175 275
rect 18145 225 18175 255
rect 18145 205 18150 225
rect 18170 205 18175 225
rect 18145 175 18175 205
rect 18145 155 18150 175
rect 18170 155 18175 175
rect 18145 125 18175 155
rect 18145 105 18150 125
rect 18170 105 18175 125
rect 18145 75 18175 105
rect 18145 55 18150 75
rect 18170 55 18175 75
rect 18145 45 18175 55
rect 18235 325 18265 335
rect 18235 305 18240 325
rect 18260 305 18265 325
rect 18235 275 18265 305
rect 18235 255 18240 275
rect 18260 255 18265 275
rect 18235 225 18265 255
rect 18235 205 18240 225
rect 18260 205 18265 225
rect 18235 175 18265 205
rect 18235 155 18240 175
rect 18260 155 18265 175
rect 18235 125 18265 155
rect 18235 105 18240 125
rect 18260 105 18265 125
rect 18235 75 18265 105
rect 18235 55 18240 75
rect 18260 55 18265 75
rect 18235 45 18265 55
rect 18325 325 18355 335
rect 18325 305 18330 325
rect 18350 305 18355 325
rect 18325 275 18355 305
rect 18325 255 18330 275
rect 18350 255 18355 275
rect 18325 225 18355 255
rect 18325 205 18330 225
rect 18350 205 18355 225
rect 18325 175 18355 205
rect 18325 155 18330 175
rect 18350 155 18355 175
rect 18325 125 18355 155
rect 18325 105 18330 125
rect 18350 105 18355 125
rect 18325 75 18355 105
rect 18325 55 18330 75
rect 18350 55 18355 75
rect 18325 45 18355 55
rect 18415 325 18445 335
rect 18415 305 18420 325
rect 18440 305 18445 325
rect 18415 275 18445 305
rect 18415 255 18420 275
rect 18440 255 18445 275
rect 18415 225 18445 255
rect 18415 205 18420 225
rect 18440 205 18445 225
rect 18415 175 18445 205
rect 18415 155 18420 175
rect 18440 155 18445 175
rect 18415 125 18445 155
rect 18415 105 18420 125
rect 18440 105 18445 125
rect 18415 75 18445 105
rect 18415 55 18420 75
rect 18440 55 18445 75
rect 18415 45 18445 55
rect 18505 325 18535 335
rect 18505 305 18510 325
rect 18530 305 18535 325
rect 18505 275 18535 305
rect 18505 255 18510 275
rect 18530 255 18535 275
rect 18505 225 18535 255
rect 18505 205 18510 225
rect 18530 205 18535 225
rect 18505 175 18535 205
rect 18505 155 18510 175
rect 18530 155 18535 175
rect 18505 125 18535 155
rect 18505 105 18510 125
rect 18530 105 18535 125
rect 18505 75 18535 105
rect 18505 55 18510 75
rect 18530 55 18535 75
rect 18505 45 18535 55
rect 18595 325 18665 335
rect 18595 305 18600 325
rect 18620 305 18640 325
rect 18660 305 18665 325
rect 18595 275 18665 305
rect 18595 255 18600 275
rect 18620 255 18640 275
rect 18660 255 18665 275
rect 18595 225 18665 255
rect 18595 205 18600 225
rect 18620 205 18640 225
rect 18660 205 18665 225
rect 18595 175 18665 205
rect 18595 155 18600 175
rect 18620 155 18640 175
rect 18660 155 18665 175
rect 18595 125 18665 155
rect 18595 105 18600 125
rect 18620 105 18640 125
rect 18660 105 18665 125
rect 18595 75 18665 105
rect 18595 55 18600 75
rect 18620 55 18640 75
rect 18660 55 18665 75
rect 18595 45 18665 55
rect 17110 15 17145 25
rect 17110 -5 17115 15
rect 17135 -5 17145 15
rect 17110 -15 17145 -5
rect 17195 15 17235 25
rect 17195 -5 17205 15
rect 17225 -5 17235 15
rect 17195 -15 17235 -5
rect 17285 15 17325 25
rect 17285 -5 17295 15
rect 17315 -5 17325 15
rect 17285 -15 17325 -5
rect 17375 15 17415 25
rect 17375 -5 17385 15
rect 17405 -5 17415 15
rect 17375 -15 17415 -5
rect 17465 15 17505 25
rect 17465 -5 17475 15
rect 17495 -5 17505 15
rect 17465 -15 17505 -5
rect 17555 15 17595 25
rect 17555 -5 17565 15
rect 17585 -5 17595 15
rect 17555 -15 17595 -5
rect 17645 15 17685 25
rect 17645 -5 17655 15
rect 17675 -5 17685 15
rect 17645 -15 17685 -5
rect 17735 15 17770 25
rect 17735 -5 17745 15
rect 17765 -5 17770 15
rect 17735 -15 17770 -5
rect 17830 15 17865 25
rect 17830 -5 17835 15
rect 17855 -5 17865 15
rect 17830 -15 17865 -5
rect 17915 15 17955 25
rect 17915 -5 17925 15
rect 17945 -5 17955 15
rect 17915 -15 17955 -5
rect 18005 15 18045 25
rect 18005 -5 18015 15
rect 18035 -5 18045 15
rect 18005 -15 18045 -5
rect 18095 15 18135 25
rect 18095 -5 18105 15
rect 18125 -5 18135 15
rect 18095 -15 18135 -5
rect 18185 15 18225 25
rect 18185 -5 18195 15
rect 18215 -5 18225 15
rect 18185 -15 18225 -5
rect 18275 15 18315 25
rect 18275 -5 18285 15
rect 18305 -5 18315 15
rect 18275 -15 18315 -5
rect 18365 15 18405 25
rect 18365 -5 18375 15
rect 18395 -5 18405 15
rect 18365 -15 18405 -5
rect 18455 15 18490 25
rect 18455 -5 18465 15
rect 18485 -5 18490 15
rect 18455 -15 18490 -5
rect 16425 -395 16455 -385
rect 16425 -415 16430 -395
rect 16450 -415 16455 -395
rect 16425 -425 16455 -415
rect 17625 -395 17655 -385
rect 17625 -415 17630 -395
rect 17650 -415 17655 -395
rect 17625 -425 17655 -415
rect 17945 -395 17975 -385
rect 17945 -415 17950 -395
rect 17970 -415 17975 -395
rect 17945 -425 17975 -415
rect 19145 -395 19175 -385
rect 19145 -415 19150 -395
rect 19170 -415 19175 -395
rect 19145 -425 19175 -415
rect 16385 -455 16455 -445
rect 16385 -475 16390 -455
rect 16410 -475 16430 -455
rect 16450 -475 16455 -455
rect 16385 -505 16455 -475
rect 16385 -525 16390 -505
rect 16410 -525 16430 -505
rect 16450 -525 16455 -505
rect 16385 -535 16455 -525
rect 16485 -455 16515 -445
rect 16485 -475 16490 -455
rect 16510 -475 16515 -455
rect 16485 -505 16515 -475
rect 16485 -525 16490 -505
rect 16510 -525 16515 -505
rect 16485 -535 16515 -525
rect 16545 -455 16575 -445
rect 16545 -475 16550 -455
rect 16570 -475 16575 -455
rect 16545 -505 16575 -475
rect 16545 -525 16550 -505
rect 16570 -525 16575 -505
rect 16545 -535 16575 -525
rect 16605 -455 16635 -445
rect 16605 -475 16610 -455
rect 16630 -475 16635 -455
rect 16605 -505 16635 -475
rect 16605 -525 16610 -505
rect 16630 -525 16635 -505
rect 16605 -535 16635 -525
rect 16665 -455 16695 -445
rect 16665 -475 16670 -455
rect 16690 -475 16695 -455
rect 16665 -505 16695 -475
rect 16665 -525 16670 -505
rect 16690 -525 16695 -505
rect 16665 -535 16695 -525
rect 16725 -455 16755 -445
rect 16725 -475 16730 -455
rect 16750 -475 16755 -455
rect 16725 -505 16755 -475
rect 16725 -525 16730 -505
rect 16750 -525 16755 -505
rect 16725 -535 16755 -525
rect 16785 -455 16815 -445
rect 16785 -475 16790 -455
rect 16810 -475 16815 -455
rect 16785 -505 16815 -475
rect 16785 -525 16790 -505
rect 16810 -525 16815 -505
rect 16785 -535 16815 -525
rect 16845 -455 16875 -445
rect 16845 -475 16850 -455
rect 16870 -475 16875 -455
rect 16845 -505 16875 -475
rect 16845 -525 16850 -505
rect 16870 -525 16875 -505
rect 16845 -535 16875 -525
rect 16905 -455 16935 -445
rect 16905 -475 16910 -455
rect 16930 -475 16935 -455
rect 16905 -505 16935 -475
rect 16905 -525 16910 -505
rect 16930 -525 16935 -505
rect 16905 -535 16935 -525
rect 16965 -455 16995 -445
rect 16965 -475 16970 -455
rect 16990 -475 16995 -455
rect 16965 -505 16995 -475
rect 16965 -525 16970 -505
rect 16990 -525 16995 -505
rect 16965 -535 16995 -525
rect 17025 -455 17055 -445
rect 17025 -475 17030 -455
rect 17050 -475 17055 -455
rect 17025 -505 17055 -475
rect 17025 -525 17030 -505
rect 17050 -525 17055 -505
rect 17025 -535 17055 -525
rect 17085 -455 17115 -445
rect 17085 -475 17090 -455
rect 17110 -475 17115 -455
rect 17085 -505 17115 -475
rect 17085 -525 17090 -505
rect 17110 -525 17115 -505
rect 17085 -535 17115 -525
rect 17145 -455 17175 -445
rect 17145 -475 17150 -455
rect 17170 -475 17175 -455
rect 17145 -505 17175 -475
rect 17145 -525 17150 -505
rect 17170 -525 17175 -505
rect 17145 -535 17175 -525
rect 17205 -455 17235 -445
rect 17205 -475 17210 -455
rect 17230 -475 17235 -455
rect 17205 -505 17235 -475
rect 17205 -525 17210 -505
rect 17230 -525 17235 -505
rect 17205 -535 17235 -525
rect 17265 -455 17295 -445
rect 17265 -475 17270 -455
rect 17290 -475 17295 -455
rect 17265 -505 17295 -475
rect 17265 -525 17270 -505
rect 17290 -525 17295 -505
rect 17265 -535 17295 -525
rect 17325 -455 17355 -445
rect 17325 -475 17330 -455
rect 17350 -475 17355 -455
rect 17325 -505 17355 -475
rect 17325 -525 17330 -505
rect 17350 -525 17355 -505
rect 17325 -535 17355 -525
rect 17385 -455 17415 -445
rect 17385 -475 17390 -455
rect 17410 -475 17415 -455
rect 17385 -505 17415 -475
rect 17385 -525 17390 -505
rect 17410 -525 17415 -505
rect 17385 -535 17415 -525
rect 17445 -455 17475 -445
rect 17445 -475 17450 -455
rect 17470 -475 17475 -455
rect 17445 -505 17475 -475
rect 17445 -525 17450 -505
rect 17470 -525 17475 -505
rect 17445 -535 17475 -525
rect 17505 -455 17535 -445
rect 17505 -475 17510 -455
rect 17530 -475 17535 -455
rect 17505 -505 17535 -475
rect 17505 -525 17510 -505
rect 17530 -525 17535 -505
rect 17505 -535 17535 -525
rect 17565 -455 17595 -445
rect 17565 -475 17570 -455
rect 17590 -475 17595 -455
rect 17565 -505 17595 -475
rect 17565 -525 17570 -505
rect 17590 -525 17595 -505
rect 17565 -535 17595 -525
rect 17625 -455 17695 -445
rect 17625 -475 17630 -455
rect 17650 -475 17670 -455
rect 17690 -475 17695 -455
rect 17625 -505 17695 -475
rect 17625 -525 17630 -505
rect 17650 -525 17670 -505
rect 17690 -525 17695 -505
rect 17625 -535 17695 -525
rect 17905 -455 17975 -445
rect 17905 -475 17910 -455
rect 17930 -475 17950 -455
rect 17970 -475 17975 -455
rect 17905 -505 17975 -475
rect 17905 -525 17910 -505
rect 17930 -525 17950 -505
rect 17970 -525 17975 -505
rect 17905 -535 17975 -525
rect 18005 -455 18035 -445
rect 18005 -475 18010 -455
rect 18030 -475 18035 -455
rect 18005 -505 18035 -475
rect 18005 -525 18010 -505
rect 18030 -525 18035 -505
rect 18005 -535 18035 -525
rect 18065 -455 18095 -445
rect 18065 -475 18070 -455
rect 18090 -475 18095 -455
rect 18065 -505 18095 -475
rect 18065 -525 18070 -505
rect 18090 -525 18095 -505
rect 18065 -535 18095 -525
rect 18125 -455 18155 -445
rect 18125 -475 18130 -455
rect 18150 -475 18155 -455
rect 18125 -505 18155 -475
rect 18125 -525 18130 -505
rect 18150 -525 18155 -505
rect 18125 -535 18155 -525
rect 18185 -455 18215 -445
rect 18185 -475 18190 -455
rect 18210 -475 18215 -455
rect 18185 -505 18215 -475
rect 18185 -525 18190 -505
rect 18210 -525 18215 -505
rect 18185 -535 18215 -525
rect 18245 -455 18275 -445
rect 18245 -475 18250 -455
rect 18270 -475 18275 -455
rect 18245 -505 18275 -475
rect 18245 -525 18250 -505
rect 18270 -525 18275 -505
rect 18245 -535 18275 -525
rect 18305 -455 18335 -445
rect 18305 -475 18310 -455
rect 18330 -475 18335 -455
rect 18305 -505 18335 -475
rect 18305 -525 18310 -505
rect 18330 -525 18335 -505
rect 18305 -535 18335 -525
rect 18365 -455 18395 -445
rect 18365 -475 18370 -455
rect 18390 -475 18395 -455
rect 18365 -505 18395 -475
rect 18365 -525 18370 -505
rect 18390 -525 18395 -505
rect 18365 -535 18395 -525
rect 18425 -455 18455 -445
rect 18425 -475 18430 -455
rect 18450 -475 18455 -455
rect 18425 -505 18455 -475
rect 18425 -525 18430 -505
rect 18450 -525 18455 -505
rect 18425 -535 18455 -525
rect 18485 -455 18515 -445
rect 18485 -475 18490 -455
rect 18510 -475 18515 -455
rect 18485 -505 18515 -475
rect 18485 -525 18490 -505
rect 18510 -525 18515 -505
rect 18485 -535 18515 -525
rect 18545 -455 18575 -445
rect 18545 -475 18550 -455
rect 18570 -475 18575 -455
rect 18545 -505 18575 -475
rect 18545 -525 18550 -505
rect 18570 -525 18575 -505
rect 18545 -535 18575 -525
rect 18605 -455 18635 -445
rect 18605 -475 18610 -455
rect 18630 -475 18635 -455
rect 18605 -505 18635 -475
rect 18605 -525 18610 -505
rect 18630 -525 18635 -505
rect 18605 -535 18635 -525
rect 18665 -455 18695 -445
rect 18665 -475 18670 -455
rect 18690 -475 18695 -455
rect 18665 -505 18695 -475
rect 18665 -525 18670 -505
rect 18690 -525 18695 -505
rect 18665 -535 18695 -525
rect 18725 -455 18755 -445
rect 18725 -475 18730 -455
rect 18750 -475 18755 -455
rect 18725 -505 18755 -475
rect 18725 -525 18730 -505
rect 18750 -525 18755 -505
rect 18725 -535 18755 -525
rect 18785 -455 18815 -445
rect 18785 -475 18790 -455
rect 18810 -475 18815 -455
rect 18785 -505 18815 -475
rect 18785 -525 18790 -505
rect 18810 -525 18815 -505
rect 18785 -535 18815 -525
rect 18845 -455 18875 -445
rect 18845 -475 18850 -455
rect 18870 -475 18875 -455
rect 18845 -505 18875 -475
rect 18845 -525 18850 -505
rect 18870 -525 18875 -505
rect 18845 -535 18875 -525
rect 18905 -455 18935 -445
rect 18905 -475 18910 -455
rect 18930 -475 18935 -455
rect 18905 -505 18935 -475
rect 18905 -525 18910 -505
rect 18930 -525 18935 -505
rect 18905 -535 18935 -525
rect 18965 -455 18995 -445
rect 18965 -475 18970 -455
rect 18990 -475 18995 -455
rect 18965 -505 18995 -475
rect 18965 -525 18970 -505
rect 18990 -525 18995 -505
rect 18965 -535 18995 -525
rect 19025 -455 19055 -445
rect 19025 -475 19030 -455
rect 19050 -475 19055 -455
rect 19025 -505 19055 -475
rect 19025 -525 19030 -505
rect 19050 -525 19055 -505
rect 19025 -535 19055 -525
rect 19085 -455 19115 -445
rect 19085 -475 19090 -455
rect 19110 -475 19115 -455
rect 19085 -505 19115 -475
rect 19085 -525 19090 -505
rect 19110 -525 19115 -505
rect 19085 -535 19115 -525
rect 19145 -455 19215 -445
rect 19145 -475 19150 -455
rect 19170 -475 19190 -455
rect 19210 -475 19215 -455
rect 19145 -505 19215 -475
rect 19145 -525 19150 -505
rect 19170 -525 19190 -505
rect 19210 -525 19215 -505
rect 19145 -535 19215 -525
rect 16515 -570 16545 -560
rect 16515 -590 16520 -570
rect 16540 -590 16545 -570
rect 16515 -600 16545 -590
rect 16600 -565 16640 -555
rect 16600 -585 16610 -565
rect 16630 -585 16640 -565
rect 16600 -595 16640 -585
rect 16845 -565 16875 -555
rect 16845 -585 16850 -565
rect 16870 -585 16875 -565
rect 16845 -595 16875 -585
rect 16960 -565 17000 -555
rect 16960 -585 16970 -565
rect 16990 -585 17000 -565
rect 16960 -595 17000 -585
rect 17205 -565 17235 -555
rect 17205 -585 17210 -565
rect 17230 -585 17235 -565
rect 17205 -595 17235 -585
rect 17320 -565 17360 -555
rect 17320 -585 17330 -565
rect 17350 -585 17360 -565
rect 17320 -595 17360 -585
rect 17535 -565 17565 -555
rect 17535 -585 17540 -565
rect 17560 -585 17565 -565
rect 17535 -595 17565 -585
rect 18035 -565 18065 -555
rect 18035 -585 18040 -565
rect 18060 -585 18065 -565
rect 18035 -595 18065 -585
rect 18240 -565 18280 -555
rect 18240 -585 18250 -565
rect 18270 -585 18280 -565
rect 18240 -595 18280 -585
rect 18365 -565 18395 -555
rect 18365 -585 18370 -565
rect 18390 -585 18395 -565
rect 18365 -595 18395 -585
rect 18600 -565 18640 -555
rect 18600 -585 18610 -565
rect 18630 -585 18640 -565
rect 18600 -595 18640 -585
rect 18725 -565 18755 -555
rect 18725 -585 18730 -565
rect 18750 -585 18755 -565
rect 18725 -595 18755 -585
rect 18960 -565 19000 -555
rect 18960 -585 18970 -565
rect 18990 -585 19000 -565
rect 18960 -595 19000 -585
rect 19055 -570 19085 -560
rect 19055 -590 19060 -570
rect 19080 -590 19085 -570
rect 19055 -600 19085 -590
rect 17007 -760 17037 -750
rect 17007 -780 17012 -760
rect 17032 -780 17037 -760
rect 17007 -790 17037 -780
rect 18563 -760 18593 -750
rect 18563 -780 18568 -760
rect 18588 -780 18593 -760
rect 18563 -790 18593 -780
rect 16965 -820 16995 -810
rect 16965 -840 16970 -820
rect 16990 -840 16995 -820
rect 16965 -870 16995 -840
rect 16965 -890 16970 -870
rect 16990 -890 16995 -870
rect 16965 -920 16995 -890
rect 16965 -940 16970 -920
rect 16990 -940 16995 -920
rect 16965 -970 16995 -940
rect 16965 -990 16970 -970
rect 16990 -990 16995 -970
rect 16965 -1020 16995 -990
rect 16965 -1040 16970 -1020
rect 16990 -1040 16995 -1020
rect 16965 -1050 16995 -1040
rect 17025 -820 17055 -810
rect 17025 -840 17030 -820
rect 17050 -840 17055 -820
rect 17025 -870 17055 -840
rect 17025 -890 17030 -870
rect 17050 -890 17055 -870
rect 17025 -920 17055 -890
rect 17025 -940 17030 -920
rect 17050 -940 17055 -920
rect 17025 -970 17055 -940
rect 17025 -990 17030 -970
rect 17050 -990 17055 -970
rect 17025 -1020 17055 -990
rect 17025 -1040 17030 -1020
rect 17050 -1040 17055 -1020
rect 17025 -1050 17055 -1040
rect 17085 -820 17115 -810
rect 17085 -840 17090 -820
rect 17110 -840 17115 -820
rect 17085 -870 17115 -840
rect 17085 -890 17090 -870
rect 17110 -890 17115 -870
rect 17085 -920 17115 -890
rect 17085 -940 17090 -920
rect 17110 -940 17115 -920
rect 17560 -820 17600 -810
rect 17560 -840 17570 -820
rect 17590 -840 17600 -820
rect 17560 -860 17600 -840
rect 17560 -880 17570 -860
rect 17590 -880 17600 -860
rect 17560 -900 17600 -880
rect 17560 -920 17570 -900
rect 17590 -920 17600 -900
rect 17560 -930 17600 -920
rect 18000 -820 18040 -810
rect 18000 -840 18010 -820
rect 18030 -840 18040 -820
rect 18000 -860 18040 -840
rect 18000 -880 18010 -860
rect 18030 -880 18040 -860
rect 18000 -900 18040 -880
rect 18000 -920 18010 -900
rect 18030 -920 18040 -900
rect 18000 -930 18040 -920
rect 18485 -820 18515 -810
rect 18485 -840 18490 -820
rect 18510 -840 18515 -820
rect 18485 -870 18515 -840
rect 18485 -890 18490 -870
rect 18510 -890 18515 -870
rect 18485 -920 18515 -890
rect 17085 -970 17115 -940
rect 17085 -990 17090 -970
rect 17110 -990 17115 -970
rect 17085 -1020 17115 -990
rect 17085 -1040 17090 -1020
rect 17110 -1040 17115 -1020
rect 17085 -1050 17115 -1040
rect 18485 -940 18490 -920
rect 18510 -940 18515 -920
rect 18485 -970 18515 -940
rect 18485 -990 18490 -970
rect 18510 -990 18515 -970
rect 18485 -1020 18515 -990
rect 18485 -1040 18490 -1020
rect 18510 -1040 18515 -1020
rect 18485 -1050 18515 -1040
rect 18545 -820 18575 -810
rect 18545 -840 18550 -820
rect 18570 -840 18575 -820
rect 18545 -870 18575 -840
rect 18545 -890 18550 -870
rect 18570 -890 18575 -870
rect 18545 -920 18575 -890
rect 18545 -940 18550 -920
rect 18570 -940 18575 -920
rect 18545 -970 18575 -940
rect 18545 -990 18550 -970
rect 18570 -990 18575 -970
rect 18545 -1020 18575 -990
rect 18545 -1040 18550 -1020
rect 18570 -1040 18575 -1020
rect 18545 -1050 18575 -1040
rect 18605 -820 18635 -810
rect 18605 -840 18610 -820
rect 18630 -840 18635 -820
rect 18605 -870 18635 -840
rect 18605 -890 18610 -870
rect 18630 -890 18635 -870
rect 18605 -920 18635 -890
rect 18605 -940 18610 -920
rect 18630 -940 18635 -920
rect 18605 -970 18635 -940
rect 18605 -990 18610 -970
rect 18630 -990 18635 -970
rect 18605 -1020 18635 -990
rect 18605 -1040 18610 -1020
rect 18630 -1040 18635 -1020
rect 18605 -1050 18635 -1040
rect 17075 -1080 17105 -1070
rect 17075 -1100 17080 -1080
rect 17100 -1100 17105 -1080
rect 17075 -1110 17105 -1100
rect 18440 -1080 18470 -1070
rect 18440 -1100 18445 -1080
rect 18465 -1100 18470 -1080
rect 18440 -1110 18470 -1100
rect 16620 -1270 16660 -1260
rect 16620 -1290 16630 -1270
rect 16650 -1290 16660 -1270
rect 16620 -1300 16660 -1290
rect 16740 -1270 16780 -1260
rect 16740 -1290 16750 -1270
rect 16770 -1290 16780 -1270
rect 16740 -1300 16780 -1290
rect 16860 -1270 16900 -1260
rect 16860 -1290 16870 -1270
rect 16890 -1290 16900 -1270
rect 16860 -1300 16900 -1290
rect 16980 -1270 17020 -1260
rect 16980 -1290 16990 -1270
rect 17010 -1290 17020 -1270
rect 16980 -1300 17020 -1290
rect 17300 -1270 17340 -1260
rect 17300 -1290 17310 -1270
rect 17330 -1290 17340 -1270
rect 17300 -1300 17340 -1290
rect 17420 -1270 17460 -1260
rect 17420 -1290 17430 -1270
rect 17450 -1290 17460 -1270
rect 17420 -1300 17460 -1290
rect 17540 -1270 17580 -1260
rect 17540 -1290 17550 -1270
rect 17570 -1290 17580 -1270
rect 18020 -1270 18060 -1260
rect 17540 -1300 17580 -1290
rect 17695 -1285 17725 -1275
rect 17695 -1305 17700 -1285
rect 17720 -1305 17725 -1285
rect 16535 -1330 16565 -1320
rect 16535 -1350 16540 -1330
rect 16560 -1350 16565 -1330
rect 16535 -1380 16565 -1350
rect 16535 -1400 16540 -1380
rect 16560 -1400 16565 -1380
rect 16535 -1430 16565 -1400
rect 16535 -1450 16540 -1430
rect 16560 -1450 16565 -1430
rect 16535 -1480 16565 -1450
rect 16535 -1500 16540 -1480
rect 16560 -1500 16565 -1480
rect 16535 -1530 16565 -1500
rect 16535 -1550 16540 -1530
rect 16560 -1550 16565 -1530
rect 16535 -1560 16565 -1550
rect 17075 -1330 17185 -1320
rect 17075 -1350 17080 -1330
rect 17100 -1350 17120 -1330
rect 17140 -1350 17160 -1330
rect 17180 -1350 17185 -1330
rect 17075 -1380 17185 -1350
rect 17075 -1400 17080 -1380
rect 17100 -1400 17120 -1380
rect 17140 -1400 17160 -1380
rect 17180 -1400 17185 -1380
rect 17075 -1430 17185 -1400
rect 17075 -1450 17080 -1430
rect 17100 -1450 17120 -1430
rect 17140 -1450 17160 -1430
rect 17180 -1450 17185 -1430
rect 17075 -1480 17185 -1450
rect 17075 -1500 17080 -1480
rect 17100 -1500 17120 -1480
rect 17140 -1500 17160 -1480
rect 17180 -1500 17185 -1480
rect 17075 -1530 17185 -1500
rect 17075 -1550 17080 -1530
rect 17100 -1550 17120 -1530
rect 17140 -1550 17160 -1530
rect 17180 -1550 17185 -1530
rect 17075 -1560 17185 -1550
rect 17695 -1330 17725 -1305
rect 17695 -1350 17700 -1330
rect 17720 -1350 17725 -1330
rect 17695 -1380 17725 -1350
rect 17695 -1400 17700 -1380
rect 17720 -1400 17725 -1380
rect 17695 -1430 17725 -1400
rect 17695 -1450 17700 -1430
rect 17720 -1450 17725 -1430
rect 17695 -1480 17725 -1450
rect 17695 -1500 17700 -1480
rect 17720 -1500 17725 -1480
rect 17695 -1530 17725 -1500
rect 17695 -1550 17700 -1530
rect 17720 -1550 17725 -1530
rect 17695 -1560 17725 -1550
rect 17875 -1285 17905 -1275
rect 17875 -1305 17880 -1285
rect 17900 -1305 17905 -1285
rect 18020 -1290 18030 -1270
rect 18050 -1290 18060 -1270
rect 18020 -1300 18060 -1290
rect 18140 -1270 18180 -1260
rect 18140 -1290 18150 -1270
rect 18170 -1290 18180 -1270
rect 18140 -1300 18180 -1290
rect 18260 -1270 18300 -1260
rect 18260 -1290 18270 -1270
rect 18290 -1290 18300 -1270
rect 18260 -1300 18300 -1290
rect 18580 -1270 18620 -1260
rect 18580 -1290 18590 -1270
rect 18610 -1290 18620 -1270
rect 18580 -1300 18620 -1290
rect 18700 -1270 18740 -1260
rect 18700 -1290 18710 -1270
rect 18730 -1290 18740 -1270
rect 18700 -1300 18740 -1290
rect 18820 -1270 18860 -1260
rect 18820 -1290 18830 -1270
rect 18850 -1290 18860 -1270
rect 18820 -1300 18860 -1290
rect 18940 -1270 18980 -1260
rect 18940 -1290 18950 -1270
rect 18970 -1290 18980 -1270
rect 18940 -1300 18980 -1290
rect 19030 -1290 19070 -1280
rect 17875 -1330 17905 -1305
rect 19030 -1310 19040 -1290
rect 19060 -1310 19070 -1290
rect 19030 -1320 19070 -1310
rect 17875 -1350 17880 -1330
rect 17900 -1350 17905 -1330
rect 17875 -1380 17905 -1350
rect 17875 -1400 17880 -1380
rect 17900 -1400 17905 -1380
rect 17875 -1430 17905 -1400
rect 17875 -1450 17880 -1430
rect 17900 -1450 17905 -1430
rect 17875 -1480 17905 -1450
rect 17875 -1500 17880 -1480
rect 17900 -1500 17905 -1480
rect 17875 -1530 17905 -1500
rect 17875 -1550 17880 -1530
rect 17900 -1550 17905 -1530
rect 17875 -1560 17905 -1550
rect 18415 -1330 18525 -1320
rect 18415 -1350 18420 -1330
rect 18440 -1350 18460 -1330
rect 18480 -1350 18500 -1330
rect 18520 -1350 18525 -1330
rect 18415 -1380 18525 -1350
rect 18415 -1400 18420 -1380
rect 18440 -1400 18460 -1380
rect 18480 -1400 18500 -1380
rect 18520 -1400 18525 -1380
rect 18415 -1430 18525 -1400
rect 18415 -1450 18420 -1430
rect 18440 -1450 18460 -1430
rect 18480 -1450 18500 -1430
rect 18520 -1450 18525 -1430
rect 18415 -1480 18525 -1450
rect 18415 -1500 18420 -1480
rect 18440 -1500 18460 -1480
rect 18480 -1500 18500 -1480
rect 18520 -1500 18525 -1480
rect 18415 -1530 18525 -1500
rect 18415 -1550 18420 -1530
rect 18440 -1550 18460 -1530
rect 18480 -1550 18500 -1530
rect 18520 -1550 18525 -1530
rect 18415 -1560 18525 -1550
rect 19035 -1330 19065 -1320
rect 19035 -1350 19040 -1330
rect 19060 -1350 19065 -1330
rect 19035 -1380 19065 -1350
rect 19035 -1400 19040 -1380
rect 19060 -1400 19065 -1380
rect 19035 -1430 19065 -1400
rect 19035 -1450 19040 -1430
rect 19060 -1450 19065 -1430
rect 19035 -1480 19065 -1450
rect 19035 -1500 19040 -1480
rect 19060 -1500 19065 -1480
rect 19035 -1530 19065 -1500
rect 19035 -1550 19040 -1530
rect 19060 -1550 19065 -1530
rect 19035 -1560 19065 -1550
rect 17120 -1580 17140 -1560
rect 18460 -1580 18480 -1560
rect 17110 -1590 17150 -1580
rect 17110 -1610 17120 -1590
rect 17140 -1610 17150 -1590
rect 17110 -1620 17150 -1610
rect 18450 -1590 18490 -1580
rect 18450 -1610 18460 -1590
rect 18480 -1610 18490 -1590
rect 18450 -1620 18490 -1610
rect 16740 -1725 16780 -1715
rect 16740 -1745 16750 -1725
rect 16770 -1745 16780 -1725
rect 16740 -1755 16780 -1745
rect 16820 -1725 16860 -1715
rect 16820 -1745 16830 -1725
rect 16850 -1745 16860 -1725
rect 16820 -1755 16860 -1745
rect 16900 -1725 16940 -1715
rect 16900 -1745 16910 -1725
rect 16930 -1745 16940 -1725
rect 16900 -1755 16940 -1745
rect 16980 -1725 17020 -1715
rect 16980 -1745 16990 -1725
rect 17010 -1745 17020 -1725
rect 16980 -1755 17020 -1745
rect 17060 -1725 17100 -1715
rect 17060 -1745 17070 -1725
rect 17090 -1745 17100 -1725
rect 17060 -1755 17100 -1745
rect 17140 -1725 17180 -1715
rect 17140 -1745 17150 -1725
rect 17170 -1745 17180 -1725
rect 17140 -1755 17180 -1745
rect 17220 -1725 17260 -1715
rect 17220 -1745 17230 -1725
rect 17250 -1745 17260 -1725
rect 17220 -1755 17260 -1745
rect 17300 -1725 17340 -1715
rect 17300 -1745 17310 -1725
rect 17330 -1745 17340 -1725
rect 17300 -1755 17340 -1745
rect 17380 -1725 17420 -1715
rect 17380 -1745 17390 -1725
rect 17410 -1745 17420 -1725
rect 17380 -1755 17420 -1745
rect 17460 -1725 17500 -1715
rect 17460 -1745 17470 -1725
rect 17490 -1745 17500 -1725
rect 17460 -1755 17500 -1745
rect 17540 -1725 17580 -1715
rect 17540 -1745 17550 -1725
rect 17570 -1745 17580 -1725
rect 17540 -1755 17580 -1745
rect 17620 -1725 17660 -1715
rect 17620 -1745 17630 -1725
rect 17650 -1745 17660 -1725
rect 17620 -1755 17660 -1745
rect 17700 -1725 17740 -1715
rect 17700 -1745 17710 -1725
rect 17730 -1745 17740 -1725
rect 17700 -1755 17740 -1745
rect 17780 -1725 17820 -1715
rect 17780 -1745 17790 -1725
rect 17810 -1745 17820 -1725
rect 17780 -1755 17820 -1745
rect 17860 -1725 17900 -1715
rect 17860 -1745 17870 -1725
rect 17890 -1745 17900 -1725
rect 17860 -1755 17900 -1745
rect 17940 -1725 17980 -1715
rect 17940 -1745 17950 -1725
rect 17970 -1745 17980 -1725
rect 17940 -1755 17980 -1745
rect 18020 -1725 18060 -1715
rect 18020 -1745 18030 -1725
rect 18050 -1745 18060 -1725
rect 18020 -1755 18060 -1745
rect 18100 -1725 18140 -1715
rect 18100 -1745 18110 -1725
rect 18130 -1745 18140 -1725
rect 18100 -1755 18140 -1745
rect 18180 -1725 18220 -1715
rect 18180 -1745 18190 -1725
rect 18210 -1745 18220 -1725
rect 18180 -1755 18220 -1745
rect 18260 -1725 18300 -1715
rect 18260 -1745 18270 -1725
rect 18290 -1745 18300 -1725
rect 18260 -1755 18300 -1745
rect 18340 -1725 18380 -1715
rect 18340 -1745 18350 -1725
rect 18370 -1745 18380 -1725
rect 18340 -1755 18380 -1745
rect 18420 -1725 18460 -1715
rect 18420 -1745 18430 -1725
rect 18450 -1745 18460 -1725
rect 18420 -1755 18460 -1745
rect 18500 -1725 18540 -1715
rect 18500 -1745 18510 -1725
rect 18530 -1745 18540 -1725
rect 18500 -1755 18540 -1745
rect 18580 -1725 18620 -1715
rect 18580 -1745 18590 -1725
rect 18610 -1745 18620 -1725
rect 18580 -1755 18620 -1745
rect 18660 -1725 18700 -1715
rect 18660 -1745 18670 -1725
rect 18690 -1745 18700 -1725
rect 18660 -1755 18700 -1745
rect 18740 -1725 18780 -1715
rect 18740 -1745 18750 -1725
rect 18770 -1745 18780 -1725
rect 18740 -1755 18780 -1745
rect 16750 -1775 16770 -1755
rect 17790 -1775 17810 -1755
rect 16745 -1785 16775 -1775
rect 16745 -1800 16750 -1785
rect 16700 -1805 16750 -1800
rect 16770 -1805 16775 -1785
rect 16700 -1810 16775 -1805
rect 16700 -1830 16710 -1810
rect 16730 -1830 16775 -1810
rect 16700 -1835 16775 -1830
rect 16700 -1840 16750 -1835
rect 16745 -1855 16750 -1840
rect 16770 -1855 16775 -1835
rect 16745 -1865 16775 -1855
rect 17785 -1785 17815 -1775
rect 17785 -1805 17790 -1785
rect 17810 -1805 17815 -1785
rect 17785 -1835 17815 -1805
rect 17785 -1855 17790 -1835
rect 17810 -1855 17815 -1835
rect 17785 -1865 17815 -1855
rect 18825 -1780 18895 -1775
rect 18825 -1785 18935 -1780
rect 18825 -1805 18830 -1785
rect 18850 -1805 18870 -1785
rect 18890 -1790 18935 -1785
rect 18890 -1805 18905 -1790
rect 18825 -1810 18905 -1805
rect 18925 -1810 18935 -1790
rect 18825 -1830 18935 -1810
rect 18825 -1835 18905 -1830
rect 18825 -1855 18830 -1835
rect 18850 -1855 18870 -1835
rect 18890 -1850 18905 -1835
rect 18925 -1850 18935 -1830
rect 18890 -1855 18935 -1850
rect 18825 -1860 18935 -1855
rect 18825 -1865 18895 -1860
rect 17425 -2005 17470 -2000
rect 17425 -2030 17435 -2005
rect 17460 -2030 17470 -2005
rect 17425 -2035 17470 -2030
rect 18124 -2005 18169 -2000
rect 18124 -2030 18134 -2005
rect 18159 -2030 18169 -2005
rect 18124 -2035 18169 -2030
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16580 -2975 16605 -2940
rect 16100 -3226 16135 -3215
rect 16100 -3251 16105 -3226
rect 16130 -3251 16135 -3226
rect 16100 -3261 16135 -3251
rect 16210 -3330 16245 -3320
rect 16210 -3355 16215 -3330
rect 16240 -3355 16245 -3330
rect 16210 -3365 16245 -3355
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19305 -3095 19340 -3085
rect 19305 -3120 19310 -3095
rect 19335 -3120 19340 -3095
rect 19305 -3130 19340 -3120
rect 19220 -3165 19245 -3130
rect 19465 -3120 19500 -3110
rect 19465 -3145 19470 -3120
rect 19495 -3145 19500 -3120
rect 19465 -3156 19500 -3145
rect 16795 -3600 18805 -3475
rect 16100 -3899 16135 -3889
rect 16100 -3924 16105 -3899
rect 16130 -3924 16135 -3899
rect 16100 -3934 16135 -3924
rect 16210 -3899 16245 -3889
rect 16210 -3924 16215 -3899
rect 16240 -3924 16245 -3899
rect 16210 -3934 16245 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4165 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19280 -3889 19305 -3854
rect 19465 -3794 19500 -3784
rect 19465 -3819 19470 -3794
rect 19495 -3819 19500 -3794
rect 19465 -3829 19500 -3819
rect 19185 -3899 19220 -3889
rect 19185 -3924 19190 -3899
rect 19215 -3924 19220 -3899
rect 19185 -3934 19220 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4185 17790 -4165
rect 17810 -4185 17820 -4165
rect 17780 -4205 17820 -4185
rect 17780 -4225 17790 -4205
rect 17810 -4225 17820 -4205
rect 17780 -4245 17820 -4225
rect 17780 -4265 17790 -4245
rect 17810 -4265 17820 -4245
rect 17780 -4275 17820 -4265
<< viali >>
rect 16985 665 17005 685
rect 17645 665 17665 685
rect 17935 665 17955 685
rect 18595 665 18615 685
rect 16945 605 16965 625
rect 16985 605 17005 625
rect 16945 555 16965 575
rect 16985 555 17005 575
rect 17040 605 17060 625
rect 17040 555 17060 575
rect 17095 605 17115 625
rect 17095 555 17115 575
rect 17150 605 17170 625
rect 17150 555 17170 575
rect 17205 605 17225 625
rect 17205 555 17225 575
rect 17260 605 17280 625
rect 17260 555 17280 575
rect 17315 605 17335 625
rect 17315 555 17335 575
rect 17370 605 17390 625
rect 17370 555 17390 575
rect 17425 605 17445 625
rect 17425 555 17445 575
rect 17480 605 17500 625
rect 17480 555 17500 575
rect 17535 605 17555 625
rect 17535 555 17555 575
rect 17590 605 17610 625
rect 17590 555 17610 575
rect 17645 605 17665 625
rect 17685 605 17705 625
rect 17645 555 17665 575
rect 17685 555 17705 575
rect 17895 605 17915 625
rect 17935 605 17955 625
rect 17895 555 17915 575
rect 17935 555 17955 575
rect 17990 605 18010 625
rect 17990 555 18010 575
rect 18045 605 18065 625
rect 18045 555 18065 575
rect 18100 605 18120 625
rect 18100 555 18120 575
rect 18155 605 18175 625
rect 18155 555 18175 575
rect 18210 605 18230 625
rect 18210 555 18230 575
rect 18265 605 18285 625
rect 18265 555 18285 575
rect 18320 605 18340 625
rect 18320 555 18340 575
rect 18375 605 18395 625
rect 18375 555 18395 575
rect 18430 605 18450 625
rect 18430 555 18450 575
rect 18485 605 18505 625
rect 18485 555 18505 575
rect 18540 605 18560 625
rect 18540 555 18560 575
rect 18595 605 18615 625
rect 18635 605 18655 625
rect 18595 555 18615 575
rect 18635 555 18655 575
rect 17069 499 17086 516
rect 17124 499 17141 516
rect 17179 499 17196 516
rect 17234 499 17251 516
rect 17289 499 17306 516
rect 17344 499 17361 516
rect 17399 499 17416 516
rect 17454 499 17471 516
rect 17509 499 17526 516
rect 17564 499 17581 516
rect 18019 499 18036 516
rect 18074 499 18091 516
rect 18129 499 18146 516
rect 18184 499 18201 516
rect 18239 499 18256 516
rect 18294 499 18311 516
rect 18349 499 18366 516
rect 18404 499 18421 516
rect 18459 499 18476 516
rect 18514 499 18531 516
rect 16980 365 17000 385
rect 17160 365 17180 385
rect 17340 365 17360 385
rect 17520 365 17540 385
rect 17700 365 17720 385
rect 17880 365 17900 385
rect 18060 365 18080 385
rect 18240 365 18260 385
rect 18420 365 18440 385
rect 18600 365 18620 385
rect 16980 305 17000 325
rect 16445 265 16465 285
rect 16555 265 16575 285
rect 16665 265 16685 285
rect 16980 255 17000 275
rect 16445 205 16465 225
rect 16445 155 16465 175
rect 16500 205 16520 225
rect 16500 155 16520 175
rect 16555 205 16575 225
rect 16555 155 16575 175
rect 16610 205 16630 225
rect 16610 155 16630 175
rect 16665 205 16685 225
rect 16665 155 16685 175
rect 16980 205 17000 225
rect 16980 155 17000 175
rect 16495 95 16515 115
rect 16555 95 16575 115
rect 16615 95 16635 115
rect 16980 105 17000 125
rect 16980 55 17000 75
rect 17070 305 17090 325
rect 17070 255 17090 275
rect 17070 205 17090 225
rect 17070 155 17090 175
rect 17070 105 17090 125
rect 17070 55 17090 75
rect 17160 305 17180 325
rect 17160 255 17180 275
rect 17160 205 17180 225
rect 17160 155 17180 175
rect 17160 105 17180 125
rect 17160 55 17180 75
rect 17250 305 17270 325
rect 17250 255 17270 275
rect 17250 205 17270 225
rect 17250 155 17270 175
rect 17250 105 17270 125
rect 17250 55 17270 75
rect 17340 305 17360 325
rect 17340 255 17360 275
rect 17340 205 17360 225
rect 17340 155 17360 175
rect 17340 105 17360 125
rect 17340 55 17360 75
rect 17430 305 17450 325
rect 17430 255 17450 275
rect 17430 205 17450 225
rect 17430 155 17450 175
rect 17430 105 17450 125
rect 17430 55 17450 75
rect 17520 305 17540 325
rect 17520 255 17540 275
rect 17520 205 17540 225
rect 17520 155 17540 175
rect 17520 105 17540 125
rect 17520 55 17540 75
rect 17610 305 17630 325
rect 17610 255 17630 275
rect 17610 205 17630 225
rect 17610 155 17630 175
rect 17610 105 17630 125
rect 17610 55 17630 75
rect 17700 305 17720 325
rect 17700 255 17720 275
rect 17700 205 17720 225
rect 17700 155 17720 175
rect 17700 105 17720 125
rect 17700 55 17720 75
rect 17790 305 17810 325
rect 17790 255 17810 275
rect 17790 205 17810 225
rect 17790 155 17810 175
rect 17790 105 17810 125
rect 17790 55 17810 75
rect 17880 305 17900 325
rect 17880 255 17900 275
rect 17880 205 17900 225
rect 17880 155 17900 175
rect 17880 105 17900 125
rect 17880 55 17900 75
rect 17970 305 17990 325
rect 17970 255 17990 275
rect 17970 205 17990 225
rect 17970 155 17990 175
rect 17970 105 17990 125
rect 17970 55 17990 75
rect 18060 305 18080 325
rect 18060 255 18080 275
rect 18060 205 18080 225
rect 18060 155 18080 175
rect 18060 105 18080 125
rect 18060 55 18080 75
rect 18150 305 18170 325
rect 18150 255 18170 275
rect 18150 205 18170 225
rect 18150 155 18170 175
rect 18150 105 18170 125
rect 18150 55 18170 75
rect 18240 305 18260 325
rect 18240 255 18260 275
rect 18240 205 18260 225
rect 18240 155 18260 175
rect 18240 105 18260 125
rect 18240 55 18260 75
rect 18330 305 18350 325
rect 18330 255 18350 275
rect 18330 205 18350 225
rect 18330 155 18350 175
rect 18330 105 18350 125
rect 18330 55 18350 75
rect 18420 305 18440 325
rect 18420 255 18440 275
rect 18420 205 18440 225
rect 18420 155 18440 175
rect 18420 105 18440 125
rect 18420 55 18440 75
rect 18510 305 18530 325
rect 18510 255 18530 275
rect 18510 205 18530 225
rect 18510 155 18530 175
rect 18510 105 18530 125
rect 18510 55 18530 75
rect 18600 305 18620 325
rect 18600 255 18620 275
rect 18600 205 18620 225
rect 18600 155 18620 175
rect 18600 105 18620 125
rect 18600 55 18620 75
rect 17115 -5 17135 15
rect 17205 -5 17225 15
rect 17295 -5 17315 15
rect 17385 -5 17405 15
rect 17475 -5 17495 15
rect 17565 -5 17585 15
rect 17655 -5 17675 15
rect 17745 -5 17765 15
rect 17835 -5 17855 15
rect 17925 -5 17945 15
rect 18015 -5 18035 15
rect 18105 -5 18125 15
rect 18195 -5 18215 15
rect 18285 -5 18305 15
rect 18375 -5 18395 15
rect 18465 -5 18485 15
rect 16430 -415 16450 -395
rect 17630 -415 17650 -395
rect 17950 -415 17970 -395
rect 19150 -415 19170 -395
rect 16430 -475 16450 -455
rect 16430 -525 16450 -505
rect 16490 -475 16510 -455
rect 16490 -525 16510 -505
rect 16550 -475 16570 -455
rect 16550 -525 16570 -505
rect 16610 -475 16630 -455
rect 16610 -525 16630 -505
rect 16670 -475 16690 -455
rect 16670 -525 16690 -505
rect 16730 -475 16750 -455
rect 16730 -525 16750 -505
rect 16790 -475 16810 -455
rect 16790 -525 16810 -505
rect 16850 -475 16870 -455
rect 16850 -525 16870 -505
rect 16910 -475 16930 -455
rect 16910 -525 16930 -505
rect 16970 -475 16990 -455
rect 16970 -525 16990 -505
rect 17030 -475 17050 -455
rect 17030 -525 17050 -505
rect 17090 -475 17110 -455
rect 17090 -525 17110 -505
rect 17150 -475 17170 -455
rect 17150 -525 17170 -505
rect 17210 -475 17230 -455
rect 17210 -525 17230 -505
rect 17270 -475 17290 -455
rect 17270 -525 17290 -505
rect 17330 -475 17350 -455
rect 17330 -525 17350 -505
rect 17390 -475 17410 -455
rect 17390 -525 17410 -505
rect 17450 -475 17470 -455
rect 17450 -525 17470 -505
rect 17510 -475 17530 -455
rect 17510 -525 17530 -505
rect 17570 -475 17590 -455
rect 17570 -525 17590 -505
rect 17630 -475 17650 -455
rect 17630 -525 17650 -505
rect 17950 -475 17970 -455
rect 17950 -525 17970 -505
rect 18010 -475 18030 -455
rect 18010 -525 18030 -505
rect 18070 -475 18090 -455
rect 18070 -525 18090 -505
rect 18130 -475 18150 -455
rect 18130 -525 18150 -505
rect 18190 -475 18210 -455
rect 18190 -525 18210 -505
rect 18250 -475 18270 -455
rect 18250 -525 18270 -505
rect 18310 -475 18330 -455
rect 18310 -525 18330 -505
rect 18370 -475 18390 -455
rect 18370 -525 18390 -505
rect 18430 -475 18450 -455
rect 18430 -525 18450 -505
rect 18490 -475 18510 -455
rect 18490 -525 18510 -505
rect 18550 -475 18570 -455
rect 18550 -525 18570 -505
rect 18610 -475 18630 -455
rect 18610 -525 18630 -505
rect 18670 -475 18690 -455
rect 18670 -525 18690 -505
rect 18730 -475 18750 -455
rect 18730 -525 18750 -505
rect 18790 -475 18810 -455
rect 18790 -525 18810 -505
rect 18850 -475 18870 -455
rect 18850 -525 18870 -505
rect 18910 -475 18930 -455
rect 18910 -525 18930 -505
rect 18970 -475 18990 -455
rect 18970 -525 18990 -505
rect 19030 -475 19050 -455
rect 19030 -525 19050 -505
rect 19090 -475 19110 -455
rect 19090 -525 19110 -505
rect 19150 -475 19170 -455
rect 19150 -525 19170 -505
rect 16520 -590 16540 -570
rect 16610 -585 16630 -565
rect 16850 -585 16870 -565
rect 16970 -585 16990 -565
rect 17210 -585 17230 -565
rect 17330 -585 17350 -565
rect 17540 -585 17560 -565
rect 18040 -585 18060 -565
rect 18250 -585 18270 -565
rect 18370 -585 18390 -565
rect 18610 -585 18630 -565
rect 18730 -585 18750 -565
rect 18970 -585 18990 -565
rect 19060 -590 19080 -570
rect 17012 -780 17032 -760
rect 18568 -780 18588 -760
rect 16970 -840 16990 -820
rect 16970 -890 16990 -870
rect 16970 -940 16990 -920
rect 16970 -990 16990 -970
rect 16970 -1040 16990 -1020
rect 17030 -840 17050 -820
rect 17030 -890 17050 -870
rect 17030 -940 17050 -920
rect 17030 -990 17050 -970
rect 17030 -1040 17050 -1020
rect 17090 -840 17110 -820
rect 17090 -890 17110 -870
rect 17090 -940 17110 -920
rect 17570 -840 17590 -820
rect 17570 -880 17590 -860
rect 17570 -920 17590 -900
rect 18010 -840 18030 -820
rect 18010 -880 18030 -860
rect 18010 -920 18030 -900
rect 18490 -840 18510 -820
rect 18490 -890 18510 -870
rect 17090 -990 17110 -970
rect 17090 -1040 17110 -1020
rect 18490 -940 18510 -920
rect 18490 -990 18510 -970
rect 18490 -1040 18510 -1020
rect 18550 -840 18570 -820
rect 18550 -890 18570 -870
rect 18550 -940 18570 -920
rect 18550 -990 18570 -970
rect 18550 -1040 18570 -1020
rect 18610 -840 18630 -820
rect 18610 -890 18630 -870
rect 18610 -940 18630 -920
rect 18610 -990 18630 -970
rect 18610 -1040 18630 -1020
rect 17080 -1100 17100 -1080
rect 18445 -1100 18465 -1080
rect 16630 -1290 16650 -1270
rect 16750 -1290 16770 -1270
rect 16870 -1290 16890 -1270
rect 16990 -1290 17010 -1270
rect 17310 -1290 17330 -1270
rect 17430 -1290 17450 -1270
rect 17550 -1290 17570 -1270
rect 17700 -1305 17720 -1285
rect 16540 -1350 16560 -1330
rect 16540 -1400 16560 -1380
rect 16540 -1450 16560 -1430
rect 16540 -1500 16560 -1480
rect 16540 -1550 16560 -1530
rect 17880 -1305 17900 -1285
rect 18030 -1290 18050 -1270
rect 18150 -1290 18170 -1270
rect 18270 -1290 18290 -1270
rect 18590 -1290 18610 -1270
rect 18710 -1290 18730 -1270
rect 18830 -1290 18850 -1270
rect 18950 -1290 18970 -1270
rect 19040 -1310 19060 -1290
rect 17120 -1610 17140 -1590
rect 18460 -1610 18480 -1590
rect 16750 -1745 16770 -1725
rect 16830 -1745 16850 -1725
rect 16910 -1745 16930 -1725
rect 16990 -1745 17010 -1725
rect 17070 -1745 17090 -1725
rect 17150 -1745 17170 -1725
rect 17230 -1745 17250 -1725
rect 17310 -1745 17330 -1725
rect 17390 -1745 17410 -1725
rect 17470 -1745 17490 -1725
rect 17550 -1745 17570 -1725
rect 17630 -1745 17650 -1725
rect 17710 -1745 17730 -1725
rect 17790 -1745 17810 -1725
rect 17870 -1745 17890 -1725
rect 17950 -1745 17970 -1725
rect 18030 -1745 18050 -1725
rect 18110 -1745 18130 -1725
rect 18190 -1745 18210 -1725
rect 18270 -1745 18290 -1725
rect 18350 -1745 18370 -1725
rect 18430 -1745 18450 -1725
rect 18510 -1745 18530 -1725
rect 18590 -1745 18610 -1725
rect 18670 -1745 18690 -1725
rect 18750 -1745 18770 -1725
rect 16710 -1830 16730 -1810
rect 18905 -1810 18925 -1790
rect 18905 -1850 18925 -1830
rect 17435 -2030 17460 -2005
rect 18134 -2030 18159 -2005
rect 16490 -2930 16515 -2905
rect 16105 -3251 16130 -3226
rect 16215 -3355 16240 -3330
rect 19085 -2930 19110 -2905
rect 19310 -3120 19335 -3095
rect 19470 -3145 19495 -3120
rect 16105 -3924 16130 -3899
rect 16215 -3924 16240 -3899
rect 16610 -3999 16635 -3974
rect 19470 -3819 19495 -3794
rect 19190 -3924 19215 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4185 17810 -4165
rect 17790 -4225 17810 -4205
rect 17790 -4265 17810 -4245
<< metal1 >>
rect 17030 745 17070 980
rect 17030 715 17035 745
rect 17065 715 17070 745
rect 17030 710 17070 715
rect 17140 745 17180 980
rect 17140 715 17145 745
rect 17175 715 17180 745
rect 17140 710 17180 715
rect 17250 745 17290 980
rect 17250 715 17255 745
rect 17285 715 17290 745
rect 17250 710 17290 715
rect 17360 745 17400 980
rect 17360 715 17365 745
rect 17395 715 17400 745
rect 17360 710 17400 715
rect 17470 745 17510 980
rect 17470 715 17475 745
rect 17505 715 17510 745
rect 17470 710 17510 715
rect 17580 745 17620 980
rect 17580 715 17585 745
rect 17615 715 17620 745
rect 17580 710 17620 715
rect 17980 745 18020 750
rect 17980 715 17985 745
rect 18015 715 18020 745
rect 17980 710 18020 715
rect 18090 745 18130 750
rect 18090 715 18095 745
rect 18125 715 18130 745
rect 18090 710 18130 715
rect 18200 745 18240 750
rect 18200 715 18205 745
rect 18235 715 18240 745
rect 18200 710 18240 715
rect 18310 745 18350 750
rect 18310 715 18315 745
rect 18345 715 18350 745
rect 18310 710 18350 715
rect 18420 745 18460 750
rect 18420 715 18425 745
rect 18455 715 18460 745
rect 18420 710 18460 715
rect 18530 745 18570 750
rect 18530 715 18535 745
rect 18565 715 18570 745
rect 18530 710 18570 715
rect 19225 745 19265 750
rect 19225 715 19230 745
rect 19260 715 19265 745
rect 16975 690 17015 695
rect 16975 660 16980 690
rect 17010 660 17015 690
rect 16975 655 17015 660
rect 16980 635 17010 655
rect 16940 625 17010 635
rect 16940 605 16945 625
rect 16965 605 16985 625
rect 17005 605 17010 625
rect 16940 575 17010 605
rect 16940 555 16945 575
rect 16965 555 16985 575
rect 17005 555 17010 575
rect 16940 545 17010 555
rect 17035 625 17065 710
rect 17085 690 17125 695
rect 17085 660 17090 690
rect 17120 660 17125 690
rect 17085 655 17125 660
rect 17035 605 17040 625
rect 17060 605 17065 625
rect 17035 575 17065 605
rect 17035 555 17040 575
rect 17060 555 17065 575
rect 17035 545 17065 555
rect 17090 625 17120 655
rect 17090 605 17095 625
rect 17115 605 17120 625
rect 17090 575 17120 605
rect 17090 555 17095 575
rect 17115 555 17120 575
rect 17090 545 17120 555
rect 17145 625 17175 710
rect 17195 690 17235 695
rect 17195 660 17200 690
rect 17230 660 17235 690
rect 17195 655 17235 660
rect 17145 605 17150 625
rect 17170 605 17175 625
rect 17145 575 17175 605
rect 17145 555 17150 575
rect 17170 555 17175 575
rect 17145 545 17175 555
rect 17200 625 17230 655
rect 17200 605 17205 625
rect 17225 605 17230 625
rect 17200 575 17230 605
rect 17200 555 17205 575
rect 17225 555 17230 575
rect 17200 545 17230 555
rect 17255 625 17285 710
rect 17305 690 17345 695
rect 17305 660 17310 690
rect 17340 660 17345 690
rect 17305 655 17345 660
rect 17255 605 17260 625
rect 17280 605 17285 625
rect 17255 575 17285 605
rect 17255 555 17260 575
rect 17280 555 17285 575
rect 17255 545 17285 555
rect 17310 625 17340 655
rect 17310 605 17315 625
rect 17335 605 17340 625
rect 17310 575 17340 605
rect 17310 555 17315 575
rect 17335 555 17340 575
rect 17310 545 17340 555
rect 17365 625 17395 710
rect 17415 690 17455 695
rect 17415 660 17420 690
rect 17450 660 17455 690
rect 17415 655 17455 660
rect 17365 605 17370 625
rect 17390 605 17395 625
rect 17365 575 17395 605
rect 17365 555 17370 575
rect 17390 555 17395 575
rect 17365 545 17395 555
rect 17420 625 17450 655
rect 17420 605 17425 625
rect 17445 605 17450 625
rect 17420 575 17450 605
rect 17420 555 17425 575
rect 17445 555 17450 575
rect 17420 545 17450 555
rect 17475 625 17505 710
rect 17525 690 17565 695
rect 17525 660 17530 690
rect 17560 660 17565 690
rect 17525 655 17565 660
rect 17475 605 17480 625
rect 17500 605 17505 625
rect 17475 575 17505 605
rect 17475 555 17480 575
rect 17500 555 17505 575
rect 17475 545 17505 555
rect 17530 625 17560 655
rect 17530 605 17535 625
rect 17555 605 17560 625
rect 17530 575 17560 605
rect 17530 555 17535 575
rect 17555 555 17560 575
rect 17530 545 17560 555
rect 17585 625 17615 710
rect 17635 690 17675 695
rect 17635 660 17640 690
rect 17670 660 17675 690
rect 17635 655 17675 660
rect 17925 690 17965 695
rect 17925 660 17930 690
rect 17960 660 17965 690
rect 17925 655 17965 660
rect 17585 605 17590 625
rect 17610 605 17615 625
rect 17585 575 17615 605
rect 17585 555 17590 575
rect 17610 555 17615 575
rect 17585 545 17615 555
rect 17640 635 17670 655
rect 17930 635 17960 655
rect 17640 625 17710 635
rect 17640 605 17645 625
rect 17665 605 17685 625
rect 17705 605 17710 625
rect 17640 575 17710 605
rect 17640 555 17645 575
rect 17665 555 17685 575
rect 17705 555 17710 575
rect 17640 545 17710 555
rect 17890 625 17960 635
rect 17890 605 17895 625
rect 17915 605 17935 625
rect 17955 605 17960 625
rect 17890 575 17960 605
rect 17890 555 17895 575
rect 17915 555 17935 575
rect 17955 555 17960 575
rect 17890 545 17960 555
rect 17985 625 18015 710
rect 18035 690 18075 695
rect 18035 660 18040 690
rect 18070 660 18075 690
rect 18035 655 18075 660
rect 17985 605 17990 625
rect 18010 605 18015 625
rect 17985 575 18015 605
rect 17985 555 17990 575
rect 18010 555 18015 575
rect 17985 545 18015 555
rect 18040 625 18070 655
rect 18040 605 18045 625
rect 18065 605 18070 625
rect 18040 575 18070 605
rect 18040 555 18045 575
rect 18065 555 18070 575
rect 18040 545 18070 555
rect 18095 625 18125 710
rect 18145 690 18185 695
rect 18145 660 18150 690
rect 18180 660 18185 690
rect 18145 655 18185 660
rect 18095 605 18100 625
rect 18120 605 18125 625
rect 18095 575 18125 605
rect 18095 555 18100 575
rect 18120 555 18125 575
rect 18095 545 18125 555
rect 18150 625 18180 655
rect 18150 605 18155 625
rect 18175 605 18180 625
rect 18150 575 18180 605
rect 18150 555 18155 575
rect 18175 555 18180 575
rect 18150 545 18180 555
rect 18205 625 18235 710
rect 18255 690 18295 695
rect 18255 660 18260 690
rect 18290 660 18295 690
rect 18255 655 18295 660
rect 18205 605 18210 625
rect 18230 605 18235 625
rect 18205 575 18235 605
rect 18205 555 18210 575
rect 18230 555 18235 575
rect 18205 545 18235 555
rect 18260 625 18290 655
rect 18260 605 18265 625
rect 18285 605 18290 625
rect 18260 575 18290 605
rect 18260 555 18265 575
rect 18285 555 18290 575
rect 18260 545 18290 555
rect 18315 625 18345 710
rect 18365 690 18405 695
rect 18365 660 18370 690
rect 18400 660 18405 690
rect 18365 655 18405 660
rect 18315 605 18320 625
rect 18340 605 18345 625
rect 18315 575 18345 605
rect 18315 555 18320 575
rect 18340 555 18345 575
rect 18315 545 18345 555
rect 18370 625 18400 655
rect 18370 605 18375 625
rect 18395 605 18400 625
rect 18370 575 18400 605
rect 18370 555 18375 575
rect 18395 555 18400 575
rect 18370 545 18400 555
rect 18425 625 18455 710
rect 18475 690 18515 695
rect 18475 660 18480 690
rect 18510 660 18515 690
rect 18475 655 18515 660
rect 18425 605 18430 625
rect 18450 605 18455 625
rect 18425 575 18455 605
rect 18425 555 18430 575
rect 18450 555 18455 575
rect 18425 545 18455 555
rect 18480 625 18510 655
rect 18480 605 18485 625
rect 18505 605 18510 625
rect 18480 575 18510 605
rect 18480 555 18485 575
rect 18505 555 18510 575
rect 18480 545 18510 555
rect 18535 625 18565 710
rect 18585 690 18625 695
rect 18585 660 18590 690
rect 18620 660 18625 690
rect 18585 655 18625 660
rect 18535 605 18540 625
rect 18560 605 18565 625
rect 18535 575 18565 605
rect 18535 555 18540 575
rect 18560 555 18565 575
rect 18535 545 18565 555
rect 18590 635 18620 655
rect 18590 625 18660 635
rect 18590 605 18595 625
rect 18615 605 18635 625
rect 18655 605 18660 625
rect 18590 575 18660 605
rect 18590 555 18595 575
rect 18615 555 18635 575
rect 18655 555 18660 575
rect 18590 545 18660 555
rect 17063 521 17092 525
rect 17063 495 17065 521
rect 17091 495 17092 521
rect 17063 490 17092 495
rect 17118 521 17147 525
rect 17118 495 17120 521
rect 17146 495 17147 521
rect 17118 490 17147 495
rect 17173 521 17202 525
rect 17173 495 17175 521
rect 17201 495 17202 521
rect 17173 490 17202 495
rect 17228 521 17257 525
rect 17228 495 17230 521
rect 17256 495 17257 521
rect 17228 490 17257 495
rect 17283 521 17312 525
rect 17283 495 17285 521
rect 17311 495 17312 521
rect 17283 490 17312 495
rect 17338 521 17367 525
rect 17338 495 17340 521
rect 17366 495 17367 521
rect 17338 490 17367 495
rect 17393 521 17422 525
rect 17393 495 17395 521
rect 17421 495 17422 521
rect 17393 490 17422 495
rect 17448 521 17477 525
rect 17448 495 17450 521
rect 17476 495 17477 521
rect 17448 490 17477 495
rect 17503 521 17532 525
rect 17503 495 17505 521
rect 17531 495 17532 521
rect 17503 490 17532 495
rect 17558 521 17587 525
rect 17558 495 17560 521
rect 17586 495 17587 521
rect 17558 490 17587 495
rect 18013 521 18042 525
rect 18013 495 18015 521
rect 18041 495 18042 521
rect 18013 490 18042 495
rect 18068 521 18097 525
rect 18068 495 18070 521
rect 18096 495 18097 521
rect 18068 490 18097 495
rect 18123 521 18152 525
rect 18123 495 18125 521
rect 18151 495 18152 521
rect 18123 490 18152 495
rect 18178 521 18207 525
rect 18178 495 18180 521
rect 18206 495 18207 521
rect 18178 490 18207 495
rect 18233 521 18262 525
rect 18233 495 18235 521
rect 18261 495 18262 521
rect 18233 490 18262 495
rect 18288 521 18317 525
rect 18288 495 18290 521
rect 18316 495 18317 521
rect 18288 490 18317 495
rect 18343 521 18372 525
rect 18343 495 18345 521
rect 18371 495 18372 521
rect 18343 490 18372 495
rect 18398 521 18427 525
rect 18398 495 18400 521
rect 18426 495 18427 521
rect 18398 490 18427 495
rect 18453 521 18482 525
rect 18453 495 18455 521
rect 18481 495 18482 521
rect 18453 490 18482 495
rect 18508 521 18537 525
rect 18508 495 18510 521
rect 18536 495 18537 521
rect 18508 490 18537 495
rect 16435 470 16475 475
rect 16435 440 16440 470
rect 16470 440 16475 470
rect 16435 430 16475 440
rect 16435 400 16440 430
rect 16470 400 16475 430
rect 16435 390 16475 400
rect 16435 360 16440 390
rect 16470 360 16475 390
rect 16435 355 16475 360
rect 16655 470 16695 475
rect 16655 440 16660 470
rect 16690 440 16695 470
rect 16655 430 16695 440
rect 16655 400 16660 430
rect 16690 400 16695 430
rect 16655 390 16695 400
rect 16655 360 16660 390
rect 16690 360 16695 390
rect 16655 355 16695 360
rect 16970 470 17010 475
rect 16970 440 16975 470
rect 17005 440 17010 470
rect 16970 430 17010 440
rect 16970 400 16975 430
rect 17005 400 17010 430
rect 16970 390 17010 400
rect 16970 360 16975 390
rect 17005 360 17010 390
rect 16970 355 17010 360
rect 17150 470 17190 475
rect 17150 440 17155 470
rect 17185 440 17190 470
rect 17150 430 17190 440
rect 17150 400 17155 430
rect 17185 400 17190 430
rect 17150 390 17190 400
rect 17150 360 17155 390
rect 17185 360 17190 390
rect 17150 355 17190 360
rect 17330 470 17370 475
rect 17330 440 17335 470
rect 17365 440 17370 470
rect 17330 430 17370 440
rect 17330 400 17335 430
rect 17365 400 17370 430
rect 17330 390 17370 400
rect 17330 360 17335 390
rect 17365 360 17370 390
rect 17330 355 17370 360
rect 17510 470 17550 475
rect 17510 440 17515 470
rect 17545 440 17550 470
rect 17510 430 17550 440
rect 17510 400 17515 430
rect 17545 400 17550 430
rect 17510 390 17550 400
rect 17510 360 17515 390
rect 17545 360 17550 390
rect 17510 355 17550 360
rect 17690 470 17730 475
rect 17690 440 17695 470
rect 17725 440 17730 470
rect 17690 430 17730 440
rect 17690 400 17695 430
rect 17725 400 17730 430
rect 17690 390 17730 400
rect 17690 360 17695 390
rect 17725 360 17730 390
rect 17690 355 17730 360
rect 17870 470 17910 475
rect 17870 440 17875 470
rect 17905 440 17910 470
rect 17870 430 17910 440
rect 17870 400 17875 430
rect 17905 400 17910 430
rect 17870 390 17910 400
rect 17870 360 17875 390
rect 17905 360 17910 390
rect 17870 355 17910 360
rect 18050 470 18090 475
rect 18050 440 18055 470
rect 18085 440 18090 470
rect 18050 430 18090 440
rect 18050 400 18055 430
rect 18085 400 18090 430
rect 18050 390 18090 400
rect 18050 360 18055 390
rect 18085 360 18090 390
rect 18050 355 18090 360
rect 18230 470 18270 475
rect 18230 440 18235 470
rect 18265 440 18270 470
rect 18230 430 18270 440
rect 18230 400 18235 430
rect 18265 400 18270 430
rect 18230 390 18270 400
rect 18230 360 18235 390
rect 18265 360 18270 390
rect 18230 355 18270 360
rect 18410 470 18450 475
rect 18410 440 18415 470
rect 18445 440 18450 470
rect 18410 430 18450 440
rect 18410 400 18415 430
rect 18445 400 18450 430
rect 18410 390 18450 400
rect 18410 360 18415 390
rect 18445 360 18450 390
rect 18410 355 18450 360
rect 18590 470 18630 475
rect 18590 440 18595 470
rect 18625 440 18630 470
rect 18590 430 18630 440
rect 18590 400 18595 430
rect 18625 400 18630 430
rect 18590 390 18630 400
rect 18590 360 18595 390
rect 18625 360 18630 390
rect 18590 355 18630 360
rect 16440 295 16470 355
rect 16660 295 16690 355
rect 16975 325 17005 335
rect 16975 305 16980 325
rect 17000 305 17005 325
rect 16435 285 16475 295
rect 16435 265 16445 285
rect 16465 265 16475 285
rect 16435 255 16475 265
rect 16545 290 16585 295
rect 16545 260 16550 290
rect 16580 260 16585 290
rect 16545 255 16585 260
rect 16655 285 16695 295
rect 16655 265 16665 285
rect 16685 265 16695 285
rect 16655 255 16695 265
rect 16780 290 16820 295
rect 16780 260 16785 290
rect 16815 260 16820 290
rect 16780 255 16820 260
rect 16975 275 17005 305
rect 16975 255 16980 275
rect 17000 255 17005 275
rect 16440 225 16470 255
rect 16440 205 16445 225
rect 16465 205 16470 225
rect 16440 175 16470 205
rect 16440 155 16445 175
rect 16465 155 16470 175
rect 16440 145 16470 155
rect 16495 225 16525 235
rect 16495 205 16500 225
rect 16520 205 16525 225
rect 16495 175 16525 205
rect 16495 155 16500 175
rect 16520 155 16525 175
rect 16495 125 16525 155
rect 16550 225 16580 255
rect 16550 205 16555 225
rect 16575 205 16580 225
rect 16550 175 16580 205
rect 16550 155 16555 175
rect 16575 155 16580 175
rect 16550 145 16580 155
rect 16605 225 16635 235
rect 16605 205 16610 225
rect 16630 205 16635 225
rect 16605 175 16635 205
rect 16605 155 16610 175
rect 16630 155 16635 175
rect 16605 125 16635 155
rect 16660 225 16690 255
rect 16660 205 16665 225
rect 16685 205 16690 225
rect 16660 175 16690 205
rect 16660 155 16665 175
rect 16685 155 16690 175
rect 16660 145 16690 155
rect 16485 120 16525 125
rect 16485 90 16490 120
rect 16520 90 16525 120
rect 16485 85 16525 90
rect 16545 115 16585 125
rect 16545 95 16555 115
rect 16575 95 16585 115
rect 16545 85 16585 95
rect 16605 120 16645 125
rect 16605 90 16610 120
rect 16640 90 16645 120
rect 16605 85 16645 90
rect 16315 -35 16355 -30
rect 16315 -65 16320 -35
rect 16350 -65 16355 -35
rect 16315 -70 16355 -65
rect 16260 -90 16300 -85
rect 16260 -120 16265 -90
rect 16295 -120 16300 -90
rect 16260 -125 16300 -120
rect 16205 -145 16245 -140
rect 16205 -175 16210 -145
rect 16240 -175 16245 -145
rect 16205 -180 16245 -175
rect 16095 -390 16135 -385
rect 16095 -420 16100 -390
rect 16130 -420 16135 -390
rect 15905 -620 16025 -615
rect 15905 -650 15910 -620
rect 15940 -650 15950 -620
rect 15980 -650 15990 -620
rect 16020 -650 16025 -620
rect 15905 -660 16025 -650
rect 15905 -690 15910 -660
rect 15940 -690 15950 -660
rect 15980 -690 15990 -660
rect 16020 -690 16025 -660
rect 15905 -700 16025 -690
rect 15905 -730 15910 -700
rect 15940 -730 15950 -700
rect 15980 -730 15990 -700
rect 16020 -730 16025 -700
rect 15905 -4370 16025 -730
rect 16095 -3215 16135 -420
rect 16215 -1800 16235 -180
rect 16270 -750 16290 -125
rect 16260 -755 16300 -750
rect 16260 -785 16265 -755
rect 16295 -785 16300 -755
rect 16260 -790 16300 -785
rect 16205 -1805 16245 -1800
rect 16205 -1835 16210 -1805
rect 16240 -1835 16245 -1805
rect 16205 -1840 16245 -1835
rect 16040 -3220 16080 -3215
rect 16040 -3250 16045 -3220
rect 16075 -3250 16080 -3220
rect 16040 -4300 16080 -3250
rect 16100 -3221 16135 -3215
rect 16100 -3261 16135 -3256
rect 16205 -1945 16245 -1940
rect 16205 -1975 16210 -1945
rect 16240 -1975 16245 -1945
rect 16205 -3320 16245 -1975
rect 16270 -2095 16290 -790
rect 16325 -1070 16345 -70
rect 16420 -255 16460 -250
rect 16420 -285 16425 -255
rect 16455 -285 16460 -255
rect 16420 -295 16460 -285
rect 16420 -325 16425 -295
rect 16455 -325 16460 -295
rect 16420 -335 16460 -325
rect 16420 -365 16425 -335
rect 16455 -365 16460 -335
rect 16420 -370 16460 -365
rect 16425 -395 16455 -370
rect 16425 -415 16430 -395
rect 16450 -415 16455 -395
rect 16425 -455 16455 -415
rect 16480 -390 16520 85
rect 16555 -140 16575 85
rect 16790 -85 16810 255
rect 16975 225 17005 255
rect 16975 205 16980 225
rect 17000 205 17005 225
rect 16975 175 17005 205
rect 16975 155 16980 175
rect 17000 155 17005 175
rect 16975 125 17005 155
rect 16975 105 16980 125
rect 17000 105 17005 125
rect 16975 75 17005 105
rect 16975 55 16980 75
rect 17000 55 17005 75
rect 16975 45 17005 55
rect 17065 325 17095 335
rect 17065 305 17070 325
rect 17090 305 17095 325
rect 17065 275 17095 305
rect 17065 255 17070 275
rect 17090 255 17095 275
rect 17065 225 17095 255
rect 17065 205 17070 225
rect 17090 205 17095 225
rect 17065 175 17095 205
rect 17065 155 17070 175
rect 17090 155 17095 175
rect 17065 125 17095 155
rect 17065 105 17070 125
rect 17090 105 17095 125
rect 17065 75 17095 105
rect 17065 55 17070 75
rect 17090 55 17095 75
rect 16780 -90 16820 -85
rect 16780 -120 16785 -90
rect 16815 -120 16820 -90
rect 16780 -125 16820 -120
rect 16545 -145 16585 -140
rect 16545 -175 16550 -145
rect 16580 -175 16585 -145
rect 16545 -180 16585 -175
rect 17065 -195 17095 55
rect 17155 325 17185 335
rect 17155 305 17160 325
rect 17180 305 17185 325
rect 17155 275 17185 305
rect 17155 255 17160 275
rect 17180 255 17185 275
rect 17155 225 17185 255
rect 17155 205 17160 225
rect 17180 205 17185 225
rect 17155 175 17185 205
rect 17155 155 17160 175
rect 17180 155 17185 175
rect 17155 125 17185 155
rect 17155 105 17160 125
rect 17180 105 17185 125
rect 17155 75 17185 105
rect 17155 55 17160 75
rect 17180 55 17185 75
rect 17155 45 17185 55
rect 17245 325 17275 335
rect 17245 305 17250 325
rect 17270 305 17275 325
rect 17245 275 17275 305
rect 17245 255 17250 275
rect 17270 255 17275 275
rect 17245 225 17275 255
rect 17245 205 17250 225
rect 17270 205 17275 225
rect 17245 175 17275 205
rect 17245 155 17250 175
rect 17270 155 17275 175
rect 17245 125 17275 155
rect 17245 105 17250 125
rect 17270 105 17275 125
rect 17245 75 17275 105
rect 17245 55 17250 75
rect 17270 55 17275 75
rect 17245 45 17275 55
rect 17335 325 17365 335
rect 17335 305 17340 325
rect 17360 305 17365 325
rect 17335 275 17365 305
rect 17335 255 17340 275
rect 17360 255 17365 275
rect 17335 225 17365 255
rect 17335 205 17340 225
rect 17360 205 17365 225
rect 17335 175 17365 205
rect 17335 155 17340 175
rect 17360 155 17365 175
rect 17335 125 17365 155
rect 17335 105 17340 125
rect 17360 105 17365 125
rect 17335 75 17365 105
rect 17335 55 17340 75
rect 17360 55 17365 75
rect 17335 45 17365 55
rect 17425 325 17455 335
rect 17425 305 17430 325
rect 17450 305 17455 325
rect 17425 275 17455 305
rect 17425 255 17430 275
rect 17450 255 17455 275
rect 17425 225 17455 255
rect 17425 205 17430 225
rect 17450 205 17455 225
rect 17425 175 17455 205
rect 17425 155 17430 175
rect 17450 155 17455 175
rect 17425 125 17455 155
rect 17425 105 17430 125
rect 17450 105 17455 125
rect 17425 75 17455 105
rect 17425 55 17430 75
rect 17450 55 17455 75
rect 17425 45 17455 55
rect 17515 325 17545 335
rect 17515 305 17520 325
rect 17540 305 17545 325
rect 17515 275 17545 305
rect 17515 255 17520 275
rect 17540 255 17545 275
rect 17515 225 17545 255
rect 17515 205 17520 225
rect 17540 205 17545 225
rect 17515 175 17545 205
rect 17515 155 17520 175
rect 17540 155 17545 175
rect 17515 125 17545 155
rect 17515 105 17520 125
rect 17540 105 17545 125
rect 17515 75 17545 105
rect 17515 55 17520 75
rect 17540 55 17545 75
rect 17515 45 17545 55
rect 17605 325 17635 335
rect 17605 305 17610 325
rect 17630 305 17635 325
rect 17605 275 17635 305
rect 17605 255 17610 275
rect 17630 255 17635 275
rect 17605 225 17635 255
rect 17605 205 17610 225
rect 17630 205 17635 225
rect 17605 175 17635 205
rect 17605 155 17610 175
rect 17630 155 17635 175
rect 17605 125 17635 155
rect 17605 105 17610 125
rect 17630 105 17635 125
rect 17605 75 17635 105
rect 17605 55 17610 75
rect 17630 55 17635 75
rect 17605 45 17635 55
rect 17695 325 17725 335
rect 17695 305 17700 325
rect 17720 305 17725 325
rect 17695 275 17725 305
rect 17695 255 17700 275
rect 17720 255 17725 275
rect 17695 225 17725 255
rect 17695 205 17700 225
rect 17720 205 17725 225
rect 17695 175 17725 205
rect 17695 155 17700 175
rect 17720 155 17725 175
rect 17695 125 17725 155
rect 17695 105 17700 125
rect 17720 105 17725 125
rect 17695 75 17725 105
rect 17695 55 17700 75
rect 17720 55 17725 75
rect 17695 45 17725 55
rect 17785 325 17815 335
rect 17785 305 17790 325
rect 17810 305 17815 325
rect 17785 275 17815 305
rect 17785 255 17790 275
rect 17810 255 17815 275
rect 17785 225 17815 255
rect 17785 205 17790 225
rect 17810 205 17815 225
rect 17785 175 17815 205
rect 17785 155 17790 175
rect 17810 155 17815 175
rect 17785 125 17815 155
rect 17785 105 17790 125
rect 17810 105 17815 125
rect 17785 75 17815 105
rect 17785 55 17790 75
rect 17810 55 17815 75
rect 17110 20 17145 25
rect 17140 -10 17145 20
rect 17110 -15 17145 -10
rect 17195 20 17235 25
rect 17195 -10 17200 20
rect 17230 -10 17235 20
rect 17195 -15 17235 -10
rect 17250 -140 17270 45
rect 17285 20 17325 25
rect 17285 -10 17290 20
rect 17320 -10 17325 20
rect 17285 -15 17325 -10
rect 17375 20 17415 25
rect 17375 -10 17380 20
rect 17410 -10 17415 20
rect 17375 -15 17415 -10
rect 17430 -85 17450 45
rect 17465 20 17505 25
rect 17465 -10 17470 20
rect 17500 -10 17505 20
rect 17465 -15 17505 -10
rect 17555 20 17595 25
rect 17555 -10 17560 20
rect 17590 -10 17595 20
rect 17555 -15 17595 -10
rect 17610 -30 17630 45
rect 17645 20 17770 25
rect 17645 -10 17650 20
rect 17680 -10 17695 20
rect 17725 -10 17740 20
rect 17645 -15 17770 -10
rect 17600 -35 17640 -30
rect 17600 -65 17605 -35
rect 17635 -65 17640 -35
rect 17600 -70 17640 -65
rect 17420 -90 17460 -85
rect 17420 -120 17425 -90
rect 17455 -120 17460 -90
rect 17420 -125 17460 -120
rect 17240 -145 17280 -140
rect 17240 -175 17245 -145
rect 17275 -175 17280 -145
rect 17240 -180 17280 -175
rect 17060 -200 17100 -195
rect 17060 -230 17065 -200
rect 17095 -230 17100 -200
rect 17060 -235 17100 -230
rect 16540 -255 16580 -250
rect 16540 -285 16545 -255
rect 16575 -285 16580 -255
rect 16540 -295 16580 -285
rect 16540 -325 16545 -295
rect 16575 -325 16580 -295
rect 16540 -335 16580 -325
rect 16540 -365 16545 -335
rect 16575 -365 16580 -335
rect 16540 -370 16580 -365
rect 16660 -255 16700 -250
rect 16660 -285 16665 -255
rect 16695 -285 16700 -255
rect 16660 -295 16700 -285
rect 16660 -325 16665 -295
rect 16695 -325 16700 -295
rect 16660 -335 16700 -325
rect 16660 -365 16665 -335
rect 16695 -365 16700 -335
rect 16660 -370 16700 -365
rect 16780 -255 16820 -250
rect 16780 -285 16785 -255
rect 16815 -285 16820 -255
rect 16780 -295 16820 -285
rect 16780 -325 16785 -295
rect 16815 -325 16820 -295
rect 16780 -335 16820 -325
rect 16780 -365 16785 -335
rect 16815 -365 16820 -335
rect 16780 -370 16820 -365
rect 16900 -255 16940 -250
rect 16900 -285 16905 -255
rect 16935 -285 16940 -255
rect 16900 -295 16940 -285
rect 16900 -325 16905 -295
rect 16935 -325 16940 -295
rect 16900 -335 16940 -325
rect 16900 -365 16905 -335
rect 16935 -365 16940 -335
rect 16900 -370 16940 -365
rect 17020 -255 17060 -250
rect 17020 -285 17025 -255
rect 17055 -285 17060 -255
rect 17020 -295 17060 -285
rect 17020 -325 17025 -295
rect 17055 -325 17060 -295
rect 17020 -335 17060 -325
rect 17020 -365 17025 -335
rect 17055 -365 17060 -335
rect 17020 -370 17060 -365
rect 17140 -255 17180 -250
rect 17140 -285 17145 -255
rect 17175 -285 17180 -255
rect 17140 -295 17180 -285
rect 17140 -325 17145 -295
rect 17175 -325 17180 -295
rect 17140 -335 17180 -325
rect 17140 -365 17145 -335
rect 17175 -365 17180 -335
rect 17140 -370 17180 -365
rect 17260 -255 17300 -250
rect 17260 -285 17265 -255
rect 17295 -285 17300 -255
rect 17260 -295 17300 -285
rect 17260 -325 17265 -295
rect 17295 -325 17300 -295
rect 17260 -335 17300 -325
rect 17260 -365 17265 -335
rect 17295 -365 17300 -335
rect 17260 -370 17300 -365
rect 17380 -255 17420 -250
rect 17380 -285 17385 -255
rect 17415 -285 17420 -255
rect 17380 -295 17420 -285
rect 17380 -325 17385 -295
rect 17415 -325 17420 -295
rect 17380 -335 17420 -325
rect 17380 -365 17385 -335
rect 17415 -365 17420 -335
rect 17380 -370 17420 -365
rect 17500 -255 17540 -250
rect 17500 -285 17505 -255
rect 17535 -285 17540 -255
rect 17500 -295 17540 -285
rect 17500 -325 17505 -295
rect 17535 -325 17540 -295
rect 17500 -335 17540 -325
rect 17500 -365 17505 -335
rect 17535 -365 17540 -335
rect 17500 -370 17540 -365
rect 17620 -255 17660 -250
rect 17620 -285 17625 -255
rect 17655 -285 17660 -255
rect 17620 -295 17660 -285
rect 17620 -325 17625 -295
rect 17655 -325 17660 -295
rect 17620 -335 17660 -325
rect 17620 -365 17625 -335
rect 17655 -365 17660 -335
rect 17620 -370 17660 -365
rect 16480 -420 16485 -390
rect 16515 -420 16520 -390
rect 16480 -425 16520 -420
rect 16425 -475 16430 -455
rect 16450 -475 16455 -455
rect 16425 -505 16455 -475
rect 16425 -525 16430 -505
rect 16450 -525 16455 -505
rect 16425 -535 16455 -525
rect 16485 -455 16515 -425
rect 16485 -475 16490 -455
rect 16510 -475 16515 -455
rect 16485 -505 16515 -475
rect 16485 -525 16490 -505
rect 16510 -525 16515 -505
rect 16485 -535 16515 -525
rect 16545 -455 16575 -370
rect 16545 -475 16550 -455
rect 16570 -475 16575 -455
rect 16545 -505 16575 -475
rect 16545 -525 16550 -505
rect 16570 -525 16575 -505
rect 16545 -535 16575 -525
rect 16605 -455 16635 -445
rect 16605 -475 16610 -455
rect 16630 -475 16635 -455
rect 16605 -505 16635 -475
rect 16605 -525 16610 -505
rect 16630 -525 16635 -505
rect 16605 -555 16635 -525
rect 16665 -455 16695 -370
rect 16665 -475 16670 -455
rect 16690 -475 16695 -455
rect 16665 -505 16695 -475
rect 16665 -525 16670 -505
rect 16690 -525 16695 -505
rect 16665 -535 16695 -525
rect 16725 -455 16755 -445
rect 16725 -475 16730 -455
rect 16750 -475 16755 -455
rect 16725 -505 16755 -475
rect 16725 -525 16730 -505
rect 16750 -525 16755 -505
rect 16600 -560 16640 -555
rect 16515 -570 16545 -560
rect 16515 -590 16520 -570
rect 16540 -590 16545 -570
rect 16515 -615 16545 -590
rect 16600 -590 16605 -560
rect 16635 -590 16640 -560
rect 16600 -595 16640 -590
rect 16725 -615 16755 -525
rect 16785 -455 16815 -370
rect 16840 -390 16880 -385
rect 16840 -420 16845 -390
rect 16875 -420 16880 -390
rect 16840 -425 16880 -420
rect 16785 -475 16790 -455
rect 16810 -475 16815 -455
rect 16785 -505 16815 -475
rect 16785 -525 16790 -505
rect 16810 -525 16815 -505
rect 16785 -535 16815 -525
rect 16845 -455 16875 -425
rect 16845 -475 16850 -455
rect 16870 -475 16875 -455
rect 16845 -505 16875 -475
rect 16845 -525 16850 -505
rect 16870 -525 16875 -505
rect 16845 -535 16875 -525
rect 16905 -455 16935 -370
rect 16905 -475 16910 -455
rect 16930 -475 16935 -455
rect 16905 -505 16935 -475
rect 16905 -525 16910 -505
rect 16930 -525 16935 -505
rect 16905 -535 16935 -525
rect 16965 -455 16995 -445
rect 16965 -475 16970 -455
rect 16990 -475 16995 -455
rect 16965 -505 16995 -475
rect 16965 -525 16970 -505
rect 16990 -525 16995 -505
rect 16965 -555 16995 -525
rect 17025 -455 17055 -370
rect 17025 -475 17030 -455
rect 17050 -475 17055 -455
rect 17025 -505 17055 -475
rect 17025 -525 17030 -505
rect 17050 -525 17055 -505
rect 17025 -535 17055 -525
rect 17085 -455 17115 -445
rect 17085 -475 17090 -455
rect 17110 -475 17115 -455
rect 17085 -505 17115 -475
rect 17085 -525 17090 -505
rect 17110 -525 17115 -505
rect 16845 -565 16875 -555
rect 16845 -585 16850 -565
rect 16870 -585 16875 -565
rect 16845 -615 16875 -585
rect 16960 -560 17000 -555
rect 16960 -590 16965 -560
rect 16995 -590 17000 -560
rect 16960 -595 17000 -590
rect 16510 -620 16550 -615
rect 16510 -650 16515 -620
rect 16545 -650 16550 -620
rect 16510 -660 16550 -650
rect 16510 -690 16515 -660
rect 16545 -690 16550 -660
rect 16510 -700 16550 -690
rect 16510 -730 16515 -700
rect 16545 -730 16550 -700
rect 16510 -735 16550 -730
rect 16720 -620 16760 -615
rect 16720 -650 16725 -620
rect 16755 -650 16760 -620
rect 16720 -660 16760 -650
rect 16720 -690 16725 -660
rect 16755 -690 16760 -660
rect 16720 -700 16760 -690
rect 16720 -730 16725 -700
rect 16755 -730 16760 -700
rect 16720 -735 16760 -730
rect 16840 -620 16880 -615
rect 16840 -650 16845 -620
rect 16875 -650 16880 -620
rect 16840 -660 16880 -650
rect 16840 -690 16845 -660
rect 16875 -690 16880 -660
rect 16840 -700 16880 -690
rect 16840 -730 16845 -700
rect 16875 -730 16880 -700
rect 16840 -735 16880 -730
rect 16970 -810 16990 -595
rect 17085 -615 17115 -525
rect 17145 -455 17175 -370
rect 17200 -390 17240 -385
rect 17200 -420 17205 -390
rect 17235 -420 17240 -390
rect 17200 -425 17240 -420
rect 17145 -475 17150 -455
rect 17170 -475 17175 -455
rect 17145 -505 17175 -475
rect 17145 -525 17150 -505
rect 17170 -525 17175 -505
rect 17145 -535 17175 -525
rect 17205 -455 17235 -425
rect 17205 -475 17210 -455
rect 17230 -475 17235 -455
rect 17205 -505 17235 -475
rect 17205 -525 17210 -505
rect 17230 -525 17235 -505
rect 17205 -535 17235 -525
rect 17265 -455 17295 -370
rect 17265 -475 17270 -455
rect 17290 -475 17295 -455
rect 17265 -505 17295 -475
rect 17265 -525 17270 -505
rect 17290 -525 17295 -505
rect 17265 -535 17295 -525
rect 17325 -455 17355 -445
rect 17325 -475 17330 -455
rect 17350 -475 17355 -455
rect 17325 -505 17355 -475
rect 17325 -525 17330 -505
rect 17350 -525 17355 -505
rect 17325 -555 17355 -525
rect 17385 -455 17415 -370
rect 17385 -475 17390 -455
rect 17410 -475 17415 -455
rect 17385 -505 17415 -475
rect 17385 -525 17390 -505
rect 17410 -525 17415 -505
rect 17385 -535 17415 -525
rect 17445 -455 17475 -445
rect 17445 -475 17450 -455
rect 17470 -475 17475 -455
rect 17445 -505 17475 -475
rect 17445 -525 17450 -505
rect 17470 -525 17475 -505
rect 17205 -565 17235 -555
rect 17205 -585 17210 -565
rect 17230 -585 17235 -565
rect 17205 -615 17235 -585
rect 17320 -560 17360 -555
rect 17320 -590 17325 -560
rect 17355 -590 17360 -560
rect 17320 -595 17360 -590
rect 17445 -615 17475 -525
rect 17505 -455 17535 -370
rect 17560 -390 17600 -385
rect 17560 -420 17565 -390
rect 17595 -420 17600 -390
rect 17560 -425 17600 -420
rect 17625 -395 17655 -370
rect 17625 -415 17630 -395
rect 17650 -415 17655 -395
rect 17505 -475 17510 -455
rect 17530 -475 17535 -455
rect 17505 -505 17535 -475
rect 17505 -525 17510 -505
rect 17530 -525 17535 -505
rect 17505 -535 17535 -525
rect 17565 -455 17595 -425
rect 17565 -475 17570 -455
rect 17590 -475 17595 -455
rect 17565 -505 17595 -475
rect 17565 -525 17570 -505
rect 17590 -525 17595 -505
rect 17565 -535 17595 -525
rect 17625 -455 17655 -415
rect 17690 -390 17730 -15
rect 17785 -195 17815 55
rect 17875 325 17905 335
rect 17875 305 17880 325
rect 17900 305 17905 325
rect 17875 275 17905 305
rect 17875 255 17880 275
rect 17900 255 17905 275
rect 17875 225 17905 255
rect 17875 205 17880 225
rect 17900 205 17905 225
rect 17875 175 17905 205
rect 17875 155 17880 175
rect 17900 155 17905 175
rect 17875 125 17905 155
rect 17875 105 17880 125
rect 17900 105 17905 125
rect 17875 75 17905 105
rect 17875 55 17880 75
rect 17900 55 17905 75
rect 17875 45 17905 55
rect 17965 325 17995 335
rect 17965 305 17970 325
rect 17990 305 17995 325
rect 17965 275 17995 305
rect 17965 255 17970 275
rect 17990 255 17995 275
rect 17965 225 17995 255
rect 17965 205 17970 225
rect 17990 205 17995 225
rect 17965 175 17995 205
rect 17965 155 17970 175
rect 17990 155 17995 175
rect 17965 125 17995 155
rect 17965 105 17970 125
rect 17990 105 17995 125
rect 17965 75 17995 105
rect 17965 55 17970 75
rect 17990 55 17995 75
rect 17965 45 17995 55
rect 18055 325 18085 335
rect 18055 305 18060 325
rect 18080 305 18085 325
rect 18055 275 18085 305
rect 18055 255 18060 275
rect 18080 255 18085 275
rect 18055 225 18085 255
rect 18055 205 18060 225
rect 18080 205 18085 225
rect 18055 175 18085 205
rect 18055 155 18060 175
rect 18080 155 18085 175
rect 18055 125 18085 155
rect 18055 105 18060 125
rect 18080 105 18085 125
rect 18055 75 18085 105
rect 18055 55 18060 75
rect 18080 55 18085 75
rect 18055 45 18085 55
rect 18145 325 18175 335
rect 18145 305 18150 325
rect 18170 305 18175 325
rect 18145 275 18175 305
rect 18145 255 18150 275
rect 18170 255 18175 275
rect 18145 225 18175 255
rect 18145 205 18150 225
rect 18170 205 18175 225
rect 18145 175 18175 205
rect 18145 155 18150 175
rect 18170 155 18175 175
rect 18145 125 18175 155
rect 18145 105 18150 125
rect 18170 105 18175 125
rect 18145 75 18175 105
rect 18145 55 18150 75
rect 18170 55 18175 75
rect 18145 45 18175 55
rect 18235 325 18265 335
rect 18235 305 18240 325
rect 18260 305 18265 325
rect 18235 275 18265 305
rect 18235 255 18240 275
rect 18260 255 18265 275
rect 18235 225 18265 255
rect 18235 205 18240 225
rect 18260 205 18265 225
rect 18235 175 18265 205
rect 18235 155 18240 175
rect 18260 155 18265 175
rect 18235 125 18265 155
rect 18235 105 18240 125
rect 18260 105 18265 125
rect 18235 75 18265 105
rect 18235 55 18240 75
rect 18260 55 18265 75
rect 18235 45 18265 55
rect 18325 325 18355 335
rect 18325 305 18330 325
rect 18350 305 18355 325
rect 18325 275 18355 305
rect 18325 255 18330 275
rect 18350 255 18355 275
rect 18325 225 18355 255
rect 18325 205 18330 225
rect 18350 205 18355 225
rect 18325 175 18355 205
rect 18325 155 18330 175
rect 18350 155 18355 175
rect 18325 125 18355 155
rect 18325 105 18330 125
rect 18350 105 18355 125
rect 18325 75 18355 105
rect 18325 55 18330 75
rect 18350 55 18355 75
rect 18325 45 18355 55
rect 18415 325 18445 335
rect 18415 305 18420 325
rect 18440 305 18445 325
rect 18415 275 18445 305
rect 18415 255 18420 275
rect 18440 255 18445 275
rect 18415 225 18445 255
rect 18415 205 18420 225
rect 18440 205 18445 225
rect 18415 175 18445 205
rect 18415 155 18420 175
rect 18440 155 18445 175
rect 18415 125 18445 155
rect 18415 105 18420 125
rect 18440 105 18445 125
rect 18415 75 18445 105
rect 18415 55 18420 75
rect 18440 55 18445 75
rect 18415 45 18445 55
rect 18505 325 18535 335
rect 18505 305 18510 325
rect 18530 305 18535 325
rect 18505 275 18535 305
rect 18505 255 18510 275
rect 18530 255 18535 275
rect 18505 225 18535 255
rect 18505 205 18510 225
rect 18530 205 18535 225
rect 18505 175 18535 205
rect 18505 155 18510 175
rect 18530 155 18535 175
rect 18505 125 18535 155
rect 18505 105 18510 125
rect 18530 105 18535 125
rect 18505 75 18535 105
rect 18505 55 18510 75
rect 18530 55 18535 75
rect 17830 20 17865 25
rect 17860 -10 17865 20
rect 17830 -15 17865 -10
rect 17915 20 17955 25
rect 17915 -10 17920 20
rect 17950 -10 17955 20
rect 17915 -15 17955 -10
rect 17970 -30 17990 45
rect 18005 20 18045 25
rect 18005 -10 18010 20
rect 18040 -10 18045 20
rect 18005 -15 18045 -10
rect 18095 20 18135 25
rect 18095 -10 18100 20
rect 18130 -10 18135 20
rect 18095 -15 18135 -10
rect 17960 -35 18000 -30
rect 17960 -65 17965 -35
rect 17995 -65 18000 -35
rect 17960 -70 18000 -65
rect 18150 -85 18170 45
rect 18185 20 18225 25
rect 18185 -10 18190 20
rect 18220 -10 18225 20
rect 18185 -15 18225 -10
rect 18275 20 18315 25
rect 18275 -10 18280 20
rect 18310 -10 18315 20
rect 18275 -15 18315 -10
rect 18140 -90 18180 -85
rect 18140 -120 18145 -90
rect 18175 -120 18180 -90
rect 18140 -125 18180 -120
rect 18330 -140 18350 45
rect 18365 20 18405 25
rect 18365 -10 18370 20
rect 18400 -10 18405 20
rect 18365 -15 18405 -10
rect 18455 20 18490 25
rect 18455 -10 18460 20
rect 18455 -15 18490 -10
rect 18320 -145 18360 -140
rect 18320 -175 18325 -145
rect 18355 -175 18360 -145
rect 18320 -180 18360 -175
rect 18505 -195 18535 55
rect 18595 325 18625 335
rect 18595 305 18600 325
rect 18620 305 18625 325
rect 18595 275 18625 305
rect 18595 255 18600 275
rect 18620 255 18625 275
rect 18595 225 18625 255
rect 18595 205 18600 225
rect 18620 205 18625 225
rect 18595 175 18625 205
rect 18595 155 18600 175
rect 18620 155 18625 175
rect 18595 125 18625 155
rect 18595 105 18600 125
rect 18620 105 18625 125
rect 18595 75 18625 105
rect 18595 55 18600 75
rect 18620 55 18625 75
rect 18595 45 18625 55
rect 17780 -200 17820 -195
rect 17780 -230 17785 -200
rect 17815 -230 17820 -200
rect 17780 -235 17820 -230
rect 18500 -200 18540 -195
rect 18500 -230 18505 -200
rect 18535 -230 18540 -200
rect 18500 -235 18540 -230
rect 17940 -255 17980 -250
rect 17940 -285 17945 -255
rect 17975 -285 17980 -255
rect 17940 -295 17980 -285
rect 17940 -325 17945 -295
rect 17975 -325 17980 -295
rect 17940 -335 17980 -325
rect 17940 -365 17945 -335
rect 17975 -365 17980 -335
rect 17940 -370 17980 -365
rect 18060 -255 18100 -250
rect 18060 -285 18065 -255
rect 18095 -285 18100 -255
rect 18060 -295 18100 -285
rect 18060 -325 18065 -295
rect 18095 -325 18100 -295
rect 18060 -335 18100 -325
rect 18060 -365 18065 -335
rect 18095 -365 18100 -335
rect 18060 -370 18100 -365
rect 18180 -255 18220 -250
rect 18180 -285 18185 -255
rect 18215 -285 18220 -255
rect 18180 -295 18220 -285
rect 18180 -325 18185 -295
rect 18215 -325 18220 -295
rect 18180 -335 18220 -325
rect 18180 -365 18185 -335
rect 18215 -365 18220 -335
rect 18180 -370 18220 -365
rect 18300 -255 18340 -250
rect 18300 -285 18305 -255
rect 18335 -285 18340 -255
rect 18300 -295 18340 -285
rect 18300 -325 18305 -295
rect 18335 -325 18340 -295
rect 18300 -335 18340 -325
rect 18300 -365 18305 -335
rect 18335 -365 18340 -335
rect 18300 -370 18340 -365
rect 18420 -255 18460 -250
rect 18420 -285 18425 -255
rect 18455 -285 18460 -255
rect 18420 -295 18460 -285
rect 18420 -325 18425 -295
rect 18455 -325 18460 -295
rect 18420 -335 18460 -325
rect 18420 -365 18425 -335
rect 18455 -365 18460 -335
rect 18420 -370 18460 -365
rect 18540 -255 18580 -250
rect 18540 -285 18545 -255
rect 18575 -285 18580 -255
rect 18540 -295 18580 -285
rect 18540 -325 18545 -295
rect 18575 -325 18580 -295
rect 18540 -335 18580 -325
rect 18540 -365 18545 -335
rect 18575 -365 18580 -335
rect 18540 -370 18580 -365
rect 18660 -255 18700 -250
rect 18660 -285 18665 -255
rect 18695 -285 18700 -255
rect 18660 -295 18700 -285
rect 18660 -325 18665 -295
rect 18695 -325 18700 -295
rect 18660 -335 18700 -325
rect 18660 -365 18665 -335
rect 18695 -365 18700 -335
rect 18660 -370 18700 -365
rect 18780 -255 18820 -250
rect 18780 -285 18785 -255
rect 18815 -285 18820 -255
rect 18780 -295 18820 -285
rect 18780 -325 18785 -295
rect 18815 -325 18820 -295
rect 18780 -335 18820 -325
rect 18780 -365 18785 -335
rect 18815 -365 18820 -335
rect 18780 -370 18820 -365
rect 18900 -255 18940 -250
rect 18900 -285 18905 -255
rect 18935 -285 18940 -255
rect 18900 -295 18940 -285
rect 18900 -325 18905 -295
rect 18935 -325 18940 -295
rect 18900 -335 18940 -325
rect 18900 -365 18905 -335
rect 18935 -365 18940 -335
rect 18900 -370 18940 -365
rect 19020 -255 19060 -250
rect 19020 -285 19025 -255
rect 19055 -285 19060 -255
rect 19020 -295 19060 -285
rect 19020 -325 19025 -295
rect 19055 -325 19060 -295
rect 19020 -335 19060 -325
rect 19020 -365 19025 -335
rect 19055 -365 19060 -335
rect 19020 -370 19060 -365
rect 19140 -255 19180 -250
rect 19140 -285 19145 -255
rect 19175 -285 19180 -255
rect 19140 -295 19180 -285
rect 19140 -325 19145 -295
rect 19175 -325 19180 -295
rect 19140 -335 19180 -325
rect 19140 -365 19145 -335
rect 19175 -365 19180 -335
rect 19140 -370 19180 -365
rect 17690 -420 17695 -390
rect 17725 -420 17730 -390
rect 17690 -425 17730 -420
rect 17870 -390 17910 -385
rect 17870 -420 17875 -390
rect 17905 -420 17910 -390
rect 17870 -425 17910 -420
rect 17945 -395 17975 -370
rect 17945 -415 17950 -395
rect 17970 -415 17975 -395
rect 17625 -475 17630 -455
rect 17650 -475 17655 -455
rect 17625 -505 17655 -475
rect 17625 -525 17630 -505
rect 17650 -525 17655 -505
rect 17625 -535 17655 -525
rect 17535 -565 17565 -555
rect 17535 -585 17540 -565
rect 17560 -585 17565 -565
rect 17535 -615 17565 -585
rect 17080 -620 17120 -615
rect 17080 -650 17085 -620
rect 17115 -650 17120 -620
rect 17080 -660 17120 -650
rect 17080 -690 17085 -660
rect 17115 -690 17120 -660
rect 17080 -700 17120 -690
rect 17080 -730 17085 -700
rect 17115 -730 17120 -700
rect 17080 -735 17120 -730
rect 17200 -620 17240 -615
rect 17200 -650 17205 -620
rect 17235 -650 17240 -620
rect 17200 -660 17240 -650
rect 17200 -690 17205 -660
rect 17235 -690 17240 -660
rect 17200 -700 17240 -690
rect 17200 -730 17205 -700
rect 17235 -730 17240 -700
rect 17200 -735 17240 -730
rect 17440 -620 17480 -615
rect 17440 -650 17445 -620
rect 17475 -650 17480 -620
rect 17440 -660 17480 -650
rect 17440 -690 17445 -660
rect 17475 -690 17480 -660
rect 17440 -700 17480 -690
rect 17440 -730 17445 -700
rect 17475 -730 17480 -700
rect 17440 -735 17480 -730
rect 17530 -620 17570 -615
rect 17530 -650 17535 -620
rect 17565 -650 17570 -620
rect 17530 -660 17570 -650
rect 17530 -690 17535 -660
rect 17565 -690 17570 -660
rect 17530 -700 17570 -690
rect 17530 -730 17535 -700
rect 17565 -730 17570 -700
rect 17530 -735 17570 -730
rect 17007 -755 17037 -750
rect 17007 -790 17037 -785
rect 17090 -810 17110 -735
rect 16965 -820 16995 -810
rect 16965 -840 16970 -820
rect 16990 -840 16995 -820
rect 16965 -870 16995 -840
rect 16965 -890 16970 -870
rect 16990 -890 16995 -870
rect 16965 -920 16995 -890
rect 16965 -940 16970 -920
rect 16990 -940 16995 -920
rect 16965 -970 16995 -940
rect 16965 -990 16970 -970
rect 16990 -990 16995 -970
rect 16965 -1020 16995 -990
rect 16965 -1040 16970 -1020
rect 16990 -1040 16995 -1020
rect 16965 -1050 16995 -1040
rect 17025 -820 17055 -810
rect 17025 -840 17030 -820
rect 17050 -840 17055 -820
rect 17025 -870 17055 -840
rect 17025 -890 17030 -870
rect 17050 -890 17055 -870
rect 17025 -920 17055 -890
rect 17025 -940 17030 -920
rect 17050 -940 17055 -920
rect 17025 -970 17055 -940
rect 17025 -990 17030 -970
rect 17050 -990 17055 -970
rect 17025 -1020 17055 -990
rect 17025 -1040 17030 -1020
rect 17050 -1040 17055 -1020
rect 16315 -1075 16355 -1070
rect 16315 -1105 16320 -1075
rect 16350 -1105 16355 -1075
rect 16315 -1110 16355 -1105
rect 16325 -1995 16345 -1110
rect 17025 -1125 17055 -1040
rect 17085 -820 17115 -810
rect 17085 -840 17090 -820
rect 17110 -840 17115 -820
rect 17085 -870 17115 -840
rect 17085 -890 17090 -870
rect 17110 -890 17115 -870
rect 17085 -920 17115 -890
rect 17085 -940 17090 -920
rect 17110 -940 17115 -920
rect 17560 -815 17600 -810
rect 17560 -845 17565 -815
rect 17595 -845 17600 -815
rect 17560 -855 17600 -845
rect 17560 -885 17565 -855
rect 17595 -885 17600 -855
rect 17560 -895 17600 -885
rect 17560 -925 17565 -895
rect 17595 -925 17600 -895
rect 17560 -930 17600 -925
rect 17085 -970 17115 -940
rect 17085 -990 17090 -970
rect 17110 -990 17115 -970
rect 17085 -1020 17115 -990
rect 17085 -1040 17090 -1020
rect 17110 -1040 17115 -1020
rect 17085 -1050 17115 -1040
rect 17075 -1075 17105 -1070
rect 17075 -1110 17105 -1105
rect 16530 -1130 16570 -1125
rect 16530 -1160 16535 -1130
rect 16565 -1160 16570 -1130
rect 16530 -1165 16570 -1160
rect 17020 -1130 17060 -1125
rect 17020 -1160 17025 -1130
rect 17055 -1160 17060 -1130
rect 17020 -1165 17060 -1160
rect 16535 -1330 16565 -1165
rect 16620 -1185 16660 -1180
rect 16620 -1215 16625 -1185
rect 16655 -1215 16660 -1185
rect 16620 -1225 16660 -1215
rect 16620 -1255 16625 -1225
rect 16655 -1255 16660 -1225
rect 16620 -1265 16660 -1255
rect 16620 -1295 16625 -1265
rect 16655 -1295 16660 -1265
rect 16620 -1300 16660 -1295
rect 16740 -1185 16780 -1180
rect 16740 -1215 16745 -1185
rect 16775 -1215 16780 -1185
rect 16740 -1225 16780 -1215
rect 16740 -1255 16745 -1225
rect 16775 -1255 16780 -1225
rect 16740 -1265 16780 -1255
rect 16740 -1295 16745 -1265
rect 16775 -1295 16780 -1265
rect 16740 -1300 16780 -1295
rect 16860 -1185 16900 -1180
rect 16860 -1215 16865 -1185
rect 16895 -1215 16900 -1185
rect 16860 -1225 16900 -1215
rect 16860 -1255 16865 -1225
rect 16895 -1255 16900 -1225
rect 16860 -1265 16900 -1255
rect 16860 -1295 16865 -1265
rect 16895 -1295 16900 -1265
rect 16860 -1300 16900 -1295
rect 16980 -1185 17020 -1180
rect 16980 -1215 16985 -1185
rect 17015 -1215 17020 -1185
rect 16980 -1225 17020 -1215
rect 16980 -1255 16985 -1225
rect 17015 -1255 17020 -1225
rect 16980 -1265 17020 -1255
rect 16980 -1295 16985 -1265
rect 17015 -1295 17020 -1265
rect 16980 -1300 17020 -1295
rect 17300 -1185 17340 -1180
rect 17300 -1215 17305 -1185
rect 17335 -1215 17340 -1185
rect 17300 -1225 17340 -1215
rect 17300 -1255 17305 -1225
rect 17335 -1255 17340 -1225
rect 17300 -1265 17340 -1255
rect 17300 -1295 17305 -1265
rect 17335 -1295 17340 -1265
rect 17300 -1300 17340 -1295
rect 17420 -1185 17460 -1180
rect 17420 -1215 17425 -1185
rect 17455 -1215 17460 -1185
rect 17420 -1225 17460 -1215
rect 17420 -1255 17425 -1225
rect 17455 -1255 17460 -1225
rect 17420 -1265 17460 -1255
rect 17420 -1295 17425 -1265
rect 17455 -1295 17460 -1265
rect 17420 -1300 17460 -1295
rect 17540 -1185 17580 -1180
rect 17540 -1215 17545 -1185
rect 17575 -1215 17580 -1185
rect 17540 -1225 17580 -1215
rect 17540 -1255 17545 -1225
rect 17575 -1255 17580 -1225
rect 17540 -1265 17580 -1255
rect 17540 -1295 17545 -1265
rect 17575 -1295 17580 -1265
rect 17540 -1300 17580 -1295
rect 17695 -1285 17725 -425
rect 17695 -1305 17700 -1285
rect 17720 -1305 17725 -1285
rect 17695 -1315 17725 -1305
rect 17740 -815 17860 -810
rect 17740 -845 17745 -815
rect 17775 -845 17785 -815
rect 17815 -845 17825 -815
rect 17855 -845 17860 -815
rect 17740 -855 17860 -845
rect 17740 -885 17745 -855
rect 17775 -885 17785 -855
rect 17815 -885 17825 -855
rect 17855 -885 17860 -855
rect 17740 -895 17860 -885
rect 17740 -925 17745 -895
rect 17775 -925 17785 -895
rect 17815 -925 17825 -895
rect 17855 -925 17860 -895
rect 16535 -1350 16540 -1330
rect 16560 -1350 16565 -1330
rect 16535 -1380 16565 -1350
rect 16535 -1400 16540 -1380
rect 16560 -1400 16565 -1380
rect 16535 -1430 16565 -1400
rect 16535 -1450 16540 -1430
rect 16560 -1450 16565 -1430
rect 16535 -1480 16565 -1450
rect 16535 -1500 16540 -1480
rect 16560 -1500 16565 -1480
rect 16535 -1530 16565 -1500
rect 16535 -1550 16540 -1530
rect 16560 -1550 16565 -1530
rect 16535 -1560 16565 -1550
rect 17110 -1585 17150 -1580
rect 17110 -1615 17115 -1585
rect 17145 -1615 17150 -1585
rect 17110 -1625 17150 -1615
rect 17110 -1655 17115 -1625
rect 17145 -1655 17150 -1625
rect 17110 -1665 17150 -1655
rect 17110 -1695 17115 -1665
rect 17145 -1695 17150 -1665
rect 17110 -1700 17150 -1695
rect 17740 -1585 17860 -925
rect 17875 -1285 17905 -425
rect 17945 -455 17975 -415
rect 18000 -390 18040 -385
rect 18000 -420 18005 -390
rect 18035 -420 18040 -390
rect 18000 -425 18040 -420
rect 17945 -475 17950 -455
rect 17970 -475 17975 -455
rect 17945 -505 17975 -475
rect 17945 -525 17950 -505
rect 17970 -525 17975 -505
rect 17945 -535 17975 -525
rect 18005 -455 18035 -425
rect 18005 -475 18010 -455
rect 18030 -475 18035 -455
rect 18005 -505 18035 -475
rect 18005 -525 18010 -505
rect 18030 -525 18035 -505
rect 18005 -535 18035 -525
rect 18065 -455 18095 -370
rect 18065 -475 18070 -455
rect 18090 -475 18095 -455
rect 18065 -505 18095 -475
rect 18065 -525 18070 -505
rect 18090 -525 18095 -505
rect 18065 -535 18095 -525
rect 18125 -455 18155 -445
rect 18125 -475 18130 -455
rect 18150 -475 18155 -455
rect 18125 -505 18155 -475
rect 18125 -525 18130 -505
rect 18150 -525 18155 -505
rect 18035 -565 18065 -555
rect 18035 -585 18040 -565
rect 18060 -585 18065 -565
rect 18035 -615 18065 -585
rect 18125 -615 18155 -525
rect 18185 -455 18215 -370
rect 18185 -475 18190 -455
rect 18210 -475 18215 -455
rect 18185 -505 18215 -475
rect 18185 -525 18190 -505
rect 18210 -525 18215 -505
rect 18185 -535 18215 -525
rect 18245 -455 18275 -445
rect 18245 -475 18250 -455
rect 18270 -475 18275 -455
rect 18245 -505 18275 -475
rect 18245 -525 18250 -505
rect 18270 -525 18275 -505
rect 18245 -555 18275 -525
rect 18305 -455 18335 -370
rect 18360 -390 18400 -385
rect 18360 -420 18365 -390
rect 18395 -420 18400 -390
rect 18360 -425 18400 -420
rect 18305 -475 18310 -455
rect 18330 -475 18335 -455
rect 18305 -505 18335 -475
rect 18305 -525 18310 -505
rect 18330 -525 18335 -505
rect 18305 -535 18335 -525
rect 18365 -455 18395 -425
rect 18365 -475 18370 -455
rect 18390 -475 18395 -455
rect 18365 -505 18395 -475
rect 18365 -525 18370 -505
rect 18390 -525 18395 -505
rect 18365 -535 18395 -525
rect 18425 -455 18455 -370
rect 18425 -475 18430 -455
rect 18450 -475 18455 -455
rect 18425 -505 18455 -475
rect 18425 -525 18430 -505
rect 18450 -525 18455 -505
rect 18425 -535 18455 -525
rect 18485 -455 18515 -445
rect 18485 -475 18490 -455
rect 18510 -475 18515 -455
rect 18485 -505 18515 -475
rect 18485 -525 18490 -505
rect 18510 -525 18515 -505
rect 18240 -560 18280 -555
rect 18240 -590 18245 -560
rect 18275 -590 18280 -560
rect 18240 -595 18280 -590
rect 18365 -565 18395 -555
rect 18365 -585 18370 -565
rect 18390 -585 18395 -565
rect 18365 -615 18395 -585
rect 18485 -615 18515 -525
rect 18545 -455 18575 -370
rect 18545 -475 18550 -455
rect 18570 -475 18575 -455
rect 18545 -505 18575 -475
rect 18545 -525 18550 -505
rect 18570 -525 18575 -505
rect 18545 -535 18575 -525
rect 18605 -455 18635 -445
rect 18605 -475 18610 -455
rect 18630 -475 18635 -455
rect 18605 -505 18635 -475
rect 18605 -525 18610 -505
rect 18630 -525 18635 -505
rect 18605 -555 18635 -525
rect 18665 -455 18695 -370
rect 18720 -390 18760 -385
rect 18720 -420 18725 -390
rect 18755 -420 18760 -390
rect 18720 -425 18760 -420
rect 18665 -475 18670 -455
rect 18690 -475 18695 -455
rect 18665 -505 18695 -475
rect 18665 -525 18670 -505
rect 18690 -525 18695 -505
rect 18665 -535 18695 -525
rect 18725 -455 18755 -425
rect 18725 -475 18730 -455
rect 18750 -475 18755 -455
rect 18725 -505 18755 -475
rect 18725 -525 18730 -505
rect 18750 -525 18755 -505
rect 18725 -535 18755 -525
rect 18785 -455 18815 -370
rect 18785 -475 18790 -455
rect 18810 -475 18815 -455
rect 18785 -505 18815 -475
rect 18785 -525 18790 -505
rect 18810 -525 18815 -505
rect 18785 -535 18815 -525
rect 18845 -455 18875 -445
rect 18845 -475 18850 -455
rect 18870 -475 18875 -455
rect 18845 -505 18875 -475
rect 18845 -525 18850 -505
rect 18870 -525 18875 -505
rect 18600 -560 18640 -555
rect 18600 -590 18605 -560
rect 18635 -590 18640 -560
rect 18600 -595 18640 -590
rect 18725 -565 18755 -555
rect 18725 -585 18730 -565
rect 18750 -585 18755 -565
rect 18030 -620 18070 -615
rect 18030 -650 18035 -620
rect 18065 -650 18070 -620
rect 18030 -655 18070 -650
rect 18120 -620 18160 -615
rect 18120 -650 18125 -620
rect 18155 -650 18160 -620
rect 18120 -655 18160 -650
rect 18360 -620 18400 -615
rect 18360 -650 18365 -620
rect 18395 -650 18400 -620
rect 18360 -655 18400 -650
rect 18480 -620 18520 -615
rect 18480 -650 18485 -620
rect 18515 -650 18520 -620
rect 18480 -655 18520 -650
rect 18000 -815 18040 -810
rect 18000 -845 18005 -815
rect 18035 -845 18040 -815
rect 18000 -855 18040 -845
rect 18000 -885 18005 -855
rect 18035 -885 18040 -855
rect 18000 -895 18040 -885
rect 18000 -925 18005 -895
rect 18035 -925 18040 -895
rect 18000 -930 18040 -925
rect 18485 -820 18515 -655
rect 18563 -755 18593 -750
rect 18563 -790 18593 -785
rect 18610 -810 18630 -595
rect 18725 -615 18755 -585
rect 18845 -615 18875 -525
rect 18905 -455 18935 -370
rect 18905 -475 18910 -455
rect 18930 -475 18935 -455
rect 18905 -505 18935 -475
rect 18905 -525 18910 -505
rect 18930 -525 18935 -505
rect 18905 -535 18935 -525
rect 18965 -455 18995 -445
rect 18965 -475 18970 -455
rect 18990 -475 18995 -455
rect 18965 -505 18995 -475
rect 18965 -525 18970 -505
rect 18990 -525 18995 -505
rect 18965 -555 18995 -525
rect 19025 -455 19055 -370
rect 19080 -390 19120 -385
rect 19080 -420 19085 -390
rect 19115 -420 19120 -390
rect 19080 -425 19120 -420
rect 19145 -395 19175 -370
rect 19145 -415 19150 -395
rect 19170 -415 19175 -395
rect 19025 -475 19030 -455
rect 19050 -475 19055 -455
rect 19025 -505 19055 -475
rect 19025 -525 19030 -505
rect 19050 -525 19055 -505
rect 19025 -535 19055 -525
rect 19085 -455 19115 -425
rect 19085 -475 19090 -455
rect 19110 -475 19115 -455
rect 19085 -505 19115 -475
rect 19085 -525 19090 -505
rect 19110 -525 19115 -505
rect 19085 -535 19115 -525
rect 19145 -455 19175 -415
rect 19145 -475 19150 -455
rect 19170 -475 19175 -455
rect 19145 -505 19175 -475
rect 19145 -525 19150 -505
rect 19170 -525 19175 -505
rect 19145 -535 19175 -525
rect 18960 -560 19000 -555
rect 18960 -590 18965 -560
rect 18995 -590 19000 -560
rect 18960 -595 19000 -590
rect 19055 -570 19085 -560
rect 19055 -590 19060 -570
rect 19080 -590 19085 -570
rect 19055 -615 19085 -590
rect 18720 -620 18760 -615
rect 18720 -650 18725 -620
rect 18755 -650 18760 -620
rect 18720 -655 18760 -650
rect 18840 -620 18880 -615
rect 18840 -650 18845 -620
rect 18875 -650 18880 -620
rect 18840 -655 18880 -650
rect 19050 -620 19130 -615
rect 19050 -650 19055 -620
rect 19085 -650 19095 -620
rect 19125 -650 19130 -620
rect 19050 -655 19130 -650
rect 18485 -840 18490 -820
rect 18510 -840 18515 -820
rect 18485 -870 18515 -840
rect 18485 -890 18490 -870
rect 18510 -890 18515 -870
rect 18485 -920 18515 -890
rect 18485 -940 18490 -920
rect 18510 -940 18515 -920
rect 18485 -970 18515 -940
rect 18485 -990 18490 -970
rect 18510 -990 18515 -970
rect 18485 -1020 18515 -990
rect 18485 -1040 18490 -1020
rect 18510 -1040 18515 -1020
rect 18485 -1050 18515 -1040
rect 18545 -820 18575 -810
rect 18545 -840 18550 -820
rect 18570 -840 18575 -820
rect 18545 -870 18575 -840
rect 18545 -890 18550 -870
rect 18570 -890 18575 -870
rect 18545 -920 18575 -890
rect 18545 -940 18550 -920
rect 18570 -940 18575 -920
rect 18545 -970 18575 -940
rect 18545 -990 18550 -970
rect 18570 -990 18575 -970
rect 18545 -1020 18575 -990
rect 18545 -1040 18550 -1020
rect 18570 -1040 18575 -1020
rect 18440 -1075 18470 -1070
rect 18440 -1110 18470 -1105
rect 18545 -1125 18575 -1040
rect 18605 -820 18635 -810
rect 18605 -840 18610 -820
rect 18630 -840 18635 -820
rect 18605 -870 18635 -840
rect 18605 -890 18610 -870
rect 18630 -890 18635 -870
rect 18605 -920 18635 -890
rect 18605 -940 18610 -920
rect 18630 -940 18635 -920
rect 18605 -970 18635 -940
rect 18605 -990 18610 -970
rect 18630 -990 18635 -970
rect 18605 -1020 18635 -990
rect 18605 -1040 18610 -1020
rect 18630 -1040 18635 -1020
rect 18605 -1050 18635 -1040
rect 18540 -1130 18580 -1125
rect 18540 -1160 18545 -1130
rect 18575 -1160 18580 -1130
rect 18540 -1165 18580 -1160
rect 19030 -1130 19070 -1125
rect 19030 -1160 19035 -1130
rect 19065 -1160 19070 -1130
rect 19030 -1165 19070 -1160
rect 17875 -1305 17880 -1285
rect 17900 -1305 17905 -1285
rect 18020 -1185 18060 -1180
rect 18020 -1215 18025 -1185
rect 18055 -1215 18060 -1185
rect 18020 -1225 18060 -1215
rect 18020 -1255 18025 -1225
rect 18055 -1255 18060 -1225
rect 18020 -1265 18060 -1255
rect 18020 -1295 18025 -1265
rect 18055 -1295 18060 -1265
rect 18020 -1300 18060 -1295
rect 18140 -1185 18180 -1180
rect 18140 -1215 18145 -1185
rect 18175 -1215 18180 -1185
rect 18140 -1225 18180 -1215
rect 18140 -1255 18145 -1225
rect 18175 -1255 18180 -1225
rect 18140 -1265 18180 -1255
rect 18140 -1295 18145 -1265
rect 18175 -1295 18180 -1265
rect 18140 -1300 18180 -1295
rect 18260 -1185 18300 -1180
rect 18260 -1215 18265 -1185
rect 18295 -1215 18300 -1185
rect 18260 -1225 18300 -1215
rect 18260 -1255 18265 -1225
rect 18295 -1255 18300 -1225
rect 18260 -1265 18300 -1255
rect 18260 -1295 18265 -1265
rect 18295 -1295 18300 -1265
rect 18260 -1300 18300 -1295
rect 18580 -1185 18620 -1180
rect 18580 -1215 18585 -1185
rect 18615 -1215 18620 -1185
rect 18580 -1225 18620 -1215
rect 18580 -1255 18585 -1225
rect 18615 -1255 18620 -1225
rect 18580 -1265 18620 -1255
rect 18580 -1295 18585 -1265
rect 18615 -1295 18620 -1265
rect 18580 -1300 18620 -1295
rect 18700 -1185 18740 -1180
rect 18700 -1215 18705 -1185
rect 18735 -1215 18740 -1185
rect 18700 -1225 18740 -1215
rect 18700 -1255 18705 -1225
rect 18735 -1255 18740 -1225
rect 18700 -1265 18740 -1255
rect 18700 -1295 18705 -1265
rect 18735 -1295 18740 -1265
rect 18700 -1300 18740 -1295
rect 18820 -1185 18860 -1180
rect 18820 -1215 18825 -1185
rect 18855 -1215 18860 -1185
rect 18820 -1225 18860 -1215
rect 18820 -1255 18825 -1225
rect 18855 -1255 18860 -1225
rect 18820 -1265 18860 -1255
rect 18820 -1295 18825 -1265
rect 18855 -1295 18860 -1265
rect 18820 -1300 18860 -1295
rect 18940 -1185 18980 -1180
rect 18940 -1215 18945 -1185
rect 18975 -1215 18980 -1185
rect 18940 -1225 18980 -1215
rect 18940 -1255 18945 -1225
rect 18975 -1255 18980 -1225
rect 18940 -1265 18980 -1255
rect 18940 -1295 18945 -1265
rect 18975 -1295 18980 -1265
rect 19040 -1280 19060 -1165
rect 18940 -1300 18980 -1295
rect 19030 -1290 19070 -1280
rect 17875 -1315 17905 -1305
rect 19030 -1310 19040 -1290
rect 19060 -1310 19070 -1290
rect 19030 -1320 19070 -1310
rect 17740 -1615 17745 -1585
rect 17775 -1615 17785 -1585
rect 17815 -1615 17825 -1585
rect 17855 -1615 17860 -1585
rect 17740 -1625 17860 -1615
rect 17740 -1655 17745 -1625
rect 17775 -1655 17785 -1625
rect 17815 -1655 17825 -1625
rect 17855 -1655 17860 -1625
rect 17740 -1665 17860 -1655
rect 17740 -1695 17745 -1665
rect 17775 -1695 17785 -1665
rect 17815 -1695 17825 -1665
rect 17855 -1695 17860 -1665
rect 17740 -1700 17860 -1695
rect 18450 -1585 18490 -1580
rect 18450 -1615 18455 -1585
rect 18485 -1615 18490 -1585
rect 18450 -1625 18490 -1615
rect 18450 -1655 18455 -1625
rect 18485 -1655 18490 -1625
rect 18450 -1665 18490 -1655
rect 18450 -1695 18455 -1665
rect 18485 -1695 18490 -1665
rect 18450 -1700 18490 -1695
rect 16740 -1720 16780 -1715
rect 16740 -1750 16745 -1720
rect 16775 -1750 16780 -1720
rect 16740 -1755 16780 -1750
rect 16820 -1720 16860 -1715
rect 16820 -1750 16825 -1720
rect 16855 -1750 16860 -1720
rect 16820 -1755 16860 -1750
rect 16900 -1720 16940 -1715
rect 16900 -1750 16905 -1720
rect 16935 -1750 16940 -1720
rect 16900 -1755 16940 -1750
rect 16980 -1720 17020 -1715
rect 16980 -1750 16985 -1720
rect 17015 -1750 17020 -1720
rect 16980 -1755 17020 -1750
rect 17060 -1720 17100 -1715
rect 17060 -1750 17065 -1720
rect 17095 -1750 17100 -1720
rect 17060 -1755 17100 -1750
rect 17140 -1720 17180 -1715
rect 17140 -1750 17145 -1720
rect 17175 -1750 17180 -1720
rect 17140 -1755 17180 -1750
rect 17220 -1720 17260 -1715
rect 17220 -1750 17225 -1720
rect 17255 -1750 17260 -1720
rect 17220 -1755 17260 -1750
rect 17300 -1720 17340 -1715
rect 17300 -1750 17305 -1720
rect 17335 -1750 17340 -1720
rect 17300 -1755 17340 -1750
rect 17380 -1720 17420 -1715
rect 17380 -1750 17385 -1720
rect 17415 -1750 17420 -1720
rect 17380 -1755 17420 -1750
rect 17460 -1720 17500 -1715
rect 17460 -1750 17465 -1720
rect 17495 -1750 17500 -1720
rect 17460 -1755 17500 -1750
rect 17540 -1720 17580 -1715
rect 17540 -1750 17545 -1720
rect 17575 -1750 17580 -1720
rect 17540 -1755 17580 -1750
rect 17620 -1720 17660 -1715
rect 17620 -1750 17625 -1720
rect 17655 -1750 17660 -1720
rect 17620 -1755 17660 -1750
rect 17700 -1720 17740 -1715
rect 17700 -1750 17705 -1720
rect 17735 -1750 17740 -1720
rect 17700 -1755 17740 -1750
rect 17780 -1720 17820 -1715
rect 17780 -1750 17785 -1720
rect 17815 -1750 17820 -1720
rect 17780 -1755 17820 -1750
rect 17860 -1720 17900 -1715
rect 17860 -1750 17865 -1720
rect 17895 -1750 17900 -1720
rect 17860 -1755 17900 -1750
rect 17940 -1720 17980 -1715
rect 17940 -1750 17945 -1720
rect 17975 -1750 17980 -1720
rect 17940 -1755 17980 -1750
rect 18020 -1720 18060 -1715
rect 18020 -1750 18025 -1720
rect 18055 -1750 18060 -1720
rect 18020 -1755 18060 -1750
rect 18100 -1720 18140 -1715
rect 18100 -1750 18105 -1720
rect 18135 -1750 18140 -1720
rect 18100 -1755 18140 -1750
rect 18180 -1720 18220 -1715
rect 18180 -1750 18185 -1720
rect 18215 -1750 18220 -1720
rect 18180 -1755 18220 -1750
rect 18260 -1720 18300 -1715
rect 18260 -1750 18265 -1720
rect 18295 -1750 18300 -1720
rect 18260 -1755 18300 -1750
rect 18340 -1720 18380 -1715
rect 18340 -1750 18345 -1720
rect 18375 -1750 18380 -1720
rect 18340 -1755 18380 -1750
rect 18420 -1720 18460 -1715
rect 18420 -1750 18425 -1720
rect 18455 -1750 18460 -1720
rect 18420 -1755 18460 -1750
rect 18500 -1720 18540 -1715
rect 18500 -1750 18505 -1720
rect 18535 -1750 18540 -1720
rect 18500 -1755 18540 -1750
rect 18580 -1720 18620 -1715
rect 18580 -1750 18585 -1720
rect 18615 -1750 18620 -1720
rect 18580 -1755 18620 -1750
rect 18660 -1720 18700 -1715
rect 18660 -1750 18665 -1720
rect 18695 -1750 18700 -1720
rect 18660 -1755 18700 -1750
rect 18740 -1720 18780 -1715
rect 18740 -1750 18745 -1720
rect 18775 -1750 18780 -1720
rect 18740 -1755 18780 -1750
rect 18895 -1785 18935 -1780
rect 16700 -1805 16740 -1800
rect 16700 -1835 16705 -1805
rect 16735 -1835 16740 -1805
rect 16700 -1840 16740 -1835
rect 18895 -1815 18900 -1785
rect 18930 -1815 18935 -1785
rect 18895 -1825 18935 -1815
rect 18895 -1855 18900 -1825
rect 18930 -1855 18935 -1825
rect 18895 -1860 18935 -1855
rect 18885 -1890 18925 -1885
rect 18885 -1920 18890 -1890
rect 18920 -1920 18925 -1890
rect 16315 -2000 16355 -1995
rect 16315 -2030 16320 -2000
rect 16350 -2030 16355 -2000
rect 16315 -2035 16355 -2030
rect 17425 -2035 17430 -2000
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2035 18169 -2000
rect 18830 -2005 18870 -2000
rect 18830 -2035 18835 -2005
rect 18865 -2035 18870 -2005
rect 17425 -2060 17465 -2035
rect 17425 -2090 17430 -2060
rect 17460 -2090 17465 -2060
rect 17425 -2095 17465 -2090
rect 16260 -2100 16300 -2095
rect 16260 -2130 16265 -2100
rect 16295 -2130 16300 -2100
rect 16260 -2135 16300 -2130
rect 16480 -2100 16520 -2095
rect 16480 -2130 16485 -2100
rect 16515 -2130 16520 -2100
rect 16480 -2135 16520 -2130
rect 16730 -2100 16770 -2095
rect 16730 -2130 16735 -2100
rect 16765 -2130 16770 -2100
rect 16730 -2135 16770 -2130
rect 16490 -2895 16510 -2135
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16740 -3100 16760 -2135
rect 16945 -2615 18655 -2265
rect 16730 -3105 16770 -3100
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 16210 -3325 16245 -3320
rect 16210 -3365 16245 -3360
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -2035
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 16040 -4330 16045 -4300
rect 16075 -4330 16080 -4300
rect 16040 -4335 16080 -4330
rect 16100 -3894 16135 -3889
rect 16210 -3894 16245 -3889
rect 15905 -4400 15910 -4370
rect 15940 -4400 15950 -4370
rect 15980 -4400 15990 -4370
rect 16020 -4400 16025 -4370
rect 15905 -4410 16025 -4400
rect 15905 -4440 15910 -4410
rect 15940 -4440 15950 -4410
rect 15980 -4440 15990 -4410
rect 16020 -4440 16025 -4410
rect 15905 -4450 16025 -4440
rect 15905 -4480 15910 -4450
rect 15940 -4480 15950 -4450
rect 15980 -4480 15990 -4450
rect 16020 -4480 16025 -4450
rect 15905 -4485 16025 -4480
rect 16100 -4505 16140 -3929
rect 16210 -4155 16245 -3929
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 16605 -4155 16640 -4004
rect 16210 -4160 16250 -4155
rect 16210 -4190 16215 -4160
rect 16245 -4190 16250 -4160
rect 16210 -4200 16250 -4190
rect 16210 -4230 16215 -4200
rect 16245 -4230 16250 -4200
rect 16210 -4240 16250 -4230
rect 16210 -4270 16215 -4240
rect 16245 -4270 16250 -4240
rect 16210 -4275 16250 -4270
rect 16605 -4160 16645 -4155
rect 16605 -4190 16610 -4160
rect 16640 -4190 16645 -4160
rect 16605 -4200 16645 -4190
rect 16605 -4230 16610 -4200
rect 16640 -4230 16645 -4200
rect 16605 -4240 16645 -4230
rect 16605 -4270 16610 -4240
rect 16640 -4270 16645 -4240
rect 16605 -4275 16645 -4270
rect 17780 -4160 17820 -4155
rect 17780 -4190 17785 -4160
rect 17815 -4190 17820 -4160
rect 17780 -4200 17820 -4190
rect 17780 -4230 17785 -4200
rect 17815 -4230 17820 -4200
rect 17780 -4240 17820 -4230
rect 17780 -4270 17785 -4240
rect 17815 -4270 17820 -4240
rect 17780 -4275 17820 -4270
rect 17250 -4300 17300 -4290
rect 17250 -4330 17260 -4300
rect 17290 -4330 17300 -4300
rect 17250 -4340 17300 -4330
rect 16900 -4360 16950 -4350
rect 16900 -4390 16910 -4360
rect 16940 -4390 16950 -4360
rect 16900 -4410 16950 -4390
rect 16900 -4440 16910 -4410
rect 16940 -4440 16950 -4410
rect 16900 -4460 16950 -4440
rect 16900 -4490 16910 -4460
rect 16940 -4490 16950 -4460
rect 18650 -4450 18700 -4440
rect 18650 -4480 18660 -4450
rect 18690 -4480 18700 -4450
rect 18650 -4490 18700 -4480
rect 18885 -4450 18925 -1920
rect 19090 -1890 19130 -655
rect 19090 -1920 19095 -1890
rect 19125 -1920 19130 -1890
rect 19090 -1925 19130 -1920
rect 19225 -1075 19265 715
rect 19465 520 19505 525
rect 19465 490 19470 520
rect 19500 490 19505 520
rect 19225 -1105 19230 -1075
rect 19260 -1105 19265 -1075
rect 19225 -1945 19265 -1105
rect 19225 -1975 19230 -1945
rect 19260 -1975 19265 -1945
rect 19225 -1980 19265 -1975
rect 19305 -200 19345 -195
rect 19305 -230 19310 -200
rect 19340 -230 19345 -200
rect 19305 -755 19345 -230
rect 19305 -785 19310 -755
rect 19340 -785 19345 -755
rect 19080 -2060 19120 -2055
rect 19080 -2090 19085 -2060
rect 19115 -2090 19120 -2060
rect 19080 -2895 19120 -2090
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19305 -3088 19345 -785
rect 19465 -390 19505 490
rect 19465 -420 19470 -390
rect 19500 -420 19505 -390
rect 19305 -3090 19340 -3088
rect 19305 -3130 19340 -3125
rect 19465 -3115 19505 -420
rect 19465 -3160 19500 -3150
rect 19465 -3789 19500 -3784
rect 19185 -3894 19220 -3889
rect 18960 -3969 18995 -3964
rect 18960 -4005 18995 -4004
rect 18955 -4160 18995 -4005
rect 18955 -4190 18960 -4160
rect 18990 -4190 18995 -4160
rect 18955 -4200 18995 -4190
rect 18955 -4230 18960 -4200
rect 18990 -4230 18995 -4200
rect 18955 -4240 18995 -4230
rect 18955 -4270 18960 -4240
rect 18990 -4270 18995 -4240
rect 18955 -4275 18995 -4270
rect 19180 -4160 19220 -3929
rect 19180 -4190 19185 -4160
rect 19215 -4190 19220 -4160
rect 19180 -4200 19220 -4190
rect 19180 -4230 19185 -4200
rect 19215 -4230 19220 -4200
rect 19180 -4240 19220 -4230
rect 19180 -4270 19185 -4240
rect 19215 -4270 19220 -4240
rect 19180 -4275 19220 -4270
rect 18885 -4480 18890 -4450
rect 18920 -4480 18925 -4450
rect 18885 -4485 18925 -4480
rect 19355 -4450 19395 -4445
rect 19355 -4480 19360 -4450
rect 19390 -4480 19395 -4450
rect 19355 -4485 19395 -4480
rect 19465 -4450 19505 -3824
rect 19465 -4480 19470 -4450
rect 19500 -4480 19505 -4450
rect 19465 -4485 19505 -4480
rect 16900 -4500 16950 -4490
rect 16100 -4535 16105 -4505
rect 16135 -4535 16140 -4505
rect 16100 -4540 16140 -4535
rect 16205 -4505 16245 -4500
rect 16205 -4535 16210 -4505
rect 16240 -4535 16245 -4505
rect 16205 -4540 16245 -4535
rect 17955 -4560 17995 -4555
rect 17955 -4590 17960 -4560
rect 17990 -4590 17995 -4560
rect 17955 -4595 17995 -4590
<< via1 >>
rect 17035 715 17065 745
rect 17145 715 17175 745
rect 17255 715 17285 745
rect 17365 715 17395 745
rect 17475 715 17505 745
rect 17585 715 17615 745
rect 17985 715 18015 745
rect 18095 715 18125 745
rect 18205 715 18235 745
rect 18315 715 18345 745
rect 18425 715 18455 745
rect 18535 715 18565 745
rect 19230 715 19260 745
rect 16980 685 17010 690
rect 16980 665 16985 685
rect 16985 665 17005 685
rect 17005 665 17010 685
rect 16980 660 17010 665
rect 17090 660 17120 690
rect 17200 660 17230 690
rect 17310 660 17340 690
rect 17420 660 17450 690
rect 17530 660 17560 690
rect 17640 685 17670 690
rect 17640 665 17645 685
rect 17645 665 17665 685
rect 17665 665 17670 685
rect 17640 660 17670 665
rect 17930 685 17960 690
rect 17930 665 17935 685
rect 17935 665 17955 685
rect 17955 665 17960 685
rect 17930 660 17960 665
rect 18040 660 18070 690
rect 18150 660 18180 690
rect 18260 660 18290 690
rect 18370 660 18400 690
rect 18480 660 18510 690
rect 18590 685 18620 690
rect 18590 665 18595 685
rect 18595 665 18615 685
rect 18615 665 18620 685
rect 18590 660 18620 665
rect 17065 516 17091 521
rect 17065 499 17069 516
rect 17069 499 17086 516
rect 17086 499 17091 516
rect 17065 495 17091 499
rect 17120 516 17146 521
rect 17120 499 17124 516
rect 17124 499 17141 516
rect 17141 499 17146 516
rect 17120 495 17146 499
rect 17175 516 17201 521
rect 17175 499 17179 516
rect 17179 499 17196 516
rect 17196 499 17201 516
rect 17175 495 17201 499
rect 17230 516 17256 521
rect 17230 499 17234 516
rect 17234 499 17251 516
rect 17251 499 17256 516
rect 17230 495 17256 499
rect 17285 516 17311 521
rect 17285 499 17289 516
rect 17289 499 17306 516
rect 17306 499 17311 516
rect 17285 495 17311 499
rect 17340 516 17366 521
rect 17340 499 17344 516
rect 17344 499 17361 516
rect 17361 499 17366 516
rect 17340 495 17366 499
rect 17395 516 17421 521
rect 17395 499 17399 516
rect 17399 499 17416 516
rect 17416 499 17421 516
rect 17395 495 17421 499
rect 17450 516 17476 521
rect 17450 499 17454 516
rect 17454 499 17471 516
rect 17471 499 17476 516
rect 17450 495 17476 499
rect 17505 516 17531 521
rect 17505 499 17509 516
rect 17509 499 17526 516
rect 17526 499 17531 516
rect 17505 495 17531 499
rect 17560 516 17586 521
rect 17560 499 17564 516
rect 17564 499 17581 516
rect 17581 499 17586 516
rect 17560 495 17586 499
rect 18015 516 18041 521
rect 18015 499 18019 516
rect 18019 499 18036 516
rect 18036 499 18041 516
rect 18015 495 18041 499
rect 18070 516 18096 521
rect 18070 499 18074 516
rect 18074 499 18091 516
rect 18091 499 18096 516
rect 18070 495 18096 499
rect 18125 516 18151 521
rect 18125 499 18129 516
rect 18129 499 18146 516
rect 18146 499 18151 516
rect 18125 495 18151 499
rect 18180 516 18206 521
rect 18180 499 18184 516
rect 18184 499 18201 516
rect 18201 499 18206 516
rect 18180 495 18206 499
rect 18235 516 18261 521
rect 18235 499 18239 516
rect 18239 499 18256 516
rect 18256 499 18261 516
rect 18235 495 18261 499
rect 18290 516 18316 521
rect 18290 499 18294 516
rect 18294 499 18311 516
rect 18311 499 18316 516
rect 18290 495 18316 499
rect 18345 516 18371 521
rect 18345 499 18349 516
rect 18349 499 18366 516
rect 18366 499 18371 516
rect 18345 495 18371 499
rect 18400 516 18426 521
rect 18400 499 18404 516
rect 18404 499 18421 516
rect 18421 499 18426 516
rect 18400 495 18426 499
rect 18455 516 18481 521
rect 18455 499 18459 516
rect 18459 499 18476 516
rect 18476 499 18481 516
rect 18455 495 18481 499
rect 18510 516 18536 521
rect 18510 499 18514 516
rect 18514 499 18531 516
rect 18531 499 18536 516
rect 18510 495 18536 499
rect 16440 440 16470 470
rect 16440 400 16470 430
rect 16440 360 16470 390
rect 16660 440 16690 470
rect 16660 400 16690 430
rect 16660 360 16690 390
rect 16975 440 17005 470
rect 16975 400 17005 430
rect 16975 385 17005 390
rect 16975 365 16980 385
rect 16980 365 17000 385
rect 17000 365 17005 385
rect 16975 360 17005 365
rect 17155 440 17185 470
rect 17155 400 17185 430
rect 17155 385 17185 390
rect 17155 365 17160 385
rect 17160 365 17180 385
rect 17180 365 17185 385
rect 17155 360 17185 365
rect 17335 440 17365 470
rect 17335 400 17365 430
rect 17335 385 17365 390
rect 17335 365 17340 385
rect 17340 365 17360 385
rect 17360 365 17365 385
rect 17335 360 17365 365
rect 17515 440 17545 470
rect 17515 400 17545 430
rect 17515 385 17545 390
rect 17515 365 17520 385
rect 17520 365 17540 385
rect 17540 365 17545 385
rect 17515 360 17545 365
rect 17695 440 17725 470
rect 17695 400 17725 430
rect 17695 385 17725 390
rect 17695 365 17700 385
rect 17700 365 17720 385
rect 17720 365 17725 385
rect 17695 360 17725 365
rect 17875 440 17905 470
rect 17875 400 17905 430
rect 17875 385 17905 390
rect 17875 365 17880 385
rect 17880 365 17900 385
rect 17900 365 17905 385
rect 17875 360 17905 365
rect 18055 440 18085 470
rect 18055 400 18085 430
rect 18055 385 18085 390
rect 18055 365 18060 385
rect 18060 365 18080 385
rect 18080 365 18085 385
rect 18055 360 18085 365
rect 18235 440 18265 470
rect 18235 400 18265 430
rect 18235 385 18265 390
rect 18235 365 18240 385
rect 18240 365 18260 385
rect 18260 365 18265 385
rect 18235 360 18265 365
rect 18415 440 18445 470
rect 18415 400 18445 430
rect 18415 385 18445 390
rect 18415 365 18420 385
rect 18420 365 18440 385
rect 18440 365 18445 385
rect 18415 360 18445 365
rect 18595 440 18625 470
rect 18595 400 18625 430
rect 18595 385 18625 390
rect 18595 365 18600 385
rect 18600 365 18620 385
rect 18620 365 18625 385
rect 18595 360 18625 365
rect 16550 285 16580 290
rect 16550 265 16555 285
rect 16555 265 16575 285
rect 16575 265 16580 285
rect 16550 260 16580 265
rect 16785 260 16815 290
rect 16490 115 16520 120
rect 16490 95 16495 115
rect 16495 95 16515 115
rect 16515 95 16520 115
rect 16490 90 16520 95
rect 16610 115 16640 120
rect 16610 95 16615 115
rect 16615 95 16635 115
rect 16635 95 16640 115
rect 16610 90 16640 95
rect 16320 -65 16350 -35
rect 16265 -120 16295 -90
rect 16210 -175 16240 -145
rect 16100 -420 16130 -390
rect 15910 -650 15940 -620
rect 15950 -650 15980 -620
rect 15990 -650 16020 -620
rect 15910 -690 15940 -660
rect 15950 -690 15980 -660
rect 15990 -690 16020 -660
rect 15910 -730 15940 -700
rect 15950 -730 15980 -700
rect 15990 -730 16020 -700
rect 16265 -785 16295 -755
rect 16210 -1835 16240 -1805
rect 16045 -3250 16075 -3220
rect 16100 -3226 16135 -3221
rect 16100 -3251 16105 -3226
rect 16105 -3251 16130 -3226
rect 16130 -3251 16135 -3226
rect 16100 -3256 16135 -3251
rect 16210 -1975 16240 -1945
rect 16425 -285 16455 -255
rect 16425 -325 16455 -295
rect 16425 -365 16455 -335
rect 16785 -120 16815 -90
rect 16550 -175 16580 -145
rect 17110 15 17140 20
rect 17110 -5 17115 15
rect 17115 -5 17135 15
rect 17135 -5 17140 15
rect 17110 -10 17140 -5
rect 17200 15 17230 20
rect 17200 -5 17205 15
rect 17205 -5 17225 15
rect 17225 -5 17230 15
rect 17200 -10 17230 -5
rect 17290 15 17320 20
rect 17290 -5 17295 15
rect 17295 -5 17315 15
rect 17315 -5 17320 15
rect 17290 -10 17320 -5
rect 17380 15 17410 20
rect 17380 -5 17385 15
rect 17385 -5 17405 15
rect 17405 -5 17410 15
rect 17380 -10 17410 -5
rect 17470 15 17500 20
rect 17470 -5 17475 15
rect 17475 -5 17495 15
rect 17495 -5 17500 15
rect 17470 -10 17500 -5
rect 17560 15 17590 20
rect 17560 -5 17565 15
rect 17565 -5 17585 15
rect 17585 -5 17590 15
rect 17560 -10 17590 -5
rect 17650 15 17680 20
rect 17650 -5 17655 15
rect 17655 -5 17675 15
rect 17675 -5 17680 15
rect 17650 -10 17680 -5
rect 17695 -10 17725 20
rect 17740 15 17770 20
rect 17740 -5 17745 15
rect 17745 -5 17765 15
rect 17765 -5 17770 15
rect 17740 -10 17770 -5
rect 17605 -65 17635 -35
rect 17425 -120 17455 -90
rect 17245 -175 17275 -145
rect 17065 -230 17095 -200
rect 16545 -285 16575 -255
rect 16545 -325 16575 -295
rect 16545 -365 16575 -335
rect 16665 -285 16695 -255
rect 16665 -325 16695 -295
rect 16665 -365 16695 -335
rect 16785 -285 16815 -255
rect 16785 -325 16815 -295
rect 16785 -365 16815 -335
rect 16905 -285 16935 -255
rect 16905 -325 16935 -295
rect 16905 -365 16935 -335
rect 17025 -285 17055 -255
rect 17025 -325 17055 -295
rect 17025 -365 17055 -335
rect 17145 -285 17175 -255
rect 17145 -325 17175 -295
rect 17145 -365 17175 -335
rect 17265 -285 17295 -255
rect 17265 -325 17295 -295
rect 17265 -365 17295 -335
rect 17385 -285 17415 -255
rect 17385 -325 17415 -295
rect 17385 -365 17415 -335
rect 17505 -285 17535 -255
rect 17505 -325 17535 -295
rect 17505 -365 17535 -335
rect 17625 -285 17655 -255
rect 17625 -325 17655 -295
rect 17625 -365 17655 -335
rect 16485 -420 16515 -390
rect 16605 -565 16635 -560
rect 16605 -585 16610 -565
rect 16610 -585 16630 -565
rect 16630 -585 16635 -565
rect 16605 -590 16635 -585
rect 16845 -420 16875 -390
rect 16965 -565 16995 -560
rect 16965 -585 16970 -565
rect 16970 -585 16990 -565
rect 16990 -585 16995 -565
rect 16965 -590 16995 -585
rect 16515 -650 16545 -620
rect 16515 -690 16545 -660
rect 16515 -730 16545 -700
rect 16725 -650 16755 -620
rect 16725 -690 16755 -660
rect 16725 -730 16755 -700
rect 16845 -650 16875 -620
rect 16845 -690 16875 -660
rect 16845 -730 16875 -700
rect 17205 -420 17235 -390
rect 17325 -565 17355 -560
rect 17325 -585 17330 -565
rect 17330 -585 17350 -565
rect 17350 -585 17355 -565
rect 17325 -590 17355 -585
rect 17565 -420 17595 -390
rect 17830 15 17860 20
rect 17830 -5 17835 15
rect 17835 -5 17855 15
rect 17855 -5 17860 15
rect 17830 -10 17860 -5
rect 17920 15 17950 20
rect 17920 -5 17925 15
rect 17925 -5 17945 15
rect 17945 -5 17950 15
rect 17920 -10 17950 -5
rect 18010 15 18040 20
rect 18010 -5 18015 15
rect 18015 -5 18035 15
rect 18035 -5 18040 15
rect 18010 -10 18040 -5
rect 18100 15 18130 20
rect 18100 -5 18105 15
rect 18105 -5 18125 15
rect 18125 -5 18130 15
rect 18100 -10 18130 -5
rect 17965 -65 17995 -35
rect 18190 15 18220 20
rect 18190 -5 18195 15
rect 18195 -5 18215 15
rect 18215 -5 18220 15
rect 18190 -10 18220 -5
rect 18280 15 18310 20
rect 18280 -5 18285 15
rect 18285 -5 18305 15
rect 18305 -5 18310 15
rect 18280 -10 18310 -5
rect 18145 -120 18175 -90
rect 18370 15 18400 20
rect 18370 -5 18375 15
rect 18375 -5 18395 15
rect 18395 -5 18400 15
rect 18370 -10 18400 -5
rect 18460 15 18490 20
rect 18460 -5 18465 15
rect 18465 -5 18485 15
rect 18485 -5 18490 15
rect 18460 -10 18490 -5
rect 18325 -175 18355 -145
rect 17785 -230 17815 -200
rect 18505 -230 18535 -200
rect 17945 -285 17975 -255
rect 17945 -325 17975 -295
rect 17945 -365 17975 -335
rect 18065 -285 18095 -255
rect 18065 -325 18095 -295
rect 18065 -365 18095 -335
rect 18185 -285 18215 -255
rect 18185 -325 18215 -295
rect 18185 -365 18215 -335
rect 18305 -285 18335 -255
rect 18305 -325 18335 -295
rect 18305 -365 18335 -335
rect 18425 -285 18455 -255
rect 18425 -325 18455 -295
rect 18425 -365 18455 -335
rect 18545 -285 18575 -255
rect 18545 -325 18575 -295
rect 18545 -365 18575 -335
rect 18665 -285 18695 -255
rect 18665 -325 18695 -295
rect 18665 -365 18695 -335
rect 18785 -285 18815 -255
rect 18785 -325 18815 -295
rect 18785 -365 18815 -335
rect 18905 -285 18935 -255
rect 18905 -325 18935 -295
rect 18905 -365 18935 -335
rect 19025 -285 19055 -255
rect 19025 -325 19055 -295
rect 19025 -365 19055 -335
rect 19145 -285 19175 -255
rect 19145 -325 19175 -295
rect 19145 -365 19175 -335
rect 17695 -420 17725 -390
rect 17875 -420 17905 -390
rect 17085 -650 17115 -620
rect 17085 -690 17115 -660
rect 17085 -730 17115 -700
rect 17205 -650 17235 -620
rect 17205 -690 17235 -660
rect 17205 -730 17235 -700
rect 17445 -650 17475 -620
rect 17445 -690 17475 -660
rect 17445 -730 17475 -700
rect 17535 -650 17565 -620
rect 17535 -690 17565 -660
rect 17535 -730 17565 -700
rect 17007 -760 17037 -755
rect 17007 -780 17012 -760
rect 17012 -780 17032 -760
rect 17032 -780 17037 -760
rect 17007 -785 17037 -780
rect 16320 -1105 16350 -1075
rect 17565 -820 17595 -815
rect 17565 -840 17570 -820
rect 17570 -840 17590 -820
rect 17590 -840 17595 -820
rect 17565 -845 17595 -840
rect 17565 -860 17595 -855
rect 17565 -880 17570 -860
rect 17570 -880 17590 -860
rect 17590 -880 17595 -860
rect 17565 -885 17595 -880
rect 17565 -900 17595 -895
rect 17565 -920 17570 -900
rect 17570 -920 17590 -900
rect 17590 -920 17595 -900
rect 17565 -925 17595 -920
rect 17075 -1080 17105 -1075
rect 17075 -1100 17080 -1080
rect 17080 -1100 17100 -1080
rect 17100 -1100 17105 -1080
rect 17075 -1105 17105 -1100
rect 16535 -1160 16565 -1130
rect 17025 -1160 17055 -1130
rect 16625 -1215 16655 -1185
rect 16625 -1255 16655 -1225
rect 16625 -1270 16655 -1265
rect 16625 -1290 16630 -1270
rect 16630 -1290 16650 -1270
rect 16650 -1290 16655 -1270
rect 16625 -1295 16655 -1290
rect 16745 -1215 16775 -1185
rect 16745 -1255 16775 -1225
rect 16745 -1270 16775 -1265
rect 16745 -1290 16750 -1270
rect 16750 -1290 16770 -1270
rect 16770 -1290 16775 -1270
rect 16745 -1295 16775 -1290
rect 16865 -1215 16895 -1185
rect 16865 -1255 16895 -1225
rect 16865 -1270 16895 -1265
rect 16865 -1290 16870 -1270
rect 16870 -1290 16890 -1270
rect 16890 -1290 16895 -1270
rect 16865 -1295 16895 -1290
rect 16985 -1215 17015 -1185
rect 16985 -1255 17015 -1225
rect 16985 -1270 17015 -1265
rect 16985 -1290 16990 -1270
rect 16990 -1290 17010 -1270
rect 17010 -1290 17015 -1270
rect 16985 -1295 17015 -1290
rect 17305 -1215 17335 -1185
rect 17305 -1255 17335 -1225
rect 17305 -1270 17335 -1265
rect 17305 -1290 17310 -1270
rect 17310 -1290 17330 -1270
rect 17330 -1290 17335 -1270
rect 17305 -1295 17335 -1290
rect 17425 -1215 17455 -1185
rect 17425 -1255 17455 -1225
rect 17425 -1270 17455 -1265
rect 17425 -1290 17430 -1270
rect 17430 -1290 17450 -1270
rect 17450 -1290 17455 -1270
rect 17425 -1295 17455 -1290
rect 17545 -1215 17575 -1185
rect 17545 -1255 17575 -1225
rect 17545 -1270 17575 -1265
rect 17545 -1290 17550 -1270
rect 17550 -1290 17570 -1270
rect 17570 -1290 17575 -1270
rect 17545 -1295 17575 -1290
rect 17745 -845 17775 -815
rect 17785 -845 17815 -815
rect 17825 -845 17855 -815
rect 17745 -885 17775 -855
rect 17785 -885 17815 -855
rect 17825 -885 17855 -855
rect 17745 -925 17775 -895
rect 17785 -925 17815 -895
rect 17825 -925 17855 -895
rect 17115 -1590 17145 -1585
rect 17115 -1610 17120 -1590
rect 17120 -1610 17140 -1590
rect 17140 -1610 17145 -1590
rect 17115 -1615 17145 -1610
rect 17115 -1655 17145 -1625
rect 17115 -1695 17145 -1665
rect 18005 -420 18035 -390
rect 18365 -420 18395 -390
rect 18245 -565 18275 -560
rect 18245 -585 18250 -565
rect 18250 -585 18270 -565
rect 18270 -585 18275 -565
rect 18245 -590 18275 -585
rect 18725 -420 18755 -390
rect 18605 -565 18635 -560
rect 18605 -585 18610 -565
rect 18610 -585 18630 -565
rect 18630 -585 18635 -565
rect 18605 -590 18635 -585
rect 18035 -650 18065 -620
rect 18125 -650 18155 -620
rect 18365 -650 18395 -620
rect 18485 -650 18515 -620
rect 18005 -820 18035 -815
rect 18005 -840 18010 -820
rect 18010 -840 18030 -820
rect 18030 -840 18035 -820
rect 18005 -845 18035 -840
rect 18005 -860 18035 -855
rect 18005 -880 18010 -860
rect 18010 -880 18030 -860
rect 18030 -880 18035 -860
rect 18005 -885 18035 -880
rect 18005 -900 18035 -895
rect 18005 -920 18010 -900
rect 18010 -920 18030 -900
rect 18030 -920 18035 -900
rect 18005 -925 18035 -920
rect 18563 -760 18593 -755
rect 18563 -780 18568 -760
rect 18568 -780 18588 -760
rect 18588 -780 18593 -760
rect 18563 -785 18593 -780
rect 19085 -420 19115 -390
rect 18965 -565 18995 -560
rect 18965 -585 18970 -565
rect 18970 -585 18990 -565
rect 18990 -585 18995 -565
rect 18965 -590 18995 -585
rect 18725 -650 18755 -620
rect 18845 -650 18875 -620
rect 19055 -650 19085 -620
rect 19095 -650 19125 -620
rect 18440 -1080 18470 -1075
rect 18440 -1100 18445 -1080
rect 18445 -1100 18465 -1080
rect 18465 -1100 18470 -1080
rect 18440 -1105 18470 -1100
rect 18545 -1160 18575 -1130
rect 19035 -1160 19065 -1130
rect 18025 -1215 18055 -1185
rect 18025 -1255 18055 -1225
rect 18025 -1270 18055 -1265
rect 18025 -1290 18030 -1270
rect 18030 -1290 18050 -1270
rect 18050 -1290 18055 -1270
rect 18025 -1295 18055 -1290
rect 18145 -1215 18175 -1185
rect 18145 -1255 18175 -1225
rect 18145 -1270 18175 -1265
rect 18145 -1290 18150 -1270
rect 18150 -1290 18170 -1270
rect 18170 -1290 18175 -1270
rect 18145 -1295 18175 -1290
rect 18265 -1215 18295 -1185
rect 18265 -1255 18295 -1225
rect 18265 -1270 18295 -1265
rect 18265 -1290 18270 -1270
rect 18270 -1290 18290 -1270
rect 18290 -1290 18295 -1270
rect 18265 -1295 18295 -1290
rect 18585 -1215 18615 -1185
rect 18585 -1255 18615 -1225
rect 18585 -1270 18615 -1265
rect 18585 -1290 18590 -1270
rect 18590 -1290 18610 -1270
rect 18610 -1290 18615 -1270
rect 18585 -1295 18615 -1290
rect 18705 -1215 18735 -1185
rect 18705 -1255 18735 -1225
rect 18705 -1270 18735 -1265
rect 18705 -1290 18710 -1270
rect 18710 -1290 18730 -1270
rect 18730 -1290 18735 -1270
rect 18705 -1295 18735 -1290
rect 18825 -1215 18855 -1185
rect 18825 -1255 18855 -1225
rect 18825 -1270 18855 -1265
rect 18825 -1290 18830 -1270
rect 18830 -1290 18850 -1270
rect 18850 -1290 18855 -1270
rect 18825 -1295 18855 -1290
rect 18945 -1215 18975 -1185
rect 18945 -1255 18975 -1225
rect 18945 -1270 18975 -1265
rect 18945 -1290 18950 -1270
rect 18950 -1290 18970 -1270
rect 18970 -1290 18975 -1270
rect 18945 -1295 18975 -1290
rect 17745 -1615 17775 -1585
rect 17785 -1615 17815 -1585
rect 17825 -1615 17855 -1585
rect 17745 -1655 17775 -1625
rect 17785 -1655 17815 -1625
rect 17825 -1655 17855 -1625
rect 17745 -1695 17775 -1665
rect 17785 -1695 17815 -1665
rect 17825 -1695 17855 -1665
rect 18455 -1590 18485 -1585
rect 18455 -1610 18460 -1590
rect 18460 -1610 18480 -1590
rect 18480 -1610 18485 -1590
rect 18455 -1615 18485 -1610
rect 18455 -1655 18485 -1625
rect 18455 -1695 18485 -1665
rect 16745 -1725 16775 -1720
rect 16745 -1745 16750 -1725
rect 16750 -1745 16770 -1725
rect 16770 -1745 16775 -1725
rect 16745 -1750 16775 -1745
rect 16825 -1725 16855 -1720
rect 16825 -1745 16830 -1725
rect 16830 -1745 16850 -1725
rect 16850 -1745 16855 -1725
rect 16825 -1750 16855 -1745
rect 16905 -1725 16935 -1720
rect 16905 -1745 16910 -1725
rect 16910 -1745 16930 -1725
rect 16930 -1745 16935 -1725
rect 16905 -1750 16935 -1745
rect 16985 -1725 17015 -1720
rect 16985 -1745 16990 -1725
rect 16990 -1745 17010 -1725
rect 17010 -1745 17015 -1725
rect 16985 -1750 17015 -1745
rect 17065 -1725 17095 -1720
rect 17065 -1745 17070 -1725
rect 17070 -1745 17090 -1725
rect 17090 -1745 17095 -1725
rect 17065 -1750 17095 -1745
rect 17145 -1725 17175 -1720
rect 17145 -1745 17150 -1725
rect 17150 -1745 17170 -1725
rect 17170 -1745 17175 -1725
rect 17145 -1750 17175 -1745
rect 17225 -1725 17255 -1720
rect 17225 -1745 17230 -1725
rect 17230 -1745 17250 -1725
rect 17250 -1745 17255 -1725
rect 17225 -1750 17255 -1745
rect 17305 -1725 17335 -1720
rect 17305 -1745 17310 -1725
rect 17310 -1745 17330 -1725
rect 17330 -1745 17335 -1725
rect 17305 -1750 17335 -1745
rect 17385 -1725 17415 -1720
rect 17385 -1745 17390 -1725
rect 17390 -1745 17410 -1725
rect 17410 -1745 17415 -1725
rect 17385 -1750 17415 -1745
rect 17465 -1725 17495 -1720
rect 17465 -1745 17470 -1725
rect 17470 -1745 17490 -1725
rect 17490 -1745 17495 -1725
rect 17465 -1750 17495 -1745
rect 17545 -1725 17575 -1720
rect 17545 -1745 17550 -1725
rect 17550 -1745 17570 -1725
rect 17570 -1745 17575 -1725
rect 17545 -1750 17575 -1745
rect 17625 -1725 17655 -1720
rect 17625 -1745 17630 -1725
rect 17630 -1745 17650 -1725
rect 17650 -1745 17655 -1725
rect 17625 -1750 17655 -1745
rect 17705 -1725 17735 -1720
rect 17705 -1745 17710 -1725
rect 17710 -1745 17730 -1725
rect 17730 -1745 17735 -1725
rect 17705 -1750 17735 -1745
rect 17785 -1725 17815 -1720
rect 17785 -1745 17790 -1725
rect 17790 -1745 17810 -1725
rect 17810 -1745 17815 -1725
rect 17785 -1750 17815 -1745
rect 17865 -1725 17895 -1720
rect 17865 -1745 17870 -1725
rect 17870 -1745 17890 -1725
rect 17890 -1745 17895 -1725
rect 17865 -1750 17895 -1745
rect 17945 -1725 17975 -1720
rect 17945 -1745 17950 -1725
rect 17950 -1745 17970 -1725
rect 17970 -1745 17975 -1725
rect 17945 -1750 17975 -1745
rect 18025 -1725 18055 -1720
rect 18025 -1745 18030 -1725
rect 18030 -1745 18050 -1725
rect 18050 -1745 18055 -1725
rect 18025 -1750 18055 -1745
rect 18105 -1725 18135 -1720
rect 18105 -1745 18110 -1725
rect 18110 -1745 18130 -1725
rect 18130 -1745 18135 -1725
rect 18105 -1750 18135 -1745
rect 18185 -1725 18215 -1720
rect 18185 -1745 18190 -1725
rect 18190 -1745 18210 -1725
rect 18210 -1745 18215 -1725
rect 18185 -1750 18215 -1745
rect 18265 -1725 18295 -1720
rect 18265 -1745 18270 -1725
rect 18270 -1745 18290 -1725
rect 18290 -1745 18295 -1725
rect 18265 -1750 18295 -1745
rect 18345 -1725 18375 -1720
rect 18345 -1745 18350 -1725
rect 18350 -1745 18370 -1725
rect 18370 -1745 18375 -1725
rect 18345 -1750 18375 -1745
rect 18425 -1725 18455 -1720
rect 18425 -1745 18430 -1725
rect 18430 -1745 18450 -1725
rect 18450 -1745 18455 -1725
rect 18425 -1750 18455 -1745
rect 18505 -1725 18535 -1720
rect 18505 -1745 18510 -1725
rect 18510 -1745 18530 -1725
rect 18530 -1745 18535 -1725
rect 18505 -1750 18535 -1745
rect 18585 -1725 18615 -1720
rect 18585 -1745 18590 -1725
rect 18590 -1745 18610 -1725
rect 18610 -1745 18615 -1725
rect 18585 -1750 18615 -1745
rect 18665 -1725 18695 -1720
rect 18665 -1745 18670 -1725
rect 18670 -1745 18690 -1725
rect 18690 -1745 18695 -1725
rect 18665 -1750 18695 -1745
rect 18745 -1725 18775 -1720
rect 18745 -1745 18750 -1725
rect 18750 -1745 18770 -1725
rect 18770 -1745 18775 -1725
rect 18745 -1750 18775 -1745
rect 16705 -1810 16735 -1805
rect 16705 -1830 16710 -1810
rect 16710 -1830 16730 -1810
rect 16730 -1830 16735 -1810
rect 16705 -1835 16735 -1830
rect 18900 -1790 18930 -1785
rect 18900 -1810 18905 -1790
rect 18905 -1810 18925 -1790
rect 18925 -1810 18930 -1790
rect 18900 -1815 18930 -1810
rect 18900 -1830 18930 -1825
rect 18900 -1850 18905 -1830
rect 18905 -1850 18925 -1830
rect 18925 -1850 18930 -1830
rect 18900 -1855 18930 -1850
rect 18890 -1920 18920 -1890
rect 16320 -2030 16350 -2000
rect 17430 -2005 17465 -2000
rect 17430 -2030 17435 -2005
rect 17435 -2030 17460 -2005
rect 17460 -2030 17465 -2005
rect 17430 -2035 17465 -2030
rect 18129 -2005 18164 -2000
rect 18129 -2030 18134 -2005
rect 18134 -2030 18159 -2005
rect 18159 -2030 18164 -2005
rect 18129 -2035 18164 -2030
rect 18835 -2035 18865 -2005
rect 17430 -2090 17460 -2060
rect 16265 -2130 16295 -2100
rect 16485 -2130 16515 -2100
rect 16735 -2130 16765 -2100
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16735 -3135 16765 -3105
rect 16210 -3330 16245 -3325
rect 16210 -3355 16215 -3330
rect 16215 -3355 16240 -3330
rect 16240 -3355 16245 -3330
rect 16210 -3360 16245 -3355
rect 17785 -3135 17815 -3105
rect 18620 -3135 18650 -3105
rect 18835 -3135 18865 -3105
rect 16045 -4330 16075 -4300
rect 16100 -3899 16135 -3894
rect 16100 -3924 16105 -3899
rect 16105 -3924 16130 -3899
rect 16130 -3924 16135 -3899
rect 16100 -3929 16135 -3924
rect 16210 -3899 16245 -3894
rect 16210 -3924 16215 -3899
rect 16215 -3924 16240 -3899
rect 16240 -3924 16245 -3899
rect 16210 -3929 16245 -3924
rect 15910 -4400 15940 -4370
rect 15950 -4400 15980 -4370
rect 15990 -4400 16020 -4370
rect 15910 -4440 15940 -4410
rect 15950 -4440 15980 -4410
rect 15990 -4440 16020 -4410
rect 15910 -4480 15940 -4450
rect 15950 -4480 15980 -4450
rect 15990 -4480 16020 -4450
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4004 16640 -3999
rect 16215 -4190 16245 -4160
rect 16215 -4230 16245 -4200
rect 16215 -4270 16245 -4240
rect 16610 -4190 16640 -4160
rect 16610 -4230 16640 -4200
rect 16610 -4270 16640 -4240
rect 17785 -4165 17815 -4160
rect 17785 -4185 17790 -4165
rect 17790 -4185 17810 -4165
rect 17810 -4185 17815 -4165
rect 17785 -4190 17815 -4185
rect 17785 -4205 17815 -4200
rect 17785 -4225 17790 -4205
rect 17790 -4225 17810 -4205
rect 17810 -4225 17815 -4205
rect 17785 -4230 17815 -4225
rect 17785 -4245 17815 -4240
rect 17785 -4265 17790 -4245
rect 17790 -4265 17810 -4245
rect 17810 -4265 17815 -4245
rect 17785 -4270 17815 -4265
rect 17260 -4330 17290 -4300
rect 16910 -4390 16940 -4360
rect 16910 -4440 16940 -4410
rect 16910 -4490 16940 -4460
rect 18660 -4480 18690 -4450
rect 19095 -1920 19125 -1890
rect 19470 490 19500 520
rect 19230 -1105 19260 -1075
rect 19230 -1975 19260 -1945
rect 19310 -230 19340 -200
rect 19310 -785 19340 -755
rect 19085 -2090 19115 -2060
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19470 -420 19500 -390
rect 19305 -3095 19340 -3090
rect 19305 -3120 19310 -3095
rect 19310 -3120 19335 -3095
rect 19335 -3120 19340 -3095
rect 19305 -3125 19340 -3120
rect 19465 -3120 19500 -3115
rect 19465 -3145 19470 -3120
rect 19470 -3145 19495 -3120
rect 19495 -3145 19500 -3120
rect 19465 -3150 19500 -3145
rect 19465 -3794 19500 -3789
rect 19465 -3819 19470 -3794
rect 19470 -3819 19495 -3794
rect 19495 -3819 19500 -3794
rect 19465 -3824 19500 -3819
rect 19185 -3899 19220 -3894
rect 19185 -3924 19190 -3899
rect 19190 -3924 19215 -3899
rect 19215 -3924 19220 -3899
rect 19185 -3929 19220 -3924
rect 18960 -3974 18995 -3969
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 18960 -4190 18990 -4160
rect 18960 -4230 18990 -4200
rect 18960 -4270 18990 -4240
rect 19185 -4190 19215 -4160
rect 19185 -4230 19215 -4200
rect 19185 -4270 19215 -4240
rect 18890 -4480 18920 -4450
rect 19360 -4480 19390 -4450
rect 19470 -4480 19500 -4450
rect 16105 -4535 16135 -4505
rect 16210 -4535 16240 -4505
rect 17960 -4590 17990 -4560
<< metal2 >>
rect 17030 745 17620 750
rect 17030 715 17035 745
rect 17065 715 17145 745
rect 17175 715 17255 745
rect 17285 715 17365 745
rect 17395 715 17475 745
rect 17505 715 17585 745
rect 17615 715 17620 745
rect 17030 710 17620 715
rect 17980 745 19265 750
rect 17980 715 17985 745
rect 18015 715 18095 745
rect 18125 715 18205 745
rect 18235 715 18315 745
rect 18345 715 18425 745
rect 18455 715 18535 745
rect 18565 715 19230 745
rect 19260 715 19265 745
rect 17980 710 19265 715
rect 15510 690 18625 695
rect 15510 660 15515 690
rect 15545 660 15560 690
rect 15590 660 15605 690
rect 15635 660 16980 690
rect 17010 660 17090 690
rect 17120 660 17200 690
rect 17230 660 17310 690
rect 17340 660 17420 690
rect 17450 660 17530 690
rect 17560 660 17640 690
rect 17670 660 17930 690
rect 17960 660 18040 690
rect 18070 660 18150 690
rect 18180 660 18260 690
rect 18290 660 18370 690
rect 18400 660 18480 690
rect 18510 660 18590 690
rect 18620 660 18625 690
rect 15510 655 18625 660
rect 17063 521 19505 525
rect 17063 495 17065 521
rect 17091 495 17120 521
rect 17146 495 17175 521
rect 17201 495 17230 521
rect 17256 495 17285 521
rect 17311 495 17340 521
rect 17366 495 17395 521
rect 17421 495 17450 521
rect 17476 495 17505 521
rect 17531 495 17560 521
rect 17586 495 18015 521
rect 18041 495 18070 521
rect 18096 495 18125 521
rect 18151 495 18180 521
rect 18206 495 18235 521
rect 18261 495 18290 521
rect 18316 495 18345 521
rect 18371 495 18400 521
rect 18426 495 18455 521
rect 18481 495 18510 521
rect 18536 520 19505 521
rect 18536 495 19470 520
rect 17063 490 19470 495
rect 19500 490 19505 520
rect 15510 470 18630 475
rect 15510 440 15515 470
rect 15545 440 15560 470
rect 15590 440 15605 470
rect 15635 440 16440 470
rect 16470 440 16660 470
rect 16690 440 16975 470
rect 17005 440 17155 470
rect 17185 440 17335 470
rect 17365 440 17515 470
rect 17545 440 17695 470
rect 17725 440 17875 470
rect 17905 440 18055 470
rect 18085 440 18235 470
rect 18265 440 18415 470
rect 18445 440 18595 470
rect 18625 440 18630 470
rect 15510 430 18630 440
rect 15510 425 16440 430
rect 15510 395 15515 425
rect 15545 395 15560 425
rect 15590 395 15605 425
rect 15635 400 16440 425
rect 16470 400 16660 430
rect 16690 400 16975 430
rect 17005 400 17155 430
rect 17185 400 17335 430
rect 17365 400 17515 430
rect 17545 400 17695 430
rect 17725 400 17875 430
rect 17905 400 18055 430
rect 18085 400 18235 430
rect 18265 400 18415 430
rect 18445 400 18595 430
rect 18625 400 18630 430
rect 15635 395 18630 400
rect 15510 390 18630 395
rect 15510 380 16440 390
rect 15510 350 15515 380
rect 15545 350 15560 380
rect 15590 350 15605 380
rect 15635 360 16440 380
rect 16470 360 16660 390
rect 16690 360 16975 390
rect 17005 360 17155 390
rect 17185 360 17335 390
rect 17365 360 17515 390
rect 17545 360 17695 390
rect 17725 360 17875 390
rect 17905 360 18055 390
rect 18085 360 18235 390
rect 18265 360 18415 390
rect 18445 360 18595 390
rect 18625 360 18630 390
rect 15635 355 18630 360
rect 15635 350 15640 355
rect 15510 345 15640 350
rect 16545 290 16585 295
rect 16545 260 16550 290
rect 16580 285 16585 290
rect 16780 290 16820 295
rect 16780 285 16785 290
rect 16580 265 16785 285
rect 16580 260 16585 265
rect 16545 255 16585 260
rect 16780 260 16785 265
rect 16815 260 16820 290
rect 16780 255 16820 260
rect 16485 120 16645 125
rect 16485 90 16490 120
rect 16520 90 16610 120
rect 16640 90 16645 120
rect 16485 85 16645 90
rect 17110 20 18490 25
rect 17140 -10 17200 20
rect 17230 -10 17290 20
rect 17320 -10 17380 20
rect 17410 -10 17470 20
rect 17500 -10 17560 20
rect 17590 -10 17650 20
rect 17680 -10 17695 20
rect 17725 -10 17740 20
rect 17770 -10 17830 20
rect 17860 -10 17920 20
rect 17950 -10 18010 20
rect 18040 -10 18100 20
rect 18130 -10 18190 20
rect 18220 -10 18280 20
rect 18310 -10 18370 20
rect 18400 -10 18460 20
rect 17110 -15 18490 -10
rect 16315 -35 18000 -30
rect 16315 -65 16320 -35
rect 16350 -65 17605 -35
rect 17635 -65 17965 -35
rect 17995 -65 18000 -35
rect 16315 -70 18000 -65
rect 16260 -90 18180 -85
rect 16260 -120 16265 -90
rect 16295 -120 16785 -90
rect 16815 -120 17425 -90
rect 17455 -120 18145 -90
rect 18175 -120 18180 -90
rect 16260 -125 18180 -120
rect 16205 -145 18360 -140
rect 16205 -175 16210 -145
rect 16240 -175 16550 -145
rect 16580 -175 17245 -145
rect 17275 -175 18325 -145
rect 18355 -175 18360 -145
rect 16205 -180 18360 -175
rect 17060 -200 19345 -195
rect 17060 -230 17065 -200
rect 17095 -230 17785 -200
rect 17815 -230 18505 -200
rect 18535 -230 19310 -200
rect 19340 -230 19345 -200
rect 17060 -235 19345 -230
rect 15510 -255 19180 -250
rect 15510 -285 15515 -255
rect 15545 -285 15560 -255
rect 15590 -285 15605 -255
rect 15635 -285 16425 -255
rect 16455 -285 16545 -255
rect 16575 -285 16665 -255
rect 16695 -285 16785 -255
rect 16815 -285 16905 -255
rect 16935 -285 17025 -255
rect 17055 -285 17145 -255
rect 17175 -285 17265 -255
rect 17295 -285 17385 -255
rect 17415 -285 17505 -255
rect 17535 -285 17625 -255
rect 17655 -285 17945 -255
rect 17975 -285 18065 -255
rect 18095 -285 18185 -255
rect 18215 -285 18305 -255
rect 18335 -285 18425 -255
rect 18455 -285 18545 -255
rect 18575 -285 18665 -255
rect 18695 -285 18785 -255
rect 18815 -285 18905 -255
rect 18935 -285 19025 -255
rect 19055 -285 19145 -255
rect 19175 -285 19180 -255
rect 15510 -295 19180 -285
rect 15510 -300 16425 -295
rect 15510 -330 15515 -300
rect 15545 -330 15560 -300
rect 15590 -330 15605 -300
rect 15635 -325 16425 -300
rect 16455 -325 16545 -295
rect 16575 -325 16665 -295
rect 16695 -325 16785 -295
rect 16815 -325 16905 -295
rect 16935 -325 17025 -295
rect 17055 -325 17145 -295
rect 17175 -325 17265 -295
rect 17295 -325 17385 -295
rect 17415 -325 17505 -295
rect 17535 -325 17625 -295
rect 17655 -325 17945 -295
rect 17975 -325 18065 -295
rect 18095 -325 18185 -295
rect 18215 -325 18305 -295
rect 18335 -325 18425 -295
rect 18455 -325 18545 -295
rect 18575 -325 18665 -295
rect 18695 -325 18785 -295
rect 18815 -325 18905 -295
rect 18935 -325 19025 -295
rect 19055 -325 19145 -295
rect 19175 -325 19180 -295
rect 15635 -330 19180 -325
rect 15510 -335 19180 -330
rect 15510 -345 16425 -335
rect 15510 -375 15515 -345
rect 15545 -375 15560 -345
rect 15590 -375 15605 -345
rect 15635 -365 16425 -345
rect 16455 -365 16545 -335
rect 16575 -365 16665 -335
rect 16695 -365 16785 -335
rect 16815 -365 16905 -335
rect 16935 -365 17025 -335
rect 17055 -365 17145 -335
rect 17175 -365 17265 -335
rect 17295 -365 17385 -335
rect 17415 -365 17505 -335
rect 17535 -365 17625 -335
rect 17655 -365 17945 -335
rect 17975 -365 18065 -335
rect 18095 -365 18185 -335
rect 18215 -365 18305 -335
rect 18335 -365 18425 -335
rect 18455 -365 18545 -335
rect 18575 -365 18665 -335
rect 18695 -365 18785 -335
rect 18815 -365 18905 -335
rect 18935 -365 19025 -335
rect 19055 -365 19145 -335
rect 19175 -365 19180 -335
rect 15635 -370 19180 -365
rect 15635 -375 15640 -370
rect 15510 -380 15640 -375
rect 16095 -390 17730 -385
rect 16095 -420 16100 -390
rect 16130 -420 16485 -390
rect 16515 -420 16845 -390
rect 16875 -420 17205 -390
rect 17235 -420 17565 -390
rect 17595 -420 17695 -390
rect 17725 -420 17730 -390
rect 16095 -425 17730 -420
rect 17870 -390 19505 -385
rect 17870 -420 17875 -390
rect 17905 -420 18005 -390
rect 18035 -420 18365 -390
rect 18395 -420 18725 -390
rect 18755 -420 19085 -390
rect 19115 -420 19470 -390
rect 19500 -420 19505 -390
rect 17870 -425 19505 -420
rect 16845 -445 16875 -425
rect 18725 -440 18755 -425
rect 16600 -560 16640 -555
rect 16600 -590 16605 -560
rect 16635 -565 16640 -560
rect 16960 -560 17000 -555
rect 16960 -565 16965 -560
rect 16635 -585 16965 -565
rect 16635 -590 16640 -585
rect 16600 -595 16640 -590
rect 16960 -590 16965 -585
rect 16995 -565 17000 -560
rect 17320 -560 17360 -555
rect 17320 -565 17325 -560
rect 16995 -585 17325 -565
rect 16995 -590 17000 -585
rect 16960 -595 17000 -590
rect 17320 -590 17325 -585
rect 17355 -590 17360 -560
rect 17320 -595 17360 -590
rect 18240 -560 18280 -555
rect 18240 -590 18245 -560
rect 18275 -565 18280 -560
rect 18600 -560 18640 -555
rect 18600 -565 18605 -560
rect 18275 -585 18605 -565
rect 18275 -590 18280 -585
rect 18240 -595 18280 -590
rect 18600 -590 18605 -585
rect 18635 -565 18640 -560
rect 18960 -560 19000 -555
rect 18960 -565 18965 -560
rect 18635 -585 18965 -565
rect 18635 -590 18640 -585
rect 18600 -595 18640 -590
rect 18960 -590 18965 -585
rect 18995 -590 19000 -560
rect 18960 -595 19000 -590
rect 15905 -620 17570 -615
rect 15905 -650 15910 -620
rect 15940 -650 15950 -620
rect 15980 -650 15990 -620
rect 16020 -650 16515 -620
rect 16545 -650 16725 -620
rect 16755 -650 16845 -620
rect 16875 -650 17085 -620
rect 17115 -650 17205 -620
rect 17235 -650 17445 -620
rect 17475 -650 17535 -620
rect 17565 -650 17570 -620
rect 15905 -660 17570 -650
rect 18030 -620 19130 -615
rect 18030 -650 18035 -620
rect 18065 -650 18125 -620
rect 18155 -650 18365 -620
rect 18395 -650 18485 -620
rect 18515 -650 18725 -620
rect 18755 -650 18845 -620
rect 18875 -650 19055 -620
rect 19085 -650 19095 -620
rect 19125 -650 19130 -620
rect 18030 -655 19130 -650
rect 15905 -690 15910 -660
rect 15940 -690 15950 -660
rect 15980 -690 15990 -660
rect 16020 -690 16515 -660
rect 16545 -690 16725 -660
rect 16755 -690 16845 -660
rect 16875 -690 17085 -660
rect 17115 -690 17205 -660
rect 17235 -690 17445 -660
rect 17475 -690 17535 -660
rect 17565 -690 17570 -660
rect 15905 -700 17570 -690
rect 15905 -730 15910 -700
rect 15940 -730 15950 -700
rect 15980 -730 15990 -700
rect 16020 -730 16515 -700
rect 16545 -730 16725 -700
rect 16755 -730 16845 -700
rect 16875 -730 17085 -700
rect 17115 -730 17205 -700
rect 17235 -730 17445 -700
rect 17475 -730 17535 -700
rect 17565 -730 17570 -700
rect 15905 -735 17570 -730
rect 16260 -755 16300 -750
rect 16260 -785 16265 -755
rect 16295 -760 16300 -755
rect 17005 -755 17037 -750
rect 17005 -760 17007 -755
rect 16295 -780 17007 -760
rect 16295 -785 16300 -780
rect 16260 -790 16300 -785
rect 17005 -785 17007 -780
rect 18563 -755 19345 -750
rect 18562 -780 18563 -760
rect 17005 -790 17037 -785
rect 18593 -785 19310 -755
rect 19340 -785 19345 -755
rect 18563 -790 19345 -785
rect 17560 -815 18040 -810
rect 17560 -845 17565 -815
rect 17595 -845 17745 -815
rect 17775 -845 17785 -815
rect 17815 -845 17825 -815
rect 17855 -845 18005 -815
rect 18035 -845 18040 -815
rect 17560 -855 18040 -845
rect 17560 -885 17565 -855
rect 17595 -885 17745 -855
rect 17775 -885 17785 -855
rect 17815 -885 17825 -855
rect 17855 -885 18005 -855
rect 18035 -885 18040 -855
rect 17560 -895 18040 -885
rect 17560 -925 17565 -895
rect 17595 -925 17745 -895
rect 17775 -925 17785 -895
rect 17815 -925 17825 -895
rect 17855 -925 18005 -895
rect 18035 -925 18040 -895
rect 17560 -930 18040 -925
rect 16315 -1075 16355 -1070
rect 16315 -1105 16320 -1075
rect 16350 -1080 16355 -1075
rect 17075 -1075 17105 -1070
rect 16350 -1100 17075 -1080
rect 16350 -1105 16355 -1100
rect 16315 -1110 16355 -1105
rect 17075 -1110 17105 -1105
rect 18440 -1075 19265 -1070
rect 18470 -1105 19230 -1075
rect 19260 -1105 19265 -1075
rect 18440 -1110 19265 -1105
rect 16530 -1130 17060 -1125
rect 16530 -1160 16535 -1130
rect 16565 -1160 17025 -1130
rect 17055 -1160 17060 -1130
rect 16530 -1165 17060 -1160
rect 18540 -1130 19070 -1125
rect 18540 -1160 18545 -1130
rect 18575 -1160 19035 -1130
rect 19065 -1160 19070 -1130
rect 18540 -1165 19070 -1160
rect 15510 -1185 18980 -1180
rect 15510 -1215 15515 -1185
rect 15545 -1215 15560 -1185
rect 15590 -1215 15605 -1185
rect 15635 -1215 16625 -1185
rect 16655 -1215 16745 -1185
rect 16775 -1215 16865 -1185
rect 16895 -1215 16985 -1185
rect 17015 -1215 17305 -1185
rect 17335 -1215 17425 -1185
rect 17455 -1215 17545 -1185
rect 17575 -1215 18025 -1185
rect 18055 -1215 18145 -1185
rect 18175 -1215 18265 -1185
rect 18295 -1215 18585 -1185
rect 18615 -1215 18705 -1185
rect 18735 -1215 18825 -1185
rect 18855 -1215 18945 -1185
rect 18975 -1215 18980 -1185
rect 15510 -1225 18980 -1215
rect 15510 -1230 16625 -1225
rect 15510 -1260 15515 -1230
rect 15545 -1260 15560 -1230
rect 15590 -1260 15605 -1230
rect 15635 -1255 16625 -1230
rect 16655 -1255 16745 -1225
rect 16775 -1255 16865 -1225
rect 16895 -1255 16985 -1225
rect 17015 -1255 17305 -1225
rect 17335 -1255 17425 -1225
rect 17455 -1255 17545 -1225
rect 17575 -1255 18025 -1225
rect 18055 -1255 18145 -1225
rect 18175 -1255 18265 -1225
rect 18295 -1255 18585 -1225
rect 18615 -1255 18705 -1225
rect 18735 -1255 18825 -1225
rect 18855 -1255 18945 -1225
rect 18975 -1255 18980 -1225
rect 15635 -1260 18980 -1255
rect 15510 -1265 18980 -1260
rect 15510 -1275 16625 -1265
rect 15510 -1305 15515 -1275
rect 15545 -1305 15560 -1275
rect 15590 -1305 15605 -1275
rect 15635 -1295 16625 -1275
rect 16655 -1295 16745 -1265
rect 16775 -1295 16865 -1265
rect 16895 -1295 16985 -1265
rect 17015 -1295 17305 -1265
rect 17335 -1295 17425 -1265
rect 17455 -1295 17545 -1265
rect 17575 -1295 18025 -1265
rect 18055 -1295 18145 -1265
rect 18175 -1295 18265 -1265
rect 18295 -1295 18585 -1265
rect 18615 -1295 18705 -1265
rect 18735 -1295 18825 -1265
rect 18855 -1295 18945 -1265
rect 18975 -1295 18980 -1265
rect 15635 -1300 18980 -1295
rect 15635 -1305 15640 -1300
rect 15510 -1310 15640 -1305
rect 17110 -1585 19675 -1580
rect 17110 -1615 17115 -1585
rect 17145 -1615 17745 -1585
rect 17775 -1615 17785 -1585
rect 17815 -1615 17825 -1585
rect 17855 -1615 18455 -1585
rect 18485 -1615 19550 -1585
rect 19580 -1615 19595 -1585
rect 19625 -1615 19640 -1585
rect 19670 -1615 19675 -1585
rect 17110 -1625 19675 -1615
rect 17110 -1655 17115 -1625
rect 17145 -1655 17745 -1625
rect 17775 -1655 17785 -1625
rect 17815 -1655 17825 -1625
rect 17855 -1655 18455 -1625
rect 18485 -1630 19675 -1625
rect 18485 -1655 19550 -1630
rect 17110 -1660 19550 -1655
rect 19580 -1660 19595 -1630
rect 19625 -1660 19640 -1630
rect 19670 -1660 19675 -1630
rect 17110 -1665 19675 -1660
rect 17110 -1695 17115 -1665
rect 17145 -1695 17745 -1665
rect 17775 -1695 17785 -1665
rect 17815 -1695 17825 -1665
rect 17855 -1695 18455 -1665
rect 18485 -1675 19675 -1665
rect 18485 -1695 19550 -1675
rect 17110 -1700 19550 -1695
rect 19545 -1705 19550 -1700
rect 19580 -1705 19595 -1675
rect 19625 -1705 19640 -1675
rect 19670 -1705 19675 -1675
rect 19545 -1710 19675 -1705
rect 16740 -1720 16780 -1715
rect 16740 -1750 16745 -1720
rect 16775 -1725 16780 -1720
rect 16820 -1720 16860 -1715
rect 16820 -1725 16825 -1720
rect 16775 -1745 16825 -1725
rect 16775 -1750 16780 -1745
rect 16740 -1755 16780 -1750
rect 16820 -1750 16825 -1745
rect 16855 -1725 16860 -1720
rect 16900 -1720 16940 -1715
rect 16900 -1725 16905 -1720
rect 16855 -1745 16905 -1725
rect 16855 -1750 16860 -1745
rect 16820 -1755 16860 -1750
rect 16900 -1750 16905 -1745
rect 16935 -1725 16940 -1720
rect 16980 -1720 17020 -1715
rect 16980 -1725 16985 -1720
rect 16935 -1745 16985 -1725
rect 16935 -1750 16940 -1745
rect 16900 -1755 16940 -1750
rect 16980 -1750 16985 -1745
rect 17015 -1725 17020 -1720
rect 17060 -1720 17100 -1715
rect 17060 -1725 17065 -1720
rect 17015 -1745 17065 -1725
rect 17015 -1750 17020 -1745
rect 16980 -1755 17020 -1750
rect 17060 -1750 17065 -1745
rect 17095 -1725 17100 -1720
rect 17140 -1720 17180 -1715
rect 17140 -1725 17145 -1720
rect 17095 -1745 17145 -1725
rect 17095 -1750 17100 -1745
rect 17060 -1755 17100 -1750
rect 17140 -1750 17145 -1745
rect 17175 -1725 17180 -1720
rect 17220 -1720 17260 -1715
rect 17220 -1725 17225 -1720
rect 17175 -1745 17225 -1725
rect 17175 -1750 17180 -1745
rect 17140 -1755 17180 -1750
rect 17220 -1750 17225 -1745
rect 17255 -1725 17260 -1720
rect 17300 -1720 17340 -1715
rect 17300 -1725 17305 -1720
rect 17255 -1745 17305 -1725
rect 17255 -1750 17260 -1745
rect 17220 -1755 17260 -1750
rect 17300 -1750 17305 -1745
rect 17335 -1725 17340 -1720
rect 17380 -1720 17420 -1715
rect 17380 -1725 17385 -1720
rect 17335 -1745 17385 -1725
rect 17335 -1750 17340 -1745
rect 17300 -1755 17340 -1750
rect 17380 -1750 17385 -1745
rect 17415 -1725 17420 -1720
rect 17460 -1720 17500 -1715
rect 17460 -1725 17465 -1720
rect 17415 -1745 17465 -1725
rect 17415 -1750 17420 -1745
rect 17380 -1755 17420 -1750
rect 17460 -1750 17465 -1745
rect 17495 -1725 17500 -1720
rect 17540 -1720 17580 -1715
rect 17540 -1725 17545 -1720
rect 17495 -1745 17545 -1725
rect 17495 -1750 17500 -1745
rect 17460 -1755 17500 -1750
rect 17540 -1750 17545 -1745
rect 17575 -1725 17580 -1720
rect 17620 -1720 17660 -1715
rect 17620 -1725 17625 -1720
rect 17575 -1745 17625 -1725
rect 17575 -1750 17580 -1745
rect 17540 -1755 17580 -1750
rect 17620 -1750 17625 -1745
rect 17655 -1725 17660 -1720
rect 17700 -1720 17740 -1715
rect 17700 -1725 17705 -1720
rect 17655 -1745 17705 -1725
rect 17655 -1750 17660 -1745
rect 17620 -1755 17660 -1750
rect 17700 -1750 17705 -1745
rect 17735 -1750 17740 -1720
rect 17700 -1755 17740 -1750
rect 17780 -1720 17820 -1715
rect 17780 -1750 17785 -1720
rect 17815 -1725 17820 -1720
rect 17860 -1720 17900 -1715
rect 17860 -1725 17865 -1720
rect 17815 -1745 17865 -1725
rect 17815 -1750 17820 -1745
rect 17780 -1755 17820 -1750
rect 17860 -1750 17865 -1745
rect 17895 -1725 17900 -1720
rect 17940 -1720 17980 -1715
rect 17940 -1725 17945 -1720
rect 17895 -1745 17945 -1725
rect 17895 -1750 17900 -1745
rect 17860 -1755 17900 -1750
rect 17940 -1750 17945 -1745
rect 17975 -1725 17980 -1720
rect 18020 -1720 18060 -1715
rect 18020 -1725 18025 -1720
rect 17975 -1745 18025 -1725
rect 17975 -1750 17980 -1745
rect 17940 -1755 17980 -1750
rect 18020 -1750 18025 -1745
rect 18055 -1725 18060 -1720
rect 18100 -1720 18140 -1715
rect 18100 -1725 18105 -1720
rect 18055 -1745 18105 -1725
rect 18055 -1750 18060 -1745
rect 18020 -1755 18060 -1750
rect 18100 -1750 18105 -1745
rect 18135 -1725 18140 -1720
rect 18180 -1720 18220 -1715
rect 18180 -1725 18185 -1720
rect 18135 -1745 18185 -1725
rect 18135 -1750 18140 -1745
rect 18100 -1755 18140 -1750
rect 18180 -1750 18185 -1745
rect 18215 -1725 18220 -1720
rect 18260 -1720 18300 -1715
rect 18260 -1725 18265 -1720
rect 18215 -1745 18265 -1725
rect 18215 -1750 18220 -1745
rect 18180 -1755 18220 -1750
rect 18260 -1750 18265 -1745
rect 18295 -1725 18300 -1720
rect 18340 -1720 18380 -1715
rect 18340 -1725 18345 -1720
rect 18295 -1745 18345 -1725
rect 18295 -1750 18300 -1745
rect 18260 -1755 18300 -1750
rect 18340 -1750 18345 -1745
rect 18375 -1725 18380 -1720
rect 18420 -1720 18460 -1715
rect 18420 -1725 18425 -1720
rect 18375 -1745 18425 -1725
rect 18375 -1750 18380 -1745
rect 18340 -1755 18380 -1750
rect 18420 -1750 18425 -1745
rect 18455 -1725 18460 -1720
rect 18500 -1720 18540 -1715
rect 18500 -1725 18505 -1720
rect 18455 -1745 18505 -1725
rect 18455 -1750 18460 -1745
rect 18420 -1755 18460 -1750
rect 18500 -1750 18505 -1745
rect 18535 -1725 18540 -1720
rect 18580 -1720 18620 -1715
rect 18580 -1725 18585 -1720
rect 18535 -1745 18585 -1725
rect 18535 -1750 18540 -1745
rect 18500 -1755 18540 -1750
rect 18580 -1750 18585 -1745
rect 18615 -1725 18620 -1720
rect 18660 -1720 18700 -1715
rect 18660 -1725 18665 -1720
rect 18615 -1745 18665 -1725
rect 18615 -1750 18620 -1745
rect 18580 -1755 18620 -1750
rect 18660 -1750 18665 -1745
rect 18695 -1725 18700 -1720
rect 18740 -1720 18780 -1715
rect 18740 -1725 18745 -1720
rect 18695 -1745 18745 -1725
rect 18695 -1750 18700 -1745
rect 18660 -1755 18700 -1750
rect 18740 -1750 18745 -1745
rect 18775 -1750 18780 -1720
rect 18740 -1755 18780 -1750
rect 18895 -1785 19675 -1780
rect 16205 -1805 16245 -1800
rect 16205 -1835 16210 -1805
rect 16240 -1810 16245 -1805
rect 16700 -1805 16740 -1800
rect 16700 -1810 16705 -1805
rect 16240 -1830 16705 -1810
rect 16240 -1835 16245 -1830
rect 16205 -1840 16245 -1835
rect 16700 -1835 16705 -1830
rect 16735 -1835 16740 -1805
rect 16700 -1840 16740 -1835
rect 18895 -1815 18900 -1785
rect 18930 -1815 19550 -1785
rect 19580 -1815 19595 -1785
rect 19625 -1815 19640 -1785
rect 19670 -1815 19675 -1785
rect 18895 -1825 19675 -1815
rect 18895 -1855 18900 -1825
rect 18930 -1830 19675 -1825
rect 18930 -1855 19550 -1830
rect 18895 -1860 19550 -1855
rect 19580 -1860 19595 -1830
rect 19625 -1860 19640 -1830
rect 19670 -1860 19675 -1830
rect 19545 -1865 19675 -1860
rect 18885 -1890 19130 -1885
rect 18885 -1920 18890 -1890
rect 18920 -1920 19095 -1890
rect 19125 -1920 19130 -1890
rect 18885 -1925 19130 -1920
rect 16205 -1945 19265 -1940
rect 16205 -1975 16210 -1945
rect 16240 -1975 19230 -1945
rect 19260 -1975 19265 -1945
rect 16205 -1980 19265 -1975
rect 16315 -2000 16355 -1995
rect 16315 -2030 16320 -2000
rect 16350 -2005 16355 -2000
rect 17425 -2005 17430 -2000
rect 16350 -2025 17430 -2005
rect 16350 -2030 16355 -2025
rect 16315 -2035 16355 -2030
rect 17425 -2035 17430 -2025
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2005 18870 -2000
rect 18164 -2035 18835 -2005
rect 18865 -2035 18870 -2005
rect 18165 -2040 18870 -2035
rect 17425 -2060 19120 -2055
rect 17425 -2090 17430 -2060
rect 17460 -2090 19085 -2060
rect 19115 -2090 19120 -2060
rect 17425 -2095 19120 -2090
rect 16260 -2100 16300 -2095
rect 16260 -2130 16265 -2100
rect 16295 -2105 16300 -2100
rect 16480 -2100 16520 -2095
rect 16480 -2105 16485 -2100
rect 16295 -2125 16485 -2105
rect 16295 -2130 16300 -2125
rect 16260 -2135 16300 -2130
rect 16480 -2130 16485 -2125
rect 16515 -2105 16520 -2100
rect 16730 -2100 16770 -2095
rect 16730 -2105 16735 -2100
rect 16515 -2125 16735 -2105
rect 16515 -2130 16520 -2125
rect 16480 -2135 16520 -2130
rect 16730 -2130 16735 -2125
rect 16765 -2130 16770 -2100
rect 16730 -2135 16770 -2130
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19305 -3090 19340 -3085
rect 16730 -3105 17820 -3100
rect 16730 -3135 16735 -3105
rect 16765 -3135 17785 -3105
rect 17815 -3135 17820 -3105
rect 16730 -3140 17820 -3135
rect 18615 -3105 18870 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 19305 -3130 19340 -3125
rect 19465 -3115 19500 -3110
rect 18615 -3140 18870 -3135
rect 19465 -3160 19500 -3150
rect 16040 -3220 16135 -3215
rect 16040 -3250 16045 -3220
rect 16075 -3221 16135 -3220
rect 16075 -3250 16100 -3221
rect 16040 -3255 16100 -3250
rect 16100 -3261 16135 -3256
rect 16210 -3325 16245 -3320
rect 16210 -3365 16245 -3360
rect 19465 -3789 19500 -3784
rect 19465 -3829 19500 -3824
rect 19475 -3830 19495 -3829
rect 16100 -3894 16135 -3889
rect 16100 -3934 16135 -3929
rect 16210 -3894 16245 -3889
rect 16210 -3934 16245 -3929
rect 19185 -3894 19220 -3889
rect 19185 -3934 19220 -3929
rect 16110 -3935 16130 -3934
rect 16220 -3935 16240 -3934
rect 19190 -3935 19210 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 19545 -4150 19675 -4145
rect 19545 -4155 19550 -4150
rect 16210 -4160 19550 -4155
rect 16210 -4190 16215 -4160
rect 16245 -4190 16610 -4160
rect 16640 -4190 17785 -4160
rect 17815 -4190 18960 -4160
rect 18990 -4190 19185 -4160
rect 19215 -4180 19550 -4160
rect 19580 -4180 19595 -4150
rect 19625 -4180 19640 -4150
rect 19670 -4180 19675 -4150
rect 19215 -4190 19675 -4180
rect 16210 -4195 19675 -4190
rect 16210 -4200 19550 -4195
rect 16210 -4230 16215 -4200
rect 16245 -4230 16610 -4200
rect 16640 -4230 17785 -4200
rect 17815 -4230 18960 -4200
rect 18990 -4230 19185 -4200
rect 19215 -4225 19550 -4200
rect 19580 -4225 19595 -4195
rect 19625 -4225 19640 -4195
rect 19670 -4225 19675 -4195
rect 19215 -4230 19675 -4225
rect 16210 -4240 19675 -4230
rect 16210 -4270 16215 -4240
rect 16245 -4270 16610 -4240
rect 16640 -4270 17785 -4240
rect 17815 -4270 18960 -4240
rect 18990 -4270 19185 -4240
rect 19215 -4270 19550 -4240
rect 19580 -4270 19595 -4240
rect 19625 -4270 19640 -4240
rect 19670 -4270 19675 -4240
rect 16210 -4275 19675 -4270
rect 17250 -4295 17300 -4290
rect 16040 -4300 17300 -4295
rect 16040 -4330 16045 -4300
rect 16075 -4330 17260 -4300
rect 17290 -4330 17300 -4300
rect 16040 -4335 17300 -4330
rect 17250 -4340 17300 -4335
rect 16900 -4360 16950 -4350
rect 16900 -4365 16910 -4360
rect 15905 -4370 16910 -4365
rect 15905 -4400 15910 -4370
rect 15940 -4400 15950 -4370
rect 15980 -4400 15990 -4370
rect 16020 -4390 16910 -4370
rect 16940 -4390 16950 -4360
rect 16020 -4400 16950 -4390
rect 15905 -4410 16950 -4400
rect 15905 -4440 15910 -4410
rect 15940 -4440 15950 -4410
rect 15980 -4440 15990 -4410
rect 16020 -4440 16910 -4410
rect 16940 -4440 16950 -4410
rect 15905 -4450 16950 -4440
rect 15905 -4480 15910 -4450
rect 15940 -4480 15950 -4450
rect 15980 -4480 15990 -4450
rect 16020 -4460 16950 -4450
rect 16020 -4480 16910 -4460
rect 15905 -4485 16910 -4480
rect 16900 -4490 16910 -4485
rect 16940 -4490 16950 -4460
rect 18650 -4445 18700 -4440
rect 18650 -4450 18925 -4445
rect 18650 -4480 18660 -4450
rect 18690 -4480 18890 -4450
rect 18920 -4480 18925 -4450
rect 18650 -4485 18925 -4480
rect 19355 -4450 19505 -4445
rect 19355 -4480 19360 -4450
rect 19390 -4480 19470 -4450
rect 19500 -4480 19505 -4450
rect 19355 -4485 19505 -4480
rect 18650 -4490 18700 -4485
rect 16900 -4500 16950 -4490
rect 16100 -4505 16245 -4500
rect 16100 -4535 16105 -4505
rect 16135 -4535 16210 -4505
rect 16240 -4535 16245 -4505
rect 16100 -4540 16245 -4535
rect 15510 -4560 17995 -4555
rect 15510 -4590 15515 -4560
rect 15545 -4590 15560 -4560
rect 15590 -4590 15605 -4560
rect 15635 -4590 17960 -4560
rect 17990 -4590 17995 -4560
rect 15510 -4595 17995 -4590
<< via2 >>
rect 15515 660 15545 690
rect 15560 660 15590 690
rect 15605 660 15635 690
rect 15515 440 15545 470
rect 15560 440 15590 470
rect 15605 440 15635 470
rect 15515 395 15545 425
rect 15560 395 15590 425
rect 15605 395 15635 425
rect 15515 350 15545 380
rect 15560 350 15590 380
rect 15605 350 15635 380
rect 15515 -285 15545 -255
rect 15560 -285 15590 -255
rect 15605 -285 15635 -255
rect 15515 -330 15545 -300
rect 15560 -330 15590 -300
rect 15605 -330 15635 -300
rect 15515 -375 15545 -345
rect 15560 -375 15590 -345
rect 15605 -375 15635 -345
rect 15515 -1215 15545 -1185
rect 15560 -1215 15590 -1185
rect 15605 -1215 15635 -1185
rect 15515 -1260 15545 -1230
rect 15560 -1260 15590 -1230
rect 15605 -1260 15635 -1230
rect 15515 -1305 15545 -1275
rect 15560 -1305 15590 -1275
rect 15605 -1305 15635 -1275
rect 19550 -1615 19580 -1585
rect 19595 -1615 19625 -1585
rect 19640 -1615 19670 -1585
rect 19550 -1660 19580 -1630
rect 19595 -1660 19625 -1630
rect 19640 -1660 19670 -1630
rect 19550 -1705 19580 -1675
rect 19595 -1705 19625 -1675
rect 19640 -1705 19670 -1675
rect 19550 -1815 19580 -1785
rect 19595 -1815 19625 -1785
rect 19640 -1815 19670 -1785
rect 19550 -1860 19580 -1830
rect 19595 -1860 19625 -1830
rect 19640 -1860 19670 -1830
rect 19550 -4180 19580 -4150
rect 19595 -4180 19625 -4150
rect 19640 -4180 19670 -4150
rect 19550 -4225 19580 -4195
rect 19595 -4225 19625 -4195
rect 19640 -4225 19670 -4195
rect 19550 -4270 19580 -4240
rect 19595 -4270 19625 -4240
rect 19640 -4270 19670 -4240
rect 17260 -4330 17290 -4300
rect 16910 -4390 16940 -4360
rect 16910 -4440 16940 -4410
rect 16910 -4490 16940 -4460
rect 18660 -4480 18690 -4450
rect 19360 -4480 19390 -4450
rect 16210 -4535 16240 -4505
rect 15515 -4590 15545 -4560
rect 15560 -4590 15590 -4560
rect 15605 -4590 15635 -4560
rect 17960 -4590 17990 -4560
<< metal3 >>
rect 15510 690 15640 695
rect 15510 660 15515 690
rect 15545 660 15560 690
rect 15590 660 15605 690
rect 15635 660 15640 690
rect 15510 470 15640 660
rect 15510 440 15515 470
rect 15545 440 15560 470
rect 15590 440 15605 470
rect 15635 440 15640 470
rect 15510 425 15640 440
rect 15510 395 15515 425
rect 15545 395 15560 425
rect 15590 395 15605 425
rect 15635 395 15640 425
rect 15510 380 15640 395
rect 15510 350 15515 380
rect 15545 350 15560 380
rect 15590 350 15605 380
rect 15635 350 15640 380
rect 15510 -255 15640 350
rect 15510 -285 15515 -255
rect 15545 -285 15560 -255
rect 15590 -285 15605 -255
rect 15635 -285 15640 -255
rect 15510 -300 15640 -285
rect 15510 -330 15515 -300
rect 15545 -330 15560 -300
rect 15590 -330 15605 -300
rect 15635 -330 15640 -300
rect 15510 -345 15640 -330
rect 15510 -375 15515 -345
rect 15545 -375 15560 -345
rect 15590 -375 15605 -345
rect 15635 -375 15640 -345
rect 15510 -1185 15640 -375
rect 15510 -1215 15515 -1185
rect 15545 -1215 15560 -1185
rect 15590 -1215 15605 -1185
rect 15635 -1215 15640 -1185
rect 15510 -1230 15640 -1215
rect 15510 -1260 15515 -1230
rect 15545 -1260 15560 -1230
rect 15590 -1260 15605 -1230
rect 15635 -1260 15640 -1230
rect 15510 -1275 15640 -1260
rect 15510 -1305 15515 -1275
rect 15545 -1305 15560 -1275
rect 15590 -1305 15605 -1275
rect 15635 -1305 15640 -1275
rect 15510 -4560 15640 -1305
rect 19545 -1585 19675 -1580
rect 19545 -1615 19550 -1585
rect 19580 -1615 19595 -1585
rect 19625 -1615 19640 -1585
rect 19670 -1615 19675 -1585
rect 19545 -1630 19675 -1615
rect 19545 -1660 19550 -1630
rect 19580 -1660 19595 -1630
rect 19625 -1660 19640 -1630
rect 19670 -1660 19675 -1630
rect 19545 -1675 19675 -1660
rect 19545 -1705 19550 -1675
rect 19580 -1705 19595 -1675
rect 19625 -1705 19640 -1675
rect 19670 -1705 19675 -1675
rect 19545 -1785 19675 -1705
rect 19545 -1815 19550 -1785
rect 19580 -1815 19595 -1785
rect 19625 -1815 19640 -1785
rect 19670 -1815 19675 -1785
rect 19545 -1830 19675 -1815
rect 19545 -1860 19550 -1830
rect 19580 -1860 19595 -1830
rect 19625 -1860 19640 -1830
rect 19670 -1860 19675 -1830
rect 19545 -4150 19675 -1860
rect 19545 -4180 19550 -4150
rect 19580 -4180 19595 -4150
rect 19625 -4180 19640 -4150
rect 19670 -4180 19675 -4150
rect 19545 -4195 19675 -4180
rect 19545 -4225 19550 -4195
rect 19580 -4225 19595 -4195
rect 19625 -4225 19640 -4195
rect 19670 -4225 19675 -4195
rect 19545 -4240 19675 -4225
rect 19545 -4270 19550 -4240
rect 19580 -4270 19595 -4240
rect 19625 -4270 19640 -4240
rect 19670 -4270 19675 -4240
rect 19545 -4275 19675 -4270
rect 17250 -4295 17300 -4290
rect 17250 -4335 17255 -4295
rect 17295 -4335 17300 -4295
rect 17250 -4340 17300 -4335
rect 16900 -4355 16950 -4350
rect 16900 -4395 16905 -4355
rect 16945 -4395 16950 -4355
rect 16900 -4405 16950 -4395
rect 16900 -4445 16905 -4405
rect 16945 -4445 16950 -4405
rect 16900 -4455 16950 -4445
rect 16900 -4495 16905 -4455
rect 16945 -4495 16950 -4455
rect 18650 -4445 18700 -4440
rect 18650 -4485 18655 -4445
rect 18695 -4485 18700 -4445
rect 18650 -4490 18700 -4485
rect 19355 -4450 19395 -4445
rect 19355 -4480 19360 -4450
rect 19390 -4480 19395 -4450
rect 16900 -4500 16950 -4495
rect 15510 -4590 15515 -4560
rect 15545 -4590 15560 -4560
rect 15590 -4590 15605 -4560
rect 15635 -4590 15640 -4560
rect 15510 -4595 15640 -4590
rect 16205 -4505 16245 -4500
rect 16205 -4535 16210 -4505
rect 16240 -4535 16245 -4505
rect 16205 -4620 16245 -4535
rect 17955 -4560 17995 -4555
rect 17955 -4590 17960 -4560
rect 17990 -4590 17995 -4560
rect 17955 -4620 17995 -4590
rect 19355 -4620 19395 -4480
rect 15760 -4715 15990 -4620
rect 16110 -4715 16340 -4620
rect 16460 -4715 16690 -4620
rect 16810 -4715 17040 -4620
rect 15760 -4765 17040 -4715
rect 15760 -4850 15990 -4765
rect 16110 -4850 16340 -4765
rect 16460 -4850 16690 -4765
rect 16810 -4850 17040 -4765
rect 17160 -4715 17390 -4620
rect 17510 -4715 17740 -4620
rect 17860 -4715 18090 -4620
rect 18210 -4715 18440 -4620
rect 17160 -4765 18440 -4715
rect 17160 -4850 17390 -4765
rect 17510 -4850 17740 -4765
rect 17860 -4850 18090 -4765
rect 18210 -4850 18440 -4765
rect 18560 -4715 18790 -4620
rect 18910 -4715 19140 -4620
rect 19260 -4715 19490 -4620
rect 19610 -4715 19840 -4620
rect 18560 -4765 19840 -4715
rect 18560 -4850 18790 -4765
rect 18910 -4850 19140 -4765
rect 19260 -4850 19490 -4765
rect 19610 -4850 19840 -4765
rect 16200 -4970 16250 -4850
rect 17950 -4970 18000 -4850
rect 19350 -4970 19400 -4850
rect 15760 -5065 15990 -4970
rect 16110 -5065 16340 -4970
rect 16460 -5065 16690 -4970
rect 16810 -5065 17040 -4970
rect 15760 -5115 17040 -5065
rect 15760 -5200 15990 -5115
rect 16110 -5200 16340 -5115
rect 16460 -5200 16690 -5115
rect 16810 -5200 17040 -5115
rect 17160 -5065 17390 -4970
rect 17510 -5065 17740 -4970
rect 17860 -5065 18090 -4970
rect 18210 -5065 18440 -4970
rect 17160 -5115 18440 -5065
rect 17160 -5200 17390 -5115
rect 17510 -5200 17740 -5115
rect 17860 -5200 18090 -5115
rect 18210 -5200 18440 -5115
rect 18560 -5065 18790 -4970
rect 18910 -5065 19140 -4970
rect 19260 -5065 19490 -4970
rect 19610 -5065 19840 -4970
rect 18560 -5115 19840 -5065
rect 18560 -5200 18790 -5115
rect 18910 -5200 19140 -5115
rect 19260 -5200 19490 -5115
rect 19610 -5200 19840 -5115
rect 16200 -5320 16250 -5200
rect 17950 -5320 18000 -5200
rect 19350 -5320 19400 -5200
rect 15760 -5415 15990 -5320
rect 16110 -5415 16340 -5320
rect 16460 -5415 16690 -5320
rect 16810 -5415 17040 -5320
rect 15760 -5465 17040 -5415
rect 15760 -5550 15990 -5465
rect 16110 -5550 16340 -5465
rect 16460 -5550 16690 -5465
rect 16810 -5550 17040 -5465
rect 17160 -5415 17390 -5320
rect 17510 -5415 17740 -5320
rect 17860 -5415 18090 -5320
rect 18210 -5415 18440 -5320
rect 17160 -5465 18440 -5415
rect 17160 -5550 17390 -5465
rect 17510 -5550 17740 -5465
rect 17860 -5550 18090 -5465
rect 18210 -5550 18440 -5465
rect 18560 -5415 18790 -5320
rect 18910 -5415 19140 -5320
rect 19260 -5415 19490 -5320
rect 19610 -5415 19840 -5320
rect 18560 -5465 19840 -5415
rect 18560 -5550 18790 -5465
rect 18910 -5550 19140 -5465
rect 19260 -5550 19490 -5465
rect 19610 -5550 19840 -5465
rect 16200 -5670 16250 -5550
rect 17950 -5670 18000 -5550
rect 19350 -5670 19400 -5550
rect 15760 -5765 15990 -5670
rect 16110 -5765 16340 -5670
rect 16460 -5765 16690 -5670
rect 16810 -5765 17040 -5670
rect 15760 -5815 17040 -5765
rect 15760 -5900 15990 -5815
rect 16110 -5900 16340 -5815
rect 16460 -5900 16690 -5815
rect 16810 -5900 17040 -5815
rect 17160 -5765 17390 -5670
rect 17510 -5765 17740 -5670
rect 17860 -5765 18090 -5670
rect 18210 -5765 18440 -5670
rect 17160 -5815 18440 -5765
rect 17160 -5900 17390 -5815
rect 17510 -5900 17740 -5815
rect 17860 -5900 18090 -5815
rect 18210 -5900 18440 -5815
rect 18560 -5765 18790 -5670
rect 18910 -5765 19140 -5670
rect 19260 -5765 19490 -5670
rect 19610 -5765 19840 -5670
rect 18560 -5815 19840 -5765
rect 18560 -5900 18790 -5815
rect 18910 -5900 19140 -5815
rect 19260 -5900 19490 -5815
rect 19610 -5900 19840 -5815
rect 16200 -6020 16250 -5900
rect 17950 -6020 18000 -5900
rect 19350 -6020 19400 -5900
rect 15760 -6115 15990 -6020
rect 16110 -6115 16340 -6020
rect 16460 -6115 16690 -6020
rect 16810 -6115 17040 -6020
rect 15760 -6165 17040 -6115
rect 15760 -6250 15990 -6165
rect 16110 -6250 16340 -6165
rect 16460 -6250 16690 -6165
rect 16810 -6250 17040 -6165
rect 17160 -6115 17390 -6020
rect 17510 -6115 17740 -6020
rect 17860 -6115 18090 -6020
rect 18210 -6115 18440 -6020
rect 17160 -6165 18440 -6115
rect 17160 -6250 17390 -6165
rect 17510 -6250 17740 -6165
rect 17860 -6250 18090 -6165
rect 18210 -6250 18440 -6165
rect 18560 -6115 18790 -6020
rect 18910 -6115 19140 -6020
rect 19260 -6115 19490 -6020
rect 19610 -6115 19840 -6020
rect 18560 -6165 19840 -6115
rect 18560 -6250 18790 -6165
rect 18910 -6250 19140 -6165
rect 19260 -6250 19490 -6165
rect 19610 -6250 19840 -6165
<< via3 >>
rect 17255 -4300 17295 -4295
rect 17255 -4330 17260 -4300
rect 17260 -4330 17290 -4300
rect 17290 -4330 17295 -4300
rect 17255 -4335 17295 -4330
rect 16905 -4360 16945 -4355
rect 16905 -4390 16910 -4360
rect 16910 -4390 16940 -4360
rect 16940 -4390 16945 -4360
rect 16905 -4395 16945 -4390
rect 16905 -4410 16945 -4405
rect 16905 -4440 16910 -4410
rect 16910 -4440 16940 -4410
rect 16940 -4440 16945 -4410
rect 16905 -4445 16945 -4440
rect 16905 -4460 16945 -4455
rect 16905 -4490 16910 -4460
rect 16910 -4490 16940 -4460
rect 16940 -4490 16945 -4460
rect 16905 -4495 16945 -4490
rect 18655 -4450 18695 -4445
rect 18655 -4480 18660 -4450
rect 18660 -4480 18690 -4450
rect 18690 -4480 18695 -4450
rect 18655 -4485 18695 -4480
<< mimcap >>
rect 15775 -4720 15975 -4635
rect 15775 -4760 15855 -4720
rect 15895 -4760 15975 -4720
rect 15775 -4835 15975 -4760
rect 16125 -4720 16325 -4635
rect 16125 -4760 16205 -4720
rect 16245 -4760 16325 -4720
rect 16125 -4835 16325 -4760
rect 16475 -4720 16675 -4635
rect 16475 -4760 16555 -4720
rect 16595 -4760 16675 -4720
rect 16475 -4835 16675 -4760
rect 16825 -4720 17025 -4635
rect 16825 -4760 16905 -4720
rect 16945 -4760 17025 -4720
rect 16825 -4835 17025 -4760
rect 17175 -4720 17375 -4635
rect 17175 -4760 17255 -4720
rect 17295 -4760 17375 -4720
rect 17175 -4835 17375 -4760
rect 17525 -4720 17725 -4635
rect 17525 -4760 17605 -4720
rect 17645 -4760 17725 -4720
rect 17525 -4835 17725 -4760
rect 17875 -4720 18075 -4635
rect 17875 -4760 17955 -4720
rect 17995 -4760 18075 -4720
rect 17875 -4835 18075 -4760
rect 18225 -4720 18425 -4635
rect 18225 -4760 18305 -4720
rect 18345 -4760 18425 -4720
rect 18225 -4835 18425 -4760
rect 18575 -4720 18775 -4635
rect 18575 -4760 18655 -4720
rect 18695 -4760 18775 -4720
rect 18575 -4835 18775 -4760
rect 18925 -4720 19125 -4635
rect 18925 -4760 19005 -4720
rect 19045 -4760 19125 -4720
rect 18925 -4835 19125 -4760
rect 19275 -4720 19475 -4635
rect 19275 -4760 19355 -4720
rect 19395 -4760 19475 -4720
rect 19275 -4835 19475 -4760
rect 19625 -4720 19825 -4635
rect 19625 -4760 19705 -4720
rect 19745 -4760 19825 -4720
rect 19625 -4835 19825 -4760
rect 15775 -5070 15975 -4985
rect 15775 -5110 15855 -5070
rect 15895 -5110 15975 -5070
rect 15775 -5185 15975 -5110
rect 16125 -5070 16325 -4985
rect 16125 -5110 16205 -5070
rect 16245 -5110 16325 -5070
rect 16125 -5185 16325 -5110
rect 16475 -5070 16675 -4985
rect 16475 -5110 16555 -5070
rect 16595 -5110 16675 -5070
rect 16475 -5185 16675 -5110
rect 16825 -5070 17025 -4985
rect 16825 -5110 16905 -5070
rect 16945 -5110 17025 -5070
rect 16825 -5185 17025 -5110
rect 17175 -5070 17375 -4985
rect 17175 -5110 17255 -5070
rect 17295 -5110 17375 -5070
rect 17175 -5185 17375 -5110
rect 17525 -5070 17725 -4985
rect 17525 -5110 17605 -5070
rect 17645 -5110 17725 -5070
rect 17525 -5185 17725 -5110
rect 17875 -5070 18075 -4985
rect 17875 -5110 17955 -5070
rect 17995 -5110 18075 -5070
rect 17875 -5185 18075 -5110
rect 18225 -5070 18425 -4985
rect 18225 -5110 18305 -5070
rect 18345 -5110 18425 -5070
rect 18225 -5185 18425 -5110
rect 18575 -5070 18775 -4985
rect 18575 -5110 18655 -5070
rect 18695 -5110 18775 -5070
rect 18575 -5185 18775 -5110
rect 18925 -5070 19125 -4985
rect 18925 -5110 19005 -5070
rect 19045 -5110 19125 -5070
rect 18925 -5185 19125 -5110
rect 19275 -5070 19475 -4985
rect 19275 -5110 19355 -5070
rect 19395 -5110 19475 -5070
rect 19275 -5185 19475 -5110
rect 19625 -5070 19825 -4985
rect 19625 -5110 19705 -5070
rect 19745 -5110 19825 -5070
rect 19625 -5185 19825 -5110
rect 15775 -5420 15975 -5335
rect 15775 -5460 15855 -5420
rect 15895 -5460 15975 -5420
rect 15775 -5535 15975 -5460
rect 16125 -5420 16325 -5335
rect 16125 -5460 16205 -5420
rect 16245 -5460 16325 -5420
rect 16125 -5535 16325 -5460
rect 16475 -5420 16675 -5335
rect 16475 -5460 16555 -5420
rect 16595 -5460 16675 -5420
rect 16475 -5535 16675 -5460
rect 16825 -5420 17025 -5335
rect 16825 -5460 16905 -5420
rect 16945 -5460 17025 -5420
rect 16825 -5535 17025 -5460
rect 17175 -5420 17375 -5335
rect 17175 -5460 17255 -5420
rect 17295 -5460 17375 -5420
rect 17175 -5535 17375 -5460
rect 17525 -5420 17725 -5335
rect 17525 -5460 17605 -5420
rect 17645 -5460 17725 -5420
rect 17525 -5535 17725 -5460
rect 17875 -5420 18075 -5335
rect 17875 -5460 17955 -5420
rect 17995 -5460 18075 -5420
rect 17875 -5535 18075 -5460
rect 18225 -5420 18425 -5335
rect 18225 -5460 18305 -5420
rect 18345 -5460 18425 -5420
rect 18225 -5535 18425 -5460
rect 18575 -5420 18775 -5335
rect 18575 -5460 18655 -5420
rect 18695 -5460 18775 -5420
rect 18575 -5535 18775 -5460
rect 18925 -5420 19125 -5335
rect 18925 -5460 19005 -5420
rect 19045 -5460 19125 -5420
rect 18925 -5535 19125 -5460
rect 19275 -5420 19475 -5335
rect 19275 -5460 19355 -5420
rect 19395 -5460 19475 -5420
rect 19275 -5535 19475 -5460
rect 19625 -5420 19825 -5335
rect 19625 -5460 19705 -5420
rect 19745 -5460 19825 -5420
rect 19625 -5535 19825 -5460
rect 15775 -5770 15975 -5685
rect 15775 -5810 15855 -5770
rect 15895 -5810 15975 -5770
rect 15775 -5885 15975 -5810
rect 16125 -5770 16325 -5685
rect 16125 -5810 16205 -5770
rect 16245 -5810 16325 -5770
rect 16125 -5885 16325 -5810
rect 16475 -5770 16675 -5685
rect 16475 -5810 16555 -5770
rect 16595 -5810 16675 -5770
rect 16475 -5885 16675 -5810
rect 16825 -5770 17025 -5685
rect 16825 -5810 16905 -5770
rect 16945 -5810 17025 -5770
rect 16825 -5885 17025 -5810
rect 17175 -5770 17375 -5685
rect 17175 -5810 17255 -5770
rect 17295 -5810 17375 -5770
rect 17175 -5885 17375 -5810
rect 17525 -5770 17725 -5685
rect 17525 -5810 17605 -5770
rect 17645 -5810 17725 -5770
rect 17525 -5885 17725 -5810
rect 17875 -5770 18075 -5685
rect 17875 -5810 17955 -5770
rect 17995 -5810 18075 -5770
rect 17875 -5885 18075 -5810
rect 18225 -5770 18425 -5685
rect 18225 -5810 18305 -5770
rect 18345 -5810 18425 -5770
rect 18225 -5885 18425 -5810
rect 18575 -5770 18775 -5685
rect 18575 -5810 18655 -5770
rect 18695 -5810 18775 -5770
rect 18575 -5885 18775 -5810
rect 18925 -5770 19125 -5685
rect 18925 -5810 19005 -5770
rect 19045 -5810 19125 -5770
rect 18925 -5885 19125 -5810
rect 19275 -5770 19475 -5685
rect 19275 -5810 19355 -5770
rect 19395 -5810 19475 -5770
rect 19275 -5885 19475 -5810
rect 19625 -5770 19825 -5685
rect 19625 -5810 19705 -5770
rect 19745 -5810 19825 -5770
rect 19625 -5885 19825 -5810
rect 15775 -6120 15975 -6035
rect 15775 -6160 15855 -6120
rect 15895 -6160 15975 -6120
rect 15775 -6235 15975 -6160
rect 16125 -6120 16325 -6035
rect 16125 -6160 16205 -6120
rect 16245 -6160 16325 -6120
rect 16125 -6235 16325 -6160
rect 16475 -6120 16675 -6035
rect 16475 -6160 16555 -6120
rect 16595 -6160 16675 -6120
rect 16475 -6235 16675 -6160
rect 16825 -6120 17025 -6035
rect 16825 -6160 16905 -6120
rect 16945 -6160 17025 -6120
rect 16825 -6235 17025 -6160
rect 17175 -6120 17375 -6035
rect 17175 -6160 17255 -6120
rect 17295 -6160 17375 -6120
rect 17175 -6235 17375 -6160
rect 17525 -6120 17725 -6035
rect 17525 -6160 17605 -6120
rect 17645 -6160 17725 -6120
rect 17525 -6235 17725 -6160
rect 17875 -6120 18075 -6035
rect 17875 -6160 17955 -6120
rect 17995 -6160 18075 -6120
rect 17875 -6235 18075 -6160
rect 18225 -6120 18425 -6035
rect 18225 -6160 18305 -6120
rect 18345 -6160 18425 -6120
rect 18225 -6235 18425 -6160
rect 18575 -6120 18775 -6035
rect 18575 -6160 18655 -6120
rect 18695 -6160 18775 -6120
rect 18575 -6235 18775 -6160
rect 18925 -6120 19125 -6035
rect 18925 -6160 19005 -6120
rect 19045 -6160 19125 -6120
rect 18925 -6235 19125 -6160
rect 19275 -6120 19475 -6035
rect 19275 -6160 19355 -6120
rect 19395 -6160 19475 -6120
rect 19275 -6235 19475 -6160
rect 19625 -6120 19825 -6035
rect 19625 -6160 19705 -6120
rect 19745 -6160 19825 -6120
rect 19625 -6235 19825 -6160
<< mimcapcontact >>
rect 15855 -4760 15895 -4720
rect 16205 -4760 16245 -4720
rect 16555 -4760 16595 -4720
rect 16905 -4760 16945 -4720
rect 17255 -4760 17295 -4720
rect 17605 -4760 17645 -4720
rect 17955 -4760 17995 -4720
rect 18305 -4760 18345 -4720
rect 18655 -4760 18695 -4720
rect 19005 -4760 19045 -4720
rect 19355 -4760 19395 -4720
rect 19705 -4760 19745 -4720
rect 15855 -5110 15895 -5070
rect 16205 -5110 16245 -5070
rect 16555 -5110 16595 -5070
rect 16905 -5110 16945 -5070
rect 17255 -5110 17295 -5070
rect 17605 -5110 17645 -5070
rect 17955 -5110 17995 -5070
rect 18305 -5110 18345 -5070
rect 18655 -5110 18695 -5070
rect 19005 -5110 19045 -5070
rect 19355 -5110 19395 -5070
rect 19705 -5110 19745 -5070
rect 15855 -5460 15895 -5420
rect 16205 -5460 16245 -5420
rect 16555 -5460 16595 -5420
rect 16905 -5460 16945 -5420
rect 17255 -5460 17295 -5420
rect 17605 -5460 17645 -5420
rect 17955 -5460 17995 -5420
rect 18305 -5460 18345 -5420
rect 18655 -5460 18695 -5420
rect 19005 -5460 19045 -5420
rect 19355 -5460 19395 -5420
rect 19705 -5460 19745 -5420
rect 15855 -5810 15895 -5770
rect 16205 -5810 16245 -5770
rect 16555 -5810 16595 -5770
rect 16905 -5810 16945 -5770
rect 17255 -5810 17295 -5770
rect 17605 -5810 17645 -5770
rect 17955 -5810 17995 -5770
rect 18305 -5810 18345 -5770
rect 18655 -5810 18695 -5770
rect 19005 -5810 19045 -5770
rect 19355 -5810 19395 -5770
rect 19705 -5810 19745 -5770
rect 15855 -6160 15895 -6120
rect 16205 -6160 16245 -6120
rect 16555 -6160 16595 -6120
rect 16905 -6160 16945 -6120
rect 17255 -6160 17295 -6120
rect 17605 -6160 17645 -6120
rect 17955 -6160 17995 -6120
rect 18305 -6160 18345 -6120
rect 18655 -6160 18695 -6120
rect 19005 -6160 19045 -6120
rect 19355 -6160 19395 -6120
rect 19705 -6160 19745 -6120
<< metal4 >>
rect 17250 -4295 17300 -4290
rect 17250 -4335 17255 -4295
rect 17295 -4335 17300 -4295
rect 16900 -4355 16950 -4350
rect 16900 -4395 16905 -4355
rect 16945 -4395 16950 -4355
rect 16900 -4405 16950 -4395
rect 16900 -4445 16905 -4405
rect 16945 -4445 16950 -4405
rect 16900 -4455 16950 -4445
rect 16900 -4495 16905 -4455
rect 16945 -4495 16950 -4455
rect 16900 -4715 16950 -4495
rect 15850 -4720 16950 -4715
rect 15850 -4760 15855 -4720
rect 15895 -4760 16205 -4720
rect 16245 -4760 16555 -4720
rect 16595 -4760 16905 -4720
rect 16945 -4760 16950 -4720
rect 15850 -4765 16950 -4760
rect 17250 -4715 17300 -4335
rect 18650 -4445 18700 -4440
rect 18650 -4485 18655 -4445
rect 18695 -4485 18700 -4445
rect 18650 -4715 18700 -4485
rect 17250 -4720 18350 -4715
rect 17250 -4760 17255 -4720
rect 17295 -4760 17605 -4720
rect 17645 -4760 17955 -4720
rect 17995 -4760 18305 -4720
rect 18345 -4760 18350 -4720
rect 17250 -4765 18350 -4760
rect 18650 -4720 19750 -4715
rect 18650 -4760 18655 -4720
rect 18695 -4760 19005 -4720
rect 19045 -4760 19355 -4720
rect 19395 -4760 19705 -4720
rect 19745 -4760 19750 -4720
rect 18650 -4765 19750 -4760
rect 16200 -5065 16250 -4765
rect 17950 -5065 18000 -4765
rect 19350 -5065 19400 -4765
rect 15850 -5070 16950 -5065
rect 15850 -5110 15855 -5070
rect 15895 -5110 16205 -5070
rect 16245 -5110 16555 -5070
rect 16595 -5110 16905 -5070
rect 16945 -5110 16950 -5070
rect 15850 -5115 16950 -5110
rect 17250 -5070 18350 -5065
rect 17250 -5110 17255 -5070
rect 17295 -5110 17605 -5070
rect 17645 -5110 17955 -5070
rect 17995 -5110 18305 -5070
rect 18345 -5110 18350 -5070
rect 17250 -5115 18350 -5110
rect 18650 -5070 19750 -5065
rect 18650 -5110 18655 -5070
rect 18695 -5110 19005 -5070
rect 19045 -5110 19355 -5070
rect 19395 -5110 19705 -5070
rect 19745 -5110 19750 -5070
rect 18650 -5115 19750 -5110
rect 16200 -5415 16250 -5115
rect 17950 -5415 18000 -5115
rect 19350 -5415 19400 -5115
rect 15850 -5420 16950 -5415
rect 15850 -5460 15855 -5420
rect 15895 -5460 16205 -5420
rect 16245 -5460 16555 -5420
rect 16595 -5460 16905 -5420
rect 16945 -5460 16950 -5420
rect 15850 -5465 16950 -5460
rect 17250 -5420 18350 -5415
rect 17250 -5460 17255 -5420
rect 17295 -5460 17605 -5420
rect 17645 -5460 17955 -5420
rect 17995 -5460 18305 -5420
rect 18345 -5460 18350 -5420
rect 17250 -5465 18350 -5460
rect 18650 -5420 19750 -5415
rect 18650 -5460 18655 -5420
rect 18695 -5460 19005 -5420
rect 19045 -5460 19355 -5420
rect 19395 -5460 19705 -5420
rect 19745 -5460 19750 -5420
rect 18650 -5465 19750 -5460
rect 16200 -5765 16250 -5465
rect 17950 -5765 18000 -5465
rect 19350 -5765 19400 -5465
rect 15850 -5770 16950 -5765
rect 15850 -5810 15855 -5770
rect 15895 -5810 16205 -5770
rect 16245 -5810 16555 -5770
rect 16595 -5810 16905 -5770
rect 16945 -5810 16950 -5770
rect 15850 -5815 16950 -5810
rect 17250 -5770 18350 -5765
rect 17250 -5810 17255 -5770
rect 17295 -5810 17605 -5770
rect 17645 -5810 17955 -5770
rect 17995 -5810 18305 -5770
rect 18345 -5810 18350 -5770
rect 17250 -5815 18350 -5810
rect 18650 -5770 19750 -5765
rect 18650 -5810 18655 -5770
rect 18695 -5810 19005 -5770
rect 19045 -5810 19355 -5770
rect 19395 -5810 19705 -5770
rect 19745 -5810 19750 -5770
rect 18650 -5815 19750 -5810
rect 16200 -6115 16250 -5815
rect 17950 -6115 18000 -5815
rect 19350 -6115 19400 -5815
rect 15850 -6120 16950 -6115
rect 15850 -6160 15855 -6120
rect 15895 -6160 16205 -6120
rect 16245 -6160 16555 -6120
rect 16595 -6160 16905 -6120
rect 16945 -6160 16950 -6120
rect 15850 -6165 16950 -6160
rect 17250 -6120 18350 -6115
rect 17250 -6160 17255 -6120
rect 17295 -6160 17605 -6120
rect 17645 -6160 17955 -6120
rect 17995 -6160 18305 -6120
rect 18345 -6160 18350 -6120
rect 17250 -6165 18350 -6160
rect 18650 -6120 19750 -6115
rect 18650 -6160 18655 -6120
rect 18695 -6160 19005 -6120
rect 19045 -6160 19355 -6120
rect 19395 -6160 19705 -6120
rect 19745 -6160 19750 -6120
rect 18650 -6165 19750 -6160
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel metal1 18780 -1735 18780 -1735 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal1 16235 -1535 16235 -1535 3 FreeSans 400 0 200 0 START_UP
flabel metal2 17060 -1165 17060 -1165 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 18580 -1165 18580 -1165 3 FreeSans 400 180 200 0 V_p_2
flabel metal2 18430 15 18430 15 5 FreeSans 400 0 0 -40 V_TOP
flabel metal2 17570 -635 17570 -635 3 FreeSans 240 0 120 0 1st_Vout_1
flabel metal2 16620 -595 16620 -595 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 18030 -635 18030 -635 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 18930 -1080 18930 -1080 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 16665 -780 16665 -780 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 16670 -1085 16670 -1085 1 FreeSans 400 0 0 80 Vin+
flabel metal1 19505 -625 19505 -625 3 FreeSans 320 0 160 0 V2
flabel metal2 19070 -195 19070 -195 1 FreeSans 320 0 0 160 V1
flabel metal3 19355 -4465 19355 -4465 7 FreeSans 400 180 -40 0 cap_res2
flabel metal2 16145 -4530 16145 -4530 5 FreeSans 400 0 0 -40 cap_res1
flabel metal3 19675 -2560 19675 -2560 3 FreeSans 800 0 400 0 GNDA
port 3 e
flabel metal3 15510 -2525 15510 -2525 7 FreeSans 800 0 -400 0 VDDA
port 1 w
flabel metal1 17380 980 17380 980 1 FreeSans 800 0 400 0 CURRENT_OUTPUT
port 2 n
<< end >>
