magic
tech sky130A
timestamp 1739788113
<< nwell >>
rect 9230 2215 10840 2505
<< nmos >>
rect 9250 1805 9310 2005
rect 9360 1805 9420 2005
rect 9470 1805 9530 2005
rect 9580 1805 9640 2005
rect 9790 1805 9850 2005
rect 9900 1805 9960 2005
rect 10010 1805 10070 2005
rect 10120 1805 10180 2005
rect 10330 1805 10390 2005
rect 10440 1805 10500 2005
rect 10550 1805 10610 2005
rect 10660 1805 10720 2005
<< pmos >>
rect 9350 2285 9410 2485
rect 9460 2285 9520 2485
rect 9570 2285 9630 2485
rect 9680 2285 9740 2485
rect 9790 2285 9850 2485
rect 9900 2285 9960 2485
rect 10110 2285 10170 2485
rect 10220 2285 10280 2485
rect 10330 2285 10390 2485
rect 10440 2285 10500 2485
rect 10550 2285 10610 2485
rect 10660 2285 10720 2485
<< ndiff >>
rect 9200 1990 9250 2005
rect 9200 1970 9215 1990
rect 9235 1970 9250 1990
rect 9200 1940 9250 1970
rect 9200 1920 9215 1940
rect 9235 1920 9250 1940
rect 9200 1890 9250 1920
rect 9200 1870 9215 1890
rect 9235 1870 9250 1890
rect 9200 1840 9250 1870
rect 9200 1820 9215 1840
rect 9235 1820 9250 1840
rect 9200 1805 9250 1820
rect 9310 1990 9360 2005
rect 9310 1970 9325 1990
rect 9345 1970 9360 1990
rect 9310 1940 9360 1970
rect 9310 1920 9325 1940
rect 9345 1920 9360 1940
rect 9310 1890 9360 1920
rect 9310 1870 9325 1890
rect 9345 1870 9360 1890
rect 9310 1840 9360 1870
rect 9310 1820 9325 1840
rect 9345 1820 9360 1840
rect 9310 1805 9360 1820
rect 9420 1990 9470 2005
rect 9420 1970 9435 1990
rect 9455 1970 9470 1990
rect 9420 1940 9470 1970
rect 9420 1920 9435 1940
rect 9455 1920 9470 1940
rect 9420 1890 9470 1920
rect 9420 1870 9435 1890
rect 9455 1870 9470 1890
rect 9420 1840 9470 1870
rect 9420 1820 9435 1840
rect 9455 1820 9470 1840
rect 9420 1805 9470 1820
rect 9530 1990 9580 2005
rect 9530 1970 9545 1990
rect 9565 1970 9580 1990
rect 9530 1940 9580 1970
rect 9530 1920 9545 1940
rect 9565 1920 9580 1940
rect 9530 1890 9580 1920
rect 9530 1870 9545 1890
rect 9565 1870 9580 1890
rect 9530 1840 9580 1870
rect 9530 1820 9545 1840
rect 9565 1820 9580 1840
rect 9530 1805 9580 1820
rect 9640 1990 9690 2005
rect 9740 1990 9790 2005
rect 9640 1970 9655 1990
rect 9675 1970 9690 1990
rect 9740 1970 9755 1990
rect 9775 1970 9790 1990
rect 9640 1940 9690 1970
rect 9740 1940 9790 1970
rect 9640 1920 9655 1940
rect 9675 1920 9690 1940
rect 9740 1920 9755 1940
rect 9775 1920 9790 1940
rect 9640 1890 9690 1920
rect 9740 1890 9790 1920
rect 9640 1870 9655 1890
rect 9675 1870 9690 1890
rect 9740 1870 9755 1890
rect 9775 1870 9790 1890
rect 9640 1840 9690 1870
rect 9740 1840 9790 1870
rect 9640 1820 9655 1840
rect 9675 1820 9690 1840
rect 9740 1820 9755 1840
rect 9775 1820 9790 1840
rect 9640 1805 9690 1820
rect 9740 1805 9790 1820
rect 9850 1990 9900 2005
rect 9850 1970 9865 1990
rect 9885 1970 9900 1990
rect 9850 1940 9900 1970
rect 9850 1920 9865 1940
rect 9885 1920 9900 1940
rect 9850 1890 9900 1920
rect 9850 1870 9865 1890
rect 9885 1870 9900 1890
rect 9850 1840 9900 1870
rect 9850 1820 9865 1840
rect 9885 1820 9900 1840
rect 9850 1805 9900 1820
rect 9960 1990 10010 2005
rect 9960 1970 9975 1990
rect 9995 1970 10010 1990
rect 9960 1940 10010 1970
rect 9960 1920 9975 1940
rect 9995 1920 10010 1940
rect 9960 1890 10010 1920
rect 9960 1870 9975 1890
rect 9995 1870 10010 1890
rect 9960 1840 10010 1870
rect 9960 1820 9975 1840
rect 9995 1820 10010 1840
rect 9960 1805 10010 1820
rect 10070 1990 10120 2005
rect 10070 1970 10085 1990
rect 10105 1970 10120 1990
rect 10070 1940 10120 1970
rect 10070 1920 10085 1940
rect 10105 1920 10120 1940
rect 10070 1890 10120 1920
rect 10070 1870 10085 1890
rect 10105 1870 10120 1890
rect 10070 1840 10120 1870
rect 10070 1820 10085 1840
rect 10105 1820 10120 1840
rect 10070 1805 10120 1820
rect 10180 1990 10230 2005
rect 10280 1990 10330 2005
rect 10180 1970 10195 1990
rect 10215 1970 10230 1990
rect 10280 1970 10295 1990
rect 10315 1970 10330 1990
rect 10180 1940 10230 1970
rect 10280 1940 10330 1970
rect 10180 1920 10195 1940
rect 10215 1920 10230 1940
rect 10280 1920 10295 1940
rect 10315 1920 10330 1940
rect 10180 1890 10230 1920
rect 10280 1890 10330 1920
rect 10180 1870 10195 1890
rect 10215 1870 10230 1890
rect 10280 1870 10295 1890
rect 10315 1870 10330 1890
rect 10180 1840 10230 1870
rect 10280 1840 10330 1870
rect 10180 1820 10195 1840
rect 10215 1820 10230 1840
rect 10280 1820 10295 1840
rect 10315 1820 10330 1840
rect 10180 1805 10230 1820
rect 10280 1805 10330 1820
rect 10390 1990 10440 2005
rect 10390 1970 10405 1990
rect 10425 1970 10440 1990
rect 10390 1940 10440 1970
rect 10390 1920 10405 1940
rect 10425 1920 10440 1940
rect 10390 1890 10440 1920
rect 10390 1870 10405 1890
rect 10425 1870 10440 1890
rect 10390 1840 10440 1870
rect 10390 1820 10405 1840
rect 10425 1820 10440 1840
rect 10390 1805 10440 1820
rect 10500 1990 10550 2005
rect 10500 1970 10515 1990
rect 10535 1970 10550 1990
rect 10500 1940 10550 1970
rect 10500 1920 10515 1940
rect 10535 1920 10550 1940
rect 10500 1890 10550 1920
rect 10500 1870 10515 1890
rect 10535 1870 10550 1890
rect 10500 1840 10550 1870
rect 10500 1820 10515 1840
rect 10535 1820 10550 1840
rect 10500 1805 10550 1820
rect 10610 1990 10660 2005
rect 10610 1970 10625 1990
rect 10645 1970 10660 1990
rect 10610 1940 10660 1970
rect 10610 1920 10625 1940
rect 10645 1920 10660 1940
rect 10610 1890 10660 1920
rect 10610 1870 10625 1890
rect 10645 1870 10660 1890
rect 10610 1840 10660 1870
rect 10610 1820 10625 1840
rect 10645 1820 10660 1840
rect 10610 1805 10660 1820
rect 10720 1990 10770 2005
rect 10720 1970 10735 1990
rect 10755 1970 10770 1990
rect 10720 1940 10770 1970
rect 10720 1920 10735 1940
rect 10755 1920 10770 1940
rect 10720 1890 10770 1920
rect 10720 1870 10735 1890
rect 10755 1870 10770 1890
rect 10720 1840 10770 1870
rect 10720 1820 10735 1840
rect 10755 1820 10770 1840
rect 10720 1805 10770 1820
<< pdiff >>
rect 9300 2470 9350 2485
rect 9300 2450 9315 2470
rect 9335 2450 9350 2470
rect 9300 2420 9350 2450
rect 9300 2400 9315 2420
rect 9335 2400 9350 2420
rect 9300 2370 9350 2400
rect 9300 2350 9315 2370
rect 9335 2350 9350 2370
rect 9300 2320 9350 2350
rect 9300 2300 9315 2320
rect 9335 2300 9350 2320
rect 9300 2285 9350 2300
rect 9410 2470 9460 2485
rect 9410 2450 9425 2470
rect 9445 2450 9460 2470
rect 9410 2420 9460 2450
rect 9410 2400 9425 2420
rect 9445 2400 9460 2420
rect 9410 2370 9460 2400
rect 9410 2350 9425 2370
rect 9445 2350 9460 2370
rect 9410 2320 9460 2350
rect 9410 2300 9425 2320
rect 9445 2300 9460 2320
rect 9410 2285 9460 2300
rect 9520 2470 9570 2485
rect 9520 2450 9535 2470
rect 9555 2450 9570 2470
rect 9520 2420 9570 2450
rect 9520 2400 9535 2420
rect 9555 2400 9570 2420
rect 9520 2370 9570 2400
rect 9520 2350 9535 2370
rect 9555 2350 9570 2370
rect 9520 2320 9570 2350
rect 9520 2300 9535 2320
rect 9555 2300 9570 2320
rect 9520 2285 9570 2300
rect 9630 2470 9680 2485
rect 9630 2450 9645 2470
rect 9665 2450 9680 2470
rect 9630 2420 9680 2450
rect 9630 2400 9645 2420
rect 9665 2400 9680 2420
rect 9630 2370 9680 2400
rect 9630 2350 9645 2370
rect 9665 2350 9680 2370
rect 9630 2320 9680 2350
rect 9630 2300 9645 2320
rect 9665 2300 9680 2320
rect 9630 2285 9680 2300
rect 9740 2470 9790 2485
rect 9740 2450 9755 2470
rect 9775 2450 9790 2470
rect 9740 2420 9790 2450
rect 9740 2400 9755 2420
rect 9775 2400 9790 2420
rect 9740 2370 9790 2400
rect 9740 2350 9755 2370
rect 9775 2350 9790 2370
rect 9740 2320 9790 2350
rect 9740 2300 9755 2320
rect 9775 2300 9790 2320
rect 9740 2285 9790 2300
rect 9850 2470 9900 2485
rect 9850 2450 9865 2470
rect 9885 2450 9900 2470
rect 9850 2420 9900 2450
rect 9850 2400 9865 2420
rect 9885 2400 9900 2420
rect 9850 2370 9900 2400
rect 9850 2350 9865 2370
rect 9885 2350 9900 2370
rect 9850 2320 9900 2350
rect 9850 2300 9865 2320
rect 9885 2300 9900 2320
rect 9850 2285 9900 2300
rect 9960 2470 10010 2485
rect 10060 2470 10110 2485
rect 9960 2450 9975 2470
rect 9995 2450 10010 2470
rect 10060 2450 10075 2470
rect 10095 2450 10110 2470
rect 9960 2420 10010 2450
rect 10060 2420 10110 2450
rect 9960 2400 9975 2420
rect 9995 2400 10010 2420
rect 10060 2400 10075 2420
rect 10095 2400 10110 2420
rect 9960 2370 10010 2400
rect 10060 2370 10110 2400
rect 9960 2350 9975 2370
rect 9995 2350 10010 2370
rect 10060 2350 10075 2370
rect 10095 2350 10110 2370
rect 9960 2320 10010 2350
rect 10060 2320 10110 2350
rect 9960 2300 9975 2320
rect 9995 2300 10010 2320
rect 10060 2300 10075 2320
rect 10095 2300 10110 2320
rect 9960 2285 10010 2300
rect 10060 2285 10110 2300
rect 10170 2470 10220 2485
rect 10170 2450 10185 2470
rect 10205 2450 10220 2470
rect 10170 2420 10220 2450
rect 10170 2400 10185 2420
rect 10205 2400 10220 2420
rect 10170 2370 10220 2400
rect 10170 2350 10185 2370
rect 10205 2350 10220 2370
rect 10170 2320 10220 2350
rect 10170 2300 10185 2320
rect 10205 2300 10220 2320
rect 10170 2285 10220 2300
rect 10280 2470 10330 2485
rect 10280 2450 10295 2470
rect 10315 2450 10330 2470
rect 10280 2420 10330 2450
rect 10280 2400 10295 2420
rect 10315 2400 10330 2420
rect 10280 2370 10330 2400
rect 10280 2350 10295 2370
rect 10315 2350 10330 2370
rect 10280 2320 10330 2350
rect 10280 2300 10295 2320
rect 10315 2300 10330 2320
rect 10280 2285 10330 2300
rect 10390 2470 10440 2485
rect 10390 2450 10405 2470
rect 10425 2450 10440 2470
rect 10390 2420 10440 2450
rect 10390 2400 10405 2420
rect 10425 2400 10440 2420
rect 10390 2370 10440 2400
rect 10390 2350 10405 2370
rect 10425 2350 10440 2370
rect 10390 2320 10440 2350
rect 10390 2300 10405 2320
rect 10425 2300 10440 2320
rect 10390 2285 10440 2300
rect 10500 2470 10550 2485
rect 10500 2450 10515 2470
rect 10535 2450 10550 2470
rect 10500 2420 10550 2450
rect 10500 2400 10515 2420
rect 10535 2400 10550 2420
rect 10500 2370 10550 2400
rect 10500 2350 10515 2370
rect 10535 2350 10550 2370
rect 10500 2320 10550 2350
rect 10500 2300 10515 2320
rect 10535 2300 10550 2320
rect 10500 2285 10550 2300
rect 10610 2470 10660 2485
rect 10610 2450 10625 2470
rect 10645 2450 10660 2470
rect 10610 2420 10660 2450
rect 10610 2400 10625 2420
rect 10645 2400 10660 2420
rect 10610 2370 10660 2400
rect 10610 2350 10625 2370
rect 10645 2350 10660 2370
rect 10610 2320 10660 2350
rect 10610 2300 10625 2320
rect 10645 2300 10660 2320
rect 10610 2285 10660 2300
rect 10720 2470 10770 2485
rect 10720 2450 10735 2470
rect 10755 2450 10770 2470
rect 10720 2420 10770 2450
rect 10720 2400 10735 2420
rect 10755 2400 10770 2420
rect 10720 2370 10770 2400
rect 10720 2350 10735 2370
rect 10755 2350 10770 2370
rect 10720 2320 10770 2350
rect 10720 2300 10735 2320
rect 10755 2300 10770 2320
rect 10720 2285 10770 2300
<< ndiffc >>
rect 9215 1970 9235 1990
rect 9215 1920 9235 1940
rect 9215 1870 9235 1890
rect 9215 1820 9235 1840
rect 9325 1970 9345 1990
rect 9325 1920 9345 1940
rect 9325 1870 9345 1890
rect 9325 1820 9345 1840
rect 9435 1970 9455 1990
rect 9435 1920 9455 1940
rect 9435 1870 9455 1890
rect 9435 1820 9455 1840
rect 9545 1970 9565 1990
rect 9545 1920 9565 1940
rect 9545 1870 9565 1890
rect 9545 1820 9565 1840
rect 9655 1970 9675 1990
rect 9755 1970 9775 1990
rect 9655 1920 9675 1940
rect 9755 1920 9775 1940
rect 9655 1870 9675 1890
rect 9755 1870 9775 1890
rect 9655 1820 9675 1840
rect 9755 1820 9775 1840
rect 9865 1970 9885 1990
rect 9865 1920 9885 1940
rect 9865 1870 9885 1890
rect 9865 1820 9885 1840
rect 9975 1970 9995 1990
rect 9975 1920 9995 1940
rect 9975 1870 9995 1890
rect 9975 1820 9995 1840
rect 10085 1970 10105 1990
rect 10085 1920 10105 1940
rect 10085 1870 10105 1890
rect 10085 1820 10105 1840
rect 10195 1970 10215 1990
rect 10295 1970 10315 1990
rect 10195 1920 10215 1940
rect 10295 1920 10315 1940
rect 10195 1870 10215 1890
rect 10295 1870 10315 1890
rect 10195 1820 10215 1840
rect 10295 1820 10315 1840
rect 10405 1970 10425 1990
rect 10405 1920 10425 1940
rect 10405 1870 10425 1890
rect 10405 1820 10425 1840
rect 10515 1970 10535 1990
rect 10515 1920 10535 1940
rect 10515 1870 10535 1890
rect 10515 1820 10535 1840
rect 10625 1970 10645 1990
rect 10625 1920 10645 1940
rect 10625 1870 10645 1890
rect 10625 1820 10645 1840
rect 10735 1970 10755 1990
rect 10735 1920 10755 1940
rect 10735 1870 10755 1890
rect 10735 1820 10755 1840
<< pdiffc >>
rect 9315 2450 9335 2470
rect 9315 2400 9335 2420
rect 9315 2350 9335 2370
rect 9315 2300 9335 2320
rect 9425 2450 9445 2470
rect 9425 2400 9445 2420
rect 9425 2350 9445 2370
rect 9425 2300 9445 2320
rect 9535 2450 9555 2470
rect 9535 2400 9555 2420
rect 9535 2350 9555 2370
rect 9535 2300 9555 2320
rect 9645 2450 9665 2470
rect 9645 2400 9665 2420
rect 9645 2350 9665 2370
rect 9645 2300 9665 2320
rect 9755 2450 9775 2470
rect 9755 2400 9775 2420
rect 9755 2350 9775 2370
rect 9755 2300 9775 2320
rect 9865 2450 9885 2470
rect 9865 2400 9885 2420
rect 9865 2350 9885 2370
rect 9865 2300 9885 2320
rect 9975 2450 9995 2470
rect 10075 2450 10095 2470
rect 9975 2400 9995 2420
rect 10075 2400 10095 2420
rect 9975 2350 9995 2370
rect 10075 2350 10095 2370
rect 9975 2300 9995 2320
rect 10075 2300 10095 2320
rect 10185 2450 10205 2470
rect 10185 2400 10205 2420
rect 10185 2350 10205 2370
rect 10185 2300 10205 2320
rect 10295 2450 10315 2470
rect 10295 2400 10315 2420
rect 10295 2350 10315 2370
rect 10295 2300 10315 2320
rect 10405 2450 10425 2470
rect 10405 2400 10425 2420
rect 10405 2350 10425 2370
rect 10405 2300 10425 2320
rect 10515 2450 10535 2470
rect 10515 2400 10535 2420
rect 10515 2350 10535 2370
rect 10515 2300 10535 2320
rect 10625 2450 10645 2470
rect 10625 2400 10645 2420
rect 10625 2350 10645 2370
rect 10625 2300 10645 2320
rect 10735 2450 10755 2470
rect 10735 2400 10755 2420
rect 10735 2350 10755 2370
rect 10735 2300 10755 2320
<< psubdiff >>
rect 9150 1990 9200 2005
rect 9150 1970 9165 1990
rect 9185 1970 9200 1990
rect 9150 1940 9200 1970
rect 9150 1920 9165 1940
rect 9185 1920 9200 1940
rect 9150 1890 9200 1920
rect 9150 1870 9165 1890
rect 9185 1870 9200 1890
rect 9150 1840 9200 1870
rect 9150 1820 9165 1840
rect 9185 1820 9200 1840
rect 9150 1805 9200 1820
rect 9690 1990 9740 2005
rect 9690 1970 9705 1990
rect 9725 1970 9740 1990
rect 9690 1940 9740 1970
rect 9690 1920 9705 1940
rect 9725 1920 9740 1940
rect 9690 1890 9740 1920
rect 9690 1870 9705 1890
rect 9725 1870 9740 1890
rect 9690 1840 9740 1870
rect 9690 1820 9705 1840
rect 9725 1820 9740 1840
rect 9690 1805 9740 1820
rect 10230 1990 10280 2005
rect 10230 1970 10245 1990
rect 10265 1970 10280 1990
rect 10230 1940 10280 1970
rect 10230 1920 10245 1940
rect 10265 1920 10280 1940
rect 10230 1890 10280 1920
rect 10230 1870 10245 1890
rect 10265 1870 10280 1890
rect 10230 1840 10280 1870
rect 10230 1820 10245 1840
rect 10265 1820 10280 1840
rect 10230 1805 10280 1820
rect 10770 1990 10820 2005
rect 10770 1970 10785 1990
rect 10805 1970 10820 1990
rect 10770 1940 10820 1970
rect 10770 1920 10785 1940
rect 10805 1920 10820 1940
rect 10770 1890 10820 1920
rect 10770 1870 10785 1890
rect 10805 1870 10820 1890
rect 10770 1840 10820 1870
rect 10770 1820 10785 1840
rect 10805 1820 10820 1840
rect 10770 1805 10820 1820
<< nsubdiff >>
rect 9250 2470 9300 2485
rect 9250 2450 9265 2470
rect 9285 2450 9300 2470
rect 9250 2420 9300 2450
rect 9250 2400 9265 2420
rect 9285 2400 9300 2420
rect 9250 2370 9300 2400
rect 9250 2350 9265 2370
rect 9285 2350 9300 2370
rect 9250 2320 9300 2350
rect 9250 2300 9265 2320
rect 9285 2300 9300 2320
rect 9250 2285 9300 2300
rect 10010 2470 10060 2485
rect 10010 2450 10025 2470
rect 10045 2450 10060 2470
rect 10010 2420 10060 2450
rect 10010 2400 10025 2420
rect 10045 2400 10060 2420
rect 10010 2370 10060 2400
rect 10010 2350 10025 2370
rect 10045 2350 10060 2370
rect 10010 2320 10060 2350
rect 10010 2300 10025 2320
rect 10045 2300 10060 2320
rect 10010 2285 10060 2300
rect 10770 2470 10820 2485
rect 10770 2450 10785 2470
rect 10805 2450 10820 2470
rect 10770 2420 10820 2450
rect 10770 2400 10785 2420
rect 10805 2400 10820 2420
rect 10770 2370 10820 2400
rect 10770 2350 10785 2370
rect 10805 2350 10820 2370
rect 10770 2320 10820 2350
rect 10770 2300 10785 2320
rect 10805 2300 10820 2320
rect 10770 2285 10820 2300
<< psubdiffcont >>
rect 9165 1970 9185 1990
rect 9165 1920 9185 1940
rect 9165 1870 9185 1890
rect 9165 1820 9185 1840
rect 9705 1970 9725 1990
rect 9705 1920 9725 1940
rect 9705 1870 9725 1890
rect 9705 1820 9725 1840
rect 10245 1970 10265 1990
rect 10245 1920 10265 1940
rect 10245 1870 10265 1890
rect 10245 1820 10265 1840
rect 10785 1970 10805 1990
rect 10785 1920 10805 1940
rect 10785 1870 10805 1890
rect 10785 1820 10805 1840
<< nsubdiffcont >>
rect 9265 2450 9285 2470
rect 9265 2400 9285 2420
rect 9265 2350 9285 2370
rect 9265 2300 9285 2320
rect 10025 2450 10045 2470
rect 10025 2400 10045 2420
rect 10025 2350 10045 2370
rect 10025 2300 10045 2320
rect 10785 2450 10805 2470
rect 10785 2400 10805 2420
rect 10785 2350 10805 2370
rect 10785 2300 10805 2320
<< poly >>
rect 9305 2530 9345 2540
rect 9305 2510 9315 2530
rect 9335 2515 9345 2530
rect 10725 2530 10765 2540
rect 10725 2515 10735 2530
rect 9335 2510 9410 2515
rect 9305 2500 9410 2510
rect 10660 2510 10735 2515
rect 10755 2510 10765 2530
rect 10660 2500 10765 2510
rect 9350 2485 9410 2500
rect 9460 2485 9520 2500
rect 9570 2485 9630 2500
rect 9680 2485 9740 2500
rect 9790 2485 9850 2500
rect 9900 2485 9960 2500
rect 10110 2485 10170 2500
rect 10220 2485 10280 2500
rect 10330 2485 10390 2500
rect 10440 2485 10500 2500
rect 10550 2485 10610 2500
rect 10660 2485 10720 2500
rect 9350 2270 9410 2285
rect 9460 2275 9520 2285
rect 9570 2275 9630 2285
rect 9680 2275 9740 2285
rect 9790 2275 9850 2285
rect 9460 2255 9850 2275
rect 9900 2275 9960 2285
rect 10110 2275 10170 2285
rect 9900 2260 10170 2275
rect 10220 2270 10280 2285
rect 10330 2270 10390 2285
rect 10440 2270 10500 2285
rect 10550 2270 10610 2285
rect 10660 2270 10720 2285
rect 10015 2240 10025 2260
rect 10045 2240 10055 2260
rect 10220 2255 10610 2270
rect 10015 2230 10055 2240
rect 10570 2245 10610 2255
rect 10570 2225 10580 2245
rect 10600 2225 10610 2245
rect 10570 2215 10610 2225
rect 9425 2115 9465 2125
rect 9425 2095 9435 2115
rect 9455 2095 9465 2115
rect 9425 2035 9465 2095
rect 10570 2065 10610 2075
rect 9695 2050 9735 2060
rect 9250 2005 9310 2020
rect 9360 2015 9530 2035
rect 9695 2030 9705 2050
rect 9725 2030 9735 2050
rect 10235 2050 10275 2060
rect 10235 2030 10245 2050
rect 10265 2030 10275 2050
rect 10570 2045 10580 2065
rect 10600 2045 10610 2065
rect 10570 2035 10610 2045
rect 9360 2005 9420 2015
rect 9470 2005 9530 2015
rect 9580 2015 9850 2030
rect 9580 2005 9640 2015
rect 9790 2005 9850 2015
rect 9900 2015 10070 2030
rect 9900 2005 9960 2015
rect 10010 2005 10070 2015
rect 10120 2015 10390 2030
rect 10120 2005 10180 2015
rect 10330 2005 10390 2015
rect 10440 2020 10610 2035
rect 10440 2005 10500 2020
rect 10550 2005 10610 2020
rect 10660 2005 10720 2020
rect 9250 1790 9310 1805
rect 9360 1790 9420 1805
rect 9205 1780 9310 1790
rect 9205 1760 9215 1780
rect 9235 1775 9310 1780
rect 9235 1760 9245 1775
rect 9205 1750 9245 1760
rect 9470 1765 9530 1805
rect 9580 1790 9640 1805
rect 9790 1790 9850 1805
rect 9900 1765 9960 1805
rect 10010 1790 10070 1805
rect 10120 1790 10180 1805
rect 10330 1790 10390 1805
rect 10440 1790 10500 1805
rect 10550 1790 10610 1805
rect 10660 1790 10720 1805
rect 10660 1780 10765 1790
rect 10660 1775 10735 1780
rect 9470 1750 9960 1765
rect 10725 1760 10735 1775
rect 10755 1760 10765 1780
rect 10725 1750 10765 1760
<< polycont >>
rect 9315 2510 9335 2530
rect 10735 2510 10755 2530
rect 10025 2240 10045 2260
rect 10580 2225 10600 2245
rect 9435 2095 9455 2115
rect 9705 2030 9725 2050
rect 10245 2030 10265 2050
rect 10580 2045 10600 2065
rect 9215 1760 9235 1780
rect 10735 1760 10755 1780
<< locali >>
rect 10890 3865 10945 3875
rect 10890 3830 10900 3865
rect 10935 3830 10945 3865
rect 10890 3820 10945 3830
rect 9150 2565 9180 2585
rect 9200 2565 9230 2585
rect 9250 2565 9280 2585
rect 9300 2565 9330 2585
rect 9350 2565 9380 2585
rect 9400 2565 9430 2585
rect 9450 2565 9480 2585
rect 9500 2565 9530 2585
rect 9550 2565 9580 2585
rect 9600 2565 9630 2585
rect 9650 2565 9680 2585
rect 9700 2565 9730 2585
rect 9750 2565 9780 2585
rect 9800 2565 9830 2585
rect 9850 2565 9880 2585
rect 9900 2565 9930 2585
rect 9950 2565 9980 2585
rect 10000 2565 10030 2585
rect 10050 2565 10080 2585
rect 10100 2565 10130 2585
rect 10150 2565 10180 2585
rect 10200 2565 10230 2585
rect 10250 2565 10280 2585
rect 10300 2565 10330 2585
rect 10350 2565 10380 2585
rect 10400 2565 10430 2585
rect 10450 2565 10480 2585
rect 10500 2565 10530 2585
rect 10550 2565 10580 2585
rect 10600 2565 10630 2585
rect 10650 2565 10680 2585
rect 10700 2565 10730 2585
rect 10750 2565 10765 2585
rect 9305 2530 9345 2565
rect 9305 2510 9315 2530
rect 9335 2510 9345 2530
rect 9305 2480 9345 2510
rect 9255 2470 9345 2480
rect 9255 2450 9265 2470
rect 9285 2450 9315 2470
rect 9335 2450 9345 2470
rect 9255 2420 9345 2450
rect 9255 2400 9265 2420
rect 9285 2400 9315 2420
rect 9335 2400 9345 2420
rect 9255 2370 9345 2400
rect 9255 2350 9265 2370
rect 9285 2350 9315 2370
rect 9335 2350 9345 2370
rect 9255 2320 9345 2350
rect 9255 2300 9265 2320
rect 9285 2300 9315 2320
rect 9335 2300 9345 2320
rect 9255 2290 9345 2300
rect 9415 2470 9455 2565
rect 9415 2450 9425 2470
rect 9445 2450 9455 2470
rect 9415 2420 9455 2450
rect 9415 2400 9425 2420
rect 9445 2400 9455 2420
rect 9415 2370 9455 2400
rect 9415 2350 9425 2370
rect 9445 2350 9455 2370
rect 9415 2320 9455 2350
rect 9415 2300 9425 2320
rect 9445 2300 9455 2320
rect 9415 2290 9455 2300
rect 9525 2470 9565 2480
rect 9525 2450 9535 2470
rect 9555 2450 9565 2470
rect 9525 2420 9565 2450
rect 9525 2400 9535 2420
rect 9555 2400 9565 2420
rect 9525 2370 9565 2400
rect 9525 2350 9535 2370
rect 9555 2350 9565 2370
rect 9525 2320 9565 2350
rect 9525 2300 9535 2320
rect 9555 2300 9565 2320
rect 9525 2270 9565 2300
rect 9635 2470 9675 2565
rect 9635 2450 9645 2470
rect 9665 2450 9675 2470
rect 9635 2420 9675 2450
rect 9635 2400 9645 2420
rect 9665 2400 9675 2420
rect 9635 2370 9675 2400
rect 9635 2350 9645 2370
rect 9665 2350 9675 2370
rect 9635 2320 9675 2350
rect 9635 2300 9645 2320
rect 9665 2300 9675 2320
rect 9635 2290 9675 2300
rect 9745 2470 9785 2480
rect 9745 2450 9755 2470
rect 9775 2450 9785 2470
rect 9745 2420 9785 2450
rect 9745 2400 9755 2420
rect 9775 2400 9785 2420
rect 9745 2370 9785 2400
rect 9745 2350 9755 2370
rect 9775 2350 9785 2370
rect 9745 2320 9785 2350
rect 9745 2300 9755 2320
rect 9775 2300 9785 2320
rect 9745 2270 9785 2300
rect 9855 2470 9895 2565
rect 10015 2480 10055 2565
rect 9855 2450 9865 2470
rect 9885 2450 9895 2470
rect 9855 2420 9895 2450
rect 9855 2400 9865 2420
rect 9885 2400 9895 2420
rect 9855 2370 9895 2400
rect 9855 2350 9865 2370
rect 9885 2350 9895 2370
rect 9855 2320 9895 2350
rect 9855 2300 9865 2320
rect 9885 2300 9895 2320
rect 9855 2290 9895 2300
rect 9965 2470 10105 2480
rect 9965 2450 9975 2470
rect 9995 2450 10025 2470
rect 10045 2450 10075 2470
rect 10095 2450 10105 2470
rect 9965 2420 10105 2450
rect 9965 2400 9975 2420
rect 9995 2400 10025 2420
rect 10045 2400 10075 2420
rect 10095 2400 10105 2420
rect 9965 2370 10105 2400
rect 9965 2350 9975 2370
rect 9995 2350 10025 2370
rect 10045 2350 10075 2370
rect 10095 2350 10105 2370
rect 9965 2320 10105 2350
rect 9965 2300 9975 2320
rect 9995 2300 10025 2320
rect 10045 2300 10075 2320
rect 10095 2300 10105 2320
rect 9965 2290 10105 2300
rect 10175 2470 10215 2565
rect 10175 2450 10185 2470
rect 10205 2450 10215 2470
rect 10175 2420 10215 2450
rect 10175 2400 10185 2420
rect 10205 2400 10215 2420
rect 10175 2370 10215 2400
rect 10175 2350 10185 2370
rect 10205 2350 10215 2370
rect 10175 2320 10215 2350
rect 10175 2300 10185 2320
rect 10205 2300 10215 2320
rect 10175 2290 10215 2300
rect 10285 2470 10325 2480
rect 10285 2450 10295 2470
rect 10315 2450 10325 2470
rect 10285 2420 10325 2450
rect 10285 2400 10295 2420
rect 10315 2400 10325 2420
rect 10285 2370 10325 2400
rect 10285 2350 10295 2370
rect 10315 2350 10325 2370
rect 10285 2320 10325 2350
rect 10285 2300 10295 2320
rect 10315 2300 10325 2320
rect 9525 2230 9785 2270
rect 10015 2260 10055 2290
rect 10015 2240 10025 2260
rect 10045 2240 10055 2260
rect 10015 2230 10055 2240
rect 10285 2270 10325 2300
rect 10395 2470 10435 2565
rect 10395 2450 10405 2470
rect 10425 2450 10435 2470
rect 10395 2420 10435 2450
rect 10395 2400 10405 2420
rect 10425 2400 10435 2420
rect 10395 2370 10435 2400
rect 10395 2350 10405 2370
rect 10425 2350 10435 2370
rect 10395 2320 10435 2350
rect 10395 2300 10405 2320
rect 10425 2300 10435 2320
rect 10395 2290 10435 2300
rect 10505 2470 10545 2480
rect 10505 2450 10515 2470
rect 10535 2450 10545 2470
rect 10505 2420 10545 2450
rect 10505 2400 10515 2420
rect 10535 2400 10545 2420
rect 10505 2370 10545 2400
rect 10505 2350 10515 2370
rect 10535 2350 10545 2370
rect 10505 2320 10545 2350
rect 10505 2300 10515 2320
rect 10535 2300 10545 2320
rect 10505 2270 10545 2300
rect 10615 2470 10655 2565
rect 10615 2450 10625 2470
rect 10645 2450 10655 2470
rect 10615 2420 10655 2450
rect 10615 2400 10625 2420
rect 10645 2400 10655 2420
rect 10615 2370 10655 2400
rect 10615 2350 10625 2370
rect 10645 2350 10655 2370
rect 10615 2320 10655 2350
rect 10615 2300 10625 2320
rect 10645 2300 10655 2320
rect 10615 2290 10655 2300
rect 10725 2530 10765 2565
rect 10725 2510 10735 2530
rect 10755 2510 10765 2530
rect 10725 2480 10765 2510
rect 10725 2470 10815 2480
rect 10725 2450 10735 2470
rect 10755 2450 10785 2470
rect 10805 2450 10815 2470
rect 10725 2420 10815 2450
rect 10725 2400 10735 2420
rect 10755 2400 10785 2420
rect 10805 2400 10815 2420
rect 10725 2370 10815 2400
rect 10725 2350 10735 2370
rect 10755 2350 10785 2370
rect 10805 2350 10815 2370
rect 10725 2320 10815 2350
rect 10725 2300 10735 2320
rect 10755 2300 10785 2320
rect 10805 2300 10815 2320
rect 10725 2290 10815 2300
rect 10285 2230 10545 2270
rect 10905 2260 10960 2270
rect 10905 2255 10915 2260
rect 9745 2165 9785 2230
rect 10505 2170 10545 2230
rect 10570 2245 10915 2255
rect 10570 2225 10580 2245
rect 10600 2225 10915 2245
rect 10950 2225 10960 2260
rect 10570 2215 10960 2225
rect 9745 2125 10005 2165
rect 9095 2115 9465 2125
rect 9095 2105 9435 2115
rect 9425 2095 9435 2105
rect 9455 2095 9465 2115
rect 9155 1990 9245 2000
rect 9155 1970 9165 1990
rect 9185 1970 9215 1990
rect 9235 1970 9245 1990
rect 9155 1940 9245 1970
rect 9155 1920 9165 1940
rect 9185 1920 9215 1940
rect 9235 1920 9245 1940
rect 9155 1890 9245 1920
rect 9155 1870 9165 1890
rect 9185 1870 9215 1890
rect 9235 1870 9245 1890
rect 9155 1840 9245 1870
rect 9155 1820 9165 1840
rect 9185 1820 9215 1840
rect 9235 1820 9245 1840
rect 9155 1810 9245 1820
rect 9205 1780 9245 1810
rect 9205 1760 9215 1780
rect 9235 1760 9245 1780
rect 9205 1735 9245 1760
rect 9315 1990 9355 2000
rect 9315 1970 9325 1990
rect 9345 1970 9355 1990
rect 9315 1940 9355 1970
rect 9315 1920 9325 1940
rect 9345 1920 9355 1940
rect 9315 1890 9355 1920
rect 9315 1870 9325 1890
rect 9345 1870 9355 1890
rect 9315 1840 9355 1870
rect 9315 1820 9325 1840
rect 9345 1820 9355 1840
rect 9315 1735 9355 1820
rect 9425 1990 9465 2095
rect 9695 2050 9735 2060
rect 9695 2030 9705 2050
rect 9725 2030 9735 2050
rect 9695 2000 9735 2030
rect 9425 1970 9435 1990
rect 9455 1970 9465 1990
rect 9425 1940 9465 1970
rect 9425 1920 9435 1940
rect 9455 1920 9465 1940
rect 9425 1890 9465 1920
rect 9425 1870 9435 1890
rect 9455 1870 9465 1890
rect 9425 1840 9465 1870
rect 9425 1820 9435 1840
rect 9455 1820 9465 1840
rect 9425 1810 9465 1820
rect 9535 1990 9575 2000
rect 9535 1970 9545 1990
rect 9565 1970 9575 1990
rect 9535 1940 9575 1970
rect 9535 1920 9545 1940
rect 9565 1920 9575 1940
rect 9535 1890 9575 1920
rect 9535 1870 9545 1890
rect 9565 1870 9575 1890
rect 9535 1840 9575 1870
rect 9535 1820 9545 1840
rect 9565 1820 9575 1840
rect 9535 1735 9575 1820
rect 9645 1990 9785 2000
rect 9645 1970 9655 1990
rect 9675 1970 9705 1990
rect 9725 1970 9755 1990
rect 9775 1970 9785 1990
rect 9645 1940 9785 1970
rect 9645 1920 9655 1940
rect 9675 1920 9705 1940
rect 9725 1920 9755 1940
rect 9775 1920 9785 1940
rect 9645 1890 9785 1920
rect 9645 1870 9655 1890
rect 9675 1870 9705 1890
rect 9725 1870 9755 1890
rect 9775 1870 9785 1890
rect 9645 1840 9785 1870
rect 9645 1820 9655 1840
rect 9675 1820 9705 1840
rect 9725 1820 9755 1840
rect 9775 1820 9785 1840
rect 9645 1810 9785 1820
rect 9855 1990 9895 2000
rect 9855 1970 9865 1990
rect 9885 1970 9895 1990
rect 9855 1940 9895 1970
rect 9855 1920 9865 1940
rect 9885 1920 9895 1940
rect 9855 1890 9895 1920
rect 9855 1870 9865 1890
rect 9885 1870 9895 1890
rect 9855 1840 9895 1870
rect 9855 1820 9865 1840
rect 9885 1820 9895 1840
rect 9695 1735 9735 1810
rect 9855 1735 9895 1820
rect 9965 1990 10005 2125
rect 10505 2130 10860 2170
rect 10235 2050 10275 2060
rect 10235 2030 10245 2050
rect 10265 2030 10275 2050
rect 10235 2000 10275 2030
rect 9965 1970 9975 1990
rect 9995 1970 10005 1990
rect 9965 1940 10005 1970
rect 9965 1920 9975 1940
rect 9995 1920 10005 1940
rect 9965 1890 10005 1920
rect 9965 1870 9975 1890
rect 9995 1870 10005 1890
rect 9965 1840 10005 1870
rect 9965 1820 9975 1840
rect 9995 1820 10005 1840
rect 9965 1810 10005 1820
rect 10075 1990 10115 2000
rect 10075 1970 10085 1990
rect 10105 1970 10115 1990
rect 10075 1940 10115 1970
rect 10075 1920 10085 1940
rect 10105 1920 10115 1940
rect 10075 1890 10115 1920
rect 10075 1870 10085 1890
rect 10105 1870 10115 1890
rect 10075 1840 10115 1870
rect 10075 1820 10085 1840
rect 10105 1820 10115 1840
rect 10075 1735 10115 1820
rect 10185 1990 10325 2000
rect 10185 1970 10195 1990
rect 10215 1970 10245 1990
rect 10265 1970 10295 1990
rect 10315 1970 10325 1990
rect 10185 1940 10325 1970
rect 10185 1920 10195 1940
rect 10215 1920 10245 1940
rect 10265 1920 10295 1940
rect 10315 1920 10325 1940
rect 10185 1890 10325 1920
rect 10185 1870 10195 1890
rect 10215 1870 10245 1890
rect 10265 1870 10295 1890
rect 10315 1870 10325 1890
rect 10185 1840 10325 1870
rect 10185 1820 10195 1840
rect 10215 1820 10245 1840
rect 10265 1820 10295 1840
rect 10315 1820 10325 1840
rect 10185 1810 10325 1820
rect 10395 1990 10435 2000
rect 10395 1970 10405 1990
rect 10425 1970 10435 1990
rect 10395 1940 10435 1970
rect 10395 1920 10405 1940
rect 10425 1920 10435 1940
rect 10395 1890 10435 1920
rect 10395 1870 10405 1890
rect 10425 1870 10435 1890
rect 10395 1840 10435 1870
rect 10395 1820 10405 1840
rect 10425 1820 10435 1840
rect 10235 1735 10275 1810
rect 10395 1735 10435 1820
rect 10505 1990 10545 2130
rect 10570 2065 10960 2075
rect 10570 2045 10580 2065
rect 10600 2045 10915 2065
rect 10570 2035 10915 2045
rect 10905 2030 10915 2035
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10505 1970 10515 1990
rect 10535 1970 10545 1990
rect 10505 1940 10545 1970
rect 10505 1920 10515 1940
rect 10535 1920 10545 1940
rect 10505 1890 10545 1920
rect 10505 1870 10515 1890
rect 10535 1870 10545 1890
rect 10505 1840 10545 1870
rect 10505 1820 10515 1840
rect 10535 1820 10545 1840
rect 10505 1810 10545 1820
rect 10615 1990 10655 2000
rect 10615 1970 10625 1990
rect 10645 1970 10655 1990
rect 10615 1940 10655 1970
rect 10615 1920 10625 1940
rect 10645 1920 10655 1940
rect 10615 1890 10655 1920
rect 10615 1870 10625 1890
rect 10645 1870 10655 1890
rect 10615 1840 10655 1870
rect 10615 1820 10625 1840
rect 10645 1820 10655 1840
rect 10615 1735 10655 1820
rect 10725 1990 10815 2000
rect 10725 1970 10735 1990
rect 10755 1970 10785 1990
rect 10805 1970 10815 1990
rect 10725 1940 10815 1970
rect 10725 1920 10735 1940
rect 10755 1920 10785 1940
rect 10805 1920 10815 1940
rect 10725 1890 10815 1920
rect 10725 1870 10735 1890
rect 10755 1870 10785 1890
rect 10805 1870 10815 1890
rect 10725 1840 10815 1870
rect 10725 1820 10735 1840
rect 10755 1820 10785 1840
rect 10805 1820 10815 1840
rect 10725 1810 10815 1820
rect 10725 1780 10765 1810
rect 10725 1760 10735 1780
rect 10755 1760 10765 1780
rect 10725 1735 10765 1760
rect 9155 1715 9185 1735
rect 9205 1715 9235 1735
rect 9255 1715 9285 1735
rect 9305 1715 9335 1735
rect 9355 1715 9385 1735
rect 9405 1715 9435 1735
rect 9455 1715 9485 1735
rect 9505 1715 9535 1735
rect 9555 1715 9585 1735
rect 9605 1715 9635 1735
rect 9655 1715 9685 1735
rect 9705 1715 9735 1735
rect 9755 1715 9785 1735
rect 9805 1715 9835 1735
rect 9855 1715 9885 1735
rect 9905 1715 9935 1735
rect 9955 1715 9985 1735
rect 10005 1715 10035 1735
rect 10055 1715 10085 1735
rect 10105 1715 10135 1735
rect 10155 1715 10185 1735
rect 10205 1715 10235 1735
rect 10255 1715 10285 1735
rect 10305 1715 10335 1735
rect 10355 1715 10385 1735
rect 10405 1715 10435 1735
rect 10455 1715 10485 1735
rect 10505 1715 10535 1735
rect 10555 1715 10585 1735
rect 10605 1715 10635 1735
rect 10655 1715 10685 1735
rect 10705 1715 10735 1735
rect 10755 1715 10765 1735
rect 10890 1560 10945 1570
rect 10890 1525 10900 1560
rect 10935 1525 10945 1560
rect 10890 1515 10945 1525
<< viali >>
rect 10900 3830 10935 3865
rect 9180 2565 9200 2585
rect 9230 2565 9250 2585
rect 9280 2565 9300 2585
rect 9330 2565 9350 2585
rect 9380 2565 9400 2585
rect 9430 2565 9450 2585
rect 9480 2565 9500 2585
rect 9530 2565 9550 2585
rect 9580 2565 9600 2585
rect 9630 2565 9650 2585
rect 9680 2565 9700 2585
rect 9730 2565 9750 2585
rect 9780 2565 9800 2585
rect 9830 2565 9850 2585
rect 9880 2565 9900 2585
rect 9930 2565 9950 2585
rect 9980 2565 10000 2585
rect 10030 2565 10050 2585
rect 10080 2565 10100 2585
rect 10130 2565 10150 2585
rect 10180 2565 10200 2585
rect 10230 2565 10250 2585
rect 10280 2565 10300 2585
rect 10330 2565 10350 2585
rect 10380 2565 10400 2585
rect 10430 2565 10450 2585
rect 10480 2565 10500 2585
rect 10530 2565 10550 2585
rect 10580 2565 10600 2585
rect 10630 2565 10650 2585
rect 10680 2565 10700 2585
rect 10730 2565 10750 2585
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
rect 9185 1715 9205 1735
rect 9235 1715 9255 1735
rect 9285 1715 9305 1735
rect 9335 1715 9355 1735
rect 9385 1715 9405 1735
rect 9435 1715 9455 1735
rect 9485 1715 9505 1735
rect 9535 1715 9555 1735
rect 9585 1715 9605 1735
rect 9635 1715 9655 1735
rect 9685 1715 9705 1735
rect 9735 1715 9755 1735
rect 9785 1715 9805 1735
rect 9835 1715 9855 1735
rect 9885 1715 9905 1735
rect 9935 1715 9955 1735
rect 9985 1715 10005 1735
rect 10035 1715 10055 1735
rect 10085 1715 10105 1735
rect 10135 1715 10155 1735
rect 10185 1715 10205 1735
rect 10235 1715 10255 1735
rect 10285 1715 10305 1735
rect 10335 1715 10355 1735
rect 10385 1715 10405 1735
rect 10435 1715 10455 1735
rect 10485 1715 10505 1735
rect 10535 1715 10555 1735
rect 10585 1715 10605 1735
rect 10635 1715 10655 1735
rect 10685 1715 10705 1735
rect 10735 1715 10755 1735
rect 10900 1525 10935 1560
<< metal1 >>
rect 9105 3865 10945 3875
rect 9105 3830 10900 3865
rect 10935 3830 10945 3865
rect 9105 3820 10945 3830
rect 9150 2585 10765 2595
rect 9150 2565 9180 2585
rect 9200 2565 9230 2585
rect 9250 2565 9280 2585
rect 9300 2565 9330 2585
rect 9350 2565 9380 2585
rect 9400 2565 9430 2585
rect 9450 2565 9480 2585
rect 9500 2565 9530 2585
rect 9550 2565 9580 2585
rect 9600 2565 9630 2585
rect 9650 2565 9680 2585
rect 9700 2565 9730 2585
rect 9750 2565 9780 2585
rect 9800 2565 9830 2585
rect 9850 2565 9880 2585
rect 9900 2565 9930 2585
rect 9950 2565 9980 2585
rect 10000 2565 10030 2585
rect 10050 2565 10080 2585
rect 10100 2565 10130 2585
rect 10150 2565 10180 2585
rect 10200 2565 10230 2585
rect 10250 2565 10280 2585
rect 10300 2565 10330 2585
rect 10350 2565 10380 2585
rect 10400 2565 10430 2585
rect 10450 2565 10480 2585
rect 10500 2565 10530 2585
rect 10550 2565 10580 2585
rect 10600 2565 10630 2585
rect 10650 2565 10680 2585
rect 10700 2565 10730 2585
rect 10750 2565 10765 2585
rect 9150 2555 10765 2565
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 9155 1735 10765 1745
rect 9155 1715 9185 1735
rect 9205 1715 9235 1735
rect 9255 1715 9285 1735
rect 9305 1715 9335 1735
rect 9355 1715 9385 1735
rect 9405 1715 9435 1735
rect 9455 1715 9485 1735
rect 9505 1715 9535 1735
rect 9555 1715 9585 1735
rect 9605 1715 9635 1735
rect 9655 1715 9685 1735
rect 9705 1715 9735 1735
rect 9755 1715 9785 1735
rect 9805 1715 9835 1735
rect 9855 1715 9885 1735
rect 9905 1715 9935 1735
rect 9955 1715 9985 1735
rect 10005 1715 10035 1735
rect 10055 1715 10085 1735
rect 10105 1715 10135 1735
rect 10155 1715 10185 1735
rect 10205 1715 10235 1735
rect 10255 1715 10285 1735
rect 10305 1715 10335 1735
rect 10355 1715 10385 1735
rect 10405 1715 10435 1735
rect 10455 1715 10485 1735
rect 10505 1715 10535 1735
rect 10555 1715 10585 1735
rect 10605 1715 10635 1735
rect 10655 1715 10685 1735
rect 10705 1715 10735 1735
rect 10755 1715 10765 1735
rect 9155 1705 10765 1715
rect 9105 1560 10945 1570
rect 9105 1525 10900 1560
rect 10935 1525 10945 1560
rect 9105 1515 10945 1525
<< via1 >>
rect 10900 3830 10935 3865
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
rect 10900 1525 10935 1560
<< metal2 >>
rect 10890 3865 10945 3875
rect 10890 3830 10900 3865
rect 10935 3830 10945 3865
rect 10890 3820 10945 3830
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10890 1560 10945 1570
rect 10890 1525 10900 1560
rect 10935 1525 10945 1560
rect 10890 1515 10945 1525
<< via2 >>
rect 10900 3830 10935 3865
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
rect 10900 1525 10935 1560
<< metal3 >>
rect 10890 3865 10945 3875
rect 10890 3830 10900 3865
rect 10935 3830 10945 3865
rect 10890 3820 10945 3830
rect 10890 2390 14620 3820
rect 10905 2260 10960 2270
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 2020 10960 2030
rect 10890 1570 14520 1900
rect 10890 1560 10945 1570
rect 10890 1525 10900 1560
rect 10935 1525 10945 1560
rect 10890 1515 10945 1525
<< via3 >>
rect 10915 2225 10950 2260
rect 10915 2030 10950 2065
<< mimcap >>
rect 10905 2450 14605 3805
rect 10905 2415 10915 2450
rect 10950 2415 14605 2450
rect 10905 2405 14605 2415
rect 10905 1875 14505 1885
rect 10905 1840 10915 1875
rect 10950 1840 14505 1875
rect 10905 1585 14505 1840
<< mimcapcontact >>
rect 10915 2415 10950 2450
rect 10915 1840 10950 1875
<< metal4 >>
rect 10905 2450 10960 2460
rect 10905 2415 10915 2450
rect 10950 2415 10960 2450
rect 10905 2260 10960 2415
rect 10905 2225 10915 2260
rect 10950 2225 10960 2260
rect 10905 2215 10960 2225
rect 10905 2065 10960 2075
rect 10905 2030 10915 2065
rect 10950 2030 10960 2065
rect 10905 1875 10960 2030
rect 10905 1840 10915 1875
rect 10950 1840 10960 1875
rect 10905 1830 10960 1840
<< labels >>
flabel locali 10545 2105 10545 2105 3 FreeSans 400 0 160 0 vout
port 4 e
flabel metal1 9155 1725 9155 1725 7 FreeSans 400 0 -200 0 GNDA
port 2 w
flabel metal1 9150 2575 9150 2575 7 FreeSans 400 0 -200 0 VDDA
port 1 w
flabel poly 10610 2020 10610 2020 3 FreeSans 400 0 200 0 DOWN_input
port 9 e
flabel poly 10610 2270 10610 2270 3 FreeSans 400 0 200 0 UP_input
port 8 e
flabel locali 9095 2115 9095 2115 7 FreeSans 400 0 -200 0 I_IN
port 7 w
flabel locali 10005 2150 10005 2150 3 FreeSans 400 0 200 0 x
port 3 e
flabel poly 9510 2255 9510 2255 5 FreeSans 400 0 0 -200 opamp_out
port 10 s
flabel metal1 9105 1540 9105 1540 7 FreeSans 400 0 -200 0 DOWN
port 6 w
flabel metal1 9105 3845 9105 3845 7 FreeSans 400 0 -200 0 UP_b
port 5 w
<< end >>
