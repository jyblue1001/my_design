* PEX produced on Mon Feb  3 06:17:36 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from current_starved_VCO_magic.ext - technology: sky130A

.subckt current_starved_VCO_magic VDDA V_OSC V_CONT GNDA
X0 a_636_n552.t1 V_CONT.t0 GNDA.t12 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 a_82_186.t1 a_50_n62.t2 V_OSC.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.16
X2 a_82_186.t2 GNDA.t14 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X3 GNDA.t11 V_CONT.t1 a_n746_764.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X4 a_636_n552.t2 a_604_n62.t2 a_50_n62.t1 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.16
X5 VDDA.t5 a_n746_764.t1 a_n746_764.t2 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X6 a_1190_n552.t2 V_OSC.t2 a_604_n62.t0 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.16
X7 a_82_n552.t0 a_50_n62.t3 V_OSC.t1 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.16
X8 a_1190_n552.t1 VDDA.t17 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X9 a_1190_n552.t0 V_CONT.t2 GNDA.t9 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X10 a_82_n552.t2 VDDA.t18 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X11 a_82_n552.t1 V_CONT.t3 GNDA.t8 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X12 a_636_186.t1 a_n746_764.t3 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X13 a_82_186.t0 a_n746_764.t4 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X14 a_636_186.t2 a_604_n62.t3 a_50_n62.t0 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.16
X15 a_1190_186.t2 V_OSC.t3 a_604_n62.t1 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.16
X16 a_1190_186.t1 a_n746_764.t5 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X17 a_636_186.t0 GNDA.t15 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X18 a_1190_186.t0 GNDA.t16 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X19 a_636_n552.t0 VDDA.t19 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
R0 V_CONT V_CONT.t1 570.367
R1 V_CONT.t1 V_CONT.n1 488.83
R2 V_CONT.n0 V_CONT.t2 486.271
R3 V_CONT.n1 V_CONT.t3 384.967
R4 V_CONT.n0 V_CONT.t0 384.967
R5 V_CONT.n1 V_CONT.n0 101.303
R6 GNDA.t7 GNDA.t10 2694.17
R7 GNDA.t13 GNDA.t2 2627.65
R8 GNDA.n2 GNDA.t4 1848.38
R9 GNDA.n5 GNDA.n2 1170
R10 GNDA.n3 GNDA.t14 1076.47
R11 GNDA.n2 GNDA.t6 779.266
R12 GNDA.n4 GNDA.n3 504.493
R13 GNDA.n4 GNDA.t16 491.64
R14 GNDA.n5 GNDA.n4 352.723
R15 GNDA.n8 GNDA.t3 264.067
R16 GNDA.n7 GNDA.t5 264.067
R17 GNDA.n1 GNDA.t1 254.768
R18 GNDA.n3 GNDA.t15 186.374
R19 GNDA.n9 GNDA.t11 127.15
R20 GNDA.n8 GNDA.t8 127.15
R21 GNDA.n7 GNDA.t12 127.15
R22 GNDA.n0 GNDA.t9 127.15
R23 GNDA.n5 GNDA.n1 14.8842
R24 GNDA.n1 GNDA.n0 9.3005
R25 GNDA.n6 GNDA.n5 9.3005
R26 GNDA.t6 GNDA.t0 4.75212
R27 GNDA.t4 GNDA.t13 4.75212
R28 GNDA.t2 GNDA.t7 4.75212
R29 GNDA.n8 GNDA.n7 0.192861
R30 GNDA.n7 GNDA.n6 0.158139
R31 GNDA.n9 GNDA.n8 0.152583
R32 GNDA GNDA.n9 0.063
R33 GNDA.n6 GNDA.n0 0.0352222
R34 a_636_n552.n0 a_636_n552.t2 289.967
R35 a_636_n552.n0 a_636_n552.t0 254.768
R36 a_636_n552.t1 a_636_n552.n0 161.701
R37 a_50_n62.n1 a_50_n62.n0 785.028
R38 a_50_n62.t0 a_50_n62.n1 374.728
R39 a_50_n62.n1 a_50_n62.t1 271.567
R40 a_50_n62.n0 a_50_n62.t2 186.775
R41 a_50_n62.n0 a_50_n62.t3 115.981
R42 V_OSC.n2 V_OSC.n0 2160.31
R43 V_OSC.n0 V_OSC.t0 374.728
R44 V_OSC.n0 V_OSC.t1 271.567
R45 V_OSC.n1 V_OSC.t3 199.686
R46 V_OSC.n2 V_OSC.n1 181.013
R47 V_OSC.n1 V_OSC.t2 128.893
R48 V_OSC V_OSC.n2 44.8005
R49 a_82_186.n0 a_82_186.t1 398.087
R50 a_82_186.t2 a_82_186.n0 349.767
R51 a_82_186.n0 a_82_186.t0 212.364
R52 VDDA.n2 VDDA.t17 1007.38
R53 VDDA.n3 VDDA.t18 618.567
R54 VDDA.t0 VDDA.t4 488.219
R55 VDDA.t12 VDDA.t2 480.288
R56 VDDA.n4 VDDA.n3 357.406
R57 VDDA.n0 VDDA.t11 354.445
R58 VDDA.n7 VDDA.t15 354.418
R59 VDDA.n4 VDDA.t13 349.767
R60 VDDA.n1 VDDA.t14 341.048
R61 VDDA.n3 VDDA.n2 308.481
R62 VDDA.n4 VDDA.n1 185
R63 VDDA.n9 VDDA.t5 143.486
R64 VDDA.n8 VDDA.t1 143.486
R65 VDDA.n6 VDDA.t9 143.486
R66 VDDA.n0 VDDA.t3 143.486
R67 VDDA.n1 VDDA.t8 139.239
R68 VDDA.n2 VDDA.t19 117.287
R69 VDDA.t2 VDDA.t16 7.05059
R70 VDDA.t8 VDDA.t7 7.05059
R71 VDDA.t6 VDDA.t0 7.05059
R72 VDDA.n5 VDDA.n4 2.32108
R73 VDDA.t16 VDDA.t10 0.881762
R74 VDDA.t7 VDDA.t12 0.881762
R75 VDDA.t14 VDDA.t6 0.881762
R76 VDDA.n5 VDDA.n0 0.0901819
R77 VDDA VDDA.n9 0.0875743
R78 VDDA.n7 VDDA.n6 0.0798344
R79 VDDA.n9 VDDA.n8 0.0302988
R80 VDDA.n8 VDDA.n7 0.0283638
R81 VDDA.n6 VDDA.n5 0.0189745
R82 a_n746_764.t0 a_n746_764.n2 466.82
R83 a_n746_764.n2 a_n746_764.t1 225.869
R84 a_n746_764.n2 a_n746_764.t2 225.786
R85 a_n746_764.t1 a_n746_764.n1 188.501
R86 a_n746_764.n0 a_n746_764.t5 188.501
R87 a_n746_764.n1 a_n746_764.n0 107.442
R88 a_n746_764.n1 a_n746_764.t4 81.0592
R89 a_n746_764.n0 a_n746_764.t3 81.0592
R90 a_604_n62.n1 a_604_n62.n0 791.453
R91 a_604_n62.t1 a_604_n62.n1 374.728
R92 a_604_n62.n1 a_604_n62.t0 271.567
R93 a_604_n62.n0 a_604_n62.t3 186.775
R94 a_604_n62.n0 a_604_n62.t2 115.981
R95 a_1190_n552.n0 a_1190_n552.t2 289.967
R96 a_1190_n552.n0 a_1190_n552.t1 254.768
R97 a_1190_n552.t0 a_1190_n552.n0 161.701
R98 a_82_n552.n0 a_82_n552.t0 289.967
R99 a_82_n552.n0 a_82_n552.t2 254.768
R100 a_82_n552.t1 a_82_n552.n0 161.701
R101 a_636_186.n0 a_636_186.t2 398.087
R102 a_636_186.t0 a_636_186.n0 349.767
R103 a_636_186.n0 a_636_186.t1 212.364
R104 a_1190_186.n0 a_1190_186.t2 398.087
R105 a_1190_186.t0 a_1190_186.n0 349.767
R106 a_1190_186.n0 a_1190_186.t1 212.364
C0 V_OSC V_CONT 0.453248f
C1 VDDA V_CONT 0.064418f
C2 VDDA V_OSC 0.257612f
C3 V_CONT GNDA 1.51368f
C4 V_OSC GNDA 1.87158f
C5 VDDA GNDA 9.996414f
C6 a_n746_764.t2 GNDA 0.153998f
C7 a_n746_764.t5 GNDA 0.465957f
C8 a_n746_764.t3 GNDA 0.365904f
C9 a_n746_764.n0 GNDA 0.27731f
C10 a_n746_764.t4 GNDA 0.365904f
C11 a_n746_764.n1 GNDA 0.276948f
C12 a_n746_764.t1 GNDA 0.518928f
C13 a_n746_764.n2 GNDA 0.237652f
C14 a_n746_764.t0 GNDA 0.137401f
C15 VDDA.t3 GNDA 0.022852f
C16 VDDA.n0 GNDA 0.320483f
C17 VDDA.t10 GNDA 0.19384f
C18 VDDA.t2 GNDA 0.193141f
C19 VDDA.t12 GNDA 0.190697f
C20 VDDA.t8 GNDA 0.057977f
C21 VDDA.t4 GNDA 0.444959f
C22 VDDA.t0 GNDA 0.196285f
C23 VDDA.t14 GNDA 0.135513f
C24 VDDA.n1 GNDA 0.184775f
C25 VDDA.n3 GNDA 0.015998f
C26 VDDA.n4 GNDA 0.023552f
C27 VDDA.n5 GNDA 0.108054f
C28 VDDA.t9 GNDA 0.022852f
C29 VDDA.n6 GNDA 0.135286f
C30 VDDA.n7 GNDA 0.117915f
C31 VDDA.t1 GNDA 0.022852f
C32 VDDA.n8 GNDA 0.086173f
C33 VDDA.t5 GNDA 0.022852f
C34 VDDA.n9 GNDA 0.150219f
.ends

