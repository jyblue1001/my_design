magic
tech sky130A
timestamp 1745563040
use sky130_fd_pr__rf_test_coil1  sky130_fd_pr__rf_test_coil1_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 0 1 7252 -1 0 7745
box -7252 -7252 7750 7252
use sky130_fd_pr__rf_test_coil2  sky130_fd_pr__rf_test_coil2_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 32420 0 1 13200
box -13250 -13250 13750 13250
use sky130_fd_pr__rf_test_coil3  sky130_fd_pr__rf_test_coil3_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 68804 0 1 18289
box -18254 -18254 18754 18254
<< end >>
