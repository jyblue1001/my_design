* NGSPICE file created from charge_pump_full.ext - technology: sky130A

.subckt charge_pump_8 w_n3090_1240# a_n2950_2110# a_n2790_310# a_n3050_2170# a_n1130_2170#
X0 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X1 a_n1130_2170# UP_input w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X2 a_n2790_310# DOWN_input a_n1130_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X3 w_n3090_1240# UP_input a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X4 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X5 DOWN_b w_n3090_1240# DOWN_b_b a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 DOWN_input DOWN_b a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X7 DOWN_b a_n2790_310# DOWN_b_b w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X8 a_n3050_2170# I_IN a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X9 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X10 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X11 UP_b UP w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X12 I_IN I_IN a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X13 a_n1130_2170# DOWN_input a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X14 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X15 UP_input UP_b a_n2950_2110# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X16 UP UP_PFD_b a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X17 a_n2790_310# I_IN I_IN a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X18 a_n2790_310# I_IN I_IN a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X19 UP_input UP w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X20 UP_PFD_b UP_PFD a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X21 a_n1130_2170# UP_input w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X22 I_IN I_IN a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X23 a_n2790_310# DOWN_PFD DOWN_b_b a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X24 DOWN_input DOWN I_IN a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X25 a_n1130_2170# UP_input w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X26 DOWN DOWN_b w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X27 w_n3090_1240# UP_input a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X28 a_n1130_2170# UP_input w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X29 UP_PFD_b UP_PFD w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X30 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X31 w_n3090_1240# DOWN_PFD DOWN_b_b w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X32 w_n3090_1240# UP_input a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X33 a_n2790_310# I_IN a_n3050_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X34 a_n3050_2170# a_n2950_2110# w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X35 UP UP_PFD_b w_n3090_1240# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X36 a_n2790_310# DOWN_input a_n1130_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X37 UP_input UP a_n2950_2110# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X38 DOWN DOWN_b a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X39 w_n3090_1240# a_n2950_2110# a_n3050_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X40 a_n3050_2170# I_IN a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X41 w_n3090_1240# UP_input a_n1130_2170# w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X42 UP_b UP a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X43 a_n1130_2170# DOWN_input a_n2790_310# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X44 DOWN_input DOWN_b I_IN w_n3090_1240# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X45 a_n2790_310# I_IN a_n3050_2170# a_n2790_310# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X46 UP_input UP_b sky130_fd_pr__cap_mim_m3_1 l=4.2 w=6
X47 DOWN_input DOWN sky130_fd_pr__cap_mim_m3_1 l=2.6 w=2.6
.ends

.subckt opamp_6_6 a_1630_200# a_3420_n350# a_1470_530# w_1980_260# a_2150_n350#
X0 a_3420_n350# n_right w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 w_1980_260# n_right a_3420_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X2 a_3420_n350# p_right a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 a_3420_n350# a_4140_1066# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 v_common_p p_bias w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X5 a_3420_n350# n_right w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 p_right p_left a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X7 w_1980_260# p_bias v_common_p w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X8 a_4140_1066# n_right a_2150_n350# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X9 a_2150_n350# p_right a_3420_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X10 a_2150_n350# p_left p_left a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X11 w_1980_260# p_bias p_bias w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X12 p_right a_1630_200# v_common_p w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 v_common_p a_1470_530# p_left w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X14 n_bias n_bias a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X15 w_1980_260# p_bias v_common_p w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X16 p_left a_1470_530# v_common_p w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X17 a_3420_n350# p_right a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X18 p_bias p_bias w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 v_common_p a_1630_200# p_right w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X20 p_left p_left a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X21 a_2150_n350# n_bias v_common_n a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X22 p_right a_4140_n1860# a_2150_n350# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X23 v_common_n a_1630_200# n_right a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X24 n_left n_left w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X25 v_common_p p_bias w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X26 n_right a_1630_200# v_common_n a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X27 w_1980_260# n_left n_right w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X28 v_common_n n_bias a_2150_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X29 v_common_n a_1470_530# n_left a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X30 n_right n_left w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X31 a_3420_n350# a_4140_n1860# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X32 p_bias p_bias w_1980_260# w_1980_260# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X33 w_1980_260# n_left n_left w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X34 a_2150_n350# p_right a_3420_n350# a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 p_bias n_bias a_2150_n350# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X36 w_1980_260# n_right a_3420_n350# w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X37 w_1980_260# p_bias p_bias w_1980_260# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X38 a_2150_n350# p_left p_right a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X39 n_left a_1470_530# v_common_n a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X40 a_2150_n350# n_bias n_bias a_2150_n350# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
.ends

**.subckt charge_pump_full
Xcharge_pump_8_0 VDDA li_1590_1640# GNDA a_n310_5360# VOUT charge_pump_8
Xopamp_6_6_0 VOUT li_1590_1640# a_n310_5360# VDDA GNDA opamp_6_6
**.ends

