magic
tech sky130A
timestamp 1740486491
<< psubdiff >>
rect 2605 245 2655 260
rect 2605 225 2620 245
rect 2640 225 2655 245
rect 2605 210 2655 225
<< psubdiffcont >>
rect 2620 225 2640 245
<< xpolycontact >>
rect 5595 295 5815 330
rect 6479 295 6699 330
<< xpolyres >>
rect 5815 295 6479 330
<< locali >>
rect 1115 320 1165 330
rect 1115 290 1125 320
rect 1155 290 1165 320
rect 5555 325 5595 330
rect 5555 300 5560 325
rect 5585 300 5595 325
rect 5555 295 5595 300
rect 6699 325 6739 330
rect 6699 300 6709 325
rect 6734 300 6739 325
rect 6699 295 6739 300
rect 1115 280 1165 290
rect 2605 245 2655 260
rect 2605 230 2620 245
rect 2475 225 2620 230
rect 2640 230 2655 245
rect 2640 225 2780 230
rect 2475 220 2780 225
rect 2475 185 2485 220
rect 2520 210 2735 220
rect 2520 185 2530 210
rect 2475 175 2530 185
rect 2725 185 2735 210
rect 2770 185 2780 220
rect 2725 175 2780 185
<< viali >>
rect 1125 290 1155 320
rect 5560 300 5585 325
rect 6709 300 6734 325
rect 2485 185 2520 220
rect 2735 185 2770 220
<< metal1 >>
rect 1115 325 5595 330
rect 1115 320 5560 325
rect 1115 290 1125 320
rect 1155 300 5560 320
rect 5585 300 5595 325
rect 1155 295 5595 300
rect 6698 325 9740 330
rect 6698 300 6709 325
rect 6734 320 9740 325
rect 6734 300 9700 320
rect 6698 295 9700 300
rect 1155 290 1165 295
rect 1115 280 1165 290
rect 9690 290 9700 295
rect 9730 290 9740 320
rect 9690 280 9740 290
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
<< via1 >>
rect 1125 290 1155 320
rect 9700 290 9730 320
rect 2485 185 2520 220
rect 2735 185 2770 220
<< metal2 >>
rect 1115 320 1165 330
rect 1115 290 1125 320
rect 1155 290 1165 320
rect 1115 280 1165 290
rect 9690 320 9740 330
rect 9690 290 9700 320
rect 9730 290 9740 320
rect 9690 280 9740 290
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
<< via2 >>
rect 1125 290 1155 320
rect 9700 290 9730 320
rect 2485 185 2520 220
rect 2735 185 2770 220
<< metal3 >>
rect 1115 320 1165 330
rect 1115 290 1125 320
rect 1155 290 1165 320
rect 1115 55 1165 290
rect 9690 320 9740 330
rect 9690 290 9700 320
rect 9730 290 9740 320
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 9690 55 9740 290
rect 1115 -6975 2545 55
rect 2710 -6975 9740 55
<< via3 >>
rect 2485 185 2520 220
rect 2735 185 2770 220
<< mimcap >>
rect 1130 30 2530 40
rect 1130 -5 2485 30
rect 2520 -5 2530 30
rect 1130 -6960 2530 -5
rect 2725 30 9725 40
rect 2725 -5 2735 30
rect 2770 -5 9725 30
rect 2725 -6960 9725 -5
<< mimcapcontact >>
rect 2485 -5 2520 30
rect 2735 -5 2770 30
<< metal4 >>
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 30 2530 185
rect 2475 -5 2485 30
rect 2520 -5 2530 30
rect 2475 -10 2530 -5
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 30 2780 185
rect 2725 -5 2735 30
rect 2770 -5 2780 30
rect 2725 -10 2780 -5
<< labels >>
flabel locali 2630 260 2630 260 1 FreeSans 800 0 0 400 GNDA
port 2 n
flabel metal1 8250 330 8250 330 1 FreeSans 800 0 0 400 R1_C1
flabel metal1 1465 330 1465 330 1 FreeSans 800 0 0 400 V_OUT
port 1 n
<< end >>
