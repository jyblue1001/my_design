* PEX produced on Tue Jul 15 03:25:46 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 GNDA.t216 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 bgr_0.V_TOP.t12 VDDA.t410 VDDA.t412 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X2 VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 GNDA.t128 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X4 two_stage_opamp_dummy_magic_0.VD1.t13 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.X.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X5 VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t25 VDDA.t84 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X7 VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 GNDA.t43 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 VOUT-.t4 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X9 VDDA.t57 bgr_0.V_TOP.t14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X10 VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 bgr_0.Vin+.t4 bgr_0.V_TOP.t15 VDDA.t419 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X12 VDDA.t293 two_stage_opamp_dummy_magic_0.Vb3.t8 two_stage_opamp_dummy_magic_0.VD3.t29 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X13 GNDA.t313 VDDA.t407 VDDA.t409 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X14 VDDA.t433 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t5 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X15 VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X18 two_stage_opamp_dummy_magic_0.VD2.t16 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.Y.t2 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X19 VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 bgr_0.1st_Vout_2.t3 bgr_0.V_CUR_REF_REG.t3 bgr_0.V_p_2.t4 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X21 VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 a_7460_23988.t0 bgr_0.Vin+.t0 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=6
X24 VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 two_stage_opamp_dummy_magic_0.V_err_gate.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X27 VDDA.t406 VDDA.t404 bgr_0.NFET_GATE_10uA.t4 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 VDDA.t403 VDDA.t401 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X29 GNDA.t68 a_6930_22564.t0 GNDA.t56 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X30 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 bgr_0.PFET_GATE_10uA.t10 VDDA.t224 VDDA.t223 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X31 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X32 GNDA.t312 GNDA.t309 GNDA.t311 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X33 VDDA.t61 bgr_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X34 VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 GNDA.t144 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_0.V_source.t27 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X36 VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 bgr_0.1st_Vout_2.t9 bgr_0.V_mir2.t17 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X41 VDDA.t421 bgr_0.V_TOP.t16 bgr_0.Vin-.t7 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X42 bgr_0.1st_Vout_1.t10 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X43 GNDA.t316 VDDA.t469 bgr_0.V_p_2.t10 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X44 VDDA.t291 two_stage_opamp_dummy_magic_0.Vb3.t9 two_stage_opamp_dummy_magic_0.VD3.t28 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X45 VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 bgr_0.cap_res2.t20 bgr_0.PFET_GATE_10uA.t6 GNDA.t121 sky130_fd_pr__res_high_po_0p35 l=2.05
X47 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_0.Y.t25 VDDA.t158 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X49 VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 two_stage_opamp_dummy_magic_0.V_source.t26 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X52 two_stage_opamp_dummy_magic_0.VD2.t3 VIN+.t0 two_stage_opamp_dummy_magic_0.V_source.t5 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X53 VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VDDA.t119 bgr_0.1st_Vout_1.t13 bgr_0.V_TOP.t4 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X56 GNDA.t97 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 two_stage_opamp_dummy_magic_0.err_amp_out.t4 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X57 GNDA.t118 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X58 bgr_0.V_TOP.t17 VDDA.t422 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 two_stage_opamp_dummy_magic_0.VD4.t11 VDDA.t398 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X61 GNDA.t308 GNDA.t306 bgr_0.NFET_GATE_10uA.t0 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X62 bgr_0.START_UP.t5 bgr_0.V_TOP.t18 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X63 VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 two_stage_opamp_dummy_magic_0.V_err_gate.t11 bgr_0.NFET_GATE_10uA.t6 GNDA.t214 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X65 bgr_0.1st_Vout_1.t8 bgr_0.Vin+.t7 bgr_0.V_p_1.t3 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X66 VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_0.X.t26 VDDA.t240 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X68 VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 bgr_0.1st_Vout_1.t14 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t395 VDDA.t397 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X71 bgr_0.V_TOP.t19 VDDA.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X73 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t392 VDDA.t394 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X74 VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VOUT-.t9 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t242 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X76 VOUT+.t5 a_5980_2720.t0 GNDA.t95 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X77 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 bgr_0.PFET_GATE_10uA.t12 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X78 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 VDDA.t380 VDDA.t382 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X79 two_stage_opamp_dummy_magic_0.VD2.t15 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.Y.t4 GNDA.t344 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X80 VDDA.t11 bgr_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X81 two_stage_opamp_dummy_magic_0.VD2.t14 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.Y.t6 GNDA.t345 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X82 VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 bgr_0.V_TOP.t20 VDDA.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 bgr_0.1st_Vout_2.t2 bgr_0.V_CUR_REF_REG.t4 bgr_0.V_p_2.t3 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X85 two_stage_opamp_dummy_magic_0.VD4.t31 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.VD4.t30 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X86 VOUT+.t9 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA.t110 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X87 VDDA.t454 two_stage_opamp_dummy_magic_0.Y.t27 VOUT+.t18 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X88 VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t289 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X90 VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VDDA.t437 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X92 two_stage_opamp_dummy_magic_0.V_err_gate.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X93 VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 VDDA.t19 two_stage_opamp_dummy_magic_0.V_err_gate.t15 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X95 two_stage_opamp_dummy_magic_0.V_err_p.t17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.err_amp_out.t9 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X96 GNDA.t337 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_0.V_source.t25 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X97 VOUT-.t17 a_14010_2720.t1 GNDA.t343 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X98 bgr_0.PFET_GATE_10uA.t5 bgr_0.1st_Vout_2.t13 VDDA.t179 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X99 GNDA.t305 GNDA.t303 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X100 two_stage_opamp_dummy_magic_0.VD1.t19 VIN-.t0 two_stage_opamp_dummy_magic_0.V_source.t37 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X101 VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 bgr_0.V_TOP.t21 VDDA.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 two_stage_opamp_dummy_magic_0.X.t28 GNDA.t142 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X104 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t352 GNDA.t351 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X105 VDDA.t391 VDDA.t389 GNDA.t314 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X106 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X107 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X108 VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t28 VDDA.t463 GNDA.t350 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X110 two_stage_opamp_dummy_magic_0.VD2.t4 VIN+.t1 two_stage_opamp_dummy_magic_0.V_source.t7 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X111 VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 two_stage_opamp_dummy_magic_0.V_source.t24 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X113 bgr_0.V_TOP.t22 VDDA.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 GNDA.t212 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X115 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 bgr_0.NFET_GATE_10uA.t8 GNDA.t210 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 two_stage_opamp_dummy_magic_0.VD4.t29 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.Y.t16 two_stage_opamp_dummy_magic_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 GNDA.t105 two_stage_opamp_dummy_magic_0.Y.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X118 VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 bgr_0.1st_Vout_2.t14 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 two_stage_opamp_dummy_magic_0.VD1.t12 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t10 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X128 VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 a_12530_23988.t0 bgr_0.Vin-.t0 GNDA.t4 sky130_fd_pr__res_xhigh_po_0p35 l=6
X130 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.Vb3.t11 VDDA.t287 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X131 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X132 VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 bgr_0.1st_Vout_2.t8 bgr_0.V_mir2.t18 VDDA.t228 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X135 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t186 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X136 VOUT-.t8 two_stage_opamp_dummy_magic_0.X.t29 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X137 two_stage_opamp_dummy_magic_0.VD2.t13 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t3 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X138 VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VDDA.t468 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X145 two_stage_opamp_dummy_magic_0.V_err_gate.t13 VDDA.t386 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X146 VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 bgr_0.1st_Vout_1.t15 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 bgr_0.V_mir1.t13 bgr_0.Vin-.t8 bgr_0.V_p_1.t9 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X151 bgr_0.V_mir1.t11 bgr_0.V_mir1.t10 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X152 two_stage_opamp_dummy_magic_0.V_err_p.t1 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X153 GNDA.t326 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA.t325 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X154 two_stage_opamp_dummy_magic_0.VD3.t26 two_stage_opamp_dummy_magic_0.Vb3.t12 VDDA.t285 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X155 GNDA.t342 a_7580_22380.t1 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=6
X156 two_stage_opamp_dummy_magic_0.V_p_mir.t1 VIN+.t2 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X157 two_stage_opamp_dummy_magic_0.VD1.t1 VIN-.t1 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X158 VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VDDA.t246 bgr_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_0.Vb1.t3 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X164 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 two_stage_opamp_dummy_magic_0.X.t30 GNDA.t141 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X165 VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 bgr_0.V_TOP.t23 VDDA.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VDDA.t385 VDDA.t383 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X168 two_stage_opamp_dummy_magic_0.VD2.t2 VIN+.t3 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X169 VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 two_stage_opamp_dummy_magic_0.V_source.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X172 GNDA.t37 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 VOUT+.t2 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X173 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 bgr_0.PFET_GATE_10uA.t15 VDDA.t115 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X174 a_5700_5524.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X175 VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 VDDA.t283 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD4.t8 VDDA.t282 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X178 VOUT+.t17 two_stage_opamp_dummy_magic_0.Y.t30 VDDA.t452 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X179 GNDA.t323 VDDA.t377 VDDA.t379 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X180 bgr_0.V_mir1.t16 bgr_0.Vin-.t9 bgr_0.V_p_1.t8 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X181 VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X184 bgr_0.START_UP.t4 bgr_0.V_TOP.t24 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X185 VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 bgr_0.PFET_GATE_10uA.t4 bgr_0.1st_Vout_2.t16 VDDA.t417 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X187 VDDA.t133 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t4 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X188 VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 two_stage_opamp_dummy_magic_0.VD1.t11 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.X.t15 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X190 VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 two_stage_opamp_dummy_magic_0.Vb2.t5 bgr_0.NFET_GATE_10uA.t9 GNDA.t208 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X194 VDDA.t281 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X195 GNDA.t206 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X196 VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_0.V_TOP.t25 VDDA.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 GNDA.t204 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X199 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.VD4.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X200 two_stage_opamp_dummy_magic_0.V_err_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t424 VDDA.t423 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X201 VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VOUT-.t7 two_stage_opamp_dummy_magic_0.X.t31 VDDA.t236 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X204 two_stage_opamp_dummy_magic_0.VD2.t12 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.Y.t9 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X205 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_0.Y.t31 GNDA.t338 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X206 VDDA.t279 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD4.t7 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X207 VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.Vb3.t16 VDDA.t277 VDDA.t276 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X212 VDDA.t74 bgr_0.V_TOP.t26 bgr_0.Vin+.t3 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X213 bgr_0.1st_Vout_2.t0 bgr_0.V_mir2.t19 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X214 VDDA.t458 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t10 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X215 VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14010_2720.t0 GNDA.t328 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X217 bgr_0.V_TOP.t1 bgr_0.1st_Vout_1.t16 VDDA.t88 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X218 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X219 bgr_0.V_CUR_REF_REG.t1 VDDA.t374 VDDA.t376 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X220 VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 bgr_0.PFET_GATE_10uA.t16 VDDA.t204 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X225 VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 GNDA.t174 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_0.V_p_mir.t3 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X227 VDDA.t120 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X228 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.VD3.t35 two_stage_opamp_dummy_magic_0.VD3.t34 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X229 two_stage_opamp_dummy_magic_0.VD1.t18 GNDA.t300 GNDA.t302 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X230 two_stage_opamp_dummy_magic_0.VD1.t15 VIN-.t2 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X231 VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 a_6810_23838.t0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t56 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X235 VDDA.t465 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X236 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 two_stage_opamp_dummy_magic_0.X.t33 GNDA.t91 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X237 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.VD4.t25 two_stage_opamp_dummy_magic_0.VD4.t24 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X238 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t129 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X239 bgr_0.Vin+.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 GNDA.t335 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X240 VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA.t297 GNDA.t299 GNDA.t298 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X243 VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 two_stage_opamp_dummy_magic_0.V_source.t21 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X247 bgr_0.Vin+.t2 bgr_0.V_TOP.t27 VDDA.t217 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X248 VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VDDA.t373 VDDA.t371 bgr_0.PFET_GATE_10uA.t9 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X250 VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 VDDA.t219 bgr_0.V_TOP.t28 bgr_0.Vin+.t1 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X252 VOUT+.t4 two_stage_opamp_dummy_magic_0.Y.t33 VDDA.t135 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X253 VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 a_5580_5524.t1 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t112 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X255 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X256 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t5 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X257 VDDA.t370 VDDA.t368 two_stage_opamp_dummy_magic_0.V_err_gate.t12 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X258 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 GNDA.t33 a_12410_22380.t0 GNDA.t32 sky130_fd_pr__res_xhigh_po_0p35 l=6
X260 GNDA.t202 bgr_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X261 VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 VDDA.t275 two_stage_opamp_dummy_magic_0.Vb3.t17 two_stage_opamp_dummy_magic_0.VD3.t24 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X264 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t94 sky130_fd_pr__res_high_po_1p41 l=1.41
X265 VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 bgr_0.cap_res1.t0 bgr_0.V_TOP.t13 GNDA.t341 sky130_fd_pr__res_high_po_0p35 l=2.05
X267 two_stage_opamp_dummy_magic_0.Vb3.t5 bgr_0.NFET_GATE_10uA.t13 GNDA.t200 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X268 bgr_0.V_mir2.t9 bgr_0.V_mir2.t8 VDDA.t147 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X269 VDDA.t367 VDDA.t365 bgr_0.V_TOP.t11 VDDA.t366 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X270 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X271 GNDA.t16 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 two_stage_opamp_dummy_magic_0.err_amp_out.t3 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X272 VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 two_stage_opamp_dummy_magic_0.VD1.t10 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.X.t14 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X275 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 bgr_0.V_TOP.t29 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X279 bgr_0.1st_Vout_2.t19 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 VOUT-.t15 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t439 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X281 VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 GNDA.t65 a_13060_22630.t0 GNDA.t64 sky130_fd_pr__res_xhigh_po_0p35 l=4
X283 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t22 VDDA.t107 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X284 VOUT-.t16 two_stage_opamp_dummy_magic_0.X.t35 VDDA.t441 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X285 VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 two_stage_opamp_dummy_magic_0.V_source.t30 two_stage_opamp_dummy_magic_0.Vb1.t1 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X287 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_0.Y.t34 GNDA.t327 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X288 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA.t6 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X289 VDDA.t364 VDDA.t362 GNDA.t324 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X290 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t19 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X291 bgr_0.1st_Vout_1.t19 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 two_stage_opamp_dummy_magic_0.X.t22 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.VD3.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X293 VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VDDA.t273 two_stage_opamp_dummy_magic_0.Vb3.t18 two_stage_opamp_dummy_magic_0.VD3.t23 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X295 bgr_0.NFET_GATE_10uA.t1 bgr_0.PFET_GATE_10uA.t17 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X296 VDDA.t59 two_stage_opamp_dummy_magic_0.V_err_gate.t23 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X297 VDDA.t443 bgr_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X298 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.VD4.t23 two_stage_opamp_dummy_magic_0.VD4.t22 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X299 VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 GNDA.t170 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 VOUT-.t10 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X303 bgr_0.V_p_2.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 bgr_0.V_mir2.t16 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X304 VDDA.t446 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t332 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X305 VDDA.t213 bgr_0.V_TOP.t30 bgr_0.START_UP.t3 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X306 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t3 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X307 VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 a_5700_5524.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA.t340 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X311 VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 bgr_0.V_TOP.t31 VDDA.t214 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 bgr_0.V_TOP.t7 bgr_0.1st_Vout_1.t21 VDDA.t250 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X315 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 two_stage_opamp_dummy_magic_0.X.t37 GNDA.t333 VDDA.t447 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X316 VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t271 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X318 two_stage_opamp_dummy_magic_0.VD2.t17 VIN+.t4 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X319 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X320 GNDA.t296 GNDA.t294 VOUT-.t12 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X321 VOUT+.t1 two_stage_opamp_dummy_magic_0.Y.t35 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X322 VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 bgr_0.V_TOP.t5 bgr_0.1st_Vout_1.t22 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X325 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X326 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t19 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X327 VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 bgr_0.NFET_GATE_10uA.t3 bgr_0.NFET_GATE_10uA.t2 GNDA.t198 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X331 GNDA.t196 bgr_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X332 VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 bgr_0.V_TOP.t32 VDDA.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 VDDA.t361 VDDA.t359 VDDA.t361 VDDA.t360 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X335 GNDA.t293 GNDA.t291 two_stage_opamp_dummy_magic_0.VD1.t17 GNDA.t292 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X336 two_stage_opamp_dummy_magic_0.VD1.t9 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X337 two_stage_opamp_dummy_magic_0.VD4.t21 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.VD4.t20 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X338 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VDDA.t75 two_stage_opamp_dummy_magic_0.Y.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X342 VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.Vb3.t20 VDDA.t269 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X345 VOUT-.t14 VDDA.t356 VDDA.t358 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X346 VDDA.t449 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X347 VDDA.t355 VDDA.t353 two_stage_opamp_dummy_magic_0.VD3.t31 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X348 VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 GNDA.t290 GNDA.t288 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X350 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GNDA.t287 GNDA.t285 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X352 bgr_0.V_mir1.t9 bgr_0.V_mir1.t8 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X353 VDDA.t53 bgr_0.V_TOP.t33 bgr_0.START_UP.t2 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X354 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X355 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t37 GNDA.t107 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X356 VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 a_7460_23988.t1 a_7580_22380.t0 GNDA.t44 sky130_fd_pr__res_xhigh_po_0p35 l=6
X361 bgr_0.V_p_2.t2 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t5 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X362 VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X365 two_stage_opamp_dummy_magic_0.err_amp_out.t1 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 GNDA.t70 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X366 two_stage_opamp_dummy_magic_0.X.t16 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.VD1.t8 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X367 VDDA.t42 two_stage_opamp_dummy_magic_0.X.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X368 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.Y.t19 two_stage_opamp_dummy_magic_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X370 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t8 bgr_0.V_p_1.t2 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X371 VDDA.t189 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t7 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X372 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_0.X.t39 GNDA.t39 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X373 VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 GNDA.t221 GNDA.t284 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X377 VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X380 GNDA.t194 bgr_0.NFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X381 two_stage_opamp_dummy_magic_0.Vb2.t1 bgr_0.NFET_GATE_10uA.t16 GNDA.t192 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X382 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t281 GNDA.t283 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X383 VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 GNDA.t221 GNDA.t280 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X385 GNDA.t279 GNDA.t277 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t278 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X386 GNDA.t276 GNDA.t274 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X387 VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 bgr_0.PFET_GATE_10uA.t8 VDDA.t350 VDDA.t352 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X390 two_stage_opamp_dummy_magic_0.VD3.t22 two_stage_opamp_dummy_magic_0.Vb3.t21 VDDA.t267 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X391 VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 bgr_0.1st_Vout_1.t2 bgr_0.V_mir1.t20 VDDA.t31 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X393 VOUT+.t7 two_stage_opamp_dummy_magic_0.Y.t38 VDDA.t156 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X394 two_stage_opamp_dummy_magic_0.Vb2_2.t9 two_stage_opamp_dummy_magic_0.Vb2.t27 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X395 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t4 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X396 VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 VOUT-.t11 GNDA.t271 GNDA.t273 GNDA.t272 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X398 two_stage_opamp_dummy_magic_0.err_amp_out.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 two_stage_opamp_dummy_magic_0.V_err_p.t14 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X399 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.Vb3.t22 VDDA.t265 VDDA.t264 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X400 two_stage_opamp_dummy_magic_0.V_source.t20 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X401 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X402 bgr_0.V_p_2.t1 bgr_0.V_CUR_REF_REG.t6 bgr_0.1st_Vout_2.t4 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X403 VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 GNDA.t221 GNDA.t263 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X406 two_stage_opamp_dummy_magic_0.V_source.t34 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t16 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X407 VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 GNDA.t221 GNDA.t264 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X410 VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VDDA.t222 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X412 GNDA.t176 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X413 VDDA.t163 bgr_0.V_mir2.t6 bgr_0.V_mir2.t7 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X414 two_stage_opamp_dummy_magic_0.V_source.t9 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X415 GNDA.t331 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X416 VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA.t99 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X420 VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t40 GNDA.t117 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X422 bgr_0.V_p_2.t0 bgr_0.V_CUR_REF_REG.t7 bgr_0.1st_Vout_2.t1 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X423 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.Y.t0 two_stage_opamp_dummy_magic_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X424 VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 a_13180_23838.t0 bgr_0.V_CUR_REF_REG.t0 GNDA.t93 sky130_fd_pr__res_xhigh_po_0p35 l=4
X426 VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 bgr_0.V_TOP.t34 VDDA.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VDDA.t26 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X433 VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 bgr_0.V_TOP.t35 VDDA.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 a_5580_5524.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t63 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X437 VDDA.t27 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X438 VDDA.t263 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD4.t3 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X439 VDDA.t233 bgr_0.1st_Vout_2.t24 bgr_0.PFET_GATE_10uA.t3 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X440 VDDA.t349 VDDA.t347 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X441 VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t344 VDDA.t346 VDDA.t345 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X443 VDDA.t7 two_stage_opamp_dummy_magic_0.X.t42 VOUT-.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X444 VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 VDDA.t343 VDDA.t341 VOUT-.t13 VDDA.t342 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X446 VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 bgr_0.PFET_GATE_10uA.t20 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X450 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X451 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X452 VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VDDA.t83 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X455 VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 VOUT+.t0 two_stage_opamp_dummy_magic_0.Y.t41 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X457 VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t2 GNDA.t51 sky130_fd_pr__res_high_po_1p41 l=1.41
X459 VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 bgr_0.V_TOP.t36 VDDA.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 two_stage_opamp_dummy_magic_0.V_err_p.t8 two_stage_opamp_dummy_magic_0.V_err_gate.t24 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X462 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t9 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X463 VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_p.t0 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X465 bgr_0.Vin-.t6 bgr_0.V_TOP.t37 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X466 two_stage_opamp_dummy_magic_0.V_source.t17 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X467 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X468 VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VDDA.t340 VDDA.t337 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X470 VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 a_14170_5524.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t120 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X472 VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 VDDA.t261 two_stage_opamp_dummy_magic_0.Vb3.t24 two_stage_opamp_dummy_magic_0.VD4.t2 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X474 VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 GNDA.t190 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA.t189 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X476 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t49 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X477 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA.t268 GNDA.t270 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X478 VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 GNDA.t81 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 VOUT+.t3 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X483 VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VDDA.t182 two_stage_opamp_dummy_magic_0.Y.t42 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X486 two_stage_opamp_dummy_magic_0.V_source.t36 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X487 VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 GNDA.t168 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X489 two_stage_opamp_dummy_magic_0.V_source.t28 VIN+.t7 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X490 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA.t265 GNDA.t267 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X491 VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VDDA.t259 two_stage_opamp_dummy_magic_0.Vb3.t25 two_stage_opamp_dummy_magic_0.VD4.t1 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X497 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 bgr_0.PFET_GATE_10uA.t22 VDDA.t202 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X498 VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 bgr_0.V_TOP.t38 VDDA.t128 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X500 VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 GNDA.t262 GNDA.t260 VOUT+.t13 GNDA.t261 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X502 VDDA.t33 bgr_0.V_mir2.t4 bgr_0.V_mir2.t5 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X503 VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 VDDA.t41 bgr_0.V_mir1.t6 bgr_0.V_mir1.t7 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X505 VDDA.t200 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X506 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.VD1.t7 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X507 bgr_0.V_p_1.t7 bgr_0.Vin-.t10 bgr_0.V_mir1.t14 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X508 VDDA.t297 GNDA.t257 GNDA.t259 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X509 two_stage_opamp_dummy_magic_0.Vb2.t8 two_stage_opamp_dummy_magic_0.Vb2_2.t4 two_stage_opamp_dummy_magic_0.Vb2_2.t6 two_stage_opamp_dummy_magic_0.Vb2_2.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X510 VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 bgr_0.1st_Vout_1.t27 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 bgr_0.1st_Vout_2.t26 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 VDDA.t103 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X515 VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 VDDA.t9 two_stage_opamp_dummy_magic_0.X.t43 VOUT-.t1 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X517 two_stage_opamp_dummy_magic_0.Y.t11 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X518 bgr_0.V_TOP.t10 VDDA.t334 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X519 VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VDDA.t333 VDDA.t331 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X523 VDDA.t330 VDDA.t328 two_stage_opamp_dummy_magic_0.Vb2_2.t0 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X524 a_14290_5524.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t339 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X525 VOUT+.t15 VDDA.t325 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X526 VDDA.t324 VDDA.t322 two_stage_opamp_dummy_magic_0.VD4.t10 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X527 bgr_0.V_p_1.t6 bgr_0.Vin-.t11 bgr_0.V_mir1.t15 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X528 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t8 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X529 VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t92 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X532 VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA.t254 GNDA.t256 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X537 VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 two_stage_opamp_dummy_magic_0.err_amp_out.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 two_stage_opamp_dummy_magic_0.V_err_p.t16 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X539 bgr_0.Vin-.t2 bgr_0.START_UP.t6 bgr_0.V_TOP.t6 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X540 two_stage_opamp_dummy_magic_0.V_source.t15 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X541 bgr_0.V_TOP.t3 bgr_0.START_UP.t7 bgr_0.Vin-.t1 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X542 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 VIN-.t5 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X543 two_stage_opamp_dummy_magic_0.V_source.t39 VIN-.t6 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t347 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X544 VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VDDA.t37 bgr_0.1st_Vout_2.t27 bgr_0.PFET_GATE_10uA.t2 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X548 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t117 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X549 VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 GNDA.t134 two_stage_opamp_dummy_magic_0.X.t44 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X552 VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 GNDA.t221 GNDA.t222 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X554 bgr_0.START_UP.t1 bgr_0.START_UP.t0 bgr_0.START_UP_NFET1.t0 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X555 bgr_0.V_p_2.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 bgr_0.V_mir2.t15 GNDA.t353 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X556 VDDA.t0 two_stage_opamp_dummy_magic_0.Y.t43 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X557 two_stage_opamp_dummy_magic_0.V_source.t2 VIN+.t8 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X558 GNDA.t166 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X559 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_0.Y.t44 GNDA.t115 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X560 VDDA.t428 two_stage_opamp_dummy_magic_0.Y.t45 VOUT+.t16 VDDA.t427 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X561 VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 VDDA.t111 bgr_0.PFET_GATE_10uA.t24 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X568 GNDA.t356 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 two_stage_opamp_dummy_magic_0.V_source.t13 GNDA.t355 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X569 VDDA.t152 bgr_0.V_mir2.t21 bgr_0.1st_Vout_2.t6 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X570 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 bgr_0.PFET_GATE_10uA.t25 VDDA.t81 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X571 VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 bgr_0.V_p_1.t5 bgr_0.Vin-.t12 bgr_0.V_mir1.t12 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X573 two_stage_opamp_dummy_magic_0.VD4.t0 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X574 GNDA.t221 GNDA.t253 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X575 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD1.t6 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X576 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 VOUT+.t12 GNDA.t250 GNDA.t252 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X581 VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 bgr_0.1st_Vout_1.t30 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 GNDA.t227 GNDA.t226 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X585 VDDA.t86 two_stage_opamp_dummy_magic_0.V_err_gate.t27 two_stage_opamp_dummy_magic_0.V_err_p.t6 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X586 VDDA.t198 two_stage_opamp_dummy_magic_0.X.t45 VOUT-.t6 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X587 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X588 a_6810_23838.t1 a_6930_22564.t1 GNDA.t56 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X589 VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X590 GNDA.t221 GNDA.t220 bgr_0.Vin-.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X591 VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 VDDA.t255 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD3.t21 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X594 VOUT+.t10 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA.t137 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X595 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 two_stage_opamp_dummy_magic_0.V_err_gate.t28 VDDA.t139 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X596 VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 GNDA.t188 bgr_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X598 bgr_0.Vin-.t5 bgr_0.V_TOP.t39 VDDA.t66 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X599 two_stage_opamp_dummy_magic_0.err_amp_out.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_p.t13 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X600 a_14290_5524.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA.t119 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X601 a_12530_23988.t1 a_12410_22380.t1 GNDA.t161 sky130_fd_pr__res_xhigh_po_0p35 l=6
X602 two_stage_opamp_dummy_magic_0.Vb3.t7 bgr_0.NFET_GATE_10uA.t19 GNDA.t186 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X603 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_0.X.t46 VDDA.t108 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X605 two_stage_opamp_dummy_magic_0.V_source.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t148 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X606 GNDA.t249 GNDA.t247 VDDA.t296 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X607 two_stage_opamp_dummy_magic_0.V_source.t8 VIN-.t7 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X608 VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 VDDA.t141 bgr_0.V_mir2.t2 bgr_0.V_mir2.t3 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X610 VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 bgr_0.1st_Vout_1.t31 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 bgr_0.1st_Vout_2.t32 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 bgr_0.V_p_1.t10 VDDA.t470 GNDA.t318 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X614 GNDA.t86 two_stage_opamp_dummy_magic_0.X.t47 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X615 VDDA.t69 two_stage_opamp_dummy_magic_0.Y.t46 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X616 VDDA.t321 VDDA.t319 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X617 VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X618 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 bgr_0.PFET_GATE_10uA.t26 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X619 VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 two_stage_opamp_dummy_magic_0.V_source.t38 VIN+.t9 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA.t346 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X622 GNDA.t124 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X623 a_13180_23838.t1 a_13060_22630.t1 GNDA.t139 sky130_fd_pr__res_xhigh_po_0p35 l=4
X624 VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 VDDA.t173 two_stage_opamp_dummy_magic_0.Y.t47 VOUT+.t8 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X628 VDDA.t318 VDDA.t316 VOUT+.t14 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X629 bgr_0.V_p_1.t1 bgr_0.Vin+.t9 bgr_0.1st_Vout_1.t6 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X630 VDDA.t51 bgr_0.V_mir1.t22 bgr_0.1st_Vout_1.t0 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X631 two_stage_opamp_dummy_magic_0.V_err_gate.t0 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X632 bgr_0.V_TOP.t40 VDDA.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 two_stage_opamp_dummy_magic_0.Vb2_2.t8 two_stage_opamp_dummy_magic_0.Vb2.t9 two_stage_opamp_dummy_magic_0.Vb2.t10 two_stage_opamp_dummy_magic_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X634 VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 GNDA.t31 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X638 two_stage_opamp_dummy_magic_0.X.t21 GNDA.t244 GNDA.t246 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X639 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X640 VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 VDDA.t105 two_stage_opamp_dummy_magic_0.V_err_gate.t29 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X642 VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 VDDA.t194 two_stage_opamp_dummy_magic_0.X.t48 VOUT-.t5 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X645 bgr_0.V_TOP.t41 VDDA.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 a_14170_5524.t0 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t104 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X647 bgr_0.V_p_1.t0 bgr_0.Vin+.t10 bgr_0.1st_Vout_1.t9 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X648 VDDA.t315 VDDA.t313 bgr_0.V_TOP.t9 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X649 two_stage_opamp_dummy_magic_0.Y.t13 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X650 VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 two_stage_opamp_dummy_magic_0.Vb2.t0 bgr_0.NFET_GATE_10uA.t20 GNDA.t184 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X652 GNDA.t182 bgr_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X653 GNDA.t240 GNDA.t238 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X654 GNDA.t354 two_stage_opamp_dummy_magic_0.Y.t48 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X655 VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 bgr_0.NFET_GATE_10uA.t22 GNDA.t180 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X658 bgr_0.V_TOP.t42 VDDA.t169 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X660 bgr_0.V_TOP.t43 VDDA.t170 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 two_stage_opamp_dummy_magic_0.V_err_p.t5 two_stage_opamp_dummy_magic_0.V_err_gate.t30 VDDA.t456 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X663 VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 VDDA.t248 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t10 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X665 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.Y.t18 two_stage_opamp_dummy_magic_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X666 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 VDDA.t310 VDDA.t312 VDDA.t311 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X667 VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 VDDA.t39 bgr_0.1st_Vout_1.t32 bgr_0.V_TOP.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X669 VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X671 VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 two_stage_opamp_dummy_magic_0.X.t49 VDDA.t195 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X674 two_stage_opamp_dummy_magic_0.V_source.t31 VIN-.t8 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X675 VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 two_stage_opamp_dummy_magic_0.V_err_p.t4 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t461 VDDA.t460 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X677 GNDA.t23 two_stage_opamp_dummy_magic_0.X.t50 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X678 bgr_0.V_TOP.t44 VDDA.t171 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VDDA.t295 GNDA.t235 GNDA.t237 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X680 two_stage_opamp_dummy_magic_0.VD3.t30 VDDA.t307 VDDA.t309 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X681 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5980_2720.t1 GNDA.t113 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X682 VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VOUT-.t18 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA.t358 GNDA.t357 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X684 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X685 bgr_0.V_TOP.t45 VDDA.t206 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 bgr_0.V_mir2.t1 bgr_0.V_mir2.t0 VDDA.t414 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X687 VDDA.t226 bgr_0.V_mir1.t2 bgr_0.V_mir1.t3 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X688 VDDA.t211 two_stage_opamp_dummy_magic_0.Y.t49 VOUT+.t11 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X689 VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 two_stage_opamp_dummy_magic_0.V_err_gate.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X692 VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 bgr_0.V_mir2.t14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 bgr_0.V_p_2.t6 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X694 VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 bgr_0.PFET_GATE_10uA.t7 VDDA.t471 GNDA.t319 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X697 two_stage_opamp_dummy_magic_0.err_amp_out.t10 GNDA.t232 GNDA.t234 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X698 VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X700 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD1.t4 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X701 VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_0.Vb1.t0 bgr_0.PFET_GATE_10uA.t27 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X703 VDDA.t208 bgr_0.V_TOP.t46 bgr_0.Vin-.t4 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X704 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_0.Y.t50 VDDA.t450 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X705 VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 VOUT-.t3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X707 VDDA.t137 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X708 VDDA.t22 two_stage_opamp_dummy_magic_0.X.t51 VOUT-.t2 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X709 VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 bgr_0.PFET_GATE_10uA.t1 bgr_0.1st_Vout_2.t33 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X711 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.Vb3.t28 VDDA.t253 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X712 VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 VDDA.t431 bgr_0.PFET_GATE_10uA.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t430 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X714 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t304 VDDA.t306 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X715 GNDA.t72 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t0 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X716 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X717 VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 GNDA.t349 two_stage_opamp_dummy_magic_0.Y.t51 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t462 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X719 VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 VDDA.t426 bgr_0.1st_Vout_2.t34 bgr_0.PFET_GATE_10uA.t0 VDDA.t425 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X722 VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t435 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X725 VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 GNDA.t231 GNDA.t229 two_stage_opamp_dummy_magic_0.X.t20 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X730 VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 bgr_0.V_mir2.t13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 bgr_0.V_p_2.t8 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X732 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t76 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X733 two_stage_opamp_dummy_magic_0.V_source.t29 VIN-.t9 two_stage_opamp_dummy_magic_0.VD1.t3 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X734 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 bgr_0.NFET_GATE_10uA.t23 GNDA.t178 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X735 GNDA.t58 two_stage_opamp_dummy_magic_0.X.t53 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X736 VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X738 GNDA.t221 GNDA.t228 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X739 VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 GNDA.t108 two_stage_opamp_dummy_magic_0.X.t54 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X741 VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 VDDA.t90 bgr_0.1st_Vout_1.t36 bgr_0.V_TOP.t2 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X745 GNDA.t225 GNDA.t223 two_stage_opamp_dummy_magic_0.Y.t12 GNDA.t224 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X746 GNDA.t322 VDDA.t472 bgr_0.V_TOP.t8 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X747 bgr_0.V_TOP.t47 VDDA.t209 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 VDDA.t167 bgr_0.V_TOP.t48 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X750 VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X752 VDDA.t154 two_stage_opamp_dummy_magic_0.Y.t52 VOUT+.t6 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X753 VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 two_stage_opamp_dummy_magic_0.Vb2_2.t3 two_stage_opamp_dummy_magic_0.Vb2_2.t1 two_stage_opamp_dummy_magic_0.Vb2_2.t3 two_stage_opamp_dummy_magic_0.Vb2_2.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X756 two_stage_opamp_dummy_magic_0.Y.t24 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X757 VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 two_stage_opamp_dummy_magic_0.V_err_gate.t1 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X759 bgr_0.V_mir2.t12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 bgr_0.V_p_2.t9 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X760 two_stage_opamp_dummy_magic_0.V_err_p.t15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t5 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X761 VDDA.t303 VDDA.t301 two_stage_opamp_dummy_magic_0.err_amp_out.t11 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X762 VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 VDDA.t445 bgr_0.PFET_GATE_10uA.t29 bgr_0.V_CUR_REF_REG.t2 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X764 VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 two_stage_opamp_dummy_magic_0.VD1.t21 VIN-.t10 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA.t348 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X768 VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X773 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 two_stage_opamp_dummy_magic_0.Y.t53 VDDA.t180 GNDA.t114 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X774 GNDA.t219 GNDA.t217 VDDA.t294 GNDA.t218 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X775 two_stage_opamp_dummy_magic_0.V_source.t10 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t164 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X776 bgr_0.V_TOP.t49 VDDA.t168 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X777 two_stage_opamp_dummy_magic_0.VD2.t0 VIN+.t10 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X778 two_stage_opamp_dummy_magic_0.V_source.t0 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X779 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 VDDA.t298 VDDA.t300 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X780 two_stage_opamp_dummy_magic_0.Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X781 two_stage_opamp_dummy_magic_0.X.t19 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X782 VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X784 VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 bgr_0.1st_Vout_2.t36 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 GNDA.t151 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X788 GNDA.t53 two_stage_opamp_dummy_magic_0.Y.t54 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X789 VDDA.t47 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X790 VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 two_stage_opamp_dummy_magic_0.Y.t20 two_stage_opamp_dummy_magic_0.Vb2.t32 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X792 VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t2 384.967
R1 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t10 369.534
R2 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t22 369.534
R3 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t7 369.534
R4 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t16 369.534
R5 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t12 369.534
R6 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.n18 369.534
R7 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 366.553
R8 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t9 192.8
R9 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t17 192.8
R10 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t23 192.8
R11 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t11 192.8
R12 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t20 192.8
R13 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t21 192.8
R14 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t8 192.8
R15 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t15 192.8
R16 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t19 192.8
R17 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t5 192.8
R18 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t13 192.8
R19 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t18 192.8
R20 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t6 192.8
R21 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t14 192.8
R22 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R23 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R24 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R25 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R26 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R27 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R28 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R29 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R30 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R31 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R32 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R33 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R34 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R35 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R36 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R37 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R38 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R39 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R40 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 39.4005
R41 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t1 39.4005
R42 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 30.6442
R43 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t0 24.0005
R44 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t3 24.0005
R45 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t14 650.511
R46 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t13 611.739
R47 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t22 611.739
R48 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t8 611.739
R49 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t16 611.739
R50 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R51 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R52 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t26 421.75
R53 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.t25 421.75
R54 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R55 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t20 421.75
R56 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R57 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R58 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t11 421.75
R59 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R60 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t21 421.75
R61 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R62 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R63 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t12 421.75
R64 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R65 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R66 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 176.185
R67 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n14 175.624
R68 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R69 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R70 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 167.094
R71 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R72 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R73 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.n17 167.094
R74 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R75 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R76 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 167.094
R77 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R78 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R79 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.n8 167.094
R80 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n5 161.631
R81 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n0 139.639
R82 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.n1 139.638
R83 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 134.577
R84 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 49.8072
R85 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n18 49.8072
R86 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n13 49.8072
R87 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.n9 49.8072
R88 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 48.0943
R89 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 41.063
R90 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R91 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R92 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R93 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R94 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R95 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R96 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.n24 13.7349
R97 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t0 11.2576
R98 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t2 11.2576
R99 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n2 4.5005
R100 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 1.438
R101 GNDA.n2426 GNDA.n2111 21305.6
R102 GNDA.n2437 GNDA.n35 21305.6
R103 GNDA.n2433 GNDA.n2109 16744.4
R104 GNDA.n2434 GNDA.n2433 16744.4
R105 GNDA.n2104 GNDA.n39 15367.3
R106 GNDA.n2431 GNDA.n2429 13534.7
R107 GNDA.n2430 GNDA.n2108 13528.5
R108 GNDA.n2433 GNDA.n2432 13200
R109 GNDA.n2427 GNDA.n2110 13120
R110 GNDA.n2437 GNDA.n34 13120
R111 GNDA.n2237 GNDA.n2236 12825.5
R112 GNDA.n2237 GNDA.n2235 12823.6
R113 GNDA.n2106 GNDA.n2105 12810.6
R114 GNDA.n2435 GNDA.n2434 12017.1
R115 GNDA.n2104 GNDA.n2103 11953.3
R116 GNDA.n2103 GNDA.n41 11890.5
R117 GNDA.n2428 GNDA.n2109 11270.3
R118 GNDA.n2432 GNDA.n2108 11178.4
R119 GNDA.n41 GNDA.n40 9950.42
R120 GNDA.n2105 GNDA.n2104 9950.42
R121 GNDA.n2435 GNDA.n2108 9632.43
R122 GNDA.n2105 GNDA.n37 9384.59
R123 GNDA.n40 GNDA.n37 9384.59
R124 GNDA.n2436 GNDA.n2435 9001.83
R125 GNDA.n2107 GNDA.n38 7427.52
R126 GNDA.n2431 GNDA.n2430 4761.61
R127 GNDA.n109 GNDA.n41 4448.89
R128 GNDA.n2103 GNDA.n2102 3974.19
R129 GNDA.n2432 GNDA.n2431 3961.87
R130 GNDA.t94 GNDA.n2436 3375.81
R131 GNDA.n2107 GNDA.n37 3105.87
R132 GNDA.n2235 GNDA.n2111 2882.18
R133 GNDA.n2236 GNDA.n35 2858
R134 GNDA.n2236 GNDA.n34 2417.58
R135 GNDA.n2235 GNDA.n2110 2393.41
R136 GNDA.n2436 GNDA.n2107 2321.1
R137 GNDA.n2430 GNDA.n2107 2315.79
R138 GNDA.n2378 GNDA.n2237 2200
R139 GNDA.n2426 GNDA.t104 2006.86
R140 GNDA.n2436 GNDA.n36 2001.83
R141 GNDA.n2429 GNDA.n2107 1779.93
R142 GNDA.n2106 GNDA.n39 1460.18
R143 GNDA.n40 GNDA.n38 1440.71
R144 GNDA.n38 GNDA.n36 1440.71
R145 GNDA.n1857 GNDA.n1856 1336.64
R146 GNDA.t315 GNDA.n109 1258.74
R147 GNDA.n341 GNDA.n219 1214.72
R148 GNDA.n342 GNDA.n341 1214.72
R149 GNDA.n342 GNDA.n334 1214.72
R150 GNDA.n348 GNDA.n334 1214.72
R151 GNDA.n348 GNDA.n151 1214.72
R152 GNDA.n355 GNDA.n150 1214.72
R153 GNDA.n355 GNDA.n327 1214.72
R154 GNDA.n361 GNDA.n327 1214.72
R155 GNDA.n362 GNDA.n361 1214.72
R156 GNDA.n362 GNDA.n149 1214.72
R157 GNDA.n1963 GNDA.n1962 1212.88
R158 GNDA.n2076 GNDA.n2075 1185.07
R159 GNDA.n2075 GNDA.n69 1185.07
R160 GNDA.n2361 GNDA.n2360 1182.8
R161 GNDA.n2346 GNDA.n2345 1182.8
R162 GNDA.n2107 GNDA.n2106 1167.58
R163 GNDA.t341 GNDA.n39 1012.83
R164 GNDA.n2428 GNDA.n2427 984.414
R165 GNDA.n2427 GNDA.t51 896.639
R166 GNDA.n109 GNDA.n36 869.924
R167 GNDA.t221 GNDA.n151 823.313
R168 GNDA.n2334 GNDA.n2111 808.163
R169 GNDA.n2366 GNDA.n35 808.163
R170 GNDA.n2412 GNDA.t257 762.534
R171 GNDA.n2414 GNDA.t247 762.534
R172 GNDA.n2551 GNDA.t217 762.534
R173 GNDA.n15 GNDA.t235 762.534
R174 GNDA.t51 GNDA.n2426 702.521
R175 GNDA.n2451 GNDA.n2450 692.506
R176 GNDA.n2547 GNDA.n2546 692.506
R177 GNDA.n2408 GNDA.n2407 692.506
R178 GNDA.n2424 GNDA.n2423 692.506
R179 GNDA.n2495 GNDA.n2494 692.506
R180 GNDA.n2535 GNDA.n2534 692.506
R181 GNDA.n2216 GNDA.n2215 692.506
R182 GNDA.n2155 GNDA.n2152 692.506
R183 GNDA.n2072 GNDA.n2071 686.717
R184 GNDA.n2365 GNDA.n2364 686.717
R185 GNDA.n2376 GNDA.n2375 686.717
R186 GNDA.n2343 GNDA.n2342 686.717
R187 GNDA.n2333 GNDA.n2332 686.717
R188 GNDA.n1964 GNDA.n1963 686.717
R189 GNDA.n1964 GNDA.n110 686.717
R190 GNDA.n2226 GNDA.n2225 686.717
R191 GNDA.n2271 GNDA.n2270 686.717
R192 GNDA.n2383 GNDA.n2382 686.717
R193 GNDA.n2396 GNDA.n2395 686.717
R194 GNDA.n2281 GNDA.n2280 686.717
R195 GNDA.n2318 GNDA.n2317 686.717
R196 GNDA.n2321 GNDA.n2320 686.717
R197 GNDA.n2284 GNDA.n2283 686.717
R198 GNDA.n2063 GNDA.n77 686.717
R199 GNDA.n167 GNDA.n160 686.717
R200 GNDA.n2285 GNDA.t309 682.201
R201 GNDA.n211 GNDA.n208 669.307
R202 GNDA.n2322 GNDA.t285 650.067
R203 GNDA.n856 GNDA.n176 585.001
R204 GNDA.n1163 GNDA.n1162 585.001
R205 GNDA.n1157 GNDA.n1156 585.001
R206 GNDA.n1036 GNDA.n1035 585.001
R207 GNDA.n1030 GNDA.n1029 585.001
R208 GNDA.n1971 GNDA.n1970 585.001
R209 GNDA.n1256 GNDA.n1255 585
R210 GNDA.n1254 GNDA.n795 585
R211 GNDA.n1253 GNDA.n1252 585
R212 GNDA.n1251 GNDA.n1250 585
R213 GNDA.n1249 GNDA.n1248 585
R214 GNDA.n1247 GNDA.n1246 585
R215 GNDA.n1245 GNDA.n1244 585
R216 GNDA.n1243 GNDA.n1242 585
R217 GNDA.n1241 GNDA.n1240 585
R218 GNDA.n1239 GNDA.n1238 585
R219 GNDA.n1237 GNDA.n790 585
R220 GNDA.n1258 GNDA.n790 585
R221 GNDA.n1236 GNDA.n798 585
R222 GNDA.n1236 GNDA.n1235 585
R223 GNDA.n184 GNDA.n182 585
R224 GNDA.n592 GNDA.n591 585
R225 GNDA.n594 GNDA.n593 585
R226 GNDA.n596 GNDA.n595 585
R227 GNDA.n598 GNDA.n597 585
R228 GNDA.n600 GNDA.n599 585
R229 GNDA.n602 GNDA.n601 585
R230 GNDA.n604 GNDA.n603 585
R231 GNDA.n606 GNDA.n605 585
R232 GNDA.n608 GNDA.n607 585
R233 GNDA.n609 GNDA.n589 585
R234 GNDA.n1258 GNDA.n589 585
R235 GNDA.n610 GNDA.n590 585
R236 GNDA.n733 GNDA.n610 585
R237 GNDA.n1258 GNDA.n581 585
R238 GNDA.n770 GNDA.n769 585
R239 GNDA.n772 GNDA.n771 585
R240 GNDA.n774 GNDA.n773 585
R241 GNDA.n776 GNDA.n775 585
R242 GNDA.n778 GNDA.n777 585
R243 GNDA.n780 GNDA.n779 585
R244 GNDA.n782 GNDA.n781 585
R245 GNDA.n784 GNDA.n783 585
R246 GNDA.n785 GNDA.n739 585
R247 GNDA.n787 GNDA.n786 585
R248 GNDA.n583 GNDA.n582 585
R249 GNDA.n1781 GNDA.n1780 585
R250 GNDA.n1780 GNDA.n149 585
R251 GNDA.n363 GNDA.n325 585
R252 GNDA.n363 GNDA.n362 585
R253 GNDA.n359 GNDA.n326 585
R254 GNDA.n361 GNDA.n326 585
R255 GNDA.n358 GNDA.n357 585
R256 GNDA.n357 GNDA.n327 585
R257 GNDA.n356 GNDA.n329 585
R258 GNDA.n356 GNDA.n355 585
R259 GNDA.n352 GNDA.n330 585
R260 GNDA.n330 GNDA.n150 585
R261 GNDA.n351 GNDA.n350 585
R262 GNDA.n350 GNDA.n151 585
R263 GNDA.n349 GNDA.n332 585
R264 GNDA.n349 GNDA.n348 585
R265 GNDA.n345 GNDA.n333 585
R266 GNDA.n334 GNDA.n333 585
R267 GNDA.n344 GNDA.n343 585
R268 GNDA.n343 GNDA.n342 585
R269 GNDA.n339 GNDA.n336 585
R270 GNDA.n341 GNDA.n339 585
R271 GNDA.n338 GNDA.n337 585
R272 GNDA.n338 GNDA.n219 585
R273 GNDA.n337 GNDA.n221 585
R274 GNDA.n221 GNDA.n219 585
R275 GNDA.n340 GNDA.n336 585
R276 GNDA.n341 GNDA.n340 585
R277 GNDA.n344 GNDA.n335 585
R278 GNDA.n342 GNDA.n335 585
R279 GNDA.n346 GNDA.n345 585
R280 GNDA.n346 GNDA.n334 585
R281 GNDA.n347 GNDA.n332 585
R282 GNDA.n348 GNDA.n347 585
R283 GNDA.n351 GNDA.n331 585
R284 GNDA.n331 GNDA.n151 585
R285 GNDA.n353 GNDA.n352 585
R286 GNDA.n353 GNDA.n150 585
R287 GNDA.n354 GNDA.n329 585
R288 GNDA.n355 GNDA.n354 585
R289 GNDA.n358 GNDA.n328 585
R290 GNDA.n328 GNDA.n327 585
R291 GNDA.n360 GNDA.n359 585
R292 GNDA.n361 GNDA.n360 585
R293 GNDA.n325 GNDA.n324 585
R294 GNDA.n362 GNDA.n324 585
R295 GNDA.n1782 GNDA.n1781 585
R296 GNDA.n1782 GNDA.n149 585
R297 GNDA.n1696 GNDA.n513 585
R298 GNDA.n1699 GNDA.n1698 585
R299 GNDA.n1695 GNDA.n515 585
R300 GNDA.n1693 GNDA.n1692 585
R301 GNDA.n517 GNDA.n516 585
R302 GNDA.n1686 GNDA.n1685 585
R303 GNDA.n1683 GNDA.n519 585
R304 GNDA.n1681 GNDA.n1680 585
R305 GNDA.n521 GNDA.n520 585
R306 GNDA.n1674 GNDA.n1673 585
R307 GNDA.n1671 GNDA.n523 585
R308 GNDA.n1669 GNDA.n1668 585
R309 GNDA.n1668 GNDA.n1667 585
R310 GNDA.n523 GNDA.n522 585
R311 GNDA.n1675 GNDA.n1674 585
R312 GNDA.n1677 GNDA.n521 585
R313 GNDA.n1680 GNDA.n1679 585
R314 GNDA.n519 GNDA.n518 585
R315 GNDA.n1687 GNDA.n1686 585
R316 GNDA.n1689 GNDA.n517 585
R317 GNDA.n1692 GNDA.n1691 585
R318 GNDA.n515 GNDA.n514 585
R319 GNDA.n1700 GNDA.n1699 585
R320 GNDA.n1702 GNDA.n513 585
R321 GNDA.n747 GNDA.n479 585
R322 GNDA.n750 GNDA.n749 585
R323 GNDA.n752 GNDA.n751 585
R324 GNDA.n754 GNDA.n745 585
R325 GNDA.n756 GNDA.n755 585
R326 GNDA.n757 GNDA.n744 585
R327 GNDA.n759 GNDA.n758 585
R328 GNDA.n761 GNDA.n742 585
R329 GNDA.n763 GNDA.n762 585
R330 GNDA.n764 GNDA.n741 585
R331 GNDA.n766 GNDA.n765 585
R332 GNDA.n768 GNDA.n740 585
R333 GNDA.n551 GNDA.n524 585
R334 GNDA.n550 GNDA.n549 585
R335 GNDA.n547 GNDA.n525 585
R336 GNDA.n545 GNDA.n544 585
R337 GNDA.n543 GNDA.n526 585
R338 GNDA.n542 GNDA.n541 585
R339 GNDA.n539 GNDA.n527 585
R340 GNDA.n537 GNDA.n536 585
R341 GNDA.n535 GNDA.n528 585
R342 GNDA.n534 GNDA.n533 585
R343 GNDA.n531 GNDA.n529 585
R344 GNDA.n483 GNDA.n480 585
R345 GNDA.n1646 GNDA.n1645 585
R346 GNDA.n1647 GNDA.n560 585
R347 GNDA.n1649 GNDA.n1648 585
R348 GNDA.n1651 GNDA.n558 585
R349 GNDA.n1653 GNDA.n1652 585
R350 GNDA.n1654 GNDA.n557 585
R351 GNDA.n1656 GNDA.n1655 585
R352 GNDA.n1658 GNDA.n555 585
R353 GNDA.n1660 GNDA.n1659 585
R354 GNDA.n1661 GNDA.n554 585
R355 GNDA.n1663 GNDA.n1662 585
R356 GNDA.n1665 GNDA.n553 585
R357 GNDA.n732 GNDA.n731 585
R358 GNDA.n729 GNDA.n728 585
R359 GNDA.n727 GNDA.n726 585
R360 GNDA.n638 GNDA.n615 585
R361 GNDA.n643 GNDA.n642 585
R362 GNDA.n645 GNDA.n637 585
R363 GNDA.n648 GNDA.n647 585
R364 GNDA.n653 GNDA.n636 585
R365 GNDA.n659 GNDA.n658 585
R366 GNDA.n661 GNDA.n635 585
R367 GNDA.n666 GNDA.n665 585
R368 GNDA.n663 GNDA.n662 585
R369 GNDA.n1779 GNDA.n323 585
R370 GNDA.n1779 GNDA.n322 585
R371 GNDA.n1735 GNDA.n1734 585
R372 GNDA.n1736 GNDA.n377 585
R373 GNDA.n1746 GNDA.n1745 585
R374 GNDA.n1748 GNDA.n376 585
R375 GNDA.n1751 GNDA.n1750 585
R376 GNDA.n1752 GNDA.n372 585
R377 GNDA.n1761 GNDA.n1760 585
R378 GNDA.n1763 GNDA.n371 585
R379 GNDA.n1766 GNDA.n1765 585
R380 GNDA.n1767 GNDA.n365 585
R381 GNDA.n1776 GNDA.n1775 585
R382 GNDA.n1778 GNDA.n364 585
R383 GNDA.n1783 GNDA.n323 585
R384 GNDA.n1783 GNDA.n322 585
R385 GNDA.n1786 GNDA.n1785 585
R386 GNDA.n1787 GNDA.n258 585
R387 GNDA.n1797 GNDA.n1796 585
R388 GNDA.n1799 GNDA.n257 585
R389 GNDA.n1802 GNDA.n1801 585
R390 GNDA.n1803 GNDA.n253 585
R391 GNDA.n1812 GNDA.n1811 585
R392 GNDA.n1814 GNDA.n252 585
R393 GNDA.n1817 GNDA.n1816 585
R394 GNDA.n1818 GNDA.n246 585
R395 GNDA.n1827 GNDA.n1826 585
R396 GNDA.n1829 GNDA.n244 585
R397 GNDA.n233 GNDA.n232 585
R398 GNDA.n1857 GNDA.n233 585
R399 GNDA.n1860 GNDA.n1859 585
R400 GNDA.n1859 GNDA.n1858 585
R401 GNDA.n1861 GNDA.n231 585
R402 GNDA.n231 GNDA.n230 585
R403 GNDA.n1863 GNDA.n1862 585
R404 GNDA.n1864 GNDA.n1863 585
R405 GNDA.n229 GNDA.n228 585
R406 GNDA.n1865 GNDA.n229 585
R407 GNDA.n1868 GNDA.n1867 585
R408 GNDA.n1867 GNDA.n1866 585
R409 GNDA.n1869 GNDA.n227 585
R410 GNDA.n227 GNDA.n226 585
R411 GNDA.n1871 GNDA.n1870 585
R412 GNDA.n1872 GNDA.n1871 585
R413 GNDA.n225 GNDA.n224 585
R414 GNDA.n1873 GNDA.n225 585
R415 GNDA.n1876 GNDA.n1875 585
R416 GNDA.n1875 GNDA.n1874 585
R417 GNDA.n1877 GNDA.n222 585
R418 GNDA.n222 GNDA.n220 585
R419 GNDA.n1879 GNDA.n1878 585
R420 GNDA.n1880 GNDA.n1879 585
R421 GNDA.n213 GNDA.n212 585
R422 GNDA.n214 GNDA.n205 585
R423 GNDA.t221 GNDA.n214 585
R424 GNDA.n218 GNDA.n217 585
R425 GNDA.n1882 GNDA.n218 585
R426 GNDA.n1885 GNDA.n1884 585
R427 GNDA.n1884 GNDA.n1883 585
R428 GNDA.n1886 GNDA.n216 585
R429 GNDA.n216 GNDA.n215 585
R430 GNDA.n1888 GNDA.n1887 585
R431 GNDA.n1889 GNDA.n1888 585
R432 GNDA.n207 GNDA.n206 585
R433 GNDA.n1890 GNDA.n207 585
R434 GNDA.n1893 GNDA.n1892 585
R435 GNDA.n1892 GNDA.n1891 585
R436 GNDA.n1895 GNDA.n204 585
R437 GNDA.n204 GNDA.n203 585
R438 GNDA.n1897 GNDA.n1896 585
R439 GNDA.n1898 GNDA.n1897 585
R440 GNDA.n201 GNDA.n200 585
R441 GNDA.n1899 GNDA.n201 585
R442 GNDA.n1902 GNDA.n1901 585
R443 GNDA.n1901 GNDA.n1900 585
R444 GNDA.n1903 GNDA.n198 585
R445 GNDA.n202 GNDA.n198 585
R446 GNDA.n1905 GNDA.n1904 585
R447 GNDA.n1905 GNDA.n143 585
R448 GNDA.n1913 GNDA.n193 585
R449 GNDA.n1913 GNDA.n144 585
R450 GNDA.n1916 GNDA.n1915 585
R451 GNDA.n1915 GNDA.n1914 585
R452 GNDA.n1917 GNDA.n192 585
R453 GNDA.n192 GNDA.n191 585
R454 GNDA.n1919 GNDA.n1918 585
R455 GNDA.n1920 GNDA.n1919 585
R456 GNDA.n190 GNDA.n189 585
R457 GNDA.n1921 GNDA.n190 585
R458 GNDA.n1924 GNDA.n1923 585
R459 GNDA.n1923 GNDA.n1922 585
R460 GNDA.n1925 GNDA.n188 585
R461 GNDA.n188 GNDA.n187 585
R462 GNDA.n1927 GNDA.n1926 585
R463 GNDA.n1928 GNDA.n1927 585
R464 GNDA.n186 GNDA.n185 585
R465 GNDA.n1929 GNDA.n186 585
R466 GNDA.n1932 GNDA.n1931 585
R467 GNDA.n1931 GNDA.n1930 585
R468 GNDA.n1933 GNDA.n183 585
R469 GNDA.n183 GNDA.n181 585
R470 GNDA.n1935 GNDA.n1934 585
R471 GNDA.n1936 GNDA.n1935 585
R472 GNDA.n477 GNDA.n476 585
R473 GNDA.n475 GNDA.n444 585
R474 GNDA.n466 GNDA.n443 585
R475 GNDA.n469 GNDA.n468 585
R476 GNDA.n465 GNDA.n446 585
R477 GNDA.n463 GNDA.n462 585
R478 GNDA.n448 GNDA.n447 585
R479 GNDA.n456 GNDA.n455 585
R480 GNDA.n453 GNDA.n451 585
R481 GNDA.n196 GNDA.n195 585
R482 GNDA.n1910 GNDA.n1909 585
R483 GNDA.n1912 GNDA.n194 585
R484 GNDA.n1731 GNDA.n478 585
R485 GNDA.n478 GNDA.n322 585
R486 GNDA.n1906 GNDA.n194 585
R487 GNDA.n1909 GNDA.n1908 585
R488 GNDA.n197 GNDA.n196 585
R489 GNDA.n451 GNDA.n450 585
R490 GNDA.n457 GNDA.n456 585
R491 GNDA.n459 GNDA.n448 585
R492 GNDA.n462 GNDA.n461 585
R493 GNDA.n446 GNDA.n445 585
R494 GNDA.n470 GNDA.n469 585
R495 GNDA.n472 GNDA.n443 585
R496 GNDA.n475 GNDA.n474 585
R497 GNDA.n476 GNDA.n441 585
R498 GNDA.n1732 GNDA.n1731 585
R499 GNDA.n1732 GNDA.n322 585
R500 GNDA.n1708 GNDA.n505 585
R501 GNDA.n1709 GNDA.n503 585
R502 GNDA.n1710 GNDA.n502 585
R503 GNDA.n500 GNDA.n498 585
R504 GNDA.n1716 GNDA.n497 585
R505 GNDA.n1717 GNDA.n495 585
R506 GNDA.n1718 GNDA.n494 585
R507 GNDA.n492 GNDA.n490 585
R508 GNDA.n1723 GNDA.n489 585
R509 GNDA.n1724 GNDA.n487 585
R510 GNDA.n486 GNDA.n482 585
R511 GNDA.n1729 GNDA.n481 585
R512 GNDA.n1729 GNDA.n1728 585
R513 GNDA.n1726 GNDA.n482 585
R514 GNDA.n1725 GNDA.n1724 585
R515 GNDA.n1723 GNDA.n1722 585
R516 GNDA.n1721 GNDA.n490 585
R517 GNDA.n1719 GNDA.n1718 585
R518 GNDA.n1717 GNDA.n491 585
R519 GNDA.n1716 GNDA.n1715 585
R520 GNDA.n1713 GNDA.n498 585
R521 GNDA.n1711 GNDA.n1710 585
R522 GNDA.n1709 GNDA.n499 585
R523 GNDA.n1708 GNDA.n1707 585
R524 GNDA.n1147 GNDA.n869 585
R525 GNDA.n1150 GNDA.n1149 585
R526 GNDA.n1145 GNDA.n872 585
R527 GNDA.n1143 GNDA.n1142 585
R528 GNDA.n874 GNDA.n873 585
R529 GNDA.n1136 GNDA.n1135 585
R530 GNDA.n1133 GNDA.n876 585
R531 GNDA.n1131 GNDA.n1130 585
R532 GNDA.n878 GNDA.n877 585
R533 GNDA.n1124 GNDA.n1123 585
R534 GNDA.n1121 GNDA.n880 585
R535 GNDA.n1119 GNDA.n1118 585
R536 GNDA.n1118 GNDA.n1117 585
R537 GNDA.n880 GNDA.n879 585
R538 GNDA.n1125 GNDA.n1124 585
R539 GNDA.n1127 GNDA.n878 585
R540 GNDA.n1130 GNDA.n1129 585
R541 GNDA.n876 GNDA.n875 585
R542 GNDA.n1137 GNDA.n1136 585
R543 GNDA.n1139 GNDA.n874 585
R544 GNDA.n1142 GNDA.n1141 585
R545 GNDA.n872 GNDA.n871 585
R546 GNDA.n1151 GNDA.n1150 585
R547 GNDA.n1153 GNDA.n869 585
R548 GNDA.n1040 GNDA.n1039 585
R549 GNDA.n939 GNDA.n938 585
R550 GNDA.n1046 GNDA.n937 585
R551 GNDA.n1047 GNDA.n935 585
R552 GNDA.n1048 GNDA.n934 585
R553 GNDA.n932 GNDA.n930 585
R554 GNDA.n1054 GNDA.n929 585
R555 GNDA.n1055 GNDA.n927 585
R556 GNDA.n1056 GNDA.n926 585
R557 GNDA.n923 GNDA.n922 585
R558 GNDA.n1092 GNDA.n1091 585
R559 GNDA.n1094 GNDA.n920 585
R560 GNDA.n1088 GNDA.n920 585
R561 GNDA.n1091 GNDA.n1090 585
R562 GNDA.n1059 GNDA.n923 585
R563 GNDA.n1057 GNDA.n1056 585
R564 GNDA.n1055 GNDA.n924 585
R565 GNDA.n1054 GNDA.n1053 585
R566 GNDA.n1051 GNDA.n930 585
R567 GNDA.n1049 GNDA.n1048 585
R568 GNDA.n1047 GNDA.n931 585
R569 GNDA.n1046 GNDA.n1045 585
R570 GNDA.n1043 GNDA.n938 585
R571 GNDA.n1041 GNDA.n1040 585
R572 GNDA.n908 GNDA.n881 585
R573 GNDA.n907 GNDA.n906 585
R574 GNDA.n904 GNDA.n882 585
R575 GNDA.n902 GNDA.n901 585
R576 GNDA.n900 GNDA.n883 585
R577 GNDA.n899 GNDA.n898 585
R578 GNDA.n896 GNDA.n884 585
R579 GNDA.n894 GNDA.n893 585
R580 GNDA.n892 GNDA.n885 585
R581 GNDA.n891 GNDA.n890 585
R582 GNDA.n888 GNDA.n886 585
R583 GNDA.n797 GNDA.n796 585
R584 GNDA.n1096 GNDA.n1095 585
R585 GNDA.n1097 GNDA.n917 585
R586 GNDA.n1099 GNDA.n1098 585
R587 GNDA.n1101 GNDA.n915 585
R588 GNDA.n1103 GNDA.n1102 585
R589 GNDA.n1104 GNDA.n914 585
R590 GNDA.n1106 GNDA.n1105 585
R591 GNDA.n1108 GNDA.n912 585
R592 GNDA.n1110 GNDA.n1109 585
R593 GNDA.n1111 GNDA.n911 585
R594 GNDA.n1113 GNDA.n1112 585
R595 GNDA.n1115 GNDA.n910 585
R596 GNDA.n141 GNDA.n140 585
R597 GNDA.n1069 GNDA.n1068 585
R598 GNDA.n1071 GNDA.n1070 585
R599 GNDA.n1073 GNDA.n1065 585
R600 GNDA.n1075 GNDA.n1074 585
R601 GNDA.n1076 GNDA.n1064 585
R602 GNDA.n1078 GNDA.n1077 585
R603 GNDA.n1080 GNDA.n1062 585
R604 GNDA.n1082 GNDA.n1081 585
R605 GNDA.n1083 GNDA.n1061 585
R606 GNDA.n1085 GNDA.n1084 585
R607 GNDA.n1087 GNDA.n1060 585
R608 GNDA.n509 GNDA.n508 585
R609 GNDA.n1704 GNDA.n509 585
R610 GNDA.n1376 GNDA.n1375 585
R611 GNDA.n1373 GNDA.n580 585
R612 GNDA.n1264 GNDA.n1263 585
R613 GNDA.n1368 GNDA.n1367 585
R614 GNDA.n1366 GNDA.n1365 585
R615 GNDA.n1292 GNDA.n1268 585
R616 GNDA.n1294 GNDA.n1293 585
R617 GNDA.n1299 GNDA.n1298 585
R618 GNDA.n1297 GNDA.n1290 585
R619 GNDA.n1305 GNDA.n1304 585
R620 GNDA.n1307 GNDA.n1306 585
R621 GNDA.n1288 GNDA.n1287 585
R622 GNDA.n511 GNDA.n510 585
R623 GNDA.n1704 GNDA.n510 585
R624 GNDA.n1705 GNDA.n508 585
R625 GNDA.n1705 GNDA.n1704 585
R626 GNDA.n1534 GNDA.n507 585
R627 GNDA.n1535 GNDA.n1468 585
R628 GNDA.n1545 GNDA.n1544 585
R629 GNDA.n1547 GNDA.n1466 585
R630 GNDA.n1550 GNDA.n1549 585
R631 GNDA.n1551 GNDA.n1462 585
R632 GNDA.n1560 GNDA.n1559 585
R633 GNDA.n1562 GNDA.n1461 585
R634 GNDA.n1565 GNDA.n1564 585
R635 GNDA.n1457 GNDA.n1456 585
R636 GNDA.n1572 GNDA.n1571 585
R637 GNDA.n1575 GNDA.n1574 585
R638 GNDA.n1703 GNDA.n511 585
R639 GNDA.n1704 GNDA.n1703 585
R640 GNDA.n1577 GNDA.n512 585
R641 GNDA.n1578 GNDA.n1392 585
R642 GNDA.n1588 GNDA.n1587 585
R643 GNDA.n1590 GNDA.n1390 585
R644 GNDA.n1593 GNDA.n1592 585
R645 GNDA.n1594 GNDA.n1386 585
R646 GNDA.n1603 GNDA.n1602 585
R647 GNDA.n1605 GNDA.n1385 585
R648 GNDA.n1608 GNDA.n1607 585
R649 GNDA.n1609 GNDA.n1379 585
R650 GNDA.n1618 GNDA.n1617 585
R651 GNDA.n1620 GNDA.n574 585
R652 GNDA.n1959 GNDA.n128 585
R653 GNDA.n1958 GNDA.n132 585
R654 GNDA.n1958 GNDA.n1957 585
R655 GNDA.n1952 GNDA.n131 585
R656 GNDA.n1956 GNDA.n131 585
R657 GNDA.n1954 GNDA.n1953 585
R658 GNDA.n1955 GNDA.n1954 585
R659 GNDA.n1951 GNDA.n134 585
R660 GNDA.n134 GNDA.n133 585
R661 GNDA.n1950 GNDA.n1949 585
R662 GNDA.n1949 GNDA.n80 585
R663 GNDA.n1948 GNDA.n135 585
R664 GNDA.n1948 GNDA.n79 585
R665 GNDA.n1947 GNDA.n137 585
R666 GNDA.n1947 GNDA.n1946 585
R667 GNDA.n1941 GNDA.n136 585
R668 GNDA.n1945 GNDA.n136 585
R669 GNDA.n1943 GNDA.n1942 585
R670 GNDA.n1944 GNDA.n1943 585
R671 GNDA.n1940 GNDA.n139 585
R672 GNDA.n139 GNDA.n138 585
R673 GNDA.n1939 GNDA.n1938 585
R674 GNDA.n1938 GNDA.n1937 585
R675 GNDA.n1962 GNDA.n1961 585
R676 GNDA.n573 GNDA.n572 585
R677 GNDA.n1625 GNDA.n1624 585
R678 GNDA.n1626 GNDA.n1625 585
R679 GNDA.n570 GNDA.n569 585
R680 GNDA.n1627 GNDA.n570 585
R681 GNDA.n1630 GNDA.n1629 585
R682 GNDA.n1629 GNDA.n1628 585
R683 GNDA.n1631 GNDA.n568 585
R684 GNDA.n571 GNDA.n568 585
R685 GNDA.n1633 GNDA.n1632 585
R686 GNDA.n1633 GNDA.n152 585
R687 GNDA.n1634 GNDA.n567 585
R688 GNDA.n1634 GNDA.n153 585
R689 GNDA.n1637 GNDA.n1636 585
R690 GNDA.n1636 GNDA.n1635 585
R691 GNDA.n1638 GNDA.n565 585
R692 GNDA.n565 GNDA.n564 585
R693 GNDA.n1640 GNDA.n1639 585
R694 GNDA.n1641 GNDA.n1640 585
R695 GNDA.n566 GNDA.n563 585
R696 GNDA.n1642 GNDA.n563 585
R697 GNDA.n1644 GNDA.n561 585
R698 GNDA.n1644 GNDA.n1643 585
R699 GNDA.n1621 GNDA.n178 585
R700 GNDA.n1833 GNDA.n1832 585
R701 GNDA.n1836 GNDA.n242 585
R702 GNDA.n242 GNDA.n241 585
R703 GNDA.n1838 GNDA.n1837 585
R704 GNDA.n1839 GNDA.n1838 585
R705 GNDA.n243 GNDA.n240 585
R706 GNDA.n1840 GNDA.n240 585
R707 GNDA.n1842 GNDA.n239 585
R708 GNDA.n1842 GNDA.n1841 585
R709 GNDA.n1844 GNDA.n1843 585
R710 GNDA.n1843 GNDA.n146 585
R711 GNDA.n1845 GNDA.n238 585
R712 GNDA.n238 GNDA.n147 585
R713 GNDA.n1847 GNDA.n1846 585
R714 GNDA.n1848 GNDA.n1847 585
R715 GNDA.n237 GNDA.n236 585
R716 GNDA.n1849 GNDA.n237 585
R717 GNDA.n1852 GNDA.n1851 585
R718 GNDA.n1851 GNDA.n1850 585
R719 GNDA.n1853 GNDA.n235 585
R720 GNDA.n235 GNDA.n234 585
R721 GNDA.n1855 GNDA.n1854 585
R722 GNDA.n1856 GNDA.n1855 585
R723 GNDA.n1831 GNDA.n1830 585
R724 GNDA.n2154 GNDA.n2153 585
R725 GNDA.n2151 GNDA.n2150 585
R726 GNDA.n2150 GNDA.n2114 585
R727 GNDA.n2159 GNDA.n2158 585
R728 GNDA.n2161 GNDA.n2149 585
R729 GNDA.n2164 GNDA.n2163 585
R730 GNDA.n2147 GNDA.n2146 585
R731 GNDA.n2169 GNDA.n2168 585
R732 GNDA.n2171 GNDA.n2145 585
R733 GNDA.n2174 GNDA.n2173 585
R734 GNDA.n2143 GNDA.n2142 585
R735 GNDA.n2179 GNDA.n2178 585
R736 GNDA.n2181 GNDA.n2141 585
R737 GNDA.n2183 GNDA.n2182 585
R738 GNDA.n2182 GNDA.n2114 585
R739 GNDA.n2316 GNDA.n2311 585
R740 GNDA.n2314 GNDA.n2310 585
R741 GNDA.n2319 GNDA.n2310 585
R742 GNDA.n2313 GNDA.n2309 585
R743 GNDA.n2279 GNDA.n2274 585
R744 GNDA.n2277 GNDA.n2273 585
R745 GNDA.n2282 GNDA.n2273 585
R746 GNDA.n2276 GNDA.n2259 585
R747 GNDA.n2130 GNDA.n2129 585
R748 GNDA.n2213 GNDA.n2128 585
R749 GNDA.n2217 GNDA.n2128 585
R750 GNDA.n2212 GNDA.n2211 585
R751 GNDA.n2210 GNDA.n2209 585
R752 GNDA.n2208 GNDA.n2207 585
R753 GNDA.n2206 GNDA.n2205 585
R754 GNDA.n2204 GNDA.n2203 585
R755 GNDA.n2202 GNDA.n2201 585
R756 GNDA.n2200 GNDA.n2199 585
R757 GNDA.n2198 GNDA.n2197 585
R758 GNDA.n2196 GNDA.n2195 585
R759 GNDA.n2194 GNDA.n2193 585
R760 GNDA.n2191 GNDA.n2127 585
R761 GNDA.n2217 GNDA.n2127 585
R762 GNDA.n2499 GNDA.n2498 585
R763 GNDA.n2532 GNDA.n2497 585
R764 GNDA.n2536 GNDA.n2497 585
R765 GNDA.n2531 GNDA.n2530 585
R766 GNDA.n2529 GNDA.n2528 585
R767 GNDA.n2527 GNDA.n2526 585
R768 GNDA.n2525 GNDA.n2524 585
R769 GNDA.n2523 GNDA.n2522 585
R770 GNDA.n2521 GNDA.n2520 585
R771 GNDA.n2519 GNDA.n2518 585
R772 GNDA.n2517 GNDA.n2516 585
R773 GNDA.n2515 GNDA.n2514 585
R774 GNDA.n2513 GNDA.n2512 585
R775 GNDA.n2510 GNDA.n25 585
R776 GNDA.n2536 GNDA.n25 585
R777 GNDA.n2455 GNDA.n2454 585
R778 GNDA.n2492 GNDA.n2453 585
R779 GNDA.n2496 GNDA.n2453 585
R780 GNDA.n2491 GNDA.n2490 585
R781 GNDA.n2489 GNDA.n2488 585
R782 GNDA.n2487 GNDA.n2486 585
R783 GNDA.n2485 GNDA.n2484 585
R784 GNDA.n2483 GNDA.n2482 585
R785 GNDA.n2481 GNDA.n2480 585
R786 GNDA.n2479 GNDA.n2478 585
R787 GNDA.n2477 GNDA.n2476 585
R788 GNDA.n2475 GNDA.n2474 585
R789 GNDA.n2473 GNDA.n2472 585
R790 GNDA.n2470 GNDA.n31 585
R791 GNDA.n2496 GNDA.n31 585
R792 GNDA.n2117 GNDA.n2116 585
R793 GNDA.n2421 GNDA.n2115 585
R794 GNDA.n2425 GNDA.n2115 585
R795 GNDA.n2420 GNDA.n2419 585
R796 GNDA.n2418 GNDA.n2417 585
R797 GNDA.n2415 GNDA.n2113 585
R798 GNDA.n2425 GNDA.n2113 585
R799 GNDA.n2394 GNDA.n2220 585
R800 GNDA.n2392 GNDA.n2219 585
R801 GNDA.n2397 GNDA.n2219 585
R802 GNDA.n2379 GNDA.n2234 585
R803 GNDA.n2386 GNDA.n2385 585
R804 GNDA.n2385 GNDA.n2384 585
R805 GNDA.n2263 GNDA.n2261 585
R806 GNDA.n2267 GNDA.n2260 585
R807 GNDA.n2272 GNDA.n2260 585
R808 GNDA.n2227 GNDA.n2223 585
R809 GNDA.n2229 GNDA.n2228 585
R810 GNDA.n2228 GNDA.n18 585
R811 GNDA.n2400 GNDA.n2399 585
R812 GNDA.n2405 GNDA.n2398 585
R813 GNDA.n2409 GNDA.n2398 585
R814 GNDA.n2404 GNDA.n2403 585
R815 GNDA.n2402 GNDA.n2121 585
R816 GNDA.n2411 GNDA.n2410 585
R817 GNDA.n2410 GNDA.n2409 585
R818 GNDA.n2539 GNDA.n2538 585
R819 GNDA.n2544 GNDA.n2537 585
R820 GNDA.n2548 GNDA.n2537 585
R821 GNDA.n2543 GNDA.n2542 585
R822 GNDA.n2541 GNDA.n17 585
R823 GNDA.n2550 GNDA.n2549 585
R824 GNDA.n2549 GNDA.n2548 585
R825 GNDA.n2440 GNDA.n2439 585
R826 GNDA.n2448 GNDA.n2438 585
R827 GNDA.n2452 GNDA.n2438 585
R828 GNDA.n2447 GNDA.n2446 585
R829 GNDA.n2445 GNDA.n2444 585
R830 GNDA.n2442 GNDA.n33 585
R831 GNDA.n2452 GNDA.n33 585
R832 GNDA.n2331 GNDA.n2245 585
R833 GNDA.n2329 GNDA.n2244 585
R834 GNDA.n2334 GNDA.n2244 585
R835 GNDA.n2341 GNDA.n2336 585
R836 GNDA.n2339 GNDA.n2335 585
R837 GNDA.n2344 GNDA.n2335 585
R838 GNDA.n2374 GNDA.n2239 585
R839 GNDA.n2372 GNDA.n2238 585
R840 GNDA.n2377 GNDA.n2238 585
R841 GNDA.n2363 GNDA.n2243 585
R842 GNDA.n2368 GNDA.n2367 585
R843 GNDA.n2367 GNDA.n2366 585
R844 GNDA.n2066 GNDA.n76 585
R845 GNDA.n2069 GNDA.n2068 585
R846 GNDA.n2070 GNDA.n2069 585
R847 GNDA.n2061 GNDA.n2060 585
R848 GNDA.n1146 GNDA.n867 585
R849 GNDA.n1146 GNDA.n855 585
R850 GNDA.n1234 GNDA.n799 585
R851 GNDA.n1234 GNDA.n1233 585
R852 GNDA.n1221 GNDA.n800 585
R853 GNDA.n1232 GNDA.n800 585
R854 GNDA.n1230 GNDA.n1229 585
R855 GNDA.n1231 GNDA.n1230 585
R856 GNDA.n803 GNDA.n801 585
R857 GNDA.n833 GNDA.n801 585
R858 GNDA.n832 GNDA.n831 585
R859 GNDA.n834 GNDA.n832 585
R860 GNDA.n837 GNDA.n836 585
R861 GNDA.n836 GNDA.n835 585
R862 GNDA.n838 GNDA.n827 585
R863 GNDA.n827 GNDA.n826 585
R864 GNDA.n849 GNDA.n848 585
R865 GNDA.n850 GNDA.n849 585
R866 GNDA.n843 GNDA.n825 585
R867 GNDA.n851 GNDA.n825 585
R868 GNDA.n853 GNDA.n824 585
R869 GNDA.n853 GNDA.n852 585
R870 GNDA.n1167 GNDA.n1166 585
R871 GNDA.n1166 GNDA.n1165 585
R872 GNDA.n942 GNDA.n854 585
R873 GNDA.n1164 GNDA.n854 585
R874 GNDA.n1038 GNDA.n1016 585
R875 GNDA.n1038 GNDA.n1037 585
R876 GNDA.n1154 GNDA.n867 585
R877 GNDA.n1155 GNDA.n1154 585
R878 GNDA.n944 GNDA.n868 585
R879 GNDA.n868 GNDA.n866 585
R880 GNDA.n67 GNDA.n65 585
R881 GNDA.n2077 GNDA.n67 585
R882 GNDA.n2092 GNDA.n2091 585
R883 GNDA.n2091 GNDA.n2090 585
R884 GNDA.n2079 GNDA.n68 585
R885 GNDA.n2089 GNDA.n68 585
R886 GNDA.n2087 GNDA.n2086 585
R887 GNDA.n2088 GNDA.n2087 585
R888 GNDA.n2082 GNDA.n42 585
R889 GNDA.n2078 GNDA.n42 585
R890 GNDA.n2100 GNDA.n2099 585
R891 GNDA.n2101 GNDA.n2100 585
R892 GNDA.n44 GNDA.n43 585
R893 GNDA.n1003 GNDA.n43 585
R894 GNDA.n1002 GNDA.n1001 585
R895 GNDA.n1004 GNDA.n1002 585
R896 GNDA.n1008 GNDA.n1007 585
R897 GNDA.n1007 GNDA.n1006 585
R898 GNDA.n1012 GNDA.n941 585
R899 GNDA.n1005 GNDA.n941 585
R900 GNDA.n1015 GNDA.n1014 585
R901 GNDA.n1017 GNDA.n1015 585
R902 GNDA.n1016 GNDA.n111 585
R903 GNDA.n1028 GNDA.n111 585
R904 GNDA.n2033 GNDA.n2032 585
R905 GNDA.n2034 GNDA.n2033 585
R906 GNDA.n106 GNDA.n104 585
R907 GNDA.n2035 GNDA.n106 585
R908 GNDA.n2050 GNDA.n2049 585
R909 GNDA.n2049 GNDA.n2048 585
R910 GNDA.n2037 GNDA.n107 585
R911 GNDA.n2047 GNDA.n107 585
R912 GNDA.n2045 GNDA.n2044 585
R913 GNDA.n2046 GNDA.n2045 585
R914 GNDA.n2040 GNDA.n81 585
R915 GNDA.n2036 GNDA.n81 585
R916 GNDA.n2058 GNDA.n2057 585
R917 GNDA.n2059 GNDA.n2058 585
R918 GNDA.n83 GNDA.n82 585
R919 GNDA.n117 GNDA.n82 585
R920 GNDA.n122 GNDA.n121 585
R921 GNDA.n123 GNDA.n122 585
R922 GNDA.n115 GNDA.n114 585
R923 GNDA.n124 GNDA.n115 585
R924 GNDA.n1975 GNDA.n1974 585
R925 GNDA.n1974 GNDA.n1973 585
R926 GNDA.n129 GNDA.n116 585
R927 GNDA.n1972 GNDA.n116 585
R928 GNDA.n173 GNDA.n70 585
R929 GNDA.n174 GNDA.n173 585
R930 GNDA.n172 GNDA.n171 585
R931 GNDA.n170 GNDA.n163 585
R932 GNDA.n165 GNDA.n164 585
R933 GNDA.t221 GNDA.n149 512.884
R934 GNDA.n2184 GNDA.t294 505.467
R935 GNDA.n2190 GNDA.t271 505.467
R936 GNDA.n2509 GNDA.t260 505.467
R937 GNDA.n2469 GNDA.t250 505.467
R938 GNDA.n2391 GNDA.t291 499.442
R939 GNDA.n2230 GNDA.t297 499.442
R940 GNDA.n2328 GNDA.t229 489.401
R941 GNDA.n2338 GNDA.t244 489.401
R942 GNDA.n2371 GNDA.t223 489.401
R943 GNDA.n2369 GNDA.t241 489.401
R944 GNDA.n2387 GNDA.t303 475.976
R945 GNDA.n2387 GNDA.t300 475.976
R946 GNDA.n2265 GNDA.t288 475.976
R947 GNDA.n2265 GNDA.t265 475.976
R948 GNDA.n2434 GNDA.n34 459.341
R949 GNDA.n2110 GNDA.n2109 459.341
R950 GNDA.n2409 GNDA.n2397 445.375
R951 GNDA.n2548 GNDA.n18 445.375
R952 GNDA.n110 GNDA.t315 433.382
R953 GNDA.n857 GNDA.t274 409.067
R954 GNDA.n1161 GNDA.t281 409.067
R955 GNDA.n1158 GNDA.t306 409.067
R956 GNDA.n1034 GNDA.t254 409.067
R957 GNDA.n1031 GNDA.t277 409.067
R958 GNDA.n1969 GNDA.t268 409.067
R959 GNDA.t230 GNDA.n2334 404.082
R960 GNDA.n2366 GNDA.t242 404.082
R961 GNDA.t221 GNDA.n150 391.411
R962 GNDA.t125 GNDA.t230 329.252
R963 GNDA.t10 GNDA.t125 329.252
R964 GNDA.t74 GNDA.t10 329.252
R965 GNDA.t77 GNDA.t74 329.252
R966 GNDA.t19 GNDA.t77 329.252
R967 GNDA.t78 GNDA.t19 329.252
R968 GNDA.t130 GNDA.t78 329.252
R969 GNDA.t157 GNDA.t130 329.252
R970 GNDA.t17 GNDA.t150 329.252
R971 GNDA.t150 GNDA.t98 329.252
R972 GNDA.t96 GNDA.t69 329.252
R973 GNDA.t69 GNDA.t127 329.252
R974 GNDA.t345 GNDA.t129 329.252
R975 GNDA.t20 GNDA.t345 329.252
R976 GNDA.t344 GNDA.t20 329.252
R977 GNDA.t75 GNDA.t344 329.252
R978 GNDA.t158 GNDA.t75 329.252
R979 GNDA.t73 GNDA.t158 329.252
R980 GNDA.t160 GNDA.t73 329.252
R981 GNDA.t242 GNDA.t160 329.252
R982 GNDA.n2359 GNDA.t232 328.733
R983 GNDA.n2347 GNDA.t238 328.733
R984 GNDA.t221 GNDA.n158 172.876
R985 GNDA.t221 GNDA.n156 172.876
R986 GNDA.t221 GNDA.n175 172.876
R987 GNDA.n921 GNDA.t221 172.876
R988 GNDA.t221 GNDA.n157 172.615
R989 GNDA.t221 GNDA.n155 172.615
R990 GNDA.n870 GNDA.t221 172.615
R991 GNDA.t221 GNDA.n78 172.615
R992 GNDA.t221 GNDA.t154 294.625
R993 GNDA.n2156 GNDA.n2155 267.125
R994 GNDA.n2177 GNDA.n2140 267.125
R995 GNDA.n2215 GNDA.n2214 267.125
R996 GNDA.n2192 GNDA.n2139 267.125
R997 GNDA.n2407 GNDA.n2406 267.125
R998 GNDA.n2401 GNDA.n2120 267.125
R999 GNDA.n2423 GNDA.n2422 267.125
R1000 GNDA.n2416 GNDA.n2118 267.125
R1001 GNDA.n2546 GNDA.n2545 267.125
R1002 GNDA.n2540 GNDA.n16 267.125
R1003 GNDA.n2450 GNDA.n2449 267.125
R1004 GNDA.n2443 GNDA.n2441 267.125
R1005 GNDA.n2534 GNDA.n2533 267.125
R1006 GNDA.n2511 GNDA.n2508 267.125
R1007 GNDA.n2494 GNDA.n2493 267.125
R1008 GNDA.n2471 GNDA.n2464 267.125
R1009 GNDA.n1258 GNDA.n789 264.301
R1010 GNDA.n1258 GNDA.n734 264.301
R1011 GNDA.n1261 GNDA.n1260 264.301
R1012 GNDA.n1960 GNDA.n130 264.301
R1013 GNDA.n1623 GNDA.n1622 264.301
R1014 GNDA.n1835 GNDA.n1834 264.301
R1015 GNDA.n1938 GNDA.n141 259.416
R1016 GNDA.n1095 GNDA.n1094 259.416
R1017 GNDA.n1913 GNDA.n1912 259.416
R1018 GNDA.n1119 GNDA.n881 259.416
R1019 GNDA.n747 GNDA.n481 259.416
R1020 GNDA.n1645 GNDA.n1644 259.416
R1021 GNDA.n1669 GNDA.n524 259.416
R1022 GNDA.n1855 GNDA.n233 259.416
R1023 GNDA.n338 GNDA.n218 259.416
R1024 GNDA.n705 GNDA.n704 258.334
R1025 GNDA.n1206 GNDA.n1205 258.334
R1026 GNDA.n1344 GNDA.n1285 258.334
R1027 GNDA.n1519 GNDA.n1474 258.334
R1028 GNDA.n1440 GNDA.n1398 258.334
R1029 GNDA.n425 GNDA.n383 258.334
R1030 GNDA.n306 GNDA.n264 258.334
R1031 GNDA.n963 GNDA.n962 258.334
R1032 GNDA.n2014 GNDA.n2013 258.334
R1033 GNDA.n2345 GNDA.t76 254.423
R1034 GNDA.t71 GNDA.n2344 254.423
R1035 GNDA.n2377 GNDA.t30 254.423
R1036 GNDA.n2361 GNDA.t11 254.423
R1037 GNDA.n1258 GNDA.n1257 254.34
R1038 GNDA.n1258 GNDA.n794 254.34
R1039 GNDA.n1258 GNDA.n793 254.34
R1040 GNDA.n1258 GNDA.n792 254.34
R1041 GNDA.n1258 GNDA.n791 254.34
R1042 GNDA.n1258 GNDA.n584 254.34
R1043 GNDA.n1258 GNDA.n585 254.34
R1044 GNDA.n1258 GNDA.n586 254.34
R1045 GNDA.n1258 GNDA.n587 254.34
R1046 GNDA.n1258 GNDA.n588 254.34
R1047 GNDA.n1258 GNDA.n735 254.34
R1048 GNDA.n1258 GNDA.n736 254.34
R1049 GNDA.n1258 GNDA.n737 254.34
R1050 GNDA.n1258 GNDA.n738 254.34
R1051 GNDA.n1258 GNDA.n788 254.34
R1052 GNDA.n1259 GNDA.n1258 254.34
R1053 GNDA.n1697 GNDA.n156 254.34
R1054 GNDA.n1694 GNDA.n156 254.34
R1055 GNDA.n1684 GNDA.n156 254.34
R1056 GNDA.n1682 GNDA.n156 254.34
R1057 GNDA.n1672 GNDA.n156 254.34
R1058 GNDA.n1670 GNDA.n156 254.34
R1059 GNDA.n1666 GNDA.n155 254.34
R1060 GNDA.n1676 GNDA.n155 254.34
R1061 GNDA.n1678 GNDA.n155 254.34
R1062 GNDA.n1688 GNDA.n155 254.34
R1063 GNDA.n1690 GNDA.n155 254.34
R1064 GNDA.n1701 GNDA.n155 254.34
R1065 GNDA.n748 GNDA.n180 254.34
R1066 GNDA.n753 GNDA.n180 254.34
R1067 GNDA.n746 GNDA.n180 254.34
R1068 GNDA.n760 GNDA.n180 254.34
R1069 GNDA.n743 GNDA.n180 254.34
R1070 GNDA.n767 GNDA.n180 254.34
R1071 GNDA.n548 GNDA.n180 254.34
R1072 GNDA.n546 GNDA.n180 254.34
R1073 GNDA.n540 GNDA.n180 254.34
R1074 GNDA.n538 GNDA.n180 254.34
R1075 GNDA.n532 GNDA.n180 254.34
R1076 GNDA.n530 GNDA.n180 254.34
R1077 GNDA.n562 GNDA.n180 254.34
R1078 GNDA.n1650 GNDA.n180 254.34
R1079 GNDA.n559 GNDA.n180 254.34
R1080 GNDA.n1657 GNDA.n180 254.34
R1081 GNDA.n556 GNDA.n180 254.34
R1082 GNDA.n1664 GNDA.n180 254.34
R1083 GNDA.n611 GNDA.n245 254.34
R1084 GNDA.n614 GNDA.n245 254.34
R1085 GNDA.n644 GNDA.n245 254.34
R1086 GNDA.n646 GNDA.n245 254.34
R1087 GNDA.n660 GNDA.n245 254.34
R1088 GNDA.n664 GNDA.n245 254.34
R1089 GNDA.n1733 GNDA.n245 254.34
R1090 GNDA.n1747 GNDA.n245 254.34
R1091 GNDA.n1749 GNDA.n245 254.34
R1092 GNDA.n1762 GNDA.n245 254.34
R1093 GNDA.n1764 GNDA.n245 254.34
R1094 GNDA.n1777 GNDA.n245 254.34
R1095 GNDA.n1784 GNDA.n245 254.34
R1096 GNDA.n1798 GNDA.n245 254.34
R1097 GNDA.n1800 GNDA.n245 254.34
R1098 GNDA.n1813 GNDA.n245 254.34
R1099 GNDA.n1815 GNDA.n245 254.34
R1100 GNDA.n1828 GNDA.n245 254.34
R1101 GNDA.n442 GNDA.n148 254.34
R1102 GNDA.n467 GNDA.n148 254.34
R1103 GNDA.n464 GNDA.n148 254.34
R1104 GNDA.n454 GNDA.n148 254.34
R1105 GNDA.n452 GNDA.n148 254.34
R1106 GNDA.n1911 GNDA.n148 254.34
R1107 GNDA.n1907 GNDA.n145 254.34
R1108 GNDA.n449 GNDA.n145 254.34
R1109 GNDA.n458 GNDA.n145 254.34
R1110 GNDA.n460 GNDA.n145 254.34
R1111 GNDA.n471 GNDA.n145 254.34
R1112 GNDA.n473 GNDA.n145 254.34
R1113 GNDA.n504 GNDA.n158 254.34
R1114 GNDA.n501 GNDA.n158 254.34
R1115 GNDA.n496 GNDA.n158 254.34
R1116 GNDA.n493 GNDA.n158 254.34
R1117 GNDA.n488 GNDA.n158 254.34
R1118 GNDA.n485 GNDA.n158 254.34
R1119 GNDA.n1727 GNDA.n157 254.34
R1120 GNDA.n484 GNDA.n157 254.34
R1121 GNDA.n1720 GNDA.n157 254.34
R1122 GNDA.n1714 GNDA.n157 254.34
R1123 GNDA.n1712 GNDA.n157 254.34
R1124 GNDA.n1706 GNDA.n157 254.34
R1125 GNDA.n1148 GNDA.n175 254.34
R1126 GNDA.n1144 GNDA.n175 254.34
R1127 GNDA.n1134 GNDA.n175 254.34
R1128 GNDA.n1132 GNDA.n175 254.34
R1129 GNDA.n1122 GNDA.n175 254.34
R1130 GNDA.n1120 GNDA.n175 254.34
R1131 GNDA.n1116 GNDA.n870 254.34
R1132 GNDA.n1126 GNDA.n870 254.34
R1133 GNDA.n1128 GNDA.n870 254.34
R1134 GNDA.n1138 GNDA.n870 254.34
R1135 GNDA.n1140 GNDA.n870 254.34
R1136 GNDA.n1152 GNDA.n870 254.34
R1137 GNDA.n940 GNDA.n921 254.34
R1138 GNDA.n936 GNDA.n921 254.34
R1139 GNDA.n933 GNDA.n921 254.34
R1140 GNDA.n928 GNDA.n921 254.34
R1141 GNDA.n925 GNDA.n921 254.34
R1142 GNDA.n1093 GNDA.n921 254.34
R1143 GNDA.n1089 GNDA.n78 254.34
R1144 GNDA.n1058 GNDA.n78 254.34
R1145 GNDA.n1052 GNDA.n78 254.34
R1146 GNDA.n1050 GNDA.n78 254.34
R1147 GNDA.n1044 GNDA.n78 254.34
R1148 GNDA.n1042 GNDA.n78 254.34
R1149 GNDA.n905 GNDA.n177 254.34
R1150 GNDA.n903 GNDA.n177 254.34
R1151 GNDA.n897 GNDA.n177 254.34
R1152 GNDA.n895 GNDA.n177 254.34
R1153 GNDA.n889 GNDA.n177 254.34
R1154 GNDA.n887 GNDA.n177 254.34
R1155 GNDA.n919 GNDA.n177 254.34
R1156 GNDA.n1100 GNDA.n177 254.34
R1157 GNDA.n916 GNDA.n177 254.34
R1158 GNDA.n1107 GNDA.n177 254.34
R1159 GNDA.n913 GNDA.n177 254.34
R1160 GNDA.n1114 GNDA.n177 254.34
R1161 GNDA.n1067 GNDA.n177 254.34
R1162 GNDA.n1072 GNDA.n177 254.34
R1163 GNDA.n1066 GNDA.n177 254.34
R1164 GNDA.n1079 GNDA.n177 254.34
R1165 GNDA.n1063 GNDA.n177 254.34
R1166 GNDA.n1086 GNDA.n177 254.34
R1167 GNDA.n1378 GNDA.n1377 254.34
R1168 GNDA.n1378 GNDA.n579 254.34
R1169 GNDA.n1378 GNDA.n578 254.34
R1170 GNDA.n1378 GNDA.n577 254.34
R1171 GNDA.n1378 GNDA.n576 254.34
R1172 GNDA.n1378 GNDA.n575 254.34
R1173 GNDA.n1467 GNDA.n1378 254.34
R1174 GNDA.n1546 GNDA.n1378 254.34
R1175 GNDA.n1548 GNDA.n1378 254.34
R1176 GNDA.n1561 GNDA.n1378 254.34
R1177 GNDA.n1563 GNDA.n1378 254.34
R1178 GNDA.n1573 GNDA.n1378 254.34
R1179 GNDA.n1391 GNDA.n1378 254.34
R1180 GNDA.n1589 GNDA.n1378 254.34
R1181 GNDA.n1591 GNDA.n1378 254.34
R1182 GNDA.n1604 GNDA.n1378 254.34
R1183 GNDA.n1606 GNDA.n1378 254.34
R1184 GNDA.n1619 GNDA.n1378 254.34
R1185 GNDA.t221 GNDA.n208 250.349
R1186 GNDA.n1088 GNDA.n1087 249.663
R1187 GNDA.n1117 GNDA.n1115 249.663
R1188 GNDA.n1935 GNDA.n182 249.663
R1189 GNDA.n1256 GNDA.n796 249.663
R1190 GNDA.n769 GNDA.n768 249.663
R1191 GNDA.n1667 GNDA.n1665 249.663
R1192 GNDA.n1728 GNDA.n483 249.663
R1193 GNDA.n1879 GNDA.n221 249.663
R1194 GNDA.n1906 GNDA.n1905 249.663
R1195 GNDA.n2069 GNDA.n76 246.25
R1196 GNDA.n2069 GNDA.n2060 246.25
R1197 GNDA.n2367 GNDA.n2243 246.25
R1198 GNDA.n2239 GNDA.n2238 246.25
R1199 GNDA.n2336 GNDA.n2335 246.25
R1200 GNDA.n2245 GNDA.n2244 246.25
R1201 GNDA.n2439 GNDA.n2438 246.25
R1202 GNDA.n2446 GNDA.n2438 246.25
R1203 GNDA.n2444 GNDA.n33 246.25
R1204 GNDA.n2538 GNDA.n2537 246.25
R1205 GNDA.n2542 GNDA.n2537 246.25
R1206 GNDA.n2549 GNDA.n17 246.25
R1207 GNDA.n2399 GNDA.n2398 246.25
R1208 GNDA.n2403 GNDA.n2398 246.25
R1209 GNDA.n2410 GNDA.n2121 246.25
R1210 GNDA.n2228 GNDA.n2227 246.25
R1211 GNDA.n2261 GNDA.n2260 246.25
R1212 GNDA.n2385 GNDA.n2234 246.25
R1213 GNDA.n2220 GNDA.n2219 246.25
R1214 GNDA.n2116 GNDA.n2115 246.25
R1215 GNDA.n2419 GNDA.n2115 246.25
R1216 GNDA.n2417 GNDA.n2113 246.25
R1217 GNDA.n2454 GNDA.n2453 246.25
R1218 GNDA.n2490 GNDA.n2453 246.25
R1219 GNDA.n2488 GNDA.n2487 246.25
R1220 GNDA.n2484 GNDA.n2483 246.25
R1221 GNDA.n2480 GNDA.n2479 246.25
R1222 GNDA.n2476 GNDA.n2475 246.25
R1223 GNDA.n2472 GNDA.n31 246.25
R1224 GNDA.n2498 GNDA.n2497 246.25
R1225 GNDA.n2530 GNDA.n2497 246.25
R1226 GNDA.n2528 GNDA.n2527 246.25
R1227 GNDA.n2524 GNDA.n2523 246.25
R1228 GNDA.n2520 GNDA.n2519 246.25
R1229 GNDA.n2516 GNDA.n2515 246.25
R1230 GNDA.n2512 GNDA.n25 246.25
R1231 GNDA.n2129 GNDA.n2128 246.25
R1232 GNDA.n2211 GNDA.n2128 246.25
R1233 GNDA.n2209 GNDA.n2208 246.25
R1234 GNDA.n2205 GNDA.n2204 246.25
R1235 GNDA.n2201 GNDA.n2200 246.25
R1236 GNDA.n2197 GNDA.n2196 246.25
R1237 GNDA.n2193 GNDA.n2127 246.25
R1238 GNDA.n2274 GNDA.n2273 246.25
R1239 GNDA.n2273 GNDA.n2259 246.25
R1240 GNDA.n2311 GNDA.n2310 246.25
R1241 GNDA.n2310 GNDA.n2309 246.25
R1242 GNDA.n2153 GNDA.n2150 246.25
R1243 GNDA.n2159 GNDA.n2150 246.25
R1244 GNDA.n2163 GNDA.n2161 246.25
R1245 GNDA.n2169 GNDA.n2146 246.25
R1246 GNDA.n2173 GNDA.n2171 246.25
R1247 GNDA.n2179 GNDA.n2142 246.25
R1248 GNDA.n2182 GNDA.n2181 246.25
R1249 GNDA.n173 GNDA.n172 246.25
R1250 GNDA.n164 GNDA.n163 246.25
R1251 GNDA.n1965 GNDA.n1964 241.643
R1252 GNDA.n2152 GNDA.n2114 241.643
R1253 GNDA.n2160 GNDA.n2114 241.643
R1254 GNDA.n2162 GNDA.n2114 241.643
R1255 GNDA.n2170 GNDA.n2114 241.643
R1256 GNDA.n2172 GNDA.n2114 241.643
R1257 GNDA.n2180 GNDA.n2114 241.643
R1258 GNDA.n2319 GNDA.n2318 241.643
R1259 GNDA.n2320 GNDA.n2319 241.643
R1260 GNDA.n2282 GNDA.n2281 241.643
R1261 GNDA.n2283 GNDA.n2282 241.643
R1262 GNDA.n2217 GNDA.n2216 241.643
R1263 GNDA.n2217 GNDA.n2122 241.643
R1264 GNDA.n2217 GNDA.n2123 241.643
R1265 GNDA.n2217 GNDA.n2124 241.643
R1266 GNDA.n2217 GNDA.n2125 241.643
R1267 GNDA.n2217 GNDA.n2126 241.643
R1268 GNDA.n2536 GNDA.n2535 241.643
R1269 GNDA.n2536 GNDA.n20 241.643
R1270 GNDA.n2536 GNDA.n21 241.643
R1271 GNDA.n2536 GNDA.n22 241.643
R1272 GNDA.n2536 GNDA.n23 241.643
R1273 GNDA.n2536 GNDA.n24 241.643
R1274 GNDA.n2496 GNDA.n2495 241.643
R1275 GNDA.n2496 GNDA.n26 241.643
R1276 GNDA.n2496 GNDA.n27 241.643
R1277 GNDA.n2496 GNDA.n28 241.643
R1278 GNDA.n2496 GNDA.n29 241.643
R1279 GNDA.n2496 GNDA.n30 241.643
R1280 GNDA.n2425 GNDA.n2424 241.643
R1281 GNDA.n2425 GNDA.n2112 241.643
R1282 GNDA.n2397 GNDA.n2396 241.643
R1283 GNDA.n2384 GNDA.n2383 241.643
R1284 GNDA.n2272 GNDA.n2271 241.643
R1285 GNDA.n2226 GNDA.n18 241.643
R1286 GNDA.n2409 GNDA.n2408 241.643
R1287 GNDA.n2409 GNDA.n2218 241.643
R1288 GNDA.n2548 GNDA.n2547 241.643
R1289 GNDA.n2548 GNDA.n19 241.643
R1290 GNDA.n2452 GNDA.n2451 241.643
R1291 GNDA.n2452 GNDA.n32 241.643
R1292 GNDA.n2334 GNDA.n2333 241.643
R1293 GNDA.n2344 GNDA.n2343 241.643
R1294 GNDA.n2377 GNDA.n2376 241.643
R1295 GNDA.n2366 GNDA.n2365 241.643
R1296 GNDA.n2071 GNDA.n2070 241.643
R1297 GNDA.n2070 GNDA.n77 241.643
R1298 GNDA.n174 GNDA.n159 241.643
R1299 GNDA.n174 GNDA.n160 241.643
R1300 GNDA.n2360 GNDA.t234 233
R1301 GNDA.n2346 GNDA.t240 233
R1302 GNDA.n2357 GNDA.n2356 226.534
R1303 GNDA.n2355 GNDA.n2354 226.534
R1304 GNDA.n2353 GNDA.n2352 226.534
R1305 GNDA.n2351 GNDA.n2350 226.534
R1306 GNDA.n2349 GNDA.n2348 226.534
R1307 GNDA.n2249 GNDA.n2247 206.052
R1308 GNDA.n5 GNDA.n3 206.052
R1309 GNDA.n2255 GNDA.n2254 205.488
R1310 GNDA.n2253 GNDA.n2252 205.488
R1311 GNDA.n2251 GNDA.n2250 205.488
R1312 GNDA.n2249 GNDA.n2248 205.488
R1313 GNDA.n11 GNDA.n10 205.488
R1314 GNDA.n9 GNDA.n8 205.488
R1315 GNDA.n7 GNDA.n6 205.488
R1316 GNDA.n5 GNDA.n4 205.488
R1317 GNDA.n2257 GNDA.n2256 200.988
R1318 GNDA.n13 GNDA.n12 200.988
R1319 GNDA.n1961 GNDA.n116 197
R1320 GNDA.n1038 GNDA.n1015 197
R1321 GNDA.n663 GNDA.n478 197
R1322 GNDA.n1146 GNDA.n854 197
R1323 GNDA.n1287 GNDA.n509 197
R1324 GNDA.n1621 GNDA.n1620 197
R1325 GNDA.n1574 GNDA.n510 197
R1326 GNDA.n1830 GNDA.n1829 197
R1327 GNDA.n1779 GNDA.n1778 197
R1328 GNDA.n214 GNDA.n213 197
R1329 GNDA.n2033 GNDA.n111 187.249
R1330 GNDA.n1154 GNDA.n868 187.249
R1331 GNDA.n733 GNDA.n732 187.249
R1332 GNDA.n1235 GNDA.n1234 187.249
R1333 GNDA.n1376 GNDA.n581 187.249
R1334 GNDA.n1703 GNDA.n512 187.249
R1335 GNDA.n1705 GNDA.n507 187.249
R1336 GNDA.n1785 GNDA.n1783 187.249
R1337 GNDA.n1734 GNDA.n1732 187.249
R1338 GNDA.n2072 GNDA.n75 185
R1339 GNDA.n2064 GNDA.n2063 185
R1340 GNDA.n706 GNDA.n705 185
R1341 GNDA.n708 GNDA.n707 185
R1342 GNDA.n710 GNDA.n709 185
R1343 GNDA.n712 GNDA.n711 185
R1344 GNDA.n714 GNDA.n713 185
R1345 GNDA.n716 GNDA.n715 185
R1346 GNDA.n718 GNDA.n717 185
R1347 GNDA.n720 GNDA.n719 185
R1348 GNDA.n721 GNDA.n612 185
R1349 GNDA.n688 GNDA.n687 185
R1350 GNDA.n690 GNDA.n689 185
R1351 GNDA.n692 GNDA.n691 185
R1352 GNDA.n694 GNDA.n693 185
R1353 GNDA.n696 GNDA.n695 185
R1354 GNDA.n698 GNDA.n697 185
R1355 GNDA.n700 GNDA.n699 185
R1356 GNDA.n702 GNDA.n701 185
R1357 GNDA.n704 GNDA.n703 185
R1358 GNDA.n670 GNDA.n669 185
R1359 GNDA.n672 GNDA.n671 185
R1360 GNDA.n674 GNDA.n673 185
R1361 GNDA.n676 GNDA.n675 185
R1362 GNDA.n678 GNDA.n677 185
R1363 GNDA.n680 GNDA.n679 185
R1364 GNDA.n682 GNDA.n681 185
R1365 GNDA.n684 GNDA.n683 185
R1366 GNDA.n686 GNDA.n685 185
R1367 GNDA.n668 GNDA.n667 185
R1368 GNDA.n657 GNDA.n656 185
R1369 GNDA.n655 GNDA.n654 185
R1370 GNDA.n652 GNDA.n651 185
R1371 GNDA.n650 GNDA.n649 185
R1372 GNDA.n641 GNDA.n640 185
R1373 GNDA.n639 GNDA.n617 185
R1374 GNDA.n725 GNDA.n724 185
R1375 GNDA.n616 GNDA.n613 185
R1376 GNDA.n1207 GNDA.n1206 185
R1377 GNDA.n1209 GNDA.n1208 185
R1378 GNDA.n1211 GNDA.n1210 185
R1379 GNDA.n1213 GNDA.n1212 185
R1380 GNDA.n1215 GNDA.n1214 185
R1381 GNDA.n1217 GNDA.n1216 185
R1382 GNDA.n1219 GNDA.n1218 185
R1383 GNDA.n1220 GNDA.n822 185
R1384 GNDA.n1224 GNDA.n1223 185
R1385 GNDA.n1189 GNDA.n1188 185
R1386 GNDA.n1191 GNDA.n1190 185
R1387 GNDA.n1193 GNDA.n1192 185
R1388 GNDA.n1195 GNDA.n1194 185
R1389 GNDA.n1197 GNDA.n1196 185
R1390 GNDA.n1199 GNDA.n1198 185
R1391 GNDA.n1201 GNDA.n1200 185
R1392 GNDA.n1203 GNDA.n1202 185
R1393 GNDA.n1205 GNDA.n1204 185
R1394 GNDA.n1171 GNDA.n1170 185
R1395 GNDA.n1173 GNDA.n1172 185
R1396 GNDA.n1175 GNDA.n1174 185
R1397 GNDA.n1177 GNDA.n1176 185
R1398 GNDA.n1179 GNDA.n1178 185
R1399 GNDA.n1181 GNDA.n1180 185
R1400 GNDA.n1183 GNDA.n1182 185
R1401 GNDA.n1185 GNDA.n1184 185
R1402 GNDA.n1187 GNDA.n1186 185
R1403 GNDA.n1169 GNDA.n1168 185
R1404 GNDA.n845 GNDA.n844 185
R1405 GNDA.n847 GNDA.n846 185
R1406 GNDA.n842 GNDA.n841 185
R1407 GNDA.n840 GNDA.n839 185
R1408 GNDA.n829 GNDA.n828 185
R1409 GNDA.n830 GNDA.n805 185
R1410 GNDA.n1228 GNDA.n1227 185
R1411 GNDA.n804 GNDA.n802 185
R1412 GNDA.n1346 GNDA.n1285 185
R1413 GNDA.n1360 GNDA.n1359 185
R1414 GNDA.n1358 GNDA.n1286 185
R1415 GNDA.n1357 GNDA.n1356 185
R1416 GNDA.n1355 GNDA.n1354 185
R1417 GNDA.n1353 GNDA.n1352 185
R1418 GNDA.n1351 GNDA.n1350 185
R1419 GNDA.n1349 GNDA.n1348 185
R1420 GNDA.n1347 GNDA.n1262 185
R1421 GNDA.n1329 GNDA.n1328 185
R1422 GNDA.n1331 GNDA.n1330 185
R1423 GNDA.n1333 GNDA.n1332 185
R1424 GNDA.n1335 GNDA.n1334 185
R1425 GNDA.n1337 GNDA.n1336 185
R1426 GNDA.n1339 GNDA.n1338 185
R1427 GNDA.n1341 GNDA.n1340 185
R1428 GNDA.n1343 GNDA.n1342 185
R1429 GNDA.n1345 GNDA.n1344 185
R1430 GNDA.n1311 GNDA.n1310 185
R1431 GNDA.n1313 GNDA.n1312 185
R1432 GNDA.n1315 GNDA.n1314 185
R1433 GNDA.n1317 GNDA.n1316 185
R1434 GNDA.n1319 GNDA.n1318 185
R1435 GNDA.n1321 GNDA.n1320 185
R1436 GNDA.n1323 GNDA.n1322 185
R1437 GNDA.n1325 GNDA.n1324 185
R1438 GNDA.n1327 GNDA.n1326 185
R1439 GNDA.n1309 GNDA.n1308 185
R1440 GNDA.n1303 GNDA.n1302 185
R1441 GNDA.n1301 GNDA.n1300 185
R1442 GNDA.n1296 GNDA.n1295 185
R1443 GNDA.n1291 GNDA.n1270 185
R1444 GNDA.n1364 GNDA.n1363 185
R1445 GNDA.n1269 GNDA.n1267 185
R1446 GNDA.n1370 GNDA.n1369 185
R1447 GNDA.n1372 GNDA.n1371 185
R1448 GNDA.n1519 GNDA.n1518 185
R1449 GNDA.n1521 GNDA.n1473 185
R1450 GNDA.n1524 GNDA.n1523 185
R1451 GNDA.n1525 GNDA.n1472 185
R1452 GNDA.n1527 GNDA.n1526 185
R1453 GNDA.n1529 GNDA.n1471 185
R1454 GNDA.n1532 GNDA.n1531 185
R1455 GNDA.n1533 GNDA.n1470 185
R1456 GNDA.n1538 GNDA.n1537 185
R1457 GNDA.n1501 GNDA.n1478 185
R1458 GNDA.n1503 GNDA.n1502 185
R1459 GNDA.n1505 GNDA.n1477 185
R1460 GNDA.n1508 GNDA.n1507 185
R1461 GNDA.n1509 GNDA.n1476 185
R1462 GNDA.n1511 GNDA.n1510 185
R1463 GNDA.n1513 GNDA.n1475 185
R1464 GNDA.n1516 GNDA.n1515 185
R1465 GNDA.n1517 GNDA.n1474 185
R1466 GNDA.n1485 GNDA.n1458 185
R1467 GNDA.n1486 GNDA.n1484 185
R1468 GNDA.n1488 GNDA.n1487 185
R1469 GNDA.n1490 GNDA.n1481 185
R1470 GNDA.n1492 GNDA.n1491 185
R1471 GNDA.n1493 GNDA.n1480 185
R1472 GNDA.n1495 GNDA.n1494 185
R1473 GNDA.n1497 GNDA.n1479 185
R1474 GNDA.n1500 GNDA.n1499 185
R1475 GNDA.n1570 GNDA.n1569 185
R1476 GNDA.n1567 GNDA.n1566 185
R1477 GNDA.n1460 GNDA.n1459 185
R1478 GNDA.n1558 GNDA.n1557 185
R1479 GNDA.n1555 GNDA.n1463 185
R1480 GNDA.n1553 GNDA.n1552 185
R1481 GNDA.n1465 GNDA.n1464 185
R1482 GNDA.n1543 GNDA.n1542 185
R1483 GNDA.n1540 GNDA.n1469 185
R1484 GNDA.n1440 GNDA.n1439 185
R1485 GNDA.n1442 GNDA.n1397 185
R1486 GNDA.n1445 GNDA.n1444 185
R1487 GNDA.n1446 GNDA.n1396 185
R1488 GNDA.n1448 GNDA.n1447 185
R1489 GNDA.n1450 GNDA.n1395 185
R1490 GNDA.n1453 GNDA.n1452 185
R1491 GNDA.n1454 GNDA.n1394 185
R1492 GNDA.n1581 GNDA.n1580 185
R1493 GNDA.n1422 GNDA.n1402 185
R1494 GNDA.n1424 GNDA.n1423 185
R1495 GNDA.n1426 GNDA.n1401 185
R1496 GNDA.n1429 GNDA.n1428 185
R1497 GNDA.n1430 GNDA.n1400 185
R1498 GNDA.n1432 GNDA.n1431 185
R1499 GNDA.n1434 GNDA.n1399 185
R1500 GNDA.n1437 GNDA.n1436 185
R1501 GNDA.n1438 GNDA.n1398 185
R1502 GNDA.n1615 GNDA.n1614 185
R1503 GNDA.n1407 GNDA.n1381 185
R1504 GNDA.n1409 GNDA.n1408 185
R1505 GNDA.n1411 GNDA.n1405 185
R1506 GNDA.n1413 GNDA.n1412 185
R1507 GNDA.n1414 GNDA.n1404 185
R1508 GNDA.n1416 GNDA.n1415 185
R1509 GNDA.n1418 GNDA.n1403 185
R1510 GNDA.n1421 GNDA.n1420 185
R1511 GNDA.n1613 GNDA.n1380 185
R1512 GNDA.n1611 GNDA.n1610 185
R1513 GNDA.n1384 GNDA.n1383 185
R1514 GNDA.n1601 GNDA.n1600 185
R1515 GNDA.n1598 GNDA.n1387 185
R1516 GNDA.n1596 GNDA.n1595 185
R1517 GNDA.n1389 GNDA.n1388 185
R1518 GNDA.n1586 GNDA.n1585 185
R1519 GNDA.n1583 GNDA.n1393 185
R1520 GNDA.n425 GNDA.n424 185
R1521 GNDA.n427 GNDA.n382 185
R1522 GNDA.n430 GNDA.n429 185
R1523 GNDA.n431 GNDA.n381 185
R1524 GNDA.n433 GNDA.n432 185
R1525 GNDA.n435 GNDA.n380 185
R1526 GNDA.n438 GNDA.n437 185
R1527 GNDA.n439 GNDA.n379 185
R1528 GNDA.n1739 GNDA.n1738 185
R1529 GNDA.n407 GNDA.n387 185
R1530 GNDA.n409 GNDA.n408 185
R1531 GNDA.n411 GNDA.n386 185
R1532 GNDA.n414 GNDA.n413 185
R1533 GNDA.n415 GNDA.n385 185
R1534 GNDA.n417 GNDA.n416 185
R1535 GNDA.n419 GNDA.n384 185
R1536 GNDA.n422 GNDA.n421 185
R1537 GNDA.n423 GNDA.n383 185
R1538 GNDA.n1773 GNDA.n1772 185
R1539 GNDA.n392 GNDA.n367 185
R1540 GNDA.n394 GNDA.n393 185
R1541 GNDA.n396 GNDA.n390 185
R1542 GNDA.n398 GNDA.n397 185
R1543 GNDA.n399 GNDA.n389 185
R1544 GNDA.n401 GNDA.n400 185
R1545 GNDA.n403 GNDA.n388 185
R1546 GNDA.n406 GNDA.n405 185
R1547 GNDA.n306 GNDA.n305 185
R1548 GNDA.n308 GNDA.n263 185
R1549 GNDA.n311 GNDA.n310 185
R1550 GNDA.n312 GNDA.n262 185
R1551 GNDA.n314 GNDA.n313 185
R1552 GNDA.n316 GNDA.n261 185
R1553 GNDA.n319 GNDA.n318 185
R1554 GNDA.n320 GNDA.n260 185
R1555 GNDA.n1790 GNDA.n1789 185
R1556 GNDA.n288 GNDA.n268 185
R1557 GNDA.n290 GNDA.n289 185
R1558 GNDA.n292 GNDA.n267 185
R1559 GNDA.n295 GNDA.n294 185
R1560 GNDA.n296 GNDA.n266 185
R1561 GNDA.n298 GNDA.n297 185
R1562 GNDA.n300 GNDA.n265 185
R1563 GNDA.n303 GNDA.n302 185
R1564 GNDA.n304 GNDA.n264 185
R1565 GNDA.n1824 GNDA.n1823 185
R1566 GNDA.n273 GNDA.n248 185
R1567 GNDA.n275 GNDA.n274 185
R1568 GNDA.n277 GNDA.n271 185
R1569 GNDA.n279 GNDA.n278 185
R1570 GNDA.n280 GNDA.n270 185
R1571 GNDA.n282 GNDA.n281 185
R1572 GNDA.n284 GNDA.n269 185
R1573 GNDA.n287 GNDA.n286 185
R1574 GNDA.n1822 GNDA.n247 185
R1575 GNDA.n1820 GNDA.n1819 185
R1576 GNDA.n251 GNDA.n250 185
R1577 GNDA.n1810 GNDA.n1809 185
R1578 GNDA.n1807 GNDA.n254 185
R1579 GNDA.n1805 GNDA.n1804 185
R1580 GNDA.n256 GNDA.n255 185
R1581 GNDA.n1795 GNDA.n1794 185
R1582 GNDA.n1792 GNDA.n259 185
R1583 GNDA.n1771 GNDA.n366 185
R1584 GNDA.n1769 GNDA.n1768 185
R1585 GNDA.n370 GNDA.n369 185
R1586 GNDA.n1759 GNDA.n1758 185
R1587 GNDA.n1756 GNDA.n373 185
R1588 GNDA.n1754 GNDA.n1753 185
R1589 GNDA.n375 GNDA.n374 185
R1590 GNDA.n1744 GNDA.n1743 185
R1591 GNDA.n1741 GNDA.n378 185
R1592 GNDA.n962 GNDA.n961 185
R1593 GNDA.n960 GNDA.n959 185
R1594 GNDA.n958 GNDA.n957 185
R1595 GNDA.n956 GNDA.n955 185
R1596 GNDA.n954 GNDA.n953 185
R1597 GNDA.n952 GNDA.n951 185
R1598 GNDA.n950 GNDA.n949 185
R1599 GNDA.n948 GNDA.n947 185
R1600 GNDA.n946 GNDA.n63 185
R1601 GNDA.n980 GNDA.n979 185
R1602 GNDA.n978 GNDA.n977 185
R1603 GNDA.n976 GNDA.n975 185
R1604 GNDA.n974 GNDA.n973 185
R1605 GNDA.n972 GNDA.n971 185
R1606 GNDA.n970 GNDA.n969 185
R1607 GNDA.n968 GNDA.n967 185
R1608 GNDA.n966 GNDA.n965 185
R1609 GNDA.n964 GNDA.n963 185
R1610 GNDA.n1009 GNDA.n997 185
R1611 GNDA.n996 GNDA.n995 185
R1612 GNDA.n994 GNDA.n993 185
R1613 GNDA.n992 GNDA.n991 185
R1614 GNDA.n990 GNDA.n989 185
R1615 GNDA.n988 GNDA.n987 185
R1616 GNDA.n986 GNDA.n985 185
R1617 GNDA.n984 GNDA.n983 185
R1618 GNDA.n982 GNDA.n981 185
R1619 GNDA.n1011 GNDA.n1010 185
R1620 GNDA.n999 GNDA.n998 185
R1621 GNDA.n1000 GNDA.n46 185
R1622 GNDA.n2098 GNDA.n2097 185
R1623 GNDA.n2081 GNDA.n45 185
R1624 GNDA.n2085 GNDA.n2084 185
R1625 GNDA.n2083 GNDA.n2080 185
R1626 GNDA.n66 GNDA.n64 185
R1627 GNDA.n2094 GNDA.n2093 185
R1628 GNDA.n2015 GNDA.n2014 185
R1629 GNDA.n2017 GNDA.n2016 185
R1630 GNDA.n2019 GNDA.n2018 185
R1631 GNDA.n2021 GNDA.n2020 185
R1632 GNDA.n2023 GNDA.n2022 185
R1633 GNDA.n2025 GNDA.n2024 185
R1634 GNDA.n2027 GNDA.n2026 185
R1635 GNDA.n2029 GNDA.n2028 185
R1636 GNDA.n2030 GNDA.n102 185
R1637 GNDA.n1997 GNDA.n1996 185
R1638 GNDA.n1999 GNDA.n1998 185
R1639 GNDA.n2001 GNDA.n2000 185
R1640 GNDA.n2003 GNDA.n2002 185
R1641 GNDA.n2005 GNDA.n2004 185
R1642 GNDA.n2007 GNDA.n2006 185
R1643 GNDA.n2009 GNDA.n2008 185
R1644 GNDA.n2011 GNDA.n2010 185
R1645 GNDA.n2013 GNDA.n2012 185
R1646 GNDA.n1979 GNDA.n1978 185
R1647 GNDA.n1981 GNDA.n1980 185
R1648 GNDA.n1983 GNDA.n1982 185
R1649 GNDA.n1985 GNDA.n1984 185
R1650 GNDA.n1987 GNDA.n1986 185
R1651 GNDA.n1989 GNDA.n1988 185
R1652 GNDA.n1991 GNDA.n1990 185
R1653 GNDA.n1993 GNDA.n1992 185
R1654 GNDA.n1995 GNDA.n1994 185
R1655 GNDA.n1977 GNDA.n1976 185
R1656 GNDA.n120 GNDA.n119 185
R1657 GNDA.n118 GNDA.n85 185
R1658 GNDA.n2056 GNDA.n2055 185
R1659 GNDA.n2039 GNDA.n84 185
R1660 GNDA.n2043 GNDA.n2042 185
R1661 GNDA.n2041 GNDA.n2038 185
R1662 GNDA.n105 GNDA.n103 185
R1663 GNDA.n2052 GNDA.n2051 185
R1664 GNDA.n2214 GNDA.n2213 185
R1665 GNDA.n2212 GNDA.n2131 185
R1666 GNDA.n2210 GNDA.n2132 185
R1667 GNDA.n2207 GNDA.n2133 185
R1668 GNDA.n2206 GNDA.n2134 185
R1669 GNDA.n2203 GNDA.n2135 185
R1670 GNDA.n2202 GNDA.n2136 185
R1671 GNDA.n2199 GNDA.n2137 185
R1672 GNDA.n2198 GNDA.n2138 185
R1673 GNDA.n2195 GNDA.n2139 185
R1674 GNDA.n2317 GNDA.n2312 185
R1675 GNDA.n2280 GNDA.n2275 185
R1676 GNDA.n2395 GNDA.n2221 185
R1677 GNDA.n2382 GNDA.n2381 185
R1678 GNDA.n2386 GNDA.n2232 185
R1679 GNDA.n2270 GNDA.n2269 185
R1680 GNDA.n2267 GNDA.n2264 185
R1681 GNDA.n2225 GNDA.n2224 185
R1682 GNDA.n2406 GNDA.n2405 185
R1683 GNDA.n2404 GNDA.n2401 185
R1684 GNDA.n2422 GNDA.n2421 185
R1685 GNDA.n2420 GNDA.n2118 185
R1686 GNDA.n2332 GNDA.n2246 185
R1687 GNDA.n2342 GNDA.n2337 185
R1688 GNDA.n2375 GNDA.n2240 185
R1689 GNDA.n2364 GNDA.n2362 185
R1690 GNDA.n2545 GNDA.n2544 185
R1691 GNDA.n2543 GNDA.n2540 185
R1692 GNDA.n2449 GNDA.n2448 185
R1693 GNDA.n2447 GNDA.n2441 185
R1694 GNDA.n2533 GNDA.n2532 185
R1695 GNDA.n2531 GNDA.n2500 185
R1696 GNDA.n2529 GNDA.n2501 185
R1697 GNDA.n2526 GNDA.n2502 185
R1698 GNDA.n2525 GNDA.n2503 185
R1699 GNDA.n2522 GNDA.n2504 185
R1700 GNDA.n2521 GNDA.n2505 185
R1701 GNDA.n2518 GNDA.n2506 185
R1702 GNDA.n2517 GNDA.n2507 185
R1703 GNDA.n2514 GNDA.n2508 185
R1704 GNDA.n2493 GNDA.n2492 185
R1705 GNDA.n2491 GNDA.n2456 185
R1706 GNDA.n2489 GNDA.n2457 185
R1707 GNDA.n2486 GNDA.n2458 185
R1708 GNDA.n2485 GNDA.n2459 185
R1709 GNDA.n2482 GNDA.n2460 185
R1710 GNDA.n2481 GNDA.n2461 185
R1711 GNDA.n2478 GNDA.n2462 185
R1712 GNDA.n2477 GNDA.n2463 185
R1713 GNDA.n2474 GNDA.n2464 185
R1714 GNDA.n2156 GNDA.n2151 185
R1715 GNDA.n2158 GNDA.n2157 185
R1716 GNDA.n2149 GNDA.n2148 185
R1717 GNDA.n2165 GNDA.n2164 185
R1718 GNDA.n2166 GNDA.n2147 185
R1719 GNDA.n2168 GNDA.n2167 185
R1720 GNDA.n2145 GNDA.n2144 185
R1721 GNDA.n2175 GNDA.n2174 185
R1722 GNDA.n2176 GNDA.n2143 185
R1723 GNDA.n2178 GNDA.n2177 185
R1724 GNDA.n162 GNDA.n70 185
R1725 GNDA.n170 GNDA.n162 185
R1726 GNDA.n168 GNDA.n70 185
R1727 GNDA.n168 GNDA.n167 185
R1728 GNDA.t221 GNDA.n144 183.948
R1729 GNDA.n1882 GNDA.n1881 183.948
R1730 GNDA.t221 GNDA.n143 180.013
R1731 GNDA.n1881 GNDA.n1880 180.013
R1732 GNDA.t239 GNDA.t159 179.593
R1733 GNDA.t5 GNDA.t245 179.593
R1734 GNDA.t15 GNDA.t224 179.593
R1735 GNDA.t233 GNDA.t126 179.593
R1736 GNDA.n1938 GNDA.n139 175.546
R1737 GNDA.n1943 GNDA.n139 175.546
R1738 GNDA.n1943 GNDA.n136 175.546
R1739 GNDA.n1947 GNDA.n136 175.546
R1740 GNDA.n1948 GNDA.n1947 175.546
R1741 GNDA.n1949 GNDA.n1948 175.546
R1742 GNDA.n1949 GNDA.n134 175.546
R1743 GNDA.n1954 GNDA.n134 175.546
R1744 GNDA.n1954 GNDA.n131 175.546
R1745 GNDA.n1958 GNDA.n131 175.546
R1746 GNDA.n1959 GNDA.n1958 175.546
R1747 GNDA.n1085 GNDA.n1061 175.546
R1748 GNDA.n1081 GNDA.n1080 175.546
R1749 GNDA.n1078 GNDA.n1064 175.546
R1750 GNDA.n1074 GNDA.n1073 175.546
R1751 GNDA.n1071 GNDA.n1068 175.546
R1752 GNDA.n2033 GNDA.n106 175.546
R1753 GNDA.n2049 GNDA.n106 175.546
R1754 GNDA.n2049 GNDA.n107 175.546
R1755 GNDA.n2045 GNDA.n107 175.546
R1756 GNDA.n2045 GNDA.n81 175.546
R1757 GNDA.n2058 GNDA.n81 175.546
R1758 GNDA.n2058 GNDA.n82 175.546
R1759 GNDA.n122 GNDA.n82 175.546
R1760 GNDA.n122 GNDA.n115 175.546
R1761 GNDA.n1974 GNDA.n115 175.546
R1762 GNDA.n1974 GNDA.n116 175.546
R1763 GNDA.n1090 GNDA.n1059 175.546
R1764 GNDA.n1057 GNDA.n924 175.546
R1765 GNDA.n1053 GNDA.n1051 175.546
R1766 GNDA.n1049 GNDA.n931 175.546
R1767 GNDA.n1045 GNDA.n1043 175.546
R1768 GNDA.n1092 GNDA.n922 175.546
R1769 GNDA.n927 GNDA.n926 175.546
R1770 GNDA.n932 GNDA.n929 175.546
R1771 GNDA.n935 GNDA.n934 175.546
R1772 GNDA.n939 GNDA.n937 175.546
R1773 GNDA.n1113 GNDA.n911 175.546
R1774 GNDA.n1109 GNDA.n1108 175.546
R1775 GNDA.n1106 GNDA.n914 175.546
R1776 GNDA.n1102 GNDA.n1101 175.546
R1777 GNDA.n1099 GNDA.n917 175.546
R1778 GNDA.n868 GNDA.n67 175.546
R1779 GNDA.n2091 GNDA.n67 175.546
R1780 GNDA.n2091 GNDA.n68 175.546
R1781 GNDA.n2087 GNDA.n68 175.546
R1782 GNDA.n2087 GNDA.n42 175.546
R1783 GNDA.n2100 GNDA.n42 175.546
R1784 GNDA.n2100 GNDA.n43 175.546
R1785 GNDA.n1002 GNDA.n43 175.546
R1786 GNDA.n1007 GNDA.n1002 175.546
R1787 GNDA.n1007 GNDA.n941 175.546
R1788 GNDA.n1015 GNDA.n941 175.546
R1789 GNDA.n1125 GNDA.n879 175.546
R1790 GNDA.n1129 GNDA.n1127 175.546
R1791 GNDA.n1137 GNDA.n875 175.546
R1792 GNDA.n1141 GNDA.n1139 175.546
R1793 GNDA.n1151 GNDA.n871 175.546
R1794 GNDA.n1910 GNDA.n195 175.546
R1795 GNDA.n455 GNDA.n453 175.546
R1796 GNDA.n463 GNDA.n447 175.546
R1797 GNDA.n468 GNDA.n465 175.546
R1798 GNDA.n466 GNDA.n444 175.546
R1799 GNDA.n1935 GNDA.n183 175.546
R1800 GNDA.n1931 GNDA.n183 175.546
R1801 GNDA.n1931 GNDA.n186 175.546
R1802 GNDA.n1927 GNDA.n186 175.546
R1803 GNDA.n1927 GNDA.n188 175.546
R1804 GNDA.n1923 GNDA.n188 175.546
R1805 GNDA.n1923 GNDA.n190 175.546
R1806 GNDA.n1919 GNDA.n190 175.546
R1807 GNDA.n1919 GNDA.n192 175.546
R1808 GNDA.n1915 GNDA.n192 175.546
R1809 GNDA.n1915 GNDA.n1913 175.546
R1810 GNDA.n728 GNDA.n727 175.546
R1811 GNDA.n643 GNDA.n638 175.546
R1812 GNDA.n647 GNDA.n645 175.546
R1813 GNDA.n659 GNDA.n636 175.546
R1814 GNDA.n665 GNDA.n661 175.546
R1815 GNDA.n593 GNDA.n592 175.546
R1816 GNDA.n597 GNDA.n596 175.546
R1817 GNDA.n601 GNDA.n600 175.546
R1818 GNDA.n605 GNDA.n604 175.546
R1819 GNDA.n607 GNDA.n589 175.546
R1820 GNDA.n590 GNDA.n589 175.546
R1821 GNDA.n1123 GNDA.n1121 175.546
R1822 GNDA.n1131 GNDA.n877 175.546
R1823 GNDA.n1135 GNDA.n1133 175.546
R1824 GNDA.n1143 GNDA.n873 175.546
R1825 GNDA.n1149 GNDA.n1145 175.546
R1826 GNDA.n890 GNDA.n888 175.546
R1827 GNDA.n894 GNDA.n885 175.546
R1828 GNDA.n898 GNDA.n896 175.546
R1829 GNDA.n902 GNDA.n883 175.546
R1830 GNDA.n906 GNDA.n904 175.546
R1831 GNDA.n1234 GNDA.n800 175.546
R1832 GNDA.n1230 GNDA.n800 175.546
R1833 GNDA.n1230 GNDA.n801 175.546
R1834 GNDA.n832 GNDA.n801 175.546
R1835 GNDA.n836 GNDA.n832 175.546
R1836 GNDA.n836 GNDA.n827 175.546
R1837 GNDA.n849 GNDA.n827 175.546
R1838 GNDA.n849 GNDA.n825 175.546
R1839 GNDA.n853 GNDA.n825 175.546
R1840 GNDA.n1166 GNDA.n853 175.546
R1841 GNDA.n1166 GNDA.n854 175.546
R1842 GNDA.n1252 GNDA.n795 175.546
R1843 GNDA.n1250 GNDA.n1249 175.546
R1844 GNDA.n1246 GNDA.n1245 175.546
R1845 GNDA.n1242 GNDA.n1241 175.546
R1846 GNDA.n1238 GNDA.n790 175.546
R1847 GNDA.n798 GNDA.n790 175.546
R1848 GNDA.n487 GNDA.n486 175.546
R1849 GNDA.n492 GNDA.n489 175.546
R1850 GNDA.n495 GNDA.n494 175.546
R1851 GNDA.n500 GNDA.n497 175.546
R1852 GNDA.n503 GNDA.n502 175.546
R1853 GNDA.n766 GNDA.n741 175.546
R1854 GNDA.n762 GNDA.n761 175.546
R1855 GNDA.n759 GNDA.n744 175.546
R1856 GNDA.n755 GNDA.n754 175.546
R1857 GNDA.n752 GNDA.n749 175.546
R1858 GNDA.n1263 GNDA.n580 175.546
R1859 GNDA.n1367 GNDA.n1366 175.546
R1860 GNDA.n1293 GNDA.n1292 175.546
R1861 GNDA.n1298 GNDA.n1297 175.546
R1862 GNDA.n1306 GNDA.n1305 175.546
R1863 GNDA.n773 GNDA.n772 175.546
R1864 GNDA.n777 GNDA.n776 175.546
R1865 GNDA.n781 GNDA.n780 175.546
R1866 GNDA.n783 GNDA.n739 175.546
R1867 GNDA.n787 GNDA.n583 175.546
R1868 GNDA.n1644 GNDA.n563 175.546
R1869 GNDA.n1640 GNDA.n563 175.546
R1870 GNDA.n1640 GNDA.n565 175.546
R1871 GNDA.n1636 GNDA.n565 175.546
R1872 GNDA.n1636 GNDA.n1634 175.546
R1873 GNDA.n1634 GNDA.n1633 175.546
R1874 GNDA.n1633 GNDA.n568 175.546
R1875 GNDA.n1629 GNDA.n568 175.546
R1876 GNDA.n1629 GNDA.n570 175.546
R1877 GNDA.n1625 GNDA.n570 175.546
R1878 GNDA.n1625 GNDA.n573 175.546
R1879 GNDA.n1663 GNDA.n554 175.546
R1880 GNDA.n1659 GNDA.n1658 175.546
R1881 GNDA.n1656 GNDA.n557 175.546
R1882 GNDA.n1652 GNDA.n1651 175.546
R1883 GNDA.n1649 GNDA.n560 175.546
R1884 GNDA.n1588 GNDA.n1392 175.546
R1885 GNDA.n1592 GNDA.n1590 175.546
R1886 GNDA.n1603 GNDA.n1386 175.546
R1887 GNDA.n1607 GNDA.n1605 175.546
R1888 GNDA.n1618 GNDA.n1379 175.546
R1889 GNDA.n1675 GNDA.n522 175.546
R1890 GNDA.n1679 GNDA.n1677 175.546
R1891 GNDA.n1687 GNDA.n518 175.546
R1892 GNDA.n1691 GNDA.n1689 175.546
R1893 GNDA.n1700 GNDA.n514 175.546
R1894 GNDA.n1726 GNDA.n1725 175.546
R1895 GNDA.n1722 GNDA.n1721 175.546
R1896 GNDA.n1719 GNDA.n491 175.546
R1897 GNDA.n1715 GNDA.n1713 175.546
R1898 GNDA.n1711 GNDA.n499 175.546
R1899 GNDA.n533 GNDA.n531 175.546
R1900 GNDA.n537 GNDA.n528 175.546
R1901 GNDA.n541 GNDA.n539 175.546
R1902 GNDA.n545 GNDA.n526 175.546
R1903 GNDA.n549 GNDA.n547 175.546
R1904 GNDA.n1545 GNDA.n1468 175.546
R1905 GNDA.n1549 GNDA.n1547 175.546
R1906 GNDA.n1560 GNDA.n1462 175.546
R1907 GNDA.n1564 GNDA.n1562 175.546
R1908 GNDA.n1572 GNDA.n1456 175.546
R1909 GNDA.n1673 GNDA.n1671 175.546
R1910 GNDA.n1681 GNDA.n520 175.546
R1911 GNDA.n1685 GNDA.n1683 175.546
R1912 GNDA.n1693 GNDA.n516 175.546
R1913 GNDA.n1698 GNDA.n1695 175.546
R1914 GNDA.n1855 GNDA.n235 175.546
R1915 GNDA.n1851 GNDA.n235 175.546
R1916 GNDA.n1851 GNDA.n237 175.546
R1917 GNDA.n1847 GNDA.n237 175.546
R1918 GNDA.n1847 GNDA.n238 175.546
R1919 GNDA.n1843 GNDA.n238 175.546
R1920 GNDA.n1843 GNDA.n1842 175.546
R1921 GNDA.n1842 GNDA.n240 175.546
R1922 GNDA.n1838 GNDA.n240 175.546
R1923 GNDA.n1838 GNDA.n242 175.546
R1924 GNDA.n1833 GNDA.n242 175.546
R1925 GNDA.n1879 GNDA.n222 175.546
R1926 GNDA.n1875 GNDA.n222 175.546
R1927 GNDA.n1875 GNDA.n225 175.546
R1928 GNDA.n1871 GNDA.n225 175.546
R1929 GNDA.n1871 GNDA.n227 175.546
R1930 GNDA.n1867 GNDA.n227 175.546
R1931 GNDA.n1867 GNDA.n229 175.546
R1932 GNDA.n1863 GNDA.n229 175.546
R1933 GNDA.n1863 GNDA.n231 175.546
R1934 GNDA.n1859 GNDA.n231 175.546
R1935 GNDA.n1859 GNDA.n233 175.546
R1936 GNDA.n1797 GNDA.n258 175.546
R1937 GNDA.n1801 GNDA.n1799 175.546
R1938 GNDA.n1812 GNDA.n253 175.546
R1939 GNDA.n1816 GNDA.n1814 175.546
R1940 GNDA.n1827 GNDA.n246 175.546
R1941 GNDA.n340 GNDA.n221 175.546
R1942 GNDA.n340 GNDA.n335 175.546
R1943 GNDA.n346 GNDA.n335 175.546
R1944 GNDA.n347 GNDA.n346 175.546
R1945 GNDA.n347 GNDA.n331 175.546
R1946 GNDA.n353 GNDA.n331 175.546
R1947 GNDA.n354 GNDA.n353 175.546
R1948 GNDA.n354 GNDA.n328 175.546
R1949 GNDA.n360 GNDA.n328 175.546
R1950 GNDA.n360 GNDA.n324 175.546
R1951 GNDA.n1782 GNDA.n324 175.546
R1952 GNDA.n1908 GNDA.n197 175.546
R1953 GNDA.n457 GNDA.n450 175.546
R1954 GNDA.n461 GNDA.n459 175.546
R1955 GNDA.n470 GNDA.n445 175.546
R1956 GNDA.n474 GNDA.n472 175.546
R1957 GNDA.n1905 GNDA.n198 175.546
R1958 GNDA.n1901 GNDA.n198 175.546
R1959 GNDA.n1901 GNDA.n201 175.546
R1960 GNDA.n1897 GNDA.n201 175.546
R1961 GNDA.n1897 GNDA.n204 175.546
R1962 GNDA.n1892 GNDA.n204 175.546
R1963 GNDA.n1892 GNDA.n207 175.546
R1964 GNDA.n1888 GNDA.n207 175.546
R1965 GNDA.n1888 GNDA.n216 175.546
R1966 GNDA.n1884 GNDA.n216 175.546
R1967 GNDA.n1884 GNDA.n218 175.546
R1968 GNDA.n1746 GNDA.n377 175.546
R1969 GNDA.n1750 GNDA.n1748 175.546
R1970 GNDA.n1761 GNDA.n372 175.546
R1971 GNDA.n1765 GNDA.n1763 175.546
R1972 GNDA.n1776 GNDA.n365 175.546
R1973 GNDA.n339 GNDA.n338 175.546
R1974 GNDA.n343 GNDA.n339 175.546
R1975 GNDA.n343 GNDA.n333 175.546
R1976 GNDA.n349 GNDA.n333 175.546
R1977 GNDA.n350 GNDA.n349 175.546
R1978 GNDA.n350 GNDA.n330 175.546
R1979 GNDA.n356 GNDA.n330 175.546
R1980 GNDA.n357 GNDA.n356 175.546
R1981 GNDA.n357 GNDA.n326 175.546
R1982 GNDA.n363 GNDA.n326 175.546
R1983 GNDA.n1780 GNDA.n363 175.546
R1984 GNDA.t221 GNDA.n148 172.876
R1985 GNDA.t221 GNDA.n145 172.615
R1986 GNDA.n2378 GNDA.t98 164.626
R1987 GNDA.n2378 GNDA.t96 164.626
R1988 GNDA.n669 GNDA.n668 163.333
R1989 GNDA.n1170 GNDA.n1169 163.333
R1990 GNDA.n1310 GNDA.n1309 163.333
R1991 GNDA.n1569 GNDA.n1458 163.333
R1992 GNDA.n1614 GNDA.n1613 163.333
R1993 GNDA.n1772 GNDA.n1771 163.333
R1994 GNDA.n1823 GNDA.n1822 163.333
R1995 GNDA.n1010 GNDA.n1009 163.333
R1996 GNDA.n1978 GNDA.n1977 163.333
R1997 GNDA.n2388 GNDA.n2387 152
R1998 GNDA.n2266 GNDA.n2265 152
R1999 GNDA.n701 GNDA.n700 150
R2000 GNDA.n697 GNDA.n696 150
R2001 GNDA.n693 GNDA.n692 150
R2002 GNDA.n689 GNDA.n688 150
R2003 GNDA.n685 GNDA.n684 150
R2004 GNDA.n681 GNDA.n680 150
R2005 GNDA.n677 GNDA.n676 150
R2006 GNDA.n673 GNDA.n672 150
R2007 GNDA.n724 GNDA.n616 150
R2008 GNDA.n640 GNDA.n617 150
R2009 GNDA.n651 GNDA.n650 150
R2010 GNDA.n656 GNDA.n655 150
R2011 GNDA.n709 GNDA.n708 150
R2012 GNDA.n713 GNDA.n712 150
R2013 GNDA.n717 GNDA.n716 150
R2014 GNDA.n721 GNDA.n720 150
R2015 GNDA.n1202 GNDA.n1201 150
R2016 GNDA.n1198 GNDA.n1197 150
R2017 GNDA.n1194 GNDA.n1193 150
R2018 GNDA.n1190 GNDA.n1189 150
R2019 GNDA.n1186 GNDA.n1185 150
R2020 GNDA.n1182 GNDA.n1181 150
R2021 GNDA.n1178 GNDA.n1177 150
R2022 GNDA.n1174 GNDA.n1173 150
R2023 GNDA.n1227 GNDA.n804 150
R2024 GNDA.n828 GNDA.n805 150
R2025 GNDA.n841 GNDA.n840 150
R2026 GNDA.n846 GNDA.n845 150
R2027 GNDA.n1210 GNDA.n1209 150
R2028 GNDA.n1214 GNDA.n1213 150
R2029 GNDA.n1218 GNDA.n1217 150
R2030 GNDA.n1224 GNDA.n822 150
R2031 GNDA.n1342 GNDA.n1341 150
R2032 GNDA.n1338 GNDA.n1337 150
R2033 GNDA.n1334 GNDA.n1333 150
R2034 GNDA.n1330 GNDA.n1329 150
R2035 GNDA.n1326 GNDA.n1325 150
R2036 GNDA.n1322 GNDA.n1321 150
R2037 GNDA.n1318 GNDA.n1317 150
R2038 GNDA.n1314 GNDA.n1313 150
R2039 GNDA.n1371 GNDA.n1370 150
R2040 GNDA.n1363 GNDA.n1269 150
R2041 GNDA.n1295 GNDA.n1270 150
R2042 GNDA.n1302 GNDA.n1301 150
R2043 GNDA.n1360 GNDA.n1286 150
R2044 GNDA.n1356 GNDA.n1355 150
R2045 GNDA.n1352 GNDA.n1351 150
R2046 GNDA.n1348 GNDA.n1347 150
R2047 GNDA.n1515 GNDA.n1513 150
R2048 GNDA.n1511 GNDA.n1476 150
R2049 GNDA.n1507 GNDA.n1505 150
R2050 GNDA.n1503 GNDA.n1478 150
R2051 GNDA.n1499 GNDA.n1497 150
R2052 GNDA.n1495 GNDA.n1480 150
R2053 GNDA.n1491 GNDA.n1490 150
R2054 GNDA.n1488 GNDA.n1484 150
R2055 GNDA.n1542 GNDA.n1540 150
R2056 GNDA.n1553 GNDA.n1464 150
R2057 GNDA.n1557 GNDA.n1555 150
R2058 GNDA.n1567 GNDA.n1459 150
R2059 GNDA.n1523 GNDA.n1521 150
R2060 GNDA.n1527 GNDA.n1472 150
R2061 GNDA.n1531 GNDA.n1529 150
R2062 GNDA.n1538 GNDA.n1470 150
R2063 GNDA.n1436 GNDA.n1434 150
R2064 GNDA.n1432 GNDA.n1400 150
R2065 GNDA.n1428 GNDA.n1426 150
R2066 GNDA.n1424 GNDA.n1402 150
R2067 GNDA.n1420 GNDA.n1418 150
R2068 GNDA.n1416 GNDA.n1404 150
R2069 GNDA.n1412 GNDA.n1411 150
R2070 GNDA.n1409 GNDA.n1407 150
R2071 GNDA.n1585 GNDA.n1583 150
R2072 GNDA.n1596 GNDA.n1388 150
R2073 GNDA.n1600 GNDA.n1598 150
R2074 GNDA.n1611 GNDA.n1383 150
R2075 GNDA.n1444 GNDA.n1442 150
R2076 GNDA.n1448 GNDA.n1396 150
R2077 GNDA.n1452 GNDA.n1450 150
R2078 GNDA.n1581 GNDA.n1394 150
R2079 GNDA.n421 GNDA.n419 150
R2080 GNDA.n417 GNDA.n385 150
R2081 GNDA.n413 GNDA.n411 150
R2082 GNDA.n409 GNDA.n387 150
R2083 GNDA.n405 GNDA.n403 150
R2084 GNDA.n401 GNDA.n389 150
R2085 GNDA.n397 GNDA.n396 150
R2086 GNDA.n394 GNDA.n392 150
R2087 GNDA.n1743 GNDA.n1741 150
R2088 GNDA.n1754 GNDA.n374 150
R2089 GNDA.n1758 GNDA.n1756 150
R2090 GNDA.n1769 GNDA.n369 150
R2091 GNDA.n429 GNDA.n427 150
R2092 GNDA.n433 GNDA.n381 150
R2093 GNDA.n437 GNDA.n435 150
R2094 GNDA.n1739 GNDA.n379 150
R2095 GNDA.n302 GNDA.n300 150
R2096 GNDA.n298 GNDA.n266 150
R2097 GNDA.n294 GNDA.n292 150
R2098 GNDA.n290 GNDA.n268 150
R2099 GNDA.n286 GNDA.n284 150
R2100 GNDA.n282 GNDA.n270 150
R2101 GNDA.n278 GNDA.n277 150
R2102 GNDA.n275 GNDA.n273 150
R2103 GNDA.n1794 GNDA.n1792 150
R2104 GNDA.n1805 GNDA.n255 150
R2105 GNDA.n1809 GNDA.n1807 150
R2106 GNDA.n1820 GNDA.n250 150
R2107 GNDA.n310 GNDA.n308 150
R2108 GNDA.n314 GNDA.n262 150
R2109 GNDA.n318 GNDA.n316 150
R2110 GNDA.n1790 GNDA.n260 150
R2111 GNDA.n967 GNDA.n966 150
R2112 GNDA.n971 GNDA.n970 150
R2113 GNDA.n975 GNDA.n974 150
R2114 GNDA.n979 GNDA.n978 150
R2115 GNDA.n983 GNDA.n982 150
R2116 GNDA.n987 GNDA.n986 150
R2117 GNDA.n991 GNDA.n990 150
R2118 GNDA.n995 GNDA.n994 150
R2119 GNDA.n2094 GNDA.n64 150
R2120 GNDA.n2084 GNDA.n2083 150
R2121 GNDA.n2097 GNDA.n45 150
R2122 GNDA.n998 GNDA.n46 150
R2123 GNDA.n959 GNDA.n958 150
R2124 GNDA.n955 GNDA.n954 150
R2125 GNDA.n951 GNDA.n950 150
R2126 GNDA.n947 GNDA.n63 150
R2127 GNDA.n2010 GNDA.n2009 150
R2128 GNDA.n2006 GNDA.n2005 150
R2129 GNDA.n2002 GNDA.n2001 150
R2130 GNDA.n1998 GNDA.n1997 150
R2131 GNDA.n1994 GNDA.n1993 150
R2132 GNDA.n1990 GNDA.n1989 150
R2133 GNDA.n1986 GNDA.n1985 150
R2134 GNDA.n1982 GNDA.n1981 150
R2135 GNDA.n2052 GNDA.n103 150
R2136 GNDA.n2042 GNDA.n2041 150
R2137 GNDA.n2055 GNDA.n84 150
R2138 GNDA.n119 GNDA.n85 150
R2139 GNDA.n2018 GNDA.n2017 150
R2140 GNDA.n2022 GNDA.n2021 150
R2141 GNDA.n2026 GNDA.n2025 150
R2142 GNDA.n2028 GNDA.n102 150
R2143 GNDA.n2157 GNDA.n2156 150
R2144 GNDA.n2157 GNDA.n2148 150
R2145 GNDA.n2165 GNDA.n2148 150
R2146 GNDA.n2166 GNDA.n2165 150
R2147 GNDA.n2167 GNDA.n2144 150
R2148 GNDA.n2175 GNDA.n2144 150
R2149 GNDA.n2176 GNDA.n2175 150
R2150 GNDA.n2177 GNDA.n2176 150
R2151 GNDA.n2214 GNDA.n2131 150
R2152 GNDA.n2132 GNDA.n2131 150
R2153 GNDA.n2133 GNDA.n2132 150
R2154 GNDA.n2134 GNDA.n2133 150
R2155 GNDA.n2136 GNDA.n2135 150
R2156 GNDA.n2137 GNDA.n2136 150
R2157 GNDA.n2138 GNDA.n2137 150
R2158 GNDA.n2139 GNDA.n2138 150
R2159 GNDA.n2533 GNDA.n2500 150
R2160 GNDA.n2501 GNDA.n2500 150
R2161 GNDA.n2502 GNDA.n2501 150
R2162 GNDA.n2503 GNDA.n2502 150
R2163 GNDA.n2505 GNDA.n2504 150
R2164 GNDA.n2506 GNDA.n2505 150
R2165 GNDA.n2507 GNDA.n2506 150
R2166 GNDA.n2508 GNDA.n2507 150
R2167 GNDA.n2493 GNDA.n2456 150
R2168 GNDA.n2457 GNDA.n2456 150
R2169 GNDA.n2458 GNDA.n2457 150
R2170 GNDA.n2459 GNDA.n2458 150
R2171 GNDA.n2461 GNDA.n2460 150
R2172 GNDA.n2462 GNDA.n2461 150
R2173 GNDA.n2463 GNDA.n2462 150
R2174 GNDA.n2464 GNDA.n2463 150
R2175 GNDA.t76 GNDA.t239 149.661
R2176 GNDA.t159 GNDA.t5 149.661
R2177 GNDA.t245 GNDA.t71 149.661
R2178 GNDA.t224 GNDA.t30 149.661
R2179 GNDA.t126 GNDA.t15 149.661
R2180 GNDA.t11 GNDA.t233 149.661
R2181 GNDA.t93 GNDA.t341 147.84
R2182 GNDA.t4 GNDA.t64 144.321
R2183 GNDA.n859 GNDA.n858 139.077
R2184 GNDA.n861 GNDA.n860 139.077
R2185 GNDA.n863 GNDA.n862 139.077
R2186 GNDA.n865 GNDA.n864 139.077
R2187 GNDA.n1019 GNDA.n1018 139.077
R2188 GNDA.n1021 GNDA.n1020 139.077
R2189 GNDA.n1023 GNDA.n1022 139.077
R2190 GNDA.n1027 GNDA.n1026 139.077
R2191 GNDA.n1025 GNDA.n1024 139.077
R2192 GNDA.n126 GNDA.n125 139.077
R2193 GNDA.t317 GNDA.t32 139.041
R2194 GNDA.n1965 GNDA.t352 135.69
R2195 GNDA.n162 GNDA.n161 134.268
R2196 GNDA.n168 GNDA.n161 134.268
R2197 GNDA.n1260 GNDA.n1259 132.721
R2198 GNDA.n1970 GNDA.t270 130.001
R2199 GNDA.n1030 GNDA.t279 130.001
R2200 GNDA.n1035 GNDA.t256 130.001
R2201 GNDA.n1157 GNDA.t308 130.001
R2202 GNDA.n1162 GNDA.t283 130.001
R2203 GNDA.n856 GNDA.t276 130.001
R2204 GNDA.n1041 GNDA.n111 124.832
R2205 GNDA.n1039 GNDA.n1038 124.832
R2206 GNDA.n1154 GNDA.n1153 124.832
R2207 GNDA.n478 GNDA.n477 124.832
R2208 GNDA.n1147 GNDA.n1146 124.832
R2209 GNDA.n509 GNDA.n505 124.832
R2210 GNDA.n1703 GNDA.n1702 124.832
R2211 GNDA.n1707 GNDA.n1705 124.832
R2212 GNDA.n1696 GNDA.n510 124.832
R2213 GNDA.n1783 GNDA.n1782 124.832
R2214 GNDA.n1732 GNDA.n441 124.832
R2215 GNDA.n1780 GNDA.n1779 124.832
R2216 GNDA.n2429 GNDA.n2428 117.394
R2217 GNDA.n71 GNDA.t33 115.948
R2218 GNDA.n209 GNDA.t68 115.105
R2219 GNDA.n71 GNDA.t65 114.635
R2220 GNDA.n210 GNDA.t342 114.635
R2221 GNDA.n2397 GNDA.t292 103.665
R2222 GNDA.t298 GNDA.n18 103.665
R2223 GNDA.n1037 GNDA.t255 101.942
R2224 GNDA.n2060 GNDA.n77 101.718
R2225 GNDA.n2446 GNDA.n32 101.718
R2226 GNDA.n2542 GNDA.n19 101.718
R2227 GNDA.n2403 GNDA.n2218 101.718
R2228 GNDA.n2419 GNDA.n2112 101.718
R2229 GNDA.n2490 GNDA.n26 101.718
R2230 GNDA.n2487 GNDA.n27 101.718
R2231 GNDA.n2483 GNDA.n28 101.718
R2232 GNDA.n2479 GNDA.n29 101.718
R2233 GNDA.n2475 GNDA.n30 101.718
R2234 GNDA.n2530 GNDA.n20 101.718
R2235 GNDA.n2527 GNDA.n21 101.718
R2236 GNDA.n2523 GNDA.n22 101.718
R2237 GNDA.n2519 GNDA.n23 101.718
R2238 GNDA.n2515 GNDA.n24 101.718
R2239 GNDA.n2211 GNDA.n2122 101.718
R2240 GNDA.n2208 GNDA.n2123 101.718
R2241 GNDA.n2204 GNDA.n2124 101.718
R2242 GNDA.n2200 GNDA.n2125 101.718
R2243 GNDA.n2196 GNDA.n2126 101.718
R2244 GNDA.n2283 GNDA.n2259 101.718
R2245 GNDA.n2320 GNDA.n2309 101.718
R2246 GNDA.n2160 GNDA.n2159 101.718
R2247 GNDA.n2163 GNDA.n2162 101.718
R2248 GNDA.n2170 GNDA.n2169 101.718
R2249 GNDA.n2173 GNDA.n2172 101.718
R2250 GNDA.n2180 GNDA.n2179 101.718
R2251 GNDA.n2153 GNDA.n2152 101.718
R2252 GNDA.n2161 GNDA.n2160 101.718
R2253 GNDA.n2162 GNDA.n2146 101.718
R2254 GNDA.n2171 GNDA.n2170 101.718
R2255 GNDA.n2172 GNDA.n2142 101.718
R2256 GNDA.n2181 GNDA.n2180 101.718
R2257 GNDA.n2318 GNDA.n2311 101.718
R2258 GNDA.n2281 GNDA.n2274 101.718
R2259 GNDA.n2216 GNDA.n2129 101.718
R2260 GNDA.n2209 GNDA.n2122 101.718
R2261 GNDA.n2205 GNDA.n2123 101.718
R2262 GNDA.n2201 GNDA.n2124 101.718
R2263 GNDA.n2197 GNDA.n2125 101.718
R2264 GNDA.n2193 GNDA.n2126 101.718
R2265 GNDA.n2535 GNDA.n2498 101.718
R2266 GNDA.n2528 GNDA.n20 101.718
R2267 GNDA.n2524 GNDA.n21 101.718
R2268 GNDA.n2520 GNDA.n22 101.718
R2269 GNDA.n2516 GNDA.n23 101.718
R2270 GNDA.n2512 GNDA.n24 101.718
R2271 GNDA.n2495 GNDA.n2454 101.718
R2272 GNDA.n2488 GNDA.n26 101.718
R2273 GNDA.n2484 GNDA.n27 101.718
R2274 GNDA.n2480 GNDA.n28 101.718
R2275 GNDA.n2476 GNDA.n29 101.718
R2276 GNDA.n2472 GNDA.n30 101.718
R2277 GNDA.n2424 GNDA.n2116 101.718
R2278 GNDA.n2417 GNDA.n2112 101.718
R2279 GNDA.n2396 GNDA.n2220 101.718
R2280 GNDA.n2383 GNDA.n2234 101.718
R2281 GNDA.n2271 GNDA.n2261 101.718
R2282 GNDA.n2227 GNDA.n2226 101.718
R2283 GNDA.n2408 GNDA.n2399 101.718
R2284 GNDA.n2218 GNDA.n2121 101.718
R2285 GNDA.n2547 GNDA.n2538 101.718
R2286 GNDA.n19 GNDA.n17 101.718
R2287 GNDA.n2451 GNDA.n2439 101.718
R2288 GNDA.n2444 GNDA.n32 101.718
R2289 GNDA.n2333 GNDA.n2245 101.718
R2290 GNDA.n2343 GNDA.n2336 101.718
R2291 GNDA.n2376 GNDA.n2239 101.718
R2292 GNDA.n2365 GNDA.n2243 101.718
R2293 GNDA.n2071 GNDA.n76 101.718
R2294 GNDA.n172 GNDA.n159 101.718
R2295 GNDA.n164 GNDA.n160 101.718
R2296 GNDA.n163 GNDA.n159 101.718
R2297 GNDA.t221 GNDA.n180 47.6748
R2298 GNDA.t221 GNDA.n177 47.6748
R2299 GNDA.n2307 GNDA.n2306 99.0842
R2300 GNDA.n2305 GNDA.n2304 99.0842
R2301 GNDA.n2303 GNDA.n2302 99.0842
R2302 GNDA.n2301 GNDA.n2300 99.0842
R2303 GNDA.n2299 GNDA.n2298 99.0842
R2304 GNDA.n2297 GNDA.n2296 99.0842
R2305 GNDA.n2295 GNDA.n2294 99.0842
R2306 GNDA.n2293 GNDA.n2292 99.0842
R2307 GNDA.n2291 GNDA.n2290 99.0842
R2308 GNDA.n2289 GNDA.n2288 99.0842
R2309 GNDA.n2287 GNDA.n2286 99.0842
R2310 GNDA.n1937 GNDA.t221 98.9756
R2311 GNDA.n1155 GNDA.n866 98.8538
R2312 GNDA.n2186 GNDA.n2185 94.601
R2313 GNDA.n2188 GNDA.n2187 94.601
R2314 GNDA.n2466 GNDA.n2465 94.601
R2315 GNDA.n2468 GNDA.n2467 94.601
R2316 GNDA.n2035 GNDA.n2034 92.6754
R2317 GNDA.t104 GNDA.t339 92.1471
R2318 GNDA.t339 GNDA.t119 92.1471
R2319 GNDA.t119 GNDA.t120 92.1471
R2320 GNDA.t328 GNDA.t343 92.1471
R2321 GNDA.n2067 GNDA.n75 91.069
R2322 GNDA.n2062 GNDA.n75 91.069
R2323 GNDA.n2064 GNDA.n74 91.069
R2324 GNDA.n2065 GNDA.n2064 91.069
R2325 GNDA.n2381 GNDA.n2233 91.069
R2326 GNDA.n2380 GNDA.n2232 91.069
R2327 GNDA.n2269 GNDA.n2268 91.069
R2328 GNDA.n2264 GNDA.n2262 91.069
R2329 GNDA.n166 GNDA.n162 91.069
R2330 GNDA.n169 GNDA.n168 91.069
R2331 GNDA.t282 GNDA.n1164 90.616
R2332 GNDA.n2393 GNDA.n2221 90.4158
R2333 GNDA.n2315 GNDA.n2312 90.2704
R2334 GNDA.n2312 GNDA.n2308 90.2704
R2335 GNDA.n2278 GNDA.n2275 90.2704
R2336 GNDA.n2275 GNDA.n2258 90.2704
R2337 GNDA.n2224 GNDA.n2222 90.2704
R2338 GNDA.n2330 GNDA.n2246 90.2704
R2339 GNDA.n2340 GNDA.n2337 90.2704
R2340 GNDA.n2373 GNDA.n2240 90.2704
R2341 GNDA.n2362 GNDA.n2242 90.2704
R2342 GNDA.n1643 GNDA.t44 89.6052
R2343 GNDA.n1936 GNDA.n181 88.5317
R2344 GNDA.n1930 GNDA.n181 88.5317
R2345 GNDA.n1930 GNDA.n1929 88.5317
R2346 GNDA.n1929 GNDA.n1928 88.5317
R2347 GNDA.n1928 GNDA.n187 88.5317
R2348 GNDA.n1922 GNDA.n1921 88.5317
R2349 GNDA.n1921 GNDA.n1920 88.5317
R2350 GNDA.n1920 GNDA.n191 88.5317
R2351 GNDA.n1914 GNDA.n191 88.5317
R2352 GNDA.n1914 GNDA.n144 88.5317
R2353 GNDA.n202 GNDA.n143 88.5317
R2354 GNDA.n1900 GNDA.n202 88.5317
R2355 GNDA.n1900 GNDA.n1899 88.5317
R2356 GNDA.n1899 GNDA.n1898 88.5317
R2357 GNDA.n1898 GNDA.n203 88.5317
R2358 GNDA.n1891 GNDA.n1890 88.5317
R2359 GNDA.n1890 GNDA.n1889 88.5317
R2360 GNDA.n1889 GNDA.n215 88.5317
R2361 GNDA.n1883 GNDA.n215 88.5317
R2362 GNDA.n1883 GNDA.n1882 88.5317
R2363 GNDA.n1880 GNDA.n220 88.5317
R2364 GNDA.n1874 GNDA.n220 88.5317
R2365 GNDA.n1874 GNDA.n1873 88.5317
R2366 GNDA.n1873 GNDA.n1872 88.5317
R2367 GNDA.n1872 GNDA.n226 88.5317
R2368 GNDA.n1866 GNDA.n1865 88.5317
R2369 GNDA.n1865 GNDA.n1864 88.5317
R2370 GNDA.n1864 GNDA.n230 88.5317
R2371 GNDA.n1858 GNDA.n230 88.5317
R2372 GNDA.n1858 GNDA.n1857 88.5317
R2373 GNDA.t343 GNDA.n2425 88.3077
R2374 GNDA.t315 GNDA.n108 85.4674
R2375 GNDA.t133 GNDA.t90 84.4682
R2376 GNDA.t57 GNDA.t332 84.4682
R2377 GNDA.t61 GNDA.t38 84.4682
R2378 GNDA.t85 GNDA.t27 84.4682
R2379 GNDA.t145 GNDA.t26 84.4682
R2380 GNDA.t348 GNDA.t292 84.4682
R2381 GNDA.t162 GNDA.t348 84.4682
R2382 GNDA.t149 GNDA.t162 84.4682
R2383 GNDA.t28 GNDA.t355 84.4682
R2384 GNDA.t21 GNDA.t346 84.4682
R2385 GNDA.t346 GNDA.t298 84.4682
R2386 GNDA.t138 GNDA.t106 84.4682
R2387 GNDA.t116 GNDA.t350 84.4682
R2388 GNDA.t2 GNDA.t334 84.4682
R2389 GNDA.t55 GNDA.t114 84.4682
R2390 GNDA.t54 GNDA.t92 84.4682
R2391 GNDA.n2088 GNDA.t195 84.4377
R2392 GNDA.n213 GNDA.n208 84.306
R2393 GNDA.t60 GNDA.t154 82.3782
R2394 GNDA.t351 GNDA.t66 82.3782
R2395 GNDA.n1881 GNDA.n219 80.9821
R2396 GNDA.t295 GNDA.t248 80.6288
R2397 GNDA.t258 GNDA.t272 80.6288
R2398 GNDA.t218 GNDA.t261 80.6288
R2399 GNDA.t251 GNDA.t236 80.6288
R2400 GNDA.n1003 GNDA.t185 80.3188
R2401 GNDA.t165 GNDA.t304 76.7893
R2402 GNDA.t7 GNDA.t146 76.7893
R2403 GNDA.t266 GNDA.t83 76.7893
R2404 GNDA.n1086 GNDA.n1085 76.3222
R2405 GNDA.n1081 GNDA.n1063 76.3222
R2406 GNDA.n1079 GNDA.n1078 76.3222
R2407 GNDA.n1074 GNDA.n1066 76.3222
R2408 GNDA.n1072 GNDA.n1071 76.3222
R2409 GNDA.n1067 GNDA.n141 76.3222
R2410 GNDA.n1089 GNDA.n1088 76.3222
R2411 GNDA.n1059 GNDA.n1058 76.3222
R2412 GNDA.n1052 GNDA.n924 76.3222
R2413 GNDA.n1051 GNDA.n1050 76.3222
R2414 GNDA.n1044 GNDA.n931 76.3222
R2415 GNDA.n1043 GNDA.n1042 76.3222
R2416 GNDA.n1093 GNDA.n1092 76.3222
R2417 GNDA.n926 GNDA.n925 76.3222
R2418 GNDA.n929 GNDA.n928 76.3222
R2419 GNDA.n934 GNDA.n933 76.3222
R2420 GNDA.n937 GNDA.n936 76.3222
R2421 GNDA.n1039 GNDA.n940 76.3222
R2422 GNDA.n1114 GNDA.n1113 76.3222
R2423 GNDA.n1109 GNDA.n913 76.3222
R2424 GNDA.n1107 GNDA.n1106 76.3222
R2425 GNDA.n1102 GNDA.n916 76.3222
R2426 GNDA.n1100 GNDA.n1099 76.3222
R2427 GNDA.n1095 GNDA.n919 76.3222
R2428 GNDA.n1117 GNDA.n1116 76.3222
R2429 GNDA.n1126 GNDA.n1125 76.3222
R2430 GNDA.n1129 GNDA.n1128 76.3222
R2431 GNDA.n1138 GNDA.n1137 76.3222
R2432 GNDA.n1141 GNDA.n1140 76.3222
R2433 GNDA.n1152 GNDA.n1151 76.3222
R2434 GNDA.n1911 GNDA.n1910 76.3222
R2435 GNDA.n453 GNDA.n452 76.3222
R2436 GNDA.n454 GNDA.n447 76.3222
R2437 GNDA.n465 GNDA.n464 76.3222
R2438 GNDA.n467 GNDA.n466 76.3222
R2439 GNDA.n477 GNDA.n442 76.3222
R2440 GNDA.n732 GNDA.n611 76.3222
R2441 GNDA.n727 GNDA.n614 76.3222
R2442 GNDA.n644 GNDA.n643 76.3222
R2443 GNDA.n647 GNDA.n646 76.3222
R2444 GNDA.n660 GNDA.n659 76.3222
R2445 GNDA.n665 GNDA.n664 76.3222
R2446 GNDA.n584 GNDA.n182 76.3222
R2447 GNDA.n593 GNDA.n585 76.3222
R2448 GNDA.n597 GNDA.n586 76.3222
R2449 GNDA.n601 GNDA.n587 76.3222
R2450 GNDA.n605 GNDA.n588 76.3222
R2451 GNDA.n1121 GNDA.n1120 76.3222
R2452 GNDA.n1122 GNDA.n877 76.3222
R2453 GNDA.n1133 GNDA.n1132 76.3222
R2454 GNDA.n1134 GNDA.n873 76.3222
R2455 GNDA.n1145 GNDA.n1144 76.3222
R2456 GNDA.n1148 GNDA.n1147 76.3222
R2457 GNDA.n888 GNDA.n887 76.3222
R2458 GNDA.n889 GNDA.n885 76.3222
R2459 GNDA.n896 GNDA.n895 76.3222
R2460 GNDA.n897 GNDA.n883 76.3222
R2461 GNDA.n904 GNDA.n903 76.3222
R2462 GNDA.n905 GNDA.n881 76.3222
R2463 GNDA.n1257 GNDA.n1256 76.3222
R2464 GNDA.n1252 GNDA.n794 76.3222
R2465 GNDA.n1249 GNDA.n793 76.3222
R2466 GNDA.n1245 GNDA.n792 76.3222
R2467 GNDA.n1241 GNDA.n791 76.3222
R2468 GNDA.n1257 GNDA.n795 76.3222
R2469 GNDA.n1250 GNDA.n794 76.3222
R2470 GNDA.n1246 GNDA.n793 76.3222
R2471 GNDA.n1242 GNDA.n792 76.3222
R2472 GNDA.n1238 GNDA.n791 76.3222
R2473 GNDA.n592 GNDA.n584 76.3222
R2474 GNDA.n596 GNDA.n585 76.3222
R2475 GNDA.n600 GNDA.n586 76.3222
R2476 GNDA.n604 GNDA.n587 76.3222
R2477 GNDA.n607 GNDA.n588 76.3222
R2478 GNDA.n486 GNDA.n485 76.3222
R2479 GNDA.n489 GNDA.n488 76.3222
R2480 GNDA.n494 GNDA.n493 76.3222
R2481 GNDA.n497 GNDA.n496 76.3222
R2482 GNDA.n502 GNDA.n501 76.3222
R2483 GNDA.n505 GNDA.n504 76.3222
R2484 GNDA.n767 GNDA.n766 76.3222
R2485 GNDA.n762 GNDA.n743 76.3222
R2486 GNDA.n760 GNDA.n759 76.3222
R2487 GNDA.n755 GNDA.n746 76.3222
R2488 GNDA.n753 GNDA.n752 76.3222
R2489 GNDA.n748 GNDA.n747 76.3222
R2490 GNDA.n1377 GNDA.n1376 76.3222
R2491 GNDA.n1263 GNDA.n579 76.3222
R2492 GNDA.n1366 GNDA.n578 76.3222
R2493 GNDA.n1293 GNDA.n577 76.3222
R2494 GNDA.n1297 GNDA.n576 76.3222
R2495 GNDA.n1306 GNDA.n575 76.3222
R2496 GNDA.n769 GNDA.n735 76.3222
R2497 GNDA.n773 GNDA.n736 76.3222
R2498 GNDA.n777 GNDA.n737 76.3222
R2499 GNDA.n781 GNDA.n738 76.3222
R2500 GNDA.n788 GNDA.n739 76.3222
R2501 GNDA.n1259 GNDA.n583 76.3222
R2502 GNDA.n772 GNDA.n735 76.3222
R2503 GNDA.n776 GNDA.n736 76.3222
R2504 GNDA.n780 GNDA.n737 76.3222
R2505 GNDA.n783 GNDA.n738 76.3222
R2506 GNDA.n788 GNDA.n787 76.3222
R2507 GNDA.n1664 GNDA.n1663 76.3222
R2508 GNDA.n1659 GNDA.n556 76.3222
R2509 GNDA.n1657 GNDA.n1656 76.3222
R2510 GNDA.n1652 GNDA.n559 76.3222
R2511 GNDA.n1650 GNDA.n1649 76.3222
R2512 GNDA.n1645 GNDA.n562 76.3222
R2513 GNDA.n1391 GNDA.n512 76.3222
R2514 GNDA.n1589 GNDA.n1588 76.3222
R2515 GNDA.n1592 GNDA.n1591 76.3222
R2516 GNDA.n1604 GNDA.n1603 76.3222
R2517 GNDA.n1607 GNDA.n1606 76.3222
R2518 GNDA.n1619 GNDA.n1618 76.3222
R2519 GNDA.n1667 GNDA.n1666 76.3222
R2520 GNDA.n1676 GNDA.n1675 76.3222
R2521 GNDA.n1679 GNDA.n1678 76.3222
R2522 GNDA.n1688 GNDA.n1687 76.3222
R2523 GNDA.n1691 GNDA.n1690 76.3222
R2524 GNDA.n1701 GNDA.n1700 76.3222
R2525 GNDA.n1728 GNDA.n1727 76.3222
R2526 GNDA.n1725 GNDA.n484 76.3222
R2527 GNDA.n1721 GNDA.n1720 76.3222
R2528 GNDA.n1714 GNDA.n491 76.3222
R2529 GNDA.n1713 GNDA.n1712 76.3222
R2530 GNDA.n1706 GNDA.n499 76.3222
R2531 GNDA.n531 GNDA.n530 76.3222
R2532 GNDA.n532 GNDA.n528 76.3222
R2533 GNDA.n539 GNDA.n538 76.3222
R2534 GNDA.n540 GNDA.n526 76.3222
R2535 GNDA.n547 GNDA.n546 76.3222
R2536 GNDA.n548 GNDA.n524 76.3222
R2537 GNDA.n1467 GNDA.n507 76.3222
R2538 GNDA.n1546 GNDA.n1545 76.3222
R2539 GNDA.n1549 GNDA.n1548 76.3222
R2540 GNDA.n1561 GNDA.n1560 76.3222
R2541 GNDA.n1564 GNDA.n1563 76.3222
R2542 GNDA.n1573 GNDA.n1572 76.3222
R2543 GNDA.n1671 GNDA.n1670 76.3222
R2544 GNDA.n1672 GNDA.n520 76.3222
R2545 GNDA.n1683 GNDA.n1682 76.3222
R2546 GNDA.n1684 GNDA.n516 76.3222
R2547 GNDA.n1695 GNDA.n1694 76.3222
R2548 GNDA.n1697 GNDA.n1696 76.3222
R2549 GNDA.n1785 GNDA.n1784 76.3222
R2550 GNDA.n1798 GNDA.n1797 76.3222
R2551 GNDA.n1801 GNDA.n1800 76.3222
R2552 GNDA.n1813 GNDA.n1812 76.3222
R2553 GNDA.n1816 GNDA.n1815 76.3222
R2554 GNDA.n1828 GNDA.n1827 76.3222
R2555 GNDA.n1907 GNDA.n1906 76.3222
R2556 GNDA.n449 GNDA.n197 76.3222
R2557 GNDA.n458 GNDA.n457 76.3222
R2558 GNDA.n461 GNDA.n460 76.3222
R2559 GNDA.n471 GNDA.n470 76.3222
R2560 GNDA.n474 GNDA.n473 76.3222
R2561 GNDA.n1734 GNDA.n1733 76.3222
R2562 GNDA.n1747 GNDA.n1746 76.3222
R2563 GNDA.n1750 GNDA.n1749 76.3222
R2564 GNDA.n1762 GNDA.n1761 76.3222
R2565 GNDA.n1765 GNDA.n1764 76.3222
R2566 GNDA.n1777 GNDA.n1776 76.3222
R2567 GNDA.n1698 GNDA.n1697 76.3222
R2568 GNDA.n1694 GNDA.n1693 76.3222
R2569 GNDA.n1685 GNDA.n1684 76.3222
R2570 GNDA.n1682 GNDA.n1681 76.3222
R2571 GNDA.n1673 GNDA.n1672 76.3222
R2572 GNDA.n1670 GNDA.n1669 76.3222
R2573 GNDA.n1666 GNDA.n522 76.3222
R2574 GNDA.n1677 GNDA.n1676 76.3222
R2575 GNDA.n1678 GNDA.n518 76.3222
R2576 GNDA.n1689 GNDA.n1688 76.3222
R2577 GNDA.n1690 GNDA.n514 76.3222
R2578 GNDA.n1702 GNDA.n1701 76.3222
R2579 GNDA.n749 GNDA.n748 76.3222
R2580 GNDA.n754 GNDA.n753 76.3222
R2581 GNDA.n746 GNDA.n744 76.3222
R2582 GNDA.n761 GNDA.n760 76.3222
R2583 GNDA.n743 GNDA.n741 76.3222
R2584 GNDA.n768 GNDA.n767 76.3222
R2585 GNDA.n549 GNDA.n548 76.3222
R2586 GNDA.n546 GNDA.n545 76.3222
R2587 GNDA.n541 GNDA.n540 76.3222
R2588 GNDA.n538 GNDA.n537 76.3222
R2589 GNDA.n533 GNDA.n532 76.3222
R2590 GNDA.n530 GNDA.n483 76.3222
R2591 GNDA.n562 GNDA.n560 76.3222
R2592 GNDA.n1651 GNDA.n1650 76.3222
R2593 GNDA.n559 GNDA.n557 76.3222
R2594 GNDA.n1658 GNDA.n1657 76.3222
R2595 GNDA.n556 GNDA.n554 76.3222
R2596 GNDA.n1665 GNDA.n1664 76.3222
R2597 GNDA.n728 GNDA.n611 76.3222
R2598 GNDA.n638 GNDA.n614 76.3222
R2599 GNDA.n645 GNDA.n644 76.3222
R2600 GNDA.n646 GNDA.n636 76.3222
R2601 GNDA.n661 GNDA.n660 76.3222
R2602 GNDA.n664 GNDA.n663 76.3222
R2603 GNDA.n1733 GNDA.n377 76.3222
R2604 GNDA.n1748 GNDA.n1747 76.3222
R2605 GNDA.n1749 GNDA.n372 76.3222
R2606 GNDA.n1763 GNDA.n1762 76.3222
R2607 GNDA.n1764 GNDA.n365 76.3222
R2608 GNDA.n1778 GNDA.n1777 76.3222
R2609 GNDA.n1784 GNDA.n258 76.3222
R2610 GNDA.n1799 GNDA.n1798 76.3222
R2611 GNDA.n1800 GNDA.n253 76.3222
R2612 GNDA.n1814 GNDA.n1813 76.3222
R2613 GNDA.n1815 GNDA.n246 76.3222
R2614 GNDA.n1829 GNDA.n1828 76.3222
R2615 GNDA.n444 GNDA.n442 76.3222
R2616 GNDA.n468 GNDA.n467 76.3222
R2617 GNDA.n464 GNDA.n463 76.3222
R2618 GNDA.n455 GNDA.n454 76.3222
R2619 GNDA.n452 GNDA.n195 76.3222
R2620 GNDA.n1912 GNDA.n1911 76.3222
R2621 GNDA.n1908 GNDA.n1907 76.3222
R2622 GNDA.n450 GNDA.n449 76.3222
R2623 GNDA.n459 GNDA.n458 76.3222
R2624 GNDA.n460 GNDA.n445 76.3222
R2625 GNDA.n472 GNDA.n471 76.3222
R2626 GNDA.n473 GNDA.n441 76.3222
R2627 GNDA.n504 GNDA.n503 76.3222
R2628 GNDA.n501 GNDA.n500 76.3222
R2629 GNDA.n496 GNDA.n495 76.3222
R2630 GNDA.n493 GNDA.n492 76.3222
R2631 GNDA.n488 GNDA.n487 76.3222
R2632 GNDA.n485 GNDA.n481 76.3222
R2633 GNDA.n1727 GNDA.n1726 76.3222
R2634 GNDA.n1722 GNDA.n484 76.3222
R2635 GNDA.n1720 GNDA.n1719 76.3222
R2636 GNDA.n1715 GNDA.n1714 76.3222
R2637 GNDA.n1712 GNDA.n1711 76.3222
R2638 GNDA.n1707 GNDA.n1706 76.3222
R2639 GNDA.n1149 GNDA.n1148 76.3222
R2640 GNDA.n1144 GNDA.n1143 76.3222
R2641 GNDA.n1135 GNDA.n1134 76.3222
R2642 GNDA.n1132 GNDA.n1131 76.3222
R2643 GNDA.n1123 GNDA.n1122 76.3222
R2644 GNDA.n1120 GNDA.n1119 76.3222
R2645 GNDA.n1116 GNDA.n879 76.3222
R2646 GNDA.n1127 GNDA.n1126 76.3222
R2647 GNDA.n1128 GNDA.n875 76.3222
R2648 GNDA.n1139 GNDA.n1138 76.3222
R2649 GNDA.n1140 GNDA.n871 76.3222
R2650 GNDA.n1153 GNDA.n1152 76.3222
R2651 GNDA.n940 GNDA.n939 76.3222
R2652 GNDA.n936 GNDA.n935 76.3222
R2653 GNDA.n933 GNDA.n932 76.3222
R2654 GNDA.n928 GNDA.n927 76.3222
R2655 GNDA.n925 GNDA.n922 76.3222
R2656 GNDA.n1094 GNDA.n1093 76.3222
R2657 GNDA.n1090 GNDA.n1089 76.3222
R2658 GNDA.n1058 GNDA.n1057 76.3222
R2659 GNDA.n1053 GNDA.n1052 76.3222
R2660 GNDA.n1050 GNDA.n1049 76.3222
R2661 GNDA.n1045 GNDA.n1044 76.3222
R2662 GNDA.n1042 GNDA.n1041 76.3222
R2663 GNDA.n906 GNDA.n905 76.3222
R2664 GNDA.n903 GNDA.n902 76.3222
R2665 GNDA.n898 GNDA.n897 76.3222
R2666 GNDA.n895 GNDA.n894 76.3222
R2667 GNDA.n890 GNDA.n889 76.3222
R2668 GNDA.n887 GNDA.n796 76.3222
R2669 GNDA.n919 GNDA.n917 76.3222
R2670 GNDA.n1101 GNDA.n1100 76.3222
R2671 GNDA.n916 GNDA.n914 76.3222
R2672 GNDA.n1108 GNDA.n1107 76.3222
R2673 GNDA.n913 GNDA.n911 76.3222
R2674 GNDA.n1115 GNDA.n1114 76.3222
R2675 GNDA.n1068 GNDA.n1067 76.3222
R2676 GNDA.n1073 GNDA.n1072 76.3222
R2677 GNDA.n1066 GNDA.n1064 76.3222
R2678 GNDA.n1080 GNDA.n1079 76.3222
R2679 GNDA.n1063 GNDA.n1061 76.3222
R2680 GNDA.n1087 GNDA.n1086 76.3222
R2681 GNDA.n1377 GNDA.n580 76.3222
R2682 GNDA.n1367 GNDA.n579 76.3222
R2683 GNDA.n1292 GNDA.n578 76.3222
R2684 GNDA.n1298 GNDA.n577 76.3222
R2685 GNDA.n1305 GNDA.n576 76.3222
R2686 GNDA.n1287 GNDA.n575 76.3222
R2687 GNDA.n1468 GNDA.n1467 76.3222
R2688 GNDA.n1547 GNDA.n1546 76.3222
R2689 GNDA.n1548 GNDA.n1462 76.3222
R2690 GNDA.n1562 GNDA.n1561 76.3222
R2691 GNDA.n1563 GNDA.n1456 76.3222
R2692 GNDA.n1574 GNDA.n1573 76.3222
R2693 GNDA.n1392 GNDA.n1391 76.3222
R2694 GNDA.n1590 GNDA.n1589 76.3222
R2695 GNDA.n1591 GNDA.n1386 76.3222
R2696 GNDA.n1605 GNDA.n1604 76.3222
R2697 GNDA.n1606 GNDA.n1379 76.3222
R2698 GNDA.n1620 GNDA.n1619 76.3222
R2699 GNDA.t296 GNDA.n2166 75.0005
R2700 GNDA.n2167 GNDA.t296 75.0005
R2701 GNDA.t273 GNDA.n2134 75.0005
R2702 GNDA.n2135 GNDA.t273 75.0005
R2703 GNDA.n2406 GNDA.t259 75.0005
R2704 GNDA.n2401 GNDA.t259 75.0005
R2705 GNDA.n2422 GNDA.t249 75.0005
R2706 GNDA.n2118 GNDA.t249 75.0005
R2707 GNDA.n2545 GNDA.t219 75.0005
R2708 GNDA.n2540 GNDA.t219 75.0005
R2709 GNDA.n2449 GNDA.t237 75.0005
R2710 GNDA.n2441 GNDA.t237 75.0005
R2711 GNDA.t262 GNDA.n2503 75.0005
R2712 GNDA.n2504 GNDA.t262 75.0005
R2713 GNDA.t252 GNDA.n2459 75.0005
R2714 GNDA.n2460 GNDA.t252 75.0005
R2715 GNDA.n2345 GNDA.t157 74.8304
R2716 GNDA.n2344 GNDA.t17 74.8304
R2717 GNDA.t127 GNDA.n2377 74.8304
R2718 GNDA.t129 GNDA.n2361 74.8304
R2719 GNDA.n688 GNDA.n623 74.5978
R2720 GNDA.n685 GNDA.n623 74.5978
R2721 GNDA.n1189 GNDA.n811 74.5978
R2722 GNDA.n1186 GNDA.n811 74.5978
R2723 GNDA.n1329 GNDA.n1275 74.5978
R2724 GNDA.n1326 GNDA.n1275 74.5978
R2725 GNDA.n1498 GNDA.n1478 74.5978
R2726 GNDA.n1499 GNDA.n1498 74.5978
R2727 GNDA.n1419 GNDA.n1402 74.5978
R2728 GNDA.n1420 GNDA.n1419 74.5978
R2729 GNDA.n404 GNDA.n387 74.5978
R2730 GNDA.n405 GNDA.n404 74.5978
R2731 GNDA.n285 GNDA.n268 74.5978
R2732 GNDA.n286 GNDA.n285 74.5978
R2733 GNDA.n979 GNDA.n52 74.5978
R2734 GNDA.n982 GNDA.n52 74.5978
R2735 GNDA.n1997 GNDA.n91 74.5978
R2736 GNDA.n1994 GNDA.n91 74.5978
R2737 GNDA.n1006 GNDA.t201 74.1404
R2738 GNDA.t143 GNDA.n2272 72.9499
R2739 GNDA.n2282 GNDA.t12 72.9499
R2740 GNDA.n2090 GNDA.t197 70.0216
R2741 GNDA.n722 GNDA.n616 69.3109
R2742 GNDA.n722 GNDA.n721 69.3109
R2743 GNDA.n1225 GNDA.n804 69.3109
R2744 GNDA.n1225 GNDA.n1224 69.3109
R2745 GNDA.n1371 GNDA.n1265 69.3109
R2746 GNDA.n1347 GNDA.n1265 69.3109
R2747 GNDA.n1540 GNDA.n1539 69.3109
R2748 GNDA.n1539 GNDA.n1538 69.3109
R2749 GNDA.n1583 GNDA.n1582 69.3109
R2750 GNDA.n1582 GNDA.n1581 69.3109
R2751 GNDA.n1741 GNDA.n1740 69.3109
R2752 GNDA.n1740 GNDA.n1739 69.3109
R2753 GNDA.n1792 GNDA.n1791 69.3109
R2754 GNDA.n1791 GNDA.n1790 69.3109
R2755 GNDA.n2095 GNDA.n2094 69.3109
R2756 GNDA.n2095 GNDA.n63 69.3109
R2757 GNDA.n2053 GNDA.n2052 69.3109
R2758 GNDA.n2053 GNDA.n102 69.3109
R2759 GNDA.t253 GNDA.n633 65.8183
R2760 GNDA.t253 GNDA.n632 65.8183
R2761 GNDA.t253 GNDA.n631 65.8183
R2762 GNDA.t253 GNDA.n630 65.8183
R2763 GNDA.t253 GNDA.n621 65.8183
R2764 GNDA.t253 GNDA.n628 65.8183
R2765 GNDA.t253 GNDA.n618 65.8183
R2766 GNDA.t253 GNDA.n629 65.8183
R2767 GNDA.t253 GNDA.n627 65.8183
R2768 GNDA.t253 GNDA.n626 65.8183
R2769 GNDA.t253 GNDA.n625 65.8183
R2770 GNDA.t253 GNDA.n624 65.8183
R2771 GNDA.t253 GNDA.n622 65.8183
R2772 GNDA.t253 GNDA.n620 65.8183
R2773 GNDA.t253 GNDA.n619 65.8183
R2774 GNDA.n723 GNDA.t253 65.8183
R2775 GNDA.t263 GNDA.n821 65.8183
R2776 GNDA.t263 GNDA.n820 65.8183
R2777 GNDA.t263 GNDA.n819 65.8183
R2778 GNDA.t263 GNDA.n818 65.8183
R2779 GNDA.t263 GNDA.n809 65.8183
R2780 GNDA.t263 GNDA.n816 65.8183
R2781 GNDA.t263 GNDA.n806 65.8183
R2782 GNDA.t263 GNDA.n817 65.8183
R2783 GNDA.t263 GNDA.n815 65.8183
R2784 GNDA.t263 GNDA.n814 65.8183
R2785 GNDA.t263 GNDA.n813 65.8183
R2786 GNDA.t263 GNDA.n812 65.8183
R2787 GNDA.t263 GNDA.n810 65.8183
R2788 GNDA.t263 GNDA.n808 65.8183
R2789 GNDA.t263 GNDA.n807 65.8183
R2790 GNDA.n1226 GNDA.t263 65.8183
R2791 GNDA.t264 GNDA.n1361 65.8183
R2792 GNDA.t264 GNDA.n1284 65.8183
R2793 GNDA.t264 GNDA.n1283 65.8183
R2794 GNDA.t264 GNDA.n1282 65.8183
R2795 GNDA.t264 GNDA.n1273 65.8183
R2796 GNDA.t264 GNDA.n1280 65.8183
R2797 GNDA.t264 GNDA.n1271 65.8183
R2798 GNDA.t264 GNDA.n1281 65.8183
R2799 GNDA.t264 GNDA.n1279 65.8183
R2800 GNDA.t264 GNDA.n1278 65.8183
R2801 GNDA.t264 GNDA.n1277 65.8183
R2802 GNDA.t264 GNDA.n1276 65.8183
R2803 GNDA.t264 GNDA.n1274 65.8183
R2804 GNDA.t264 GNDA.n1272 65.8183
R2805 GNDA.n1362 GNDA.t264 65.8183
R2806 GNDA.t264 GNDA.n1266 65.8183
R2807 GNDA.n1520 GNDA.t220 65.8183
R2808 GNDA.n1522 GNDA.t220 65.8183
R2809 GNDA.n1528 GNDA.t220 65.8183
R2810 GNDA.n1530 GNDA.t220 65.8183
R2811 GNDA.n1504 GNDA.t220 65.8183
R2812 GNDA.n1506 GNDA.t220 65.8183
R2813 GNDA.n1512 GNDA.t220 65.8183
R2814 GNDA.n1514 GNDA.t220 65.8183
R2815 GNDA.n1483 GNDA.t220 65.8183
R2816 GNDA.n1489 GNDA.t220 65.8183
R2817 GNDA.n1482 GNDA.t220 65.8183
R2818 GNDA.n1496 GNDA.t220 65.8183
R2819 GNDA.n1568 GNDA.t220 65.8183
R2820 GNDA.n1556 GNDA.t220 65.8183
R2821 GNDA.n1554 GNDA.t220 65.8183
R2822 GNDA.n1541 GNDA.t220 65.8183
R2823 GNDA.n1441 GNDA.t280 65.8183
R2824 GNDA.n1443 GNDA.t280 65.8183
R2825 GNDA.n1449 GNDA.t280 65.8183
R2826 GNDA.n1451 GNDA.t280 65.8183
R2827 GNDA.n1425 GNDA.t280 65.8183
R2828 GNDA.n1427 GNDA.t280 65.8183
R2829 GNDA.n1433 GNDA.t280 65.8183
R2830 GNDA.n1435 GNDA.t280 65.8183
R2831 GNDA.t280 GNDA.n1382 65.8183
R2832 GNDA.n1410 GNDA.t280 65.8183
R2833 GNDA.n1406 GNDA.t280 65.8183
R2834 GNDA.n1417 GNDA.t280 65.8183
R2835 GNDA.n1612 GNDA.t280 65.8183
R2836 GNDA.n1599 GNDA.t280 65.8183
R2837 GNDA.n1597 GNDA.t280 65.8183
R2838 GNDA.n1584 GNDA.t280 65.8183
R2839 GNDA.n426 GNDA.t228 65.8183
R2840 GNDA.n428 GNDA.t228 65.8183
R2841 GNDA.n434 GNDA.t228 65.8183
R2842 GNDA.n436 GNDA.t228 65.8183
R2843 GNDA.n410 GNDA.t228 65.8183
R2844 GNDA.n412 GNDA.t228 65.8183
R2845 GNDA.n418 GNDA.t228 65.8183
R2846 GNDA.n420 GNDA.t228 65.8183
R2847 GNDA.t228 GNDA.n368 65.8183
R2848 GNDA.n395 GNDA.t228 65.8183
R2849 GNDA.n391 GNDA.t228 65.8183
R2850 GNDA.n402 GNDA.t228 65.8183
R2851 GNDA.n307 GNDA.t222 65.8183
R2852 GNDA.n309 GNDA.t222 65.8183
R2853 GNDA.n315 GNDA.t222 65.8183
R2854 GNDA.n317 GNDA.t222 65.8183
R2855 GNDA.n291 GNDA.t222 65.8183
R2856 GNDA.n293 GNDA.t222 65.8183
R2857 GNDA.n299 GNDA.t222 65.8183
R2858 GNDA.n301 GNDA.t222 65.8183
R2859 GNDA.t222 GNDA.n249 65.8183
R2860 GNDA.n276 GNDA.t222 65.8183
R2861 GNDA.n272 GNDA.t222 65.8183
R2862 GNDA.n283 GNDA.t222 65.8183
R2863 GNDA.n1821 GNDA.t222 65.8183
R2864 GNDA.n1808 GNDA.t222 65.8183
R2865 GNDA.n1806 GNDA.t222 65.8183
R2866 GNDA.n1793 GNDA.t222 65.8183
R2867 GNDA.n1770 GNDA.t228 65.8183
R2868 GNDA.n1757 GNDA.t228 65.8183
R2869 GNDA.n1755 GNDA.t228 65.8183
R2870 GNDA.n1742 GNDA.t228 65.8183
R2871 GNDA.t226 GNDA.n62 65.8183
R2872 GNDA.t226 GNDA.n61 65.8183
R2873 GNDA.t226 GNDA.n60 65.8183
R2874 GNDA.t226 GNDA.n59 65.8183
R2875 GNDA.t226 GNDA.n50 65.8183
R2876 GNDA.t226 GNDA.n57 65.8183
R2877 GNDA.t226 GNDA.n48 65.8183
R2878 GNDA.t226 GNDA.n58 65.8183
R2879 GNDA.t226 GNDA.n56 65.8183
R2880 GNDA.t226 GNDA.n55 65.8183
R2881 GNDA.t226 GNDA.n54 65.8183
R2882 GNDA.t226 GNDA.n53 65.8183
R2883 GNDA.t226 GNDA.n51 65.8183
R2884 GNDA.n2096 GNDA.t226 65.8183
R2885 GNDA.t226 GNDA.n49 65.8183
R2886 GNDA.t226 GNDA.n47 65.8183
R2887 GNDA.t284 GNDA.n101 65.8183
R2888 GNDA.t284 GNDA.n100 65.8183
R2889 GNDA.t284 GNDA.n99 65.8183
R2890 GNDA.t284 GNDA.n98 65.8183
R2891 GNDA.t284 GNDA.n89 65.8183
R2892 GNDA.t284 GNDA.n96 65.8183
R2893 GNDA.t284 GNDA.n87 65.8183
R2894 GNDA.t284 GNDA.n97 65.8183
R2895 GNDA.t284 GNDA.n95 65.8183
R2896 GNDA.t284 GNDA.n94 65.8183
R2897 GNDA.t284 GNDA.n93 65.8183
R2898 GNDA.t284 GNDA.n92 65.8183
R2899 GNDA.t284 GNDA.n90 65.8183
R2900 GNDA.n2054 GNDA.t284 65.8183
R2901 GNDA.t284 GNDA.n88 65.8183
R2902 GNDA.t284 GNDA.n86 65.8183
R2903 GNDA.t40 GNDA.t133 65.271
R2904 GNDA.t26 GNDA.t42 65.271
R2905 GNDA.t106 GNDA.t109 65.271
R2906 GNDA.t36 GNDA.t54 65.271
R2907 GNDA.t221 GNDA.n178 65.0078
R2908 GNDA.n1231 GNDA.t191 63.8432
R2909 GNDA.n2089 GNDA.t213 63.8432
R2910 GNDA.n2046 GNDA.t207 63.8432
R2911 GNDA.t95 GNDA.t113 62.9326
R2912 GNDA.t63 GNDA.t340 62.9326
R2913 GNDA.t340 GNDA.t3 62.9326
R2914 GNDA.t3 GNDA.t112 62.9326
R2915 GNDA.n2452 GNDA.n2437 61.4316
R2916 GNDA.n850 GNDA.t193 59.7243
R2917 GNDA.n1004 GNDA.t215 59.7243
R2918 GNDA.n124 GNDA.t205 59.7243
R2919 GNDA.n1233 GNDA.t103 58.6946
R2920 GNDA.t89 GNDA.n834 58.6946
R2921 GNDA.t87 GNDA.n851 58.6946
R2922 GNDA.t253 GNDA.n722 57.8461
R2923 GNDA.t263 GNDA.n1225 57.8461
R2924 GNDA.t264 GNDA.n1265 57.8461
R2925 GNDA.n1539 GNDA.t220 57.8461
R2926 GNDA.n1582 GNDA.t280 57.8461
R2927 GNDA.n1791 GNDA.t222 57.8461
R2928 GNDA.n1740 GNDA.t228 57.8461
R2929 GNDA.t226 GNDA.n2095 57.8461
R2930 GNDA.t284 GNDA.n2053 57.8461
R2931 GNDA.t248 GNDA.n2114 57.5921
R2932 GNDA.n2217 GNDA.t258 57.5921
R2933 GNDA.n2319 GNDA.t132 57.5921
R2934 GNDA.n2384 GNDA.t45 57.5921
R2935 GNDA.n2536 GNDA.t218 57.5921
R2936 GNDA.t236 GNDA.n2496 57.5921
R2937 GNDA.t181 GNDA.t321 56.6352
R2938 GNDA.n2076 GNDA.t307 56.6352
R2939 GNDA.t353 GNDA.t177 56.6352
R2940 GNDA.n1960 GNDA.n1959 56.3995
R2941 GNDA.n734 GNDA.n590 56.3995
R2942 GNDA.n798 GNDA.n789 56.3995
R2943 GNDA.n1235 GNDA.n789 56.3995
R2944 GNDA.n734 GNDA.n733 56.3995
R2945 GNDA.n1260 GNDA.n581 56.3995
R2946 GNDA.n1622 GNDA.n573 56.3995
R2947 GNDA.n1834 GNDA.n1833 56.3995
R2948 GNDA.n1961 GNDA.n1960 56.3995
R2949 GNDA.n1622 GNDA.n1621 56.3995
R2950 GNDA.n1834 GNDA.n1830 56.3995
R2951 GNDA.n1163 GNDA.n855 55.6055
R2952 GNDA.t253 GNDA.n623 55.2026
R2953 GNDA.t263 GNDA.n811 55.2026
R2954 GNDA.t264 GNDA.n1275 55.2026
R2955 GNDA.n1498 GNDA.t220 55.2026
R2956 GNDA.n1419 GNDA.t280 55.2026
R2957 GNDA.n404 GNDA.t228 55.2026
R2958 GNDA.n285 GNDA.t222 55.2026
R2959 GNDA.t226 GNDA.n52 55.2026
R2960 GNDA.t284 GNDA.n91 55.2026
R2961 GNDA.n1017 GNDA.n69 54.5757
R2962 GNDA.n1029 GNDA.n1028 54.5757
R2963 GNDA.t25 GNDA.n2047 54.5757
R2964 GNDA.n117 GNDA.t14 54.5757
R2965 GNDA.t67 GNDA.n1972 54.5757
R2966 GNDA.t171 GNDA.t289 53.7527
R2967 GNDA.t336 GNDA.t9 53.7527
R2968 GNDA.t155 GNDA.t62 53.7527
R2969 GNDA.t325 GNDA.t34 53.7527
R2970 GNDA.t147 GNDA.t82 53.7527
R2971 GNDA.t173 GNDA.t140 53.7527
R2972 GNDA.t47 GNDA.t320 53.7527
R2973 GNDA.t310 GNDA.t49 53.7527
R2974 GNDA.t199 GNDA.n1004 53.546
R2975 GNDA.n704 GNDA.n629 53.3664
R2976 GNDA.n700 GNDA.n618 53.3664
R2977 GNDA.n696 GNDA.n628 53.3664
R2978 GNDA.n692 GNDA.n621 53.3664
R2979 GNDA.n681 GNDA.n624 53.3664
R2980 GNDA.n677 GNDA.n625 53.3664
R2981 GNDA.n673 GNDA.n626 53.3664
R2982 GNDA.n669 GNDA.n627 53.3664
R2983 GNDA.n724 GNDA.n723 53.3664
R2984 GNDA.n640 GNDA.n619 53.3664
R2985 GNDA.n651 GNDA.n620 53.3664
R2986 GNDA.n656 GNDA.n622 53.3664
R2987 GNDA.n708 GNDA.n633 53.3664
R2988 GNDA.n709 GNDA.n632 53.3664
R2989 GNDA.n713 GNDA.n631 53.3664
R2990 GNDA.n717 GNDA.n630 53.3664
R2991 GNDA.n705 GNDA.n633 53.3664
R2992 GNDA.n712 GNDA.n632 53.3664
R2993 GNDA.n716 GNDA.n631 53.3664
R2994 GNDA.n720 GNDA.n630 53.3664
R2995 GNDA.n689 GNDA.n621 53.3664
R2996 GNDA.n693 GNDA.n628 53.3664
R2997 GNDA.n697 GNDA.n618 53.3664
R2998 GNDA.n701 GNDA.n629 53.3664
R2999 GNDA.n672 GNDA.n627 53.3664
R3000 GNDA.n676 GNDA.n626 53.3664
R3001 GNDA.n680 GNDA.n625 53.3664
R3002 GNDA.n684 GNDA.n624 53.3664
R3003 GNDA.n668 GNDA.n622 53.3664
R3004 GNDA.n655 GNDA.n620 53.3664
R3005 GNDA.n650 GNDA.n619 53.3664
R3006 GNDA.n723 GNDA.n617 53.3664
R3007 GNDA.n1205 GNDA.n817 53.3664
R3008 GNDA.n1201 GNDA.n806 53.3664
R3009 GNDA.n1197 GNDA.n816 53.3664
R3010 GNDA.n1193 GNDA.n809 53.3664
R3011 GNDA.n1182 GNDA.n812 53.3664
R3012 GNDA.n1178 GNDA.n813 53.3664
R3013 GNDA.n1174 GNDA.n814 53.3664
R3014 GNDA.n1170 GNDA.n815 53.3664
R3015 GNDA.n1227 GNDA.n1226 53.3664
R3016 GNDA.n828 GNDA.n807 53.3664
R3017 GNDA.n841 GNDA.n808 53.3664
R3018 GNDA.n845 GNDA.n810 53.3664
R3019 GNDA.n1209 GNDA.n821 53.3664
R3020 GNDA.n1210 GNDA.n820 53.3664
R3021 GNDA.n1214 GNDA.n819 53.3664
R3022 GNDA.n1218 GNDA.n818 53.3664
R3023 GNDA.n1206 GNDA.n821 53.3664
R3024 GNDA.n1213 GNDA.n820 53.3664
R3025 GNDA.n1217 GNDA.n819 53.3664
R3026 GNDA.n822 GNDA.n818 53.3664
R3027 GNDA.n1190 GNDA.n809 53.3664
R3028 GNDA.n1194 GNDA.n816 53.3664
R3029 GNDA.n1198 GNDA.n806 53.3664
R3030 GNDA.n1202 GNDA.n817 53.3664
R3031 GNDA.n1173 GNDA.n815 53.3664
R3032 GNDA.n1177 GNDA.n814 53.3664
R3033 GNDA.n1181 GNDA.n813 53.3664
R3034 GNDA.n1185 GNDA.n812 53.3664
R3035 GNDA.n1169 GNDA.n810 53.3664
R3036 GNDA.n846 GNDA.n808 53.3664
R3037 GNDA.n840 GNDA.n807 53.3664
R3038 GNDA.n1226 GNDA.n805 53.3664
R3039 GNDA.n1344 GNDA.n1281 53.3664
R3040 GNDA.n1341 GNDA.n1271 53.3664
R3041 GNDA.n1337 GNDA.n1280 53.3664
R3042 GNDA.n1333 GNDA.n1273 53.3664
R3043 GNDA.n1322 GNDA.n1276 53.3664
R3044 GNDA.n1318 GNDA.n1277 53.3664
R3045 GNDA.n1314 GNDA.n1278 53.3664
R3046 GNDA.n1310 GNDA.n1279 53.3664
R3047 GNDA.n1370 GNDA.n1266 53.3664
R3048 GNDA.n1363 GNDA.n1362 53.3664
R3049 GNDA.n1295 GNDA.n1272 53.3664
R3050 GNDA.n1302 GNDA.n1274 53.3664
R3051 GNDA.n1361 GNDA.n1360 53.3664
R3052 GNDA.n1286 GNDA.n1284 53.3664
R3053 GNDA.n1355 GNDA.n1283 53.3664
R3054 GNDA.n1351 GNDA.n1282 53.3664
R3055 GNDA.n1361 GNDA.n1285 53.3664
R3056 GNDA.n1356 GNDA.n1284 53.3664
R3057 GNDA.n1352 GNDA.n1283 53.3664
R3058 GNDA.n1348 GNDA.n1282 53.3664
R3059 GNDA.n1330 GNDA.n1273 53.3664
R3060 GNDA.n1334 GNDA.n1280 53.3664
R3061 GNDA.n1338 GNDA.n1271 53.3664
R3062 GNDA.n1342 GNDA.n1281 53.3664
R3063 GNDA.n1313 GNDA.n1279 53.3664
R3064 GNDA.n1317 GNDA.n1278 53.3664
R3065 GNDA.n1321 GNDA.n1277 53.3664
R3066 GNDA.n1325 GNDA.n1276 53.3664
R3067 GNDA.n1309 GNDA.n1274 53.3664
R3068 GNDA.n1301 GNDA.n1272 53.3664
R3069 GNDA.n1362 GNDA.n1270 53.3664
R3070 GNDA.n1269 GNDA.n1266 53.3664
R3071 GNDA.n1514 GNDA.n1474 53.3664
R3072 GNDA.n1513 GNDA.n1512 53.3664
R3073 GNDA.n1506 GNDA.n1476 53.3664
R3074 GNDA.n1505 GNDA.n1504 53.3664
R3075 GNDA.n1496 GNDA.n1495 53.3664
R3076 GNDA.n1491 GNDA.n1482 53.3664
R3077 GNDA.n1489 GNDA.n1488 53.3664
R3078 GNDA.n1483 GNDA.n1458 53.3664
R3079 GNDA.n1542 GNDA.n1541 53.3664
R3080 GNDA.n1554 GNDA.n1553 53.3664
R3081 GNDA.n1557 GNDA.n1556 53.3664
R3082 GNDA.n1568 GNDA.n1567 53.3664
R3083 GNDA.n1521 GNDA.n1520 53.3664
R3084 GNDA.n1523 GNDA.n1522 53.3664
R3085 GNDA.n1528 GNDA.n1527 53.3664
R3086 GNDA.n1531 GNDA.n1530 53.3664
R3087 GNDA.n1520 GNDA.n1519 53.3664
R3088 GNDA.n1522 GNDA.n1472 53.3664
R3089 GNDA.n1529 GNDA.n1528 53.3664
R3090 GNDA.n1530 GNDA.n1470 53.3664
R3091 GNDA.n1504 GNDA.n1503 53.3664
R3092 GNDA.n1507 GNDA.n1506 53.3664
R3093 GNDA.n1512 GNDA.n1511 53.3664
R3094 GNDA.n1515 GNDA.n1514 53.3664
R3095 GNDA.n1484 GNDA.n1483 53.3664
R3096 GNDA.n1490 GNDA.n1489 53.3664
R3097 GNDA.n1482 GNDA.n1480 53.3664
R3098 GNDA.n1497 GNDA.n1496 53.3664
R3099 GNDA.n1569 GNDA.n1568 53.3664
R3100 GNDA.n1556 GNDA.n1459 53.3664
R3101 GNDA.n1555 GNDA.n1554 53.3664
R3102 GNDA.n1541 GNDA.n1464 53.3664
R3103 GNDA.n1435 GNDA.n1398 53.3664
R3104 GNDA.n1434 GNDA.n1433 53.3664
R3105 GNDA.n1427 GNDA.n1400 53.3664
R3106 GNDA.n1426 GNDA.n1425 53.3664
R3107 GNDA.n1417 GNDA.n1416 53.3664
R3108 GNDA.n1412 GNDA.n1406 53.3664
R3109 GNDA.n1410 GNDA.n1409 53.3664
R3110 GNDA.n1614 GNDA.n1382 53.3664
R3111 GNDA.n1585 GNDA.n1584 53.3664
R3112 GNDA.n1597 GNDA.n1596 53.3664
R3113 GNDA.n1600 GNDA.n1599 53.3664
R3114 GNDA.n1612 GNDA.n1611 53.3664
R3115 GNDA.n1442 GNDA.n1441 53.3664
R3116 GNDA.n1444 GNDA.n1443 53.3664
R3117 GNDA.n1449 GNDA.n1448 53.3664
R3118 GNDA.n1452 GNDA.n1451 53.3664
R3119 GNDA.n1441 GNDA.n1440 53.3664
R3120 GNDA.n1443 GNDA.n1396 53.3664
R3121 GNDA.n1450 GNDA.n1449 53.3664
R3122 GNDA.n1451 GNDA.n1394 53.3664
R3123 GNDA.n1425 GNDA.n1424 53.3664
R3124 GNDA.n1428 GNDA.n1427 53.3664
R3125 GNDA.n1433 GNDA.n1432 53.3664
R3126 GNDA.n1436 GNDA.n1435 53.3664
R3127 GNDA.n1407 GNDA.n1382 53.3664
R3128 GNDA.n1411 GNDA.n1410 53.3664
R3129 GNDA.n1406 GNDA.n1404 53.3664
R3130 GNDA.n1418 GNDA.n1417 53.3664
R3131 GNDA.n1613 GNDA.n1612 53.3664
R3132 GNDA.n1599 GNDA.n1383 53.3664
R3133 GNDA.n1598 GNDA.n1597 53.3664
R3134 GNDA.n1584 GNDA.n1388 53.3664
R3135 GNDA.n420 GNDA.n383 53.3664
R3136 GNDA.n419 GNDA.n418 53.3664
R3137 GNDA.n412 GNDA.n385 53.3664
R3138 GNDA.n411 GNDA.n410 53.3664
R3139 GNDA.n402 GNDA.n401 53.3664
R3140 GNDA.n397 GNDA.n391 53.3664
R3141 GNDA.n395 GNDA.n394 53.3664
R3142 GNDA.n1772 GNDA.n368 53.3664
R3143 GNDA.n1743 GNDA.n1742 53.3664
R3144 GNDA.n1755 GNDA.n1754 53.3664
R3145 GNDA.n1758 GNDA.n1757 53.3664
R3146 GNDA.n1770 GNDA.n1769 53.3664
R3147 GNDA.n427 GNDA.n426 53.3664
R3148 GNDA.n429 GNDA.n428 53.3664
R3149 GNDA.n434 GNDA.n433 53.3664
R3150 GNDA.n437 GNDA.n436 53.3664
R3151 GNDA.n426 GNDA.n425 53.3664
R3152 GNDA.n428 GNDA.n381 53.3664
R3153 GNDA.n435 GNDA.n434 53.3664
R3154 GNDA.n436 GNDA.n379 53.3664
R3155 GNDA.n410 GNDA.n409 53.3664
R3156 GNDA.n413 GNDA.n412 53.3664
R3157 GNDA.n418 GNDA.n417 53.3664
R3158 GNDA.n421 GNDA.n420 53.3664
R3159 GNDA.n392 GNDA.n368 53.3664
R3160 GNDA.n396 GNDA.n395 53.3664
R3161 GNDA.n391 GNDA.n389 53.3664
R3162 GNDA.n403 GNDA.n402 53.3664
R3163 GNDA.n301 GNDA.n264 53.3664
R3164 GNDA.n300 GNDA.n299 53.3664
R3165 GNDA.n293 GNDA.n266 53.3664
R3166 GNDA.n292 GNDA.n291 53.3664
R3167 GNDA.n283 GNDA.n282 53.3664
R3168 GNDA.n278 GNDA.n272 53.3664
R3169 GNDA.n276 GNDA.n275 53.3664
R3170 GNDA.n1823 GNDA.n249 53.3664
R3171 GNDA.n1794 GNDA.n1793 53.3664
R3172 GNDA.n1806 GNDA.n1805 53.3664
R3173 GNDA.n1809 GNDA.n1808 53.3664
R3174 GNDA.n1821 GNDA.n1820 53.3664
R3175 GNDA.n308 GNDA.n307 53.3664
R3176 GNDA.n310 GNDA.n309 53.3664
R3177 GNDA.n315 GNDA.n314 53.3664
R3178 GNDA.n318 GNDA.n317 53.3664
R3179 GNDA.n307 GNDA.n306 53.3664
R3180 GNDA.n309 GNDA.n262 53.3664
R3181 GNDA.n316 GNDA.n315 53.3664
R3182 GNDA.n317 GNDA.n260 53.3664
R3183 GNDA.n291 GNDA.n290 53.3664
R3184 GNDA.n294 GNDA.n293 53.3664
R3185 GNDA.n299 GNDA.n298 53.3664
R3186 GNDA.n302 GNDA.n301 53.3664
R3187 GNDA.n273 GNDA.n249 53.3664
R3188 GNDA.n277 GNDA.n276 53.3664
R3189 GNDA.n272 GNDA.n270 53.3664
R3190 GNDA.n284 GNDA.n283 53.3664
R3191 GNDA.n1822 GNDA.n1821 53.3664
R3192 GNDA.n1808 GNDA.n250 53.3664
R3193 GNDA.n1807 GNDA.n1806 53.3664
R3194 GNDA.n1793 GNDA.n255 53.3664
R3195 GNDA.n1771 GNDA.n1770 53.3664
R3196 GNDA.n1757 GNDA.n369 53.3664
R3197 GNDA.n1756 GNDA.n1755 53.3664
R3198 GNDA.n1742 GNDA.n374 53.3664
R3199 GNDA.n963 GNDA.n58 53.3664
R3200 GNDA.n967 GNDA.n48 53.3664
R3201 GNDA.n971 GNDA.n57 53.3664
R3202 GNDA.n975 GNDA.n50 53.3664
R3203 GNDA.n986 GNDA.n53 53.3664
R3204 GNDA.n990 GNDA.n54 53.3664
R3205 GNDA.n994 GNDA.n55 53.3664
R3206 GNDA.n1009 GNDA.n56 53.3664
R3207 GNDA.n64 GNDA.n47 53.3664
R3208 GNDA.n2084 GNDA.n49 53.3664
R3209 GNDA.n2097 GNDA.n2096 53.3664
R3210 GNDA.n998 GNDA.n51 53.3664
R3211 GNDA.n959 GNDA.n62 53.3664
R3212 GNDA.n958 GNDA.n61 53.3664
R3213 GNDA.n954 GNDA.n60 53.3664
R3214 GNDA.n950 GNDA.n59 53.3664
R3215 GNDA.n962 GNDA.n62 53.3664
R3216 GNDA.n955 GNDA.n61 53.3664
R3217 GNDA.n951 GNDA.n60 53.3664
R3218 GNDA.n947 GNDA.n59 53.3664
R3219 GNDA.n978 GNDA.n50 53.3664
R3220 GNDA.n974 GNDA.n57 53.3664
R3221 GNDA.n970 GNDA.n48 53.3664
R3222 GNDA.n966 GNDA.n58 53.3664
R3223 GNDA.n995 GNDA.n56 53.3664
R3224 GNDA.n991 GNDA.n55 53.3664
R3225 GNDA.n987 GNDA.n54 53.3664
R3226 GNDA.n983 GNDA.n53 53.3664
R3227 GNDA.n1010 GNDA.n51 53.3664
R3228 GNDA.n2096 GNDA.n46 53.3664
R3229 GNDA.n49 GNDA.n45 53.3664
R3230 GNDA.n2083 GNDA.n47 53.3664
R3231 GNDA.n2013 GNDA.n97 53.3664
R3232 GNDA.n2009 GNDA.n87 53.3664
R3233 GNDA.n2005 GNDA.n96 53.3664
R3234 GNDA.n2001 GNDA.n89 53.3664
R3235 GNDA.n1990 GNDA.n92 53.3664
R3236 GNDA.n1986 GNDA.n93 53.3664
R3237 GNDA.n1982 GNDA.n94 53.3664
R3238 GNDA.n1978 GNDA.n95 53.3664
R3239 GNDA.n103 GNDA.n86 53.3664
R3240 GNDA.n2042 GNDA.n88 53.3664
R3241 GNDA.n2055 GNDA.n2054 53.3664
R3242 GNDA.n119 GNDA.n90 53.3664
R3243 GNDA.n2017 GNDA.n101 53.3664
R3244 GNDA.n2018 GNDA.n100 53.3664
R3245 GNDA.n2022 GNDA.n99 53.3664
R3246 GNDA.n2026 GNDA.n98 53.3664
R3247 GNDA.n2014 GNDA.n101 53.3664
R3248 GNDA.n2021 GNDA.n100 53.3664
R3249 GNDA.n2025 GNDA.n99 53.3664
R3250 GNDA.n2028 GNDA.n98 53.3664
R3251 GNDA.n1998 GNDA.n89 53.3664
R3252 GNDA.n2002 GNDA.n96 53.3664
R3253 GNDA.n2006 GNDA.n87 53.3664
R3254 GNDA.n2010 GNDA.n97 53.3664
R3255 GNDA.n1981 GNDA.n95 53.3664
R3256 GNDA.n1985 GNDA.n94 53.3664
R3257 GNDA.n1989 GNDA.n93 53.3664
R3258 GNDA.n1993 GNDA.n92 53.3664
R3259 GNDA.n1977 GNDA.n90 53.3664
R3260 GNDA.n2054 GNDA.n85 53.3664
R3261 GNDA.n88 GNDA.n84 53.3664
R3262 GNDA.n2041 GNDA.n86 53.3664
R3263 GNDA.n1856 GNDA.n234 52.7091
R3264 GNDA.n1850 GNDA.n234 52.7091
R3265 GNDA.n1850 GNDA.n1849 52.7091
R3266 GNDA.n1849 GNDA.n1848 52.7091
R3267 GNDA.n1848 GNDA.n147 52.7091
R3268 GNDA.n1841 GNDA.n146 52.7091
R3269 GNDA.n1841 GNDA.n1840 52.7091
R3270 GNDA.n1840 GNDA.n1839 52.7091
R3271 GNDA.n1839 GNDA.n241 52.7091
R3272 GNDA.n1832 GNDA.n241 52.7091
R3273 GNDA.n1832 GNDA.n1831 52.7091
R3274 GNDA.n1831 GNDA.t121 52.7091
R3275 GNDA.n1643 GNDA.n1642 52.7091
R3276 GNDA.n1642 GNDA.n1641 52.7091
R3277 GNDA.n1641 GNDA.n564 52.7091
R3278 GNDA.n1635 GNDA.n564 52.7091
R3279 GNDA.n1635 GNDA.n153 52.7091
R3280 GNDA.n571 GNDA.n152 52.7091
R3281 GNDA.n1628 GNDA.n571 52.7091
R3282 GNDA.n1628 GNDA.n1627 52.7091
R3283 GNDA.n1627 GNDA.n1626 52.7091
R3284 GNDA.n1626 GNDA.n572 52.7091
R3285 GNDA.n572 GNDA.n178 52.7091
R3286 GNDA.n1937 GNDA.n138 52.7091
R3287 GNDA.n1944 GNDA.n138 52.7091
R3288 GNDA.n1945 GNDA.n1944 52.7091
R3289 GNDA.n1946 GNDA.n1945 52.7091
R3290 GNDA.n1946 GNDA.n79 52.7091
R3291 GNDA.n133 GNDA.n80 52.7091
R3292 GNDA.n1955 GNDA.n133 52.7091
R3293 GNDA.n1956 GNDA.n1955 52.7091
R3294 GNDA.n1957 GNDA.n1956 52.7091
R3295 GNDA.n1957 GNDA.n128 52.7091
R3296 GNDA.n1962 GNDA.n128 52.7091
R3297 GNDA.n1156 GNDA.t221 51.4866
R3298 GNDA.n1036 GNDA.t221 51.4866
R3299 GNDA.t169 GNDA.t57 49.9132
R3300 GNDA.t27 GNDA.t357 49.9132
R3301 GNDA.t350 GNDA.t80 49.9132
R3302 GNDA.t136 GNDA.t55 49.9132
R3303 GNDA.t187 GNDA.n2089 49.4271
R3304 GNDA.n1028 GNDA.t100 48.3974
R3305 GNDA.n2356 GNDA.t31 48.0005
R3306 GNDA.n2356 GNDA.t16 48.0005
R3307 GNDA.n2354 GNDA.t70 48.0005
R3308 GNDA.n2354 GNDA.t128 48.0005
R3309 GNDA.n2352 GNDA.t99 48.0005
R3310 GNDA.n2352 GNDA.t97 48.0005
R3311 GNDA.n2350 GNDA.t18 48.0005
R3312 GNDA.n2350 GNDA.t151 48.0005
R3313 GNDA.n2348 GNDA.t6 48.0005
R3314 GNDA.n2348 GNDA.t72 48.0005
R3315 GNDA.t24 GNDA.n855 47.3677
R3316 GNDA.t275 GNDA.t122 46.338
R3317 GNDA.t269 GNDA.t135 46.338
R3318 GNDA.t221 GNDA.n187 46.2335
R3319 GNDA.t221 GNDA.n203 46.2335
R3320 GNDA.t221 GNDA.n226 46.2335
R3321 GNDA.n2425 GNDA.n2114 46.0738
R3322 GNDA.n2409 GNDA.n2217 46.0738
R3323 GNDA.t132 GNDA.t286 46.0738
R3324 GNDA.t22 GNDA.t0 46.0738
R3325 GNDA.t111 GNDA.t330 46.0738
R3326 GNDA.t329 GNDA.t163 46.0738
R3327 GNDA.t347 GNDA.t175 46.0738
R3328 GNDA.t35 GNDA.t152 46.0738
R3329 GNDA.t50 GNDA.t167 46.0738
R3330 GNDA.t301 GNDA.t45 46.0738
R3331 GNDA.n2548 GNDA.n2536 46.0738
R3332 GNDA.n2496 GNDA.n2452 46.0738
R3333 GNDA.n1232 GNDA.t275 43.2488
R3334 GNDA.n2090 GNDA.t187 43.2488
R3335 GNDA.n2047 GNDA.t203 43.2488
R3336 GNDA.n1922 GNDA.t221 42.2987
R3337 GNDA.n1891 GNDA.t221 42.2987
R3338 GNDA.n1866 GNDA.t221 42.2987
R3339 GNDA.t139 GNDA.t93 42.2405
R3340 GNDA.t64 GNDA.t139 42.2405
R3341 GNDA.t161 GNDA.t4 42.2405
R3342 GNDA.t32 GNDA.t161 42.2405
R3343 GNDA.n2378 GNDA.t52 42.2344
R3344 GNDA.n2078 GNDA.t335 42.2191
R3345 GNDA.t221 GNDA.t24 41.1894
R3346 GNDA.t100 GNDA.t221 41.1894
R3347 GNDA.t112 GNDA.t94 39.8575
R3348 GNDA.n2074 GNDA.n70 39.3903
R3349 GNDA.n851 GNDA.t183 39.1299
R3350 GNDA.n2102 GNDA.n2101 39.1299
R3351 GNDA.n1006 GNDA.t199 39.1299
R3352 GNDA.n1973 GNDA.t269 39.1299
R3353 GNDA.t286 GNDA.t22 38.3949
R3354 GNDA.t0 GNDA.t111 38.3949
R3355 GNDA.t330 GNDA.t329 38.3949
R3356 GNDA.t163 GNDA.t347 38.3949
R3357 GNDA.t175 GNDA.t35 38.3949
R3358 GNDA.t152 GNDA.t50 38.3949
R3359 GNDA.t167 GNDA.t301 38.3949
R3360 GNDA.n1156 GNDA.n1155 38.1002
R3361 GNDA.n1005 GNDA.n69 38.1002
R3362 GNDA.n2059 GNDA.t14 38.1002
R3363 GNDA.n1973 GNDA.t67 38.1002
R3364 GNDA.n1037 GNDA.n1036 37.0705
R3365 GNDA.t221 GNDA.t209 36.0408
R3366 GNDA.t221 GNDA.t189 36.0408
R3367 GNDA.t221 GNDA.n147 35.7252
R3368 GNDA.t221 GNDA.n153 35.7252
R3369 GNDA.t221 GNDA.n79 35.7252
R3370 GNDA.n2073 GNDA.n2072 35.3278
R3371 GNDA.t38 GNDA.t169 34.5555
R3372 GNDA.t357 GNDA.t61 34.5555
R3373 GNDA.t80 GNDA.t2 34.5555
R3374 GNDA.t334 GNDA.t136 34.5555
R3375 GNDA.t103 GNDA.n1232 33.9813
R3376 GNDA.n835 GNDA.t89 33.9813
R3377 GNDA.n2077 GNDA.n2076 33.9813
R3378 GNDA.n826 GNDA.t193 32.9516
R3379 GNDA.t215 GNDA.n1003 32.9516
R3380 GNDA.t205 GNDA.n123 32.9516
R3381 GNDA.t221 GNDA.n154 32.9056
R3382 GNDA.t221 GNDA.n179 32.9056
R3383 GNDA.n1966 GNDA.n1965 32.3063
R3384 GNDA.t120 GNDA.t328 30.716
R3385 GNDA.t289 GNDA.t143 30.716
R3386 GNDA.t9 GNDA.t171 30.716
R3387 GNDA.t62 GNDA.t336 30.716
R3388 GNDA.t34 GNDA.t155 30.716
R3389 GNDA.t82 GNDA.t325 30.716
R3390 GNDA.t140 GNDA.t147 30.716
R3391 GNDA.t320 GNDA.t173 30.716
R3392 GNDA.t49 GNDA.t47 30.716
R3393 GNDA.t12 GNDA.t310 30.716
R3394 GNDA.n2556 GNDA.n0 29.8047
R3395 GNDA.t351 GNDA.n110 29.2831
R3396 GNDA.n833 GNDA.t191 28.8327
R3397 GNDA.t213 GNDA.n2088 28.8327
R3398 GNDA.t207 GNDA.n2036 28.8327
R3399 GNDA.t321 GNDA.n833 27.803
R3400 GNDA.t88 GNDA.n850 27.803
R3401 GNDA.n1164 GNDA.t59 27.803
R3402 GNDA.n706 GNDA.n703 27.5561
R3403 GNDA.n1207 GNDA.n1204 27.5561
R3404 GNDA.n1346 GNDA.n1345 27.5561
R3405 GNDA.n1518 GNDA.n1517 27.5561
R3406 GNDA.n1439 GNDA.n1438 27.5561
R3407 GNDA.n424 GNDA.n423 27.5561
R3408 GNDA.n305 GNDA.n304 27.5561
R3409 GNDA.n964 GNDA.n961 27.5561
R3410 GNDA.n2015 GNDA.n2012 27.5561
R3411 GNDA.n2319 GNDA.t149 26.8766
R3412 GNDA.n2384 GNDA.t165 26.8766
R3413 GNDA.t123 GNDA.t131 26.8766
R3414 GNDA.n687 GNDA.n686 26.6672
R3415 GNDA.n1188 GNDA.n1187 26.6672
R3416 GNDA.n1328 GNDA.n1327 26.6672
R3417 GNDA.n1501 GNDA.n1500 26.6672
R3418 GNDA.n1422 GNDA.n1421 26.6672
R3419 GNDA.n407 GNDA.n406 26.6672
R3420 GNDA.n288 GNDA.n287 26.6672
R3421 GNDA.n981 GNDA.n980 26.6672
R3422 GNDA.n1996 GNDA.n1995 26.6672
R3423 GNDA.t183 GNDA.t88 25.7435
R3424 GNDA.t203 GNDA.t101 25.7435
R3425 GNDA.n171 GNDA.n161 25.3679
R3426 GNDA.n2230 GNDA.n2229 24.991
R3427 GNDA.n2392 GNDA.n2391 24.7472
R3428 GNDA.n2556 GNDA.n2555 24.133
R3429 GNDA.n858 GNDA.t192 24.0005
R3430 GNDA.n858 GNDA.t182 24.0005
R3431 GNDA.n860 GNDA.t210 24.0005
R3432 GNDA.n860 GNDA.t194 24.0005
R3433 GNDA.n862 GNDA.t184 24.0005
R3434 GNDA.n862 GNDA.t212 24.0005
R3435 GNDA.n864 GNDA.t198 24.0005
R3436 GNDA.n864 GNDA.t188 24.0005
R3437 GNDA.n1018 GNDA.t214 24.0005
R3438 GNDA.n1018 GNDA.t196 24.0005
R3439 GNDA.n1020 GNDA.t186 24.0005
R3440 GNDA.n1020 GNDA.t216 24.0005
R3441 GNDA.n1022 GNDA.t200 24.0005
R3442 GNDA.n1022 GNDA.t202 24.0005
R3443 GNDA.n1026 GNDA.t180 24.0005
R3444 GNDA.n1026 GNDA.t204 24.0005
R3445 GNDA.n1024 GNDA.t208 24.0005
R3446 GNDA.n1024 GNDA.t190 24.0005
R3447 GNDA.n125 GNDA.t178 24.0005
R3448 GNDA.n125 GNDA.t206 24.0005
R3449 GNDA.n2034 GNDA.t79 23.6841
R3450 GNDA.t101 GNDA.n2046 23.6841
R3451 GNDA.n123 GNDA.t353 23.6841
R3452 GNDA.n2388 GNDA.n2386 23.6611
R3453 GNDA.n2267 GNDA.n2266 23.6611
R3454 GNDA.n2191 GNDA.n2190 22.8576
R3455 GNDA.n2322 GNDA.n2321 22.8576
R3456 GNDA.n2285 GNDA.n2284 22.8576
R3457 GNDA.n2412 GNDA.n2411 22.8576
R3458 GNDA.n2415 GNDA.n2414 22.8576
R3459 GNDA.n2329 GNDA.n2328 22.8576
R3460 GNDA.n2339 GNDA.n2338 22.8576
R3461 GNDA.n2372 GNDA.n2371 22.8576
R3462 GNDA.n2369 GNDA.n2368 22.8576
R3463 GNDA.n2551 GNDA.n2550 22.8576
R3464 GNDA.n2442 GNDA.n15 22.8576
R3465 GNDA.n2510 GNDA.n2509 22.8576
R3466 GNDA.n2470 GNDA.n2469 22.8576
R3467 GNDA.n2184 GNDA.n2183 22.8576
R3468 GNDA.t197 GNDA.n2077 22.6544
R3469 GNDA.n2048 GNDA.t179 22.6544
R3470 GNDA.t351 GNDA.n108 21.084
R3471 GNDA.n211 GNDA.n210 21.0192
R3472 GNDA.t113 GNDA.t63 20.9779
R3473 GNDA.n857 GNDA.n856 20.8233
R3474 GNDA.n1162 GNDA.n1161 20.8233
R3475 GNDA.n1158 GNDA.n1157 20.8233
R3476 GNDA.n1035 GNDA.n1034 20.8233
R3477 GNDA.n1031 GNDA.n1030 20.8233
R3478 GNDA.n1970 GNDA.n1969 20.8233
R3479 GNDA.t221 GNDA.n174 20.5949
R3480 GNDA.t102 GNDA.n174 20.5949
R3481 GNDA.t59 GNDA.n1163 20.5949
R3482 GNDA.n1029 GNDA.t79 20.5949
R3483 GNDA.n2070 GNDA.t13 20.5949
R3484 GNDA.n2070 GNDA.t221 20.5949
R3485 GNDA.t221 GNDA.n142 19.9378
R3486 GNDA.n2256 GNDA.t39 19.7005
R3487 GNDA.n2256 GNDA.t313 19.7005
R3488 GNDA.n2254 GNDA.t142 19.7005
R3489 GNDA.n2254 GNDA.t58 19.7005
R3490 GNDA.n2252 GNDA.t333 19.7005
R3491 GNDA.n2252 GNDA.t108 19.7005
R3492 GNDA.n2250 GNDA.t91 19.7005
R3493 GNDA.n2250 GNDA.t23 19.7005
R3494 GNDA.n2248 GNDA.t141 19.7005
R3495 GNDA.n2248 GNDA.t86 19.7005
R3496 GNDA.n2247 GNDA.t314 19.7005
R3497 GNDA.n2247 GNDA.t134 19.7005
R3498 GNDA.n12 GNDA.t324 19.7005
R3499 GNDA.n12 GNDA.t349 19.7005
R3500 GNDA.n10 GNDA.t107 19.7005
R3501 GNDA.n10 GNDA.t53 19.7005
R3502 GNDA.n8 GNDA.t117 19.7005
R3503 GNDA.n8 GNDA.t118 19.7005
R3504 GNDA.n6 GNDA.t338 19.7005
R3505 GNDA.n6 GNDA.t354 19.7005
R3506 GNDA.n4 GNDA.t327 19.7005
R3507 GNDA.n4 GNDA.t105 19.7005
R3508 GNDA.n3 GNDA.t115 19.7005
R3509 GNDA.n3 GNDA.t323 19.7005
R3510 GNDA.t221 GNDA.n1936 19.6741
R3511 GNDA.n2360 GNDA.n2359 19.2005
R3512 GNDA.n2347 GNDA.n2346 19.2005
R3513 GNDA.t332 GNDA.t40 19.1977
R3514 GNDA.t42 GNDA.t85 19.1977
R3515 GNDA.t109 GNDA.t116 19.1977
R3516 GNDA.t114 GNDA.t36 19.1977
R3517 GNDA.n2231 GNDA.n2230 18.5713
R3518 GNDA.n1894 GNDA.n205 18.5605
R3519 GNDA.n852 GNDA.t211 18.5355
R3520 GNDA.t201 GNDA.n1005 18.5355
R3521 GNDA.n2437 GNDA.t95 18.3557
R3522 GNDA GNDA.n72 18.1546
R3523 GNDA.n2414 GNDA.n2413 18.1442
R3524 GNDA.n2552 GNDA.n15 18.1442
R3525 GNDA.n2370 GNDA.n2369 17.8005
R3526 GNDA.n1646 GNDA.n561 17.5843
R3527 GNDA.n1854 GNDA.n232 17.5843
R3528 GNDA.n1939 GNDA.n140 17.5843
R3529 GNDA.t221 GNDA.n176 17.5058
R3530 GNDA.n1971 GNDA.n108 17.5058
R3531 GNDA.t221 GNDA.n146 16.9844
R3532 GNDA.t221 GNDA.n152 16.9844
R3533 GNDA.t221 GNDA.n80 16.9844
R3534 GNDA.n1934 GNDA.n184 16.9379
R3535 GNDA.n1255 GNDA.n797 16.9379
R3536 GNDA.n770 GNDA.n740 16.9379
R3537 GNDA.n552 GNDA.n323 16.7709
R3538 GNDA.n918 GNDA.n511 16.7709
R3539 GNDA.n1731 GNDA.n1730 16.7709
R3540 GNDA.n909 GNDA.n508 16.7709
R3541 GNDA.n707 GNDA.n706 16.0005
R3542 GNDA.n710 GNDA.n707 16.0005
R3543 GNDA.n711 GNDA.n710 16.0005
R3544 GNDA.n714 GNDA.n711 16.0005
R3545 GNDA.n715 GNDA.n714 16.0005
R3546 GNDA.n718 GNDA.n715 16.0005
R3547 GNDA.n719 GNDA.n718 16.0005
R3548 GNDA.n719 GNDA.n612 16.0005
R3549 GNDA.n703 GNDA.n702 16.0005
R3550 GNDA.n702 GNDA.n699 16.0005
R3551 GNDA.n699 GNDA.n698 16.0005
R3552 GNDA.n698 GNDA.n695 16.0005
R3553 GNDA.n695 GNDA.n694 16.0005
R3554 GNDA.n694 GNDA.n691 16.0005
R3555 GNDA.n691 GNDA.n690 16.0005
R3556 GNDA.n690 GNDA.n687 16.0005
R3557 GNDA.n686 GNDA.n683 16.0005
R3558 GNDA.n683 GNDA.n682 16.0005
R3559 GNDA.n682 GNDA.n679 16.0005
R3560 GNDA.n679 GNDA.n678 16.0005
R3561 GNDA.n678 GNDA.n675 16.0005
R3562 GNDA.n675 GNDA.n674 16.0005
R3563 GNDA.n674 GNDA.n671 16.0005
R3564 GNDA.n671 GNDA.n670 16.0005
R3565 GNDA.n1208 GNDA.n1207 16.0005
R3566 GNDA.n1211 GNDA.n1208 16.0005
R3567 GNDA.n1212 GNDA.n1211 16.0005
R3568 GNDA.n1215 GNDA.n1212 16.0005
R3569 GNDA.n1216 GNDA.n1215 16.0005
R3570 GNDA.n1219 GNDA.n1216 16.0005
R3571 GNDA.n1220 GNDA.n1219 16.0005
R3572 GNDA.n1223 GNDA.n1220 16.0005
R3573 GNDA.n1204 GNDA.n1203 16.0005
R3574 GNDA.n1203 GNDA.n1200 16.0005
R3575 GNDA.n1200 GNDA.n1199 16.0005
R3576 GNDA.n1199 GNDA.n1196 16.0005
R3577 GNDA.n1196 GNDA.n1195 16.0005
R3578 GNDA.n1195 GNDA.n1192 16.0005
R3579 GNDA.n1192 GNDA.n1191 16.0005
R3580 GNDA.n1191 GNDA.n1188 16.0005
R3581 GNDA.n1187 GNDA.n1184 16.0005
R3582 GNDA.n1184 GNDA.n1183 16.0005
R3583 GNDA.n1183 GNDA.n1180 16.0005
R3584 GNDA.n1180 GNDA.n1179 16.0005
R3585 GNDA.n1179 GNDA.n1176 16.0005
R3586 GNDA.n1176 GNDA.n1175 16.0005
R3587 GNDA.n1175 GNDA.n1172 16.0005
R3588 GNDA.n1172 GNDA.n1171 16.0005
R3589 GNDA.n1359 GNDA.n1346 16.0005
R3590 GNDA.n1359 GNDA.n1358 16.0005
R3591 GNDA.n1358 GNDA.n1357 16.0005
R3592 GNDA.n1357 GNDA.n1354 16.0005
R3593 GNDA.n1354 GNDA.n1353 16.0005
R3594 GNDA.n1353 GNDA.n1350 16.0005
R3595 GNDA.n1350 GNDA.n1349 16.0005
R3596 GNDA.n1349 GNDA.n1262 16.0005
R3597 GNDA.n1345 GNDA.n1343 16.0005
R3598 GNDA.n1343 GNDA.n1340 16.0005
R3599 GNDA.n1340 GNDA.n1339 16.0005
R3600 GNDA.n1339 GNDA.n1336 16.0005
R3601 GNDA.n1336 GNDA.n1335 16.0005
R3602 GNDA.n1335 GNDA.n1332 16.0005
R3603 GNDA.n1332 GNDA.n1331 16.0005
R3604 GNDA.n1331 GNDA.n1328 16.0005
R3605 GNDA.n1327 GNDA.n1324 16.0005
R3606 GNDA.n1324 GNDA.n1323 16.0005
R3607 GNDA.n1323 GNDA.n1320 16.0005
R3608 GNDA.n1320 GNDA.n1319 16.0005
R3609 GNDA.n1319 GNDA.n1316 16.0005
R3610 GNDA.n1316 GNDA.n1315 16.0005
R3611 GNDA.n1315 GNDA.n1312 16.0005
R3612 GNDA.n1312 GNDA.n1311 16.0005
R3613 GNDA.n1518 GNDA.n1473 16.0005
R3614 GNDA.n1524 GNDA.n1473 16.0005
R3615 GNDA.n1525 GNDA.n1524 16.0005
R3616 GNDA.n1526 GNDA.n1525 16.0005
R3617 GNDA.n1526 GNDA.n1471 16.0005
R3618 GNDA.n1532 GNDA.n1471 16.0005
R3619 GNDA.n1533 GNDA.n1532 16.0005
R3620 GNDA.n1537 GNDA.n1533 16.0005
R3621 GNDA.n1517 GNDA.n1516 16.0005
R3622 GNDA.n1516 GNDA.n1475 16.0005
R3623 GNDA.n1510 GNDA.n1475 16.0005
R3624 GNDA.n1510 GNDA.n1509 16.0005
R3625 GNDA.n1509 GNDA.n1508 16.0005
R3626 GNDA.n1508 GNDA.n1477 16.0005
R3627 GNDA.n1502 GNDA.n1477 16.0005
R3628 GNDA.n1502 GNDA.n1501 16.0005
R3629 GNDA.n1500 GNDA.n1479 16.0005
R3630 GNDA.n1494 GNDA.n1479 16.0005
R3631 GNDA.n1494 GNDA.n1493 16.0005
R3632 GNDA.n1493 GNDA.n1492 16.0005
R3633 GNDA.n1492 GNDA.n1481 16.0005
R3634 GNDA.n1487 GNDA.n1481 16.0005
R3635 GNDA.n1487 GNDA.n1486 16.0005
R3636 GNDA.n1486 GNDA.n1485 16.0005
R3637 GNDA.n1439 GNDA.n1397 16.0005
R3638 GNDA.n1445 GNDA.n1397 16.0005
R3639 GNDA.n1446 GNDA.n1445 16.0005
R3640 GNDA.n1447 GNDA.n1446 16.0005
R3641 GNDA.n1447 GNDA.n1395 16.0005
R3642 GNDA.n1453 GNDA.n1395 16.0005
R3643 GNDA.n1454 GNDA.n1453 16.0005
R3644 GNDA.n1580 GNDA.n1454 16.0005
R3645 GNDA.n1438 GNDA.n1437 16.0005
R3646 GNDA.n1437 GNDA.n1399 16.0005
R3647 GNDA.n1431 GNDA.n1399 16.0005
R3648 GNDA.n1431 GNDA.n1430 16.0005
R3649 GNDA.n1430 GNDA.n1429 16.0005
R3650 GNDA.n1429 GNDA.n1401 16.0005
R3651 GNDA.n1423 GNDA.n1401 16.0005
R3652 GNDA.n1423 GNDA.n1422 16.0005
R3653 GNDA.n1421 GNDA.n1403 16.0005
R3654 GNDA.n1415 GNDA.n1403 16.0005
R3655 GNDA.n1415 GNDA.n1414 16.0005
R3656 GNDA.n1414 GNDA.n1413 16.0005
R3657 GNDA.n1413 GNDA.n1405 16.0005
R3658 GNDA.n1408 GNDA.n1405 16.0005
R3659 GNDA.n1408 GNDA.n1381 16.0005
R3660 GNDA.n1615 GNDA.n1381 16.0005
R3661 GNDA.n424 GNDA.n382 16.0005
R3662 GNDA.n430 GNDA.n382 16.0005
R3663 GNDA.n431 GNDA.n430 16.0005
R3664 GNDA.n432 GNDA.n431 16.0005
R3665 GNDA.n432 GNDA.n380 16.0005
R3666 GNDA.n438 GNDA.n380 16.0005
R3667 GNDA.n439 GNDA.n438 16.0005
R3668 GNDA.n1738 GNDA.n439 16.0005
R3669 GNDA.n423 GNDA.n422 16.0005
R3670 GNDA.n422 GNDA.n384 16.0005
R3671 GNDA.n416 GNDA.n384 16.0005
R3672 GNDA.n416 GNDA.n415 16.0005
R3673 GNDA.n415 GNDA.n414 16.0005
R3674 GNDA.n414 GNDA.n386 16.0005
R3675 GNDA.n408 GNDA.n386 16.0005
R3676 GNDA.n408 GNDA.n407 16.0005
R3677 GNDA.n406 GNDA.n388 16.0005
R3678 GNDA.n400 GNDA.n388 16.0005
R3679 GNDA.n400 GNDA.n399 16.0005
R3680 GNDA.n399 GNDA.n398 16.0005
R3681 GNDA.n398 GNDA.n390 16.0005
R3682 GNDA.n393 GNDA.n390 16.0005
R3683 GNDA.n393 GNDA.n367 16.0005
R3684 GNDA.n1773 GNDA.n367 16.0005
R3685 GNDA.n305 GNDA.n263 16.0005
R3686 GNDA.n311 GNDA.n263 16.0005
R3687 GNDA.n312 GNDA.n311 16.0005
R3688 GNDA.n313 GNDA.n312 16.0005
R3689 GNDA.n313 GNDA.n261 16.0005
R3690 GNDA.n319 GNDA.n261 16.0005
R3691 GNDA.n320 GNDA.n319 16.0005
R3692 GNDA.n1789 GNDA.n320 16.0005
R3693 GNDA.n304 GNDA.n303 16.0005
R3694 GNDA.n303 GNDA.n265 16.0005
R3695 GNDA.n297 GNDA.n265 16.0005
R3696 GNDA.n297 GNDA.n296 16.0005
R3697 GNDA.n296 GNDA.n295 16.0005
R3698 GNDA.n295 GNDA.n267 16.0005
R3699 GNDA.n289 GNDA.n267 16.0005
R3700 GNDA.n289 GNDA.n288 16.0005
R3701 GNDA.n287 GNDA.n269 16.0005
R3702 GNDA.n281 GNDA.n269 16.0005
R3703 GNDA.n281 GNDA.n280 16.0005
R3704 GNDA.n280 GNDA.n279 16.0005
R3705 GNDA.n279 GNDA.n271 16.0005
R3706 GNDA.n274 GNDA.n271 16.0005
R3707 GNDA.n274 GNDA.n248 16.0005
R3708 GNDA.n1824 GNDA.n248 16.0005
R3709 GNDA.n961 GNDA.n960 16.0005
R3710 GNDA.n960 GNDA.n957 16.0005
R3711 GNDA.n957 GNDA.n956 16.0005
R3712 GNDA.n956 GNDA.n953 16.0005
R3713 GNDA.n953 GNDA.n952 16.0005
R3714 GNDA.n952 GNDA.n949 16.0005
R3715 GNDA.n949 GNDA.n948 16.0005
R3716 GNDA.n948 GNDA.n946 16.0005
R3717 GNDA.n965 GNDA.n964 16.0005
R3718 GNDA.n968 GNDA.n965 16.0005
R3719 GNDA.n969 GNDA.n968 16.0005
R3720 GNDA.n972 GNDA.n969 16.0005
R3721 GNDA.n973 GNDA.n972 16.0005
R3722 GNDA.n976 GNDA.n973 16.0005
R3723 GNDA.n977 GNDA.n976 16.0005
R3724 GNDA.n980 GNDA.n977 16.0005
R3725 GNDA.n984 GNDA.n981 16.0005
R3726 GNDA.n985 GNDA.n984 16.0005
R3727 GNDA.n988 GNDA.n985 16.0005
R3728 GNDA.n989 GNDA.n988 16.0005
R3729 GNDA.n992 GNDA.n989 16.0005
R3730 GNDA.n993 GNDA.n992 16.0005
R3731 GNDA.n996 GNDA.n993 16.0005
R3732 GNDA.n997 GNDA.n996 16.0005
R3733 GNDA.n2016 GNDA.n2015 16.0005
R3734 GNDA.n2019 GNDA.n2016 16.0005
R3735 GNDA.n2020 GNDA.n2019 16.0005
R3736 GNDA.n2023 GNDA.n2020 16.0005
R3737 GNDA.n2024 GNDA.n2023 16.0005
R3738 GNDA.n2027 GNDA.n2024 16.0005
R3739 GNDA.n2029 GNDA.n2027 16.0005
R3740 GNDA.n2030 GNDA.n2029 16.0005
R3741 GNDA.n2012 GNDA.n2011 16.0005
R3742 GNDA.n2011 GNDA.n2008 16.0005
R3743 GNDA.n2008 GNDA.n2007 16.0005
R3744 GNDA.n2007 GNDA.n2004 16.0005
R3745 GNDA.n2004 GNDA.n2003 16.0005
R3746 GNDA.n2003 GNDA.n2000 16.0005
R3747 GNDA.n2000 GNDA.n1999 16.0005
R3748 GNDA.n1999 GNDA.n1996 16.0005
R3749 GNDA.n1995 GNDA.n1992 16.0005
R3750 GNDA.n1992 GNDA.n1991 16.0005
R3751 GNDA.n1991 GNDA.n1988 16.0005
R3752 GNDA.n1988 GNDA.n1987 16.0005
R3753 GNDA.n1987 GNDA.n1984 16.0005
R3754 GNDA.n1984 GNDA.n1983 16.0005
R3755 GNDA.n1983 GNDA.n1980 16.0005
R3756 GNDA.n1980 GNDA.n1979 16.0005
R3757 GNDA.n212 GNDA.n211 16.0005
R3758 GNDA.n212 GNDA.n205 16.0005
R3759 GNDA.n2221 GNDA.t293 16.0005
R3760 GNDA.n2232 GNDA.t305 16.0005
R3761 GNDA.n2381 GNDA.t302 16.0005
R3762 GNDA.n2264 GNDA.t290 16.0005
R3763 GNDA.n2269 GNDA.t267 16.0005
R3764 GNDA.n2224 GNDA.t299 16.0005
R3765 GNDA.n2246 GNDA.t231 16.0005
R3766 GNDA.n2337 GNDA.t246 16.0005
R3767 GNDA.n2240 GNDA.t225 16.0005
R3768 GNDA.n2362 GNDA.t243 16.0005
R3769 GNDA.t211 GNDA.t87 15.4463
R3770 GNDA.t179 GNDA.t25 15.4463
R3771 GNDA.n2469 GNDA.n2468 14.9255
R3772 GNDA.n2186 GNDA.n2184 14.9255
R3773 GNDA.n1378 GNDA.n154 14.555
R3774 GNDA.n245 GNDA.n179 14.555
R3775 GNDA.n859 GNDA.n857 14.363
R3776 GNDA.n2349 GNDA.n2347 14.363
R3777 GNDA.n2391 GNDA.n2390 14.3213
R3778 GNDA.n2389 GNDA.n2388 14.3213
R3779 GNDA.n2266 GNDA.n2231 14.3213
R3780 GNDA.n2287 GNDA.n2285 14.0818
R3781 GNDA.n2413 GNDA.n2412 14.0193
R3782 GNDA.n2552 GNDA.n2551 14.0193
R3783 GNDA.n1161 GNDA.n1160 13.8005
R3784 GNDA.n1159 GNDA.n1158 13.8005
R3785 GNDA.n1034 GNDA.n1033 13.8005
R3786 GNDA.n1032 GNDA.n1031 13.8005
R3787 GNDA.n1969 GNDA.n1968 13.8005
R3788 GNDA.n2190 GNDA.n2189 13.8005
R3789 GNDA.n2323 GNDA.n2322 13.8005
R3790 GNDA.n2328 GNDA.n2327 13.8005
R3791 GNDA.n2338 GNDA.n2241 13.8005
R3792 GNDA.n2371 GNDA.n2370 13.8005
R3793 GNDA.n2359 GNDA.n2358 13.8005
R3794 GNDA.n2509 GNDA.n2 13.8005
R3795 GNDA.n2326 GNDA.n2257 12.8807
R3796 GNDA.n2073 GNDA.n73 12.7542
R3797 GNDA.n835 GNDA.t209 12.3572
R3798 GNDA.n2101 GNDA.t185 12.3572
R3799 GNDA.t177 GNDA.n117 12.3572
R3800 GNDA.n2075 GNDA.n2074 12.2193
R3801 GNDA.t121 GNDA.t56 11.7135
R3802 GNDA.n591 GNDA.n184 11.6369
R3803 GNDA.n594 GNDA.n591 11.6369
R3804 GNDA.n595 GNDA.n594 11.6369
R3805 GNDA.n598 GNDA.n595 11.6369
R3806 GNDA.n599 GNDA.n598 11.6369
R3807 GNDA.n602 GNDA.n599 11.6369
R3808 GNDA.n603 GNDA.n602 11.6369
R3809 GNDA.n606 GNDA.n603 11.6369
R3810 GNDA.n608 GNDA.n606 11.6369
R3811 GNDA.n609 GNDA.n608 11.6369
R3812 GNDA.n886 GNDA.n797 11.6369
R3813 GNDA.n891 GNDA.n886 11.6369
R3814 GNDA.n892 GNDA.n891 11.6369
R3815 GNDA.n893 GNDA.n892 11.6369
R3816 GNDA.n893 GNDA.n884 11.6369
R3817 GNDA.n899 GNDA.n884 11.6369
R3818 GNDA.n900 GNDA.n899 11.6369
R3819 GNDA.n901 GNDA.n900 11.6369
R3820 GNDA.n901 GNDA.n882 11.6369
R3821 GNDA.n907 GNDA.n882 11.6369
R3822 GNDA.n908 GNDA.n907 11.6369
R3823 GNDA.n1255 GNDA.n1254 11.6369
R3824 GNDA.n1254 GNDA.n1253 11.6369
R3825 GNDA.n1253 GNDA.n1251 11.6369
R3826 GNDA.n1251 GNDA.n1248 11.6369
R3827 GNDA.n1248 GNDA.n1247 11.6369
R3828 GNDA.n1247 GNDA.n1244 11.6369
R3829 GNDA.n1244 GNDA.n1243 11.6369
R3830 GNDA.n1243 GNDA.n1240 11.6369
R3831 GNDA.n1240 GNDA.n1239 11.6369
R3832 GNDA.n1239 GNDA.n1237 11.6369
R3833 GNDA.n771 GNDA.n770 11.6369
R3834 GNDA.n774 GNDA.n771 11.6369
R3835 GNDA.n775 GNDA.n774 11.6369
R3836 GNDA.n778 GNDA.n775 11.6369
R3837 GNDA.n779 GNDA.n778 11.6369
R3838 GNDA.n782 GNDA.n779 11.6369
R3839 GNDA.n784 GNDA.n782 11.6369
R3840 GNDA.n785 GNDA.n784 11.6369
R3841 GNDA.n786 GNDA.n785 11.6369
R3842 GNDA.n786 GNDA.n582 11.6369
R3843 GNDA.n765 GNDA.n740 11.6369
R3844 GNDA.n765 GNDA.n764 11.6369
R3845 GNDA.n764 GNDA.n763 11.6369
R3846 GNDA.n763 GNDA.n742 11.6369
R3847 GNDA.n758 GNDA.n742 11.6369
R3848 GNDA.n758 GNDA.n757 11.6369
R3849 GNDA.n757 GNDA.n756 11.6369
R3850 GNDA.n756 GNDA.n745 11.6369
R3851 GNDA.n751 GNDA.n745 11.6369
R3852 GNDA.n751 GNDA.n750 11.6369
R3853 GNDA.n750 GNDA.n479 11.6369
R3854 GNDA.n566 GNDA.n561 11.6369
R3855 GNDA.n1639 GNDA.n566 11.6369
R3856 GNDA.n1639 GNDA.n1638 11.6369
R3857 GNDA.n1638 GNDA.n1637 11.6369
R3858 GNDA.n1637 GNDA.n567 11.6369
R3859 GNDA.n1632 GNDA.n567 11.6369
R3860 GNDA.n1632 GNDA.n1631 11.6369
R3861 GNDA.n1631 GNDA.n1630 11.6369
R3862 GNDA.n1630 GNDA.n569 11.6369
R3863 GNDA.n1624 GNDA.n569 11.6369
R3864 GNDA.n1662 GNDA.n553 11.6369
R3865 GNDA.n1662 GNDA.n1661 11.6369
R3866 GNDA.n1661 GNDA.n1660 11.6369
R3867 GNDA.n1660 GNDA.n555 11.6369
R3868 GNDA.n1655 GNDA.n555 11.6369
R3869 GNDA.n1655 GNDA.n1654 11.6369
R3870 GNDA.n1654 GNDA.n1653 11.6369
R3871 GNDA.n1653 GNDA.n558 11.6369
R3872 GNDA.n1648 GNDA.n558 11.6369
R3873 GNDA.n1648 GNDA.n1647 11.6369
R3874 GNDA.n1647 GNDA.n1646 11.6369
R3875 GNDA.n529 GNDA.n480 11.6369
R3876 GNDA.n534 GNDA.n529 11.6369
R3877 GNDA.n535 GNDA.n534 11.6369
R3878 GNDA.n536 GNDA.n535 11.6369
R3879 GNDA.n536 GNDA.n527 11.6369
R3880 GNDA.n542 GNDA.n527 11.6369
R3881 GNDA.n543 GNDA.n542 11.6369
R3882 GNDA.n544 GNDA.n543 11.6369
R3883 GNDA.n544 GNDA.n525 11.6369
R3884 GNDA.n550 GNDA.n525 11.6369
R3885 GNDA.n551 GNDA.n550 11.6369
R3886 GNDA.n1878 GNDA.n1877 11.6369
R3887 GNDA.n1877 GNDA.n1876 11.6369
R3888 GNDA.n1876 GNDA.n224 11.6369
R3889 GNDA.n1870 GNDA.n224 11.6369
R3890 GNDA.n1870 GNDA.n1869 11.6369
R3891 GNDA.n1869 GNDA.n1868 11.6369
R3892 GNDA.n1868 GNDA.n228 11.6369
R3893 GNDA.n1862 GNDA.n228 11.6369
R3894 GNDA.n1862 GNDA.n1861 11.6369
R3895 GNDA.n1861 GNDA.n1860 11.6369
R3896 GNDA.n1860 GNDA.n232 11.6369
R3897 GNDA.n1854 GNDA.n1853 11.6369
R3898 GNDA.n1853 GNDA.n1852 11.6369
R3899 GNDA.n1852 GNDA.n236 11.6369
R3900 GNDA.n1846 GNDA.n236 11.6369
R3901 GNDA.n1846 GNDA.n1845 11.6369
R3902 GNDA.n1845 GNDA.n1844 11.6369
R3903 GNDA.n1844 GNDA.n239 11.6369
R3904 GNDA.n243 GNDA.n239 11.6369
R3905 GNDA.n1837 GNDA.n243 11.6369
R3906 GNDA.n1837 GNDA.n1836 11.6369
R3907 GNDA.n1940 GNDA.n1939 11.6369
R3908 GNDA.n1942 GNDA.n1940 11.6369
R3909 GNDA.n1942 GNDA.n1941 11.6369
R3910 GNDA.n1941 GNDA.n137 11.6369
R3911 GNDA.n137 GNDA.n135 11.6369
R3912 GNDA.n1950 GNDA.n135 11.6369
R3913 GNDA.n1951 GNDA.n1950 11.6369
R3914 GNDA.n1953 GNDA.n1951 11.6369
R3915 GNDA.n1953 GNDA.n1952 11.6369
R3916 GNDA.n1952 GNDA.n132 11.6369
R3917 GNDA.n1084 GNDA.n1060 11.6369
R3918 GNDA.n1084 GNDA.n1083 11.6369
R3919 GNDA.n1083 GNDA.n1082 11.6369
R3920 GNDA.n1082 GNDA.n1062 11.6369
R3921 GNDA.n1077 GNDA.n1062 11.6369
R3922 GNDA.n1077 GNDA.n1076 11.6369
R3923 GNDA.n1076 GNDA.n1075 11.6369
R3924 GNDA.n1075 GNDA.n1065 11.6369
R3925 GNDA.n1070 GNDA.n1065 11.6369
R3926 GNDA.n1070 GNDA.n1069 11.6369
R3927 GNDA.n1069 GNDA.n140 11.6369
R3928 GNDA.n1112 GNDA.n910 11.6369
R3929 GNDA.n1112 GNDA.n1111 11.6369
R3930 GNDA.n1111 GNDA.n1110 11.6369
R3931 GNDA.n1110 GNDA.n912 11.6369
R3932 GNDA.n1105 GNDA.n912 11.6369
R3933 GNDA.n1105 GNDA.n1104 11.6369
R3934 GNDA.n1104 GNDA.n1103 11.6369
R3935 GNDA.n1103 GNDA.n915 11.6369
R3936 GNDA.n1098 GNDA.n915 11.6369
R3937 GNDA.n1098 GNDA.n1097 11.6369
R3938 GNDA.n1097 GNDA.n1096 11.6369
R3939 GNDA.n1904 GNDA.n1903 11.6369
R3940 GNDA.n1903 GNDA.n1902 11.6369
R3941 GNDA.n1902 GNDA.n200 11.6369
R3942 GNDA.n1896 GNDA.n200 11.6369
R3943 GNDA.n1896 GNDA.n1895 11.6369
R3944 GNDA.n1893 GNDA.n206 11.6369
R3945 GNDA.n1887 GNDA.n206 11.6369
R3946 GNDA.n1887 GNDA.n1886 11.6369
R3947 GNDA.n1886 GNDA.n1885 11.6369
R3948 GNDA.n1885 GNDA.n217 11.6369
R3949 GNDA.n1934 GNDA.n1933 11.6369
R3950 GNDA.n1933 GNDA.n1932 11.6369
R3951 GNDA.n1932 GNDA.n185 11.6369
R3952 GNDA.n1926 GNDA.n185 11.6369
R3953 GNDA.n1926 GNDA.n1925 11.6369
R3954 GNDA.n1925 GNDA.n1924 11.6369
R3955 GNDA.n1924 GNDA.n189 11.6369
R3956 GNDA.n1918 GNDA.n189 11.6369
R3957 GNDA.n1918 GNDA.n1917 11.6369
R3958 GNDA.n1917 GNDA.n1916 11.6369
R3959 GNDA.n1916 GNDA.n193 11.6369
R3960 GNDA.n2272 GNDA.t28 11.5188
R3961 GNDA.n2282 GNDA.t21 11.5188
R3962 GNDA.n1968 GNDA.n1967 11.3792
R3963 GNDA.n2554 GNDA.n2553 10.2036
R3964 GNDA.n2553 GNDA.n14 10.0943
R3965 GNDA.n127 GNDA.n0 9.75668
R3966 GNDA.n168 GNDA.t318 9.6005
R3967 GNDA.n162 GNDA.t322 9.6005
R3968 GNDA.n2064 GNDA.t316 9.6005
R3969 GNDA.n75 GNDA.t319 9.6005
R3970 GNDA.n2312 GNDA.t287 9.6005
R3971 GNDA.n2306 GNDA.t1 9.6005
R3972 GNDA.n2306 GNDA.t331 9.6005
R3973 GNDA.n2304 GNDA.t164 9.6005
R3974 GNDA.n2304 GNDA.t176 9.6005
R3975 GNDA.n2302 GNDA.t153 9.6005
R3976 GNDA.n2302 GNDA.t168 9.6005
R3977 GNDA.n2300 GNDA.t46 9.6005
R3978 GNDA.n2300 GNDA.t166 9.6005
R3979 GNDA.n2298 GNDA.t8 9.6005
R3980 GNDA.n2298 GNDA.t124 9.6005
R3981 GNDA.n2296 GNDA.t84 9.6005
R3982 GNDA.n2296 GNDA.t356 9.6005
R3983 GNDA.n2294 GNDA.t29 9.6005
R3984 GNDA.n2294 GNDA.t144 9.6005
R3985 GNDA.n2292 GNDA.t172 9.6005
R3986 GNDA.n2292 GNDA.t337 9.6005
R3987 GNDA.n2290 GNDA.t156 9.6005
R3988 GNDA.n2290 GNDA.t326 9.6005
R3989 GNDA.n2288 GNDA.t148 9.6005
R3990 GNDA.n2288 GNDA.t174 9.6005
R3991 GNDA.n2286 GNDA.t48 9.6005
R3992 GNDA.n2286 GNDA.t311 9.6005
R3993 GNDA.n2275 GNDA.t312 9.6005
R3994 GNDA.t221 GNDA.t44 9.37093
R3995 GNDA.n2213 GNDA.n2130 9.14336
R3996 GNDA.n2213 GNDA.n2212 9.14336
R3997 GNDA.n2212 GNDA.n2210 9.14336
R3998 GNDA.n2210 GNDA.n2207 9.14336
R3999 GNDA.n2207 GNDA.n2206 9.14336
R4000 GNDA.n2206 GNDA.n2203 9.14336
R4001 GNDA.n2203 GNDA.n2202 9.14336
R4002 GNDA.n2202 GNDA.n2199 9.14336
R4003 GNDA.n2199 GNDA.n2198 9.14336
R4004 GNDA.n2198 GNDA.n2195 9.14336
R4005 GNDA.n2195 GNDA.n2194 9.14336
R4006 GNDA.n2317 GNDA.n2316 9.14336
R4007 GNDA.n2314 GNDA.n2313 9.14336
R4008 GNDA.n2280 GNDA.n2279 9.14336
R4009 GNDA.n2277 GNDA.n2276 9.14336
R4010 GNDA.n2225 GNDA.n2223 9.14336
R4011 GNDA.n2405 GNDA.n2400 9.14336
R4012 GNDA.n2405 GNDA.n2404 9.14336
R4013 GNDA.n2404 GNDA.n2402 9.14336
R4014 GNDA.n2421 GNDA.n2117 9.14336
R4015 GNDA.n2421 GNDA.n2420 9.14336
R4016 GNDA.n2420 GNDA.n2418 9.14336
R4017 GNDA.n2332 GNDA.n2331 9.14336
R4018 GNDA.n2342 GNDA.n2341 9.14336
R4019 GNDA.n2375 GNDA.n2374 9.14336
R4020 GNDA.n2364 GNDA.n2363 9.14336
R4021 GNDA.n2544 GNDA.n2539 9.14336
R4022 GNDA.n2544 GNDA.n2543 9.14336
R4023 GNDA.n2543 GNDA.n2541 9.14336
R4024 GNDA.n2448 GNDA.n2440 9.14336
R4025 GNDA.n2448 GNDA.n2447 9.14336
R4026 GNDA.n2447 GNDA.n2445 9.14336
R4027 GNDA.n2532 GNDA.n2499 9.14336
R4028 GNDA.n2532 GNDA.n2531 9.14336
R4029 GNDA.n2531 GNDA.n2529 9.14336
R4030 GNDA.n2529 GNDA.n2526 9.14336
R4031 GNDA.n2526 GNDA.n2525 9.14336
R4032 GNDA.n2525 GNDA.n2522 9.14336
R4033 GNDA.n2522 GNDA.n2521 9.14336
R4034 GNDA.n2521 GNDA.n2518 9.14336
R4035 GNDA.n2518 GNDA.n2517 9.14336
R4036 GNDA.n2517 GNDA.n2514 9.14336
R4037 GNDA.n2514 GNDA.n2513 9.14336
R4038 GNDA.n2492 GNDA.n2455 9.14336
R4039 GNDA.n2492 GNDA.n2491 9.14336
R4040 GNDA.n2491 GNDA.n2489 9.14336
R4041 GNDA.n2489 GNDA.n2486 9.14336
R4042 GNDA.n2486 GNDA.n2485 9.14336
R4043 GNDA.n2485 GNDA.n2482 9.14336
R4044 GNDA.n2482 GNDA.n2481 9.14336
R4045 GNDA.n2481 GNDA.n2478 9.14336
R4046 GNDA.n2478 GNDA.n2477 9.14336
R4047 GNDA.n2477 GNDA.n2474 9.14336
R4048 GNDA.n2474 GNDA.n2473 9.14336
R4049 GNDA.n2154 GNDA.n2151 9.14336
R4050 GNDA.n2158 GNDA.n2151 9.14336
R4051 GNDA.n2158 GNDA.n2149 9.14336
R4052 GNDA.n2164 GNDA.n2149 9.14336
R4053 GNDA.n2164 GNDA.n2147 9.14336
R4054 GNDA.n2168 GNDA.n2147 9.14336
R4055 GNDA.n2168 GNDA.n2145 9.14336
R4056 GNDA.n2174 GNDA.n2145 9.14336
R4057 GNDA.n2174 GNDA.n2143 9.14336
R4058 GNDA.n2178 GNDA.n2143 9.14336
R4059 GNDA.n2178 GNDA.n2141 9.14336
R4060 GNDA.n1704 GNDA.n154 8.60107
R4061 GNDA.n322 GNDA.n179 8.60107
R4062 GNDA.n2395 GNDA.n2394 8.53383
R4063 GNDA.n834 GNDA.t181 8.23827
R4064 GNDA.t195 GNDA.n2078 8.23827
R4065 GNDA.t189 GNDA.n2059 8.23827
R4066 GNDA.n1963 GNDA.n108 8.19962
R4067 GNDA.t304 GNDA.t7 7.67938
R4068 GNDA.t146 GNDA.t123 7.67938
R4069 GNDA.t131 GNDA.n2378 7.67938
R4070 GNDA.t83 GNDA.t52 7.67938
R4071 GNDA.t355 GNDA.t266 7.67938
R4072 GNDA.n72 GNDA.n71 7.56675
R4073 GNDA.n209 GNDA.n127 7.56675
R4074 GNDA.n852 GNDA.t154 7.20855
R4075 GNDA.n2036 GNDA.t13 7.20855
R4076 GNDA.t135 GNDA.n124 7.20855
R4077 GNDA.n1972 GNDA.n1971 7.20855
R4078 GNDA.n2324 GNDA.n2323 7.03175
R4079 GNDA.n2324 GNDA.n1 6.8755
R4080 GNDA.n909 GNDA.n908 6.72373
R4081 GNDA.n1730 GNDA.n479 6.72373
R4082 GNDA.n552 GNDA.n551 6.72373
R4083 GNDA.n1096 GNDA.n918 6.72373
R4084 GNDA.n223 GNDA.n217 6.72373
R4085 GNDA.n199 GNDA.n193 6.72373
R4086 GNDA.n14 GNDA.n13 6.39112
R4087 GNDA.n2555 GNDA.n2554 6.28175
R4088 GNDA.n2555 GNDA.n1 6.28175
R4089 GNDA.n553 GNDA.n552 6.20656
R4090 GNDA.n1730 GNDA.n480 6.20656
R4091 GNDA.n1878 GNDA.n223 6.20656
R4092 GNDA.n1060 GNDA.n918 6.20656
R4093 GNDA.n910 GNDA.n909 6.20656
R4094 GNDA.n1904 GNDA.n199 6.20656
R4095 GNDA.t335 GNDA.t221 6.17883
R4096 GNDA.n1895 GNDA.n1894 6.07727
R4097 GNDA.n171 GNDA.n70 5.81868
R4098 GNDA.n171 GNDA.n170 5.81868
R4099 GNDA.n2192 GNDA.n2191 5.78934
R4100 GNDA.n2411 GNDA.n2120 5.78934
R4101 GNDA.n2416 GNDA.n2415 5.78934
R4102 GNDA.n2550 GNDA.n16 5.78934
R4103 GNDA.n2443 GNDA.n2442 5.78934
R4104 GNDA.n2511 GNDA.n2510 5.78934
R4105 GNDA.n2471 GNDA.n2470 5.78934
R4106 GNDA.n2183 GNDA.n2140 5.78934
R4107 GNDA.n72 GNDA.n0 5.737
R4108 GNDA.n1894 GNDA.n1893 5.5601
R4109 GNDA.n2553 GNDA.n2552 5.54068
R4110 GNDA.n670 GNDA.n634 5.51161
R4111 GNDA.n1171 GNDA.n823 5.51161
R4112 GNDA.n1311 GNDA.n1289 5.51161
R4113 GNDA.n1485 GNDA.n1455 5.51161
R4114 GNDA.n1616 GNDA.n1615 5.51161
R4115 GNDA.n1774 GNDA.n1773 5.51161
R4116 GNDA.n1825 GNDA.n1824 5.51161
R4117 GNDA.n1013 GNDA.n997 5.51161
R4118 GNDA.n1979 GNDA.n113 5.51161
R4119 GNDA.n2327 GNDA.n2326 5.46925
R4120 GNDA.n1623 GNDA.n574 5.1717
R4121 GNDA.n1835 GNDA.n244 5.1717
R4122 GNDA.n130 GNDA.n129 5.1717
R4123 GNDA.n2102 GNDA.t221 5.14911
R4124 GNDA.t66 GNDA.t278 5.14911
R4125 GNDA.n2257 GNDA.n2255 5.063
R4126 GNDA.n13 GNDA.n11 5.063
R4127 GNDA.n731 GNDA.n610 4.9157
R4128 GNDA.n1236 GNDA.n799 4.9157
R4129 GNDA.n1375 GNDA.n1261 4.9157
R4130 GNDA.n2325 GNDA.n2119 4.5005
R4131 GNDA.n2316 GNDA.n2315 4.46219
R4132 GNDA.n2313 GNDA.n2308 4.46219
R4133 GNDA.n2315 GNDA.n2314 4.46219
R4134 GNDA.n2321 GNDA.n2308 4.46219
R4135 GNDA.n2279 GNDA.n2278 4.46219
R4136 GNDA.n2276 GNDA.n2258 4.46219
R4137 GNDA.n2278 GNDA.n2277 4.46219
R4138 GNDA.n2284 GNDA.n2258 4.46219
R4139 GNDA.n2223 GNDA.n2222 4.46219
R4140 GNDA.n2229 GNDA.n2222 4.46219
R4141 GNDA.n2331 GNDA.n2330 4.46219
R4142 GNDA.n2330 GNDA.n2329 4.46219
R4143 GNDA.n2341 GNDA.n2340 4.46219
R4144 GNDA.n2340 GNDA.n2339 4.46219
R4145 GNDA.n2374 GNDA.n2373 4.46219
R4146 GNDA.n2373 GNDA.n2372 4.46219
R4147 GNDA.n2363 GNDA.n2242 4.46219
R4148 GNDA.n2368 GNDA.n2242 4.46219
R4149 GNDA.n337 GNDA.n336 4.26717
R4150 GNDA.n344 GNDA.n336 4.26717
R4151 GNDA.n345 GNDA.n344 4.26717
R4152 GNDA.n345 GNDA.n332 4.26717
R4153 GNDA.n351 GNDA.n332 4.26717
R4154 GNDA.n352 GNDA.n351 4.26717
R4155 GNDA.n352 GNDA.n329 4.26717
R4156 GNDA.n358 GNDA.n329 4.26717
R4157 GNDA.n359 GNDA.n358 4.26717
R4158 GNDA.n359 GNDA.n325 4.26717
R4159 GNDA.n1781 GNDA.n325 4.26717
R4160 GNDA.n1091 GNDA.n920 4.26717
R4161 GNDA.n1091 GNDA.n923 4.26717
R4162 GNDA.n1056 GNDA.n923 4.26717
R4163 GNDA.n1056 GNDA.n1055 4.26717
R4164 GNDA.n1055 GNDA.n1054 4.26717
R4165 GNDA.n1054 GNDA.n930 4.26717
R4166 GNDA.n1048 GNDA.n930 4.26717
R4167 GNDA.n1048 GNDA.n1047 4.26717
R4168 GNDA.n1047 GNDA.n1046 4.26717
R4169 GNDA.n1046 GNDA.n938 4.26717
R4170 GNDA.n1040 GNDA.n938 4.26717
R4171 GNDA.n1668 GNDA.n523 4.26717
R4172 GNDA.n1674 GNDA.n523 4.26717
R4173 GNDA.n1674 GNDA.n521 4.26717
R4174 GNDA.n1680 GNDA.n521 4.26717
R4175 GNDA.n1680 GNDA.n519 4.26717
R4176 GNDA.n1686 GNDA.n519 4.26717
R4177 GNDA.n1686 GNDA.n517 4.26717
R4178 GNDA.n1692 GNDA.n517 4.26717
R4179 GNDA.n1692 GNDA.n515 4.26717
R4180 GNDA.n1699 GNDA.n515 4.26717
R4181 GNDA.n1699 GNDA.n513 4.26717
R4182 GNDA.n1909 GNDA.n194 4.26717
R4183 GNDA.n1909 GNDA.n196 4.26717
R4184 GNDA.n451 GNDA.n196 4.26717
R4185 GNDA.n456 GNDA.n451 4.26717
R4186 GNDA.n456 GNDA.n448 4.26717
R4187 GNDA.n462 GNDA.n448 4.26717
R4188 GNDA.n462 GNDA.n446 4.26717
R4189 GNDA.n469 GNDA.n446 4.26717
R4190 GNDA.n469 GNDA.n443 4.26717
R4191 GNDA.n475 GNDA.n443 4.26717
R4192 GNDA.n476 GNDA.n475 4.26717
R4193 GNDA.n1729 GNDA.n482 4.26717
R4194 GNDA.n1724 GNDA.n482 4.26717
R4195 GNDA.n1724 GNDA.n1723 4.26717
R4196 GNDA.n1723 GNDA.n490 4.26717
R4197 GNDA.n1718 GNDA.n490 4.26717
R4198 GNDA.n1718 GNDA.n1717 4.26717
R4199 GNDA.n1717 GNDA.n1716 4.26717
R4200 GNDA.n1716 GNDA.n498 4.26717
R4201 GNDA.n1710 GNDA.n498 4.26717
R4202 GNDA.n1710 GNDA.n1709 4.26717
R4203 GNDA.n1709 GNDA.n1708 4.26717
R4204 GNDA.n1118 GNDA.n880 4.26717
R4205 GNDA.n1124 GNDA.n880 4.26717
R4206 GNDA.n1124 GNDA.n878 4.26717
R4207 GNDA.n1130 GNDA.n878 4.26717
R4208 GNDA.n1130 GNDA.n876 4.26717
R4209 GNDA.n1136 GNDA.n876 4.26717
R4210 GNDA.n1136 GNDA.n874 4.26717
R4211 GNDA.n1142 GNDA.n874 4.26717
R4212 GNDA.n1142 GNDA.n872 4.26717
R4213 GNDA.n1150 GNDA.n872 4.26717
R4214 GNDA.n1150 GNDA.n869 4.26717
R4215 GNDA.n2390 GNDA.n2389 4.2505
R4216 GNDA GNDA.n2556 4.2117
R4217 GNDA.n2358 GNDA.n14 4.19842
R4218 GNDA.n2394 GNDA.n2393 4.17148
R4219 GNDA.n2393 GNDA.n2392 4.17148
R4220 GNDA.n2074 GNDA.n2073 4.063
R4221 GNDA.n2327 GNDA.n2241 4.0005
R4222 GNDA.n337 GNDA.n223 3.93531
R4223 GNDA.n920 GNDA.n918 3.93531
R4224 GNDA.n1668 GNDA.n552 3.93531
R4225 GNDA.n199 GNDA.n194 3.93531
R4226 GNDA.n1730 GNDA.n1729 3.93531
R4227 GNDA.n1118 GNDA.n909 3.93531
R4228 GNDA.t90 GNDA.t295 3.83994
R4229 GNDA.t272 GNDA.t145 3.83994
R4230 GNDA.t261 GNDA.t138 3.83994
R4231 GNDA.t92 GNDA.t251 3.83994
R4232 GNDA.n729 GNDA.n613 3.7893
R4233 GNDA.n726 GNDA.n725 3.7893
R4234 GNDA.n639 GNDA.n615 3.7893
R4235 GNDA.n642 GNDA.n641 3.7893
R4236 GNDA.n649 GNDA.n637 3.7893
R4237 GNDA.n654 GNDA.n653 3.7893
R4238 GNDA.n658 GNDA.n657 3.7893
R4239 GNDA.n667 GNDA.n635 3.7893
R4240 GNDA.n1221 GNDA.n802 3.7893
R4241 GNDA.n1229 GNDA.n1228 3.7893
R4242 GNDA.n830 GNDA.n803 3.7893
R4243 GNDA.n831 GNDA.n829 3.7893
R4244 GNDA.n839 GNDA.n837 3.7893
R4245 GNDA.n848 GNDA.n847 3.7893
R4246 GNDA.n844 GNDA.n843 3.7893
R4247 GNDA.n1168 GNDA.n824 3.7893
R4248 GNDA.n1373 GNDA.n1372 3.7893
R4249 GNDA.n1369 GNDA.n1264 3.7893
R4250 GNDA.n1368 GNDA.n1267 3.7893
R4251 GNDA.n1365 GNDA.n1364 3.7893
R4252 GNDA.n1291 GNDA.n1268 3.7893
R4253 GNDA.n1300 GNDA.n1299 3.7893
R4254 GNDA.n1303 GNDA.n1290 3.7893
R4255 GNDA.n1308 GNDA.n1304 3.7893
R4256 GNDA.n1535 GNDA.n1469 3.7893
R4257 GNDA.n1544 GNDA.n1543 3.7893
R4258 GNDA.n1466 GNDA.n1465 3.7893
R4259 GNDA.n1552 GNDA.n1550 3.7893
R4260 GNDA.n1551 GNDA.n1463 3.7893
R4261 GNDA.n1461 GNDA.n1460 3.7893
R4262 GNDA.n1566 GNDA.n1565 3.7893
R4263 GNDA.n1570 GNDA.n1457 3.7893
R4264 GNDA.n1578 GNDA.n1393 3.7893
R4265 GNDA.n1587 GNDA.n1586 3.7893
R4266 GNDA.n1390 GNDA.n1389 3.7893
R4267 GNDA.n1595 GNDA.n1593 3.7893
R4268 GNDA.n1594 GNDA.n1387 3.7893
R4269 GNDA.n1385 GNDA.n1384 3.7893
R4270 GNDA.n1610 GNDA.n1608 3.7893
R4271 GNDA.n1609 GNDA.n1380 3.7893
R4272 GNDA.n1787 GNDA.n259 3.7893
R4273 GNDA.n1796 GNDA.n1795 3.7893
R4274 GNDA.n257 GNDA.n256 3.7893
R4275 GNDA.n1804 GNDA.n1802 3.7893
R4276 GNDA.n1803 GNDA.n254 3.7893
R4277 GNDA.n252 GNDA.n251 3.7893
R4278 GNDA.n1819 GNDA.n1817 3.7893
R4279 GNDA.n1818 GNDA.n247 3.7893
R4280 GNDA.n1736 GNDA.n378 3.7893
R4281 GNDA.n1745 GNDA.n1744 3.7893
R4282 GNDA.n376 GNDA.n375 3.7893
R4283 GNDA.n1753 GNDA.n1751 3.7893
R4284 GNDA.n1752 GNDA.n373 3.7893
R4285 GNDA.n371 GNDA.n370 3.7893
R4286 GNDA.n1768 GNDA.n1766 3.7893
R4287 GNDA.n1767 GNDA.n366 3.7893
R4288 GNDA.n2093 GNDA.n65 3.7893
R4289 GNDA.n2092 GNDA.n66 3.7893
R4290 GNDA.n2080 GNDA.n2079 3.7893
R4291 GNDA.n2086 GNDA.n2085 3.7893
R4292 GNDA.n2082 GNDA.n2081 3.7893
R4293 GNDA.n1000 GNDA.n44 3.7893
R4294 GNDA.n1001 GNDA.n999 3.7893
R4295 GNDA.n1011 GNDA.n1008 3.7893
R4296 GNDA.n2051 GNDA.n104 3.7893
R4297 GNDA.n2050 GNDA.n105 3.7893
R4298 GNDA.n2038 GNDA.n2037 3.7893
R4299 GNDA.n2044 GNDA.n2043 3.7893
R4300 GNDA.n2040 GNDA.n2039 3.7893
R4301 GNDA.n118 GNDA.n83 3.7893
R4302 GNDA.n121 GNDA.n120 3.7893
R4303 GNDA.n1976 GNDA.n114 3.7893
R4304 GNDA.n652 GNDA 3.7381
R4305 GNDA.n842 GNDA 3.7381
R4306 GNDA.n1296 GNDA 3.7381
R4307 GNDA GNDA.n1558 3.7381
R4308 GNDA GNDA.n1601 3.7381
R4309 GNDA GNDA.n1810 3.7381
R4310 GNDA GNDA.n1759 3.7381
R4311 GNDA GNDA.n2098 3.7381
R4312 GNDA GNDA.n2056 3.7381
R4313 GNDA.n1967 GNDA.n127 3.51962
R4314 GNDA.n2326 GNDA.n2325 3.5005
R4315 GNDA.n2185 GNDA.t41 3.42907
R4316 GNDA.n2185 GNDA.t170 3.42907
R4317 GNDA.n2187 GNDA.t358 3.42907
R4318 GNDA.n2187 GNDA.t43 3.42907
R4319 GNDA.n2465 GNDA.t110 3.42907
R4320 GNDA.n2465 GNDA.t81 3.42907
R4321 GNDA.n2467 GNDA.t137 3.42907
R4322 GNDA.n2467 GNDA.t37 3.42907
R4323 GNDA.n2325 GNDA.n2324 3.20362
R4324 GNDA.n2215 GNDA.n2130 3.19754
R4325 GNDA.n2194 GNDA.n2192 3.19754
R4326 GNDA.n2407 GNDA.n2400 3.19754
R4327 GNDA.n2402 GNDA.n2120 3.19754
R4328 GNDA.n2423 GNDA.n2117 3.19754
R4329 GNDA.n2418 GNDA.n2416 3.19754
R4330 GNDA.n2546 GNDA.n2539 3.19754
R4331 GNDA.n2541 GNDA.n16 3.19754
R4332 GNDA.n2450 GNDA.n2440 3.19754
R4333 GNDA.n2445 GNDA.n2443 3.19754
R4334 GNDA.n2534 GNDA.n2499 3.19754
R4335 GNDA.n2513 GNDA.n2511 3.19754
R4336 GNDA.n2494 GNDA.n2455 3.19754
R4337 GNDA.n2473 GNDA.n2471 3.19754
R4338 GNDA.n2155 GNDA.n2154 3.19754
R4339 GNDA.n2141 GNDA.n2140 3.19754
R4340 GNDA.n1233 GNDA.n176 3.08966
R4341 GNDA.t122 GNDA.n1231 3.08966
R4342 GNDA.n826 GNDA.t102 3.08966
R4343 GNDA.n1165 GNDA.t60 3.08966
R4344 GNDA.n2048 GNDA.t351 3.08966
R4345 GNDA.n2066 GNDA.n74 2.86505
R4346 GNDA.n2067 GNDA.n2066 2.86505
R4347 GNDA.n2065 GNDA.n2061 2.86505
R4348 GNDA.n2062 GNDA.n2061 2.86505
R4349 GNDA.n2068 GNDA.n2067 2.86505
R4350 GNDA.n2063 GNDA.n2062 2.86505
R4351 GNDA.n2072 GNDA.n74 2.86505
R4352 GNDA.n2068 GNDA.n2065 2.86505
R4353 GNDA.n2380 GNDA.n2379 2.86505
R4354 GNDA.n2379 GNDA.n2233 2.86505
R4355 GNDA.n2386 GNDA.n2233 2.86505
R4356 GNDA.n2382 GNDA.n2380 2.86505
R4357 GNDA.n2263 GNDA.n2262 2.86505
R4358 GNDA.n2268 GNDA.n2263 2.86505
R4359 GNDA.n2268 GNDA.n2267 2.86505
R4360 GNDA.n2270 GNDA.n2262 2.86505
R4361 GNDA.n169 GNDA.n165 2.86505
R4362 GNDA.n166 GNDA.n165 2.86505
R4363 GNDA.n167 GNDA.n166 2.86505
R4364 GNDA.n170 GNDA.n169 2.86505
R4365 GNDA.n731 GNDA.n730 2.6629
R4366 GNDA.n662 GNDA.n440 2.6629
R4367 GNDA.n1222 GNDA.n799 2.6629
R4368 GNDA.n943 GNDA.n942 2.6629
R4369 GNDA.n1375 GNDA.n1374 2.6629
R4370 GNDA.n1288 GNDA.n506 2.6629
R4371 GNDA.n1536 GNDA.n1534 2.6629
R4372 GNDA.n1576 GNDA.n1575 2.6629
R4373 GNDA.n1579 GNDA.n1577 2.6629
R4374 GNDA.n1788 GNDA.n1786 2.6629
R4375 GNDA.n1737 GNDA.n1735 2.6629
R4376 GNDA.n364 GNDA.n321 2.6629
R4377 GNDA.n945 GNDA.n944 2.6629
R4378 GNDA.n1014 GNDA.n112 2.6629
R4379 GNDA.n2032 GNDA.n2031 2.6629
R4380 GNDA.n662 GNDA.n634 2.4581
R4381 GNDA.n942 GNDA.n823 2.4581
R4382 GNDA.n1289 GNDA.n1288 2.4581
R4383 GNDA.n1534 GNDA.n506 2.4581
R4384 GNDA.n1575 GNDA.n1455 2.4581
R4385 GNDA.n1577 GNDA.n1576 2.4581
R4386 GNDA.n1616 GNDA.n574 2.4581
R4387 GNDA.n1786 GNDA.n321 2.4581
R4388 GNDA.n1825 GNDA.n244 2.4581
R4389 GNDA.n1735 GNDA.n440 2.4581
R4390 GNDA.n1774 GNDA.n364 2.4581
R4391 GNDA.n944 GNDA.n943 2.4581
R4392 GNDA.n1014 GNDA.n1013 2.4581
R4393 GNDA.n2032 GNDA.n112 2.4581
R4394 GNDA.n129 GNDA.n113 2.4581
R4395 GNDA.n2370 GNDA.n2241 2.2505
R4396 GNDA.n1781 GNDA.n321 2.18124
R4397 GNDA.n1040 GNDA.n112 2.18124
R4398 GNDA.n1576 GNDA.n513 2.18124
R4399 GNDA.n476 GNDA.n440 2.18124
R4400 GNDA.n1708 GNDA.n506 2.18124
R4401 GNDA.n943 GNDA.n869 2.18124
R4402 GNDA.n666 GNDA.n634 2.1509
R4403 GNDA.n1167 GNDA.n823 2.1509
R4404 GNDA.n1307 GNDA.n1289 2.1509
R4405 GNDA.n1571 GNDA.n1455 2.1509
R4406 GNDA.n1617 GNDA.n1616 2.1509
R4407 GNDA.n1826 GNDA.n1825 2.1509
R4408 GNDA.n1775 GNDA.n1774 2.1509
R4409 GNDA.n1013 GNDA.n1012 2.1509
R4410 GNDA.n1975 GNDA.n113 2.1509
R4411 GNDA.n730 GNDA.n612 2.13383
R4412 GNDA.n1223 GNDA.n1222 2.13383
R4413 GNDA.n1374 GNDA.n1262 2.13383
R4414 GNDA.n1537 GNDA.n1536 2.13383
R4415 GNDA.n1580 GNDA.n1579 2.13383
R4416 GNDA.n1738 GNDA.n1737 2.13383
R4417 GNDA.n1789 GNDA.n1788 2.13383
R4418 GNDA.n946 GNDA.n945 2.13383
R4419 GNDA.n2031 GNDA.n2030 2.13383
R4420 GNDA.n73 GNDA 2.09787
R4421 GNDA.n323 GNDA.n321 2.08643
R4422 GNDA.n1016 GNDA.n112 2.08643
R4423 GNDA.n1576 GNDA.n511 2.08643
R4424 GNDA.n1731 GNDA.n440 2.08643
R4425 GNDA.n508 GNDA.n506 2.08643
R4426 GNDA.n943 GNDA.n867 2.08643
R4427 GNDA.n1165 GNDA.t282 2.05994
R4428 GNDA.n866 GNDA.t307 2.05994
R4429 GNDA.t255 GNDA.n1017 2.05994
R4430 GNDA.t278 GNDA.n2035 2.05994
R4431 GNDA.n730 GNDA.n729 1.9461
R4432 GNDA.n1222 GNDA.n1221 1.9461
R4433 GNDA.n1374 GNDA.n1373 1.9461
R4434 GNDA.n1536 GNDA.n1535 1.9461
R4435 GNDA.n1579 GNDA.n1578 1.9461
R4436 GNDA.n1788 GNDA.n1787 1.9461
R4437 GNDA.n1737 GNDA.n1736 1.9461
R4438 GNDA.n945 GNDA.n65 1.9461
R4439 GNDA.n2031 GNDA.n104 1.9461
R4440 GNDA.n210 GNDA.n209 1.90675
R4441 GNDA.n142 GNDA.t317 1.83728
R4442 GNDA.n2389 GNDA.n2231 1.7505
R4443 GNDA.n610 GNDA.n609 1.47392
R4444 GNDA.n1237 GNDA.n1236 1.47392
R4445 GNDA.n1261 GNDA.n582 1.47392
R4446 GNDA.n1624 GNDA.n1623 1.47392
R4447 GNDA.n1836 GNDA.n1835 1.47392
R4448 GNDA.n132 GNDA.n130 1.47392
R4449 GNDA.n2554 GNDA.n2 1.28175
R4450 GNDA.n2189 GNDA.n1 1.28175
R4451 GNDA.n2468 GNDA.n2466 1.1255
R4452 GNDA.n2466 GNDA.n2 1.1255
R4453 GNDA.n2189 GNDA.n2188 1.1255
R4454 GNDA.n2188 GNDA.n2186 1.1255
R4455 GNDA.n2413 GNDA.n2119 1.04068
R4456 GNDA.n2390 GNDA.n2119 0.978179
R4457 GNDA.n1033 GNDA.n1032 0.96925
R4458 GNDA.n1160 GNDA.n1159 0.96925
R4459 GNDA.n726 GNDA.n613 0.8197
R4460 GNDA.n725 GNDA.n615 0.8197
R4461 GNDA.n642 GNDA.n639 0.8197
R4462 GNDA.n641 GNDA.n637 0.8197
R4463 GNDA.n653 GNDA.n652 0.8197
R4464 GNDA.n658 GNDA.n654 0.8197
R4465 GNDA.n657 GNDA.n635 0.8197
R4466 GNDA.n667 GNDA.n666 0.8197
R4467 GNDA.n1229 GNDA.n802 0.8197
R4468 GNDA.n1228 GNDA.n803 0.8197
R4469 GNDA.n831 GNDA.n830 0.8197
R4470 GNDA.n837 GNDA.n829 0.8197
R4471 GNDA.n848 GNDA.n842 0.8197
R4472 GNDA.n847 GNDA.n843 0.8197
R4473 GNDA.n844 GNDA.n824 0.8197
R4474 GNDA.n1168 GNDA.n1167 0.8197
R4475 GNDA.n1372 GNDA.n1264 0.8197
R4476 GNDA.n1369 GNDA.n1368 0.8197
R4477 GNDA.n1365 GNDA.n1267 0.8197
R4478 GNDA.n1364 GNDA.n1268 0.8197
R4479 GNDA.n1299 GNDA.n1296 0.8197
R4480 GNDA.n1300 GNDA.n1290 0.8197
R4481 GNDA.n1304 GNDA.n1303 0.8197
R4482 GNDA.n1308 GNDA.n1307 0.8197
R4483 GNDA.n1544 GNDA.n1469 0.8197
R4484 GNDA.n1543 GNDA.n1466 0.8197
R4485 GNDA.n1550 GNDA.n1465 0.8197
R4486 GNDA.n1552 GNDA.n1551 0.8197
R4487 GNDA.n1558 GNDA.n1461 0.8197
R4488 GNDA.n1565 GNDA.n1460 0.8197
R4489 GNDA.n1566 GNDA.n1457 0.8197
R4490 GNDA.n1571 GNDA.n1570 0.8197
R4491 GNDA.n1587 GNDA.n1393 0.8197
R4492 GNDA.n1586 GNDA.n1390 0.8197
R4493 GNDA.n1593 GNDA.n1389 0.8197
R4494 GNDA.n1595 GNDA.n1594 0.8197
R4495 GNDA.n1601 GNDA.n1385 0.8197
R4496 GNDA.n1608 GNDA.n1384 0.8197
R4497 GNDA.n1610 GNDA.n1609 0.8197
R4498 GNDA.n1617 GNDA.n1380 0.8197
R4499 GNDA.n1796 GNDA.n259 0.8197
R4500 GNDA.n1795 GNDA.n257 0.8197
R4501 GNDA.n1802 GNDA.n256 0.8197
R4502 GNDA.n1804 GNDA.n1803 0.8197
R4503 GNDA.n1810 GNDA.n252 0.8197
R4504 GNDA.n1817 GNDA.n251 0.8197
R4505 GNDA.n1819 GNDA.n1818 0.8197
R4506 GNDA.n1826 GNDA.n247 0.8197
R4507 GNDA.n1745 GNDA.n378 0.8197
R4508 GNDA.n1744 GNDA.n376 0.8197
R4509 GNDA.n1751 GNDA.n375 0.8197
R4510 GNDA.n1753 GNDA.n1752 0.8197
R4511 GNDA.n1759 GNDA.n371 0.8197
R4512 GNDA.n1766 GNDA.n370 0.8197
R4513 GNDA.n1768 GNDA.n1767 0.8197
R4514 GNDA.n1775 GNDA.n366 0.8197
R4515 GNDA.n2093 GNDA.n2092 0.8197
R4516 GNDA.n2079 GNDA.n66 0.8197
R4517 GNDA.n2086 GNDA.n2080 0.8197
R4518 GNDA.n2085 GNDA.n2082 0.8197
R4519 GNDA.n2098 GNDA.n44 0.8197
R4520 GNDA.n1001 GNDA.n1000 0.8197
R4521 GNDA.n1008 GNDA.n999 0.8197
R4522 GNDA.n1012 GNDA.n1011 0.8197
R4523 GNDA.n2051 GNDA.n2050 0.8197
R4524 GNDA.n2037 GNDA.n105 0.8197
R4525 GNDA.n2044 GNDA.n2038 0.8197
R4526 GNDA.n2043 GNDA.n2040 0.8197
R4527 GNDA.n2056 GNDA.n83 0.8197
R4528 GNDA.n121 GNDA.n118 0.8197
R4529 GNDA.n120 GNDA.n114 0.8197
R4530 GNDA.n1976 GNDA.n1975 0.8197
R4531 GNDA.t221 GNDA.t56 0.586152
R4532 GNDA.n1258 GNDA.n142 0.575776
R4533 GNDA.n649 GNDA 0.5637
R4534 GNDA.n839 GNDA 0.5637
R4535 GNDA GNDA.n1291 0.5637
R4536 GNDA.n1463 GNDA 0.5637
R4537 GNDA.n1387 GNDA 0.5637
R4538 GNDA.n254 GNDA 0.5637
R4539 GNDA.n373 GNDA 0.5637
R4540 GNDA.n2081 GNDA 0.5637
R4541 GNDA.n2039 GNDA 0.5637
R4542 GNDA.n1968 GNDA.n126 0.563
R4543 GNDA.n1025 GNDA.n126 0.563
R4544 GNDA.n1027 GNDA.n1025 0.563
R4545 GNDA.n1032 GNDA.n1027 0.563
R4546 GNDA.n1033 GNDA.n1023 0.563
R4547 GNDA.n1023 GNDA.n1021 0.563
R4548 GNDA.n1021 GNDA.n1019 0.563
R4549 GNDA.n1019 GNDA.n865 0.563
R4550 GNDA.n1159 GNDA.n865 0.563
R4551 GNDA.n1160 GNDA.n863 0.563
R4552 GNDA.n863 GNDA.n861 0.563
R4553 GNDA.n861 GNDA.n859 0.563
R4554 GNDA.n2289 GNDA.n2287 0.563
R4555 GNDA.n2291 GNDA.n2289 0.563
R4556 GNDA.n2293 GNDA.n2291 0.563
R4557 GNDA.n2295 GNDA.n2293 0.563
R4558 GNDA.n2297 GNDA.n2295 0.563
R4559 GNDA.n2299 GNDA.n2297 0.563
R4560 GNDA.n2301 GNDA.n2299 0.563
R4561 GNDA.n2303 GNDA.n2301 0.563
R4562 GNDA.n2305 GNDA.n2303 0.563
R4563 GNDA.n2307 GNDA.n2305 0.563
R4564 GNDA.n2323 GNDA.n2307 0.563
R4565 GNDA.n2251 GNDA.n2249 0.563
R4566 GNDA.n2253 GNDA.n2251 0.563
R4567 GNDA.n2255 GNDA.n2253 0.563
R4568 GNDA.n7 GNDA.n5 0.563
R4569 GNDA.n9 GNDA.n7 0.563
R4570 GNDA.n11 GNDA.n9 0.563
R4571 GNDA.n2351 GNDA.n2349 0.563
R4572 GNDA.n2353 GNDA.n2351 0.563
R4573 GNDA.n2355 GNDA.n2353 0.563
R4574 GNDA.n2357 GNDA.n2355 0.563
R4575 GNDA.n2358 GNDA.n2357 0.563
R4576 GNDA.n1966 GNDA.n73 0.276625
R4577 GNDA GNDA.n648 0.2565
R4578 GNDA GNDA.n838 0.2565
R4579 GNDA.n1294 GNDA 0.2565
R4580 GNDA.n1559 GNDA 0.2565
R4581 GNDA.n1602 GNDA 0.2565
R4582 GNDA.n1811 GNDA 0.2565
R4583 GNDA.n1760 GNDA 0.2565
R4584 GNDA.n2099 GNDA 0.2565
R4585 GNDA.n2057 GNDA 0.2565
R4586 GNDA.n1967 GNDA.n1966 0.22375
R4587 GNDA.n648 GNDA 0.0517
R4588 GNDA.n838 GNDA 0.0517
R4589 GNDA GNDA.n1294 0.0517
R4590 GNDA.n1559 GNDA 0.0517
R4591 GNDA.n1602 GNDA 0.0517
R4592 GNDA.n1811 GNDA 0.0517
R4593 GNDA.n1760 GNDA 0.0517
R4594 GNDA.n2099 GNDA 0.0517
R4595 GNDA.n2057 GNDA 0.0517
R4596 VDDA.n322 VDDA.t325 1212.4
R4597 VDDA.n386 VDDA.t316 1212.4
R4598 VDDA.n109 VDDA.t341 1212.4
R4599 VDDA.n178 VDDA.t356 1212.4
R4600 VDDA.n203 VDDA.t402 1095.3
R4601 VDDA.t396 VDDA.n202 1095.3
R4602 VDDA.t369 VDDA.n295 1093.7
R4603 VDDA.t311 VDDA.n86 1093.7
R4604 VDDA.n296 VDDA.t387 1082.5
R4605 VDDA.n88 VDDA.t302 1082.5
R4606 VDDA.n395 VDDA.t330 905.125
R4607 VDDA.n394 VDDA.t340 905.125
R4608 VDDA.n503 VDDA.t373 708.125
R4609 VDDA.t373 VDDA.n459 708.125
R4610 VDDA.n480 VDDA.t315 708.125
R4611 VDDA.t315 VDDA.n462 708.125
R4612 VDDA.n392 VDDA.n391 682
R4613 VDDA.n525 VDDA.t411 676.966
R4614 VDDA.n395 VDDA.t329 672.274
R4615 VDDA.t338 VDDA.n394 672.274
R4616 VDDA.n295 VDDA.t370 665.4
R4617 VDDA.n294 VDDA.t388 665.4
R4618 VDDA.n87 VDDA.t303 665.4
R4619 VDDA.n86 VDDA.t312 665.4
R4620 VDDA.n203 VDDA.t403 663.801
R4621 VDDA.n202 VDDA.t397 663.801
R4622 VDDA.n482 VDDA.t335 660.001
R4623 VDDA.t372 VDDA.n504 657.76
R4624 VDDA.t314 VDDA.n481 657.76
R4625 VDDA.n407 VDDA.t359 652.076
R4626 VDDA.n441 VDDA.t380 652.076
R4627 VDDA.n219 VDDA.t322 652.076
R4628 VDDA.n252 VDDA.t398 652.076
R4629 VDDA.n11 VDDA.t353 652.076
R4630 VDDA.n44 VDDA.t307 652.076
R4631 VDDA.t405 VDDA.n602 645.231
R4632 VDDA.n603 VDDA.t375 645.231
R4633 VDDA.t348 VDDA.n571 643.038
R4634 VDDA.t366 VDDA.n524 643.038
R4635 VDDA.n572 VDDA.t345 643.038
R4636 VDDA.t320 VDDA.n610 643.037
R4637 VDDA.n611 VDDA.t393 643.037
R4638 VDDA.t384 VDDA.n588 643.037
R4639 VDDA.n589 VDDA.t305 643.037
R4640 VDDA.n182 VDDA.n181 626.534
R4641 VDDA.n184 VDDA.n183 626.534
R4642 VDDA.n186 VDDA.n185 626.534
R4643 VDDA.n188 VDDA.n187 626.534
R4644 VDDA.n190 VDDA.n189 626.534
R4645 VDDA.n192 VDDA.n191 626.534
R4646 VDDA.n194 VDDA.n193 626.534
R4647 VDDA.n196 VDDA.n195 626.534
R4648 VDDA.n198 VDDA.n197 626.534
R4649 VDDA.n200 VDDA.n199 626.534
R4650 VDDA.n282 VDDA.t377 624.725
R4651 VDDA.n72 VDDA.t389 624.725
R4652 VDDA.n292 VDDA.t362 601.867
R4653 VDDA.n84 VDDA.t407 601.867
R4654 VDDA.n357 VDDA.n300 587.407
R4655 VDDA.n365 VDDA.n364 587.407
R4656 VDDA.n351 VDDA.n350 587.407
R4657 VDDA.n331 VDDA.n330 587.407
R4658 VDDA.n138 VDDA.n110 587.407
R4659 VDDA.n123 VDDA.n119 587.407
R4660 VDDA.n149 VDDA.n92 587.407
R4661 VDDA.n157 VDDA.n156 587.407
R4662 VDDA.n550 VDDA.n518 587.407
R4663 VDDA.n546 VDDA.n545 587.407
R4664 VDDA.n563 VDDA.n562 587.407
R4665 VDDA.n557 VDDA.n512 587.407
R4666 VDDA.n440 VDDA.n400 585
R4667 VDDA.n422 VDDA.n421 585
R4668 VDDA.n381 VDDA.n357 585
R4669 VDDA.n380 VDDA.n358 585
R4670 VDDA.n379 VDDA.n359 585
R4671 VDDA.n376 VDDA.n360 585
R4672 VDDA.n375 VDDA.n361 585
R4673 VDDA.n372 VDDA.n362 585
R4674 VDDA.n371 VDDA.n363 585
R4675 VDDA.n368 VDDA.n364 585
R4676 VDDA.n350 VDDA.n349 585
R4677 VDDA.n346 VDDA.n324 585
R4678 VDDA.n345 VDDA.n325 585
R4679 VDDA.n342 VDDA.n326 585
R4680 VDDA.n341 VDDA.n327 585
R4681 VDDA.n338 VDDA.n328 585
R4682 VDDA.n337 VDDA.n329 585
R4683 VDDA.n334 VDDA.n330 585
R4684 VDDA.n251 VDDA.n210 585
R4685 VDDA.n233 VDDA.n232 585
R4686 VDDA.n173 VDDA.n149 585
R4687 VDDA.n172 VDDA.n150 585
R4688 VDDA.n171 VDDA.n151 585
R4689 VDDA.n168 VDDA.n152 585
R4690 VDDA.n167 VDDA.n153 585
R4691 VDDA.n164 VDDA.n154 585
R4692 VDDA.n163 VDDA.n155 585
R4693 VDDA.n160 VDDA.n156 585
R4694 VDDA.n136 VDDA.n110 585
R4695 VDDA.n135 VDDA.n134 585
R4696 VDDA.n133 VDDA.n113 585
R4697 VDDA.n132 VDDA.n131 585
R4698 VDDA.n130 VDDA.n129 585
R4699 VDDA.n128 VDDA.n118 585
R4700 VDDA.n127 VDDA.n126 585
R4701 VDDA.n125 VDDA.n119 585
R4702 VDDA.n43 VDDA.n2 585
R4703 VDDA.n25 VDDA.n24 585
R4704 VDDA.n562 VDDA.n561 585
R4705 VDDA.n560 VDDA.n557 585
R4706 VDDA.n548 VDDA.n518 585
R4707 VDDA.n547 VDDA.n546 585
R4708 VDDA.t150 VDDA.t369 580.557
R4709 VDDA.t94 VDDA.t150 580.557
R4710 VDDA.t25 VDDA.t94 580.557
R4711 VDDA.t205 VDDA.t25 580.557
R4712 VDDA.t145 VDDA.t205 580.557
R4713 VDDA.t243 VDDA.t145 580.557
R4714 VDDA.t13 VDDA.t243 580.557
R4715 VDDA.t161 VDDA.t13 580.557
R4716 VDDA.t415 VDDA.t161 580.557
R4717 VDDA.t187 VDDA.t415 580.557
R4718 VDDA.t387 VDDA.t187 580.557
R4719 VDDA.t402 VDDA.t34 580.557
R4720 VDDA.t34 VDDA.t18 580.557
R4721 VDDA.t18 VDDA.t159 580.557
R4722 VDDA.t159 VDDA.t436 580.557
R4723 VDDA.t436 VDDA.t91 580.557
R4724 VDDA.t91 VDDA.t467 580.557
R4725 VDDA.t467 VDDA.t138 580.557
R4726 VDDA.t138 VDDA.t457 580.557
R4727 VDDA.t457 VDDA.t455 580.557
R4728 VDDA.t455 VDDA.t58 580.557
R4729 VDDA.t58 VDDA.t434 580.557
R4730 VDDA.t434 VDDA.t464 580.557
R4731 VDDA.t464 VDDA.t460 580.557
R4732 VDDA.t460 VDDA.t102 580.557
R4733 VDDA.t102 VDDA.t185 580.557
R4734 VDDA.t185 VDDA.t85 580.557
R4735 VDDA.t85 VDDA.t423 580.557
R4736 VDDA.t423 VDDA.t104 580.557
R4737 VDDA.t104 VDDA.t106 580.557
R4738 VDDA.t106 VDDA.t136 580.557
R4739 VDDA.t136 VDDA.t396 580.557
R4740 VDDA.t302 VDDA.t149 580.557
R4741 VDDA.t149 VDDA.t63 580.557
R4742 VDDA.t63 VDDA.t3 580.557
R4743 VDDA.t3 VDDA.t62 580.557
R4744 VDDA.t62 VDDA.t148 580.557
R4745 VDDA.t148 VDDA.t12 580.557
R4746 VDDA.t12 VDDA.t251 580.557
R4747 VDDA.t251 VDDA.t142 580.557
R4748 VDDA.t142 VDDA.t229 580.557
R4749 VDDA.t229 VDDA.t192 580.557
R4750 VDDA.t192 VDDA.t311 580.557
R4751 VDDA.n505 VDDA.t351 540.818
R4752 VDDA.n290 VDDA.t364 464.281
R4753 VDDA.n287 VDDA.t364 464.281
R4754 VDDA.n281 VDDA.t379 464.281
R4755 VDDA.t379 VDDA.n280 464.281
R4756 VDDA.n71 VDDA.t391 464.281
R4757 VDDA.t391 VDDA.n70 464.281
R4758 VDDA.t409 VDDA.n63 464.281
R4759 VDDA.n79 VDDA.t409 464.281
R4760 VDDA.n393 VDDA.t337 447.226
R4761 VDDA.n396 VDDA.t328 447.226
R4762 VDDA.n570 VDDA.t347 419.108
R4763 VDDA.n573 VDDA.t344 419.108
R4764 VDDA.n523 VDDA.t365 413.084
R4765 VDDA.n526 VDDA.t410 413.084
R4766 VDDA.n609 VDDA.t319 409.067
R4767 VDDA.n612 VDDA.t392 409.067
R4768 VDDA.n601 VDDA.t404 409.067
R4769 VDDA.n604 VDDA.t374 409.067
R4770 VDDA.n587 VDDA.t383 409.067
R4771 VDDA.t143 VDDA.t372 407.144
R4772 VDDA.t188 VDDA.t143 407.144
R4773 VDDA.t230 VDDA.t188 407.144
R4774 VDDA.t32 VDDA.t230 407.144
R4775 VDDA.t413 VDDA.t32 407.144
R4776 VDDA.t232 VDDA.t413 407.144
R4777 VDDA.t178 VDDA.t232 407.144
R4778 VDDA.t151 VDDA.t178 407.144
R4779 VDDA.t1 VDDA.t151 407.144
R4780 VDDA.t162 VDDA.t1 407.144
R4781 VDDA.t122 VDDA.t162 407.144
R4782 VDDA.t36 VDDA.t122 407.144
R4783 VDDA.t416 VDDA.t36 407.144
R4784 VDDA.t247 VDDA.t416 407.144
R4785 VDDA.t227 VDDA.t247 407.144
R4786 VDDA.t140 VDDA.t227 407.144
R4787 VDDA.t146 VDDA.t140 407.144
R4788 VDDA.t425 VDDA.t146 407.144
R4789 VDDA.t351 VDDA.t425 407.144
R4790 VDDA.t249 VDDA.t314 407.144
R4791 VDDA.t40 VDDA.t249 407.144
R4792 VDDA.t4 VDDA.t40 407.144
R4793 VDDA.t50 VDDA.t4 407.144
R4794 VDDA.t130 VDDA.t50 407.144
R4795 VDDA.t89 VDDA.t130 407.144
R4796 VDDA.t87 VDDA.t89 407.144
R4797 VDDA.t225 VDDA.t87 407.144
R4798 VDDA.t164 VDDA.t225 407.144
R4799 VDDA.t432 VDDA.t164 407.144
R4800 VDDA.t48 VDDA.t432 407.144
R4801 VDDA.t38 VDDA.t48 407.144
R4802 VDDA.t176 VDDA.t38 407.144
R4803 VDDA.t46 VDDA.t176 407.144
R4804 VDDA.t116 VDDA.t46 407.144
R4805 VDDA.t132 VDDA.t116 407.144
R4806 VDDA.t30 VDDA.t132 407.144
R4807 VDDA.t118 VDDA.t30 407.144
R4808 VDDA.t335 VDDA.t118 407.144
R4809 VDDA.n590 VDDA.t304 390.322
R4810 VDDA.n503 VDDA.t371 379.582
R4811 VDDA.n480 VDDA.t313 379.582
R4812 VDDA.t350 VDDA.n506 379.277
R4813 VDDA.t23 VDDA.t348 373.214
R4814 VDDA.t245 VDDA.t23 373.214
R4815 VDDA.t345 VDDA.t245 373.214
R4816 VDDA.t93 VDDA.t366 373.214
R4817 VDDA.t244 VDDA.t93 373.214
R4818 VDDA.t411 VDDA.t244 373.214
R4819 VDDA.t28 VDDA.t320 373.214
R4820 VDDA.t448 VDDA.t28 373.214
R4821 VDDA.t78 VDDA.t448 373.214
R4822 VDDA.t10 VDDA.t78 373.214
R4823 VDDA.t393 VDDA.t10 373.214
R4824 VDDA.t112 VDDA.t405 373.214
R4825 VDDA.t110 VDDA.t112 373.214
R4826 VDDA.t223 VDDA.t110 373.214
R4827 VDDA.t442 VDDA.t223 373.214
R4828 VDDA.t80 VDDA.t442 373.214
R4829 VDDA.t60 VDDA.t80 373.214
R4830 VDDA.t203 VDDA.t60 373.214
R4831 VDDA.t199 VDDA.t203 373.214
R4832 VDDA.t201 VDDA.t199 373.214
R4833 VDDA.t444 VDDA.t201 373.214
R4834 VDDA.t375 VDDA.t444 373.214
R4835 VDDA.t44 VDDA.t384 373.214
R4836 VDDA.t430 VDDA.t44 373.214
R4837 VDDA.t114 VDDA.t430 373.214
R4838 VDDA.t82 VDDA.t114 373.214
R4839 VDDA.t305 VDDA.t82 373.214
R4840 VDDA.n295 VDDA.t368 365.884
R4841 VDDA.n294 VDDA.t386 365.884
R4842 VDDA.n86 VDDA.t310 365.884
R4843 VDDA.n87 VDDA.t301 365.884
R4844 VDDA.n543 VDDA.t331 360.868
R4845 VDDA.n568 VDDA.t298 360.868
R4846 VDDA.n507 VDDA.t350 358.858
R4847 VDDA.t371 VDDA.n502 358.858
R4848 VDDA.n483 VDDA.t334 358.858
R4849 VDDA.t313 VDDA.n479 358.858
R4850 VDDA.n602 VDDA.t406 354.154
R4851 VDDA.n603 VDDA.t376 354.154
R4852 VDDA.n482 VDDA.t336 354.065
R4853 VDDA.n572 VDDA.t346 354.065
R4854 VDDA.n571 VDDA.t349 354.063
R4855 VDDA.n524 VDDA.t367 354.063
R4856 VDDA.n458 VDDA.t352 351.793
R4857 VDDA.n525 VDDA.t412 347.224
R4858 VDDA.n584 VDDA.n583 345.127
R4859 VDDA.n586 VDDA.n585 345.127
R4860 VDDA.n580 VDDA.n579 344.7
R4861 VDDA.n607 VDDA.n606 344.7
R4862 VDDA.n456 VDDA.n455 341.675
R4863 VDDA.n486 VDDA.n485 341.675
R4864 VDDA.n488 VDDA.n487 341.675
R4865 VDDA.n490 VDDA.n489 341.675
R4866 VDDA.n492 VDDA.n491 341.675
R4867 VDDA.n494 VDDA.n493 341.675
R4868 VDDA.n496 VDDA.n495 341.675
R4869 VDDA.n498 VDDA.n497 341.675
R4870 VDDA.n500 VDDA.n499 341.675
R4871 VDDA.n461 VDDA.n460 341.675
R4872 VDDA.n464 VDDA.n463 341.675
R4873 VDDA.n466 VDDA.n465 341.675
R4874 VDDA.n468 VDDA.n467 341.675
R4875 VDDA.n470 VDDA.n469 341.675
R4876 VDDA.n472 VDDA.n471 341.675
R4877 VDDA.n474 VDDA.n473 341.675
R4878 VDDA.n476 VDDA.n475 341.675
R4879 VDDA.n478 VDDA.n477 341.675
R4880 VDDA.n582 VDDA.n581 339.272
R4881 VDDA.n593 VDDA.n592 339.272
R4882 VDDA.n595 VDDA.n594 339.272
R4883 VDDA.n597 VDDA.n596 339.272
R4884 VDDA.n599 VDDA.n598 339.272
R4885 VDDA.n576 VDDA.n575 334.772
R4886 VDDA.n588 VDDA.t385 332.267
R4887 VDDA.n589 VDDA.t306 332.267
R4888 VDDA.n610 VDDA.t321 332.084
R4889 VDDA.n611 VDDA.t394 332.084
R4890 VDDA.n201 VDDA.t395 328.733
R4891 VDDA.n204 VDDA.t401 328.733
R4892 VDDA.n428 VDDA.n400 290.233
R4893 VDDA.n434 VDDA.n400 290.233
R4894 VDDA.n429 VDDA.n400 290.233
R4895 VDDA.n421 VDDA.n409 290.233
R4896 VDDA.n421 VDDA.n414 290.233
R4897 VDDA.n421 VDDA.n419 290.233
R4898 VDDA.n239 VDDA.n210 290.233
R4899 VDDA.n245 VDDA.n210 290.233
R4900 VDDA.n240 VDDA.n210 290.233
R4901 VDDA.n232 VDDA.n221 290.233
R4902 VDDA.n232 VDDA.n226 290.233
R4903 VDDA.n232 VDDA.n231 290.233
R4904 VDDA.n31 VDDA.n2 290.233
R4905 VDDA.n37 VDDA.n2 290.233
R4906 VDDA.n32 VDDA.n2 290.233
R4907 VDDA.n24 VDDA.n13 290.233
R4908 VDDA.n24 VDDA.n18 290.233
R4909 VDDA.n24 VDDA.n23 290.233
R4910 VDDA.n285 VDDA.t363 267.188
R4911 VDDA.t378 VDDA.n284 267.188
R4912 VDDA.t390 VDDA.n74 267.188
R4913 VDDA.n81 VDDA.t408 267.188
R4914 VDDA.t329 VDDA.t190 259.091
R4915 VDDA.t190 VDDA.t338 259.091
R4916 VDDA.t220 VDDA.t332 251.471
R4917 VDDA.t212 VDDA.t220 251.471
R4918 VDDA.t95 VDDA.t212 251.471
R4919 VDDA.t207 VDDA.t95 251.471
R4920 VDDA.t125 VDDA.t207 251.471
R4921 VDDA.t73 VDDA.t125 251.471
R4922 VDDA.t216 VDDA.t73 251.471
R4923 VDDA.t56 VDDA.t216 251.471
R4924 VDDA.t127 VDDA.t56 251.471
R4925 VDDA.t218 VDDA.t127 251.471
R4926 VDDA.t418 VDDA.t218 251.471
R4927 VDDA.t420 VDDA.t418 251.471
R4928 VDDA.t65 VDDA.t420 251.471
R4929 VDDA.t52 VDDA.t65 251.471
R4930 VDDA.t70 VDDA.t52 251.471
R4931 VDDA.t166 VDDA.t70 251.471
R4932 VDDA.t299 VDDA.t166 251.471
R4933 VDDA.n358 VDDA.n357 246.25
R4934 VDDA.n359 VDDA.n358 246.25
R4935 VDDA.n360 VDDA.n359 246.25
R4936 VDDA.n362 VDDA.n361 246.25
R4937 VDDA.n363 VDDA.n362 246.25
R4938 VDDA.n364 VDDA.n363 246.25
R4939 VDDA.n350 VDDA.n324 246.25
R4940 VDDA.n325 VDDA.n324 246.25
R4941 VDDA.n326 VDDA.n325 246.25
R4942 VDDA.n328 VDDA.n327 246.25
R4943 VDDA.n329 VDDA.n328 246.25
R4944 VDDA.n330 VDDA.n329 246.25
R4945 VDDA.n134 VDDA.n110 246.25
R4946 VDDA.n134 VDDA.n133 246.25
R4947 VDDA.n133 VDDA.n132 246.25
R4948 VDDA.n129 VDDA.n128 246.25
R4949 VDDA.n128 VDDA.n127 246.25
R4950 VDDA.n127 VDDA.n119 246.25
R4951 VDDA.n150 VDDA.n149 246.25
R4952 VDDA.n151 VDDA.n150 246.25
R4953 VDDA.n152 VDDA.n151 246.25
R4954 VDDA.n154 VDDA.n153 246.25
R4955 VDDA.n155 VDDA.n154 246.25
R4956 VDDA.n156 VDDA.n155 246.25
R4957 VDDA.n280 VDDA.n275 243.698
R4958 VDDA.n70 VDDA.n65 243.698
R4959 VDDA.n564 VDDA.n563 243.698
R4960 VDDA.n429 VDDA.n426 242.903
R4961 VDDA.n419 VDDA.n405 242.903
R4962 VDDA.n240 VDDA.n237 242.903
R4963 VDDA.n231 VDDA.n215 242.903
R4964 VDDA.n32 VDDA.n29 242.903
R4965 VDDA.n23 VDDA.n7 242.903
R4966 VDDA.n440 VDDA.n439 238.367
R4967 VDDA.n385 VDDA.n384 238.367
R4968 VDDA.n283 VDDA.n282 238.367
R4969 VDDA.n251 VDDA.n250 238.367
R4970 VDDA.n177 VDDA.n176 238.367
R4971 VDDA.n73 VDDA.n72 238.367
R4972 VDDA.n43 VDDA.n42 238.367
R4973 VDDA.n506 VDDA.n505 238.367
R4974 VDDA.n505 VDDA.n457 238.367
R4975 VDDA.t332 VDDA.n552 237.5
R4976 VDDA.n565 VDDA.t299 237.5
R4977 VDDA.t363 VDDA.t462 217.708
R4978 VDDA.t462 VDDA.t174 217.708
R4979 VDDA.t174 VDDA.t64 217.708
R4980 VDDA.t64 VDDA.t183 217.708
R4981 VDDA.t183 VDDA.t184 217.708
R4982 VDDA.t184 VDDA.t459 217.708
R4983 VDDA.t459 VDDA.t466 217.708
R4984 VDDA.t466 VDDA.t429 217.708
R4985 VDDA.t429 VDDA.t157 217.708
R4986 VDDA.t157 VDDA.t181 217.708
R4987 VDDA.t181 VDDA.t378 217.708
R4988 VDDA.t196 VDDA.t390 217.708
R4989 VDDA.t234 VDDA.t196 217.708
R4990 VDDA.t109 VDDA.t234 217.708
R4991 VDDA.t121 VDDA.t109 217.708
R4992 VDDA.t20 VDDA.t121 217.708
R4993 VDDA.t447 VDDA.t20 217.708
R4994 VDDA.t175 VDDA.t447 217.708
R4995 VDDA.t237 VDDA.t175 217.708
R4996 VDDA.t77 VDDA.t237 217.708
R4997 VDDA.t43 VDDA.t77 217.708
R4998 VDDA.t408 VDDA.t43 217.708
R4999 VDDA.n365 VDDA.n306 190.333
R5000 VDDA.n331 VDDA.n312 190.333
R5001 VDDA.n287 VDDA.n286 190.333
R5002 VDDA.n157 VDDA.n146 190.333
R5003 VDDA.n123 VDDA.n99 190.333
R5004 VDDA.n80 VDDA.n79 190.333
R5005 VDDA.n551 VDDA.n550 190.333
R5006 VDDA.n402 VDDA.n401 185
R5007 VDDA.n437 VDDA.n436 185
R5008 VDDA.n438 VDDA.n437 185
R5009 VDDA.n435 VDDA.n427 185
R5010 VDDA.n433 VDDA.n432 185
R5011 VDDA.n431 VDDA.n430 185
R5012 VDDA.n423 VDDA.n422 185
R5013 VDDA.n424 VDDA.n423 185
R5014 VDDA.n408 VDDA.n406 185
R5015 VDDA.n411 VDDA.n410 185
R5016 VDDA.n413 VDDA.n412 185
R5017 VDDA.n416 VDDA.n415 185
R5018 VDDA.n418 VDDA.n417 185
R5019 VDDA.n356 VDDA.n301 185
R5020 VDDA.n382 VDDA.n381 185
R5021 VDDA.n383 VDDA.n382 185
R5022 VDDA.n380 VDDA.n355 185
R5023 VDDA.n379 VDDA.n378 185
R5024 VDDA.n377 VDDA.n376 185
R5025 VDDA.n375 VDDA.n374 185
R5026 VDDA.n373 VDDA.n372 185
R5027 VDDA.n371 VDDA.n370 185
R5028 VDDA.n369 VDDA.n368 185
R5029 VDDA.n367 VDDA.n366 185
R5030 VDDA.n383 VDDA.n306 185
R5031 VDDA.n353 VDDA.n352 185
R5032 VDDA.n354 VDDA.n353 185
R5033 VDDA.n323 VDDA.n313 185
R5034 VDDA.n349 VDDA.n348 185
R5035 VDDA.n347 VDDA.n346 185
R5036 VDDA.n345 VDDA.n344 185
R5037 VDDA.n343 VDDA.n342 185
R5038 VDDA.n341 VDDA.n340 185
R5039 VDDA.n339 VDDA.n338 185
R5040 VDDA.n337 VDDA.n336 185
R5041 VDDA.n335 VDDA.n334 185
R5042 VDDA.n333 VDDA.n332 185
R5043 VDDA.n354 VDDA.n312 185
R5044 VDDA.n277 VDDA.n276 185
R5045 VDDA.n279 VDDA.n278 185
R5046 VDDA.n291 VDDA.n271 185
R5047 VDDA.n285 VDDA.n271 185
R5048 VDDA.n289 VDDA.n272 185
R5049 VDDA.n288 VDDA.n273 185
R5050 VDDA.n286 VDDA.n285 185
R5051 VDDA.n212 VDDA.n211 185
R5052 VDDA.n248 VDDA.n247 185
R5053 VDDA.n249 VDDA.n248 185
R5054 VDDA.n246 VDDA.n238 185
R5055 VDDA.n244 VDDA.n243 185
R5056 VDDA.n242 VDDA.n241 185
R5057 VDDA.n234 VDDA.n233 185
R5058 VDDA.n235 VDDA.n234 185
R5059 VDDA.n220 VDDA.n216 185
R5060 VDDA.n223 VDDA.n222 185
R5061 VDDA.n225 VDDA.n224 185
R5062 VDDA.n228 VDDA.n227 185
R5063 VDDA.n230 VDDA.n229 185
R5064 VDDA.n148 VDDA.n93 185
R5065 VDDA.n174 VDDA.n173 185
R5066 VDDA.n175 VDDA.n174 185
R5067 VDDA.n172 VDDA.n147 185
R5068 VDDA.n171 VDDA.n170 185
R5069 VDDA.n169 VDDA.n168 185
R5070 VDDA.n167 VDDA.n166 185
R5071 VDDA.n165 VDDA.n164 185
R5072 VDDA.n163 VDDA.n162 185
R5073 VDDA.n161 VDDA.n160 185
R5074 VDDA.n159 VDDA.n158 185
R5075 VDDA.n175 VDDA.n146 185
R5076 VDDA.n140 VDDA.n139 185
R5077 VDDA.n141 VDDA.n140 185
R5078 VDDA.n137 VDDA.n100 185
R5079 VDDA.n136 VDDA.n111 185
R5080 VDDA.n135 VDDA.n112 185
R5081 VDDA.n114 VDDA.n113 185
R5082 VDDA.n131 VDDA.n115 185
R5083 VDDA.n130 VDDA.n116 185
R5084 VDDA.n118 VDDA.n117 185
R5085 VDDA.n126 VDDA.n120 185
R5086 VDDA.n125 VDDA.n121 185
R5087 VDDA.n124 VDDA.n122 185
R5088 VDDA.n141 VDDA.n99 185
R5089 VDDA.n67 VDDA.n66 185
R5090 VDDA.n69 VDDA.n68 185
R5091 VDDA.n83 VDDA.n82 185
R5092 VDDA.n82 VDDA.n81 185
R5093 VDDA.n77 VDDA.n64 185
R5094 VDDA.n78 VDDA.n76 185
R5095 VDDA.n81 VDDA.n80 185
R5096 VDDA.n4 VDDA.n3 185
R5097 VDDA.n40 VDDA.n39 185
R5098 VDDA.n41 VDDA.n40 185
R5099 VDDA.n38 VDDA.n30 185
R5100 VDDA.n36 VDDA.n35 185
R5101 VDDA.n34 VDDA.n33 185
R5102 VDDA.n26 VDDA.n25 185
R5103 VDDA.n27 VDDA.n26 185
R5104 VDDA.n12 VDDA.n8 185
R5105 VDDA.n15 VDDA.n14 185
R5106 VDDA.n17 VDDA.n16 185
R5107 VDDA.n20 VDDA.n19 185
R5108 VDDA.n22 VDDA.n21 185
R5109 VDDA.n556 VDDA.n555 185
R5110 VDDA.n561 VDDA.n554 185
R5111 VDDA.n565 VDDA.n554 185
R5112 VDDA.n560 VDDA.n559 185
R5113 VDDA.n558 VDDA.n513 185
R5114 VDDA.n567 VDDA.n566 185
R5115 VDDA.n566 VDDA.n565 185
R5116 VDDA.n552 VDDA.n551 185
R5117 VDDA.n549 VDDA.n517 185
R5118 VDDA.n548 VDDA.n519 185
R5119 VDDA.n547 VDDA.n520 185
R5120 VDDA.n522 VDDA.n521 185
R5121 VDDA.n544 VDDA.n516 185
R5122 VDDA.n552 VDDA.n516 185
R5123 VDDA.t360 VDDA.n424 170.513
R5124 VDDA.n438 VDDA.t381 170.513
R5125 VDDA.t323 VDDA.n235 170.513
R5126 VDDA.n249 VDDA.t399 170.513
R5127 VDDA.t354 VDDA.n27 170.513
R5128 VDDA.n41 VDDA.t308 170.513
R5129 VDDA.n511 VDDA.n510 168.435
R5130 VDDA.n529 VDDA.n528 168.435
R5131 VDDA.n531 VDDA.n530 168.435
R5132 VDDA.n533 VDDA.n532 168.435
R5133 VDDA.n535 VDDA.n534 168.435
R5134 VDDA.n537 VDDA.n536 168.435
R5135 VDDA.n539 VDDA.n538 168.435
R5136 VDDA.n541 VDDA.n540 168.435
R5137 VDDA.n420 VDDA.n399 159.803
R5138 VDDA.n209 VDDA.n208 159.803
R5139 VDDA.n218 VDDA.n217 159.803
R5140 VDDA.n254 VDDA.n253 159.803
R5141 VDDA.n256 VDDA.n255 159.803
R5142 VDDA.n1 VDDA.n0 159.803
R5143 VDDA.n10 VDDA.n9 159.803
R5144 VDDA.n46 VDDA.n45 159.803
R5145 VDDA.n48 VDDA.n47 159.803
R5146 VDDA.n259 VDDA.n258 155.303
R5147 VDDA.n51 VDDA.n50 155.303
R5148 VDDA.n437 VDDA.n402 150
R5149 VDDA.n437 VDDA.n427 150
R5150 VDDA.n432 VDDA.n431 150
R5151 VDDA.n423 VDDA.n406 150
R5152 VDDA.n412 VDDA.n411 150
R5153 VDDA.n417 VDDA.n416 150
R5154 VDDA.n382 VDDA.n301 150
R5155 VDDA.n382 VDDA.n355 150
R5156 VDDA.n378 VDDA.n377 150
R5157 VDDA.n374 VDDA.n373 150
R5158 VDDA.n370 VDDA.n369 150
R5159 VDDA.n366 VDDA.n306 150
R5160 VDDA.n353 VDDA.n313 150
R5161 VDDA.n348 VDDA.n347 150
R5162 VDDA.n344 VDDA.n343 150
R5163 VDDA.n340 VDDA.n339 150
R5164 VDDA.n336 VDDA.n335 150
R5165 VDDA.n332 VDDA.n312 150
R5166 VDDA.n278 VDDA.n276 150
R5167 VDDA.n272 VDDA.n271 150
R5168 VDDA.n286 VDDA.n273 150
R5169 VDDA.n248 VDDA.n212 150
R5170 VDDA.n248 VDDA.n238 150
R5171 VDDA.n243 VDDA.n242 150
R5172 VDDA.n234 VDDA.n216 150
R5173 VDDA.n224 VDDA.n223 150
R5174 VDDA.n229 VDDA.n228 150
R5175 VDDA.n174 VDDA.n93 150
R5176 VDDA.n174 VDDA.n147 150
R5177 VDDA.n170 VDDA.n169 150
R5178 VDDA.n166 VDDA.n165 150
R5179 VDDA.n162 VDDA.n161 150
R5180 VDDA.n158 VDDA.n146 150
R5181 VDDA.n140 VDDA.n100 150
R5182 VDDA.n112 VDDA.n111 150
R5183 VDDA.n115 VDDA.n114 150
R5184 VDDA.n117 VDDA.n116 150
R5185 VDDA.n121 VDDA.n120 150
R5186 VDDA.n122 VDDA.n99 150
R5187 VDDA.n68 VDDA.n66 150
R5188 VDDA.n82 VDDA.n64 150
R5189 VDDA.n80 VDDA.n76 150
R5190 VDDA.n40 VDDA.n4 150
R5191 VDDA.n40 VDDA.n30 150
R5192 VDDA.n35 VDDA.n34 150
R5193 VDDA.n26 VDDA.n8 150
R5194 VDDA.n16 VDDA.n15 150
R5195 VDDA.n21 VDDA.n20 150
R5196 VDDA.n555 VDDA.n554 150
R5197 VDDA.n559 VDDA.n554 150
R5198 VDDA.n566 VDDA.n513 150
R5199 VDDA.n551 VDDA.n517 150
R5200 VDDA.n520 VDDA.n519 150
R5201 VDDA.n521 VDDA.n516 150
R5202 VDDA.t280 VDDA.t360 146.155
R5203 VDDA.t381 VDDA.t280 146.155
R5204 VDDA.t264 VDDA.t323 146.155
R5205 VDDA.t260 VDDA.t264 146.155
R5206 VDDA.t268 VDDA.t260 146.155
R5207 VDDA.t278 VDDA.t268 146.155
R5208 VDDA.t288 VDDA.t278 146.155
R5209 VDDA.t258 VDDA.t288 146.155
R5210 VDDA.t256 VDDA.t258 146.155
R5211 VDDA.t262 VDDA.t256 146.155
R5212 VDDA.t270 VDDA.t262 146.155
R5213 VDDA.t282 VDDA.t270 146.155
R5214 VDDA.t399 VDDA.t282 146.155
R5215 VDDA.t276 VDDA.t354 146.155
R5216 VDDA.t272 VDDA.t276 146.155
R5217 VDDA.t284 VDDA.t272 146.155
R5218 VDDA.t290 VDDA.t284 146.155
R5219 VDDA.t252 VDDA.t290 146.155
R5220 VDDA.t254 VDDA.t252 146.155
R5221 VDDA.t266 VDDA.t254 146.155
R5222 VDDA.t274 VDDA.t266 146.155
R5223 VDDA.t286 VDDA.t274 146.155
R5224 VDDA.t292 VDDA.t286 146.155
R5225 VDDA.t308 VDDA.t292 146.155
R5226 VDDA.n299 VDDA.n298 145.429
R5227 VDDA.n315 VDDA.n314 145.429
R5228 VDDA.n317 VDDA.n316 145.429
R5229 VDDA.n319 VDDA.n318 145.429
R5230 VDDA.n321 VDDA.n320 145.429
R5231 VDDA.n91 VDDA.n90 145.429
R5232 VDDA.n102 VDDA.n101 145.429
R5233 VDDA.n104 VDDA.n103 145.429
R5234 VDDA.n106 VDDA.n105 145.429
R5235 VDDA.n108 VDDA.n107 145.429
R5236 VDDA.t318 VDDA.n360 123.126
R5237 VDDA.n361 VDDA.t318 123.126
R5238 VDDA.t327 VDDA.n326 123.126
R5239 VDDA.n327 VDDA.t327 123.126
R5240 VDDA.n132 VDDA.t343 123.126
R5241 VDDA.n129 VDDA.t343 123.126
R5242 VDDA.t358 VDDA.n152 123.126
R5243 VDDA.n153 VDDA.t358 123.126
R5244 VDDA.t333 VDDA.n518 123.126
R5245 VDDA.n546 VDDA.t333 123.126
R5246 VDDA.n562 VDDA.t300 123.126
R5247 VDDA.n557 VDDA.t300 123.126
R5248 VDDA.n383 VDDA.t317 100.195
R5249 VDDA.t326 VDDA.n354 100.195
R5250 VDDA.t342 VDDA.n141 100.195
R5251 VDDA.n175 VDDA.t357 100.195
R5252 VDDA.n262 VDDA.n260 97.4002
R5253 VDDA.n54 VDDA.n52 97.4002
R5254 VDDA.n270 VDDA.n269 96.8377
R5255 VDDA.n268 VDDA.n267 96.8377
R5256 VDDA.n266 VDDA.n265 96.8377
R5257 VDDA.n264 VDDA.n263 96.8377
R5258 VDDA.n262 VDDA.n261 96.8377
R5259 VDDA.n62 VDDA.n61 96.8377
R5260 VDDA.n60 VDDA.n59 96.8377
R5261 VDDA.n58 VDDA.n57 96.8377
R5262 VDDA.n56 VDDA.n55 96.8377
R5263 VDDA.n54 VDDA.n53 96.8377
R5264 VDDA.t317 VDDA.t134 81.6411
R5265 VDDA.t134 VDDA.t210 81.6411
R5266 VDDA.t210 VDDA.t16 81.6411
R5267 VDDA.t16 VDDA.t153 81.6411
R5268 VDDA.t153 VDDA.t155 81.6411
R5269 VDDA.t155 VDDA.t427 81.6411
R5270 VDDA.t427 VDDA.t451 81.6411
R5271 VDDA.t451 VDDA.t172 81.6411
R5272 VDDA.t172 VDDA.t14 81.6411
R5273 VDDA.t14 VDDA.t453 81.6411
R5274 VDDA.t453 VDDA.t326 81.6411
R5275 VDDA.t241 VDDA.t342 81.6411
R5276 VDDA.t8 VDDA.t241 81.6411
R5277 VDDA.t238 VDDA.t8 81.6411
R5278 VDDA.t197 VDDA.t238 81.6411
R5279 VDDA.t235 VDDA.t197 81.6411
R5280 VDDA.t193 VDDA.t235 81.6411
R5281 VDDA.t440 VDDA.t193 81.6411
R5282 VDDA.t6 VDDA.t440 81.6411
R5283 VDDA.t438 VDDA.t6 81.6411
R5284 VDDA.t21 VDDA.t438 81.6411
R5285 VDDA.t357 VDDA.t21 81.6411
R5286 VDDA.n181 VDDA.t35 78.8005
R5287 VDDA.n181 VDDA.t19 78.8005
R5288 VDDA.n183 VDDA.t160 78.8005
R5289 VDDA.n183 VDDA.t437 78.8005
R5290 VDDA.n185 VDDA.t92 78.8005
R5291 VDDA.n185 VDDA.t468 78.8005
R5292 VDDA.n187 VDDA.t139 78.8005
R5293 VDDA.n187 VDDA.t458 78.8005
R5294 VDDA.n189 VDDA.t456 78.8005
R5295 VDDA.n189 VDDA.t59 78.8005
R5296 VDDA.n191 VDDA.t435 78.8005
R5297 VDDA.n191 VDDA.t465 78.8005
R5298 VDDA.n193 VDDA.t461 78.8005
R5299 VDDA.n193 VDDA.t103 78.8005
R5300 VDDA.n195 VDDA.t186 78.8005
R5301 VDDA.n195 VDDA.t86 78.8005
R5302 VDDA.n197 VDDA.t424 78.8005
R5303 VDDA.n197 VDDA.t105 78.8005
R5304 VDDA.n199 VDDA.t107 78.8005
R5305 VDDA.n199 VDDA.t137 78.8005
R5306 VDDA.n439 VDDA.n438 65.8183
R5307 VDDA.n438 VDDA.n425 65.8183
R5308 VDDA.n438 VDDA.n426 65.8183
R5309 VDDA.n424 VDDA.n403 65.8183
R5310 VDDA.n424 VDDA.n404 65.8183
R5311 VDDA.n424 VDDA.n405 65.8183
R5312 VDDA.n384 VDDA.n383 65.8183
R5313 VDDA.n383 VDDA.n302 65.8183
R5314 VDDA.n383 VDDA.n303 65.8183
R5315 VDDA.n383 VDDA.n304 65.8183
R5316 VDDA.n383 VDDA.n305 65.8183
R5317 VDDA.n354 VDDA.n307 65.8183
R5318 VDDA.n354 VDDA.n308 65.8183
R5319 VDDA.n354 VDDA.n309 65.8183
R5320 VDDA.n354 VDDA.n310 65.8183
R5321 VDDA.n354 VDDA.n311 65.8183
R5322 VDDA.n284 VDDA.n283 65.8183
R5323 VDDA.n284 VDDA.n275 65.8183
R5324 VDDA.n285 VDDA.n274 65.8183
R5325 VDDA.n250 VDDA.n249 65.8183
R5326 VDDA.n249 VDDA.n236 65.8183
R5327 VDDA.n249 VDDA.n237 65.8183
R5328 VDDA.n235 VDDA.n213 65.8183
R5329 VDDA.n235 VDDA.n214 65.8183
R5330 VDDA.n235 VDDA.n215 65.8183
R5331 VDDA.n176 VDDA.n175 65.8183
R5332 VDDA.n175 VDDA.n142 65.8183
R5333 VDDA.n175 VDDA.n143 65.8183
R5334 VDDA.n175 VDDA.n144 65.8183
R5335 VDDA.n175 VDDA.n145 65.8183
R5336 VDDA.n141 VDDA.n94 65.8183
R5337 VDDA.n141 VDDA.n95 65.8183
R5338 VDDA.n141 VDDA.n96 65.8183
R5339 VDDA.n141 VDDA.n97 65.8183
R5340 VDDA.n141 VDDA.n98 65.8183
R5341 VDDA.n74 VDDA.n73 65.8183
R5342 VDDA.n74 VDDA.n65 65.8183
R5343 VDDA.n81 VDDA.n75 65.8183
R5344 VDDA.n42 VDDA.n41 65.8183
R5345 VDDA.n41 VDDA.n28 65.8183
R5346 VDDA.n41 VDDA.n29 65.8183
R5347 VDDA.n27 VDDA.n5 65.8183
R5348 VDDA.n27 VDDA.n6 65.8183
R5349 VDDA.n27 VDDA.n7 65.8183
R5350 VDDA.n565 VDDA.n564 65.8183
R5351 VDDA.n565 VDDA.n553 65.8183
R5352 VDDA.n552 VDDA.n514 65.8183
R5353 VDDA.n552 VDDA.n515 65.8183
R5354 VDDA.n452 VDDA.t471 59.5681
R5355 VDDA.n451 VDDA.t472 59.5681
R5356 VDDA.n427 VDDA.n425 53.3664
R5357 VDDA.n431 VDDA.n426 53.3664
R5358 VDDA.n439 VDDA.n402 53.3664
R5359 VDDA.n432 VDDA.n425 53.3664
R5360 VDDA.n406 VDDA.n403 53.3664
R5361 VDDA.n412 VDDA.n404 53.3664
R5362 VDDA.n417 VDDA.n405 53.3664
R5363 VDDA.n411 VDDA.n403 53.3664
R5364 VDDA.n416 VDDA.n404 53.3664
R5365 VDDA.n355 VDDA.n302 53.3664
R5366 VDDA.n377 VDDA.n303 53.3664
R5367 VDDA.n373 VDDA.n304 53.3664
R5368 VDDA.n369 VDDA.n305 53.3664
R5369 VDDA.n384 VDDA.n301 53.3664
R5370 VDDA.n378 VDDA.n302 53.3664
R5371 VDDA.n374 VDDA.n303 53.3664
R5372 VDDA.n370 VDDA.n304 53.3664
R5373 VDDA.n366 VDDA.n305 53.3664
R5374 VDDA.n313 VDDA.n307 53.3664
R5375 VDDA.n347 VDDA.n308 53.3664
R5376 VDDA.n343 VDDA.n309 53.3664
R5377 VDDA.n339 VDDA.n310 53.3664
R5378 VDDA.n335 VDDA.n311 53.3664
R5379 VDDA.n348 VDDA.n307 53.3664
R5380 VDDA.n344 VDDA.n308 53.3664
R5381 VDDA.n340 VDDA.n309 53.3664
R5382 VDDA.n336 VDDA.n310 53.3664
R5383 VDDA.n332 VDDA.n311 53.3664
R5384 VDDA.n283 VDDA.n276 53.3664
R5385 VDDA.n278 VDDA.n275 53.3664
R5386 VDDA.n274 VDDA.n272 53.3664
R5387 VDDA.n274 VDDA.n273 53.3664
R5388 VDDA.n238 VDDA.n236 53.3664
R5389 VDDA.n242 VDDA.n237 53.3664
R5390 VDDA.n250 VDDA.n212 53.3664
R5391 VDDA.n243 VDDA.n236 53.3664
R5392 VDDA.n216 VDDA.n213 53.3664
R5393 VDDA.n224 VDDA.n214 53.3664
R5394 VDDA.n229 VDDA.n215 53.3664
R5395 VDDA.n223 VDDA.n213 53.3664
R5396 VDDA.n228 VDDA.n214 53.3664
R5397 VDDA.n147 VDDA.n142 53.3664
R5398 VDDA.n169 VDDA.n143 53.3664
R5399 VDDA.n165 VDDA.n144 53.3664
R5400 VDDA.n161 VDDA.n145 53.3664
R5401 VDDA.n176 VDDA.n93 53.3664
R5402 VDDA.n170 VDDA.n142 53.3664
R5403 VDDA.n166 VDDA.n143 53.3664
R5404 VDDA.n162 VDDA.n144 53.3664
R5405 VDDA.n158 VDDA.n145 53.3664
R5406 VDDA.n100 VDDA.n94 53.3664
R5407 VDDA.n112 VDDA.n95 53.3664
R5408 VDDA.n115 VDDA.n96 53.3664
R5409 VDDA.n117 VDDA.n97 53.3664
R5410 VDDA.n121 VDDA.n98 53.3664
R5411 VDDA.n111 VDDA.n94 53.3664
R5412 VDDA.n114 VDDA.n95 53.3664
R5413 VDDA.n116 VDDA.n96 53.3664
R5414 VDDA.n120 VDDA.n97 53.3664
R5415 VDDA.n122 VDDA.n98 53.3664
R5416 VDDA.n73 VDDA.n66 53.3664
R5417 VDDA.n68 VDDA.n65 53.3664
R5418 VDDA.n75 VDDA.n64 53.3664
R5419 VDDA.n76 VDDA.n75 53.3664
R5420 VDDA.n30 VDDA.n28 53.3664
R5421 VDDA.n34 VDDA.n29 53.3664
R5422 VDDA.n42 VDDA.n4 53.3664
R5423 VDDA.n35 VDDA.n28 53.3664
R5424 VDDA.n8 VDDA.n5 53.3664
R5425 VDDA.n16 VDDA.n6 53.3664
R5426 VDDA.n21 VDDA.n7 53.3664
R5427 VDDA.n15 VDDA.n5 53.3664
R5428 VDDA.n20 VDDA.n6 53.3664
R5429 VDDA.n559 VDDA.n553 53.3664
R5430 VDDA.n564 VDDA.n555 53.3664
R5431 VDDA.n553 VDDA.n513 53.3664
R5432 VDDA.n517 VDDA.n514 53.3664
R5433 VDDA.n520 VDDA.n515 53.3664
R5434 VDDA.n519 VDDA.n514 53.3664
R5435 VDDA.n521 VDDA.n515 53.3664
R5436 VDDA.n451 VDDA.t470 52.3888
R5437 VDDA.n453 VDDA.t469 48.9557
R5438 VDDA.n396 VDDA.n395 46.6291
R5439 VDDA.n394 VDDA.n393 46.6291
R5440 VDDA.n455 VDDA.t147 39.4005
R5441 VDDA.n455 VDDA.t426 39.4005
R5442 VDDA.n485 VDDA.t228 39.4005
R5443 VDDA.n485 VDDA.t141 39.4005
R5444 VDDA.n487 VDDA.t417 39.4005
R5445 VDDA.n487 VDDA.t248 39.4005
R5446 VDDA.n489 VDDA.t123 39.4005
R5447 VDDA.n489 VDDA.t37 39.4005
R5448 VDDA.n491 VDDA.t2 39.4005
R5449 VDDA.n491 VDDA.t163 39.4005
R5450 VDDA.n493 VDDA.t179 39.4005
R5451 VDDA.n493 VDDA.t152 39.4005
R5452 VDDA.n495 VDDA.t414 39.4005
R5453 VDDA.n495 VDDA.t233 39.4005
R5454 VDDA.n497 VDDA.t231 39.4005
R5455 VDDA.n497 VDDA.t33 39.4005
R5456 VDDA.n499 VDDA.t144 39.4005
R5457 VDDA.n499 VDDA.t189 39.4005
R5458 VDDA.n460 VDDA.t31 39.4005
R5459 VDDA.n460 VDDA.t119 39.4005
R5460 VDDA.n463 VDDA.t117 39.4005
R5461 VDDA.n463 VDDA.t133 39.4005
R5462 VDDA.n465 VDDA.t177 39.4005
R5463 VDDA.n465 VDDA.t47 39.4005
R5464 VDDA.n467 VDDA.t49 39.4005
R5465 VDDA.n467 VDDA.t39 39.4005
R5466 VDDA.n469 VDDA.t165 39.4005
R5467 VDDA.n469 VDDA.t433 39.4005
R5468 VDDA.n471 VDDA.t88 39.4005
R5469 VDDA.n471 VDDA.t226 39.4005
R5470 VDDA.n473 VDDA.t131 39.4005
R5471 VDDA.n473 VDDA.t90 39.4005
R5472 VDDA.n475 VDDA.t5 39.4005
R5473 VDDA.n475 VDDA.t51 39.4005
R5474 VDDA.n477 VDDA.t250 39.4005
R5475 VDDA.n477 VDDA.t41 39.4005
R5476 VDDA.n575 VDDA.t24 39.4005
R5477 VDDA.n575 VDDA.t246 39.4005
R5478 VDDA.n579 VDDA.t79 39.4005
R5479 VDDA.n579 VDDA.t11 39.4005
R5480 VDDA.n606 VDDA.t29 39.4005
R5481 VDDA.n606 VDDA.t449 39.4005
R5482 VDDA.n581 VDDA.t202 39.4005
R5483 VDDA.n581 VDDA.t445 39.4005
R5484 VDDA.n592 VDDA.t204 39.4005
R5485 VDDA.n592 VDDA.t200 39.4005
R5486 VDDA.n594 VDDA.t81 39.4005
R5487 VDDA.n594 VDDA.t61 39.4005
R5488 VDDA.n596 VDDA.t224 39.4005
R5489 VDDA.n596 VDDA.t443 39.4005
R5490 VDDA.n598 VDDA.t113 39.4005
R5491 VDDA.n598 VDDA.t111 39.4005
R5492 VDDA.n583 VDDA.t115 39.4005
R5493 VDDA.n583 VDDA.t83 39.4005
R5494 VDDA.n585 VDDA.t45 39.4005
R5495 VDDA.n585 VDDA.t431 39.4005
R5496 VDDA.n450 VDDA.n444 27.9413
R5497 VDDA.n612 VDDA.n611 27.2462
R5498 VDDA.n610 VDDA.n609 27.2462
R5499 VDDA.n590 VDDA.n589 27.2462
R5500 VDDA.n588 VDDA.n587 27.2462
R5501 VDDA.n571 VDDA.n570 25.087
R5502 VDDA.n573 VDDA.n572 25.087
R5503 VDDA.n604 VDDA.n603 25.0384
R5504 VDDA.n602 VDDA.n601 25.0384
R5505 VDDA.n524 VDDA.n523 22.9536
R5506 VDDA.n483 VDDA.n482 22.9536
R5507 VDDA.n441 VDDA.n440 22.8576
R5508 VDDA.n422 VDDA.n407 22.8576
R5509 VDDA.n386 VDDA.n385 22.8576
R5510 VDDA.n352 VDDA.n322 22.8576
R5511 VDDA.n292 VDDA.n291 22.8576
R5512 VDDA.n252 VDDA.n251 22.8576
R5513 VDDA.n233 VDDA.n219 22.8576
R5514 VDDA.n178 VDDA.n177 22.8576
R5515 VDDA.n139 VDDA.n109 22.8576
R5516 VDDA.n84 VDDA.n83 22.8576
R5517 VDDA.n44 VDDA.n43 22.8576
R5518 VDDA.n25 VDDA.n11 22.8576
R5519 VDDA.n568 VDDA.n567 22.8576
R5520 VDDA.n544 VDDA.n543 22.8576
R5521 VDDA.n391 VDDA.t191 21.8894
R5522 VDDA.n391 VDDA.t339 21.8894
R5523 VDDA.n444 VDDA.n443 20.883
R5524 VDDA.n507 VDDA.n457 20.7243
R5525 VDDA.n502 VDDA.n459 20.7243
R5526 VDDA.n479 VDDA.n462 20.7243
R5527 VDDA.n526 VDDA.n525 20.4312
R5528 VDDA.n450 VDDA.t68 19.9244
R5529 VDDA.n293 VDDA.n292 19.613
R5530 VDDA.n85 VDDA.n84 19.613
R5531 VDDA.n204 VDDA.n203 19.2005
R5532 VDDA.n202 VDDA.n201 19.2005
R5533 VDDA.n297 VDDA.n296 18.863
R5534 VDDA.n89 VDDA.n88 18.863
R5535 VDDA.n527 VDDA.n523 15.488
R5536 VDDA.n479 VDDA.n478 14.6963
R5537 VDDA.n254 VDDA.n252 14.4255
R5538 VDDA.n219 VDDA.n218 14.4255
R5539 VDDA.n46 VDDA.n44 14.4255
R5540 VDDA.n11 VDDA.n10 14.4255
R5541 VDDA.n322 VDDA.n321 14.363
R5542 VDDA.n201 VDDA.n200 14.363
R5543 VDDA.n109 VDDA.n108 14.363
R5544 VDDA.n574 VDDA.n573 14.363
R5545 VDDA.n574 VDDA.n570 14.363
R5546 VDDA.n587 VDDA.n586 14.363
R5547 VDDA.n527 VDDA.n526 14.238
R5548 VDDA.n502 VDDA.n501 14.0713
R5549 VDDA.n508 VDDA.n507 14.0713
R5550 VDDA.n484 VDDA.n483 14.0713
R5551 VDDA.n407 VDDA.n399 14.0505
R5552 VDDA.n393 VDDA.n392 14.0505
R5553 VDDA.n442 VDDA.n441 13.8005
R5554 VDDA.n397 VDDA.n396 13.8005
R5555 VDDA.n387 VDDA.n386 13.8005
R5556 VDDA.n205 VDDA.n204 13.8005
R5557 VDDA.n179 VDDA.n178 13.8005
R5558 VDDA.n543 VDDA.n542 13.8005
R5559 VDDA.n569 VDDA.n568 13.8005
R5560 VDDA.n609 VDDA.n608 13.8005
R5561 VDDA.n601 VDDA.n600 13.8005
R5562 VDDA.n591 VDDA.n590 13.8005
R5563 VDDA.n605 VDDA.n604 13.8005
R5564 VDDA.n613 VDDA.n612 13.8005
R5565 VDDA.n510 VDDA.t71 13.1338
R5566 VDDA.n510 VDDA.t167 13.1338
R5567 VDDA.n528 VDDA.t66 13.1338
R5568 VDDA.n528 VDDA.t53 13.1338
R5569 VDDA.n530 VDDA.t419 13.1338
R5570 VDDA.n530 VDDA.t421 13.1338
R5571 VDDA.n532 VDDA.t128 13.1338
R5572 VDDA.n532 VDDA.t219 13.1338
R5573 VDDA.n534 VDDA.t217 13.1338
R5574 VDDA.n534 VDDA.t57 13.1338
R5575 VDDA.n536 VDDA.t126 13.1338
R5576 VDDA.n536 VDDA.t74 13.1338
R5577 VDDA.n538 VDDA.t96 13.1338
R5578 VDDA.n538 VDDA.t208 13.1338
R5579 VDDA.n540 VDDA.t221 13.1338
R5580 VDDA.n540 VDDA.t213 13.1338
R5581 VDDA.n614 VDDA.n613 11.4105
R5582 VDDA.t361 VDDA.n420 11.2576
R5583 VDDA.n420 VDDA.t281 11.2576
R5584 VDDA.n421 VDDA.t361 11.2576
R5585 VDDA.n400 VDDA.t382 11.2576
R5586 VDDA.n258 VDDA.t289 11.2576
R5587 VDDA.n258 VDDA.t259 11.2576
R5588 VDDA.n208 VDDA.t269 11.2576
R5589 VDDA.n208 VDDA.t279 11.2576
R5590 VDDA.n217 VDDA.t265 11.2576
R5591 VDDA.n217 VDDA.t261 11.2576
R5592 VDDA.n232 VDDA.t324 11.2576
R5593 VDDA.n210 VDDA.t400 11.2576
R5594 VDDA.n253 VDDA.t271 11.2576
R5595 VDDA.n253 VDDA.t283 11.2576
R5596 VDDA.n255 VDDA.t257 11.2576
R5597 VDDA.n255 VDDA.t263 11.2576
R5598 VDDA.n50 VDDA.t253 11.2576
R5599 VDDA.n50 VDDA.t255 11.2576
R5600 VDDA.n0 VDDA.t285 11.2576
R5601 VDDA.n0 VDDA.t291 11.2576
R5602 VDDA.n9 VDDA.t277 11.2576
R5603 VDDA.n9 VDDA.t273 11.2576
R5604 VDDA.n24 VDDA.t355 11.2576
R5605 VDDA.n2 VDDA.t309 11.2576
R5606 VDDA.n45 VDDA.t287 11.2576
R5607 VDDA.n45 VDDA.t293 11.2576
R5608 VDDA.n47 VDDA.t267 11.2576
R5609 VDDA.n47 VDDA.t275 11.2576
R5610 VDDA.n296 VDDA.n294 11.2005
R5611 VDDA.n88 VDDA.n87 11.2005
R5612 VDDA.n454 VDDA.n453 11.1572
R5613 VDDA.n293 VDDA.n270 10.8443
R5614 VDDA.n85 VDDA.n62 10.8443
R5615 VDDA.n578 VDDA.n577 9.7855
R5616 VDDA.n440 VDDA.n401 9.14336
R5617 VDDA.n436 VDDA.n435 9.14336
R5618 VDDA.n433 VDDA.n430 9.14336
R5619 VDDA.n422 VDDA.n408 9.14336
R5620 VDDA.n413 VDDA.n410 9.14336
R5621 VDDA.n418 VDDA.n415 9.14336
R5622 VDDA.n381 VDDA.n356 9.14336
R5623 VDDA.n381 VDDA.n380 9.14336
R5624 VDDA.n380 VDDA.n379 9.14336
R5625 VDDA.n379 VDDA.n376 9.14336
R5626 VDDA.n376 VDDA.n375 9.14336
R5627 VDDA.n375 VDDA.n372 9.14336
R5628 VDDA.n372 VDDA.n371 9.14336
R5629 VDDA.n371 VDDA.n368 9.14336
R5630 VDDA.n368 VDDA.n367 9.14336
R5631 VDDA.n349 VDDA.n323 9.14336
R5632 VDDA.n349 VDDA.n346 9.14336
R5633 VDDA.n346 VDDA.n345 9.14336
R5634 VDDA.n345 VDDA.n342 9.14336
R5635 VDDA.n342 VDDA.n341 9.14336
R5636 VDDA.n341 VDDA.n338 9.14336
R5637 VDDA.n338 VDDA.n337 9.14336
R5638 VDDA.n337 VDDA.n334 9.14336
R5639 VDDA.n334 VDDA.n333 9.14336
R5640 VDDA.n279 VDDA.n277 9.14336
R5641 VDDA.n289 VDDA.n288 9.14336
R5642 VDDA.n251 VDDA.n211 9.14336
R5643 VDDA.n247 VDDA.n246 9.14336
R5644 VDDA.n244 VDDA.n241 9.14336
R5645 VDDA.n233 VDDA.n220 9.14336
R5646 VDDA.n225 VDDA.n222 9.14336
R5647 VDDA.n230 VDDA.n227 9.14336
R5648 VDDA.n173 VDDA.n148 9.14336
R5649 VDDA.n173 VDDA.n172 9.14336
R5650 VDDA.n172 VDDA.n171 9.14336
R5651 VDDA.n171 VDDA.n168 9.14336
R5652 VDDA.n168 VDDA.n167 9.14336
R5653 VDDA.n167 VDDA.n164 9.14336
R5654 VDDA.n164 VDDA.n163 9.14336
R5655 VDDA.n163 VDDA.n160 9.14336
R5656 VDDA.n160 VDDA.n159 9.14336
R5657 VDDA.n137 VDDA.n136 9.14336
R5658 VDDA.n136 VDDA.n135 9.14336
R5659 VDDA.n135 VDDA.n113 9.14336
R5660 VDDA.n131 VDDA.n113 9.14336
R5661 VDDA.n131 VDDA.n130 9.14336
R5662 VDDA.n130 VDDA.n118 9.14336
R5663 VDDA.n126 VDDA.n118 9.14336
R5664 VDDA.n126 VDDA.n125 9.14336
R5665 VDDA.n125 VDDA.n124 9.14336
R5666 VDDA.n69 VDDA.n67 9.14336
R5667 VDDA.n78 VDDA.n77 9.14336
R5668 VDDA.n43 VDDA.n3 9.14336
R5669 VDDA.n39 VDDA.n38 9.14336
R5670 VDDA.n36 VDDA.n33 9.14336
R5671 VDDA.n25 VDDA.n12 9.14336
R5672 VDDA.n17 VDDA.n14 9.14336
R5673 VDDA.n22 VDDA.n19 9.14336
R5674 VDDA.n561 VDDA.n556 9.14336
R5675 VDDA.n561 VDDA.n560 9.14336
R5676 VDDA.n560 VDDA.n558 9.14336
R5677 VDDA.n549 VDDA.n548 9.14336
R5678 VDDA.n548 VDDA.n547 9.14336
R5679 VDDA.n547 VDDA.n522 9.14336
R5680 VDDA.n509 VDDA.n508 8.973
R5681 VDDA.n389 VDDA.n388 8.8755
R5682 VDDA.n207 VDDA.n206 8.28175
R5683 VDDA.n389 VDDA.n259 8.15675
R5684 VDDA.n207 VDDA.n51 8.15675
R5685 VDDA.n269 VDDA.t294 8.0005
R5686 VDDA.n269 VDDA.t222 8.0005
R5687 VDDA.n267 VDDA.t158 8.0005
R5688 VDDA.n267 VDDA.t182 8.0005
R5689 VDDA.n265 VDDA.t463 8.0005
R5690 VDDA.n265 VDDA.t0 8.0005
R5691 VDDA.n263 VDDA.t450 8.0005
R5692 VDDA.n263 VDDA.t75 8.0005
R5693 VDDA.n261 VDDA.t180 8.0005
R5694 VDDA.n261 VDDA.t69 8.0005
R5695 VDDA.n260 VDDA.t129 8.0005
R5696 VDDA.n260 VDDA.t295 8.0005
R5697 VDDA.n61 VDDA.t240 8.0005
R5698 VDDA.n61 VDDA.t297 8.0005
R5699 VDDA.n59 VDDA.t108 8.0005
R5700 VDDA.n59 VDDA.t26 8.0005
R5701 VDDA.n57 VDDA.t84 8.0005
R5702 VDDA.n57 VDDA.t27 8.0005
R5703 VDDA.n55 VDDA.t76 8.0005
R5704 VDDA.n55 VDDA.t42 8.0005
R5705 VDDA.n53 VDDA.t195 8.0005
R5706 VDDA.n53 VDDA.t446 8.0005
R5707 VDDA.n52 VDDA.t296 8.0005
R5708 VDDA.n52 VDDA.t120 8.0005
R5709 VDDA.n206 VDDA.n205 6.71925
R5710 VDDA.n298 VDDA.t135 6.56717
R5711 VDDA.n298 VDDA.t211 6.56717
R5712 VDDA.n314 VDDA.t17 6.56717
R5713 VDDA.n314 VDDA.t154 6.56717
R5714 VDDA.n316 VDDA.t156 6.56717
R5715 VDDA.n316 VDDA.t428 6.56717
R5716 VDDA.n318 VDDA.t452 6.56717
R5717 VDDA.n318 VDDA.t173 6.56717
R5718 VDDA.n320 VDDA.t15 6.56717
R5719 VDDA.n320 VDDA.t454 6.56717
R5720 VDDA.n90 VDDA.t439 6.56717
R5721 VDDA.n90 VDDA.t22 6.56717
R5722 VDDA.n101 VDDA.t441 6.56717
R5723 VDDA.n101 VDDA.t7 6.56717
R5724 VDDA.n103 VDDA.t236 6.56717
R5725 VDDA.n103 VDDA.t194 6.56717
R5726 VDDA.n105 VDDA.t239 6.56717
R5727 VDDA.n105 VDDA.t198 6.56717
R5728 VDDA.n107 VDDA.t242 6.56717
R5729 VDDA.n107 VDDA.t9 6.56717
R5730 VDDA.n398 VDDA.n390 6.563
R5731 VDDA.n390 VDDA.n389 6.0005
R5732 VDDA.n390 VDDA.n207 6.0005
R5733 VDDA.n388 VDDA.n387 5.8755
R5734 VDDA.n180 VDDA.n179 5.8755
R5735 VDDA.n385 VDDA.n300 5.33286
R5736 VDDA.n352 VDDA.n351 5.33286
R5737 VDDA.n291 VDDA.n290 5.33286
R5738 VDDA.n282 VDDA.n281 5.33286
R5739 VDDA.n139 VDDA.n138 5.33286
R5740 VDDA.n177 VDDA.n92 5.33286
R5741 VDDA.n72 VDDA.n71 5.33286
R5742 VDDA.n83 VDDA.n63 5.33286
R5743 VDDA.n567 VDDA.n512 5.33286
R5744 VDDA.n545 VDDA.n544 5.33286
R5745 VDDA.n443 VDDA.n442 5.28175
R5746 VDDA.n398 VDDA.n397 5.28175
R5747 VDDA.n577 VDDA.n576 5.0005
R5748 VDDA.n454 VDDA.n450 4.5595
R5749 VDDA.n458 VDDA.n457 4.54311
R5750 VDDA.n506 VDDA.n458 4.54311
R5751 VDDA.n428 VDDA.n401 4.53698
R5752 VDDA.n435 VDDA.n434 4.53698
R5753 VDDA.n430 VDDA.n429 4.53698
R5754 VDDA.n436 VDDA.n428 4.53698
R5755 VDDA.n434 VDDA.n433 4.53698
R5756 VDDA.n409 VDDA.n408 4.53698
R5757 VDDA.n414 VDDA.n413 4.53698
R5758 VDDA.n419 VDDA.n418 4.53698
R5759 VDDA.n410 VDDA.n409 4.53698
R5760 VDDA.n415 VDDA.n414 4.53698
R5761 VDDA.n239 VDDA.n211 4.53698
R5762 VDDA.n246 VDDA.n245 4.53698
R5763 VDDA.n241 VDDA.n240 4.53698
R5764 VDDA.n247 VDDA.n239 4.53698
R5765 VDDA.n245 VDDA.n244 4.53698
R5766 VDDA.n221 VDDA.n220 4.53698
R5767 VDDA.n226 VDDA.n225 4.53698
R5768 VDDA.n231 VDDA.n230 4.53698
R5769 VDDA.n222 VDDA.n221 4.53698
R5770 VDDA.n227 VDDA.n226 4.53698
R5771 VDDA.n31 VDDA.n3 4.53698
R5772 VDDA.n38 VDDA.n37 4.53698
R5773 VDDA.n33 VDDA.n32 4.53698
R5774 VDDA.n39 VDDA.n31 4.53698
R5775 VDDA.n37 VDDA.n36 4.53698
R5776 VDDA.n13 VDDA.n12 4.53698
R5777 VDDA.n18 VDDA.n17 4.53698
R5778 VDDA.n23 VDDA.n22 4.53698
R5779 VDDA.n14 VDDA.n13 4.53698
R5780 VDDA.n19 VDDA.n18 4.53698
R5781 VDDA.n259 VDDA.n257 4.5005
R5782 VDDA.n51 VDDA.n49 4.5005
R5783 VDDA.n576 VDDA.n574 4.5005
R5784 VDDA.n504 VDDA.n459 4.48641
R5785 VDDA.n504 VDDA.n503 4.48641
R5786 VDDA.n481 VDDA.n462 4.48641
R5787 VDDA.n481 VDDA.n480 4.48641
R5788 VDDA.n452 VDDA.n451 4.12334
R5789 VDDA.n356 VDDA.n300 3.75335
R5790 VDDA.n367 VDDA.n365 3.75335
R5791 VDDA.n351 VDDA.n323 3.75335
R5792 VDDA.n333 VDDA.n331 3.75335
R5793 VDDA.n281 VDDA.n277 3.75335
R5794 VDDA.n280 VDDA.n279 3.75335
R5795 VDDA.n290 VDDA.n289 3.75335
R5796 VDDA.n288 VDDA.n287 3.75335
R5797 VDDA.n148 VDDA.n92 3.75335
R5798 VDDA.n159 VDDA.n157 3.75335
R5799 VDDA.n138 VDDA.n137 3.75335
R5800 VDDA.n124 VDDA.n123 3.75335
R5801 VDDA.n71 VDDA.n67 3.75335
R5802 VDDA.n70 VDDA.n69 3.75335
R5803 VDDA.n77 VDDA.n63 3.75335
R5804 VDDA.n79 VDDA.n78 3.75335
R5805 VDDA.n563 VDDA.n556 3.75335
R5806 VDDA.n558 VDDA.n512 3.75335
R5807 VDDA.n550 VDDA.n549 3.75335
R5808 VDDA.n545 VDDA.n522 3.75335
R5809 VDDA.n615 VDDA.n614 3.71013
R5810 VDDA.n453 VDDA.n452 3.43377
R5811 VDDA.n297 VDDA.n293 3.15675
R5812 VDDA.n89 VDDA.n85 3.15675
R5813 VDDA.n577 VDDA.n569 2.5005
R5814 VDDA.n615 VDDA.n444 2.1343
R5815 VDDA VDDA.n615 2.0779
R5816 VDDA.n501 VDDA.n484 1.8755
R5817 VDDA.n542 VDDA.n527 1.84425
R5818 VDDA.n600 VDDA.n591 1.813
R5819 VDDA.n608 VDDA.n605 1.813
R5820 VDDA.n388 VDDA.n297 1.688
R5821 VDDA.n180 VDDA.n89 1.688
R5822 VDDA.n542 VDDA.n541 1.0005
R5823 VDDA.n541 VDDA.n539 1.0005
R5824 VDDA.n539 VDDA.n537 1.0005
R5825 VDDA.n537 VDDA.n535 1.0005
R5826 VDDA.n535 VDDA.n533 1.0005
R5827 VDDA.n533 VDDA.n531 1.0005
R5828 VDDA.n531 VDDA.n529 1.0005
R5829 VDDA.n529 VDDA.n511 1.0005
R5830 VDDA.n569 VDDA.n511 1.0005
R5831 VDDA.n443 VDDA.n398 0.938
R5832 VDDA.n509 VDDA.n454 0.840625
R5833 VDDA.n578 VDDA.n509 0.74075
R5834 VDDA.n442 VDDA.n399 0.6255
R5835 VDDA.n397 VDDA.n392 0.6255
R5836 VDDA.n257 VDDA.n256 0.6255
R5837 VDDA.n256 VDDA.n254 0.6255
R5838 VDDA.n218 VDDA.n209 0.6255
R5839 VDDA.n257 VDDA.n209 0.6255
R5840 VDDA.n49 VDDA.n48 0.6255
R5841 VDDA.n48 VDDA.n46 0.6255
R5842 VDDA.n10 VDDA.n1 0.6255
R5843 VDDA.n49 VDDA.n1 0.6255
R5844 VDDA.n478 VDDA.n476 0.6255
R5845 VDDA.n476 VDDA.n474 0.6255
R5846 VDDA.n474 VDDA.n472 0.6255
R5847 VDDA.n472 VDDA.n470 0.6255
R5848 VDDA.n470 VDDA.n468 0.6255
R5849 VDDA.n468 VDDA.n466 0.6255
R5850 VDDA.n466 VDDA.n464 0.6255
R5851 VDDA.n464 VDDA.n461 0.6255
R5852 VDDA.n484 VDDA.n461 0.6255
R5853 VDDA.n501 VDDA.n500 0.6255
R5854 VDDA.n500 VDDA.n498 0.6255
R5855 VDDA.n498 VDDA.n496 0.6255
R5856 VDDA.n496 VDDA.n494 0.6255
R5857 VDDA.n494 VDDA.n492 0.6255
R5858 VDDA.n492 VDDA.n490 0.6255
R5859 VDDA.n490 VDDA.n488 0.6255
R5860 VDDA.n488 VDDA.n486 0.6255
R5861 VDDA.n486 VDDA.n456 0.6255
R5862 VDDA.n508 VDDA.n456 0.6255
R5863 VDDA.n321 VDDA.n319 0.563
R5864 VDDA.n319 VDDA.n317 0.563
R5865 VDDA.n317 VDDA.n315 0.563
R5866 VDDA.n315 VDDA.n299 0.563
R5867 VDDA.n387 VDDA.n299 0.563
R5868 VDDA.n264 VDDA.n262 0.563
R5869 VDDA.n266 VDDA.n264 0.563
R5870 VDDA.n268 VDDA.n266 0.563
R5871 VDDA.n270 VDDA.n268 0.563
R5872 VDDA.n200 VDDA.n198 0.563
R5873 VDDA.n198 VDDA.n196 0.563
R5874 VDDA.n196 VDDA.n194 0.563
R5875 VDDA.n194 VDDA.n192 0.563
R5876 VDDA.n192 VDDA.n190 0.563
R5877 VDDA.n190 VDDA.n188 0.563
R5878 VDDA.n188 VDDA.n186 0.563
R5879 VDDA.n186 VDDA.n184 0.563
R5880 VDDA.n184 VDDA.n182 0.563
R5881 VDDA.n205 VDDA.n182 0.563
R5882 VDDA.n108 VDDA.n106 0.563
R5883 VDDA.n106 VDDA.n104 0.563
R5884 VDDA.n104 VDDA.n102 0.563
R5885 VDDA.n102 VDDA.n91 0.563
R5886 VDDA.n179 VDDA.n91 0.563
R5887 VDDA.n56 VDDA.n54 0.563
R5888 VDDA.n58 VDDA.n56 0.563
R5889 VDDA.n60 VDDA.n58 0.563
R5890 VDDA.n62 VDDA.n60 0.563
R5891 VDDA.n586 VDDA.n584 0.563
R5892 VDDA.n591 VDDA.n584 0.563
R5893 VDDA.n600 VDDA.n599 0.563
R5894 VDDA.n599 VDDA.n597 0.563
R5895 VDDA.n597 VDDA.n595 0.563
R5896 VDDA.n595 VDDA.n593 0.563
R5897 VDDA.n593 VDDA.n582 0.563
R5898 VDDA.n605 VDDA.n582 0.563
R5899 VDDA.n608 VDDA.n607 0.563
R5900 VDDA.n607 VDDA.n580 0.563
R5901 VDDA.n613 VDDA.n580 0.563
R5902 VDDA.n206 VDDA.n180 0.46925
R5903 VDDA VDDA.n578 0.41175
R5904 VDDA.t209 VDDA.t67 0.1603
R5905 VDDA.t101 VDDA.t422 0.1603
R5906 VDDA.t168 VDDA.t169 0.1603
R5907 VDDA.t72 VDDA.t98 0.1603
R5908 VDDA.t55 VDDA.t214 0.1603
R5909 VDDA.n446 VDDA.t215 0.159278
R5910 VDDA.n447 VDDA.t99 0.159278
R5911 VDDA.n448 VDDA.t171 0.159278
R5912 VDDA.n449 VDDA.t97 0.159278
R5913 VDDA.n449 VDDA.t54 0.1368
R5914 VDDA.n449 VDDA.t209 0.1368
R5915 VDDA.n448 VDDA.t170 0.1368
R5916 VDDA.n448 VDDA.t101 0.1368
R5917 VDDA.n447 VDDA.t124 0.1368
R5918 VDDA.n447 VDDA.t168 0.1368
R5919 VDDA.n446 VDDA.t206 0.1368
R5920 VDDA.n446 VDDA.t72 0.1368
R5921 VDDA.n445 VDDA.t100 0.1368
R5922 VDDA.n445 VDDA.t55 0.1368
R5923 VDDA.n614 VDDA 0.135625
R5924 VDDA.t215 VDDA.n445 0.00152174
R5925 VDDA.t99 VDDA.n446 0.00152174
R5926 VDDA.t171 VDDA.n447 0.00152174
R5927 VDDA.t97 VDDA.n448 0.00152174
R5928 VDDA.t68 VDDA.n449 0.00152174
R5929 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 369.534
R5930 bgr_0.V_TOP.n23 bgr_0.V_TOP.n21 339.961
R5931 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 339.272
R5932 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 339.272
R5933 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 339.272
R5934 bgr_0.V_TOP.n29 bgr_0.V_TOP.n28 339.272
R5935 bgr_0.V_TOP.n24 bgr_0.V_TOP.n20 334.772
R5936 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 224.934
R5937 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 224.934
R5938 bgr_0.V_TOP.n37 bgr_0.V_TOP.n36 224.934
R5939 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 224.934
R5940 bgr_0.V_TOP.n35 bgr_0.V_TOP.n34 224.934
R5941 bgr_0.V_TOP.n34 bgr_0.V_TOP.n33 224.934
R5942 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 224.934
R5943 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R5944 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R5945 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R5946 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R5947 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R5948 bgr_0.V_TOP bgr_0.V_TOP.t48 214.222
R5949 bgr_0.V_TOP.n31 bgr_0.V_TOP.n30 163.175
R5950 bgr_0.V_TOP.n39 bgr_0.V_TOP.t24 144.601
R5951 bgr_0.V_TOP.n38 bgr_0.V_TOP.t33 144.601
R5952 bgr_0.V_TOP.n37 bgr_0.V_TOP.t39 144.601
R5953 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 144.601
R5954 bgr_0.V_TOP.n35 bgr_0.V_TOP.t15 144.601
R5955 bgr_0.V_TOP.n34 bgr_0.V_TOP.t28 144.601
R5956 bgr_0.V_TOP.n33 bgr_0.V_TOP.t38 144.601
R5957 bgr_0.V_TOP.n32 bgr_0.V_TOP.t14 144.601
R5958 bgr_0.V_TOP.n0 bgr_0.V_TOP.t30 144.601
R5959 bgr_0.V_TOP.n1 bgr_0.V_TOP.t18 144.601
R5960 bgr_0.V_TOP.n2 bgr_0.V_TOP.t46 144.601
R5961 bgr_0.V_TOP.n3 bgr_0.V_TOP.t37 144.601
R5962 bgr_0.V_TOP.n4 bgr_0.V_TOP.t26 144.601
R5963 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R5964 bgr_0.V_TOP.n17 bgr_0.V_TOP.t13 108.424
R5965 bgr_0.V_TOP.n30 bgr_0.V_TOP.t8 95.4467
R5966 bgr_0.V_TOP bgr_0.V_TOP.n39 69.6227
R5967 bgr_0.V_TOP.n32 bgr_0.V_TOP.n31 69.6227
R5968 bgr_0.V_TOP.n31 bgr_0.V_TOP.n5 69.6227
R5969 bgr_0.V_TOP.n18 bgr_0.V_TOP.t9 39.4005
R5970 bgr_0.V_TOP.n18 bgr_0.V_TOP.t7 39.4005
R5971 bgr_0.V_TOP.n20 bgr_0.V_TOP.t2 39.4005
R5972 bgr_0.V_TOP.n20 bgr_0.V_TOP.t1 39.4005
R5973 bgr_0.V_TOP.n22 bgr_0.V_TOP.t6 39.4005
R5974 bgr_0.V_TOP.n22 bgr_0.V_TOP.t12 39.4005
R5975 bgr_0.V_TOP.n21 bgr_0.V_TOP.t11 39.4005
R5976 bgr_0.V_TOP.n21 bgr_0.V_TOP.t3 39.4005
R5977 bgr_0.V_TOP.n26 bgr_0.V_TOP.t0 39.4005
R5978 bgr_0.V_TOP.n26 bgr_0.V_TOP.t5 39.4005
R5979 bgr_0.V_TOP.n28 bgr_0.V_TOP.t4 39.4005
R5980 bgr_0.V_TOP.n28 bgr_0.V_TOP.t10 39.4005
R5981 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 37.1479
R5982 bgr_0.V_TOP.n19 bgr_0.V_TOP.n17 27.8371
R5983 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 8.313
R5984 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 5.188
R5985 bgr_0.V_TOP.n6 bgr_0.V_TOP.t31 4.8295
R5986 bgr_0.V_TOP.n7 bgr_0.V_TOP.t22 4.8295
R5987 bgr_0.V_TOP.n8 bgr_0.V_TOP.t20 4.8295
R5988 bgr_0.V_TOP.n9 bgr_0.V_TOP.t45 4.8295
R5989 bgr_0.V_TOP.n10 bgr_0.V_TOP.t42 4.8295
R5990 bgr_0.V_TOP.n11 bgr_0.V_TOP.t36 4.8295
R5991 bgr_0.V_TOP.n12 bgr_0.V_TOP.t17 4.8295
R5992 bgr_0.V_TOP.n13 bgr_0.V_TOP.t43 4.8295
R5993 bgr_0.V_TOP.n14 bgr_0.V_TOP.t34 4.8295
R5994 bgr_0.V_TOP.n6 bgr_0.V_TOP.t35 4.5005
R5995 bgr_0.V_TOP.n7 bgr_0.V_TOP.t32 4.5005
R5996 bgr_0.V_TOP.n8 bgr_0.V_TOP.t25 4.5005
R5997 bgr_0.V_TOP.n9 bgr_0.V_TOP.t21 4.5005
R5998 bgr_0.V_TOP.n10 bgr_0.V_TOP.t49 4.5005
R5999 bgr_0.V_TOP.n11 bgr_0.V_TOP.t44 4.5005
R6000 bgr_0.V_TOP.n12 bgr_0.V_TOP.t23 4.5005
R6001 bgr_0.V_TOP.n13 bgr_0.V_TOP.t19 4.5005
R6002 bgr_0.V_TOP.n16 bgr_0.V_TOP.t40 4.5005
R6003 bgr_0.V_TOP.n15 bgr_0.V_TOP.t47 4.5005
R6004 bgr_0.V_TOP.n14 bgr_0.V_TOP.t41 4.5005
R6005 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 4.5005
R6006 bgr_0.V_TOP.n29 bgr_0.V_TOP.n27 2.1255
R6007 bgr_0.V_TOP.n27 bgr_0.V_TOP.n25 2.1255
R6008 bgr_0.V_TOP.n25 bgr_0.V_TOP.n19 2.1255
R6009 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 0.3295
R6010 bgr_0.V_TOP.n9 bgr_0.V_TOP.n8 0.3295
R6011 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 0.3295
R6012 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 0.3295
R6013 bgr_0.V_TOP.n16 bgr_0.V_TOP.n15 0.3295
R6014 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 0.3295
R6015 bgr_0.V_TOP.n9 bgr_0.V_TOP.n7 0.2825
R6016 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 0.2825
R6017 bgr_0.V_TOP.n13 bgr_0.V_TOP.n11 0.2825
R6018 bgr_0.V_TOP.n14 bgr_0.V_TOP.n13 0.2825
R6019 VOUT-.n8 VOUT-.n0 149.19
R6020 VOUT-.n3 VOUT-.n1 149.19
R6021 VOUT-.n7 VOUT-.n6 148.626
R6022 VOUT-.n5 VOUT-.n4 148.626
R6023 VOUT-.n3 VOUT-.n2 148.626
R6024 VOUT-.n10 VOUT-.n9 144.126
R6025 VOUT-.n91 VOUT-.t17 112.184
R6026 VOUT-.n88 VOUT-.n86 98.9303
R6027 VOUT-.n90 VOUT-.n89 97.8053
R6028 VOUT-.n88 VOUT-.n87 97.8053
R6029 VOUT-.n85 VOUT-.n10 15.5682
R6030 VOUT-.n85 VOUT-.n84 11.5649
R6031 VOUT- VOUT-.n85 9.46925
R6032 VOUT-.n9 VOUT-.t1 6.56717
R6033 VOUT-.n9 VOUT-.t8 6.56717
R6034 VOUT-.n6 VOUT-.t6 6.56717
R6035 VOUT-.n6 VOUT-.t7 6.56717
R6036 VOUT-.n4 VOUT-.t5 6.56717
R6037 VOUT-.n4 VOUT-.t16 6.56717
R6038 VOUT-.n2 VOUT-.t0 6.56717
R6039 VOUT-.n2 VOUT-.t15 6.56717
R6040 VOUT-.n1 VOUT-.t2 6.56717
R6041 VOUT-.n1 VOUT-.t14 6.56717
R6042 VOUT-.n0 VOUT-.t13 6.56717
R6043 VOUT-.n0 VOUT-.t9 6.56717
R6044 VOUT-.n39 VOUT-.t68 4.8295
R6045 VOUT-.n47 VOUT-.t66 4.8295
R6046 VOUT-.n45 VOUT-.t115 4.8295
R6047 VOUT-.n43 VOUT-.t150 4.8295
R6048 VOUT-.n42 VOUT-.t132 4.8295
R6049 VOUT-.n41 VOUT-.t29 4.8295
R6050 VOUT-.n59 VOUT-.t125 4.8295
R6051 VOUT-.n60 VOUT-.t73 4.8295
R6052 VOUT-.n61 VOUT-.t23 4.8295
R6053 VOUT-.n62 VOUT-.t109 4.8295
R6054 VOUT-.n63 VOUT-.t76 4.8295
R6055 VOUT-.n64 VOUT-.t44 4.8295
R6056 VOUT-.n66 VOUT-.t37 4.8295
R6057 VOUT-.n67 VOUT-.t143 4.8295
R6058 VOUT-.n69 VOUT-.t70 4.8295
R6059 VOUT-.n70 VOUT-.t39 4.8295
R6060 VOUT-.n72 VOUT-.t32 4.8295
R6061 VOUT-.n73 VOUT-.t138 4.8295
R6062 VOUT-.n75 VOUT-.t131 4.8295
R6063 VOUT-.n76 VOUT-.t101 4.8295
R6064 VOUT-.n78 VOUT-.t28 4.8295
R6065 VOUT-.n79 VOUT-.t133 4.8295
R6066 VOUT-.n11 VOUT-.t26 4.8295
R6067 VOUT-.n13 VOUT-.t36 4.8295
R6068 VOUT-.n24 VOUT-.t140 4.8295
R6069 VOUT-.n25 VOUT-.t111 4.8295
R6070 VOUT-.n27 VOUT-.t41 4.8295
R6071 VOUT-.n28 VOUT-.t151 4.8295
R6072 VOUT-.n30 VOUT-.t80 4.8295
R6073 VOUT-.n31 VOUT-.t51 4.8295
R6074 VOUT-.n33 VOUT-.t49 4.8295
R6075 VOUT-.n34 VOUT-.t19 4.8295
R6076 VOUT-.n36 VOUT-.t85 4.8295
R6077 VOUT-.n37 VOUT-.t55 4.8295
R6078 VOUT-.n81 VOUT-.t124 4.8295
R6079 VOUT-.n49 VOUT-.t91 4.8154
R6080 VOUT-.n50 VOUT-.t69 4.8154
R6081 VOUT-.n51 VOUT-.t107 4.8154
R6082 VOUT-.n49 VOUT-.t31 4.806
R6083 VOUT-.n50 VOUT-.t149 4.806
R6084 VOUT-.n51 VOUT-.t50 4.806
R6085 VOUT-.n52 VOUT-.t144 4.806
R6086 VOUT-.n52 VOUT-.t83 4.806
R6087 VOUT-.n53 VOUT-.t120 4.806
R6088 VOUT-.n54 VOUT-.t104 4.806
R6089 VOUT-.n55 VOUT-.t137 4.806
R6090 VOUT-.n56 VOUT-.t35 4.806
R6091 VOUT-.n57 VOUT-.t156 4.806
R6092 VOUT-.n14 VOUT-.t71 4.806
R6093 VOUT-.n14 VOUT-.t113 4.806
R6094 VOUT-.n15 VOUT-.t114 4.806
R6095 VOUT-.n15 VOUT-.t24 4.806
R6096 VOUT-.n16 VOUT-.t65 4.806
R6097 VOUT-.n16 VOUT-.t62 4.806
R6098 VOUT-.n17 VOUT-.t154 4.806
R6099 VOUT-.n17 VOUT-.t95 4.806
R6100 VOUT-.n18 VOUT-.t105 4.806
R6101 VOUT-.n18 VOUT-.t126 4.806
R6102 VOUT-.n19 VOUT-.t141 4.806
R6103 VOUT-.n19 VOUT-.t38 4.806
R6104 VOUT-.n20 VOUT-.t92 4.806
R6105 VOUT-.n20 VOUT-.t74 4.806
R6106 VOUT-.n21 VOUT-.t42 4.806
R6107 VOUT-.n22 VOUT-.t82 4.806
R6108 VOUT-.n39 VOUT-.t86 4.5005
R6109 VOUT-.n40 VOUT-.t54 4.5005
R6110 VOUT-.n47 VOUT-.t77 4.5005
R6111 VOUT-.n48 VOUT-.t43 4.5005
R6112 VOUT-.n45 VOUT-.t58 4.5005
R6113 VOUT-.n46 VOUT-.t22 4.5005
R6114 VOUT-.n43 VOUT-.t94 4.5005
R6115 VOUT-.n44 VOUT-.t61 4.5005
R6116 VOUT-.n42 VOUT-.t99 4.5005
R6117 VOUT-.n41 VOUT-.t52 4.5005
R6118 VOUT-.n58 VOUT-.t155 4.5005
R6119 VOUT-.n57 VOUT-.t116 4.5005
R6120 VOUT-.n56 VOUT-.t136 4.5005
R6121 VOUT-.n55 VOUT-.t100 4.5005
R6122 VOUT-.n54 VOUT-.t64 4.5005
R6123 VOUT-.n53 VOUT-.t81 4.5005
R6124 VOUT-.n52 VOUT-.t45 4.5005
R6125 VOUT-.n51 VOUT-.t146 4.5005
R6126 VOUT-.n50 VOUT-.t108 4.5005
R6127 VOUT-.n49 VOUT-.t130 4.5005
R6128 VOUT-.n59 VOUT-.t152 4.5005
R6129 VOUT-.n60 VOUT-.t112 4.5005
R6130 VOUT-.n61 VOUT-.t47 4.5005
R6131 VOUT-.n62 VOUT-.t147 4.5005
R6132 VOUT-.n63 VOUT-.t27 4.5005
R6133 VOUT-.n65 VOUT-.t128 4.5005
R6134 VOUT-.n64 VOUT-.t97 4.5005
R6135 VOUT-.n66 VOUT-.t123 4.5005
R6136 VOUT-.n68 VOUT-.t88 4.5005
R6137 VOUT-.n67 VOUT-.t57 4.5005
R6138 VOUT-.n69 VOUT-.t20 4.5005
R6139 VOUT-.n71 VOUT-.t121 4.5005
R6140 VOUT-.n70 VOUT-.t87 4.5005
R6141 VOUT-.n72 VOUT-.t118 4.5005
R6142 VOUT-.n74 VOUT-.t84 4.5005
R6143 VOUT-.n73 VOUT-.t53 4.5005
R6144 VOUT-.n75 VOUT-.t79 4.5005
R6145 VOUT-.n77 VOUT-.t48 4.5005
R6146 VOUT-.n76 VOUT-.t153 4.5005
R6147 VOUT-.n78 VOUT-.t117 4.5005
R6148 VOUT-.n80 VOUT-.t78 4.5005
R6149 VOUT-.n79 VOUT-.t46 4.5005
R6150 VOUT-.n11 VOUT-.t119 4.5005
R6151 VOUT-.n12 VOUT-.t33 4.5005
R6152 VOUT-.n13 VOUT-.t122 4.5005
R6153 VOUT-.n23 VOUT-.t90 4.5005
R6154 VOUT-.n22 VOUT-.t56 4.5005
R6155 VOUT-.n21 VOUT-.t142 4.5005
R6156 VOUT-.n20 VOUT-.t110 4.5005
R6157 VOUT-.n19 VOUT-.t72 4.5005
R6158 VOUT-.n18 VOUT-.t25 4.5005
R6159 VOUT-.n17 VOUT-.t127 4.5005
R6160 VOUT-.n16 VOUT-.t93 4.5005
R6161 VOUT-.n15 VOUT-.t60 4.5005
R6162 VOUT-.n14 VOUT-.t148 4.5005
R6163 VOUT-.n24 VOUT-.t89 4.5005
R6164 VOUT-.n26 VOUT-.t59 4.5005
R6165 VOUT-.n25 VOUT-.t21 4.5005
R6166 VOUT-.n27 VOUT-.t129 4.5005
R6167 VOUT-.n29 VOUT-.t98 4.5005
R6168 VOUT-.n28 VOUT-.t63 4.5005
R6169 VOUT-.n30 VOUT-.t30 4.5005
R6170 VOUT-.n32 VOUT-.t134 4.5005
R6171 VOUT-.n31 VOUT-.t103 4.5005
R6172 VOUT-.n33 VOUT-.t135 4.5005
R6173 VOUT-.n35 VOUT-.t102 4.5005
R6174 VOUT-.n34 VOUT-.t67 4.5005
R6175 VOUT-.n36 VOUT-.t34 4.5005
R6176 VOUT-.n38 VOUT-.t139 4.5005
R6177 VOUT-.n37 VOUT-.t106 4.5005
R6178 VOUT-.n81 VOUT-.t75 4.5005
R6179 VOUT-.n82 VOUT-.t40 4.5005
R6180 VOUT-.n83 VOUT-.t145 4.5005
R6181 VOUT-.n84 VOUT-.t96 4.5005
R6182 VOUT-.n10 VOUT-.n8 4.5005
R6183 VOUT-.n89 VOUT-.t12 3.42907
R6184 VOUT-.n89 VOUT-.t3 3.42907
R6185 VOUT-.n87 VOUT-.t10 3.42907
R6186 VOUT-.n87 VOUT-.t18 3.42907
R6187 VOUT-.n86 VOUT-.t4 3.42907
R6188 VOUT-.n86 VOUT-.t11 3.42907
R6189 VOUT-.n91 VOUT-.n90 1.30519
R6190 VOUT- VOUT-.n91 1.24269
R6191 VOUT-.n90 VOUT-.n88 1.1255
R6192 VOUT-.n5 VOUT-.n3 0.563
R6193 VOUT-.n7 VOUT-.n5 0.563
R6194 VOUT-.n8 VOUT-.n7 0.563
R6195 VOUT-.n40 VOUT-.n39 0.3295
R6196 VOUT-.n48 VOUT-.n47 0.3295
R6197 VOUT-.n46 VOUT-.n45 0.3295
R6198 VOUT-.n44 VOUT-.n43 0.3295
R6199 VOUT-.n58 VOUT-.n41 0.3295
R6200 VOUT-.n58 VOUT-.n57 0.3295
R6201 VOUT-.n57 VOUT-.n56 0.3295
R6202 VOUT-.n56 VOUT-.n55 0.3295
R6203 VOUT-.n55 VOUT-.n54 0.3295
R6204 VOUT-.n54 VOUT-.n53 0.3295
R6205 VOUT-.n53 VOUT-.n52 0.3295
R6206 VOUT-.n52 VOUT-.n51 0.3295
R6207 VOUT-.n51 VOUT-.n50 0.3295
R6208 VOUT-.n50 VOUT-.n49 0.3295
R6209 VOUT-.n60 VOUT-.n59 0.3295
R6210 VOUT-.n62 VOUT-.n61 0.3295
R6211 VOUT-.n65 VOUT-.n63 0.3295
R6212 VOUT-.n65 VOUT-.n64 0.3295
R6213 VOUT-.n68 VOUT-.n66 0.3295
R6214 VOUT-.n68 VOUT-.n67 0.3295
R6215 VOUT-.n71 VOUT-.n69 0.3295
R6216 VOUT-.n71 VOUT-.n70 0.3295
R6217 VOUT-.n74 VOUT-.n72 0.3295
R6218 VOUT-.n74 VOUT-.n73 0.3295
R6219 VOUT-.n77 VOUT-.n75 0.3295
R6220 VOUT-.n77 VOUT-.n76 0.3295
R6221 VOUT-.n80 VOUT-.n78 0.3295
R6222 VOUT-.n80 VOUT-.n79 0.3295
R6223 VOUT-.n12 VOUT-.n11 0.3295
R6224 VOUT-.n23 VOUT-.n13 0.3295
R6225 VOUT-.n23 VOUT-.n22 0.3295
R6226 VOUT-.n22 VOUT-.n21 0.3295
R6227 VOUT-.n21 VOUT-.n20 0.3295
R6228 VOUT-.n20 VOUT-.n19 0.3295
R6229 VOUT-.n19 VOUT-.n18 0.3295
R6230 VOUT-.n18 VOUT-.n17 0.3295
R6231 VOUT-.n17 VOUT-.n16 0.3295
R6232 VOUT-.n16 VOUT-.n15 0.3295
R6233 VOUT-.n15 VOUT-.n14 0.3295
R6234 VOUT-.n26 VOUT-.n24 0.3295
R6235 VOUT-.n26 VOUT-.n25 0.3295
R6236 VOUT-.n29 VOUT-.n27 0.3295
R6237 VOUT-.n29 VOUT-.n28 0.3295
R6238 VOUT-.n32 VOUT-.n30 0.3295
R6239 VOUT-.n32 VOUT-.n31 0.3295
R6240 VOUT-.n35 VOUT-.n33 0.3295
R6241 VOUT-.n35 VOUT-.n34 0.3295
R6242 VOUT-.n38 VOUT-.n36 0.3295
R6243 VOUT-.n38 VOUT-.n37 0.3295
R6244 VOUT-.n82 VOUT-.n81 0.3295
R6245 VOUT-.n83 VOUT-.n82 0.3295
R6246 VOUT-.n84 VOUT-.n83 0.3295
R6247 VOUT-.n53 VOUT-.n48 0.306
R6248 VOUT-.n54 VOUT-.n46 0.306
R6249 VOUT-.n55 VOUT-.n44 0.306
R6250 VOUT-.n56 VOUT-.n42 0.306
R6251 VOUT-.n58 VOUT-.n40 0.2825
R6252 VOUT-.n60 VOUT-.n58 0.2825
R6253 VOUT-.n62 VOUT-.n60 0.2825
R6254 VOUT-.n65 VOUT-.n62 0.2825
R6255 VOUT-.n68 VOUT-.n65 0.2825
R6256 VOUT-.n71 VOUT-.n68 0.2825
R6257 VOUT-.n74 VOUT-.n71 0.2825
R6258 VOUT-.n77 VOUT-.n74 0.2825
R6259 VOUT-.n80 VOUT-.n77 0.2825
R6260 VOUT-.n23 VOUT-.n12 0.2825
R6261 VOUT-.n26 VOUT-.n23 0.2825
R6262 VOUT-.n29 VOUT-.n26 0.2825
R6263 VOUT-.n32 VOUT-.n29 0.2825
R6264 VOUT-.n35 VOUT-.n32 0.2825
R6265 VOUT-.n38 VOUT-.n35 0.2825
R6266 VOUT-.n82 VOUT-.n38 0.2825
R6267 VOUT-.n82 VOUT-.n80 0.2825
R6268 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.197
R6269 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.87
R6270 two_stage_opamp_dummy_magic_0.cap_res_X.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R6271 two_stage_opamp_dummy_magic_0.cap_res_X.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R6272 two_stage_opamp_dummy_magic_0.cap_res_X.t11 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R6273 two_stage_opamp_dummy_magic_0.cap_res_X.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R6274 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R6275 two_stage_opamp_dummy_magic_0.cap_res_X.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.1603
R6276 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R6277 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1603
R6278 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.1603
R6279 two_stage_opamp_dummy_magic_0.cap_res_X.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.1603
R6280 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R6281 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R6282 two_stage_opamp_dummy_magic_0.cap_res_X.t5 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R6283 two_stage_opamp_dummy_magic_0.cap_res_X.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R6284 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R6285 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R6286 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R6287 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1603
R6288 two_stage_opamp_dummy_magic_0.cap_res_X.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1603
R6289 two_stage_opamp_dummy_magic_0.cap_res_X.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1603
R6290 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R6291 two_stage_opamp_dummy_magic_0.cap_res_X.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R6292 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.1603
R6293 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R6294 two_stage_opamp_dummy_magic_0.cap_res_X.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1603
R6295 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R6296 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.1603
R6297 two_stage_opamp_dummy_magic_0.cap_res_X.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.1603
R6298 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.1603
R6299 two_stage_opamp_dummy_magic_0.cap_res_X.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.1603
R6300 two_stage_opamp_dummy_magic_0.cap_res_X.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1603
R6301 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1603
R6302 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.1603
R6303 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1603
R6304 two_stage_opamp_dummy_magic_0.cap_res_X.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1603
R6305 two_stage_opamp_dummy_magic_0.cap_res_X.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R6306 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.1603
R6307 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.1603
R6308 two_stage_opamp_dummy_magic_0.cap_res_X.t9 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R6309 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.1603
R6310 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1603
R6311 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1603
R6312 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.1603
R6313 two_stage_opamp_dummy_magic_0.cap_res_X.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1603
R6314 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1603
R6315 two_stage_opamp_dummy_magic_0.cap_res_X.t15 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1603
R6316 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.1603
R6317 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R6318 two_stage_opamp_dummy_magic_0.cap_res_X.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R6319 two_stage_opamp_dummy_magic_0.cap_res_X.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.1603
R6320 two_stage_opamp_dummy_magic_0.cap_res_X.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R6321 two_stage_opamp_dummy_magic_0.cap_res_X.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1603
R6322 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.1603
R6323 two_stage_opamp_dummy_magic_0.cap_res_X.t7 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1603
R6324 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.159278
R6325 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.159278
R6326 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.159278
R6327 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.159278
R6328 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.159278
R6329 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.159278
R6330 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.159278
R6331 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.159278
R6332 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.159278
R6333 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.159278
R6334 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.159278
R6335 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.159278
R6336 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.159278
R6337 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.159278
R6338 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.159278
R6339 two_stage_opamp_dummy_magic_0.cap_res_X.t98 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.159278
R6340 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.159278
R6341 two_stage_opamp_dummy_magic_0.cap_res_X.t23 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.159278
R6342 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.159278
R6343 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.159278
R6344 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R6345 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R6346 two_stage_opamp_dummy_magic_0.cap_res_X.t109 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R6347 two_stage_opamp_dummy_magic_0.cap_res_X.t73 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R6348 two_stage_opamp_dummy_magic_0.cap_res_X.t36 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R6349 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R6350 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R6351 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R6352 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R6353 two_stage_opamp_dummy_magic_0.cap_res_X.t2 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R6354 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.159278
R6355 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.159278
R6356 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.159278
R6357 two_stage_opamp_dummy_magic_0.cap_res_X.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.137822
R6358 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R6359 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1368
R6360 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1368
R6361 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1368
R6362 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1368
R6363 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.1368
R6364 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.1368
R6365 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1368
R6366 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.1368
R6367 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.1368
R6368 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1368
R6369 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.1368
R6370 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1368
R6371 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.1368
R6372 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R6373 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1368
R6374 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1368
R6375 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.1368
R6376 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.1368
R6377 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1368
R6378 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1368
R6379 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1368
R6380 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R6381 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1368
R6382 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R6383 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.1368
R6384 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1368
R6385 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1368
R6386 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R6387 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1368
R6388 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.1368
R6389 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.1133
R6390 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.1133
R6391 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.1133
R6392 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R6393 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R6394 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R6395 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R6396 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R6397 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R6398 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R6399 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R6400 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R6401 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R6402 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R6403 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.1133
R6404 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.1133
R6405 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.1133
R6406 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R6407 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.00152174
R6408 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.00152174
R6409 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.00152174
R6410 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.00152174
R6411 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.00152174
R6412 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.00152174
R6413 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.00152174
R6414 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.00152174
R6415 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.00152174
R6416 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R6417 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R6418 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.00152174
R6419 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R6420 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.00152174
R6421 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.00152174
R6422 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.00152174
R6423 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.00152174
R6424 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.00152174
R6425 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.00152174
R6426 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.00152174
R6427 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.00152174
R6428 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R6429 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.00152174
R6430 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.00152174
R6431 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.00152174
R6432 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.00152174
R6433 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.00152174
R6434 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.00152174
R6435 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R6436 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.00152174
R6437 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.00152174
R6438 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.00152174
R6439 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.00152174
R6440 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.00152174
R6441 two_stage_opamp_dummy_magic_0.cap_res_X.t57 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.00152174
R6442 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 631.202
R6443 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 629.952
R6444 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 625.452
R6445 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 289.2
R6446 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 289.2
R6447 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 227.002
R6448 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 212.733
R6449 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 212.733
R6450 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 176.733
R6451 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 176.733
R6452 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 176.733
R6453 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 176.733
R6454 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 176.733
R6455 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 152
R6456 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 152
R6457 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 112.468
R6458 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 112.468
R6459 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R6460 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R6461 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 112.468
R6462 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 112.468
R6463 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R6464 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 112.468
R6465 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 78.8005
R6466 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 78.8005
R6467 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 78.8005
R6468 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 78.8005
R6469 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 78.8005
R6470 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 78.8005
R6471 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 48.0005
R6472 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 48.0005
R6473 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 48.0005
R6474 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 48.0005
R6475 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 48.0005
R6476 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 48.0005
R6477 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 45.5227
R6478 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 45.5227
R6479 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 45.5227
R6480 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 45.5227
R6481 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 15.2693
R6482 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 14.0193
R6483 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 5.7505
R6484 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 4.938
R6485 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 0.8755
R6486 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R6487 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R6488 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t12 449.868
R6489 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t16 449.868
R6490 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R6491 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R6492 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R6493 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R6494 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R6495 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R6496 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R6497 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R6498 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t18 273.134
R6499 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R6500 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t21 273.134
R6501 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R6502 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R6503 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R6504 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R6505 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t14 273.134
R6506 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R6507 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R6508 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 176.733
R6509 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R6510 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R6511 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R6512 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R6513 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.n15 176.733
R6514 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 176.733
R6515 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R6516 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R6517 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R6518 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R6519 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.n6 176.733
R6520 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t2 175.553
R6521 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n12 172.207
R6522 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.n21 165.8
R6523 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t1 62.3283
R6524 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 54.6272
R6525 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n16 54.6272
R6526 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n11 54.6272
R6527 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.n7 54.6272
R6528 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 43.0005
R6529 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t3 39.4005
R6530 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R6531 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R6532 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R6533 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n3 22.5312
R6534 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 12.1255
R6535 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 6.92238
R6536 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t51 1172.87
R6537 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t27 1172.87
R6538 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.t48 996.134
R6539 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.t35 996.134
R6540 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t42 996.134
R6541 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t34 996.134
R6542 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t43 996.134
R6543 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t29 996.134
R6544 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t45 996.134
R6545 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t31 996.134
R6546 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t26 690.867
R6547 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.t32 690.867
R6548 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t39 530.201
R6549 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t44 530.201
R6550 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t40 514.134
R6551 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t46 514.134
R6552 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t41 514.134
R6553 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t25 514.134
R6554 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t38 514.134
R6555 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t52 514.134
R6556 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t36 514.134
R6557 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.t49 514.134
R6558 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.t54 353.467
R6559 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t28 353.467
R6560 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t53 353.467
R6561 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t30 353.467
R6562 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t47 353.467
R6563 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t33 353.467
R6564 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t50 353.467
R6565 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6566 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 176.733
R6567 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n48 176.733
R6568 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.n47 176.733
R6569 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R6570 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R6571 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R6572 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 176.733
R6573 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 176.733
R6574 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 176.733
R6575 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.n23 176.733
R6576 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6577 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6578 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6579 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R6580 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.n31 176.733
R6581 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 176.733
R6582 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6583 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6584 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 166.258
R6585 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.n11 163.626
R6586 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 163.001
R6587 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 163.001
R6588 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 163.001
R6589 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.n12 163.001
R6590 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n30 161.541
R6591 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 161.541
R6592 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n20 158.501
R6593 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n0 117.888
R6594 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 117.326
R6595 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 117.326
R6596 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 117.326
R6597 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 117.326
R6598 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.n1 117.326
R6599 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 54.6272
R6600 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n26 54.6272
R6601 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 54.6272
R6602 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n35 54.6272
R6603 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 53.3126
R6604 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n46 53.3126
R6605 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.X.n52 50.3023
R6606 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n21 16.8755
R6607 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t20 16.0005
R6608 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.t16 16.0005
R6609 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t11 16.0005
R6610 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t13 16.0005
R6611 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R6612 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t12 16.0005
R6613 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R6614 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t9 16.0005
R6615 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t10 16.0005
R6616 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t8 16.0005
R6617 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R6618 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R6619 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.n40 13.4693
R6620 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t3 11.2576
R6621 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R6622 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t4 11.2576
R6623 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R6624 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R6625 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R6626 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t24 11.2576
R6627 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t22 11.2576
R6628 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t18 11.2576
R6629 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t23 11.2576
R6630 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R6631 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t19 11.2576
R6632 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.n19 5.1255
R6633 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 4.5005
R6634 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n42 2.59425
R6635 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n10 1.8755
R6636 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n13 0.6255
R6637 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n15 0.6255
R6638 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n17 0.6255
R6639 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 0.563
R6640 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.563
R6641 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.563
R6642 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n8 0.563
R6643 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n9 146.47
R6644 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 146.47
R6645 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 145.906
R6646 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 145.906
R6647 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n7 145.906
R6648 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 145.906
R6649 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 114.719
R6650 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.n18 114.719
R6651 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 114.156
R6652 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 114.156
R6653 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R6654 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R6655 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R6656 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R6657 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R6658 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R6659 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R6660 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R6661 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R6662 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R6663 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R6664 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R6665 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R6666 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R6667 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R6668 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R6669 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R6670 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R6671 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R6672 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R6673 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R6674 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R6675 two_stage_opamp_dummy_magic_0.VD1.t13 two_stage_opamp_dummy_magic_0.VD1.n19 16.0005
R6676 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.n14 5.24008
R6677 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 4.5005
R6678 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.563
R6679 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R6680 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n2 0.563
R6681 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 0.563
R6682 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 0.234875
R6683 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n8 0.234875
R6684 VOUT+.n8 VOUT+.n6 149.19
R6685 VOUT+.n14 VOUT+.n13 149.19
R6686 VOUT+.n12 VOUT+.n11 148.626
R6687 VOUT+.n10 VOUT+.n9 148.626
R6688 VOUT+.n8 VOUT+.n7 148.626
R6689 VOUT+.n16 VOUT+.n15 144.126
R6690 VOUT+.n5 VOUT+.t5 112.184
R6691 VOUT+.n2 VOUT+.n0 98.9303
R6692 VOUT+.n4 VOUT+.n3 97.8053
R6693 VOUT+.n2 VOUT+.n1 97.8053
R6694 VOUT+.n91 VOUT+.n16 15.5682
R6695 VOUT+.n91 VOUT+.n90 11.5649
R6696 VOUT+ VOUT+.n91 9.2505
R6697 VOUT+.n15 VOUT+.t8 6.56717
R6698 VOUT+.n15 VOUT+.t0 6.56717
R6699 VOUT+.n13 VOUT+.t18 6.56717
R6700 VOUT+.n13 VOUT+.t15 6.56717
R6701 VOUT+.n11 VOUT+.t16 6.56717
R6702 VOUT+.n11 VOUT+.t17 6.56717
R6703 VOUT+.n9 VOUT+.t6 6.56717
R6704 VOUT+.n9 VOUT+.t7 6.56717
R6705 VOUT+.n7 VOUT+.t11 6.56717
R6706 VOUT+.n7 VOUT+.t1 6.56717
R6707 VOUT+.n6 VOUT+.t14 6.56717
R6708 VOUT+.n6 VOUT+.t4 6.56717
R6709 VOUT+.n45 VOUT+.t56 4.8295
R6710 VOUT+.n47 VOUT+.t105 4.8295
R6711 VOUT+.n48 VOUT+.t29 4.8295
R6712 VOUT+.n50 VOUT+.t60 4.8295
R6713 VOUT+.n52 VOUT+.t115 4.8295
R6714 VOUT+.n63 VOUT+.t20 4.8295
R6715 VOUT+.n66 VOUT+.t31 4.8295
R6716 VOUT+.n65 VOUT+.t121 4.8295
R6717 VOUT+.n68 VOUT+.t67 4.8295
R6718 VOUT+.n67 VOUT+.t152 4.8295
R6719 VOUT+.n69 VOUT+.t131 4.8295
R6720 VOUT+.n70 VOUT+.t118 4.8295
R6721 VOUT+.n72 VOUT+.t89 4.8295
R6722 VOUT+.n73 VOUT+.t76 4.8295
R6723 VOUT+.n75 VOUT+.t127 4.8295
R6724 VOUT+.n76 VOUT+.t110 4.8295
R6725 VOUT+.n78 VOUT+.t84 4.8295
R6726 VOUT+.n79 VOUT+.t68 4.8295
R6727 VOUT+.n81 VOUT+.t42 4.8295
R6728 VOUT+.n82 VOUT+.t30 4.8295
R6729 VOUT+.n84 VOUT+.t81 4.8295
R6730 VOUT+.n85 VOUT+.t64 4.8295
R6731 VOUT+.n17 VOUT+.t150 4.8295
R6732 VOUT+.n28 VOUT+.t75 4.8295
R6733 VOUT+.n30 VOUT+.t54 4.8295
R6734 VOUT+.n31 VOUT+.t34 4.8295
R6735 VOUT+.n33 VOUT+.t95 4.8295
R6736 VOUT+.n34 VOUT+.t79 4.8295
R6737 VOUT+.n36 VOUT+.t134 4.8295
R6738 VOUT+.n37 VOUT+.t122 4.8295
R6739 VOUT+.n39 VOUT+.t102 4.8295
R6740 VOUT+.n40 VOUT+.t82 4.8295
R6741 VOUT+.n42 VOUT+.t137 4.8295
R6742 VOUT+.n43 VOUT+.t126 4.8295
R6743 VOUT+.n87 VOUT+.t28 4.8295
R6744 VOUT+.n56 VOUT+.t57 4.8154
R6745 VOUT+.n55 VOUT+.t33 4.8154
R6746 VOUT+.n54 VOUT+.t77 4.8154
R6747 VOUT+.n62 VOUT+.t116 4.806
R6748 VOUT+.n61 VOUT+.t147 4.806
R6749 VOUT+.n60 VOUT+.t43 4.806
R6750 VOUT+.n59 VOUT+.t83 4.806
R6751 VOUT+.n58 VOUT+.t63 4.806
R6752 VOUT+.n57 VOUT+.t26 4.806
R6753 VOUT+.n57 VOUT+.t103 4.806
R6754 VOUT+.n56 VOUT+.t135 4.806
R6755 VOUT+.n55 VOUT+.t120 4.806
R6756 VOUT+.n54 VOUT+.t155 4.806
R6757 VOUT+.n27 VOUT+.t91 4.806
R6758 VOUT+.n26 VOUT+.t38 4.806
R6759 VOUT+.n25 VOUT+.t130 4.806
R6760 VOUT+.n25 VOUT+.t90 4.806
R6761 VOUT+.n24 VOUT+.t80 4.806
R6762 VOUT+.n24 VOUT+.t128 4.806
R6763 VOUT+.n23 VOUT+.t124 4.806
R6764 VOUT+.n23 VOUT+.t32 4.806
R6765 VOUT+.n22 VOUT+.t70 4.806
R6766 VOUT+.n22 VOUT+.t73 4.806
R6767 VOUT+.n21 VOUT+.t23 4.806
R6768 VOUT+.n21 VOUT+.t108 4.806
R6769 VOUT+.n20 VOUT+.t62 4.806
R6770 VOUT+.n20 VOUT+.t19 4.806
R6771 VOUT+.n19 VOUT+.t151 4.806
R6772 VOUT+.n19 VOUT+.t49 4.806
R6773 VOUT+.n46 VOUT+.t132 4.5005
R6774 VOUT+.n45 VOUT+.t96 4.5005
R6775 VOUT+.n47 VOUT+.t69 4.5005
R6776 VOUT+.n48 VOUT+.t139 4.5005
R6777 VOUT+.n49 VOUT+.t109 4.5005
R6778 VOUT+.n50 VOUT+.t37 4.5005
R6779 VOUT+.n51 VOUT+.t144 4.5005
R6780 VOUT+.n52 VOUT+.t21 4.5005
R6781 VOUT+.n53 VOUT+.t125 4.5005
R6782 VOUT+.n54 VOUT+.t119 4.5005
R6783 VOUT+.n55 VOUT+.t78 4.5005
R6784 VOUT+.n56 VOUT+.t97 4.5005
R6785 VOUT+.n57 VOUT+.t61 4.5005
R6786 VOUT+.n58 VOUT+.t27 4.5005
R6787 VOUT+.n59 VOUT+.t41 4.5005
R6788 VOUT+.n60 VOUT+.t145 4.5005
R6789 VOUT+.n61 VOUT+.t113 4.5005
R6790 VOUT+.n62 VOUT+.t72 4.5005
R6791 VOUT+.n64 VOUT+.t92 4.5005
R6792 VOUT+.n63 VOUT+.t55 4.5005
R6793 VOUT+.n66 VOUT+.t50 4.5005
R6794 VOUT+.n65 VOUT+.t156 4.5005
R6795 VOUT+.n68 VOUT+.t86 4.5005
R6796 VOUT+.n67 VOUT+.t47 4.5005
R6797 VOUT+.n69 VOUT+.t94 4.5005
R6798 VOUT+.n71 VOUT+.t39 4.5005
R6799 VOUT+.n70 VOUT+.t146 4.5005
R6800 VOUT+.n72 VOUT+.t53 4.5005
R6801 VOUT+.n74 VOUT+.t142 4.5005
R6802 VOUT+.n73 VOUT+.t112 4.5005
R6803 VOUT+.n75 VOUT+.t88 4.5005
R6804 VOUT+.n77 VOUT+.t35 4.5005
R6805 VOUT+.n76 VOUT+.t140 4.5005
R6806 VOUT+.n78 VOUT+.t46 4.5005
R6807 VOUT+.n80 VOUT+.t136 4.5005
R6808 VOUT+.n79 VOUT+.t104 4.5005
R6809 VOUT+.n81 VOUT+.t149 4.5005
R6810 VOUT+.n83 VOUT+.t99 4.5005
R6811 VOUT+.n82 VOUT+.t65 4.5005
R6812 VOUT+.n84 VOUT+.t40 4.5005
R6813 VOUT+.n86 VOUT+.t133 4.5005
R6814 VOUT+.n85 VOUT+.t98 4.5005
R6815 VOUT+.n18 VOUT+.t45 4.5005
R6816 VOUT+.n17 VOUT+.t101 4.5005
R6817 VOUT+.n19 VOUT+.t85 4.5005
R6818 VOUT+.n20 VOUT+.t48 4.5005
R6819 VOUT+.n21 VOUT+.t138 4.5005
R6820 VOUT+.n22 VOUT+.t107 4.5005
R6821 VOUT+.n23 VOUT+.t71 4.5005
R6822 VOUT+.n24 VOUT+.t25 4.5005
R6823 VOUT+.n25 VOUT+.t129 4.5005
R6824 VOUT+.n26 VOUT+.t87 4.5005
R6825 VOUT+.n27 VOUT+.t52 4.5005
R6826 VOUT+.n29 VOUT+.t141 4.5005
R6827 VOUT+.n28 VOUT+.t111 4.5005
R6828 VOUT+.n30 VOUT+.t24 4.5005
R6829 VOUT+.n32 VOUT+.t114 4.5005
R6830 VOUT+.n31 VOUT+.t74 4.5005
R6831 VOUT+.n33 VOUT+.t59 4.5005
R6832 VOUT+.n35 VOUT+.t148 4.5005
R6833 VOUT+.n34 VOUT+.t117 4.5005
R6834 VOUT+.n36 VOUT+.t100 4.5005
R6835 VOUT+.n38 VOUT+.t44 4.5005
R6836 VOUT+.n37 VOUT+.t153 4.5005
R6837 VOUT+.n39 VOUT+.t66 4.5005
R6838 VOUT+.n41 VOUT+.t154 4.5005
R6839 VOUT+.n40 VOUT+.t123 4.5005
R6840 VOUT+.n42 VOUT+.t106 4.5005
R6841 VOUT+.n44 VOUT+.t51 4.5005
R6842 VOUT+.n43 VOUT+.t22 4.5005
R6843 VOUT+.n90 VOUT+.t36 4.5005
R6844 VOUT+.n89 VOUT+.t143 4.5005
R6845 VOUT+.n88 VOUT+.t93 4.5005
R6846 VOUT+.n87 VOUT+.t58 4.5005
R6847 VOUT+.n16 VOUT+.n14 4.5005
R6848 VOUT+.n3 VOUT+.t2 3.42907
R6849 VOUT+.n3 VOUT+.t12 3.42907
R6850 VOUT+.n1 VOUT+.t3 3.42907
R6851 VOUT+.n1 VOUT+.t10 3.42907
R6852 VOUT+.n0 VOUT+.t13 3.42907
R6853 VOUT+.n0 VOUT+.t9 3.42907
R6854 VOUT+ VOUT+.n5 1.46144
R6855 VOUT+.n5 VOUT+.n4 1.30519
R6856 VOUT+.n4 VOUT+.n2 1.1255
R6857 VOUT+.n10 VOUT+.n8 0.563
R6858 VOUT+.n12 VOUT+.n10 0.563
R6859 VOUT+.n14 VOUT+.n12 0.563
R6860 VOUT+.n46 VOUT+.n45 0.3295
R6861 VOUT+.n49 VOUT+.n48 0.3295
R6862 VOUT+.n51 VOUT+.n50 0.3295
R6863 VOUT+.n53 VOUT+.n52 0.3295
R6864 VOUT+.n55 VOUT+.n54 0.3295
R6865 VOUT+.n56 VOUT+.n55 0.3295
R6866 VOUT+.n57 VOUT+.n56 0.3295
R6867 VOUT+.n58 VOUT+.n57 0.3295
R6868 VOUT+.n59 VOUT+.n58 0.3295
R6869 VOUT+.n60 VOUT+.n59 0.3295
R6870 VOUT+.n61 VOUT+.n60 0.3295
R6871 VOUT+.n62 VOUT+.n61 0.3295
R6872 VOUT+.n64 VOUT+.n62 0.3295
R6873 VOUT+.n64 VOUT+.n63 0.3295
R6874 VOUT+.n66 VOUT+.n65 0.3295
R6875 VOUT+.n68 VOUT+.n67 0.3295
R6876 VOUT+.n71 VOUT+.n69 0.3295
R6877 VOUT+.n71 VOUT+.n70 0.3295
R6878 VOUT+.n74 VOUT+.n72 0.3295
R6879 VOUT+.n74 VOUT+.n73 0.3295
R6880 VOUT+.n77 VOUT+.n75 0.3295
R6881 VOUT+.n77 VOUT+.n76 0.3295
R6882 VOUT+.n80 VOUT+.n78 0.3295
R6883 VOUT+.n80 VOUT+.n79 0.3295
R6884 VOUT+.n83 VOUT+.n81 0.3295
R6885 VOUT+.n83 VOUT+.n82 0.3295
R6886 VOUT+.n86 VOUT+.n84 0.3295
R6887 VOUT+.n86 VOUT+.n85 0.3295
R6888 VOUT+.n18 VOUT+.n17 0.3295
R6889 VOUT+.n20 VOUT+.n19 0.3295
R6890 VOUT+.n21 VOUT+.n20 0.3295
R6891 VOUT+.n22 VOUT+.n21 0.3295
R6892 VOUT+.n23 VOUT+.n22 0.3295
R6893 VOUT+.n24 VOUT+.n23 0.3295
R6894 VOUT+.n25 VOUT+.n24 0.3295
R6895 VOUT+.n26 VOUT+.n25 0.3295
R6896 VOUT+.n27 VOUT+.n26 0.3295
R6897 VOUT+.n29 VOUT+.n27 0.3295
R6898 VOUT+.n29 VOUT+.n28 0.3295
R6899 VOUT+.n32 VOUT+.n30 0.3295
R6900 VOUT+.n32 VOUT+.n31 0.3295
R6901 VOUT+.n35 VOUT+.n33 0.3295
R6902 VOUT+.n35 VOUT+.n34 0.3295
R6903 VOUT+.n38 VOUT+.n36 0.3295
R6904 VOUT+.n38 VOUT+.n37 0.3295
R6905 VOUT+.n41 VOUT+.n39 0.3295
R6906 VOUT+.n41 VOUT+.n40 0.3295
R6907 VOUT+.n44 VOUT+.n42 0.3295
R6908 VOUT+.n44 VOUT+.n43 0.3295
R6909 VOUT+.n90 VOUT+.n89 0.3295
R6910 VOUT+.n89 VOUT+.n88 0.3295
R6911 VOUT+.n88 VOUT+.n87 0.3295
R6912 VOUT+.n61 VOUT+.n47 0.306
R6913 VOUT+.n60 VOUT+.n49 0.306
R6914 VOUT+.n59 VOUT+.n51 0.306
R6915 VOUT+.n58 VOUT+.n53 0.306
R6916 VOUT+.n64 VOUT+.n46 0.2825
R6917 VOUT+.n66 VOUT+.n64 0.2825
R6918 VOUT+.n68 VOUT+.n66 0.2825
R6919 VOUT+.n71 VOUT+.n68 0.2825
R6920 VOUT+.n74 VOUT+.n71 0.2825
R6921 VOUT+.n77 VOUT+.n74 0.2825
R6922 VOUT+.n80 VOUT+.n77 0.2825
R6923 VOUT+.n83 VOUT+.n80 0.2825
R6924 VOUT+.n86 VOUT+.n83 0.2825
R6925 VOUT+.n29 VOUT+.n18 0.2825
R6926 VOUT+.n32 VOUT+.n29 0.2825
R6927 VOUT+.n35 VOUT+.n32 0.2825
R6928 VOUT+.n38 VOUT+.n35 0.2825
R6929 VOUT+.n41 VOUT+.n38 0.2825
R6930 VOUT+.n44 VOUT+.n41 0.2825
R6931 VOUT+.n88 VOUT+.n44 0.2825
R6932 VOUT+.n88 VOUT+.n86 0.2825
R6933 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 50.3211
R6934 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R6935 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R6936 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1603
R6937 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1603
R6938 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R6939 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1603
R6940 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.1603
R6941 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1603
R6942 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1603
R6943 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1603
R6944 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R6945 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1603
R6946 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1603
R6947 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R6948 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R6949 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R6950 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1603
R6951 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R6952 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1603
R6953 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1603
R6954 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.1603
R6955 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R6956 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1603
R6957 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.1603
R6958 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1603
R6959 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1603
R6960 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1603
R6961 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.1603
R6962 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.1603
R6963 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1603
R6964 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R6965 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1603
R6966 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R6967 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.1603
R6968 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1603
R6969 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1603
R6970 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1603
R6971 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1603
R6972 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.1603
R6973 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R6974 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R6975 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R6976 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1603
R6977 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1603
R6978 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1603
R6979 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1603
R6980 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R6981 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.1603
R6982 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R6983 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R6984 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R6985 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R6986 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R6987 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.1603
R6988 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.159278
R6989 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.159278
R6990 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.159278
R6991 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.159278
R6992 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.159278
R6993 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.159278
R6994 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.159278
R6995 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.159278
R6996 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R6997 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R6998 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R6999 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7000 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7001 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7002 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7003 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7004 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7005 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7006 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.159278
R7007 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.159278
R7008 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.159278
R7009 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.159278
R7010 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.159278
R7011 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.159278
R7012 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.159278
R7013 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.159278
R7014 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.159278
R7015 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.159278
R7016 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.159278
R7017 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.159278
R7018 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.159278
R7019 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.159278
R7020 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.159278
R7021 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.137822
R7022 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.1368
R7023 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.1368
R7024 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.1368
R7025 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.1368
R7026 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1368
R7027 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1368
R7028 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.1368
R7029 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.1368
R7030 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1368
R7031 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.1368
R7032 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.1368
R7033 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1368
R7034 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.1368
R7035 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1368
R7036 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1368
R7037 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.1368
R7038 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7039 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1368
R7040 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1368
R7041 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1368
R7042 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1368
R7043 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1368
R7044 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1368
R7045 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1368
R7046 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R7047 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1368
R7048 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1368
R7049 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1368
R7050 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1368
R7051 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.1368
R7052 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1368
R7053 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7054 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7055 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7056 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.1133
R7057 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.1133
R7058 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.1133
R7059 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.1133
R7060 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.1133
R7061 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.1133
R7062 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7063 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7064 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7065 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7066 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7067 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7068 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7069 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7070 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7071 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.00152174
R7072 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.00152174
R7073 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R7074 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.00152174
R7075 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.00152174
R7076 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.00152174
R7077 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.00152174
R7078 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.00152174
R7079 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.00152174
R7080 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.00152174
R7081 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.00152174
R7082 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.00152174
R7083 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.00152174
R7084 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.00152174
R7085 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.00152174
R7086 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R7087 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.00152174
R7088 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.00152174
R7089 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.00152174
R7090 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.00152174
R7091 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.00152174
R7092 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.00152174
R7093 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.00152174
R7094 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.00152174
R7095 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.00152174
R7096 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.00152174
R7097 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.00152174
R7098 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R7099 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R7100 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.00152174
R7101 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R7102 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.00152174
R7103 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.00152174
R7104 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.00152174
R7105 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.00152174
R7106 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 144.827
R7107 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 134.577
R7108 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 118.986
R7109 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 100.6
R7110 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 100.038
R7111 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 100.038
R7112 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 100.038
R7113 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 100.038
R7114 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 43.284
R7115 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 37.4067
R7116 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 24.0005
R7117 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 24.0005
R7118 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 24.0005
R7119 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R7120 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R7121 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 8.0005
R7122 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R7123 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 8.0005
R7124 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R7125 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R7126 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R7127 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 8.0005
R7128 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R7129 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R7130 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 5.6255
R7131 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 0.563
R7132 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 0.563
R7133 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 0.563
R7134 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 0.047375
R7135 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 525.38
R7136 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 525.38
R7137 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 358.288
R7138 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 358.288
R7139 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 281.168
R7140 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 281.168
R7141 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 281.168
R7142 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 281.168
R7143 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7144 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7145 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.05
R7146 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.05
R7147 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 116.038
R7148 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 116.038
R7149 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 77.1205
R7150 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 77.1205
R7151 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 18.0005
R7152 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 688.859
R7153 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 514.134
R7154 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 321.024
R7155 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 320.229
R7156 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 274.716
R7157 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 274.716
R7158 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 245.82
R7159 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 245.82
R7160 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 245.018
R7161 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 245.018
R7162 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 214.056
R7163 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 197.939
R7164 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 197.939
R7165 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 174.726
R7166 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 174.726
R7167 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 174.726
R7168 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 174.726
R7169 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 173.591
R7170 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 169.216
R7171 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 169.216
R7172 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 128.534
R7173 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 128.534
R7174 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 125.736
R7175 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 123.573
R7176 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 123.573
R7177 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 112.468
R7178 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 112.468
R7179 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 44.3599
R7180 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R7181 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R7182 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R7183 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R7184 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R7185 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R7186 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 10.0317
R7187 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 4.3755
R7188 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 3.89425
R7189 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 3.03175
R7190 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 1.88487
R7191 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 1.28175
R7192 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 1.28175
R7193 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 0.79425
R7194 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7195 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7196 bgr_0.Vin+.n0 bgr_0.Vin+.t8 303.259
R7197 bgr_0.Vin+.n5 bgr_0.Vin+.n3 227.169
R7198 bgr_0.Vin+.n0 bgr_0.Vin+.t9 174.726
R7199 bgr_0.Vin+.n1 bgr_0.Vin+.t6 174.726
R7200 bgr_0.Vin+.n2 bgr_0.Vin+.t10 174.726
R7201 bgr_0.Vin+.n7 bgr_0.Vin+.n6 168.435
R7202 bgr_0.Vin+.n5 bgr_0.Vin+.n4 168.435
R7203 bgr_0.Vin+.n8 bgr_0.Vin+.t5 158.989
R7204 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7205 bgr_0.Vin+.t0 bgr_0.Vin+.n8 119.067
R7206 bgr_0.Vin+.n3 bgr_0.Vin+.t7 96.4005
R7207 bgr_0.Vin+.n8 bgr_0.Vin+.n7 35.0317
R7208 bgr_0.Vin+.n6 bgr_0.Vin+.t1 13.1338
R7209 bgr_0.Vin+.n6 bgr_0.Vin+.t4 13.1338
R7210 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R7211 bgr_0.Vin+.n4 bgr_0.Vin+.t2 13.1338
R7212 bgr_0.Vin+.n7 bgr_0.Vin+.n5 2.1255
R7213 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t12 652.076
R7214 two_stage_opamp_dummy_magic_0.VD3.n59 two_stage_opamp_dummy_magic_0.VD3.t15 652.076
R7215 two_stage_opamp_dummy_magic_0.VD3.n58 two_stage_opamp_dummy_magic_0.VD3.n11 585
R7216 two_stage_opamp_dummy_magic_0.VD3.n42 two_stage_opamp_dummy_magic_0.VD3.n29 585
R7217 two_stage_opamp_dummy_magic_0.VD3.n46 two_stage_opamp_dummy_magic_0.VD3.n11 290.233
R7218 two_stage_opamp_dummy_magic_0.VD3.n52 two_stage_opamp_dummy_magic_0.VD3.n11 290.233
R7219 two_stage_opamp_dummy_magic_0.VD3.n47 two_stage_opamp_dummy_magic_0.VD3.n11 290.233
R7220 two_stage_opamp_dummy_magic_0.VD3.n40 two_stage_opamp_dummy_magic_0.VD3.n29 290.233
R7221 two_stage_opamp_dummy_magic_0.VD3.n35 two_stage_opamp_dummy_magic_0.VD3.n29 290.233
R7222 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n29 290.233
R7223 two_stage_opamp_dummy_magic_0.VD3.n47 two_stage_opamp_dummy_magic_0.VD3.n15 242.903
R7224 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n18 242.903
R7225 two_stage_opamp_dummy_magic_0.VD3.n58 two_stage_opamp_dummy_magic_0.VD3.n57 238.367
R7226 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 185
R7227 two_stage_opamp_dummy_magic_0.VD3.n55 two_stage_opamp_dummy_magic_0.VD3.n54 185
R7228 two_stage_opamp_dummy_magic_0.VD3.n56 two_stage_opamp_dummy_magic_0.VD3.n55 185
R7229 two_stage_opamp_dummy_magic_0.VD3.n53 two_stage_opamp_dummy_magic_0.VD3.n45 185
R7230 two_stage_opamp_dummy_magic_0.VD3.n51 two_stage_opamp_dummy_magic_0.VD3.n50 185
R7231 two_stage_opamp_dummy_magic_0.VD3.n49 two_stage_opamp_dummy_magic_0.VD3.n48 185
R7232 two_stage_opamp_dummy_magic_0.VD3.n43 two_stage_opamp_dummy_magic_0.VD3.n42 185
R7233 two_stage_opamp_dummy_magic_0.VD3.n44 two_stage_opamp_dummy_magic_0.VD3.n43 185
R7234 two_stage_opamp_dummy_magic_0.VD3.n41 two_stage_opamp_dummy_magic_0.VD3.n19 185
R7235 two_stage_opamp_dummy_magic_0.VD3.n39 two_stage_opamp_dummy_magic_0.VD3.n38 185
R7236 two_stage_opamp_dummy_magic_0.VD3.n37 two_stage_opamp_dummy_magic_0.VD3.n36 185
R7237 two_stage_opamp_dummy_magic_0.VD3.n34 two_stage_opamp_dummy_magic_0.VD3.n33 185
R7238 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n31 185
R7239 two_stage_opamp_dummy_magic_0.VD3.n56 two_stage_opamp_dummy_magic_0.VD3.t16 170.513
R7240 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.VD3.n44 170.513
R7241 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 163.626
R7242 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 163.001
R7243 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 163.001
R7244 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n3 163.001
R7245 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 163.001
R7246 two_stage_opamp_dummy_magic_0.VD3.n62 two_stage_opamp_dummy_magic_0.VD3.n61 162.999
R7247 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n9 159.803
R7248 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 159.803
R7249 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 159.803
R7250 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 159.803
R7251 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n26 159.803
R7252 two_stage_opamp_dummy_magic_0.VD3.n55 two_stage_opamp_dummy_magic_0.VD3.n13 150
R7253 two_stage_opamp_dummy_magic_0.VD3.n55 two_stage_opamp_dummy_magic_0.VD3.n45 150
R7254 two_stage_opamp_dummy_magic_0.VD3.n50 two_stage_opamp_dummy_magic_0.VD3.n49 150
R7255 two_stage_opamp_dummy_magic_0.VD3.n43 two_stage_opamp_dummy_magic_0.VD3.n19 150
R7256 two_stage_opamp_dummy_magic_0.VD3.n38 two_stage_opamp_dummy_magic_0.VD3.n37 150
R7257 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 150
R7258 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t2 146.155
R7259 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.VD3.t4 146.155
R7260 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.t10 146.155
R7261 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t6 146.155
R7262 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.VD3.t8 146.155
R7263 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t36 146.155
R7264 two_stage_opamp_dummy_magic_0.VD3.t36 two_stage_opamp_dummy_magic_0.VD3.t32 146.155
R7265 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.VD3.t18 146.155
R7266 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.t34 146.155
R7267 two_stage_opamp_dummy_magic_0.VD3.t34 two_stage_opamp_dummy_magic_0.VD3.t0 146.155
R7268 two_stage_opamp_dummy_magic_0.VD3.t0 two_stage_opamp_dummy_magic_0.VD3.t13 146.155
R7269 two_stage_opamp_dummy_magic_0.VD3.n57 two_stage_opamp_dummy_magic_0.VD3.n56 65.8183
R7270 two_stage_opamp_dummy_magic_0.VD3.n56 two_stage_opamp_dummy_magic_0.VD3.n14 65.8183
R7271 two_stage_opamp_dummy_magic_0.VD3.n56 two_stage_opamp_dummy_magic_0.VD3.n15 65.8183
R7272 two_stage_opamp_dummy_magic_0.VD3.n44 two_stage_opamp_dummy_magic_0.VD3.n16 65.8183
R7273 two_stage_opamp_dummy_magic_0.VD3.n44 two_stage_opamp_dummy_magic_0.VD3.n17 65.8183
R7274 two_stage_opamp_dummy_magic_0.VD3.n44 two_stage_opamp_dummy_magic_0.VD3.n18 65.8183
R7275 two_stage_opamp_dummy_magic_0.VD3.n45 two_stage_opamp_dummy_magic_0.VD3.n14 53.3664
R7276 two_stage_opamp_dummy_magic_0.VD3.n49 two_stage_opamp_dummy_magic_0.VD3.n15 53.3664
R7277 two_stage_opamp_dummy_magic_0.VD3.n57 two_stage_opamp_dummy_magic_0.VD3.n13 53.3664
R7278 two_stage_opamp_dummy_magic_0.VD3.n50 two_stage_opamp_dummy_magic_0.VD3.n14 53.3664
R7279 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n16 53.3664
R7280 two_stage_opamp_dummy_magic_0.VD3.n37 two_stage_opamp_dummy_magic_0.VD3.n17 53.3664
R7281 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n18 53.3664
R7282 two_stage_opamp_dummy_magic_0.VD3.n38 two_stage_opamp_dummy_magic_0.VD3.n16 53.3664
R7283 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n17 53.3664
R7284 two_stage_opamp_dummy_magic_0.VD3.n59 two_stage_opamp_dummy_magic_0.VD3.n58 22.8576
R7285 two_stage_opamp_dummy_magic_0.VD3.n42 two_stage_opamp_dummy_magic_0.VD3.n28 22.8576
R7286 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.n27 14.4255
R7287 two_stage_opamp_dummy_magic_0.VD3.n60 two_stage_opamp_dummy_magic_0.VD3.n59 13.8005
R7288 two_stage_opamp_dummy_magic_0.VD3.n61 two_stage_opamp_dummy_magic_0.VD3.n60 13.688
R7289 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R7290 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R7291 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R7292 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R7293 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R7294 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R7295 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t33 11.2576
R7296 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t19 11.2576
R7297 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t35 11.2576
R7298 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R7299 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R7300 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t14 11.2576
R7301 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R7302 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t27 11.2576
R7303 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R7304 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R7305 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t28 11.2576
R7306 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R7307 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R7308 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t26 11.2576
R7309 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R7310 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t25 11.2576
R7311 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.VD3.n62 11.2576
R7312 two_stage_opamp_dummy_magic_0.VD3.n62 two_stage_opamp_dummy_magic_0.VD3.t30 11.2576
R7313 two_stage_opamp_dummy_magic_0.VD3.n58 two_stage_opamp_dummy_magic_0.VD3.n12 9.14336
R7314 two_stage_opamp_dummy_magic_0.VD3.n54 two_stage_opamp_dummy_magic_0.VD3.n53 9.14336
R7315 two_stage_opamp_dummy_magic_0.VD3.n51 two_stage_opamp_dummy_magic_0.VD3.n48 9.14336
R7316 two_stage_opamp_dummy_magic_0.VD3.n42 two_stage_opamp_dummy_magic_0.VD3.n41 9.14336
R7317 two_stage_opamp_dummy_magic_0.VD3.n39 two_stage_opamp_dummy_magic_0.VD3.n36 9.14336
R7318 two_stage_opamp_dummy_magic_0.VD3.n34 two_stage_opamp_dummy_magic_0.VD3.n31 9.14336
R7319 two_stage_opamp_dummy_magic_0.VD3.n46 two_stage_opamp_dummy_magic_0.VD3.n12 4.53698
R7320 two_stage_opamp_dummy_magic_0.VD3.n53 two_stage_opamp_dummy_magic_0.VD3.n52 4.53698
R7321 two_stage_opamp_dummy_magic_0.VD3.n48 two_stage_opamp_dummy_magic_0.VD3.n47 4.53698
R7322 two_stage_opamp_dummy_magic_0.VD3.n54 two_stage_opamp_dummy_magic_0.VD3.n46 4.53698
R7323 two_stage_opamp_dummy_magic_0.VD3.n52 two_stage_opamp_dummy_magic_0.VD3.n51 4.53698
R7324 two_stage_opamp_dummy_magic_0.VD3.n41 two_stage_opamp_dummy_magic_0.VD3.n40 4.53698
R7325 two_stage_opamp_dummy_magic_0.VD3.n36 two_stage_opamp_dummy_magic_0.VD3.n35 4.53698
R7326 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 4.53698
R7327 two_stage_opamp_dummy_magic_0.VD3.n40 two_stage_opamp_dummy_magic_0.VD3.n39 4.53698
R7328 two_stage_opamp_dummy_magic_0.VD3.n35 two_stage_opamp_dummy_magic_0.VD3.n34 4.53698
R7329 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n25 0.6255
R7330 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n23 0.6255
R7331 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n21 0.6255
R7332 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n10 0.6255
R7333 two_stage_opamp_dummy_magic_0.VD3.n60 two_stage_opamp_dummy_magic_0.VD3.n10 0.6255
R7334 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R7335 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R7336 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n6 0.6255
R7337 two_stage_opamp_dummy_magic_0.VD3.n61 two_stage_opamp_dummy_magic_0.VD3.n8 0.6255
R7338 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7339 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7340 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7341 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 310.488
R7342 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7343 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7344 bgr_0.V_mir1.n7 bgr_0.V_mir1.t12 278.312
R7345 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7346 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7347 bgr_0.V_mir1.n18 bgr_0.V_mir1.t6 184.097
R7348 bgr_0.V_mir1.n11 bgr_0.V_mir1.t2 184.097
R7349 bgr_0.V_mir1.n2 bgr_0.V_mir1.t0 184.097
R7350 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7351 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7352 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7353 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7354 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7355 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7356 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 120.501
R7357 bgr_0.V_mir1.n17 bgr_0.V_mir1.t10 120.501
R7358 bgr_0.V_mir1.n9 bgr_0.V_mir1.t17 120.501
R7359 bgr_0.V_mir1.n10 bgr_0.V_mir1.t8 120.501
R7360 bgr_0.V_mir1.n0 bgr_0.V_mir1.t18 120.501
R7361 bgr_0.V_mir1.n1 bgr_0.V_mir1.t4 120.501
R7362 bgr_0.V_mir1.n6 bgr_0.V_mir1.t14 48.0005
R7363 bgr_0.V_mir1.n6 bgr_0.V_mir1.t13 48.0005
R7364 bgr_0.V_mir1.n5 bgr_0.V_mir1.t15 48.0005
R7365 bgr_0.V_mir1.n5 bgr_0.V_mir1.t16 48.0005
R7366 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7367 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7368 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7369 bgr_0.V_mir1.n12 bgr_0.V_mir1.t3 39.4005
R7370 bgr_0.V_mir1.n12 bgr_0.V_mir1.t9 39.4005
R7371 bgr_0.V_mir1.n3 bgr_0.V_mir1.t1 39.4005
R7372 bgr_0.V_mir1.n3 bgr_0.V_mir1.t5 39.4005
R7373 bgr_0.V_mir1.n20 bgr_0.V_mir1.t7 39.4005
R7374 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7375 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7376 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7377 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7378 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7379 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7380 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7381 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t13 354.854
R7382 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t21 346.8
R7383 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n19 339.522
R7384 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 339.522
R7385 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n14 335.022
R7386 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t8 275.909
R7387 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.n10 227.909
R7388 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n12 222.034
R7389 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t22 184.097
R7390 bgr_0.1st_Vout_1.n17 bgr_0.1st_Vout_1.t32 184.097
R7391 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t16 184.097
R7392 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t36 184.097
R7393 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n17 166.05
R7394 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n8 166.05
R7395 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.n4 54.2759
R7396 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t9 48.0005
R7397 bgr_0.1st_Vout_1.n12 bgr_0.1st_Vout_1.t10 48.0005
R7398 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t6 48.0005
R7399 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t7 48.0005
R7400 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t4 39.4005
R7401 bgr_0.1st_Vout_1.n19 bgr_0.1st_Vout_1.t2 39.4005
R7402 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t0 39.4005
R7403 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 39.4005
R7404 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t5 39.4005
R7405 bgr_0.1st_Vout_1.n14 bgr_0.1st_Vout_1.t1 39.4005
R7406 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t11 4.8295
R7407 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t29 4.8295
R7408 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t31 4.8295
R7409 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R7410 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.8295
R7411 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t14 4.8295
R7412 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t30 4.8295
R7413 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t18 4.8295
R7414 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t23 4.8295
R7415 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t15 4.5005
R7416 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t35 4.5005
R7417 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t34 4.5005
R7418 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t28 4.5005
R7419 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t27 4.5005
R7420 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t19 4.5005
R7421 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t33 4.5005
R7422 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t26 4.5005
R7423 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.t25 4.5005
R7424 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t17 4.5005
R7425 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t12 4.5005
R7426 bgr_0.1st_Vout_1.n13 bgr_0.1st_Vout_1.n11 4.5005
R7427 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n15 4.5005
R7428 bgr_0.1st_Vout_1.n20 bgr_0.1st_Vout_1.n18 1.3755
R7429 bgr_0.1st_Vout_1.n16 bgr_0.1st_Vout_1.n9 1.3755
R7430 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n5 1.188
R7431 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n2 0.8935
R7432 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n0 0.8935
R7433 bgr_0.1st_Vout_1.n15 bgr_0.1st_Vout_1.n13 0.78175
R7434 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.n3 0.6585
R7435 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 0.6585
R7436 bgr_0.1st_Vout_1.n18 bgr_0.1st_Vout_1.n16 0.6255
R7437 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.n7 0.6255
R7438 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n20 0.438
R7439 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t33 355.293
R7440 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t34 346.8
R7441 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n10 339.522
R7442 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n8 339.522
R7443 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.n3 335.022
R7444 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t4 275.909
R7445 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.n5 227.909
R7446 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n7 222.034
R7447 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t16 184.097
R7448 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t27 184.097
R7449 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t13 184.097
R7450 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.t24 184.097
R7451 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n11 166.05
R7452 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n9 166.05
R7453 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n4 52.9634
R7454 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t1 48.0005
R7455 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t2 48.0005
R7456 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t5 48.0005
R7457 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t3 48.0005
R7458 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t10 39.4005
R7459 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t8 39.4005
R7460 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t7 39.4005
R7461 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t9 39.4005
R7462 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t6 39.4005
R7463 bgr_0.1st_Vout_2.t0 bgr_0.1st_Vout_2.n12 39.4005
R7464 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n1 5.28175
R7465 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.n0 5.188
R7466 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t17 4.8295
R7467 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t35 4.8295
R7468 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t11 4.8295
R7469 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t26 4.8295
R7470 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t30 4.8295
R7471 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t19 4.8295
R7472 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t36 4.8295
R7473 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.8295
R7474 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t18 4.8295
R7475 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t12 4.5005
R7476 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t32 4.5005
R7477 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R7478 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t23 4.5005
R7479 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t22 4.5005
R7480 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t15 4.5005
R7481 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t29 4.5005
R7482 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t21 4.5005
R7483 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t28 4.5005
R7484 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R7485 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t14 4.5005
R7486 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.n6 4.5005
R7487 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 3.1025
R7488 bgr_0.cap_res2.t20 bgr_0.cap_res2.t17 121.245
R7489 bgr_0.cap_res2.t12 bgr_0.cap_res2.t6 0.1603
R7490 bgr_0.cap_res2.t5 bgr_0.cap_res2.t0 0.1603
R7491 bgr_0.cap_res2.t10 bgr_0.cap_res2.t4 0.1603
R7492 bgr_0.cap_res2.t3 bgr_0.cap_res2.t19 0.1603
R7493 bgr_0.cap_res2.t18 bgr_0.cap_res2.t15 0.1603
R7494 bgr_0.cap_res2.n1 bgr_0.cap_res2.t2 0.159278
R7495 bgr_0.cap_res2.n2 bgr_0.cap_res2.t9 0.159278
R7496 bgr_0.cap_res2.n3 bgr_0.cap_res2.t16 0.159278
R7497 bgr_0.cap_res2.n4 bgr_0.cap_res2.t11 0.159278
R7498 bgr_0.cap_res2.n4 bgr_0.cap_res2.t14 0.1368
R7499 bgr_0.cap_res2.n4 bgr_0.cap_res2.t12 0.1368
R7500 bgr_0.cap_res2.n3 bgr_0.cap_res2.t8 0.1368
R7501 bgr_0.cap_res2.n3 bgr_0.cap_res2.t5 0.1368
R7502 bgr_0.cap_res2.n2 bgr_0.cap_res2.t13 0.1368
R7503 bgr_0.cap_res2.n2 bgr_0.cap_res2.t10 0.1368
R7504 bgr_0.cap_res2.n1 bgr_0.cap_res2.t7 0.1368
R7505 bgr_0.cap_res2.n1 bgr_0.cap_res2.t3 0.1368
R7506 bgr_0.cap_res2.n0 bgr_0.cap_res2.t1 0.1368
R7507 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R7508 bgr_0.cap_res2.t2 bgr_0.cap_res2.n0 0.00152174
R7509 bgr_0.cap_res2.t9 bgr_0.cap_res2.n1 0.00152174
R7510 bgr_0.cap_res2.t16 bgr_0.cap_res2.n2 0.00152174
R7511 bgr_0.cap_res2.t11 bgr_0.cap_res2.n3 0.00152174
R7512 bgr_0.cap_res2.t17 bgr_0.cap_res2.n4 0.00152174
R7513 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t31 650.273
R7514 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t9 650.273
R7515 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t12 611.739
R7516 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R7517 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t13 611.739
R7518 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t23 611.739
R7519 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.t27 445.423
R7520 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R7521 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t24 421.75
R7522 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t28 421.75
R7523 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R7524 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R7525 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t19 421.75
R7526 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R7527 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t32 421.75
R7528 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t18 421.75
R7529 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R7530 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R7531 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R7532 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t16 421.75
R7533 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R7534 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R7535 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R7536 two_stage_opamp_dummy_magic_0.Vb2.n30 two_stage_opamp_dummy_magic_0.Vb2.n17 169.352
R7537 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R7538 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.n5 167.094
R7539 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R7540 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 167.094
R7541 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.n1 167.094
R7542 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R7543 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R7544 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.n14 167.094
R7545 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R7546 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 167.094
R7547 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.n10 167.094
R7548 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R7549 two_stage_opamp_dummy_magic_0.Vb2 two_stage_opamp_dummy_magic_0.Vb2.n8 161.477
R7550 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n26 160.06
R7551 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n18 140.857
R7552 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 139.608
R7553 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n23 139.608
R7554 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 139.608
R7555 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 61.3349
R7556 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 49.8072
R7557 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n3 49.8072
R7558 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 49.8072
R7559 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n12 49.8072
R7560 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R7561 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R7562 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R7563 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.t0 24.0005
R7564 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R7565 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t1 24.0005
R7566 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R7567 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R7568 two_stage_opamp_dummy_magic_0.Vb2.n30 two_stage_opamp_dummy_magic_0.Vb2.n29 12.8443
R7569 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t10 11.2576
R7570 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t8 11.2576
R7571 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n20 7.563
R7572 two_stage_opamp_dummy_magic_0.Vb2 two_stage_opamp_dummy_magic_0.Vb2.n30 7.2505
R7573 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n25 4.54113
R7574 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 2.84425
R7575 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.n22 1.2505
R7576 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 0.928625
R7577 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t27 1172.87
R7578 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t33 1172.87
R7579 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t45 996.134
R7580 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t30 996.134
R7581 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t47 996.134
R7582 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t41 996.134
R7583 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t49 996.134
R7584 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t35 996.134
R7585 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t52 996.134
R7586 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t38 996.134
R7587 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t32 690.867
R7588 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t39 690.867
R7589 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t44 530.201
R7590 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t51 530.201
R7591 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t46 514.134
R7592 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t53 514.134
R7593 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t36 514.134
R7594 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t50 514.134
R7595 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t43 514.134
R7596 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t28 514.134
R7597 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t42 514.134
R7598 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t25 514.134
R7599 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t26 353.467
R7600 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t31 353.467
R7601 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t48 353.467
R7602 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t34 353.467
R7603 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t29 353.467
R7604 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t37 353.467
R7605 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t54 353.467
R7606 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t40 353.467
R7607 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 176.733
R7608 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.n48 176.733
R7609 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R7610 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R7611 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R7612 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R7613 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n28 176.733
R7614 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R7615 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R7616 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R7617 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R7618 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R7619 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 176.733
R7620 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R7621 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R7622 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R7623 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R7624 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R7625 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n51 166.258
R7626 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n11 163.626
R7627 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 163.001
R7628 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 163.001
R7629 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 163.001
R7630 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n12 163.001
R7631 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.541
R7632 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.541
R7633 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 158.501
R7634 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n0 117.888
R7635 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 117.326
R7636 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n7 117.326
R7637 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 117.326
R7638 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 117.326
R7639 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.n1 117.326
R7640 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 54.6272
R7641 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n24 54.6272
R7642 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 54.6272
R7643 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n33 54.6272
R7644 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 53.3126
R7645 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n46 53.3126
R7646 two_stage_opamp_dummy_magic_0.Y.t1 two_stage_opamp_dummy_magic_0.Y.n52 50.3031
R7647 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n21 16.8755
R7648 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R7649 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.t13 16.0005
R7650 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t3 16.0005
R7651 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t10 16.0005
R7652 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R7653 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R7654 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R7655 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t8 16.0005
R7656 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t2 16.0005
R7657 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t7 16.0005
R7658 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t12 16.0005
R7659 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R7660 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 13.4693
R7661 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t22 11.2576
R7662 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t24 11.2576
R7663 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t14 11.2576
R7664 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t21 11.2576
R7665 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t18 11.2576
R7666 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t17 11.2576
R7667 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t16 11.2576
R7668 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t20 11.2576
R7669 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t19 11.2576
R7670 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t23 11.2576
R7671 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t0 11.2576
R7672 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t15 11.2576
R7673 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n19 5.1255
R7674 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 4.5005
R7675 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n42 2.59425
R7676 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n10 1.8755
R7677 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n13 0.6255
R7678 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n15 0.6255
R7679 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n17 0.6255
R7680 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n2 0.563
R7681 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n4 0.563
R7682 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n6 0.563
R7683 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n8 0.563
R7684 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n14 146.47
R7685 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 146.47
R7686 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 145.906
R7687 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 145.906
R7688 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 145.906
R7689 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 145.906
R7690 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.n4 114.719
R7691 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.n1 114.719
R7692 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.n2 114.156
R7693 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.n5 114.156
R7694 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n0 109.656
R7695 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R7696 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R7697 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R7698 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R7699 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R7700 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R7701 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R7702 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R7703 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R7704 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R7705 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R7706 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R7707 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R7708 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R7709 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R7710 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R7711 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R7712 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R7713 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R7714 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R7715 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R7716 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R7717 two_stage_opamp_dummy_magic_0.VD2 two_stage_opamp_dummy_magic_0.VD2.n19 4.92758
R7718 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.n7 4.5005
R7719 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 0.563
R7720 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R7721 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.n6 0.563
R7722 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.n3 0.563
R7723 two_stage_opamp_dummy_magic_0.VD2 two_stage_opamp_dummy_magic_0.VD2.n8 0.313
R7724 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 0.234875
R7725 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n13 0.234875
R7726 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.n3 526.183
R7727 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 514.134
R7728 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n0 360.586
R7729 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 303.259
R7730 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 210.169
R7731 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t3 174.726
R7732 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t7 174.726
R7733 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 174.726
R7734 bgr_0.V_CUR_REF_REG.t0 bgr_0.V_CUR_REF_REG.n5 153.474
R7735 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 128.534
R7736 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t6 96.4005
R7737 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t2 39.4005
R7738 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t1 39.4005
R7739 bgr_0.V_p_2.n1 bgr_0.V_p_2.n2 229.562
R7740 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7741 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7742 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7743 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7744 bgr_0.V_p_2.n0 bgr_0.V_p_2.t10 98.7279
R7745 bgr_0.V_p_2.n5 bgr_0.V_p_2.t9 48.0005
R7746 bgr_0.V_p_2.n5 bgr_0.V_p_2.t0 48.0005
R7747 bgr_0.V_p_2.n4 bgr_0.V_p_2.t3 48.0005
R7748 bgr_0.V_p_2.n4 bgr_0.V_p_2.t5 48.0005
R7749 bgr_0.V_p_2.n3 bgr_0.V_p_2.t8 48.0005
R7750 bgr_0.V_p_2.n3 bgr_0.V_p_2.t1 48.0005
R7751 bgr_0.V_p_2.n2 bgr_0.V_p_2.t6 48.0005
R7752 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R7753 bgr_0.V_p_2.t4 bgr_0.V_p_2.n6 48.0005
R7754 bgr_0.V_p_2.n6 bgr_0.V_p_2.t7 48.0005
R7755 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7756 a_7460_23988.t0 a_7460_23988.t1 178.133
R7757 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 631.202
R7758 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 631.202
R7759 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 629.952
R7760 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 629.952
R7761 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 629.407
R7762 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 628.907
R7763 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 628.907
R7764 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 628.907
R7765 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 625.432
R7766 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 624.385
R7767 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R7768 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R7769 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R7770 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R7771 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R7772 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R7773 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R7774 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R7775 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R7776 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R7777 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R7778 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R7779 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R7780 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R7781 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R7782 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R7783 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R7784 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R7785 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R7786 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R7787 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 7.39633
R7788 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 6.188
R7789 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.n27 632.106
R7790 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n22 630.515
R7791 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n24 629.952
R7792 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n23 629.952
R7793 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 629.952
R7794 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n25 629.952
R7795 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t32 289.2
R7796 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t24 289.2
R7797 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R7798 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R7799 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R7800 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R7801 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R7802 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R7803 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R7804 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R7805 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R7806 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.n2 176.733
R7807 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.n3 176.733
R7808 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.n4 176.733
R7809 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R7810 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R7811 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R7812 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R7813 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n21 175.013
R7814 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n20 161.821
R7815 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R7816 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R7817 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R7818 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R7819 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R7820 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R7821 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R7822 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R7823 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t29 112.468
R7824 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R7825 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R7826 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R7827 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R7828 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R7829 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t17 112.468
R7830 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R7831 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R7832 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R7833 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R7834 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R7835 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R7836 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R7837 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t8 78.8005
R7838 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R7839 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R7840 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R7841 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R7842 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R7843 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R7844 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R7845 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 54.6272
R7846 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n9 54.6272
R7847 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t10 24.0005
R7848 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t11 24.0005
R7849 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 7.7505
R7850 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.n1 1.1255
R7851 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 1.1255
R7852 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.n1 630.984
R7853 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.n0 630.984
R7854 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 629.734
R7855 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 629.734
R7856 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.n2 629.734
R7857 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n10 629.47
R7858 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.n15 628.907
R7859 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.n13 628.907
R7860 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 628.907
R7861 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 625.234
R7862 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n9 624.385
R7863 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7864 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7865 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7866 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7867 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7868 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7869 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7870 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7871 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7872 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7873 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7874 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7875 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7876 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7877 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7878 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7879 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7880 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7881 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7882 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7883 two_stage_opamp_dummy_magic_0.V_err_p.t12 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7884 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7885 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 5.0005
R7886 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n8 4.5005
R7887 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 1.2505
R7888 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 1.2505
R7889 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.n7 1.2505
R7890 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 0.760917
R7891 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.n12 0.563
R7892 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.n14 0.563
R7893 a_6930_22564.t0 a_6930_22564.t1 178.133
R7894 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t13 369.534
R7895 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t12 369.534
R7896 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t29 369.534
R7897 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t17 369.534
R7898 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t21 369.534
R7899 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t20 369.534
R7900 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7901 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7902 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7903 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7904 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t14 238.322
R7905 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t27 238.322
R7906 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t26 192.8
R7907 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t19 192.8
R7908 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t16 192.8
R7909 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t23 192.8
R7910 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t22 192.8
R7911 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t24 192.8
R7912 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t10 192.8
R7913 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t18 192.8
R7914 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t25 192.8
R7915 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t11 192.8
R7916 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t15 192.8
R7917 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t28 192.8
R7918 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7919 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7920 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7921 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7922 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7923 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7924 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7925 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7926 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.n14 167.519
R7927 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7928 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t6 137.48
R7929 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t7 100.635
R7930 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7931 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7932 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7933 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7934 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7935 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7936 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t9 39.4005
R7937 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t1 39.4005
R7938 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t3 39.4005
R7939 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t5 39.4005
R7940 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t2 39.4005
R7941 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t4 39.4005
R7942 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t0 39.4005
R7943 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t8 39.4005
R7944 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 27.5005
R7945 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n13 9.53175
R7946 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7947 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 2.34425
R7948 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7949 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7950 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 1.688
R7951 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 610.534
R7952 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 610.534
R7953 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R7954 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R7955 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R7956 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R7957 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 433.8
R7958 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 433.8
R7959 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 433.8
R7960 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R7961 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R7962 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R7963 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R7964 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R7965 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R7966 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R7967 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R7968 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R7969 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R7970 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 433.8
R7971 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 339.836
R7972 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.834
R7973 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R7974 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 287.264
R7975 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 176.733
R7976 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R7977 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R7978 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R7979 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R7980 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R7981 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R7982 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R7983 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R7984 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R7985 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R7986 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R7987 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R7988 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R7989 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R7990 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 176.733
R7991 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 162.791
R7992 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 111.779
R7993 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 68.223
R7994 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.V_tail_gate.n29 58.7539
R7995 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 54.6272
R7996 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 54.6272
R7997 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 53.2453
R7998 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 52.01
R7999 two_stage_opamp_dummy_magic_0.V_tail_gate two_stage_opamp_dummy_magic_0.V_tail_gate.n6 51.6642
R8000 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R8001 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 39.4005
R8002 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R8003 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R8004 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R8005 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R8006 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R8007 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R8008 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R8009 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 16.0005
R8010 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R8011 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R8012 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R8013 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.t11 323.632
R8014 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t6 323.632
R8015 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.t12 168.701
R8016 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R8017 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t13 168.701
R8018 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t7 168.701
R8019 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.t8 168.701
R8020 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.t5 168.701
R8021 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R8022 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t4 168.701
R8023 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 165.8
R8024 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.n6 165.8
R8025 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 165.8
R8026 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.n1 165.8
R8027 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 116.546
R8028 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 116.546
R8029 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t2 107.328
R8030 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t1 107.328
R8031 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.n0 32.49
R8032 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 31.9025
R8033 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.n5 3.50675
R8034 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n2 1.28175
R8035 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n7 1.28175
R8036 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.n4 1.18175
R8037 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 1.18175
R8038 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.t30 217.776
R8039 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n10 114.469
R8040 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n3 114.469
R8041 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.n17 113.906
R8042 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n15 113.906
R8043 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n13 113.906
R8044 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n11 113.906
R8045 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.n8 113.906
R8046 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n6 113.906
R8047 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n4 113.906
R8048 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n20 109.406
R8049 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.n0 102.941
R8050 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.n37 102.285
R8051 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n35 102.284
R8052 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n33 102.284
R8053 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n31 102.284
R8054 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.n29 102.284
R8055 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n27 102.284
R8056 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.n25 102.284
R8057 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.n1 102.284
R8058 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n22 97.7845
R8059 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t6 16.0005
R8060 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t8 16.0005
R8061 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.t1 16.0005
R8062 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.t9 16.0005
R8063 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t5 16.0005
R8064 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t28 16.0005
R8065 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t32 16.0005
R8066 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t36 16.0005
R8067 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t7 16.0005
R8068 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t2 16.0005
R8069 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.t3 16.0005
R8070 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.t38 16.0005
R8071 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t37 16.0005
R8072 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t39 16.0005
R8073 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t4 16.0005
R8074 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t29 16.0005
R8075 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t33 16.0005
R8076 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t31 16.0005
R8077 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t40 16.0005
R8078 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t34 16.0005
R8079 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.t25 9.6005
R8080 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.t15 9.6005
R8081 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.t23 9.6005
R8082 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.t12 9.6005
R8083 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.t13 9.6005
R8084 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.t20 9.6005
R8085 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.t11 9.6005
R8086 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.t21 9.6005
R8087 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t14 9.6005
R8088 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t22 9.6005
R8089 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.t16 9.6005
R8090 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.t24 9.6005
R8091 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t19 9.6005
R8092 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t26 9.6005
R8093 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t18 9.6005
R8094 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t10 9.6005
R8095 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t35 9.6005
R8096 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t0 9.6005
R8097 two_stage_opamp_dummy_magic_0.V_source.t27 two_stage_opamp_dummy_magic_0.V_source.n38 9.6005
R8098 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.t17 9.6005
R8099 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n19 4.5005
R8100 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.n23 4.5005
R8101 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.n18 3.6255
R8102 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n21 1.80606
R8103 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n34 0.563
R8104 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.n36 0.563
R8105 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n12 0.563
R8106 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n14 0.563
R8107 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.n16 0.563
R8108 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n5 0.563
R8109 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.n7 0.563
R8110 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.n9 0.563
R8111 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.n2 0.563
R8112 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.n24 0.563
R8113 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n26 0.563
R8114 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.n28 0.563
R8115 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n30 0.563
R8116 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.n32 0.563
R8117 bgr_0.cap_res1.t0 bgr_0.cap_res1.t10 121.245
R8118 bgr_0.cap_res1.t16 bgr_0.cap_res1.t19 0.1603
R8119 bgr_0.cap_res1.t9 bgr_0.cap_res1.t15 0.1603
R8120 bgr_0.cap_res1.t14 bgr_0.cap_res1.t18 0.1603
R8121 bgr_0.cap_res1.t7 bgr_0.cap_res1.t13 0.1603
R8122 bgr_0.cap_res1.t1 bgr_0.cap_res1.t6 0.1603
R8123 bgr_0.cap_res1.n1 bgr_0.cap_res1.t17 0.159278
R8124 bgr_0.cap_res1.n2 bgr_0.cap_res1.t2 0.159278
R8125 bgr_0.cap_res1.n3 bgr_0.cap_res1.t8 0.159278
R8126 bgr_0.cap_res1.n4 bgr_0.cap_res1.t3 0.159278
R8127 bgr_0.cap_res1.n4 bgr_0.cap_res1.t16 0.1368
R8128 bgr_0.cap_res1.n4 bgr_0.cap_res1.t12 0.1368
R8129 bgr_0.cap_res1.n3 bgr_0.cap_res1.t9 0.1368
R8130 bgr_0.cap_res1.n3 bgr_0.cap_res1.t5 0.1368
R8131 bgr_0.cap_res1.n2 bgr_0.cap_res1.t14 0.1368
R8132 bgr_0.cap_res1.n2 bgr_0.cap_res1.t11 0.1368
R8133 bgr_0.cap_res1.n1 bgr_0.cap_res1.t7 0.1368
R8134 bgr_0.cap_res1.n1 bgr_0.cap_res1.t4 0.1368
R8135 bgr_0.cap_res1.n0 bgr_0.cap_res1.t1 0.1368
R8136 bgr_0.cap_res1.n0 bgr_0.cap_res1.t20 0.1368
R8137 bgr_0.cap_res1.t17 bgr_0.cap_res1.n0 0.00152174
R8138 bgr_0.cap_res1.t2 bgr_0.cap_res1.n1 0.00152174
R8139 bgr_0.cap_res1.t8 bgr_0.cap_res1.n2 0.00152174
R8140 bgr_0.cap_res1.t3 bgr_0.cap_res1.n3 0.00152174
R8141 bgr_0.cap_res1.t10 bgr_0.cap_res1.n4 0.00152174
R8142 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R8143 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R8144 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 325.473
R8145 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 310.488
R8146 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R8147 bgr_0.V_mir2.n4 bgr_0.V_mir2.t20 310.488
R8148 bgr_0.V_mir2.n2 bgr_0.V_mir2.t14 278.312
R8149 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 228.939
R8150 bgr_0.V_mir2.n3 bgr_0.V_mir2.n0 224.439
R8151 bgr_0.V_mir2.n18 bgr_0.V_mir2.t10 184.097
R8152 bgr_0.V_mir2.n11 bgr_0.V_mir2.t8 184.097
R8153 bgr_0.V_mir2.n6 bgr_0.V_mir2.t0 184.097
R8154 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R8155 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R8156 bgr_0.V_mir2.n5 bgr_0.V_mir2.n4 167.094
R8157 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R8158 bgr_0.V_mir2.n8 bgr_0.V_mir2.n6 152
R8159 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R8160 bgr_0.V_mir2.n16 bgr_0.V_mir2.t19 120.501
R8161 bgr_0.V_mir2.n17 bgr_0.V_mir2.t6 120.501
R8162 bgr_0.V_mir2.n9 bgr_0.V_mir2.t18 120.501
R8163 bgr_0.V_mir2.n10 bgr_0.V_mir2.t2 120.501
R8164 bgr_0.V_mir2.n4 bgr_0.V_mir2.t17 120.501
R8165 bgr_0.V_mir2.n5 bgr_0.V_mir2.t4 120.501
R8166 bgr_0.V_mir2.n1 bgr_0.V_mir2.t16 48.0005
R8167 bgr_0.V_mir2.n1 bgr_0.V_mir2.t12 48.0005
R8168 bgr_0.V_mir2.n0 bgr_0.V_mir2.t15 48.0005
R8169 bgr_0.V_mir2.n0 bgr_0.V_mir2.t13 48.0005
R8170 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R8171 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R8172 bgr_0.V_mir2.n6 bgr_0.V_mir2.n5 40.7027
R8173 bgr_0.V_mir2.n12 bgr_0.V_mir2.t3 39.4005
R8174 bgr_0.V_mir2.n12 bgr_0.V_mir2.t9 39.4005
R8175 bgr_0.V_mir2.n7 bgr_0.V_mir2.t5 39.4005
R8176 bgr_0.V_mir2.n7 bgr_0.V_mir2.t1 39.4005
R8177 bgr_0.V_mir2.n20 bgr_0.V_mir2.t7 39.4005
R8178 bgr_0.V_mir2.t11 bgr_0.V_mir2.n20 39.4005
R8179 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 15.8005
R8180 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 15.8005
R8181 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 9.3005
R8182 bgr_0.V_mir2.n3 bgr_0.V_mir2.n2 5.8755
R8183 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R8184 bgr_0.V_mir2.n15 bgr_0.V_mir2.n3 0.78175
R8185 bgr_0.Vin-.n7 bgr_0.Vin-.t12 688.859
R8186 bgr_0.Vin-.n9 bgr_0.Vin-.n8 514.134
R8187 bgr_0.Vin-.n6 bgr_0.Vin-.n5 351.522
R8188 bgr_0.Vin-.n11 bgr_0.Vin-.n10 213.4
R8189 bgr_0.Vin-.n7 bgr_0.Vin-.t8 174.726
R8190 bgr_0.Vin-.n8 bgr_0.Vin-.t10 174.726
R8191 bgr_0.Vin-.n9 bgr_0.Vin-.t9 174.726
R8192 bgr_0.Vin-.n10 bgr_0.Vin-.t11 174.726
R8193 bgr_0.Vin-.n4 bgr_0.Vin-.n2 173.029
R8194 bgr_0.Vin-.n4 bgr_0.Vin-.n3 168.654
R8195 bgr_0.Vin-.n8 bgr_0.Vin-.n7 128.534
R8196 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R8197 bgr_0.Vin-.n12 bgr_0.Vin-.t0 119.099
R8198 bgr_0.Vin-.n16 bgr_0.Vin-.n15 83.5719
R8199 bgr_0.Vin-.n1 bgr_0.Vin-.n0 83.5719
R8200 bgr_0.Vin-.n19 bgr_0.Vin-.n1 73.8495
R8201 bgr_0.Vin-.t3 bgr_0.Vin-.n14 65.0341
R8202 bgr_0.Vin-.n5 bgr_0.Vin-.t1 39.4005
R8203 bgr_0.Vin-.n5 bgr_0.Vin-.t2 39.4005
R8204 bgr_0.Vin-.n13 bgr_0.Vin-.n12 28.813
R8205 bgr_0.Vin-.n15 bgr_0.Vin-.n1 26.074
R8206 bgr_0.Vin-.n12 bgr_0.Vin-.n11 16.188
R8207 bgr_0.Vin-.n3 bgr_0.Vin-.t4 13.1338
R8208 bgr_0.Vin-.n3 bgr_0.Vin-.t6 13.1338
R8209 bgr_0.Vin-.n2 bgr_0.Vin-.t7 13.1338
R8210 bgr_0.Vin-.n2 bgr_0.Vin-.t5 13.1338
R8211 bgr_0.Vin-.n11 bgr_0.Vin-.n6 11.2193
R8212 bgr_0.Vin-.n6 bgr_0.Vin-.n4 3.8755
R8213 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56483
R8214 bgr_0.Vin-.n18 bgr_0.Vin-.n17 1.5505
R8215 bgr_0.Vin-.n17 bgr_0.Vin-.n0 0.885803
R8216 bgr_0.Vin-.n17 bgr_0.Vin-.n16 0.77514
R8217 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n0 0.756696
R8218 bgr_0.Vin-.n19 bgr_0.Vin-.n18 0.711459
R8219 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_0.Vin-.n19 0.576566
R8220 bgr_0.Vin-.n14 bgr_0.Vin-.n13 0.531499
R8221 bgr_0.Vin-.n15 bgr_0.Vin-.t3 0.290206
R8222 bgr_0.Vin-.n18 bgr_0.Vin-.n13 0.00817857
R8223 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 229.562
R8224 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R8225 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R8226 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R8227 bgr_0.V_p_1.n6 bgr_0.V_p_1.n0 228.938
R8228 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.7279
R8229 bgr_0.V_p_1.n5 bgr_0.V_p_1.t9 48.0005
R8230 bgr_0.V_p_1.n5 bgr_0.V_p_1.t1 48.0005
R8231 bgr_0.V_p_1.n4 bgr_0.V_p_1.t2 48.0005
R8232 bgr_0.V_p_1.n4 bgr_0.V_p_1.t5 48.0005
R8233 bgr_0.V_p_1.n3 bgr_0.V_p_1.t8 48.0005
R8234 bgr_0.V_p_1.n3 bgr_0.V_p_1.t0 48.0005
R8235 bgr_0.V_p_1.n2 bgr_0.V_p_1.t3 48.0005
R8236 bgr_0.V_p_1.n2 bgr_0.V_p_1.t6 48.0005
R8237 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8238 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R8239 bgr_0.V_p_1.n0 bgr_0.V_p_1.n1 1.8755
R8240 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 144.827
R8241 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 134.577
R8242 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 118.986
R8243 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 100.6
R8244 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 100.038
R8245 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 100.038
R8246 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 100.038
R8247 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 100.038
R8248 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 43.284
R8249 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 37.4067
R8250 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 24.0005
R8251 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 24.0005
R8252 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R8253 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 24.0005
R8254 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 8.0005
R8255 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R8256 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R8257 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 8.0005
R8258 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 8.0005
R8259 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 8.0005
R8260 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R8261 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R8262 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R8263 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R8264 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 5.6255
R8265 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 0.563
R8266 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 0.563
R8267 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 0.563
R8268 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 0.047375
R8269 VIN+.n9 VIN+.t2 490.072
R8270 VIN+.n4 VIN+.t9 449.868
R8271 VIN+.n0 VIN+.t10 449.868
R8272 VIN+.n4 VIN+.t3 273.134
R8273 VIN+.n5 VIN+.t8 273.134
R8274 VIN+.n6 VIN+.t1 273.134
R8275 VIN+.n7 VIN+.t6 273.134
R8276 VIN+.n3 VIN+.t4 273.134
R8277 VIN+.n2 VIN+.t7 273.134
R8278 VIN+.n1 VIN+.t0 273.134
R8279 VIN+.n0 VIN+.t5 273.134
R8280 VIN+.n7 VIN+.n6 176.733
R8281 VIN+.n6 VIN+.n5 176.733
R8282 VIN+.n5 VIN+.n4 176.733
R8283 VIN+.n1 VIN+.n0 176.733
R8284 VIN+.n2 VIN+.n1 176.733
R8285 VIN+.n3 VIN+.n2 176.733
R8286 VIN+.n9 VIN+.n8 165.8
R8287 VIN+.n8 VIN+.n7 56.2338
R8288 VIN+.n8 VIN+.n3 56.2338
R8289 VIN+ VIN+.n9 2.14112
R8290 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t12 685.053
R8291 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n2 633.639
R8292 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 630.234
R8293 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.n3 630.234
R8294 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.n0 226.534
R8295 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.n9 226.534
R8296 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 222.034
R8297 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t5 78.8005
R8298 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t6 78.8005
R8299 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t9 78.8005
R8300 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t7 78.8005
R8301 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.t11 78.8005
R8302 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.t8 78.8005
R8303 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t3 48.0005
R8304 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t10 48.0005
R8305 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t0 48.0005
R8306 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t2 48.0005
R8307 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.err_amp_out.n10 48.0005
R8308 two_stage_opamp_dummy_magic_0.err_amp_out.n10 two_stage_opamp_dummy_magic_0.err_amp_out.t1 48.0005
R8309 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 8.6255
R8310 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 5.7505
R8311 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n4 1.2505
R8312 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n1 1.2505
R8313 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R8314 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R8315 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 292.5
R8316 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 209.251
R8317 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 208.689
R8318 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 208.689
R8319 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 208.689
R8320 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 208.689
R8321 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 120.305
R8322 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 52.763
R8323 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 51.7297
R8324 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 50.813
R8325 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R8326 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 39.4005
R8327 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 39.4005
R8328 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 39.4005
R8329 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 39.4005
R8330 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R8331 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R8332 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 19.7005
R8333 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 19.7005
R8334 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R8335 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R8336 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R8337 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 19.7005
R8338 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R8339 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 19.7005
R8340 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R8341 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 5.90675
R8342 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R8343 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R8344 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R8345 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t35 652.076
R8346 two_stage_opamp_dummy_magic_0.VD4.n61 two_stage_opamp_dummy_magic_0.VD4.t32 652.076
R8347 two_stage_opamp_dummy_magic_0.VD4.n60 two_stage_opamp_dummy_magic_0.VD4.n13 585
R8348 two_stage_opamp_dummy_magic_0.VD4.n42 two_stage_opamp_dummy_magic_0.VD4.n41 585
R8349 two_stage_opamp_dummy_magic_0.VD4.n48 two_stage_opamp_dummy_magic_0.VD4.n13 290.233
R8350 two_stage_opamp_dummy_magic_0.VD4.n54 two_stage_opamp_dummy_magic_0.VD4.n13 290.233
R8351 two_stage_opamp_dummy_magic_0.VD4.n49 two_stage_opamp_dummy_magic_0.VD4.n13 290.233
R8352 two_stage_opamp_dummy_magic_0.VD4.n41 two_stage_opamp_dummy_magic_0.VD4.n30 290.233
R8353 two_stage_opamp_dummy_magic_0.VD4.n41 two_stage_opamp_dummy_magic_0.VD4.n35 290.233
R8354 two_stage_opamp_dummy_magic_0.VD4.n41 two_stage_opamp_dummy_magic_0.VD4.n40 290.233
R8355 two_stage_opamp_dummy_magic_0.VD4.n49 two_stage_opamp_dummy_magic_0.VD4.n46 242.903
R8356 two_stage_opamp_dummy_magic_0.VD4.n40 two_stage_opamp_dummy_magic_0.VD4.n18 242.903
R8357 two_stage_opamp_dummy_magic_0.VD4.n60 two_stage_opamp_dummy_magic_0.VD4.n59 238.367
R8358 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n14 185
R8359 two_stage_opamp_dummy_magic_0.VD4.n57 two_stage_opamp_dummy_magic_0.VD4.n56 185
R8360 two_stage_opamp_dummy_magic_0.VD4.n58 two_stage_opamp_dummy_magic_0.VD4.n57 185
R8361 two_stage_opamp_dummy_magic_0.VD4.n55 two_stage_opamp_dummy_magic_0.VD4.n47 185
R8362 two_stage_opamp_dummy_magic_0.VD4.n53 two_stage_opamp_dummy_magic_0.VD4.n52 185
R8363 two_stage_opamp_dummy_magic_0.VD4.n51 two_stage_opamp_dummy_magic_0.VD4.n50 185
R8364 two_stage_opamp_dummy_magic_0.VD4.n43 two_stage_opamp_dummy_magic_0.VD4.n42 185
R8365 two_stage_opamp_dummy_magic_0.VD4.n44 two_stage_opamp_dummy_magic_0.VD4.n43 185
R8366 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n19 185
R8367 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n31 185
R8368 two_stage_opamp_dummy_magic_0.VD4.n34 two_stage_opamp_dummy_magic_0.VD4.n33 185
R8369 two_stage_opamp_dummy_magic_0.VD4.n37 two_stage_opamp_dummy_magic_0.VD4.n36 185
R8370 two_stage_opamp_dummy_magic_0.VD4.n39 two_stage_opamp_dummy_magic_0.VD4.n38 185
R8371 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.VD4.n44 170.513
R8372 two_stage_opamp_dummy_magic_0.VD4.n58 two_stage_opamp_dummy_magic_0.VD4.t33 170.513
R8373 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n0 163.626
R8374 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n9 163.001
R8375 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 163.001
R8376 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 163.001
R8377 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.n3 163.001
R8378 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n1 163.001
R8379 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n11 159.804
R8380 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n20 159.803
R8381 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.n22 159.803
R8382 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 159.803
R8383 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.803
R8384 two_stage_opamp_dummy_magic_0.VD4.n57 two_stage_opamp_dummy_magic_0.VD4.n15 150
R8385 two_stage_opamp_dummy_magic_0.VD4.n57 two_stage_opamp_dummy_magic_0.VD4.n47 150
R8386 two_stage_opamp_dummy_magic_0.VD4.n52 two_stage_opamp_dummy_magic_0.VD4.n51 150
R8387 two_stage_opamp_dummy_magic_0.VD4.n43 two_stage_opamp_dummy_magic_0.VD4.n19 150
R8388 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 150
R8389 two_stage_opamp_dummy_magic_0.VD4.n38 two_stage_opamp_dummy_magic_0.VD4.n37 150
R8390 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.VD4.t36 146.155
R8391 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t22 146.155
R8392 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.VD4.t18 146.155
R8393 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.VD4.t24 146.155
R8394 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t28 146.155
R8395 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.VD4.t12 146.155
R8396 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.VD4.t14 146.155
R8397 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t16 146.155
R8398 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.VD4.t20 146.155
R8399 two_stage_opamp_dummy_magic_0.VD4.t30 two_stage_opamp_dummy_magic_0.VD4.t26 146.155
R8400 two_stage_opamp_dummy_magic_0.VD4.t33 two_stage_opamp_dummy_magic_0.VD4.t30 146.155
R8401 two_stage_opamp_dummy_magic_0.VD4.n59 two_stage_opamp_dummy_magic_0.VD4.n58 65.8183
R8402 two_stage_opamp_dummy_magic_0.VD4.n58 two_stage_opamp_dummy_magic_0.VD4.n45 65.8183
R8403 two_stage_opamp_dummy_magic_0.VD4.n58 two_stage_opamp_dummy_magic_0.VD4.n46 65.8183
R8404 two_stage_opamp_dummy_magic_0.VD4.n44 two_stage_opamp_dummy_magic_0.VD4.n16 65.8183
R8405 two_stage_opamp_dummy_magic_0.VD4.n44 two_stage_opamp_dummy_magic_0.VD4.n17 65.8183
R8406 two_stage_opamp_dummy_magic_0.VD4.n44 two_stage_opamp_dummy_magic_0.VD4.n18 65.8183
R8407 two_stage_opamp_dummy_magic_0.VD4.n47 two_stage_opamp_dummy_magic_0.VD4.n45 53.3664
R8408 two_stage_opamp_dummy_magic_0.VD4.n51 two_stage_opamp_dummy_magic_0.VD4.n46 53.3664
R8409 two_stage_opamp_dummy_magic_0.VD4.n59 two_stage_opamp_dummy_magic_0.VD4.n15 53.3664
R8410 two_stage_opamp_dummy_magic_0.VD4.n52 two_stage_opamp_dummy_magic_0.VD4.n45 53.3664
R8411 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n16 53.3664
R8412 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n17 53.3664
R8413 two_stage_opamp_dummy_magic_0.VD4.n38 two_stage_opamp_dummy_magic_0.VD4.n18 53.3664
R8414 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.n16 53.3664
R8415 two_stage_opamp_dummy_magic_0.VD4.n37 two_stage_opamp_dummy_magic_0.VD4.n17 53.3664
R8416 two_stage_opamp_dummy_magic_0.VD4.n61 two_stage_opamp_dummy_magic_0.VD4.n60 22.8576
R8417 two_stage_opamp_dummy_magic_0.VD4.n42 two_stage_opamp_dummy_magic_0.VD4.n28 22.8576
R8418 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.n27 14.4255
R8419 two_stage_opamp_dummy_magic_0.VD4.n62 two_stage_opamp_dummy_magic_0.VD4.n61 13.8005
R8420 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R8421 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R8422 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R8423 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R8424 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R8425 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R8426 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R8427 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t19 11.2576
R8428 two_stage_opamp_dummy_magic_0.VD4.n41 two_stage_opamp_dummy_magic_0.VD4.t37 11.2576
R8429 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t34 11.2576
R8430 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R8431 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t4 11.2576
R8432 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t2 11.2576
R8433 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t5 11.2576
R8434 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8435 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R8436 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R8437 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R8438 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t3 11.2576
R8439 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R8440 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R8441 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R8442 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R8443 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R8444 two_stage_opamp_dummy_magic_0.VD4.n60 two_stage_opamp_dummy_magic_0.VD4.n14 9.14336
R8445 two_stage_opamp_dummy_magic_0.VD4.n56 two_stage_opamp_dummy_magic_0.VD4.n55 9.14336
R8446 two_stage_opamp_dummy_magic_0.VD4.n53 two_stage_opamp_dummy_magic_0.VD4.n50 9.14336
R8447 two_stage_opamp_dummy_magic_0.VD4.n42 two_stage_opamp_dummy_magic_0.VD4.n29 9.14336
R8448 two_stage_opamp_dummy_magic_0.VD4.n34 two_stage_opamp_dummy_magic_0.VD4.n31 9.14336
R8449 two_stage_opamp_dummy_magic_0.VD4.n39 two_stage_opamp_dummy_magic_0.VD4.n36 9.14336
R8450 two_stage_opamp_dummy_magic_0.VD4.n63 two_stage_opamp_dummy_magic_0.VD4.n10 8.2505
R8451 two_stage_opamp_dummy_magic_0.VD4.n63 two_stage_opamp_dummy_magic_0.VD4.n62 5.3755
R8452 two_stage_opamp_dummy_magic_0.VD4.n48 two_stage_opamp_dummy_magic_0.VD4.n14 4.53698
R8453 two_stage_opamp_dummy_magic_0.VD4.n55 two_stage_opamp_dummy_magic_0.VD4.n54 4.53698
R8454 two_stage_opamp_dummy_magic_0.VD4.n50 two_stage_opamp_dummy_magic_0.VD4.n49 4.53698
R8455 two_stage_opamp_dummy_magic_0.VD4.n56 two_stage_opamp_dummy_magic_0.VD4.n48 4.53698
R8456 two_stage_opamp_dummy_magic_0.VD4.n54 two_stage_opamp_dummy_magic_0.VD4.n53 4.53698
R8457 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.n29 4.53698
R8458 two_stage_opamp_dummy_magic_0.VD4.n35 two_stage_opamp_dummy_magic_0.VD4.n34 4.53698
R8459 two_stage_opamp_dummy_magic_0.VD4.n40 two_stage_opamp_dummy_magic_0.VD4.n39 4.53698
R8460 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 4.53698
R8461 two_stage_opamp_dummy_magic_0.VD4.n36 two_stage_opamp_dummy_magic_0.VD4.n35 4.53698
R8462 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.n2 0.6255
R8463 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n4 0.6255
R8464 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n6 0.6255
R8465 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n8 0.6255
R8466 two_stage_opamp_dummy_magic_0.VD4.n62 two_stage_opamp_dummy_magic_0.VD4.n12 0.6255
R8467 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.6255
R8468 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n23 0.6255
R8469 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.n21 0.6255
R8470 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.n12 0.6255
R8471 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n63 0.063
R8472 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8473 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8474 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8475 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8476 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8477 bgr_0.START_UP.n0 bgr_0.START_UP.t1 130.001
R8478 bgr_0.START_UP.n0 bgr_0.START_UP.t0 81.7074
R8479 bgr_0.START_UP bgr_0.START_UP.n0 36.9489
R8480 bgr_0.START_UP bgr_0.START_UP.n5 13.4693
R8481 bgr_0.START_UP.n1 bgr_0.START_UP.t2 13.1338
R8482 bgr_0.START_UP.n1 bgr_0.START_UP.t4 13.1338
R8483 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8484 bgr_0.START_UP.n2 bgr_0.START_UP.t5 13.1338
R8485 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8486 a_5980_2720.t0 a_5980_2720.t1 169.905
R8487 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 652.076
R8488 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 652.076
R8489 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n27 585
R8490 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 585
R8491 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 290.233
R8492 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n21 290.233
R8493 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n26 290.233
R8494 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n43 290.233
R8495 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 290.233
R8496 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n44 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 290.233
R8497 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 242.903
R8498 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 242.903
R8499 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n41 238.367
R8500 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n28 185
R8501 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n29 185
R8502 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 185
R8503 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 185
R8504 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n19 185
R8505 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n22 185
R8506 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n24 185
R8507 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 185
R8508 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 185
R8509 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n39 185
R8510 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n37 185
R8511 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n32 185
R8512 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n34 185
R8513 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n30 170.513
R8514 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 170.513
R8515 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 169.694
R8516 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 155.303
R8517 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 150
R8518 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n39 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n38 150
R8519 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n35 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n32 150
R8520 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n29 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 150
R8521 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 150
R8522 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n23 150
R8523 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 146.155
R8524 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 146.155
R8525 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 65.8183
R8526 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 65.8183
R8527 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n30 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 65.8183
R8528 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n40 65.8183
R8529 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n31 65.8183
R8530 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n40 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n36 65.8183
R8531 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n38 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n31 53.3664
R8532 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n36 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n35 53.3664
R8533 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 53.3664
R8534 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 53.3664
R8535 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n24 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 53.3664
R8536 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 53.3664
R8537 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n23 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 53.3664
R8538 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n41 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 53.3664
R8539 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n32 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n31 53.3664
R8540 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 22.8576
R8541 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n42 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 22.8576
R8542 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 14.4255
R8543 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 14.0505
R8544 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 11.2576
R8545 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 11.2576
R8546 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 11.2576
R8547 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 11.2576
R8548 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n27 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 11.2576
R8549 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n44 11.2576
R8550 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n28 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 9.14336
R8551 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 9.14336
R8552 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n25 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n22 9.14336
R8553 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 9.14336
R8554 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 9.14336
R8555 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n33 9.14336
R8556 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 4.53698
R8557 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n21 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n20 4.53698
R8558 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n26 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n25 4.53698
R8559 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.53698
R8560 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n22 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n21 4.53698
R8561 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n42 4.53698
R8562 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n37 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 4.53698
R8563 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n34 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 4.53698
R8564 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n43 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 4.53698
R8565 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n33 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 4.53698
R8566 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 4.5005
R8567 a_14010_2720.t0 a_14010_2720.t1 169.905
R8568 VIN-.n9 VIN-.t5 490.075
R8569 VIN-.n4 VIN-.t7 449.868
R8570 VIN-.n0 VIN-.t10 449.868
R8571 VIN-.n4 VIN-.t1 273.134
R8572 VIN-.n5 VIN-.t6 273.134
R8573 VIN-.n6 VIN-.t0 273.134
R8574 VIN-.n7 VIN-.t9 273.134
R8575 VIN-.n3 VIN-.t3 273.134
R8576 VIN-.n2 VIN-.t8 273.134
R8577 VIN-.n1 VIN-.t2 273.134
R8578 VIN-.n0 VIN-.t4 273.134
R8579 VIN-.n7 VIN-.n6 176.733
R8580 VIN-.n6 VIN-.n5 176.733
R8581 VIN-.n5 VIN-.n4 176.733
R8582 VIN-.n1 VIN-.n0 176.733
R8583 VIN-.n2 VIN-.n1 176.733
R8584 VIN-.n3 VIN-.n2 176.733
R8585 VIN-.n9 VIN-.n8 165.8
R8586 VIN-.n8 VIN-.n7 56.2338
R8587 VIN-.n8 VIN-.n3 56.2338
R8588 VIN- VIN-.n9 2.14112
R8589 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R8590 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R8591 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R8592 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 209.251
R8593 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 208.689
R8594 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 208.689
R8595 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 208.689
R8596 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 208.689
R8597 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 120.305
R8598 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R8599 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 52.1563
R8600 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 50.813
R8601 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R8602 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R8603 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R8604 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 39.4005
R8605 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R8606 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 39.4005
R8607 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R8608 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 19.7005
R8609 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R8610 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R8611 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R8612 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R8613 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R8614 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 19.7005
R8615 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R8616 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R8617 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 5.90675
R8618 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R8619 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R8620 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R8621 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R8622 a_12530_23988.t0 a_12530_23988.t1 178.133
R8623 a_7580_22380.t0 a_7580_22380.t1 178.133
R8624 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 223.377
R8625 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R8626 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t1 16.0005
R8627 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t3 9.6005
R8628 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R8629 a_5700_5524.t0 a_5700_5524.t1 169.905
R8630 a_6810_23838.t0 a_6810_23838.t1 178.133
R8631 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 195.608
R8632 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 84.0884
R8633 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 83.5719
R8634 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 83.5719
R8635 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 83.5719
R8636 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 83.5719
R8637 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 83.5719
R8638 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 83.5719
R8639 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 83.5719
R8640 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 83.5719
R8641 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 83.5719
R8642 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 83.5719
R8643 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 83.5719
R8644 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 83.5719
R8645 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 83.5719
R8646 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 83.5719
R8647 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 83.5719
R8648 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 83.5719
R8649 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 83.5719
R8650 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R8651 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 83.5719
R8652 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 83.5719
R8653 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R8654 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 83.5719
R8655 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 83.5719
R8656 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 73.8495
R8657 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 73.3165
R8658 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 73.3165
R8659 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 73.3165
R8660 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 73.3165
R8661 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R8662 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 73.3165
R8663 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 73.19
R8664 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 73.19
R8665 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 73.19
R8666 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 73.19
R8667 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R8668 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 73.19
R8669 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 65.0299
R8670 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 65.0299
R8671 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 26.074
R8672 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 26.074
R8673 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 26.074
R8674 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 26.074
R8675 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 26.074
R8676 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 26.074
R8677 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 26.074
R8678 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 26.074
R8679 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 26.074
R8680 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n142 26.074
R8681 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 25.7843
R8682 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 25.7843
R8683 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 25.7843
R8684 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 25.7843
R8685 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 25.7843
R8686 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 25.7843
R8687 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n144 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n143 19.9902
R8688 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 9.3005
R8689 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 9.3005
R8690 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 9.3005
R8691 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R8692 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 9.3005
R8693 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 9.3005
R8694 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R8695 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R8696 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 9.3005
R8697 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R8698 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 9.3005
R8699 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R8700 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R8701 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R8702 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R8703 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 9.3005
R8704 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R8705 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R8706 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 9.3005
R8707 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 9.3005
R8708 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R8709 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 9.3005
R8710 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 9.3005
R8711 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 9.3005
R8712 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 9.3005
R8713 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 9.3005
R8714 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 9.3005
R8715 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R8716 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R8717 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 9.3005
R8718 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 9.3005
R8719 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R8720 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R8721 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 9.3005
R8722 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 9.3005
R8723 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R8724 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R8725 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 9.3005
R8726 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R8727 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 9.3005
R8728 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 9.3005
R8729 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R8730 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 9.3005
R8731 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R8732 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 9.3005
R8733 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R8734 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 9.3005
R8735 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R8736 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 9.3005
R8737 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 9.3005
R8738 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 9.3005
R8739 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 9.3005
R8740 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 9.3005
R8741 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 9.3005
R8742 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 4.64654
R8743 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 4.64654
R8744 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 4.64654
R8745 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 4.64654
R8746 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 4.64654
R8747 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 4.64654
R8748 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 4.64654
R8749 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 4.64654
R8750 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 4.64654
R8751 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 2.36206
R8752 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 2.36206
R8753 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 2.36206
R8754 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 2.36206
R8755 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 2.19742
R8756 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 2.19742
R8757 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 2.19742
R8758 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 2.19742
R8759 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n146 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 1.56836
R8760 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 1.56363
R8761 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 1.56363
R8762 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 1.5505
R8763 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 1.5505
R8764 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 1.5505
R8765 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.5505
R8766 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 1.5505
R8767 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 1.5505
R8768 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 1.5505
R8769 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R8770 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 1.5505
R8771 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.5505
R8772 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 1.5505
R8773 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.5505
R8774 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 1.5505
R8775 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 1.5505
R8776 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 1.5505
R8777 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n147 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n146 1.5505
R8778 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R8779 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.5505
R8780 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 1.5505
R8781 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 1.25468
R8782 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.25468
R8783 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 1.25468
R8784 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 1.25468
R8785 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 1.25468
R8786 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.25468
R8787 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 1.19225
R8788 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 1.19225
R8789 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.19225
R8790 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 1.19225
R8791 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.19225
R8792 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.19225
R8793 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n145 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.14402
R8794 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R8795 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.07024
R8796 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 1.07024
R8797 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 1.07024
R8798 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 1.07024
R8799 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 1.07024
R8800 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 1.0237
R8801 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.0237
R8802 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.0237
R8803 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 1.0237
R8804 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 1.0237
R8805 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 1.0237
R8806 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 0.885803
R8807 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 0.885803
R8808 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.885803
R8809 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 0.885803
R8810 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.885803
R8811 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 0.885803
R8812 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.885803
R8813 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R8814 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.812055
R8815 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 0.812055
R8816 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.77514
R8817 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.77514
R8818 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.77514
R8819 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.77514
R8820 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R8821 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.77514
R8822 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.77514
R8823 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.77514
R8824 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8825 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8826 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8827 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R8828 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 0.756696
R8829 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.756696
R8830 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.756696
R8831 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R8832 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.711459
R8833 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n147 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 0.701365
R8834 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 0.647417
R8835 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.647417
R8836 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 0.590702
R8837 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.590702
R8838 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.590702
R8839 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.590702
R8840 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.590702
R8841 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.590702
R8842 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.576566
R8843 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 0.530034
R8844 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.530034
R8845 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R8846 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R8847 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R8848 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 0.290206
R8849 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 0.290206
R8850 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.290206
R8851 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 0.290206
R8852 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 0.290206
R8853 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8854 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8855 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.203382
R8856 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8857 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8858 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R8859 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n147 0.203382
R8860 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 0.154071
R8861 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 0.154071
R8862 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 0.154071
R8863 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.154071
R8864 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.137464
R8865 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.137464
R8866 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 0.134964
R8867 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.134964
R8868 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.0183571
R8869 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.0183571
R8870 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.0183571
R8871 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.0183571
R8872 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.0183571
R8873 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.0183571
R8874 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.0183571
R8875 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.0183571
R8876 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.0183571
R8877 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.0183571
R8878 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.0183571
R8879 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.0183571
R8880 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.0183571
R8881 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.0183571
R8882 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.0183571
R8883 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.0183571
R8884 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.0183571
R8885 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 0.0183571
R8886 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n146 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R8887 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.0106786
R8888 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 0.0106786
R8889 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.0106786
R8890 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8891 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.00992001
R8892 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.00992001
R8893 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.00992001
R8894 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.00992001
R8895 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.00992001
R8896 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.00992001
R8897 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 0.00992001
R8898 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R8899 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.00992001
R8900 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.00992001
R8901 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.00992001
R8902 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.00992001
R8903 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.00992001
R8904 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 0.00992001
R8905 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.00992001
R8906 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 0.00992001
R8907 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.00992001
R8908 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 0.00817857
R8909 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.00817857
R8910 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 0.00817857
R8911 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.00817857
R8912 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R8913 a_5580_5524.t0 a_5580_5524.t1 262.248
R8914 a_12410_22380.t0 a_12410_22380.t1 178.133
R8915 a_13060_22630.t0 a_13060_22630.t1 178.133
R8916 two_stage_opamp_dummy_magic_0.Vb2_2.n32 two_stage_opamp_dummy_magic_0.Vb2_2.n31 692.967
R8917 two_stage_opamp_dummy_magic_0.Vb2_2.n34 two_stage_opamp_dummy_magic_0.Vb2_2.t1 652.076
R8918 two_stage_opamp_dummy_magic_0.Vb2_2.n30 two_stage_opamp_dummy_magic_0.Vb2_2.t4 652.076
R8919 two_stage_opamp_dummy_magic_0.Vb2_2.n36 two_stage_opamp_dummy_magic_0.Vb2_2.n0 587.407
R8920 two_stage_opamp_dummy_magic_0.Vb2_2.n41 two_stage_opamp_dummy_magic_0.Vb2_2.n2 587.407
R8921 two_stage_opamp_dummy_magic_0.Vb2_2.n29 two_stage_opamp_dummy_magic_0.Vb2_2.n11 585
R8922 two_stage_opamp_dummy_magic_0.Vb2_2.n3 two_stage_opamp_dummy_magic_0.Vb2_2.n0 585
R8923 two_stage_opamp_dummy_magic_0.Vb2_2.t3 two_stage_opamp_dummy_magic_0.Vb2_2.n44 585
R8924 two_stage_opamp_dummy_magic_0.Vb2_2.n43 two_stage_opamp_dummy_magic_0.Vb2_2.n2 585
R8925 two_stage_opamp_dummy_magic_0.Vb2_2.n17 two_stage_opamp_dummy_magic_0.Vb2_2.n11 290.233
R8926 two_stage_opamp_dummy_magic_0.Vb2_2.n23 two_stage_opamp_dummy_magic_0.Vb2_2.n11 290.233
R8927 two_stage_opamp_dummy_magic_0.Vb2_2.n18 two_stage_opamp_dummy_magic_0.Vb2_2.n11 290.233
R8928 two_stage_opamp_dummy_magic_0.Vb2_2.t3 two_stage_opamp_dummy_magic_0.Vb2_2.n0 246.25
R8929 two_stage_opamp_dummy_magic_0.Vb2_2.t3 two_stage_opamp_dummy_magic_0.Vb2_2.n2 246.25
R8930 two_stage_opamp_dummy_magic_0.Vb2_2.n41 two_stage_opamp_dummy_magic_0.Vb2_2.n40 243.698
R8931 two_stage_opamp_dummy_magic_0.Vb2_2.n18 two_stage_opamp_dummy_magic_0.Vb2_2.n15 242.903
R8932 two_stage_opamp_dummy_magic_0.Vb2_2.n29 two_stage_opamp_dummy_magic_0.Vb2_2.n28 238.367
R8933 two_stage_opamp_dummy_magic_0.Vb2_2.n13 two_stage_opamp_dummy_magic_0.Vb2_2.n12 185
R8934 two_stage_opamp_dummy_magic_0.Vb2_2.n26 two_stage_opamp_dummy_magic_0.Vb2_2.n25 185
R8935 two_stage_opamp_dummy_magic_0.Vb2_2.n27 two_stage_opamp_dummy_magic_0.Vb2_2.n26 185
R8936 two_stage_opamp_dummy_magic_0.Vb2_2.n24 two_stage_opamp_dummy_magic_0.Vb2_2.n16 185
R8937 two_stage_opamp_dummy_magic_0.Vb2_2.n22 two_stage_opamp_dummy_magic_0.Vb2_2.n21 185
R8938 two_stage_opamp_dummy_magic_0.Vb2_2.n20 two_stage_opamp_dummy_magic_0.Vb2_2.n19 185
R8939 two_stage_opamp_dummy_magic_0.Vb2_2.n38 two_stage_opamp_dummy_magic_0.Vb2_2.n37 185
R8940 two_stage_opamp_dummy_magic_0.Vb2_2.n39 two_stage_opamp_dummy_magic_0.Vb2_2.n38 185
R8941 two_stage_opamp_dummy_magic_0.Vb2_2.n35 two_stage_opamp_dummy_magic_0.Vb2_2.n10 185
R8942 two_stage_opamp_dummy_magic_0.Vb2_2.n7 two_stage_opamp_dummy_magic_0.Vb2_2.n3 185
R8943 two_stage_opamp_dummy_magic_0.Vb2_2.n44 two_stage_opamp_dummy_magic_0.Vb2_2.n4 185
R8944 two_stage_opamp_dummy_magic_0.Vb2_2.n43 two_stage_opamp_dummy_magic_0.Vb2_2.n5 185
R8945 two_stage_opamp_dummy_magic_0.Vb2_2.n42 two_stage_opamp_dummy_magic_0.Vb2_2.n6 185
R8946 two_stage_opamp_dummy_magic_0.Vb2_2.n39 two_stage_opamp_dummy_magic_0.Vb2_2.t2 170.513
R8947 two_stage_opamp_dummy_magic_0.Vb2_2.n27 two_stage_opamp_dummy_magic_0.Vb2_2.t5 170.513
R8948 two_stage_opamp_dummy_magic_0.Vb2_2.n32 two_stage_opamp_dummy_magic_0.Vb2_2.n1 155.304
R8949 two_stage_opamp_dummy_magic_0.Vb2_2.n26 two_stage_opamp_dummy_magic_0.Vb2_2.n13 150
R8950 two_stage_opamp_dummy_magic_0.Vb2_2.n26 two_stage_opamp_dummy_magic_0.Vb2_2.n16 150
R8951 two_stage_opamp_dummy_magic_0.Vb2_2.n21 two_stage_opamp_dummy_magic_0.Vb2_2.n20 150
R8952 two_stage_opamp_dummy_magic_0.Vb2_2.n38 two_stage_opamp_dummy_magic_0.Vb2_2.n10 150
R8953 two_stage_opamp_dummy_magic_0.Vb2_2.n7 two_stage_opamp_dummy_magic_0.Vb2_2.n4 150
R8954 two_stage_opamp_dummy_magic_0.Vb2_2.n6 two_stage_opamp_dummy_magic_0.Vb2_2.n5 150
R8955 two_stage_opamp_dummy_magic_0.Vb2_2.t7 two_stage_opamp_dummy_magic_0.Vb2_2.t2 146.155
R8956 two_stage_opamp_dummy_magic_0.Vb2_2.t5 two_stage_opamp_dummy_magic_0.Vb2_2.t7 146.155
R8957 two_stage_opamp_dummy_magic_0.Vb2_2.n28 two_stage_opamp_dummy_magic_0.Vb2_2.n27 65.8183
R8958 two_stage_opamp_dummy_magic_0.Vb2_2.n27 two_stage_opamp_dummy_magic_0.Vb2_2.n14 65.8183
R8959 two_stage_opamp_dummy_magic_0.Vb2_2.n27 two_stage_opamp_dummy_magic_0.Vb2_2.n15 65.8183
R8960 two_stage_opamp_dummy_magic_0.Vb2_2.n39 two_stage_opamp_dummy_magic_0.Vb2_2.n8 65.8183
R8961 two_stage_opamp_dummy_magic_0.Vb2_2.n39 two_stage_opamp_dummy_magic_0.Vb2_2.n9 65.8183
R8962 two_stage_opamp_dummy_magic_0.Vb2_2.n40 two_stage_opamp_dummy_magic_0.Vb2_2.n39 65.8183
R8963 two_stage_opamp_dummy_magic_0.Vb2_2.n16 two_stage_opamp_dummy_magic_0.Vb2_2.n14 53.3664
R8964 two_stage_opamp_dummy_magic_0.Vb2_2.n20 two_stage_opamp_dummy_magic_0.Vb2_2.n15 53.3664
R8965 two_stage_opamp_dummy_magic_0.Vb2_2.n28 two_stage_opamp_dummy_magic_0.Vb2_2.n13 53.3664
R8966 two_stage_opamp_dummy_magic_0.Vb2_2.n21 two_stage_opamp_dummy_magic_0.Vb2_2.n14 53.3664
R8967 two_stage_opamp_dummy_magic_0.Vb2_2.n10 two_stage_opamp_dummy_magic_0.Vb2_2.n8 53.3664
R8968 two_stage_opamp_dummy_magic_0.Vb2_2.n9 two_stage_opamp_dummy_magic_0.Vb2_2.n4 53.3664
R8969 two_stage_opamp_dummy_magic_0.Vb2_2.n40 two_stage_opamp_dummy_magic_0.Vb2_2.n6 53.3664
R8970 two_stage_opamp_dummy_magic_0.Vb2_2.n8 two_stage_opamp_dummy_magic_0.Vb2_2.n7 53.3664
R8971 two_stage_opamp_dummy_magic_0.Vb2_2.n9 two_stage_opamp_dummy_magic_0.Vb2_2.n5 53.3664
R8972 two_stage_opamp_dummy_magic_0.Vb2_2.n30 two_stage_opamp_dummy_magic_0.Vb2_2.n29 22.8576
R8973 two_stage_opamp_dummy_magic_0.Vb2_2.n37 two_stage_opamp_dummy_magic_0.Vb2_2.n34 22.8576
R8974 two_stage_opamp_dummy_magic_0.Vb2_2.n31 two_stage_opamp_dummy_magic_0.Vb2_2.t0 21.8894
R8975 two_stage_opamp_dummy_magic_0.Vb2_2.n31 two_stage_opamp_dummy_magic_0.Vb2_2.t9 21.8894
R8976 two_stage_opamp_dummy_magic_0.Vb2_2.n33 two_stage_opamp_dummy_magic_0.Vb2_2.n30 14.4255
R8977 two_stage_opamp_dummy_magic_0.Vb2_2.n34 two_stage_opamp_dummy_magic_0.Vb2_2.n33 14.0505
R8978 two_stage_opamp_dummy_magic_0.Vb2_2.n11 two_stage_opamp_dummy_magic_0.Vb2_2.t6 11.2576
R8979 two_stage_opamp_dummy_magic_0.Vb2_2.t3 two_stage_opamp_dummy_magic_0.Vb2_2.n1 11.2576
R8980 two_stage_opamp_dummy_magic_0.Vb2_2.n1 two_stage_opamp_dummy_magic_0.Vb2_2.t8 11.2576
R8981 two_stage_opamp_dummy_magic_0.Vb2_2.n29 two_stage_opamp_dummy_magic_0.Vb2_2.n12 9.14336
R8982 two_stage_opamp_dummy_magic_0.Vb2_2.n25 two_stage_opamp_dummy_magic_0.Vb2_2.n24 9.14336
R8983 two_stage_opamp_dummy_magic_0.Vb2_2.n22 two_stage_opamp_dummy_magic_0.Vb2_2.n19 9.14336
R8984 two_stage_opamp_dummy_magic_0.Vb2_2.n35 two_stage_opamp_dummy_magic_0.Vb2_2.n3 9.14336
R8985 two_stage_opamp_dummy_magic_0.Vb2_2.n44 two_stage_opamp_dummy_magic_0.Vb2_2.n3 9.14336
R8986 two_stage_opamp_dummy_magic_0.Vb2_2.n44 two_stage_opamp_dummy_magic_0.Vb2_2.n43 9.14336
R8987 two_stage_opamp_dummy_magic_0.Vb2_2.n43 two_stage_opamp_dummy_magic_0.Vb2_2.n42 9.14336
R8988 two_stage_opamp_dummy_magic_0.Vb2_2.n37 two_stage_opamp_dummy_magic_0.Vb2_2.n36 5.33286
R8989 two_stage_opamp_dummy_magic_0.Vb2_2.n17 two_stage_opamp_dummy_magic_0.Vb2_2.n12 4.53698
R8990 two_stage_opamp_dummy_magic_0.Vb2_2.n24 two_stage_opamp_dummy_magic_0.Vb2_2.n23 4.53698
R8991 two_stage_opamp_dummy_magic_0.Vb2_2.n19 two_stage_opamp_dummy_magic_0.Vb2_2.n18 4.53698
R8992 two_stage_opamp_dummy_magic_0.Vb2_2.n25 two_stage_opamp_dummy_magic_0.Vb2_2.n17 4.53698
R8993 two_stage_opamp_dummy_magic_0.Vb2_2.n23 two_stage_opamp_dummy_magic_0.Vb2_2.n22 4.53698
R8994 two_stage_opamp_dummy_magic_0.Vb2_2.n33 two_stage_opamp_dummy_magic_0.Vb2_2.n32 4.5005
R8995 two_stage_opamp_dummy_magic_0.Vb2_2.n36 two_stage_opamp_dummy_magic_0.Vb2_2.n35 3.75335
R8996 two_stage_opamp_dummy_magic_0.Vb2_2.n42 two_stage_opamp_dummy_magic_0.Vb2_2.n41 3.75335
R8997 a_13180_23838.t0 a_13180_23838.t1 178.133
R8998 a_14170_5524.t0 a_14170_5524.t1 262.248
R8999 a_14290_5524.t0 a_14290_5524.t1 169.905
C0 m1_10050_19490# two_stage_opamp_dummy_magic_0.V_err_gate 0.091711f
C1 two_stage_opamp_dummy_magic_0.cap_res_X VDDA 0.39294f
C2 two_stage_opamp_dummy_magic_0.V_tail_gate VOUT- 0.020003f
C3 VIN+ VIN- 0.141796f
C4 two_stage_opamp_dummy_magic_0.VD4 VDDA 4.4335f
C5 two_stage_opamp_dummy_magic_0.Vb2 two_stage_opamp_dummy_magic_0.V_err_gate 2.11965f
C6 bgr_0.PFET_GATE_10uA VDDA 7.97055f
C7 m1_4880_3600# m2_4880_3600# 0.016063f
C8 bgr_0.V_TOP VDDA 13.2374f
C9 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C10 two_stage_opamp_dummy_magic_0.V_tail_gate VIN+ 0.054588f
C11 two_stage_opamp_dummy_magic_0.Vb2 bgr_0.START_UP 0.08188f
C12 bgr_0.V_TOP bgr_0.1st_Vout_1 2.47405f
C13 two_stage_opamp_dummy_magic_0.V_err_gate VOUT- 0.040291f
C14 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.Vb2 0.615754f
C15 two_stage_opamp_dummy_magic_0.V_tail_gate VIN- 0.158715f
C16 two_stage_opamp_dummy_magic_0.cap_res_X VOUT+ 0.037134f
C17 two_stage_opamp_dummy_magic_0.VD2 li_9020_5340# 0.070041f
C18 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.Vb2 1.23597f
C19 li_11100_5340# VIN- 0.024834f
C20 two_stage_opamp_dummy_magic_0.VD4 VOUT+ 0.023279f
C21 bgr_0.PFET_GATE_10uA m2_9370_16580# 0.012f
C22 bgr_0.PFET_GATE_10uA bgr_0.START_UP_NFET1 0.0108f
C23 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_tail_gate 0.038519f
C24 bgr_0.1st_Vout_1 VDDA 0.896465f
C25 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.Vb2 0.936691f
C26 two_stage_opamp_dummy_magic_0.cap_res_X VOUT- 51.0174f
C27 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_gate 1.39954f
C28 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.START_UP 1.36583f
C29 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 3.50895f
C30 bgr_0.START_UP_NFET1 VDDA 0.167059f
C31 two_stage_opamp_dummy_magic_0.Vb2 VDDA 1.51759f
C32 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_tail_gate 0.252494f
C33 VDDA VOUT+ 5.84986f
C34 bgr_0.NFET_GATE_10uA bgr_0.START_UP 1.64177f
C35 two_stage_opamp_dummy_magic_0.Vb2 bgr_0.1st_Vout_1 0.042752f
C36 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_0.V_TOP 0.055802f
C37 m1_10050_19490# two_stage_opamp_dummy_magic_0.Vb2 0.08176f
C38 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.506358f
C39 VDDA VOUT- 5.85294f
C40 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.V_tail_gate 0.241309f
C41 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.67032f
C42 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.583702f
C43 two_stage_opamp_dummy_magic_0.VD2 VIN+ 1.00457f
C44 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.046803f
C45 bgr_0.NFET_GATE_10uA bgr_0.PFET_GATE_10uA 0.012365f
C46 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.052756f
C47 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_tail_gate 0.269369f
C48 li_9020_5340# VIN+ 0.024834f
C49 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter m1_10050_19490# 0.013969f
C50 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.V_err_gate 0.333809f
C51 two_stage_opamp_dummy_magic_0.V_err_amp_ref VDDA 2.94626f
C52 two_stage_opamp_dummy_magic_0.Vb2 VOUT- 0.058721f
C53 VOUT+ VOUT- 0.397591f
C54 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.V_err_gate 0.010508f
C55 two_stage_opamp_dummy_magic_0.VD2 two_stage_opamp_dummy_magic_0.V_tail_gate 0.028539f
C56 bgr_0.NFET_GATE_10uA VDDA 0.818988f
C57 two_stage_opamp_dummy_magic_0.V_tail_gate VDDA 3.59138f
C58 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter two_stage_opamp_dummy_magic_0.Vb2 0.01158f
C59 bgr_0.NFET_GATE_10uA bgr_0.1st_Vout_1 0.03875f
C60 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_gate 0.08195f
C61 bgr_0.V_TOP m2_10730_16580# 0.012f
C62 bgr_0.V_TOP bgr_0.START_UP 0.792764f
C63 two_stage_opamp_dummy_magic_0.cap_res_X bgr_0.PFET_GATE_10uA 0.011459f
C64 two_stage_opamp_dummy_magic_0.V_err_amp_ref VOUT+ 0.042098f
C65 two_stage_opamp_dummy_magic_0.V_err_gate VDDA 2.00665f
C66 bgr_0.NFET_GATE_10uA bgr_0.START_UP_NFET1 0.351171f
C67 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.Vb2 0.538556f
C68 two_stage_opamp_dummy_magic_0.V_err_gate bgr_0.1st_Vout_1 0.041119f
C69 two_stage_opamp_dummy_magic_0.Vb2 two_stage_opamp_dummy_magic_0.V_tail_gate 0.084214f
C70 bgr_0.START_UP VDDA 1.09181f
C71 bgr_0.V_TOP bgr_0.PFET_GATE_10uA 0.221314f
C72 m2_10730_16580# bgr_0.1st_Vout_1 0.075543f
C73 bgr_0.START_UP bgr_0.1st_Vout_1 0.04354f
C74 VIN- GNDA 1.45233f
C75 VIN+ GNDA 1.46001f
C76 VOUT- GNDA 15.844832f
C77 VOUT+ GNDA 15.878867f
C78 VDDA GNDA 0.121269p
C79 m2_4880_3600# GNDA 0.05269f $ **FLOATING
C80 m2_10730_16580# GNDA 0.0105f $ **FLOATING
C81 m2_9370_16580# GNDA 0.010002f $ **FLOATING
C82 m1_4880_3600# GNDA 0.059696f $ **FLOATING
C83 m1_10050_19490# GNDA 0.259273f $ **FLOATING
C84 li_11100_5340# GNDA 0.022196f $ **FLOATING
C85 li_9020_5340# GNDA 0.022196f $ **FLOATING
C86 two_stage_opamp_dummy_magic_0.VD2 GNDA 2.13193f
C87 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 32.98453f
C88 two_stage_opamp_dummy_magic_0.V_tail_gate GNDA 8.285028f
C89 bgr_0.1st_Vout_1 GNDA 7.823503f
C90 bgr_0.START_UP GNDA 5.877827f
C91 bgr_0.START_UP_NFET1 GNDA 4.29564f
C92 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 10.25024f
C93 two_stage_opamp_dummy_magic_0.Vb2 GNDA 7.300634f
C94 bgr_0.NFET_GATE_10uA GNDA 7.92412f
C95 bgr_0.V_TOP GNDA 9.96016f
C96 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.8955f
C97 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 7.313879f
C98 bgr_0.PFET_GATE_10uA GNDA 6.602193f
C99 two_stage_opamp_dummy_magic_0.VD4 GNDA 4.871677f
C100 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.01637f
C101 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.01637f
C102 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.041034f
C103 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.01637f
C104 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.01637f
C105 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.040818f
C106 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.362787f
C107 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.01637f
C108 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.01637f
C109 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.03274f
C110 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.060887f
C111 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.206157f
C112 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.03274f
C113 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.03274f
C114 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.097293f
C115 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.03274f
C116 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.03274f
C117 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.096862f
C118 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.331325f
C119 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.03274f
C120 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.03274f
C121 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.096862f
C122 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.171607f
C123 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.03274f
C124 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.03274f
C125 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.096862f
C126 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.171607f
C127 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.03274f
C128 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.03274f
C129 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.096862f
C130 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.239231f
C131 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 1.32734f
C132 bgr_0.V_CMFB_S1 GNDA 1.1041f
C133 bgr_0.START_UP.t0 GNDA 1.06745f
C134 bgr_0.START_UP.t1 GNDA 0.02806f
C135 bgr_0.START_UP.n0 GNDA 0.714928f
C136 bgr_0.START_UP.t2 GNDA 0.026778f
C137 bgr_0.START_UP.t4 GNDA 0.026778f
C138 bgr_0.START_UP.n1 GNDA 0.097147f
C139 bgr_0.START_UP.t3 GNDA 0.026778f
C140 bgr_0.START_UP.t5 GNDA 0.026778f
C141 bgr_0.START_UP.n2 GNDA 0.08937f
C142 bgr_0.START_UP.n3 GNDA 0.462855f
C143 bgr_0.START_UP.t7 GNDA 0.010062f
C144 bgr_0.START_UP.t6 GNDA 0.010062f
C145 bgr_0.START_UP.n4 GNDA 0.028407f
C146 bgr_0.START_UP.n5 GNDA 0.260836f
C147 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.030951f
C148 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.030951f
C149 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.108702f
C150 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.030951f
C151 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.030951f
C152 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.108329f
C153 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.202138f
C154 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.030951f
C155 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.030951f
C156 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.108329f
C157 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.104793f
C158 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.030951f
C159 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.030951f
C160 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.108329f
C161 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.104793f
C162 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.030951f
C163 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.030951f
C164 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.108329f
C165 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.104793f
C166 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.030951f
C167 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.030951f
C168 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.108329f
C169 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.153987f
C170 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.030951f
C171 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.030951f
C172 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.10726f
C173 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.104977f
C174 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.030951f
C175 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.092854f
C176 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.030951f
C177 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.017686f
C178 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.014321f
C179 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.017686f
C180 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.054268f
C181 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.030951f
C182 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.030951f
C183 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.10726f
C184 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.104977f
C185 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.030951f
C186 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.030951f
C187 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.10726f
C188 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.104977f
C189 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.030951f
C190 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.030951f
C191 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.10726f
C192 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.104977f
C193 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.030951f
C194 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.030951f
C195 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.10726f
C196 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.134403f
C197 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.046089f
C198 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.030951f
C199 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.030951f
C200 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.017686f
C201 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.017686f
C202 two_stage_opamp_dummy_magic_0.VD4.n34 GNDA 0.030951f
C203 two_stage_opamp_dummy_magic_0.VD4.n36 GNDA 0.030951f
C204 two_stage_opamp_dummy_magic_0.VD4.n37 GNDA 0.017686f
C205 two_stage_opamp_dummy_magic_0.VD4.n38 GNDA 0.017686f
C206 two_stage_opamp_dummy_magic_0.VD4.n39 GNDA 0.030951f
C207 two_stage_opamp_dummy_magic_0.VD4.n40 GNDA 0.031222f
C208 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.030951f
C209 two_stage_opamp_dummy_magic_0.VD4.n41 GNDA 0.092854f
C210 two_stage_opamp_dummy_magic_0.VD4.n42 GNDA 0.029837f
C211 two_stage_opamp_dummy_magic_0.VD4.n43 GNDA 0.017686f
C212 two_stage_opamp_dummy_magic_0.VD4.n44 GNDA 0.258664f
C213 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.224175f
C214 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.206931f
C215 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.206931f
C216 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.206931f
C217 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.206931f
C218 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.206931f
C219 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.206931f
C220 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.206931f
C221 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.206931f
C222 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.206931f
C223 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.206931f
C224 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.224175f
C225 two_stage_opamp_dummy_magic_0.VD4.n46 GNDA 0.014321f
C226 two_stage_opamp_dummy_magic_0.VD4.n47 GNDA 0.017686f
C227 two_stage_opamp_dummy_magic_0.VD4.n49 GNDA 0.031222f
C228 two_stage_opamp_dummy_magic_0.VD4.n50 GNDA 0.030951f
C229 two_stage_opamp_dummy_magic_0.VD4.n51 GNDA 0.017686f
C230 two_stage_opamp_dummy_magic_0.VD4.n52 GNDA 0.017686f
C231 two_stage_opamp_dummy_magic_0.VD4.n53 GNDA 0.030951f
C232 two_stage_opamp_dummy_magic_0.VD4.n55 GNDA 0.030951f
C233 two_stage_opamp_dummy_magic_0.VD4.n56 GNDA 0.030951f
C234 two_stage_opamp_dummy_magic_0.VD4.n57 GNDA 0.017686f
C235 two_stage_opamp_dummy_magic_0.VD4.n58 GNDA 0.258664f
C236 two_stage_opamp_dummy_magic_0.VD4.n59 GNDA 0.013727f
C237 two_stage_opamp_dummy_magic_0.VD4.n60 GNDA 0.033797f
C238 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.054268f
C239 two_stage_opamp_dummy_magic_0.VD4.n61 GNDA 0.044756f
C240 two_stage_opamp_dummy_magic_0.VD4.n62 GNDA 0.062101f
C241 two_stage_opamp_dummy_magic_0.VD4.n63 GNDA 0.087485f
C242 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.01637f
C243 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.01637f
C244 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.041052f
C245 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.01637f
C246 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.01637f
C247 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.040835f
C248 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.363013f
C249 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.01637f
C250 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.01637f
C251 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.03274f
C252 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.060861f
C253 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.206157f
C254 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.03274f
C255 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.03274f
C256 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.097293f
C257 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.03274f
C258 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.03274f
C259 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.096862f
C260 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.331325f
C261 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.03274f
C262 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.03274f
C263 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.096862f
C264 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.171607f
C265 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.03274f
C266 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.03274f
C267 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.096862f
C268 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.171607f
C269 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.03274f
C270 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.03274f
C271 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.096862f
C272 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.239231f
C273 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 1.32734f
C274 bgr_0.V_CMFB_S3 GNDA 1.10386f
C275 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.066308f
C276 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.020237f
C277 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.966965f
C278 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.017268f
C279 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.017079f
C280 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.330906f
C281 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 0.017079f
C282 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 0.303032f
C283 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.018944f
C284 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.157213f
C285 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.177766f
C286 two_stage_opamp_dummy_magic_0.err_amp_out.n10 GNDA 0.020237f
C287 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.020156f
C288 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.020156f
C289 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.073261f
C290 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.020156f
C291 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.020156f
C292 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.060879f
C293 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 1.18743f
C294 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.247627f
C295 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.060467f
C296 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.060467f
C297 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.252232f
C298 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.060467f
C299 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.060467f
C300 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.251304f
C301 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.345024f
C302 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.060467f
C303 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.060467f
C304 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.251304f
C305 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.18003f
C306 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.060467f
C307 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.060467f
C308 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.251304f
C309 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 0.18003f
C310 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.060467f
C311 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.060467f
C312 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.251304f
C313 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.249769f
C314 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 1.34239f
C315 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n13 GNDA 1.98073f
C316 bgr_0.V_CMFB_S4 GNDA 0.010078f
C317 bgr_0.Vin-.n0 GNDA 0.069747f
C318 bgr_0.Vin-.n1 GNDA 0.316148f
C319 bgr_0.Vin-.t7 GNDA 0.027101f
C320 bgr_0.Vin-.t5 GNDA 0.027101f
C321 bgr_0.Vin-.n2 GNDA 0.094346f
C322 bgr_0.Vin-.t4 GNDA 0.027101f
C323 bgr_0.Vin-.t6 GNDA 0.027101f
C324 bgr_0.Vin-.n3 GNDA 0.090091f
C325 bgr_0.Vin-.n4 GNDA 0.386489f
C326 bgr_0.Vin-.n5 GNDA 0.027681f
C327 bgr_0.Vin-.n6 GNDA 0.366254f
C328 bgr_0.Vin-.t12 GNDA 0.022346f
C329 bgr_0.Vin-.n7 GNDA 0.026209f
C330 bgr_0.Vin-.n8 GNDA 0.021455f
C331 bgr_0.Vin-.n9 GNDA 0.021455f
C332 bgr_0.Vin-.n10 GNDA 0.036491f
C333 bgr_0.Vin-.n11 GNDA 0.497932f
C334 bgr_0.Vin-.t0 GNDA 0.117924f
C335 bgr_0.Vin-.n12 GNDA 0.655831f
C336 bgr_0.Vin-.n13 GNDA 1.07297f
C337 bgr_0.Vin-.n14 GNDA 0.471323f
C338 bgr_0.Vin-.t3 GNDA 0.261631f
C339 bgr_0.Vin-.n15 GNDA 0.069875f
C340 bgr_0.Vin-.n16 GNDA 0.119593f
C341 bgr_0.Vin-.n17 GNDA 0.07053f
C342 bgr_0.Vin-.n18 GNDA 0.579028f
C343 bgr_0.Vin-.n19 GNDA 0.358216f
C344 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.086538f
C345 bgr_0.V_mir2.t7 GNDA 0.019293f
C346 bgr_0.V_mir2.n0 GNDA 0.025223f
C347 bgr_0.V_mir2.t14 GNDA 0.041163f
C348 bgr_0.V_mir2.n1 GNDA 0.027381f
C349 bgr_0.V_mir2.n2 GNDA 0.451535f
C350 bgr_0.V_mir2.n3 GNDA 0.146338f
C351 bgr_0.V_mir2.t4 GNDA 0.023151f
C352 bgr_0.V_mir2.t17 GNDA 0.023151f
C353 bgr_0.V_mir2.t20 GNDA 0.037369f
C354 bgr_0.V_mir2.n4 GNDA 0.041731f
C355 bgr_0.V_mir2.n5 GNDA 0.028507f
C356 bgr_0.V_mir2.t0 GNDA 0.02939f
C357 bgr_0.V_mir2.n6 GNDA 0.044354f
C358 bgr_0.V_mir2.t5 GNDA 0.019293f
C359 bgr_0.V_mir2.t1 GNDA 0.019293f
C360 bgr_0.V_mir2.n7 GNDA 0.044166f
C361 bgr_0.V_mir2.n8 GNDA 0.109943f
C362 bgr_0.V_mir2.t2 GNDA 0.023151f
C363 bgr_0.V_mir2.t18 GNDA 0.023151f
C364 bgr_0.V_mir2.t22 GNDA 0.037369f
C365 bgr_0.V_mir2.n9 GNDA 0.041731f
C366 bgr_0.V_mir2.n10 GNDA 0.028507f
C367 bgr_0.V_mir2.t8 GNDA 0.02939f
C368 bgr_0.V_mir2.n11 GNDA 0.044354f
C369 bgr_0.V_mir2.t3 GNDA 0.019293f
C370 bgr_0.V_mir2.t9 GNDA 0.019293f
C371 bgr_0.V_mir2.n12 GNDA 0.044166f
C372 bgr_0.V_mir2.n13 GNDA 0.111042f
C373 bgr_0.V_mir2.n14 GNDA 0.381359f
C374 bgr_0.V_mir2.n15 GNDA 0.051125f
C375 bgr_0.V_mir2.t6 GNDA 0.023151f
C376 bgr_0.V_mir2.t19 GNDA 0.023151f
C377 bgr_0.V_mir2.t21 GNDA 0.037369f
C378 bgr_0.V_mir2.n16 GNDA 0.041731f
C379 bgr_0.V_mir2.n17 GNDA 0.028507f
C380 bgr_0.V_mir2.t10 GNDA 0.02939f
C381 bgr_0.V_mir2.n18 GNDA 0.044354f
C382 bgr_0.V_mir2.n19 GNDA 0.085095f
C383 bgr_0.V_mir2.n20 GNDA 0.044166f
C384 bgr_0.V_mir2.t11 GNDA 0.019293f
C385 bgr_0.cap_res1.t12 GNDA 0.331712f
C386 bgr_0.cap_res1.t19 GNDA 0.349187f
C387 bgr_0.cap_res1.t16 GNDA 0.350452f
C388 bgr_0.cap_res1.t5 GNDA 0.331712f
C389 bgr_0.cap_res1.t15 GNDA 0.349187f
C390 bgr_0.cap_res1.t9 GNDA 0.350452f
C391 bgr_0.cap_res1.t11 GNDA 0.331712f
C392 bgr_0.cap_res1.t18 GNDA 0.349187f
C393 bgr_0.cap_res1.t14 GNDA 0.350452f
C394 bgr_0.cap_res1.t4 GNDA 0.331712f
C395 bgr_0.cap_res1.t13 GNDA 0.349187f
C396 bgr_0.cap_res1.t7 GNDA 0.350452f
C397 bgr_0.cap_res1.t20 GNDA 0.331712f
C398 bgr_0.cap_res1.t6 GNDA 0.349187f
C399 bgr_0.cap_res1.t1 GNDA 0.350452f
C400 bgr_0.cap_res1.n0 GNDA 0.23406f
C401 bgr_0.cap_res1.t17 GNDA 0.186395f
C402 bgr_0.cap_res1.n1 GNDA 0.253961f
C403 bgr_0.cap_res1.t2 GNDA 0.186395f
C404 bgr_0.cap_res1.n2 GNDA 0.253961f
C405 bgr_0.cap_res1.t8 GNDA 0.186395f
C406 bgr_0.cap_res1.n3 GNDA 0.253961f
C407 bgr_0.cap_res1.t3 GNDA 0.186395f
C408 bgr_0.cap_res1.n4 GNDA 0.253961f
C409 bgr_0.cap_res1.t10 GNDA 0.363549f
C410 bgr_0.cap_res1.t0 GNDA 0.08421f
C411 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.011089f
C412 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.011089f
C413 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.027759f
C414 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.011089f
C415 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.011089f
C416 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.027759f
C417 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.011089f
C418 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.011089f
C419 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.02761f
C420 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.187477f
C421 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.157474f
C422 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.011089f
C423 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.011089f
C424 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.022178f
C425 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.039374f
C426 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.016633f
C427 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.016633f
C428 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.056318f
C429 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.029524f
C430 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.029524f
C431 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.029524f
C432 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.029524f
C433 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.029524f
C434 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.029524f
C435 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.029524f
C436 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.029524f
C437 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.029524f
C438 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.034459f
C439 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.03249f
C440 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.020376f
C441 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.020376f
C442 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.020376f
C443 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.020376f
C444 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.020376f
C445 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.020376f
C446 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.020376f
C447 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.018217f
C448 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.029524f
C449 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.029524f
C450 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.029524f
C451 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.029524f
C452 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.029524f
C453 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.029524f
C454 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.029524f
C455 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.029524f
C456 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.029524f
C457 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.034459f
C458 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.03249f
C459 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.020376f
C460 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.020376f
C461 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.020376f
C462 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.020376f
C463 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.020376f
C464 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.020376f
C465 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.020376f
C466 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.018217f
C467 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.017179f
C468 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.247131f
C469 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.016633f
C470 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.016633f
C471 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.033267f
C472 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 0.053323f
C473 bgr_0.PFET_GATE_10uA.t28 GNDA 0.020856f
C474 bgr_0.PFET_GATE_10uA.t20 GNDA 0.030831f
C475 bgr_0.PFET_GATE_10uA.n0 GNDA 0.033972f
C476 bgr_0.PFET_GATE_10uA.t15 GNDA 0.020856f
C477 bgr_0.PFET_GATE_10uA.t21 GNDA 0.030831f
C478 bgr_0.PFET_GATE_10uA.n1 GNDA 0.033972f
C479 bgr_0.PFET_GATE_10uA.n2 GNDA 0.040878f
C480 bgr_0.PFET_GATE_10uA.t19 GNDA 0.020856f
C481 bgr_0.PFET_GATE_10uA.t12 GNDA 0.030831f
C482 bgr_0.PFET_GATE_10uA.n3 GNDA 0.033972f
C483 bgr_0.PFET_GATE_10uA.t26 GNDA 0.020856f
C484 bgr_0.PFET_GATE_10uA.t13 GNDA 0.030831f
C485 bgr_0.PFET_GATE_10uA.n4 GNDA 0.033972f
C486 bgr_0.PFET_GATE_10uA.n5 GNDA 0.034081f
C487 bgr_0.PFET_GATE_10uA.t7 GNDA 0.312465f
C488 bgr_0.PFET_GATE_10uA.t0 GNDA 0.021391f
C489 bgr_0.PFET_GATE_10uA.t8 GNDA 0.021391f
C490 bgr_0.PFET_GATE_10uA.n6 GNDA 0.054673f
C491 bgr_0.PFET_GATE_10uA.t2 GNDA 0.021391f
C492 bgr_0.PFET_GATE_10uA.t4 GNDA 0.021391f
C493 bgr_0.PFET_GATE_10uA.n7 GNDA 0.05326f
C494 bgr_0.PFET_GATE_10uA.n8 GNDA 0.520952f
C495 bgr_0.PFET_GATE_10uA.t3 GNDA 0.021391f
C496 bgr_0.PFET_GATE_10uA.t5 GNDA 0.021391f
C497 bgr_0.PFET_GATE_10uA.n9 GNDA 0.05326f
C498 bgr_0.PFET_GATE_10uA.n10 GNDA 0.295408f
C499 bgr_0.PFET_GATE_10uA.n11 GNDA 0.603055f
C500 bgr_0.PFET_GATE_10uA.t9 GNDA 0.021391f
C501 bgr_0.PFET_GATE_10uA.t1 GNDA 0.021391f
C502 bgr_0.PFET_GATE_10uA.n12 GNDA 0.05159f
C503 bgr_0.PFET_GATE_10uA.n13 GNDA 0.275411f
C504 bgr_0.PFET_GATE_10uA.t6 GNDA 0.464967f
C505 bgr_0.PFET_GATE_10uA.t27 GNDA 0.024114f
C506 bgr_0.PFET_GATE_10uA.t14 GNDA 0.024114f
C507 bgr_0.PFET_GATE_10uA.n14 GNDA 0.069715f
C508 bgr_0.PFET_GATE_10uA.n15 GNDA 1.91969f
C509 bgr_0.PFET_GATE_10uA.n16 GNDA 0.771508f
C510 bgr_0.PFET_GATE_10uA.n17 GNDA 0.759224f
C511 bgr_0.PFET_GATE_10uA.t11 GNDA 0.020856f
C512 bgr_0.PFET_GATE_10uA.t25 GNDA 0.020856f
C513 bgr_0.PFET_GATE_10uA.t18 GNDA 0.020856f
C514 bgr_0.PFET_GATE_10uA.t10 GNDA 0.020856f
C515 bgr_0.PFET_GATE_10uA.t24 GNDA 0.020856f
C516 bgr_0.PFET_GATE_10uA.t17 GNDA 0.030831f
C517 bgr_0.PFET_GATE_10uA.n18 GNDA 0.038154f
C518 bgr_0.PFET_GATE_10uA.n19 GNDA 0.027273f
C519 bgr_0.PFET_GATE_10uA.n20 GNDA 0.027273f
C520 bgr_0.PFET_GATE_10uA.n21 GNDA 0.027273f
C521 bgr_0.PFET_GATE_10uA.n22 GNDA 0.023091f
C522 bgr_0.PFET_GATE_10uA.t16 GNDA 0.020856f
C523 bgr_0.PFET_GATE_10uA.t23 GNDA 0.020856f
C524 bgr_0.PFET_GATE_10uA.t22 GNDA 0.020856f
C525 bgr_0.PFET_GATE_10uA.t29 GNDA 0.030831f
C526 bgr_0.PFET_GATE_10uA.n23 GNDA 0.038154f
C527 bgr_0.PFET_GATE_10uA.n24 GNDA 0.027273f
C528 bgr_0.PFET_GATE_10uA.n25 GNDA 0.023091f
C529 bgr_0.PFET_GATE_10uA.n26 GNDA 0.031695f
C530 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 0.425161f
C531 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 0.662076f
C532 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.020481f
C533 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.031939f
C534 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.024921f
C535 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.024921f
C536 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.024921f
C537 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.024921f
C538 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.024921f
C539 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.024921f
C540 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.02046f
C541 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.020481f
C542 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.031939f
C543 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.024921f
C544 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.024921f
C545 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.024921f
C546 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.024921f
C547 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.024921f
C548 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.024921f
C549 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.024921f
C550 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.024921f
C551 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.02046f
C552 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.034783f
C553 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.022916f
C554 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.022916f
C555 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.348451f
C556 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.011458f
C557 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.011458f
C558 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.02698f
C559 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.011458f
C560 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.011458f
C561 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.026798f
C562 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.011458f
C563 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.011458f
C564 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.026798f
C565 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.011458f
C566 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.011458f
C567 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.026798f
C568 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.011458f
C569 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.011458f
C570 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.026798f
C571 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.011458f
C572 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.011458f
C573 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.026647f
C574 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.331264f
C575 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.013493f
C576 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.013493f
C577 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.049393f
C578 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.013493f
C579 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.013493f
C580 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.048979f
C581 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.179573f
C582 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.013493f
C583 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.013493f
C584 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.048979f
C585 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.093142f
C586 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.013493f
C587 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.013493f
C588 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.048979f
C589 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.093142f
C590 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.013493f
C591 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.013493f
C592 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.048979f
C593 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.093142f
C594 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.013493f
C595 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.013493f
C596 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.048979f
C597 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.112031f
C598 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.031482f
C599 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.031482f
C600 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.110568f
C601 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.031482f
C602 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.031482f
C603 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.110188f
C604 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.205607f
C605 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.031482f
C606 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.031482f
C607 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.110188f
C608 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.106591f
C609 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.031482f
C610 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.031482f
C611 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.110188f
C612 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.106591f
C613 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.031482f
C614 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.031482f
C615 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.110188f
C616 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.125547f
C617 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.031482f
C618 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.031482f
C619 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.107979f
C620 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.184593f
C621 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.018889f
C622 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.018889f
C623 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.018889f
C624 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.022937f
C625 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.022937f
C626 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.014842f
C627 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.013091f
C628 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.018889f
C629 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.018889f
C630 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.018889f
C631 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.018889f
C632 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.018889f
C633 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.022937f
C634 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.022937f
C635 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.014842f
C636 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.014842f
C637 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.014842f
C638 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.013091f
C639 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.013602f
C640 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.029009f
C641 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.029009f
C642 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.029009f
C643 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.032978f
C644 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.029762f
C645 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.018215f
C646 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.016464f
C647 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.029009f
C648 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.029009f
C649 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.029009f
C650 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.029009f
C651 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.029009f
C652 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.032978f
C653 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.029762f
C654 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.018215f
C655 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.018215f
C656 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.018215f
C657 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.016464f
C658 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.013602f
C659 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.121373f
C660 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.290786f
C661 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.075108f
C662 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.059367f
C663 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.059367f
C664 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.059367f
C665 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.059367f
C666 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.06323f
C667 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.050107f
C668 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.028334f
C669 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.028334f
C670 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.02659f
C671 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.059367f
C672 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.059367f
C673 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.059367f
C674 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.059367f
C675 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.06323f
C676 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.050107f
C677 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.028334f
C678 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.028334f
C679 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 0.02659f
C680 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.016175f
C681 two_stage_opamp_dummy_magic_0.Y.n52 GNDA 0.478888f
C682 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.437339f
C683 two_stage_opamp_dummy_magic_0.Vb2.t32 GNDA 0.043632f
C684 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.043632f
C685 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.043632f
C686 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.043632f
C687 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.050351f
C688 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.04088f
C689 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.025122f
C690 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.025122f
C691 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.023309f
C692 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.043632f
C693 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.043632f
C694 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.043632f
C695 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.043632f
C696 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.050351f
C697 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.04088f
C698 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.025122f
C699 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.025122f
C700 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.023309f
C701 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.013512f
C702 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.043632f
C703 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.043632f
C704 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.043632f
C705 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.043632f
C706 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.050351f
C707 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.04088f
C708 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.025122f
C709 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.025122f
C710 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.023309f
C711 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.043632f
C712 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.043632f
C713 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.043632f
C714 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.043632f
C715 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.050351f
C716 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.04088f
C717 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.025122f
C718 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.025122f
C719 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.023309f
C720 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.016397f
C721 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.03003f
C722 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.029147f
C723 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.303104f
C724 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.029147f
C725 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 0.204441f
C726 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.029147f
C727 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.808923f
C728 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.053353f
C729 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.723168f
C730 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.030851f
C731 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.030851f
C732 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.107063f
C733 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.053353f
C734 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.18525f
C735 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.031502f
C736 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.094361f
C737 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.154162f
C738 two_stage_opamp_dummy_magic_0.Vb2.n30 GNDA 0.287807f
C739 bgr_0.cap_res2.t6 GNDA 0.358376f
C740 bgr_0.cap_res2.t12 GNDA 0.359675f
C741 bgr_0.cap_res2.t14 GNDA 0.340442f
C742 bgr_0.cap_res2.t0 GNDA 0.358376f
C743 bgr_0.cap_res2.t5 GNDA 0.359675f
C744 bgr_0.cap_res2.t8 GNDA 0.340442f
C745 bgr_0.cap_res2.t4 GNDA 0.358376f
C746 bgr_0.cap_res2.t10 GNDA 0.359675f
C747 bgr_0.cap_res2.t13 GNDA 0.340442f
C748 bgr_0.cap_res2.t19 GNDA 0.358376f
C749 bgr_0.cap_res2.t3 GNDA 0.359675f
C750 bgr_0.cap_res2.t7 GNDA 0.340442f
C751 bgr_0.cap_res2.t15 GNDA 0.358376f
C752 bgr_0.cap_res2.t18 GNDA 0.359675f
C753 bgr_0.cap_res2.t1 GNDA 0.340442f
C754 bgr_0.cap_res2.n0 GNDA 0.24022f
C755 bgr_0.cap_res2.t2 GNDA 0.1913f
C756 bgr_0.cap_res2.n1 GNDA 0.260644f
C757 bgr_0.cap_res2.t9 GNDA 0.1913f
C758 bgr_0.cap_res2.n2 GNDA 0.260644f
C759 bgr_0.cap_res2.t16 GNDA 0.1913f
C760 bgr_0.cap_res2.n3 GNDA 0.260644f
C761 bgr_0.cap_res2.t11 GNDA 0.1913f
C762 bgr_0.cap_res2.n4 GNDA 0.260644f
C763 bgr_0.cap_res2.t17 GNDA 0.373116f
C764 bgr_0.cap_res2.t20 GNDA 0.086426f
C765 bgr_0.1st_Vout_2.n0 GNDA 0.723004f
C766 bgr_0.1st_Vout_2.n1 GNDA 0.237573f
C767 bgr_0.1st_Vout_2.n2 GNDA 1.43086f
C768 bgr_0.1st_Vout_2.n3 GNDA 0.104399f
C769 bgr_0.1st_Vout_2.n4 GNDA 1.45767f
C770 bgr_0.1st_Vout_2.n5 GNDA 0.010417f
C771 bgr_0.1st_Vout_2.t4 GNDA 0.015189f
C772 bgr_0.1st_Vout_2.n6 GNDA 0.157567f
C773 bgr_0.1st_Vout_2.t33 GNDA 0.017308f
C774 bgr_0.1st_Vout_2.n8 GNDA 0.018179f
C775 bgr_0.1st_Vout_2.t24 GNDA 0.010986f
C776 bgr_0.1st_Vout_2.t13 GNDA 0.010986f
C777 bgr_0.1st_Vout_2.n9 GNDA 0.024439f
C778 bgr_0.1st_Vout_2.t28 GNDA 0.288462f
C779 bgr_0.1st_Vout_2.t17 GNDA 0.293375f
C780 bgr_0.1st_Vout_2.t12 GNDA 0.288462f
C781 bgr_0.1st_Vout_2.t32 GNDA 0.288462f
C782 bgr_0.1st_Vout_2.t35 GNDA 0.293375f
C783 bgr_0.1st_Vout_2.t11 GNDA 0.293375f
C784 bgr_0.1st_Vout_2.t31 GNDA 0.288462f
C785 bgr_0.1st_Vout_2.t23 GNDA 0.288462f
C786 bgr_0.1st_Vout_2.t26 GNDA 0.293375f
C787 bgr_0.1st_Vout_2.t30 GNDA 0.293375f
C788 bgr_0.1st_Vout_2.t22 GNDA 0.288462f
C789 bgr_0.1st_Vout_2.t15 GNDA 0.288462f
C790 bgr_0.1st_Vout_2.t19 GNDA 0.293375f
C791 bgr_0.1st_Vout_2.t36 GNDA 0.293375f
C792 bgr_0.1st_Vout_2.t29 GNDA 0.288462f
C793 bgr_0.1st_Vout_2.t21 GNDA 0.288462f
C794 bgr_0.1st_Vout_2.t25 GNDA 0.293375f
C795 bgr_0.1st_Vout_2.t18 GNDA 0.293375f
C796 bgr_0.1st_Vout_2.t14 GNDA 0.288462f
C797 bgr_0.1st_Vout_2.t20 GNDA 0.288462f
C798 bgr_0.1st_Vout_2.t34 GNDA 0.018845f
C799 bgr_0.1st_Vout_2.n10 GNDA 0.018179f
C800 bgr_0.1st_Vout_2.t27 GNDA 0.010986f
C801 bgr_0.1st_Vout_2.t16 GNDA 0.010986f
C802 bgr_0.1st_Vout_2.n11 GNDA 0.024439f
C803 bgr_0.1st_Vout_2.n12 GNDA 0.017425f
C804 bgr_0.1st_Vout_1.n0 GNDA 0.538712f
C805 bgr_0.1st_Vout_1.n1 GNDA 0.236313f
C806 bgr_0.1st_Vout_1.n2 GNDA 0.973284f
C807 bgr_0.1st_Vout_1.n3 GNDA 0.907198f
C808 bgr_0.1st_Vout_1.n4 GNDA 0.891647f
C809 bgr_0.1st_Vout_1.t11 GNDA 0.358463f
C810 bgr_0.1st_Vout_1.t15 GNDA 0.35246f
C811 bgr_0.1st_Vout_1.t29 GNDA 0.358463f
C812 bgr_0.1st_Vout_1.t35 GNDA 0.35246f
C813 bgr_0.1st_Vout_1.t31 GNDA 0.358463f
C814 bgr_0.1st_Vout_1.t34 GNDA 0.35246f
C815 bgr_0.1st_Vout_1.t20 GNDA 0.358463f
C816 bgr_0.1st_Vout_1.t28 GNDA 0.35246f
C817 bgr_0.1st_Vout_1.t24 GNDA 0.358463f
C818 bgr_0.1st_Vout_1.t27 GNDA 0.35246f
C819 bgr_0.1st_Vout_1.t14 GNDA 0.358463f
C820 bgr_0.1st_Vout_1.t19 GNDA 0.35246f
C821 bgr_0.1st_Vout_1.t30 GNDA 0.358463f
C822 bgr_0.1st_Vout_1.t33 GNDA 0.35246f
C823 bgr_0.1st_Vout_1.t18 GNDA 0.358463f
C824 bgr_0.1st_Vout_1.t26 GNDA 0.35246f
C825 bgr_0.1st_Vout_1.t23 GNDA 0.358463f
C826 bgr_0.1st_Vout_1.t25 GNDA 0.35246f
C827 bgr_0.1st_Vout_1.t17 GNDA 0.35246f
C828 bgr_0.1st_Vout_1.t12 GNDA 0.35246f
C829 bgr_0.1st_Vout_1.t21 GNDA 0.023025f
C830 bgr_0.1st_Vout_1.n5 GNDA 0.715456f
C831 bgr_0.1st_Vout_1.n6 GNDA 0.022212f
C832 bgr_0.1st_Vout_1.n7 GNDA 0.104674f
C833 bgr_0.1st_Vout_1.t36 GNDA 0.013423f
C834 bgr_0.1st_Vout_1.t16 GNDA 0.013423f
C835 bgr_0.1st_Vout_1.n8 GNDA 0.029862f
C836 bgr_0.1st_Vout_1.n9 GNDA 0.082514f
C837 bgr_0.1st_Vout_1.t8 GNDA 0.018559f
C838 bgr_0.1st_Vout_1.n10 GNDA 0.012728f
C839 bgr_0.1st_Vout_1.n11 GNDA 0.192525f
C840 bgr_0.1st_Vout_1.n12 GNDA 0.011517f
C841 bgr_0.1st_Vout_1.n13 GNDA 0.048842f
C842 bgr_0.1st_Vout_1.n14 GNDA 0.021291f
C843 bgr_0.1st_Vout_1.n15 GNDA 0.078719f
C844 bgr_0.1st_Vout_1.n16 GNDA 0.038771f
C845 bgr_0.1st_Vout_1.t32 GNDA 0.013423f
C846 bgr_0.1st_Vout_1.t22 GNDA 0.013423f
C847 bgr_0.1st_Vout_1.n17 GNDA 0.029862f
C848 bgr_0.1st_Vout_1.n18 GNDA 0.082514f
C849 bgr_0.1st_Vout_1.n19 GNDA 0.022212f
C850 bgr_0.1st_Vout_1.n20 GNDA 0.104674f
C851 bgr_0.1st_Vout_1.t13 GNDA 0.021069f
C852 bgr_0.V_mir1.t7 GNDA 0.019293f
C853 bgr_0.V_mir1.t0 GNDA 0.02939f
C854 bgr_0.V_mir1.t4 GNDA 0.023151f
C855 bgr_0.V_mir1.t18 GNDA 0.023151f
C856 bgr_0.V_mir1.t20 GNDA 0.037369f
C857 bgr_0.V_mir1.n0 GNDA 0.041731f
C858 bgr_0.V_mir1.n1 GNDA 0.028507f
C859 bgr_0.V_mir1.n2 GNDA 0.044354f
C860 bgr_0.V_mir1.t1 GNDA 0.019293f
C861 bgr_0.V_mir1.t5 GNDA 0.019293f
C862 bgr_0.V_mir1.n3 GNDA 0.044166f
C863 bgr_0.V_mir1.n4 GNDA 0.109943f
C864 bgr_0.V_mir1.n5 GNDA 0.025223f
C865 bgr_0.V_mir1.t12 GNDA 0.041163f
C866 bgr_0.V_mir1.n6 GNDA 0.027381f
C867 bgr_0.V_mir1.n7 GNDA 0.451535f
C868 bgr_0.V_mir1.n8 GNDA 0.146338f
C869 bgr_0.V_mir1.t2 GNDA 0.02939f
C870 bgr_0.V_mir1.t8 GNDA 0.023151f
C871 bgr_0.V_mir1.t17 GNDA 0.023151f
C872 bgr_0.V_mir1.t21 GNDA 0.037369f
C873 bgr_0.V_mir1.n9 GNDA 0.041731f
C874 bgr_0.V_mir1.n10 GNDA 0.028507f
C875 bgr_0.V_mir1.n11 GNDA 0.044354f
C876 bgr_0.V_mir1.t3 GNDA 0.019293f
C877 bgr_0.V_mir1.t9 GNDA 0.019293f
C878 bgr_0.V_mir1.n12 GNDA 0.044166f
C879 bgr_0.V_mir1.n13 GNDA 0.085095f
C880 bgr_0.V_mir1.n14 GNDA 0.051125f
C881 bgr_0.V_mir1.n15 GNDA 0.381359f
C882 bgr_0.V_mir1.t6 GNDA 0.02939f
C883 bgr_0.V_mir1.t10 GNDA 0.023151f
C884 bgr_0.V_mir1.t22 GNDA 0.023151f
C885 bgr_0.V_mir1.t19 GNDA 0.037369f
C886 bgr_0.V_mir1.n16 GNDA 0.041731f
C887 bgr_0.V_mir1.n17 GNDA 0.028507f
C888 bgr_0.V_mir1.n18 GNDA 0.044354f
C889 bgr_0.V_mir1.n19 GNDA 0.111042f
C890 bgr_0.V_mir1.n20 GNDA 0.044166f
C891 bgr_0.V_mir1.t11 GNDA 0.019293f
C892 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.030951f
C893 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.030951f
C894 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.030951f
C895 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.108702f
C896 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.030951f
C897 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.030951f
C898 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.108329f
C899 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.202138f
C900 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.030951f
C901 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.030951f
C902 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.108329f
C903 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.104793f
C904 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.030951f
C905 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.030951f
C906 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.108329f
C907 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.104793f
C908 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.030951f
C909 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.030951f
C910 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.108329f
C911 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.104793f
C912 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.030951f
C913 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.030951f
C914 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.10726f
C915 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.104977f
C916 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.030951f
C917 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.092854f
C918 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.030951f
C919 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.017686f
C920 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.014321f
C921 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.014321f
C922 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.017686f
C923 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.054268f
C924 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.030951f
C925 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.030951f
C926 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.10726f
C927 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.104977f
C928 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.030951f
C929 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.030951f
C930 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.10726f
C931 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.104977f
C932 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.030951f
C933 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.030951f
C934 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.10726f
C935 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.104977f
C936 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.030951f
C937 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.030951f
C938 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.10726f
C939 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.134403f
C940 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.046089f
C941 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.030951f
C942 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.092854f
C943 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.031222f
C944 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.030951f
C945 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.017686f
C946 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.017686f
C947 two_stage_opamp_dummy_magic_0.VD3.n34 GNDA 0.030951f
C948 two_stage_opamp_dummy_magic_0.VD3.n36 GNDA 0.030951f
C949 two_stage_opamp_dummy_magic_0.VD3.n37 GNDA 0.017686f
C950 two_stage_opamp_dummy_magic_0.VD3.n38 GNDA 0.017686f
C951 two_stage_opamp_dummy_magic_0.VD3.n39 GNDA 0.030951f
C952 two_stage_opamp_dummy_magic_0.VD3.n41 GNDA 0.030951f
C953 two_stage_opamp_dummy_magic_0.VD3.n42 GNDA 0.029837f
C954 two_stage_opamp_dummy_magic_0.VD3.n43 GNDA 0.017686f
C955 two_stage_opamp_dummy_magic_0.VD3.n44 GNDA 0.258664f
C956 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.224175f
C957 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.206931f
C958 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.206931f
C959 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.206931f
C960 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.206931f
C961 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.206931f
C962 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.206931f
C963 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.206931f
C964 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.206931f
C965 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.206931f
C966 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.206931f
C967 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.224175f
C968 two_stage_opamp_dummy_magic_0.VD3.n45 GNDA 0.017686f
C969 two_stage_opamp_dummy_magic_0.VD3.n47 GNDA 0.031222f
C970 two_stage_opamp_dummy_magic_0.VD3.n48 GNDA 0.030951f
C971 two_stage_opamp_dummy_magic_0.VD3.n49 GNDA 0.017686f
C972 two_stage_opamp_dummy_magic_0.VD3.n50 GNDA 0.017686f
C973 two_stage_opamp_dummy_magic_0.VD3.n51 GNDA 0.030951f
C974 two_stage_opamp_dummy_magic_0.VD3.n53 GNDA 0.030951f
C975 two_stage_opamp_dummy_magic_0.VD3.n54 GNDA 0.030951f
C976 two_stage_opamp_dummy_magic_0.VD3.n55 GNDA 0.017686f
C977 two_stage_opamp_dummy_magic_0.VD3.n56 GNDA 0.258664f
C978 two_stage_opamp_dummy_magic_0.VD3.n57 GNDA 0.013727f
C979 two_stage_opamp_dummy_magic_0.VD3.n58 GNDA 0.033797f
C980 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.054268f
C981 two_stage_opamp_dummy_magic_0.VD3.n59 GNDA 0.044756f
C982 two_stage_opamp_dummy_magic_0.VD3.n60 GNDA 0.117031f
C983 two_stage_opamp_dummy_magic_0.VD3.n61 GNDA 0.19008f
C984 two_stage_opamp_dummy_magic_0.VD3.n62 GNDA 0.108328f
C985 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.030951f
C986 bgr_0.Vin+.t5 GNDA 0.173951f
C987 bgr_0.Vin+.t7 GNDA 0.010696f
C988 bgr_0.Vin+.t8 GNDA 0.025367f
C989 bgr_0.Vin+.t9 GNDA 0.01649f
C990 bgr_0.Vin+.n0 GNDA 0.054406f
C991 bgr_0.Vin+.t6 GNDA 0.01649f
C992 bgr_0.Vin+.n1 GNDA 0.042338f
C993 bgr_0.Vin+.t10 GNDA 0.01649f
C994 bgr_0.Vin+.n2 GNDA 0.042909f
C995 bgr_0.Vin+.n3 GNDA 0.130793f
C996 bgr_0.Vin+.t3 GNDA 0.05348f
C997 bgr_0.Vin+.t2 GNDA 0.05348f
C998 bgr_0.Vin+.n4 GNDA 0.176679f
C999 bgr_0.Vin+.n5 GNDA 1.27851f
C1000 bgr_0.Vin+.t1 GNDA 0.05348f
C1001 bgr_0.Vin+.t4 GNDA 0.05348f
C1002 bgr_0.Vin+.n6 GNDA 0.176679f
C1003 bgr_0.Vin+.n7 GNDA 1.06525f
C1004 bgr_0.Vin+.n8 GNDA 1.7265f
C1005 bgr_0.Vin+.t0 GNDA 0.232527f
C1006 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.017554f
C1007 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.011801f
C1008 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.030621f
C1009 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.15121f
C1010 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.010848f
C1011 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.024352f
C1012 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.149641f
C1013 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.017387f
C1014 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.144462f
C1015 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.011801f
C1016 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 0.030621f
C1017 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.083799f
C1018 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.010848f
C1019 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.024352f
C1020 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.108915f
C1021 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.200033f
C1022 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.031281f
C1023 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.011697f
C1024 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 0.036688f
C1025 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.011697f
C1026 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 0.030033f
C1027 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.011697f
C1028 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.030033f
C1029 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.011697f
C1030 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.052058f
C1031 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 1.04078f
C1032 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.037936f
C1033 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.037936f
C1034 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.13361f
C1035 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.037936f
C1036 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.037936f
C1037 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.127125f
C1038 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.594097f
C1039 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.037936f
C1040 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.037936f
C1041 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.127125f
C1042 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.424825f
C1043 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.839127f
C1044 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.105955f
C1045 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.265252f
C1046 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.265252f
C1047 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.314813f
C1048 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.166282f
C1049 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.105267f
C1050 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.287351f
C1051 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.102656f
C1052 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.487173f
C1053 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.287351f
C1054 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.265252f
C1055 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.265252f
C1056 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.314813f
C1057 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.166282f
C1058 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.105267f
C1059 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.102656f
C1060 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.487173f
C1061 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.105955f
C1062 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.019639f
C1063 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.019639f
C1064 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.071382f
C1065 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.019639f
C1066 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.019639f
C1067 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.059318f
C1068 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 1.15698f
C1069 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.241277f
C1070 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.058917f
C1071 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.058917f
C1072 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.245765f
C1073 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.058917f
C1074 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.058917f
C1075 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.244861f
C1076 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.336177f
C1077 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.058917f
C1078 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.058917f
C1079 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.244861f
C1080 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.175414f
C1081 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.058917f
C1082 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.058917f
C1083 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.244861f
C1084 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 0.175414f
C1085 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.058917f
C1086 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.058917f
C1087 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.244861f
C1088 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.243365f
C1089 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 1.30797f
C1090 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n13 GNDA 1.92994f
C1091 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.345142f
C1092 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.346293f
C1093 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.186001f
C1094 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.198613f
C1095 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.345142f
C1096 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.346293f
C1097 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.186001f
C1098 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.217197f
C1099 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.345142f
C1100 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.346293f
C1101 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.186001f
C1102 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.217197f
C1103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.345142f
C1104 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.346293f
C1105 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.186001f
C1106 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.217197f
C1107 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.345142f
C1108 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.346293f
C1109 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.364878f
C1110 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.364878f
C1111 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.186001f
C1112 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.217197f
C1113 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.345142f
C1114 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.346293f
C1115 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.364878f
C1116 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.364878f
C1117 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.186001f
C1118 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.217197f
C1119 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.346293f
C1120 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.347548f
C1121 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.346293f
C1122 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.349008f
C1123 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.379597f
C1124 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.328964f
C1125 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.346293f
C1126 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.347548f
C1127 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.328964f
C1128 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.346293f
C1129 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.347548f
C1130 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.346293f
C1131 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.347548f
C1132 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.346293f
C1133 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.347548f
C1134 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.346293f
C1135 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.347548f
C1136 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.346293f
C1137 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.347548f
C1138 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.346293f
C1139 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.347548f
C1140 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.346293f
C1141 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.347548f
C1142 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.346293f
C1143 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.347548f
C1144 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.346293f
C1145 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.347548f
C1146 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.346293f
C1147 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.347548f
C1148 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.346293f
C1149 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.347548f
C1150 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.346293f
C1151 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.347548f
C1152 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.346293f
C1153 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.347548f
C1154 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.346293f
C1155 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.347548f
C1156 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.346293f
C1157 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.347548f
C1158 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.346293f
C1159 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.347548f
C1160 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.346293f
C1161 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.347548f
C1162 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.346293f
C1163 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.347548f
C1164 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.346293f
C1165 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.347548f
C1166 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.346293f
C1167 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.347548f
C1168 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.346293f
C1169 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.347548f
C1170 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.346293f
C1171 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.347548f
C1172 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.346293f
C1173 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.347548f
C1174 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.346293f
C1175 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.347548f
C1176 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.346293f
C1177 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.347548f
C1178 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.345142f
C1179 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.346293f
C1180 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.186001f
C1181 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.198613f
C1182 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.345142f
C1183 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.346293f
C1184 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.186001f
C1185 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.217197f
C1186 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.345142f
C1187 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.346293f
C1188 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.186001f
C1189 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.217197f
C1190 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.345142f
C1191 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.346293f
C1192 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.186001f
C1193 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.217197f
C1194 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.345142f
C1195 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.346293f
C1196 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.186001f
C1197 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.217197f
C1198 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.345142f
C1199 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.346293f
C1200 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.186001f
C1201 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.217197f
C1202 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.345142f
C1203 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.346293f
C1204 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.186001f
C1205 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.217197f
C1206 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.346293f
C1207 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.186001f
C1208 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.197462f
C1209 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.346293f
C1210 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.186001f
C1211 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.197462f
C1212 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.346293f
C1213 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.347548f
C1214 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.346293f
C1215 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.347548f
C1216 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.167416f
C1217 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.215942f
C1218 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.18485f
C1219 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.234527f
C1220 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.18485f
C1221 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.251856f
C1222 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.18485f
C1223 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.251856f
C1224 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.18485f
C1225 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.251856f
C1226 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.18485f
C1227 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.251856f
C1228 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.18485f
C1229 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.251856f
C1230 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.18485f
C1231 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.251856f
C1232 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.18485f
C1233 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.251856f
C1234 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.18485f
C1235 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.251856f
C1236 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.18485f
C1237 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.251856f
C1238 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.18485f
C1239 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.251856f
C1240 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.18485f
C1241 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.251856f
C1242 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.18485f
C1243 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.251856f
C1244 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.18485f
C1245 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.251856f
C1246 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.18485f
C1247 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.251856f
C1248 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.18485f
C1249 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.234527f
C1250 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.345142f
C1251 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.167416f
C1252 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.217197f
C1253 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.345142f
C1254 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.346293f
C1255 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.364878f
C1256 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.186001f
C1257 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.217197f
C1258 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.345142f
C1259 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.217197f
C1260 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.186001f
C1261 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.364878f
C1262 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.364878f
C1263 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.730561f
C1264 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.29977f
C1265 VOUT+.t13 GNDA 0.048668f
C1266 VOUT+.t9 GNDA 0.048668f
C1267 VOUT+.n0 GNDA 0.225914f
C1268 VOUT+.t3 GNDA 0.048668f
C1269 VOUT+.t10 GNDA 0.048668f
C1270 VOUT+.n1 GNDA 0.225185f
C1271 VOUT+.n2 GNDA 0.138481f
C1272 VOUT+.t2 GNDA 0.048668f
C1273 VOUT+.t12 GNDA 0.048668f
C1274 VOUT+.n3 GNDA 0.225185f
C1275 VOUT+.n4 GNDA 0.077142f
C1276 VOUT+.t5 GNDA 0.081011f
C1277 VOUT+.n5 GNDA 0.091611f
C1278 VOUT+.t14 GNDA 0.041716f
C1279 VOUT+.t4 GNDA 0.041716f
C1280 VOUT+.n6 GNDA 0.168663f
C1281 VOUT+.t11 GNDA 0.041716f
C1282 VOUT+.t1 GNDA 0.041716f
C1283 VOUT+.n7 GNDA 0.168362f
C1284 VOUT+.n8 GNDA 0.164256f
C1285 VOUT+.t6 GNDA 0.041716f
C1286 VOUT+.t7 GNDA 0.041716f
C1287 VOUT+.n9 GNDA 0.168362f
C1288 VOUT+.n10 GNDA 0.084712f
C1289 VOUT+.t16 GNDA 0.041716f
C1290 VOUT+.t17 GNDA 0.041716f
C1291 VOUT+.n11 GNDA 0.168362f
C1292 VOUT+.n12 GNDA 0.084712f
C1293 VOUT+.t18 GNDA 0.041716f
C1294 VOUT+.t15 GNDA 0.041716f
C1295 VOUT+.n13 GNDA 0.168663f
C1296 VOUT+.n14 GNDA 0.100402f
C1297 VOUT+.t8 GNDA 0.041716f
C1298 VOUT+.t0 GNDA 0.041716f
C1299 VOUT+.n15 GNDA 0.166369f
C1300 VOUT+.n16 GNDA 0.14091f
C1301 VOUT+.t45 GNDA 0.278104f
C1302 VOUT+.t150 GNDA 0.28284f
C1303 VOUT+.t101 GNDA 0.278104f
C1304 VOUT+.n17 GNDA 0.186459f
C1305 VOUT+.n18 GNDA 0.12167f
C1306 VOUT+.t91 GNDA 0.282247f
C1307 VOUT+.t38 GNDA 0.282247f
C1308 VOUT+.t130 GNDA 0.282247f
C1309 VOUT+.t90 GNDA 0.282247f
C1310 VOUT+.t80 GNDA 0.282247f
C1311 VOUT+.t128 GNDA 0.282247f
C1312 VOUT+.t124 GNDA 0.282247f
C1313 VOUT+.t32 GNDA 0.282247f
C1314 VOUT+.t70 GNDA 0.282247f
C1315 VOUT+.t73 GNDA 0.282247f
C1316 VOUT+.t23 GNDA 0.282247f
C1317 VOUT+.t108 GNDA 0.282247f
C1318 VOUT+.t62 GNDA 0.282247f
C1319 VOUT+.t19 GNDA 0.282247f
C1320 VOUT+.t151 GNDA 0.282247f
C1321 VOUT+.t49 GNDA 0.282247f
C1322 VOUT+.t85 GNDA 0.278104f
C1323 VOUT+.n19 GNDA 0.304579f
C1324 VOUT+.t48 GNDA 0.278104f
C1325 VOUT+.n20 GNDA 0.356724f
C1326 VOUT+.t138 GNDA 0.278104f
C1327 VOUT+.n21 GNDA 0.356724f
C1328 VOUT+.t107 GNDA 0.278104f
C1329 VOUT+.n22 GNDA 0.356724f
C1330 VOUT+.t71 GNDA 0.278104f
C1331 VOUT+.n23 GNDA 0.356724f
C1332 VOUT+.t25 GNDA 0.278104f
C1333 VOUT+.n24 GNDA 0.356724f
C1334 VOUT+.t129 GNDA 0.278104f
C1335 VOUT+.n25 GNDA 0.356724f
C1336 VOUT+.t87 GNDA 0.278104f
C1337 VOUT+.n26 GNDA 0.239197f
C1338 VOUT+.t52 GNDA 0.278104f
C1339 VOUT+.n27 GNDA 0.239197f
C1340 VOUT+.t141 GNDA 0.278104f
C1341 VOUT+.t75 GNDA 0.28284f
C1342 VOUT+.t111 GNDA 0.278104f
C1343 VOUT+.n28 GNDA 0.186459f
C1344 VOUT+.n29 GNDA 0.225959f
C1345 VOUT+.t54 GNDA 0.28284f
C1346 VOUT+.t24 GNDA 0.278104f
C1347 VOUT+.n30 GNDA 0.186459f
C1348 VOUT+.t114 GNDA 0.278104f
C1349 VOUT+.t34 GNDA 0.28284f
C1350 VOUT+.t74 GNDA 0.278104f
C1351 VOUT+.n31 GNDA 0.186459f
C1352 VOUT+.n32 GNDA 0.225959f
C1353 VOUT+.t95 GNDA 0.28284f
C1354 VOUT+.t59 GNDA 0.278104f
C1355 VOUT+.n33 GNDA 0.186459f
C1356 VOUT+.t148 GNDA 0.278104f
C1357 VOUT+.t79 GNDA 0.28284f
C1358 VOUT+.t117 GNDA 0.278104f
C1359 VOUT+.n34 GNDA 0.186459f
C1360 VOUT+.n35 GNDA 0.225959f
C1361 VOUT+.t134 GNDA 0.28284f
C1362 VOUT+.t100 GNDA 0.278104f
C1363 VOUT+.n36 GNDA 0.186459f
C1364 VOUT+.t44 GNDA 0.278104f
C1365 VOUT+.t122 GNDA 0.28284f
C1366 VOUT+.t153 GNDA 0.278104f
C1367 VOUT+.n37 GNDA 0.186459f
C1368 VOUT+.n38 GNDA 0.225959f
C1369 VOUT+.t102 GNDA 0.28284f
C1370 VOUT+.t66 GNDA 0.278104f
C1371 VOUT+.n39 GNDA 0.186459f
C1372 VOUT+.t154 GNDA 0.278104f
C1373 VOUT+.t82 GNDA 0.28284f
C1374 VOUT+.t123 GNDA 0.278104f
C1375 VOUT+.n40 GNDA 0.186459f
C1376 VOUT+.n41 GNDA 0.225959f
C1377 VOUT+.t137 GNDA 0.28284f
C1378 VOUT+.t106 GNDA 0.278104f
C1379 VOUT+.n42 GNDA 0.186459f
C1380 VOUT+.t51 GNDA 0.278104f
C1381 VOUT+.t126 GNDA 0.28284f
C1382 VOUT+.t22 GNDA 0.278104f
C1383 VOUT+.n43 GNDA 0.186459f
C1384 VOUT+.n44 GNDA 0.225959f
C1385 VOUT+.t132 GNDA 0.278104f
C1386 VOUT+.t56 GNDA 0.28284f
C1387 VOUT+.t96 GNDA 0.278104f
C1388 VOUT+.n45 GNDA 0.186459f
C1389 VOUT+.n46 GNDA 0.12167f
C1390 VOUT+.t116 GNDA 0.282247f
C1391 VOUT+.t105 GNDA 0.28284f
C1392 VOUT+.t69 GNDA 0.278104f
C1393 VOUT+.n47 GNDA 0.182114f
C1394 VOUT+.t147 GNDA 0.282247f
C1395 VOUT+.t29 GNDA 0.28284f
C1396 VOUT+.t139 GNDA 0.278104f
C1397 VOUT+.n48 GNDA 0.186459f
C1398 VOUT+.t109 GNDA 0.278104f
C1399 VOUT+.n49 GNDA 0.117325f
C1400 VOUT+.t43 GNDA 0.282247f
C1401 VOUT+.t60 GNDA 0.28284f
C1402 VOUT+.t37 GNDA 0.278104f
C1403 VOUT+.n50 GNDA 0.186459f
C1404 VOUT+.t144 GNDA 0.278104f
C1405 VOUT+.n51 GNDA 0.117325f
C1406 VOUT+.t83 GNDA 0.282247f
C1407 VOUT+.t115 GNDA 0.28284f
C1408 VOUT+.t21 GNDA 0.278104f
C1409 VOUT+.n52 GNDA 0.186459f
C1410 VOUT+.t125 GNDA 0.278104f
C1411 VOUT+.n53 GNDA 0.117325f
C1412 VOUT+.t63 GNDA 0.282247f
C1413 VOUT+.t26 GNDA 0.282247f
C1414 VOUT+.t103 GNDA 0.282247f
C1415 VOUT+.t57 GNDA 0.28248f
C1416 VOUT+.t135 GNDA 0.282247f
C1417 VOUT+.t33 GNDA 0.28248f
C1418 VOUT+.t120 GNDA 0.282247f
C1419 VOUT+.t77 GNDA 0.28248f
C1420 VOUT+.t155 GNDA 0.282247f
C1421 VOUT+.t119 GNDA 0.278104f
C1422 VOUT+.n54 GNDA 0.307823f
C1423 VOUT+.t78 GNDA 0.278104f
C1424 VOUT+.n55 GNDA 0.359967f
C1425 VOUT+.t97 GNDA 0.278104f
C1426 VOUT+.n56 GNDA 0.359967f
C1427 VOUT+.t61 GNDA 0.278104f
C1428 VOUT+.n57 GNDA 0.356724f
C1429 VOUT+.t27 GNDA 0.278104f
C1430 VOUT+.n58 GNDA 0.295687f
C1431 VOUT+.t41 GNDA 0.278104f
C1432 VOUT+.n59 GNDA 0.295687f
C1433 VOUT+.t145 GNDA 0.278104f
C1434 VOUT+.n60 GNDA 0.295687f
C1435 VOUT+.t113 GNDA 0.278104f
C1436 VOUT+.n61 GNDA 0.295687f
C1437 VOUT+.t72 GNDA 0.278104f
C1438 VOUT+.n62 GNDA 0.239197f
C1439 VOUT+.t92 GNDA 0.278104f
C1440 VOUT+.t20 GNDA 0.28284f
C1441 VOUT+.t55 GNDA 0.278104f
C1442 VOUT+.n63 GNDA 0.186459f
C1443 VOUT+.n64 GNDA 0.225959f
C1444 VOUT+.t31 GNDA 0.28284f
C1445 VOUT+.t50 GNDA 0.278104f
C1446 VOUT+.t121 GNDA 0.28284f
C1447 VOUT+.t156 GNDA 0.278104f
C1448 VOUT+.n65 GNDA 0.186459f
C1449 VOUT+.n66 GNDA 0.290748f
C1450 VOUT+.t67 GNDA 0.28284f
C1451 VOUT+.t86 GNDA 0.278104f
C1452 VOUT+.t152 GNDA 0.28284f
C1453 VOUT+.t47 GNDA 0.278104f
C1454 VOUT+.n67 GNDA 0.186459f
C1455 VOUT+.n68 GNDA 0.290748f
C1456 VOUT+.t131 GNDA 0.28284f
C1457 VOUT+.t94 GNDA 0.278104f
C1458 VOUT+.n69 GNDA 0.186459f
C1459 VOUT+.t39 GNDA 0.278104f
C1460 VOUT+.t118 GNDA 0.28284f
C1461 VOUT+.t146 GNDA 0.278104f
C1462 VOUT+.n70 GNDA 0.186459f
C1463 VOUT+.n71 GNDA 0.225959f
C1464 VOUT+.t89 GNDA 0.28284f
C1465 VOUT+.t53 GNDA 0.278104f
C1466 VOUT+.n72 GNDA 0.186459f
C1467 VOUT+.t142 GNDA 0.278104f
C1468 VOUT+.t76 GNDA 0.28284f
C1469 VOUT+.t112 GNDA 0.278104f
C1470 VOUT+.n73 GNDA 0.186459f
C1471 VOUT+.n74 GNDA 0.225959f
C1472 VOUT+.t127 GNDA 0.28284f
C1473 VOUT+.t88 GNDA 0.278104f
C1474 VOUT+.n75 GNDA 0.186459f
C1475 VOUT+.t35 GNDA 0.278104f
C1476 VOUT+.t110 GNDA 0.28284f
C1477 VOUT+.t140 GNDA 0.278104f
C1478 VOUT+.n76 GNDA 0.186459f
C1479 VOUT+.n77 GNDA 0.225959f
C1480 VOUT+.t84 GNDA 0.28284f
C1481 VOUT+.t46 GNDA 0.278104f
C1482 VOUT+.n78 GNDA 0.186459f
C1483 VOUT+.t136 GNDA 0.278104f
C1484 VOUT+.t68 GNDA 0.28284f
C1485 VOUT+.t104 GNDA 0.278104f
C1486 VOUT+.n79 GNDA 0.186459f
C1487 VOUT+.n80 GNDA 0.225959f
C1488 VOUT+.t42 GNDA 0.28284f
C1489 VOUT+.t149 GNDA 0.278104f
C1490 VOUT+.n81 GNDA 0.186459f
C1491 VOUT+.t99 GNDA 0.278104f
C1492 VOUT+.t30 GNDA 0.28284f
C1493 VOUT+.t65 GNDA 0.278104f
C1494 VOUT+.n82 GNDA 0.186459f
C1495 VOUT+.n83 GNDA 0.225959f
C1496 VOUT+.t81 GNDA 0.28284f
C1497 VOUT+.t40 GNDA 0.278104f
C1498 VOUT+.n84 GNDA 0.186459f
C1499 VOUT+.t133 GNDA 0.278104f
C1500 VOUT+.t64 GNDA 0.28284f
C1501 VOUT+.t98 GNDA 0.278104f
C1502 VOUT+.n85 GNDA 0.186459f
C1503 VOUT+.n86 GNDA 0.225959f
C1504 VOUT+.t28 GNDA 0.28284f
C1505 VOUT+.t58 GNDA 0.278104f
C1506 VOUT+.n87 GNDA 0.186459f
C1507 VOUT+.t93 GNDA 0.278104f
C1508 VOUT+.n88 GNDA 0.225959f
C1509 VOUT+.t143 GNDA 0.278104f
C1510 VOUT+.n89 GNDA 0.12167f
C1511 VOUT+.t36 GNDA 0.278104f
C1512 VOUT+.n90 GNDA 0.177423f
C1513 VOUT+.n91 GNDA 0.210673f
C1514 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.013493f
C1515 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.013493f
C1516 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.049393f
C1517 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.013493f
C1518 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.013493f
C1519 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.048979f
C1520 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.179573f
C1521 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.013493f
C1522 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.013493f
C1523 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.048979f
C1524 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.093142f
C1525 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.013493f
C1526 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.013493f
C1527 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.048979f
C1528 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.093142f
C1529 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.013493f
C1530 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.013493f
C1531 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.048979f
C1532 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.093142f
C1533 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.013493f
C1534 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.013493f
C1535 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.048979f
C1536 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.112031f
C1537 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.031482f
C1538 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.031482f
C1539 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.110567f
C1540 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.031482f
C1541 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.031482f
C1542 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.110188f
C1543 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.205608f
C1544 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.031482f
C1545 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.031482f
C1546 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.110188f
C1547 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.106591f
C1548 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.031482f
C1549 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.031482f
C1550 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.110188f
C1551 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.106591f
C1552 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.031482f
C1553 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.031482f
C1554 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.110188f
C1555 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.125547f
C1556 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.031482f
C1557 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.031482f
C1558 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.107979f
C1559 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.184593f
C1560 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.018889f
C1561 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.018889f
C1562 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.018889f
C1563 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.018889f
C1564 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.018889f
C1565 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.022937f
C1566 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.022937f
C1567 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.014842f
C1568 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.014842f
C1569 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.014842f
C1570 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.013091f
C1571 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.018889f
C1572 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.018889f
C1573 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.018889f
C1574 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.022937f
C1575 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.022937f
C1576 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.014842f
C1577 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.013091f
C1578 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.013602f
C1579 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.029009f
C1580 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.029009f
C1581 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.029009f
C1582 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.029009f
C1583 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.029009f
C1584 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.032978f
C1585 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.029762f
C1586 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.018215f
C1587 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.018215f
C1588 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.018215f
C1589 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.016464f
C1590 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.029009f
C1591 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.029009f
C1592 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.029009f
C1593 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.032978f
C1594 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.029762f
C1595 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.018215f
C1596 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.016464f
C1597 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.013602f
C1598 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.121373f
C1599 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.290786f
C1600 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.075108f
C1601 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.059367f
C1602 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.059367f
C1603 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.059367f
C1604 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.059367f
C1605 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.06323f
C1606 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.050107f
C1607 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.028334f
C1608 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.028334f
C1609 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.02659f
C1610 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.059367f
C1611 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.059367f
C1612 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.059367f
C1613 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.059367f
C1614 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.06323f
C1615 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.050107f
C1616 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.028334f
C1617 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.028334f
C1618 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.02659f
C1619 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.016175f
C1620 two_stage_opamp_dummy_magic_0.X.n52 GNDA 0.47889f
C1621 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.437337f
C1622 two_stage_opamp_dummy_magic_0.Vb1.n0 GNDA 0.020805f
C1623 two_stage_opamp_dummy_magic_0.Vb1.n1 GNDA 0.020666f
C1624 two_stage_opamp_dummy_magic_0.Vb1.n2 GNDA 0.226929f
C1625 two_stage_opamp_dummy_magic_0.Vb1.t1 GNDA 0.236522f
C1626 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA 0.038084f
C1627 two_stage_opamp_dummy_magic_0.Vb1.n3 GNDA 0.347531f
C1628 two_stage_opamp_dummy_magic_0.Vb1.t24 GNDA 0.012761f
C1629 two_stage_opamp_dummy_magic_0.Vb1.t14 GNDA 0.012761f
C1630 two_stage_opamp_dummy_magic_0.Vb1.t23 GNDA 0.012761f
C1631 two_stage_opamp_dummy_magic_0.Vb1.t6 GNDA 0.012761f
C1632 two_stage_opamp_dummy_magic_0.Vb1.t16 GNDA 0.016552f
C1633 two_stage_opamp_dummy_magic_0.Vb1.n4 GNDA 0.017997f
C1634 two_stage_opamp_dummy_magic_0.Vb1.n5 GNDA 0.012139f
C1635 two_stage_opamp_dummy_magic_0.Vb1.n6 GNDA 0.012139f
C1636 two_stage_opamp_dummy_magic_0.Vb1.n7 GNDA 0.010523f
C1637 two_stage_opamp_dummy_magic_0.Vb1.t15 GNDA 0.012761f
C1638 two_stage_opamp_dummy_magic_0.Vb1.t19 GNDA 0.012761f
C1639 two_stage_opamp_dummy_magic_0.Vb1.t10 GNDA 0.012761f
C1640 two_stage_opamp_dummy_magic_0.Vb1.t21 GNDA 0.012761f
C1641 two_stage_opamp_dummy_magic_0.Vb1.t12 GNDA 0.016552f
C1642 two_stage_opamp_dummy_magic_0.Vb1.n8 GNDA 0.017997f
C1643 two_stage_opamp_dummy_magic_0.Vb1.n9 GNDA 0.012139f
C1644 two_stage_opamp_dummy_magic_0.Vb1.n10 GNDA 0.012139f
C1645 two_stage_opamp_dummy_magic_0.Vb1.n11 GNDA 0.010523f
C1646 two_stage_opamp_dummy_magic_0.Vb1.n12 GNDA 0.017235f
C1647 two_stage_opamp_dummy_magic_0.Vb1.t25 GNDA 0.012761f
C1648 two_stage_opamp_dummy_magic_0.Vb1.t9 GNDA 0.012761f
C1649 two_stage_opamp_dummy_magic_0.Vb1.t18 GNDA 0.012761f
C1650 two_stage_opamp_dummy_magic_0.Vb1.t7 GNDA 0.012761f
C1651 two_stage_opamp_dummy_magic_0.Vb1.t17 GNDA 0.016552f
C1652 two_stage_opamp_dummy_magic_0.Vb1.n13 GNDA 0.017997f
C1653 two_stage_opamp_dummy_magic_0.Vb1.n14 GNDA 0.012139f
C1654 two_stage_opamp_dummy_magic_0.Vb1.n15 GNDA 0.012139f
C1655 two_stage_opamp_dummy_magic_0.Vb1.n16 GNDA 0.010523f
C1656 two_stage_opamp_dummy_magic_0.Vb1.t8 GNDA 0.012761f
C1657 two_stage_opamp_dummy_magic_0.Vb1.t20 GNDA 0.012761f
C1658 two_stage_opamp_dummy_magic_0.Vb1.t11 GNDA 0.012761f
C1659 two_stage_opamp_dummy_magic_0.Vb1.t22 GNDA 0.012761f
C1660 two_stage_opamp_dummy_magic_0.Vb1.t13 GNDA 0.016552f
C1661 two_stage_opamp_dummy_magic_0.Vb1.n17 GNDA 0.017997f
C1662 two_stage_opamp_dummy_magic_0.Vb1.n18 GNDA 0.012139f
C1663 two_stage_opamp_dummy_magic_0.Vb1.n19 GNDA 0.012139f
C1664 two_stage_opamp_dummy_magic_0.Vb1.n20 GNDA 0.010523f
C1665 two_stage_opamp_dummy_magic_0.Vb1.n21 GNDA 0.013046f
C1666 two_stage_opamp_dummy_magic_0.Vb1.n22 GNDA 0.280421f
C1667 two_stage_opamp_dummy_magic_0.Vb1.n23 GNDA 0.723357f
C1668 bgr_0.VB1_CUR_BIAS GNDA 0.46063f
C1669 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 GNDA 0.011375f
C1670 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 GNDA 0.011375f
C1671 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA 0.011375f
C1672 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 GNDA 0.032925f
C1673 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 GNDA 0.011375f
C1674 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA 0.011375f
C1675 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 GNDA 0.025519f
C1676 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA 0.011375f
C1677 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 GNDA 0.011375f
C1678 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 GNDA 0.027057f
C1679 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA 0.011375f
C1680 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA 0.011375f
C1681 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 GNDA 0.026605f
C1682 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 GNDA 0.557444f
C1683 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 GNDA 0.223671f
C1684 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 GNDA 0.255693f
C1685 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 GNDA 0.27819f
C1686 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 GNDA 0.020334f
C1687 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 GNDA 0.031709f
C1688 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 GNDA 0.024742f
C1689 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 GNDA 0.022056f
C1690 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 GNDA 0.011375f
C1691 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 GNDA 0.011375f
C1692 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 GNDA 0.026858f
C1693 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 GNDA 0.094877f
C1694 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 GNDA 0.032671f
C1695 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 GNDA 0.022056f
C1696 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 GNDA 0.024742f
C1697 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 GNDA 0.024742f
C1698 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 GNDA 0.022056f
C1699 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA 0.020334f
C1700 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 GNDA 0.029024f
C1701 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 GNDA 0.032671f
C1702 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 GNDA 0.105585f
C1703 two_stage_opamp_dummy_magic_0.err_amp_mir.n21 GNDA 0.026858f
C1704 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA 0.011375f
C1705 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.346251f
C1706 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.347506f
C1707 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.346251f
C1708 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.348966f
C1709 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.379551f
C1710 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.346251f
C1711 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.347506f
C1712 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.328924f
C1713 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.346251f
C1714 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.347506f
C1715 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.328924f
C1716 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.346251f
C1717 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.347506f
C1718 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.346251f
C1719 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.347506f
C1720 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.346251f
C1721 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.347506f
C1722 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.346251f
C1723 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.347506f
C1724 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.346251f
C1725 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.347506f
C1726 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.346251f
C1727 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.347506f
C1728 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.346251f
C1729 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.347506f
C1730 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.346251f
C1731 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.347506f
C1732 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.346251f
C1733 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.347506f
C1734 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.346251f
C1735 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.347506f
C1736 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.346251f
C1737 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.347506f
C1738 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.346251f
C1739 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.347506f
C1740 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.346251f
C1741 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.347506f
C1742 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.346251f
C1743 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.347506f
C1744 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.346251f
C1745 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.347506f
C1746 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.346251f
C1747 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.347506f
C1748 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.346251f
C1749 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.347506f
C1750 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.346251f
C1751 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.347506f
C1752 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.346251f
C1753 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.347506f
C1754 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.346251f
C1755 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.347506f
C1756 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.346251f
C1757 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.347506f
C1758 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.346251f
C1759 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.347506f
C1760 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.346251f
C1761 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.347506f
C1762 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.346251f
C1763 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.347506f
C1764 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.346251f
C1765 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.347506f
C1766 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.3451f
C1767 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.346251f
C1768 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.185978f
C1769 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.198589f
C1770 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.3451f
C1771 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.346251f
C1772 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.185978f
C1773 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.217171f
C1774 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.3451f
C1775 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.346251f
C1776 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.185978f
C1777 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.217171f
C1778 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.3451f
C1779 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.346251f
C1780 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.185978f
C1781 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.217171f
C1782 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.3451f
C1783 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.346251f
C1784 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185978f
C1785 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.217171f
C1786 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.3451f
C1787 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.346251f
C1788 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.185978f
C1789 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.217171f
C1790 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.3451f
C1791 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.346251f
C1792 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.185978f
C1793 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.217171f
C1794 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.346251f
C1795 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.185978f
C1796 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.197438f
C1797 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.346251f
C1798 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.185978f
C1799 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.197438f
C1800 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.346251f
C1801 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.347506f
C1802 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.167396f
C1803 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.215916f
C1804 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.184828f
C1805 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.234498f
C1806 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.184828f
C1807 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.251826f
C1808 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.184828f
C1809 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.251826f
C1810 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.184828f
C1811 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.251826f
C1812 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.184828f
C1813 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.251826f
C1814 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.184828f
C1815 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.251826f
C1816 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.184828f
C1817 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.251826f
C1818 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.184828f
C1819 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.251826f
C1820 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.184828f
C1821 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.251826f
C1822 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.184828f
C1823 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.251826f
C1824 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.184828f
C1825 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.251826f
C1826 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.184828f
C1827 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.251826f
C1828 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.184828f
C1829 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.251826f
C1830 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.184828f
C1831 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.251826f
C1832 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.184828f
C1833 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.251826f
C1834 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.184828f
C1835 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.234498f
C1836 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.3451f
C1837 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.167396f
C1838 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.217171f
C1839 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.3451f
C1840 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.346251f
C1841 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.364834f
C1842 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.185978f
C1843 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.217171f
C1844 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.3451f
C1845 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.346251f
C1846 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.185978f
C1847 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.198589f
C1848 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.3451f
C1849 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.346251f
C1850 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.185978f
C1851 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.217171f
C1852 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.3451f
C1853 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.346251f
C1854 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.185978f
C1855 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.217171f
C1856 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.3451f
C1857 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.346251f
C1858 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.185978f
C1859 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.217171f
C1860 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.3451f
C1861 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.346251f
C1862 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.364834f
C1863 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.364834f
C1864 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.185978f
C1865 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.217171f
C1866 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.3451f
C1867 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.346251f
C1868 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.364834f
C1869 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.364834f
C1870 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.185978f
C1871 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.217171f
C1872 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.3451f
C1873 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.217171f
C1874 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.185978f
C1875 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.364834f
C1876 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.364834f
C1877 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.430822f
C1878 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.292647f
C1879 VOUT-.t13 GNDA 0.041786f
C1880 VOUT-.t9 GNDA 0.041786f
C1881 VOUT-.n0 GNDA 0.16895f
C1882 VOUT-.t2 GNDA 0.041786f
C1883 VOUT-.t14 GNDA 0.041786f
C1884 VOUT-.n1 GNDA 0.168949f
C1885 VOUT-.t0 GNDA 0.041786f
C1886 VOUT-.t15 GNDA 0.041786f
C1887 VOUT-.n2 GNDA 0.168648f
C1888 VOUT-.n3 GNDA 0.164536f
C1889 VOUT-.t5 GNDA 0.041786f
C1890 VOUT-.t16 GNDA 0.041786f
C1891 VOUT-.n4 GNDA 0.168648f
C1892 VOUT-.n5 GNDA 0.084856f
C1893 VOUT-.t6 GNDA 0.041786f
C1894 VOUT-.t7 GNDA 0.041786f
C1895 VOUT-.n6 GNDA 0.168648f
C1896 VOUT-.n7 GNDA 0.084856f
C1897 VOUT-.n8 GNDA 0.100572f
C1898 VOUT-.t1 GNDA 0.041786f
C1899 VOUT-.t8 GNDA 0.041786f
C1900 VOUT-.n9 GNDA 0.166651f
C1901 VOUT-.n10 GNDA 0.141149f
C1902 VOUT-.t26 GNDA 0.283321f
C1903 VOUT-.t119 GNDA 0.278576f
C1904 VOUT-.n11 GNDA 0.186776f
C1905 VOUT-.t33 GNDA 0.278576f
C1906 VOUT-.n12 GNDA 0.121877f
C1907 VOUT-.t36 GNDA 0.283321f
C1908 VOUT-.t122 GNDA 0.278576f
C1909 VOUT-.n13 GNDA 0.186776f
C1910 VOUT-.t90 GNDA 0.278576f
C1911 VOUT-.t82 GNDA 0.282727f
C1912 VOUT-.t42 GNDA 0.282727f
C1913 VOUT-.t92 GNDA 0.282727f
C1914 VOUT-.t74 GNDA 0.282727f
C1915 VOUT-.t141 GNDA 0.282727f
C1916 VOUT-.t38 GNDA 0.282727f
C1917 VOUT-.t105 GNDA 0.282727f
C1918 VOUT-.t126 GNDA 0.282727f
C1919 VOUT-.t154 GNDA 0.282727f
C1920 VOUT-.t95 GNDA 0.282727f
C1921 VOUT-.t65 GNDA 0.282727f
C1922 VOUT-.t62 GNDA 0.282727f
C1923 VOUT-.t114 GNDA 0.282727f
C1924 VOUT-.t24 GNDA 0.282727f
C1925 VOUT-.t71 GNDA 0.282727f
C1926 VOUT-.t113 GNDA 0.282727f
C1927 VOUT-.t148 GNDA 0.278576f
C1928 VOUT-.n14 GNDA 0.305096f
C1929 VOUT-.t60 GNDA 0.278576f
C1930 VOUT-.n15 GNDA 0.357329f
C1931 VOUT-.t93 GNDA 0.278576f
C1932 VOUT-.n16 GNDA 0.357329f
C1933 VOUT-.t127 GNDA 0.278576f
C1934 VOUT-.n17 GNDA 0.357329f
C1935 VOUT-.t25 GNDA 0.278576f
C1936 VOUT-.n18 GNDA 0.357329f
C1937 VOUT-.t72 GNDA 0.278576f
C1938 VOUT-.n19 GNDA 0.357329f
C1939 VOUT-.t110 GNDA 0.278576f
C1940 VOUT-.n20 GNDA 0.357329f
C1941 VOUT-.t142 GNDA 0.278576f
C1942 VOUT-.n21 GNDA 0.239603f
C1943 VOUT-.t56 GNDA 0.278576f
C1944 VOUT-.n22 GNDA 0.239603f
C1945 VOUT-.n23 GNDA 0.226343f
C1946 VOUT-.t140 GNDA 0.283321f
C1947 VOUT-.t89 GNDA 0.278576f
C1948 VOUT-.n24 GNDA 0.186776f
C1949 VOUT-.t59 GNDA 0.278576f
C1950 VOUT-.t111 GNDA 0.283321f
C1951 VOUT-.t21 GNDA 0.278576f
C1952 VOUT-.n25 GNDA 0.186776f
C1953 VOUT-.n26 GNDA 0.226343f
C1954 VOUT-.t41 GNDA 0.283321f
C1955 VOUT-.t129 GNDA 0.278576f
C1956 VOUT-.n27 GNDA 0.186776f
C1957 VOUT-.t98 GNDA 0.278576f
C1958 VOUT-.t151 GNDA 0.283321f
C1959 VOUT-.t63 GNDA 0.278576f
C1960 VOUT-.n28 GNDA 0.186776f
C1961 VOUT-.n29 GNDA 0.226343f
C1962 VOUT-.t80 GNDA 0.283321f
C1963 VOUT-.t30 GNDA 0.278576f
C1964 VOUT-.n30 GNDA 0.186776f
C1965 VOUT-.t134 GNDA 0.278576f
C1966 VOUT-.t51 GNDA 0.283321f
C1967 VOUT-.t103 GNDA 0.278576f
C1968 VOUT-.n31 GNDA 0.186776f
C1969 VOUT-.n32 GNDA 0.226343f
C1970 VOUT-.t49 GNDA 0.283321f
C1971 VOUT-.t135 GNDA 0.278576f
C1972 VOUT-.n33 GNDA 0.186776f
C1973 VOUT-.t102 GNDA 0.278576f
C1974 VOUT-.t19 GNDA 0.283321f
C1975 VOUT-.t67 GNDA 0.278576f
C1976 VOUT-.n34 GNDA 0.186776f
C1977 VOUT-.n35 GNDA 0.226343f
C1978 VOUT-.t85 GNDA 0.283321f
C1979 VOUT-.t34 GNDA 0.278576f
C1980 VOUT-.n36 GNDA 0.186776f
C1981 VOUT-.t139 GNDA 0.278576f
C1982 VOUT-.t55 GNDA 0.283321f
C1983 VOUT-.t106 GNDA 0.278576f
C1984 VOUT-.n37 GNDA 0.186776f
C1985 VOUT-.n38 GNDA 0.226343f
C1986 VOUT-.t68 GNDA 0.283321f
C1987 VOUT-.t86 GNDA 0.278576f
C1988 VOUT-.n39 GNDA 0.186776f
C1989 VOUT-.t54 GNDA 0.278576f
C1990 VOUT-.n40 GNDA 0.121877f
C1991 VOUT-.t29 GNDA 0.283321f
C1992 VOUT-.t52 GNDA 0.278576f
C1993 VOUT-.n41 GNDA 0.186776f
C1994 VOUT-.t155 GNDA 0.278576f
C1995 VOUT-.t156 GNDA 0.282727f
C1996 VOUT-.t132 GNDA 0.283321f
C1997 VOUT-.t99 GNDA 0.278576f
C1998 VOUT-.n42 GNDA 0.182423f
C1999 VOUT-.t35 GNDA 0.282727f
C2000 VOUT-.t150 GNDA 0.283321f
C2001 VOUT-.t94 GNDA 0.278576f
C2002 VOUT-.n43 GNDA 0.186776f
C2003 VOUT-.t61 GNDA 0.278576f
C2004 VOUT-.n44 GNDA 0.117524f
C2005 VOUT-.t137 GNDA 0.282727f
C2006 VOUT-.t115 GNDA 0.283321f
C2007 VOUT-.t58 GNDA 0.278576f
C2008 VOUT-.n45 GNDA 0.186776f
C2009 VOUT-.t22 GNDA 0.278576f
C2010 VOUT-.n46 GNDA 0.117524f
C2011 VOUT-.t104 GNDA 0.282727f
C2012 VOUT-.t66 GNDA 0.283321f
C2013 VOUT-.t77 GNDA 0.278576f
C2014 VOUT-.n47 GNDA 0.186776f
C2015 VOUT-.t43 GNDA 0.278576f
C2016 VOUT-.n48 GNDA 0.117524f
C2017 VOUT-.t120 GNDA 0.282727f
C2018 VOUT-.t144 GNDA 0.282727f
C2019 VOUT-.t83 GNDA 0.282727f
C2020 VOUT-.t107 GNDA 0.28296f
C2021 VOUT-.t50 GNDA 0.282727f
C2022 VOUT-.t69 GNDA 0.28296f
C2023 VOUT-.t149 GNDA 0.282727f
C2024 VOUT-.t91 GNDA 0.28296f
C2025 VOUT-.t31 GNDA 0.282727f
C2026 VOUT-.t130 GNDA 0.278576f
C2027 VOUT-.n49 GNDA 0.308345f
C2028 VOUT-.t108 GNDA 0.278576f
C2029 VOUT-.n50 GNDA 0.360578f
C2030 VOUT-.t146 GNDA 0.278576f
C2031 VOUT-.n51 GNDA 0.360578f
C2032 VOUT-.t45 GNDA 0.278576f
C2033 VOUT-.n52 GNDA 0.357329f
C2034 VOUT-.t81 GNDA 0.278576f
C2035 VOUT-.n53 GNDA 0.296189f
C2036 VOUT-.t64 GNDA 0.278576f
C2037 VOUT-.n54 GNDA 0.296189f
C2038 VOUT-.t100 GNDA 0.278576f
C2039 VOUT-.n55 GNDA 0.296189f
C2040 VOUT-.t136 GNDA 0.278576f
C2041 VOUT-.n56 GNDA 0.296189f
C2042 VOUT-.t116 GNDA 0.278576f
C2043 VOUT-.n57 GNDA 0.239603f
C2044 VOUT-.n58 GNDA 0.226343f
C2045 VOUT-.t125 GNDA 0.283321f
C2046 VOUT-.t152 GNDA 0.278576f
C2047 VOUT-.n59 GNDA 0.186776f
C2048 VOUT-.t112 GNDA 0.278576f
C2049 VOUT-.t73 GNDA 0.283321f
C2050 VOUT-.n60 GNDA 0.291242f
C2051 VOUT-.t23 GNDA 0.283321f
C2052 VOUT-.t47 GNDA 0.278576f
C2053 VOUT-.n61 GNDA 0.186776f
C2054 VOUT-.t147 GNDA 0.278576f
C2055 VOUT-.t109 GNDA 0.283321f
C2056 VOUT-.n62 GNDA 0.291242f
C2057 VOUT-.t76 GNDA 0.283321f
C2058 VOUT-.t27 GNDA 0.278576f
C2059 VOUT-.n63 GNDA 0.186776f
C2060 VOUT-.t128 GNDA 0.278576f
C2061 VOUT-.t44 GNDA 0.283321f
C2062 VOUT-.t97 GNDA 0.278576f
C2063 VOUT-.n64 GNDA 0.186776f
C2064 VOUT-.n65 GNDA 0.226343f
C2065 VOUT-.t37 GNDA 0.283321f
C2066 VOUT-.t123 GNDA 0.278576f
C2067 VOUT-.n66 GNDA 0.186776f
C2068 VOUT-.t88 GNDA 0.278576f
C2069 VOUT-.t143 GNDA 0.283321f
C2070 VOUT-.t57 GNDA 0.278576f
C2071 VOUT-.n67 GNDA 0.186776f
C2072 VOUT-.n68 GNDA 0.226343f
C2073 VOUT-.t70 GNDA 0.283321f
C2074 VOUT-.t20 GNDA 0.278576f
C2075 VOUT-.n69 GNDA 0.186776f
C2076 VOUT-.t121 GNDA 0.278576f
C2077 VOUT-.t39 GNDA 0.283321f
C2078 VOUT-.t87 GNDA 0.278576f
C2079 VOUT-.n70 GNDA 0.186776f
C2080 VOUT-.n71 GNDA 0.226343f
C2081 VOUT-.t32 GNDA 0.283321f
C2082 VOUT-.t118 GNDA 0.278576f
C2083 VOUT-.n72 GNDA 0.186776f
C2084 VOUT-.t84 GNDA 0.278576f
C2085 VOUT-.t138 GNDA 0.283321f
C2086 VOUT-.t53 GNDA 0.278576f
C2087 VOUT-.n73 GNDA 0.186776f
C2088 VOUT-.n74 GNDA 0.226343f
C2089 VOUT-.t131 GNDA 0.283321f
C2090 VOUT-.t79 GNDA 0.278576f
C2091 VOUT-.n75 GNDA 0.186776f
C2092 VOUT-.t48 GNDA 0.278576f
C2093 VOUT-.t101 GNDA 0.283321f
C2094 VOUT-.t153 GNDA 0.278576f
C2095 VOUT-.n76 GNDA 0.186776f
C2096 VOUT-.n77 GNDA 0.226343f
C2097 VOUT-.t28 GNDA 0.283321f
C2098 VOUT-.t117 GNDA 0.278576f
C2099 VOUT-.n78 GNDA 0.186776f
C2100 VOUT-.t78 GNDA 0.278576f
C2101 VOUT-.t133 GNDA 0.283321f
C2102 VOUT-.t46 GNDA 0.278576f
C2103 VOUT-.n79 GNDA 0.186776f
C2104 VOUT-.n80 GNDA 0.226343f
C2105 VOUT-.t124 GNDA 0.283321f
C2106 VOUT-.t75 GNDA 0.278576f
C2107 VOUT-.n81 GNDA 0.186776f
C2108 VOUT-.t40 GNDA 0.278576f
C2109 VOUT-.n82 GNDA 0.226343f
C2110 VOUT-.t145 GNDA 0.278576f
C2111 VOUT-.n83 GNDA 0.121877f
C2112 VOUT-.t96 GNDA 0.278576f
C2113 VOUT-.n84 GNDA 0.177725f
C2114 VOUT-.n85 GNDA 0.212227f
C2115 VOUT-.t4 GNDA 0.048751f
C2116 VOUT-.t11 GNDA 0.048751f
C2117 VOUT-.n86 GNDA 0.226297f
C2118 VOUT-.t10 GNDA 0.048751f
C2119 VOUT-.t18 GNDA 0.048751f
C2120 VOUT-.n87 GNDA 0.225568f
C2121 VOUT-.n88 GNDA 0.138716f
C2122 VOUT-.t12 GNDA 0.048751f
C2123 VOUT-.t3 GNDA 0.048751f
C2124 VOUT-.n89 GNDA 0.225568f
C2125 VOUT-.n90 GNDA 0.077273f
C2126 VOUT-.t17 GNDA 0.081149f
C2127 VOUT-.n91 GNDA 0.089317f
C2128 bgr_0.V_TOP.t24 GNDA 0.095448f
C2129 bgr_0.V_TOP.t33 GNDA 0.095448f
C2130 bgr_0.V_TOP.t39 GNDA 0.095448f
C2131 bgr_0.V_TOP.t16 GNDA 0.095448f
C2132 bgr_0.V_TOP.t15 GNDA 0.095448f
C2133 bgr_0.V_TOP.t28 GNDA 0.095448f
C2134 bgr_0.V_TOP.t38 GNDA 0.095448f
C2135 bgr_0.V_TOP.t14 GNDA 0.095448f
C2136 bgr_0.V_TOP.t27 GNDA 0.095448f
C2137 bgr_0.V_TOP.t26 GNDA 0.095448f
C2138 bgr_0.V_TOP.t37 GNDA 0.095448f
C2139 bgr_0.V_TOP.t46 GNDA 0.095448f
C2140 bgr_0.V_TOP.t18 GNDA 0.095448f
C2141 bgr_0.V_TOP.t30 GNDA 0.095448f
C2142 bgr_0.V_TOP.t29 GNDA 0.124774f
C2143 bgr_0.V_TOP.n0 GNDA 0.069758f
C2144 bgr_0.V_TOP.n1 GNDA 0.050905f
C2145 bgr_0.V_TOP.n2 GNDA 0.050905f
C2146 bgr_0.V_TOP.n3 GNDA 0.050905f
C2147 bgr_0.V_TOP.n4 GNDA 0.050905f
C2148 bgr_0.V_TOP.n5 GNDA 0.04747f
C2149 bgr_0.V_TOP.t8 GNDA 0.122745f
C2150 bgr_0.V_TOP.t40 GNDA 0.36361f
C2151 bgr_0.V_TOP.t31 GNDA 0.369803f
C2152 bgr_0.V_TOP.t35 GNDA 0.36361f
C2153 bgr_0.V_TOP.n6 GNDA 0.243789f
C2154 bgr_0.V_TOP.t32 GNDA 0.36361f
C2155 bgr_0.V_TOP.t22 GNDA 0.369803f
C2156 bgr_0.V_TOP.n7 GNDA 0.311966f
C2157 bgr_0.V_TOP.t20 GNDA 0.369803f
C2158 bgr_0.V_TOP.t25 GNDA 0.36361f
C2159 bgr_0.V_TOP.n8 GNDA 0.243789f
C2160 bgr_0.V_TOP.t21 GNDA 0.36361f
C2161 bgr_0.V_TOP.t45 GNDA 0.369803f
C2162 bgr_0.V_TOP.n9 GNDA 0.380142f
C2163 bgr_0.V_TOP.t42 GNDA 0.369803f
C2164 bgr_0.V_TOP.t49 GNDA 0.36361f
C2165 bgr_0.V_TOP.n10 GNDA 0.243789f
C2166 bgr_0.V_TOP.t44 GNDA 0.36361f
C2167 bgr_0.V_TOP.t36 GNDA 0.369803f
C2168 bgr_0.V_TOP.n11 GNDA 0.380142f
C2169 bgr_0.V_TOP.t17 GNDA 0.369803f
C2170 bgr_0.V_TOP.t23 GNDA 0.36361f
C2171 bgr_0.V_TOP.n12 GNDA 0.243789f
C2172 bgr_0.V_TOP.t19 GNDA 0.36361f
C2173 bgr_0.V_TOP.t43 GNDA 0.369803f
C2174 bgr_0.V_TOP.n13 GNDA 0.380142f
C2175 bgr_0.V_TOP.t34 GNDA 0.369803f
C2176 bgr_0.V_TOP.t41 GNDA 0.36361f
C2177 bgr_0.V_TOP.n14 GNDA 0.311966f
C2178 bgr_0.V_TOP.t47 GNDA 0.36361f
C2179 bgr_0.V_TOP.n15 GNDA 0.159079f
C2180 bgr_0.V_TOP.n16 GNDA 0.544408f
C2181 bgr_0.V_TOP.t13 GNDA 0.102288f
C2182 bgr_0.V_TOP.n17 GNDA 0.724299f
C2183 bgr_0.V_TOP.n18 GNDA 0.022634f
C2184 bgr_0.V_TOP.n19 GNDA 0.414649f
C2185 bgr_0.V_TOP.n20 GNDA 0.021924f
C2186 bgr_0.V_TOP.n21 GNDA 0.022786f
C2187 bgr_0.V_TOP.n22 GNDA 0.022634f
C2188 bgr_0.V_TOP.n23 GNDA 0.209756f
C2189 bgr_0.V_TOP.n24 GNDA 0.127416f
C2190 bgr_0.V_TOP.n25 GNDA 0.072722f
C2191 bgr_0.V_TOP.n26 GNDA 0.022634f
C2192 bgr_0.V_TOP.n27 GNDA 0.125537f
C2193 bgr_0.V_TOP.n28 GNDA 0.022634f
C2194 bgr_0.V_TOP.n29 GNDA 0.124344f
C2195 bgr_0.V_TOP.n30 GNDA 0.273328f
C2196 bgr_0.V_TOP.n31 GNDA 0.019234f
C2197 bgr_0.V_TOP.n32 GNDA 0.04747f
C2198 bgr_0.V_TOP.n33 GNDA 0.050905f
C2199 bgr_0.V_TOP.n34 GNDA 0.050905f
C2200 bgr_0.V_TOP.n35 GNDA 0.050905f
C2201 bgr_0.V_TOP.n36 GNDA 0.050905f
C2202 bgr_0.V_TOP.n37 GNDA 0.050905f
C2203 bgr_0.V_TOP.n38 GNDA 0.050905f
C2204 bgr_0.V_TOP.n39 GNDA 0.04747f
C2205 bgr_0.V_TOP.t48 GNDA 0.109989f
C2206 VDDA.t285 GNDA 0.022433f
C2207 VDDA.t291 GNDA 0.022433f
C2208 VDDA.n0 GNDA 0.077741f
C2209 VDDA.n1 GNDA 0.076086f
C2210 VDDA.t309 GNDA 0.022433f
C2211 VDDA.n2 GNDA 0.067299f
C2212 VDDA.n3 GNDA 0.022433f
C2213 VDDA.n4 GNDA 0.012819f
C2214 VDDA.n7 GNDA 0.01038f
C2215 VDDA.n8 GNDA 0.012819f
C2216 VDDA.t353 GNDA 0.039332f
C2217 VDDA.t277 GNDA 0.022433f
C2218 VDDA.t273 GNDA 0.022433f
C2219 VDDA.n9 GNDA 0.077741f
C2220 VDDA.n10 GNDA 0.097414f
C2221 VDDA.n11 GNDA 0.033405f
C2222 VDDA.n12 GNDA 0.022433f
C2223 VDDA.n14 GNDA 0.022433f
C2224 VDDA.n15 GNDA 0.012819f
C2225 VDDA.n16 GNDA 0.012819f
C2226 VDDA.n17 GNDA 0.022433f
C2227 VDDA.n19 GNDA 0.022433f
C2228 VDDA.n20 GNDA 0.012819f
C2229 VDDA.n21 GNDA 0.012819f
C2230 VDDA.n22 GNDA 0.022433f
C2231 VDDA.n23 GNDA 0.022629f
C2232 VDDA.t355 GNDA 0.022433f
C2233 VDDA.n24 GNDA 0.067299f
C2234 VDDA.n25 GNDA 0.021625f
C2235 VDDA.n26 GNDA 0.012819f
C2236 VDDA.n27 GNDA 0.187476f
C2237 VDDA.t354 GNDA 0.162479f
C2238 VDDA.t276 GNDA 0.149981f
C2239 VDDA.t272 GNDA 0.149981f
C2240 VDDA.t284 GNDA 0.149981f
C2241 VDDA.t290 GNDA 0.149981f
C2242 VDDA.t252 GNDA 0.149981f
C2243 VDDA.t254 GNDA 0.149981f
C2244 VDDA.t266 GNDA 0.149981f
C2245 VDDA.t274 GNDA 0.149981f
C2246 VDDA.t286 GNDA 0.149981f
C2247 VDDA.t292 GNDA 0.149981f
C2248 VDDA.t308 GNDA 0.162479f
C2249 VDDA.n29 GNDA 0.01038f
C2250 VDDA.n30 GNDA 0.012819f
C2251 VDDA.n32 GNDA 0.022629f
C2252 VDDA.n33 GNDA 0.022433f
C2253 VDDA.n34 GNDA 0.012819f
C2254 VDDA.n35 GNDA 0.012819f
C2255 VDDA.n36 GNDA 0.022433f
C2256 VDDA.n38 GNDA 0.022433f
C2257 VDDA.n39 GNDA 0.022433f
C2258 VDDA.n40 GNDA 0.012819f
C2259 VDDA.n41 GNDA 0.187476f
C2260 VDDA.n43 GNDA 0.024495f
C2261 VDDA.t307 GNDA 0.039332f
C2262 VDDA.n44 GNDA 0.033405f
C2263 VDDA.t287 GNDA 0.022433f
C2264 VDDA.t293 GNDA 0.022433f
C2265 VDDA.n45 GNDA 0.077741f
C2266 VDDA.n46 GNDA 0.097414f
C2267 VDDA.t267 GNDA 0.022433f
C2268 VDDA.t275 GNDA 0.022433f
C2269 VDDA.n47 GNDA 0.077741f
C2270 VDDA.n48 GNDA 0.076086f
C2271 VDDA.n49 GNDA 0.02051f
C2272 VDDA.t253 GNDA 0.022433f
C2273 VDDA.t255 GNDA 0.022433f
C2274 VDDA.n50 GNDA 0.076131f
C2275 VDDA.n51 GNDA 0.087702f
C2276 VDDA.t296 GNDA 0.019228f
C2277 VDDA.t120 GNDA 0.019228f
C2278 VDDA.n52 GNDA 0.079517f
C2279 VDDA.t195 GNDA 0.019228f
C2280 VDDA.t446 GNDA 0.019228f
C2281 VDDA.n53 GNDA 0.079212f
C2282 VDDA.n54 GNDA 0.109827f
C2283 VDDA.t76 GNDA 0.019228f
C2284 VDDA.t42 GNDA 0.019228f
C2285 VDDA.n55 GNDA 0.079212f
C2286 VDDA.n56 GNDA 0.057309f
C2287 VDDA.t84 GNDA 0.019228f
C2288 VDDA.t27 GNDA 0.019228f
C2289 VDDA.n57 GNDA 0.079212f
C2290 VDDA.n58 GNDA 0.057309f
C2291 VDDA.t108 GNDA 0.019228f
C2292 VDDA.t26 GNDA 0.019228f
C2293 VDDA.n59 GNDA 0.079212f
C2294 VDDA.n60 GNDA 0.057309f
C2295 VDDA.t240 GNDA 0.019228f
C2296 VDDA.t297 GNDA 0.019228f
C2297 VDDA.n61 GNDA 0.079212f
C2298 VDDA.n62 GNDA 0.115606f
C2299 VDDA.t407 GNDA 0.019376f
C2300 VDDA.n64 GNDA 0.012819f
C2301 VDDA.n65 GNDA 0.010537f
C2302 VDDA.n66 GNDA 0.012819f
C2303 VDDA.t389 GNDA 0.02025f
C2304 VDDA.n67 GNDA 0.022433f
C2305 VDDA.n68 GNDA 0.012819f
C2306 VDDA.n69 GNDA 0.022433f
C2307 VDDA.n70 GNDA 0.031211f
C2308 VDDA.t391 GNDA 0.033797f
C2309 VDDA.n72 GNDA 0.051313f
C2310 VDDA.n74 GNDA 0.113447f
C2311 VDDA.t390 GNDA 0.094219f
C2312 VDDA.t196 GNDA 0.084605f
C2313 VDDA.t234 GNDA 0.084605f
C2314 VDDA.t109 GNDA 0.084605f
C2315 VDDA.t121 GNDA 0.084605f
C2316 VDDA.t20 GNDA 0.084605f
C2317 VDDA.t447 GNDA 0.084605f
C2318 VDDA.t175 GNDA 0.084605f
C2319 VDDA.t237 GNDA 0.084605f
C2320 VDDA.t77 GNDA 0.084605f
C2321 VDDA.t43 GNDA 0.084605f
C2322 VDDA.t408 GNDA 0.094219f
C2323 VDDA.n76 GNDA 0.012819f
C2324 VDDA.n77 GNDA 0.022433f
C2325 VDDA.n78 GNDA 0.022433f
C2326 VDDA.t409 GNDA 0.033797f
C2327 VDDA.n79 GNDA 0.028257f
C2328 VDDA.n80 GNDA 0.013491f
C2329 VDDA.n81 GNDA 0.113447f
C2330 VDDA.n82 GNDA 0.012819f
C2331 VDDA.n83 GNDA 0.025423f
C2332 VDDA.n84 GNDA 0.041082f
C2333 VDDA.n85 GNDA 0.161985f
C2334 VDDA.t312 GNDA 0.011691f
C2335 VDDA.n86 GNDA 0.053162f
C2336 VDDA.t311 GNDA 0.047946f
C2337 VDDA.t192 GNDA 0.031727f
C2338 VDDA.t229 GNDA 0.031727f
C2339 VDDA.t142 GNDA 0.031727f
C2340 VDDA.t251 GNDA 0.031727f
C2341 VDDA.t12 GNDA 0.031727f
C2342 VDDA.t148 GNDA 0.031727f
C2343 VDDA.t62 GNDA 0.031727f
C2344 VDDA.t3 GNDA 0.031727f
C2345 VDDA.t63 GNDA 0.031727f
C2346 VDDA.t149 GNDA 0.031727f
C2347 VDDA.t302 GNDA 0.047682f
C2348 VDDA.t303 GNDA 0.011691f
C2349 VDDA.n87 GNDA 0.02772f
C2350 VDDA.n88 GNDA 0.03966f
C2351 VDDA.n89 GNDA 0.084431f
C2352 VDDA.t439 GNDA 0.038457f
C2353 VDDA.t22 GNDA 0.038457f
C2354 VDDA.n90 GNDA 0.154283f
C2355 VDDA.n91 GNDA 0.07838f
C2356 VDDA.n93 GNDA 0.012819f
C2357 VDDA.n99 GNDA 0.013491f
C2358 VDDA.n100 GNDA 0.012819f
C2359 VDDA.t341 GNDA 0.046596f
C2360 VDDA.t441 GNDA 0.038457f
C2361 VDDA.t7 GNDA 0.038457f
C2362 VDDA.n101 GNDA 0.154283f
C2363 VDDA.n102 GNDA 0.07838f
C2364 VDDA.t236 GNDA 0.038457f
C2365 VDDA.t194 GNDA 0.038457f
C2366 VDDA.n103 GNDA 0.154283f
C2367 VDDA.n104 GNDA 0.07838f
C2368 VDDA.t239 GNDA 0.038457f
C2369 VDDA.t198 GNDA 0.038457f
C2370 VDDA.n105 GNDA 0.154283f
C2371 VDDA.n106 GNDA 0.07838f
C2372 VDDA.t242 GNDA 0.038457f
C2373 VDDA.t9 GNDA 0.038457f
C2374 VDDA.n107 GNDA 0.154283f
C2375 VDDA.n108 GNDA 0.099184f
C2376 VDDA.n109 GNDA 0.038361f
C2377 VDDA.n110 GNDA 0.025503f
C2378 VDDA.n111 GNDA 0.012819f
C2379 VDDA.n112 GNDA 0.012819f
C2380 VDDA.n113 GNDA 0.022433f
C2381 VDDA.n114 GNDA 0.012819f
C2382 VDDA.n115 GNDA 0.012819f
C2383 VDDA.n116 GNDA 0.012819f
C2384 VDDA.n117 GNDA 0.012819f
C2385 VDDA.n118 GNDA 0.022433f
C2386 VDDA.n119 GNDA 0.025503f
C2387 VDDA.n120 GNDA 0.012819f
C2388 VDDA.n121 GNDA 0.012819f
C2389 VDDA.n122 GNDA 0.012819f
C2390 VDDA.n123 GNDA 0.032471f
C2391 VDDA.n124 GNDA 0.022433f
C2392 VDDA.n125 GNDA 0.022433f
C2393 VDDA.n126 GNDA 0.022433f
C2394 VDDA.n127 GNDA 0.012819f
C2395 VDDA.n128 GNDA 0.012819f
C2396 VDDA.n130 GNDA 0.022433f
C2397 VDDA.n131 GNDA 0.022433f
C2398 VDDA.n133 GNDA 0.012819f
C2399 VDDA.n134 GNDA 0.012819f
C2400 VDDA.n135 GNDA 0.022433f
C2401 VDDA.n136 GNDA 0.022433f
C2402 VDDA.n137 GNDA 0.022433f
C2403 VDDA.n139 GNDA 0.025423f
C2404 VDDA.n140 GNDA 0.012819f
C2405 VDDA.n141 GNDA 0.302526f
C2406 VDDA.t342 GNDA 0.25125f
C2407 VDDA.t241 GNDA 0.225612f
C2408 VDDA.t8 GNDA 0.225612f
C2409 VDDA.t238 GNDA 0.225612f
C2410 VDDA.t197 GNDA 0.225612f
C2411 VDDA.t235 GNDA 0.225612f
C2412 VDDA.t193 GNDA 0.225612f
C2413 VDDA.t440 GNDA 0.225612f
C2414 VDDA.t6 GNDA 0.225612f
C2415 VDDA.t438 GNDA 0.225612f
C2416 VDDA.t21 GNDA 0.225612f
C2417 VDDA.t357 GNDA 0.25125f
C2418 VDDA.n146 GNDA 0.013491f
C2419 VDDA.n147 GNDA 0.012819f
C2420 VDDA.n148 GNDA 0.022433f
C2421 VDDA.n149 GNDA 0.025503f
C2422 VDDA.n150 GNDA 0.012819f
C2423 VDDA.n151 GNDA 0.012819f
C2424 VDDA.n154 GNDA 0.012819f
C2425 VDDA.n155 GNDA 0.012819f
C2426 VDDA.n156 GNDA 0.025503f
C2427 VDDA.n157 GNDA 0.032471f
C2428 VDDA.n158 GNDA 0.012819f
C2429 VDDA.n159 GNDA 0.022433f
C2430 VDDA.n160 GNDA 0.022433f
C2431 VDDA.n161 GNDA 0.012819f
C2432 VDDA.n162 GNDA 0.012819f
C2433 VDDA.n163 GNDA 0.022433f
C2434 VDDA.n164 GNDA 0.022433f
C2435 VDDA.n165 GNDA 0.012819f
C2436 VDDA.n166 GNDA 0.012819f
C2437 VDDA.n167 GNDA 0.022433f
C2438 VDDA.n168 GNDA 0.022433f
C2439 VDDA.n169 GNDA 0.012819f
C2440 VDDA.n170 GNDA 0.012819f
C2441 VDDA.n171 GNDA 0.022433f
C2442 VDDA.n172 GNDA 0.022433f
C2443 VDDA.n173 GNDA 0.022433f
C2444 VDDA.n174 GNDA 0.012819f
C2445 VDDA.n175 GNDA 0.302526f
C2446 VDDA.n177 GNDA 0.028293f
C2447 VDDA.t356 GNDA 0.046596f
C2448 VDDA.n178 GNDA 0.037513f
C2449 VDDA.n179 GNDA 0.052145f
C2450 VDDA.n180 GNDA 0.035204f
C2451 VDDA.n182 GNDA 0.049075f
C2452 VDDA.t397 GNDA 0.011678f
C2453 VDDA.n184 GNDA 0.049075f
C2454 VDDA.n186 GNDA 0.049075f
C2455 VDDA.n188 GNDA 0.049075f
C2456 VDDA.n190 GNDA 0.049075f
C2457 VDDA.n192 GNDA 0.049075f
C2458 VDDA.n194 GNDA 0.049075f
C2459 VDDA.n196 GNDA 0.049075f
C2460 VDDA.n198 GNDA 0.049075f
C2461 VDDA.n200 GNDA 0.06988f
C2462 VDDA.n201 GNDA 0.021167f
C2463 VDDA.n202 GNDA 0.038717f
C2464 VDDA.t396 GNDA 0.04799f
C2465 VDDA.t136 GNDA 0.031727f
C2466 VDDA.t106 GNDA 0.031727f
C2467 VDDA.t104 GNDA 0.031727f
C2468 VDDA.t423 GNDA 0.031727f
C2469 VDDA.t85 GNDA 0.031727f
C2470 VDDA.t185 GNDA 0.031727f
C2471 VDDA.t102 GNDA 0.031727f
C2472 VDDA.t460 GNDA 0.031727f
C2473 VDDA.t464 GNDA 0.031727f
C2474 VDDA.t434 GNDA 0.031727f
C2475 VDDA.t58 GNDA 0.031727f
C2476 VDDA.t455 GNDA 0.031727f
C2477 VDDA.t457 GNDA 0.031727f
C2478 VDDA.t138 GNDA 0.031727f
C2479 VDDA.t467 GNDA 0.031727f
C2480 VDDA.t91 GNDA 0.031727f
C2481 VDDA.t436 GNDA 0.031727f
C2482 VDDA.t159 GNDA 0.031727f
C2483 VDDA.t18 GNDA 0.031727f
C2484 VDDA.t34 GNDA 0.031727f
C2485 VDDA.t402 GNDA 0.04603f
C2486 VDDA.t403 GNDA 0.011678f
C2487 VDDA.n203 GNDA 0.035069f
C2488 VDDA.n204 GNDA 0.020319f
C2489 VDDA.n205 GNDA 0.064374f
C2490 VDDA.n206 GNDA 0.0877f
C2491 VDDA.n207 GNDA 0.152164f
C2492 VDDA.t269 GNDA 0.022433f
C2493 VDDA.t279 GNDA 0.022433f
C2494 VDDA.n208 GNDA 0.077741f
C2495 VDDA.n209 GNDA 0.076086f
C2496 VDDA.t400 GNDA 0.022433f
C2497 VDDA.n210 GNDA 0.067299f
C2498 VDDA.n211 GNDA 0.022433f
C2499 VDDA.n212 GNDA 0.012819f
C2500 VDDA.n215 GNDA 0.01038f
C2501 VDDA.n216 GNDA 0.012819f
C2502 VDDA.t322 GNDA 0.039332f
C2503 VDDA.t265 GNDA 0.022433f
C2504 VDDA.t261 GNDA 0.022433f
C2505 VDDA.n217 GNDA 0.077741f
C2506 VDDA.n218 GNDA 0.097414f
C2507 VDDA.n219 GNDA 0.033405f
C2508 VDDA.n220 GNDA 0.022433f
C2509 VDDA.n222 GNDA 0.022433f
C2510 VDDA.n223 GNDA 0.012819f
C2511 VDDA.n224 GNDA 0.012819f
C2512 VDDA.n225 GNDA 0.022433f
C2513 VDDA.n227 GNDA 0.022433f
C2514 VDDA.n228 GNDA 0.012819f
C2515 VDDA.n229 GNDA 0.012819f
C2516 VDDA.n230 GNDA 0.022433f
C2517 VDDA.n231 GNDA 0.022629f
C2518 VDDA.t324 GNDA 0.022433f
C2519 VDDA.n232 GNDA 0.067299f
C2520 VDDA.n233 GNDA 0.021625f
C2521 VDDA.n234 GNDA 0.012819f
C2522 VDDA.n235 GNDA 0.187476f
C2523 VDDA.t323 GNDA 0.162479f
C2524 VDDA.t264 GNDA 0.149981f
C2525 VDDA.t260 GNDA 0.149981f
C2526 VDDA.t268 GNDA 0.149981f
C2527 VDDA.t278 GNDA 0.149981f
C2528 VDDA.t288 GNDA 0.149981f
C2529 VDDA.t258 GNDA 0.149981f
C2530 VDDA.t256 GNDA 0.149981f
C2531 VDDA.t262 GNDA 0.149981f
C2532 VDDA.t270 GNDA 0.149981f
C2533 VDDA.t282 GNDA 0.149981f
C2534 VDDA.t399 GNDA 0.162479f
C2535 VDDA.n237 GNDA 0.01038f
C2536 VDDA.n238 GNDA 0.012819f
C2537 VDDA.n240 GNDA 0.022629f
C2538 VDDA.n241 GNDA 0.022433f
C2539 VDDA.n242 GNDA 0.012819f
C2540 VDDA.n243 GNDA 0.012819f
C2541 VDDA.n244 GNDA 0.022433f
C2542 VDDA.n246 GNDA 0.022433f
C2543 VDDA.n247 GNDA 0.022433f
C2544 VDDA.n248 GNDA 0.012819f
C2545 VDDA.n249 GNDA 0.187476f
C2546 VDDA.n251 GNDA 0.024495f
C2547 VDDA.t398 GNDA 0.039332f
C2548 VDDA.n252 GNDA 0.033405f
C2549 VDDA.t271 GNDA 0.022433f
C2550 VDDA.t283 GNDA 0.022433f
C2551 VDDA.n253 GNDA 0.077741f
C2552 VDDA.n254 GNDA 0.097414f
C2553 VDDA.t257 GNDA 0.022433f
C2554 VDDA.t263 GNDA 0.022433f
C2555 VDDA.n255 GNDA 0.077741f
C2556 VDDA.n256 GNDA 0.076086f
C2557 VDDA.n257 GNDA 0.02051f
C2558 VDDA.t289 GNDA 0.022433f
C2559 VDDA.t259 GNDA 0.022433f
C2560 VDDA.n258 GNDA 0.076131f
C2561 VDDA.n259 GNDA 0.087702f
C2562 VDDA.t129 GNDA 0.019228f
C2563 VDDA.t295 GNDA 0.019228f
C2564 VDDA.n260 GNDA 0.079517f
C2565 VDDA.t180 GNDA 0.019228f
C2566 VDDA.t69 GNDA 0.019228f
C2567 VDDA.n261 GNDA 0.079212f
C2568 VDDA.n262 GNDA 0.109827f
C2569 VDDA.t450 GNDA 0.019228f
C2570 VDDA.t75 GNDA 0.019228f
C2571 VDDA.n263 GNDA 0.079212f
C2572 VDDA.n264 GNDA 0.057309f
C2573 VDDA.t463 GNDA 0.019228f
C2574 VDDA.t0 GNDA 0.019228f
C2575 VDDA.n265 GNDA 0.079212f
C2576 VDDA.n266 GNDA 0.057309f
C2577 VDDA.t158 GNDA 0.019228f
C2578 VDDA.t182 GNDA 0.019228f
C2579 VDDA.n267 GNDA 0.079212f
C2580 VDDA.n268 GNDA 0.057309f
C2581 VDDA.t294 GNDA 0.019228f
C2582 VDDA.t222 GNDA 0.019228f
C2583 VDDA.n269 GNDA 0.079212f
C2584 VDDA.n270 GNDA 0.115606f
C2585 VDDA.t362 GNDA 0.019376f
C2586 VDDA.n271 GNDA 0.012819f
C2587 VDDA.t364 GNDA 0.033797f
C2588 VDDA.n272 GNDA 0.012819f
C2589 VDDA.n273 GNDA 0.012819f
C2590 VDDA.n275 GNDA 0.010537f
C2591 VDDA.n276 GNDA 0.012819f
C2592 VDDA.t377 GNDA 0.02025f
C2593 VDDA.n277 GNDA 0.022433f
C2594 VDDA.n278 GNDA 0.012819f
C2595 VDDA.n279 GNDA 0.022433f
C2596 VDDA.n280 GNDA 0.031211f
C2597 VDDA.t379 GNDA 0.033797f
C2598 VDDA.n282 GNDA 0.051313f
C2599 VDDA.n284 GNDA 0.113447f
C2600 VDDA.t378 GNDA 0.094219f
C2601 VDDA.t181 GNDA 0.084605f
C2602 VDDA.t157 GNDA 0.084605f
C2603 VDDA.t429 GNDA 0.084605f
C2604 VDDA.t466 GNDA 0.084605f
C2605 VDDA.t459 GNDA 0.084605f
C2606 VDDA.t184 GNDA 0.084605f
C2607 VDDA.t183 GNDA 0.084605f
C2608 VDDA.t64 GNDA 0.084605f
C2609 VDDA.t174 GNDA 0.084605f
C2610 VDDA.t462 GNDA 0.084605f
C2611 VDDA.t363 GNDA 0.094219f
C2612 VDDA.n285 GNDA 0.113447f
C2613 VDDA.n286 GNDA 0.013491f
C2614 VDDA.n287 GNDA 0.028257f
C2615 VDDA.n288 GNDA 0.022433f
C2616 VDDA.n289 GNDA 0.022433f
C2617 VDDA.n291 GNDA 0.025423f
C2618 VDDA.n292 GNDA 0.041082f
C2619 VDDA.n293 GNDA 0.161985f
C2620 VDDA.t388 GNDA 0.011691f
C2621 VDDA.n294 GNDA 0.02772f
C2622 VDDA.t370 GNDA 0.011691f
C2623 VDDA.n295 GNDA 0.053162f
C2624 VDDA.t369 GNDA 0.047946f
C2625 VDDA.t150 GNDA 0.031727f
C2626 VDDA.t94 GNDA 0.031727f
C2627 VDDA.t25 GNDA 0.031727f
C2628 VDDA.t205 GNDA 0.031727f
C2629 VDDA.t145 GNDA 0.031727f
C2630 VDDA.t243 GNDA 0.031727f
C2631 VDDA.t13 GNDA 0.031727f
C2632 VDDA.t161 GNDA 0.031727f
C2633 VDDA.t415 GNDA 0.031727f
C2634 VDDA.t187 GNDA 0.031727f
C2635 VDDA.t387 GNDA 0.047682f
C2636 VDDA.n296 GNDA 0.03966f
C2637 VDDA.n297 GNDA 0.084431f
C2638 VDDA.t135 GNDA 0.038457f
C2639 VDDA.t211 GNDA 0.038457f
C2640 VDDA.n298 GNDA 0.154283f
C2641 VDDA.n299 GNDA 0.07838f
C2642 VDDA.n301 GNDA 0.012819f
C2643 VDDA.n306 GNDA 0.013491f
C2644 VDDA.n312 GNDA 0.013491f
C2645 VDDA.n313 GNDA 0.012819f
C2646 VDDA.t325 GNDA 0.046596f
C2647 VDDA.t17 GNDA 0.038457f
C2648 VDDA.t154 GNDA 0.038457f
C2649 VDDA.n314 GNDA 0.154283f
C2650 VDDA.n315 GNDA 0.07838f
C2651 VDDA.t156 GNDA 0.038457f
C2652 VDDA.t428 GNDA 0.038457f
C2653 VDDA.n316 GNDA 0.154283f
C2654 VDDA.n317 GNDA 0.07838f
C2655 VDDA.t452 GNDA 0.038457f
C2656 VDDA.t173 GNDA 0.038457f
C2657 VDDA.n318 GNDA 0.154283f
C2658 VDDA.n319 GNDA 0.07838f
C2659 VDDA.t15 GNDA 0.038457f
C2660 VDDA.t454 GNDA 0.038457f
C2661 VDDA.n320 GNDA 0.154283f
C2662 VDDA.n321 GNDA 0.099184f
C2663 VDDA.n322 GNDA 0.038361f
C2664 VDDA.n323 GNDA 0.022433f
C2665 VDDA.n324 GNDA 0.012819f
C2666 VDDA.n325 GNDA 0.012819f
C2667 VDDA.n328 GNDA 0.012819f
C2668 VDDA.n329 GNDA 0.012819f
C2669 VDDA.n330 GNDA 0.025503f
C2670 VDDA.n331 GNDA 0.032471f
C2671 VDDA.n332 GNDA 0.012819f
C2672 VDDA.n333 GNDA 0.022433f
C2673 VDDA.n334 GNDA 0.022433f
C2674 VDDA.n335 GNDA 0.012819f
C2675 VDDA.n336 GNDA 0.012819f
C2676 VDDA.n337 GNDA 0.022433f
C2677 VDDA.n338 GNDA 0.022433f
C2678 VDDA.n339 GNDA 0.012819f
C2679 VDDA.n340 GNDA 0.012819f
C2680 VDDA.n341 GNDA 0.022433f
C2681 VDDA.n342 GNDA 0.022433f
C2682 VDDA.n343 GNDA 0.012819f
C2683 VDDA.n344 GNDA 0.012819f
C2684 VDDA.n345 GNDA 0.022433f
C2685 VDDA.n346 GNDA 0.022433f
C2686 VDDA.n347 GNDA 0.012819f
C2687 VDDA.n348 GNDA 0.012819f
C2688 VDDA.n349 GNDA 0.022433f
C2689 VDDA.n350 GNDA 0.025503f
C2690 VDDA.n352 GNDA 0.025423f
C2691 VDDA.n353 GNDA 0.012819f
C2692 VDDA.n354 GNDA 0.302526f
C2693 VDDA.t326 GNDA 0.25125f
C2694 VDDA.t453 GNDA 0.225612f
C2695 VDDA.t14 GNDA 0.225612f
C2696 VDDA.t172 GNDA 0.225612f
C2697 VDDA.t451 GNDA 0.225612f
C2698 VDDA.t427 GNDA 0.225612f
C2699 VDDA.t155 GNDA 0.225612f
C2700 VDDA.t153 GNDA 0.225612f
C2701 VDDA.t16 GNDA 0.225612f
C2702 VDDA.t210 GNDA 0.225612f
C2703 VDDA.t134 GNDA 0.225612f
C2704 VDDA.t317 GNDA 0.25125f
C2705 VDDA.n355 GNDA 0.012819f
C2706 VDDA.n356 GNDA 0.022433f
C2707 VDDA.n357 GNDA 0.025503f
C2708 VDDA.n358 GNDA 0.012819f
C2709 VDDA.n359 GNDA 0.012819f
C2710 VDDA.n362 GNDA 0.012819f
C2711 VDDA.n363 GNDA 0.012819f
C2712 VDDA.n364 GNDA 0.025503f
C2713 VDDA.n365 GNDA 0.032471f
C2714 VDDA.n366 GNDA 0.012819f
C2715 VDDA.n367 GNDA 0.022433f
C2716 VDDA.n368 GNDA 0.022433f
C2717 VDDA.n369 GNDA 0.012819f
C2718 VDDA.n370 GNDA 0.012819f
C2719 VDDA.n371 GNDA 0.022433f
C2720 VDDA.n372 GNDA 0.022433f
C2721 VDDA.n373 GNDA 0.012819f
C2722 VDDA.n374 GNDA 0.012819f
C2723 VDDA.n375 GNDA 0.022433f
C2724 VDDA.n376 GNDA 0.022433f
C2725 VDDA.n377 GNDA 0.012819f
C2726 VDDA.n378 GNDA 0.012819f
C2727 VDDA.n379 GNDA 0.022433f
C2728 VDDA.n380 GNDA 0.022433f
C2729 VDDA.n381 GNDA 0.022433f
C2730 VDDA.n382 GNDA 0.012819f
C2731 VDDA.n383 GNDA 0.302526f
C2732 VDDA.n385 GNDA 0.028293f
C2733 VDDA.t316 GNDA 0.046596f
C2734 VDDA.n386 GNDA 0.037513f
C2735 VDDA.n387 GNDA 0.052145f
C2736 VDDA.n388 GNDA 0.102562f
C2737 VDDA.n389 GNDA 0.156901f
C2738 VDDA.n390 GNDA 0.14022f
C2739 VDDA.t191 GNDA 0.011537f
C2740 VDDA.t339 GNDA 0.011537f
C2741 VDDA.n391 GNDA 0.026769f
C2742 VDDA.n392 GNDA 0.086851f
C2743 VDDA.t330 GNDA 0.040934f
C2744 VDDA.t337 GNDA 0.023666f
C2745 VDDA.n393 GNDA 0.046815f
C2746 VDDA.t340 GNDA 0.040934f
C2747 VDDA.n394 GNDA 0.07685f
C2748 VDDA.t338 GNDA 0.137161f
C2749 VDDA.t190 GNDA 0.084605f
C2750 VDDA.t329 GNDA 0.137161f
C2751 VDDA.n395 GNDA 0.07685f
C2752 VDDA.t328 GNDA 0.023666f
C2753 VDDA.n396 GNDA 0.046487f
C2754 VDDA.n397 GNDA 0.043496f
C2755 VDDA.n398 GNDA 0.061626f
C2756 VDDA.n399 GNDA 0.09036f
C2757 VDDA.t382 GNDA 0.022433f
C2758 VDDA.n400 GNDA 0.067299f
C2759 VDDA.n401 GNDA 0.022433f
C2760 VDDA.n402 GNDA 0.012819f
C2761 VDDA.n405 GNDA 0.01038f
C2762 VDDA.n406 GNDA 0.012819f
C2763 VDDA.t359 GNDA 0.039332f
C2764 VDDA.n407 GNDA 0.032767f
C2765 VDDA.n408 GNDA 0.022433f
C2766 VDDA.n410 GNDA 0.022433f
C2767 VDDA.n411 GNDA 0.012819f
C2768 VDDA.n412 GNDA 0.012819f
C2769 VDDA.n413 GNDA 0.022433f
C2770 VDDA.n415 GNDA 0.022433f
C2771 VDDA.n416 GNDA 0.012819f
C2772 VDDA.n417 GNDA 0.012819f
C2773 VDDA.n418 GNDA 0.022433f
C2774 VDDA.n419 GNDA 0.022629f
C2775 VDDA.t281 GNDA 0.022433f
C2776 VDDA.n420 GNDA 0.077741f
C2777 VDDA.t361 GNDA 0.044866f
C2778 VDDA.n421 GNDA 0.067299f
C2779 VDDA.n422 GNDA 0.021625f
C2780 VDDA.n423 GNDA 0.012819f
C2781 VDDA.n424 GNDA 0.187476f
C2782 VDDA.t360 GNDA 0.162479f
C2783 VDDA.t280 GNDA 0.149981f
C2784 VDDA.t381 GNDA 0.162479f
C2785 VDDA.n426 GNDA 0.01038f
C2786 VDDA.n427 GNDA 0.012819f
C2787 VDDA.n429 GNDA 0.022629f
C2788 VDDA.n430 GNDA 0.022433f
C2789 VDDA.n431 GNDA 0.012819f
C2790 VDDA.n432 GNDA 0.012819f
C2791 VDDA.n433 GNDA 0.022433f
C2792 VDDA.n435 GNDA 0.022433f
C2793 VDDA.n436 GNDA 0.022433f
C2794 VDDA.n437 GNDA 0.012819f
C2795 VDDA.n438 GNDA 0.187476f
C2796 VDDA.n440 GNDA 0.024495f
C2797 VDDA.t380 GNDA 0.039332f
C2798 VDDA.n441 GNDA 0.032439f
C2799 VDDA.n442 GNDA 0.043496f
C2800 VDDA.n443 GNDA 0.181871f
C2801 VDDA.n444 GNDA 3.444f
C2802 VDDA.t67 GNDA 0.358288f
C2803 VDDA.t209 GNDA 0.359586f
C2804 VDDA.t54 GNDA 0.340358f
C2805 VDDA.t422 GNDA 0.358288f
C2806 VDDA.t101 GNDA 0.359586f
C2807 VDDA.t170 GNDA 0.340358f
C2808 VDDA.t169 GNDA 0.358288f
C2809 VDDA.t168 GNDA 0.359586f
C2810 VDDA.t124 GNDA 0.340358f
C2811 VDDA.t98 GNDA 0.358288f
C2812 VDDA.t72 GNDA 0.359586f
C2813 VDDA.t206 GNDA 0.340358f
C2814 VDDA.t214 GNDA 0.358288f
C2815 VDDA.t55 GNDA 0.359586f
C2816 VDDA.t100 GNDA 0.340358f
C2817 VDDA.n445 GNDA 0.240161f
C2818 VDDA.t215 GNDA 0.191253f
C2819 VDDA.n446 GNDA 0.26058f
C2820 VDDA.t99 GNDA 0.191253f
C2821 VDDA.n447 GNDA 0.26058f
C2822 VDDA.t171 GNDA 0.191253f
C2823 VDDA.n448 GNDA 0.26058f
C2824 VDDA.t97 GNDA 0.191253f
C2825 VDDA.n449 GNDA 0.26058f
C2826 VDDA.t68 GNDA 0.335043f
C2827 VDDA.n450 GNDA 2.97549f
C2828 VDDA.t469 GNDA 0.708591f
C2829 VDDA.t471 GNDA 0.755222f
C2830 VDDA.t472 GNDA 0.754926f
C2831 VDDA.t470 GNDA 0.726508f
C2832 VDDA.n451 GNDA 0.505724f
C2833 VDDA.n452 GNDA 0.24835f
C2834 VDDA.n453 GNDA 0.360996f
C2835 VDDA.n454 GNDA 0.658955f
C2836 VDDA.n455 GNDA 0.016121f
C2837 VDDA.n456 GNDA 0.065279f
C2838 VDDA.n457 GNDA 0.027107f
C2839 VDDA.t352 GNDA 0.022294f
C2840 VDDA.n459 GNDA 0.027107f
C2841 VDDA.n460 GNDA 0.016121f
C2842 VDDA.n461 GNDA 0.065279f
C2843 VDDA.t336 GNDA 0.02245f
C2844 VDDA.n462 GNDA 0.027107f
C2845 VDDA.n463 GNDA 0.016121f
C2846 VDDA.n464 GNDA 0.065279f
C2847 VDDA.n465 GNDA 0.016121f
C2848 VDDA.n466 GNDA 0.065279f
C2849 VDDA.n467 GNDA 0.016121f
C2850 VDDA.n468 GNDA 0.065279f
C2851 VDDA.n469 GNDA 0.016121f
C2852 VDDA.n470 GNDA 0.065279f
C2853 VDDA.n471 GNDA 0.016121f
C2854 VDDA.n472 GNDA 0.065279f
C2855 VDDA.n473 GNDA 0.016121f
C2856 VDDA.n474 GNDA 0.065279f
C2857 VDDA.n475 GNDA 0.016121f
C2858 VDDA.n476 GNDA 0.065279f
C2859 VDDA.n477 GNDA 0.016121f
C2860 VDDA.n478 GNDA 0.09381f
C2861 VDDA.n479 GNDA 0.024854f
C2862 VDDA.t313 GNDA 0.02366f
C2863 VDDA.t315 GNDA 0.022294f
C2864 VDDA.n480 GNDA 0.042734f
C2865 VDDA.n481 GNDA 0.06496f
C2866 VDDA.t314 GNDA 0.080563f
C2867 VDDA.t249 GNDA 0.053839f
C2868 VDDA.t40 GNDA 0.053839f
C2869 VDDA.t4 GNDA 0.053839f
C2870 VDDA.t50 GNDA 0.053839f
C2871 VDDA.t130 GNDA 0.053839f
C2872 VDDA.t89 GNDA 0.053839f
C2873 VDDA.t87 GNDA 0.053839f
C2874 VDDA.t225 GNDA 0.053839f
C2875 VDDA.t164 GNDA 0.053839f
C2876 VDDA.t432 GNDA 0.053839f
C2877 VDDA.t48 GNDA 0.053839f
C2878 VDDA.t38 GNDA 0.053839f
C2879 VDDA.t176 GNDA 0.053839f
C2880 VDDA.t46 GNDA 0.053839f
C2881 VDDA.t116 GNDA 0.053839f
C2882 VDDA.t132 GNDA 0.053839f
C2883 VDDA.t30 GNDA 0.053839f
C2884 VDDA.t118 GNDA 0.053839f
C2885 VDDA.t335 GNDA 0.082124f
C2886 VDDA.n482 GNDA 0.116935f
C2887 VDDA.t334 GNDA 0.015866f
C2888 VDDA.n483 GNDA 0.026219f
C2889 VDDA.n484 GNDA 0.047745f
C2890 VDDA.n485 GNDA 0.016121f
C2891 VDDA.n486 GNDA 0.065279f
C2892 VDDA.n487 GNDA 0.016121f
C2893 VDDA.n488 GNDA 0.065279f
C2894 VDDA.n489 GNDA 0.016121f
C2895 VDDA.n490 GNDA 0.065279f
C2896 VDDA.n491 GNDA 0.016121f
C2897 VDDA.n492 GNDA 0.065279f
C2898 VDDA.n493 GNDA 0.016121f
C2899 VDDA.n494 GNDA 0.065279f
C2900 VDDA.n495 GNDA 0.016121f
C2901 VDDA.n496 GNDA 0.065279f
C2902 VDDA.n497 GNDA 0.016121f
C2903 VDDA.n498 GNDA 0.065279f
C2904 VDDA.n499 GNDA 0.016121f
C2905 VDDA.n500 GNDA 0.065279f
C2906 VDDA.n501 GNDA 0.047745f
C2907 VDDA.n502 GNDA 0.023587f
C2908 VDDA.t371 GNDA 0.02366f
C2909 VDDA.t373 GNDA 0.022294f
C2910 VDDA.n503 GNDA 0.042734f
C2911 VDDA.n504 GNDA 0.06496f
C2912 VDDA.t372 GNDA 0.080563f
C2913 VDDA.t143 GNDA 0.053839f
C2914 VDDA.t188 GNDA 0.053839f
C2915 VDDA.t230 GNDA 0.053839f
C2916 VDDA.t32 GNDA 0.053839f
C2917 VDDA.t413 GNDA 0.053839f
C2918 VDDA.t232 GNDA 0.053839f
C2919 VDDA.t178 GNDA 0.053839f
C2920 VDDA.t151 GNDA 0.053839f
C2921 VDDA.t1 GNDA 0.053839f
C2922 VDDA.t162 GNDA 0.053839f
C2923 VDDA.t122 GNDA 0.053839f
C2924 VDDA.t36 GNDA 0.053839f
C2925 VDDA.t416 GNDA 0.053839f
C2926 VDDA.t247 GNDA 0.053839f
C2927 VDDA.t227 GNDA 0.053839f
C2928 VDDA.t140 GNDA 0.053839f
C2929 VDDA.t146 GNDA 0.053839f
C2930 VDDA.t425 GNDA 0.053839f
C2931 VDDA.t351 GNDA 0.066516f
C2932 VDDA.n505 GNDA 0.079007f
C2933 VDDA.n506 GNDA 0.042907f
C2934 VDDA.t350 GNDA 0.023648f
C2935 VDDA.n507 GNDA 0.023587f
C2936 VDDA.n508 GNDA 0.11065f
C2937 VDDA.n509 GNDA 0.213341f
C2938 VDDA.t71 GNDA 0.019228f
C2939 VDDA.t167 GNDA 0.019228f
C2940 VDDA.n510 GNDA 0.063524f
C2941 VDDA.n511 GNDA 0.08197f
C2942 VDDA.n513 GNDA 0.012819f
C2943 VDDA.n516 GNDA 0.012819f
C2944 VDDA.n517 GNDA 0.012819f
C2945 VDDA.n518 GNDA 0.022299f
C2946 VDDA.n519 GNDA 0.012819f
C2947 VDDA.n520 GNDA 0.012819f
C2948 VDDA.n521 GNDA 0.012819f
C2949 VDDA.n522 GNDA 0.022433f
C2950 VDDA.t331 GNDA 0.091688f
C2951 VDDA.t365 GNDA 0.012151f
C2952 VDDA.n523 GNDA 0.031486f
C2953 VDDA.t412 GNDA 0.025591f
C2954 VDDA.t367 GNDA 0.02245f
C2955 VDDA.n524 GNDA 0.112312f
C2956 VDDA.t366 GNDA 0.077774f
C2957 VDDA.t93 GNDA 0.049353f
C2958 VDDA.t244 GNDA 0.049353f
C2959 VDDA.t411 GNDA 0.079486f
C2960 VDDA.n525 GNDA 0.117627f
C2961 VDDA.t410 GNDA 0.012151f
C2962 VDDA.n526 GNDA 0.031246f
C2963 VDDA.n527 GNDA 0.093994f
C2964 VDDA.t66 GNDA 0.019228f
C2965 VDDA.t53 GNDA 0.019228f
C2966 VDDA.n528 GNDA 0.063524f
C2967 VDDA.n529 GNDA 0.08197f
C2968 VDDA.t419 GNDA 0.019228f
C2969 VDDA.t421 GNDA 0.019228f
C2970 VDDA.n530 GNDA 0.063524f
C2971 VDDA.n531 GNDA 0.08197f
C2972 VDDA.t128 GNDA 0.019228f
C2973 VDDA.t219 GNDA 0.019228f
C2974 VDDA.n532 GNDA 0.063524f
C2975 VDDA.n533 GNDA 0.08197f
C2976 VDDA.t217 GNDA 0.019228f
C2977 VDDA.t57 GNDA 0.019228f
C2978 VDDA.n534 GNDA 0.063524f
C2979 VDDA.n535 GNDA 0.08197f
C2980 VDDA.t126 GNDA 0.019228f
C2981 VDDA.t74 GNDA 0.019228f
C2982 VDDA.n536 GNDA 0.063524f
C2983 VDDA.n537 GNDA 0.08197f
C2984 VDDA.t96 GNDA 0.019228f
C2985 VDDA.t208 GNDA 0.019228f
C2986 VDDA.n538 GNDA 0.063524f
C2987 VDDA.n539 GNDA 0.08197f
C2988 VDDA.t221 GNDA 0.019228f
C2989 VDDA.t213 GNDA 0.019228f
C2990 VDDA.n540 GNDA 0.063524f
C2991 VDDA.n541 GNDA 0.08197f
C2992 VDDA.n542 GNDA 0.043765f
C2993 VDDA.n543 GNDA 0.034243f
C2994 VDDA.n544 GNDA 0.025423f
C2995 VDDA.n546 GNDA 0.022299f
C2996 VDDA.n547 GNDA 0.022433f
C2997 VDDA.n548 GNDA 0.022433f
C2998 VDDA.n549 GNDA 0.022433f
C2999 VDDA.n550 GNDA 0.032471f
C3000 VDDA.n551 GNDA 0.013491f
C3001 VDDA.n552 GNDA 0.179785f
C3002 VDDA.t332 GNDA 0.190681f
C3003 VDDA.t220 GNDA 0.196129f
C3004 VDDA.t212 GNDA 0.196129f
C3005 VDDA.t95 GNDA 0.196129f
C3006 VDDA.t207 GNDA 0.196129f
C3007 VDDA.t125 GNDA 0.196129f
C3008 VDDA.t73 GNDA 0.196129f
C3009 VDDA.t216 GNDA 0.196129f
C3010 VDDA.t56 GNDA 0.196129f
C3011 VDDA.t127 GNDA 0.196129f
C3012 VDDA.t218 GNDA 0.196129f
C3013 VDDA.t418 GNDA 0.196129f
C3014 VDDA.t420 GNDA 0.196129f
C3015 VDDA.t65 GNDA 0.196129f
C3016 VDDA.t52 GNDA 0.196129f
C3017 VDDA.t70 GNDA 0.196129f
C3018 VDDA.t166 GNDA 0.196129f
C3019 VDDA.t299 GNDA 0.190681f
C3020 VDDA.n554 GNDA 0.012819f
C3021 VDDA.n555 GNDA 0.012819f
C3022 VDDA.n556 GNDA 0.022433f
C3023 VDDA.n557 GNDA 0.022299f
C3024 VDDA.n558 GNDA 0.022433f
C3025 VDDA.n559 GNDA 0.012819f
C3026 VDDA.n560 GNDA 0.022433f
C3027 VDDA.n561 GNDA 0.022433f
C3028 VDDA.n562 GNDA 0.022299f
C3029 VDDA.n563 GNDA 0.035425f
C3030 VDDA.n564 GNDA 0.010537f
C3031 VDDA.n565 GNDA 0.179785f
C3032 VDDA.n566 GNDA 0.012819f
C3033 VDDA.n567 GNDA 0.025423f
C3034 VDDA.t298 GNDA 0.091688f
C3035 VDDA.n568 GNDA 0.034243f
C3036 VDDA.n569 GNDA 0.050495f
C3037 VDDA.t347 GNDA 0.011836f
C3038 VDDA.n570 GNDA 0.025293f
C3039 VDDA.t346 GNDA 0.02245f
C3040 VDDA.t349 GNDA 0.02245f
C3041 VDDA.n571 GNDA 0.11168f
C3042 VDDA.t348 GNDA 0.077774f
C3043 VDDA.t23 GNDA 0.049353f
C3044 VDDA.t245 GNDA 0.049353f
C3045 VDDA.t345 GNDA 0.077774f
C3046 VDDA.n572 GNDA 0.11168f
C3047 VDDA.t344 GNDA 0.011836f
C3048 VDDA.n573 GNDA 0.025293f
C3049 VDDA.n574 GNDA 0.060838f
C3050 VDDA.n575 GNDA 0.015458f
C3051 VDDA.n576 GNDA 0.054277f
C3052 VDDA.n577 GNDA 0.126026f
C3053 VDDA.n578 GNDA 0.174064f
C3054 VDDA.n579 GNDA 0.015988f
C3055 VDDA.n580 GNDA 0.056438f
C3056 VDDA.t394 GNDA 0.023368f
C3057 VDDA.t321 GNDA 0.023368f
C3058 VDDA.t319 GNDA 0.012622f
C3059 VDDA.n581 GNDA 0.015959f
C3060 VDDA.n582 GNDA 0.056468f
C3061 VDDA.t404 GNDA 0.012622f
C3062 VDDA.n583 GNDA 0.015995f
C3063 VDDA.n584 GNDA 0.056432f
C3064 VDDA.t306 GNDA 0.02338f
C3065 VDDA.t385 GNDA 0.02338f
C3066 VDDA.t383 GNDA 0.012622f
C3067 VDDA.n585 GNDA 0.015995f
C3068 VDDA.n586 GNDA 0.077236f
C3069 VDDA.n587 GNDA 0.026808f
C3070 VDDA.n588 GNDA 0.066718f
C3071 VDDA.t384 GNDA 0.070312f
C3072 VDDA.t44 GNDA 0.049353f
C3073 VDDA.t430 GNDA 0.049353f
C3074 VDDA.t114 GNDA 0.049353f
C3075 VDDA.t82 GNDA 0.049353f
C3076 VDDA.t305 GNDA 0.070312f
C3077 VDDA.n589 GNDA 0.066718f
C3078 VDDA.t304 GNDA 0.013023f
C3079 VDDA.n590 GNDA 0.026361f
C3080 VDDA.n591 GNDA 0.038958f
C3081 VDDA.n592 GNDA 0.015959f
C3082 VDDA.n593 GNDA 0.056468f
C3083 VDDA.n594 GNDA 0.015959f
C3084 VDDA.n595 GNDA 0.056468f
C3085 VDDA.n596 GNDA 0.015959f
C3086 VDDA.n597 GNDA 0.056468f
C3087 VDDA.n598 GNDA 0.015959f
C3088 VDDA.n599 GNDA 0.056468f
C3089 VDDA.n600 GNDA 0.038958f
C3090 VDDA.n601 GNDA 0.024937f
C3091 VDDA.t406 GNDA 0.022404f
C3092 VDDA.n602 GNDA 0.068536f
C3093 VDDA.t405 GNDA 0.070492f
C3094 VDDA.t112 GNDA 0.049353f
C3095 VDDA.t110 GNDA 0.049353f
C3096 VDDA.t223 GNDA 0.049353f
C3097 VDDA.t442 GNDA 0.049353f
C3098 VDDA.t80 GNDA 0.049353f
C3099 VDDA.t60 GNDA 0.049353f
C3100 VDDA.t203 GNDA 0.049353f
C3101 VDDA.t199 GNDA 0.049353f
C3102 VDDA.t201 GNDA 0.049353f
C3103 VDDA.t444 GNDA 0.049353f
C3104 VDDA.t375 GNDA 0.070492f
C3105 VDDA.t376 GNDA 0.022404f
C3106 VDDA.n603 GNDA 0.068536f
C3107 VDDA.t374 GNDA 0.012622f
C3108 VDDA.n604 GNDA 0.024937f
C3109 VDDA.n605 GNDA 0.038958f
C3110 VDDA.n606 GNDA 0.015988f
C3111 VDDA.n607 GNDA 0.056438f
C3112 VDDA.n608 GNDA 0.038958f
C3113 VDDA.n609 GNDA 0.02596f
C3114 VDDA.n610 GNDA 0.06673f
C3115 VDDA.t320 GNDA 0.070312f
C3116 VDDA.t28 GNDA 0.049353f
C3117 VDDA.t448 GNDA 0.049353f
C3118 VDDA.t78 GNDA 0.049353f
C3119 VDDA.t10 GNDA 0.049353f
C3120 VDDA.t393 GNDA 0.070312f
C3121 VDDA.n611 GNDA 0.06673f
C3122 VDDA.t392 GNDA 0.012622f
C3123 VDDA.n612 GNDA 0.02596f
C3124 VDDA.n613 GNDA 0.129612f
C3125 VDDA.n614 GNDA 0.151316f
C3126 VDDA.n615 GNDA 0.721369f
C3127 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.015146f
C3128 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.015146f
C3129 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.048787f
C3130 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.015146f
C3131 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.015146f
C3132 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.048787f
C3133 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.268962f
C3134 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.015146f
C3135 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.015146f
C3136 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.045748f
C3137 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.814637f
C3138 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.053011f
C3139 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.053011f
C3140 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.18689f
C3141 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.074973f
C3142 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.074973f
C3143 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.074973f
C3144 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.074973f
C3145 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.086519f
C3146 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.070244f
C3147 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.043166f
C3148 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.043166f
C3149 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.040052f
C3150 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.074973f
C3151 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.074973f
C3152 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.074973f
C3153 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.074973f
C3154 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.086519f
C3155 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.070244f
C3156 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.043166f
C3157 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.043166f
C3158 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.040052f
C3159 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.042481f
C3160 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.074973f
C3161 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.074973f
C3162 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.074973f
C3163 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.074973f
C3164 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.086519f
C3165 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.070244f
C3166 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.043166f
C3167 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.043166f
C3168 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.040052f
C3169 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.074973f
C3170 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.074973f
C3171 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.074973f
C3172 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.074973f
C3173 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.086519f
C3174 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.070244f
C3175 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.043166f
C3176 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.043166f
C3177 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.040052f
C3178 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 0.044218f
C3179 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 1.21734f
C3180 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.091901f
C3181 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.319469f
C3182 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 0.946702f
C3183 bgr_0.VB3_CUR_BIAS GNDA 1.69501f
C3184 bgr_0.NFET_GATE_10uA.t0 GNDA 0.01496f
C3185 bgr_0.NFET_GATE_10uA.t3 GNDA 0.01496f
C3186 bgr_0.NFET_GATE_10uA.n0 GNDA 0.042091f
C3187 bgr_0.NFET_GATE_10uA.t18 GNDA 0.014586f
C3188 bgr_0.NFET_GATE_10uA.t6 GNDA 0.014586f
C3189 bgr_0.NFET_GATE_10uA.t14 GNDA 0.014586f
C3190 bgr_0.NFET_GATE_10uA.t19 GNDA 0.014586f
C3191 bgr_0.NFET_GATE_10uA.t5 GNDA 0.014586f
C3192 bgr_0.NFET_GATE_10uA.t13 GNDA 0.014586f
C3193 bgr_0.NFET_GATE_10uA.t12 GNDA 0.021563f
C3194 bgr_0.NFET_GATE_10uA.n1 GNDA 0.026685f
C3195 bgr_0.NFET_GATE_10uA.n2 GNDA 0.019075f
C3196 bgr_0.NFET_GATE_10uA.n3 GNDA 0.016149f
C3197 bgr_0.NFET_GATE_10uA.t15 GNDA 0.014586f
C3198 bgr_0.NFET_GATE_10uA.t8 GNDA 0.014586f
C3199 bgr_0.NFET_GATE_10uA.t21 GNDA 0.014586f
C3200 bgr_0.NFET_GATE_10uA.t16 GNDA 0.021563f
C3201 bgr_0.NFET_GATE_10uA.n4 GNDA 0.026685f
C3202 bgr_0.NFET_GATE_10uA.n5 GNDA 0.019075f
C3203 bgr_0.NFET_GATE_10uA.n6 GNDA 0.016149f
C3204 bgr_0.NFET_GATE_10uA.t20 GNDA 0.014586f
C3205 bgr_0.NFET_GATE_10uA.t7 GNDA 0.021563f
C3206 bgr_0.NFET_GATE_10uA.n7 GNDA 0.02376f
C3207 bgr_0.NFET_GATE_10uA.n8 GNDA 0.026114f
C3208 bgr_0.NFET_GATE_10uA.t11 GNDA 0.014586f
C3209 bgr_0.NFET_GATE_10uA.t22 GNDA 0.021563f
C3210 bgr_0.NFET_GATE_10uA.n9 GNDA 0.02376f
C3211 bgr_0.NFET_GATE_10uA.t9 GNDA 0.014586f
C3212 bgr_0.NFET_GATE_10uA.t17 GNDA 0.014586f
C3213 bgr_0.NFET_GATE_10uA.t23 GNDA 0.014586f
C3214 bgr_0.NFET_GATE_10uA.t10 GNDA 0.021563f
C3215 bgr_0.NFET_GATE_10uA.n10 GNDA 0.026685f
C3216 bgr_0.NFET_GATE_10uA.n11 GNDA 0.019075f
C3217 bgr_0.NFET_GATE_10uA.n12 GNDA 0.016149f
C3218 bgr_0.NFET_GATE_10uA.n13 GNDA 0.026114f
C3219 bgr_0.NFET_GATE_10uA.n14 GNDA 0.605807f
C3220 bgr_0.NFET_GATE_10uA.n15 GNDA 0.022264f
C3221 bgr_0.NFET_GATE_10uA.n16 GNDA 0.016149f
C3222 bgr_0.NFET_GATE_10uA.n17 GNDA 0.019075f
C3223 bgr_0.NFET_GATE_10uA.n18 GNDA 0.026685f
C3224 bgr_0.NFET_GATE_10uA.t2 GNDA 0.034164f
C3225 bgr_0.NFET_GATE_10uA.n19 GNDA 0.327308f
C3226 bgr_0.NFET_GATE_10uA.t4 GNDA 0.01496f
C3227 bgr_0.NFET_GATE_10uA.t1 GNDA 0.01496f
C3228 bgr_0.NFET_GATE_10uA.n20 GNDA 0.088541f
.ends

