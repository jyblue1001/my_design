** sch_path: /foss/designs/my_design/projects/pll/bandgapref/xschem_ngspice/test_inverter_speed.sch
**.subckt test_inverter_speed
XM1 osc2 osc GND GND sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 osc2 GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC2 net1 GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XC3 osc GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM2 osc2 osc VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 osc2 GND GND sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 osc2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 osc net1 GND GND sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 osc net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdd VDD GND pwl(0.0 1.8327163051845377 1e-12 1.827150722564271 2e-12 1.8876464291669526 3e-12 1.8202667600561389 4e-12 1.8127049038133833 5e-12 1.8198545732105111 6e-12 1.811375372220331 7e-12 1.7980088332918194 8e-12 1.6985618111425342 9e-12 1.8039984489818213 1e-11 1.8436861317641091 1.0999999999999999e-11 1.7242481449842257 1.2e-11 1.74465448117946 1.3e-11 1.779977046226712 1.4e-11 1.7654321474659338 1.5e-11 1.7457109778607447 1.6e-11 1.734077282159694 1.7e-11 1.8047726152800552 1.8e-11 1.7947853528159656 1.9e-11 1.880322241904439 2e-11 1.81520340985055 2.1e-11 1.797257058363057 2.1999999999999998e-11 1.8429975132421361 2.2999999999999998e-11 1.8129058639024833 2.4e-11 1.873786698609793 2.5e-11 1.8738382328660022 2.6e-11 1.7980182393626367 2.7e-11 1.794646553649616 2.8e-11 1.800480187092507 2.9e-11 1.8126723401508396 3e-11 1.8415158703042316 3.0999999999999996e-11 1.7860117694425384 3.2e-11 1.9183980760348054 3.3e-11 1.9146084384181121 3.4e-11 1.8085188476706282 3.5e-11 1.8030216766837042 3.6e-11 1.8218751124857824 3.7e-11 1.7994970598589757 3.8e-11 1.7619410749303062 3.9e-11 1.7716910702781905 4e-11 1.7617258662469193 4.1e-11 1.8035733451621732 4.2e-11 1.74288737654952 4.3e-11 1.7523137462652534 4.3999999999999997e-11 1.8019499239134829 4.5e-11 1.797432047520622 4.5999999999999996e-11 1.7794026875360538 4.7e-11 1.8296039029812214 4.8e-11 1.8290052193898894 4.9e-11 1.8660871233256664 5e-11 1.8453094698367798 5.1e-11 1.7736432107102071 5.2e-11 1.771398856588518 5.3e-11 1.7762419727765941 5.4e-11 1.7809855653489972 5.5e-11 1.8344639860810346 5.6e-11 1.7903709284055143 5.7e-11 1.7393791983651332 5.8e-11 1.8457352685251858 5.9e-11 1.8299948394126697 6e-11 1.7257636016843345 6.1e-11 1.8673062038010133 6.199999999999999e-11 1.762676761815815 6.3e-11 1.7952771188210894 6.4e-11 1.9344724663194366 6.5e-11 1.8251606735451913 6.6e-11 1.8070142198778365 6.7e-11 1.822581794950495 6.8e-11 1.8433577434055992 6.9e-11 1.8586440173766894 7e-11 1.7425359813992904 7.1e-11 1.908620640745165 7.2e-11 1.809265471687075 7.299999999999999e-11 1.844092011535034 7.4e-11 1.815814443978189 7.5e-11 1.8174549087939922 7.6e-11 1.8287526526198765 7.699999999999999e-11 1.8631080043146955 7.8e-11 1.8740262721701177 7.9e-11 1.8399547186028353 8e-11 1.8081440203655703 8.1e-11 1.7704822848666333 8.2e-11 1.8660169054545077 8.3e-11 1.7710966578621177 8.4e-11 1.7318553616796206 8.5e-11 1.875550956593855 8.6e-11 1.8543217730065096 8.7e-11 1.7397375772838228 8.799999999999999e-11 1.7790413917046584 8.9e-11 1.7138392857590918 9e-11 1.8094626979028263 9.1e-11 1.7758694168721911 9.199999999999999e-11 1.865294402245647 9.3e-11 1.8123795933580056 9.4e-11 1.8584406078309548 9.5e-11 1.8203795966909146 9.6e-11 1.8178487287873468 9.7e-11 1.840061141763086 9.8e-11 1.810236469328369 9.9e-11 1.834747653214371 1e-10 1.7666772180902084 1.01e-10 1.8087590761371912 1.02e-10 1.8563767022233388 1.0299999999999999e-10 1.8130697940285188 1.04e-10 1.6895555487883662 1.05e-10 1.8087338310604508 1.06e-10 1.7540745386880878 1.0699999999999999e-10 1.8675103460919664 1.08e-10 1.7738438132242673 1.09e-10 1.8584599146746883 1.1e-10 1.8529599305652158 1.1099999999999999e-10 1.8012818479235302 1.12e-10 1.7435015924492512 1.13e-10 1.8142981271385161 1.14e-10 1.8168733588171588 1.15e-10 1.736323185007797 1.16e-10 1.7698746000291739 1.17e-10 1.7043762614875524 1.18e-10 1.8490234073031433 1.19e-10 1.7893660424350661 1.2e-10 1.8299550896087775 1.21e-10 1.7682521891554293 1.22e-10 1.8249636686114266 1.23e-10 1.8035102004820962 1.2399999999999999e-10 1.8631913929211772 1.25e-10 1.8247753649882044 1.26e-10 1.729842720329594 1.27e-10 1.8474062857114282 1.28e-10 1.8980464136902777 1.29e-10 1.7756414755971017 1.3e-10 1.8602163851492055 1.3099999999999999e-10 1.839373040237761 1.32e-10 1.6919714693796637 1.33e-10 1.7587745979458784 1.34e-10 1.7772445295072739 1.35e-10 1.8194947604226803 1.36e-10 1.8214205989932994 1.37e-10 1.796676872737809 1.38e-10 1.6611047099965506 1.3899999999999999e-10 1.7753040942362022 1.4e-10 1.789923447186002 1.41e-10 1.852785759262784 1.42e-10 1.772254482917616 1.43e-10 1.8642870186214546 1.44e-10 1.9347324173058447 1.45e-10 1.7373192320136581 1.4599999999999999e-10 1.782007285700916 1.47e-10 1.7769120182112843 1.48e-10 1.7299175052672497 1.49e-10 1.8099256977227507 1.5e-10 1.81258345437525 1.51e-10 1.7175717443739735 1.52e-10 1.875958495052148 1.53e-10 1.7143257509104879 1.5399999999999999e-10 1.7554870717803346 1.55e-10 1.7114560908048528 1.56e-10 1.7785807150851236 1.57e-10 1.814927416852382 1.58e-10 1.920141092598495 1.59e-10 1.8318528243949899 1.6e-10 1.8928977903367257 1.6099999999999999e-10 1.7367926150394395 1.62e-10 1.8015987104376114 1.63e-10 1.831131476372892 1.64e-10 1.8110945830559895 1.65e-10 1.8274505911427714 1.66e-10 1.840632084390052 1.67e-10 1.7926623546669853 1.68e-10 1.7543338959632977 1.6899999999999999e-10 1.8112472279815335 1.7e-10 1.892847611496924 1.71e-10 1.8356475030886137 1.72e-10 1.8194375824388276 1.73e-10 1.8635047639391793 1.74e-10 1.8512658674280962 1.75e-10 1.739939426288583 1.7599999999999999e-10 1.7394318964443 1.77e-10 1.784372051580798 1.78e-10 1.7733712748329675 1.79e-10 1.7437075992682964 1.8e-10 1.7797065637555363 1.81e-10 1.775782669509666 1.82e-10 1.7674352393604331 1.83e-10 1.8320641689700579 1.8399999999999998e-10 1.7515451852029589 1.85e-10 1.7907335914133466 1.86e-10 1.7619570970322196 1.87e-10 1.7606457104889137 1.88e-10 1.767291897882778 1.89e-10 1.8308038749605262 1.9e-10 1.8060057668893026 1.9099999999999999e-10 1.8038307340594935 1.92e-10 1.7942232997201708 1.93e-10 1.7753041272411356 1.94e-10 1.8820891809039575 1.95e-10 1.736481815052756 1.96e-10 1.7839690857544812 1.97e-10 1.780820651883771 1.98e-10 1.7510035305165252 1.9899999999999998e-10 1.802346838405276 2e-10 1.790709793261867 2.01e-10 1.7810931910078376 2.02e-10 1.764024699612373 2.03e-10 1.8613974171287135 2.04e-10 1.7346341405753394 2.05e-10 1.7958649619438924 2.0599999999999999e-10 1.7930651016880403 2.0699999999999998e-10 1.7671243362540134 2.08e-10 1.7295170568155256 2.09e-10 1.8873202440666708 2.1e-10 1.8131174498940459 2.11e-10 1.7793823573439829 2.12e-10 1.7707309828575886 2.13e-10 1.8070857144790426 2.1399999999999998e-10 1.9103031465033133 2.15e-10 1.7520335621287375 2.16e-10 1.7495553351840465 2.17e-10 1.8792339142293186 2.18e-10 1.7873648389806545 2.19e-10 1.738971562048089 2.2e-10 1.7673587817321181 2.2099999999999999e-10 1.8359129265294811 2.2199999999999998e-10 1.7785325822148348 2.23e-10 1.8472501140719813 2.24e-10 1.7227493837506547 2.25e-10 1.80520149489594 2.26e-10 1.8550738359721042 2.27e-10 1.7788619433261934 2.28e-10 1.7809275320837539 2.2899999999999998e-10 1.8131550714963651 2.3e-10 1.8927200163280187 2.31e-10 1.8174313280437118 2.32e-10 1.7809101505568816 2.3299999999999997e-10 1.8438652865012009 2.34e-10 1.7352870719310767 2.35e-10 1.724461276433924 2.36e-10 1.8646636098479699 2.37e-10 1.724577243702446 2.38e-10 1.8643364131764497 2.39e-10 1.8793716611795215 2.4e-10 1.814649273202232 2.41e-10 1.8641452959260896 2.42e-10 1.8186258370160142 2.43e-10 1.7353990523265796 2.44e-10 1.8385102708004288 2.45e-10 1.8226079209882364 2.46e-10 1.8116134868681137 2.47e-10 1.7560684440252738 2.4799999999999997e-10 1.698745518195347 2.49e-10 1.8356789212116196 2.5e-10 1.873349046369865 2.51e-10 1.7855092411869902 2.52e-10 1.7284146395947466 2.53e-10 1.859024104315031 2.54e-10 1.8089708870459844 2.55e-10 1.8296133863256758 2.56e-10 1.7689105373547749 2.57e-10 1.7524662977463255 2.58e-10 1.8357262558721041 2.59e-10 1.8168405716747036 2.6e-10 1.869501670571628 2.61e-10 1.704914165125521 2.6199999999999997e-10 1.7242081384202792 2.6299999999999997e-10 1.8670133127728823 2.64e-10 1.723501923166897 2.65e-10 1.8150874661067185 2.66e-10 1.8923877218318341 2.67e-10 1.7489654202743217 2.68e-10 1.8381260620763389 2.69e-10 1.892944231201272 2.7e-10 1.8040969117366228 2.71e-10 1.7901917882218121 2.72e-10 1.8384620535472656 2.73e-10 1.8280530991865374 2.74e-10 1.7983780674303693 2.75e-10 1.8390920586298152 2.76e-10 1.9241346219269726 2.7699999999999997e-10 1.834940547731193 2.7799999999999997e-10 1.8360359084954947 2.79e-10 1.7735112917552498 2.8e-10 1.7608496394533457 2.81e-10 1.754972781584991 2.82e-10 1.78282596142972 2.83e-10 1.8104270312509942 2.84e-10 1.8357740297572214 2.85e-10 1.740709667793627 2.86e-10 1.6840868627708734 2.87e-10 1.8083184881754923 2.88e-10 1.7610959558789234 2.89e-10 1.8439445977971005 2.9e-10 1.782610089067769 2.91e-10 1.8620604992971905 2.9199999999999997e-10 1.7952068826409717 2.9299999999999997e-10 1.9477332379013066 2.94e-10 1.753457388738422 2.95e-10 1.8068204123977625 2.96e-10 1.773307131721585 2.97e-10 1.7685648812945667 2.98e-10 1.8546707952390522 2.99e-10 1.7257405371251675 3e-10 1.8988203653557014 3.01e-10 1.8200388150343114 3.02e-10 1.8820099979233094 3.03e-10 1.7296527251999512 3.04e-10 1.7938752338443889 3.05e-10 1.7763063372771595 3.06e-10 1.8216643439068592 3.0699999999999997e-10 1.7563903100987515 3.0799999999999997e-10 1.7668474801145486 3.09e-10 1.8364885944862954 3.1e-10 1.7579814281502697 3.11e-10 1.8398511064690457 3.12e-10 1.7835301518909021 3.13e-10 1.811704013326776 3.14e-10 1.8486673110723217 3.15e-10 1.7486833518282747 3.16e-10 1.8320573808321057 3.17e-10 1.9134720987863332 3.18e-10 1.8572132752075319 3.19e-10 1.7631667475342458 3.2e-10 1.795006729072496 3.21e-10 1.7845579333857007 3.2199999999999997e-10 1.7960236359322488 3.2299999999999997e-10 1.7829808631513566 3.24e-10 1.831407629204796 3.25e-10 1.8563554585453705 3.26e-10 1.700593223315943 3.27e-10 1.884505667281176 3.28e-10 1.7560276747581218 3.29e-10 1.88368404750047 3.3e-10 1.8641994131912827 3.31e-10 1.7722060553445471 3.32e-10 1.7466836186633004 3.33e-10 1.8154194563909472 3.34e-10 1.803668692204579 3.35e-10 1.9002857302240792 3.36e-10 1.7923129022928002 3.3699999999999997e-10 1.9471947066231405 3.3799999999999997e-10 1.8320028643202053 3.39e-10 1.8352222243536254 3.4e-10 1.8244011307238228 3.41e-10 1.7724897037472318 3.42e-10 1.7667339430834805 3.43e-10 1.7734681633752418 3.44e-10 1.8377575754498814 3.45e-10 1.7659442408673907 3.46e-10 1.8217388503548337 3.47e-10 1.7997890164417105 3.48e-10 1.8338911980521408 3.49e-10 1.7841707433738108 3.5e-10 1.8615548767092047 3.51e-10 1.7428581043966662 3.5199999999999997e-10 1.8331480010031411 3.5299999999999997e-10 1.807109481193172 3.54e-10 1.8206008397425344 3.55e-10 1.8041557573322764 3.56e-10 1.825492066676335 3.57e-10 1.7896191164442812 3.58e-10 1.7839017541963487 3.59e-10 1.8416279496865868 3.6e-10 1.7918204453036897 3.61e-10 1.7848263840531606 3.62e-10 1.8303478450903783 3.63e-10 1.849044806708202 3.64e-10 1.6682611899650235 3.65e-10 1.8556407080955277 3.66e-10 1.7320227958952024 3.6699999999999997e-10 1.7265963425003084 3.6799999999999997e-10 1.7165601567027915 3.69e-10 1.786014462448796 3.7e-10 1.777109222326703 3.71e-10 1.8714263257349597 3.72e-10 1.7501933900535693 3.73e-10 1.7566761995966051 3.74e-10 1.7879596334506376 3.75e-10 1.8119625098203347 3.76e-10 1.8508563759329681 3.77e-10 1.7761801911999764 3.78e-10 1.851257806510909 3.79e-10 1.8416360830088212 3.8e-10 1.697188274435075 3.81e-10 1.7437655195570514 3.8199999999999997e-10 1.818099583055236 3.8299999999999997e-10 1.7293408240742143 3.84e-10 1.8102787061938104 3.85e-10 1.7285085547259962 3.86e-10 1.7971177259192832 3.87e-10 1.751071015979872 3.88e-10 1.7257109465867175 3.89e-10 1.7533497913901763 3.9e-10 1.8938389385466667 3.91e-10 1.8086591607372908 3.92e-10 1.69508316190296 3.93e-10 1.8043552033250916 3.94e-10 1.8369296923052258 3.95e-10 1.8910064888880596 3.96e-10 1.7853143163078573 3.9699999999999997e-10 1.692284968738109 3.9799999999999997e-10 1.8365333901965408 3.9899999999999997e-10 1.8332999986095653 4e-10 1.815257311169251 4.01e-10 1.8079666627603568 4.02e-10 1.7370943374717904 4.03e-10 1.828333883395394 4.04e-10 1.861367527155647 4.05e-10 1.7819570981310726 4.06e-10 1.7525854148742044 4.07e-10 1.7346040493313455 4.08e-10 1.8098654903828404 4.09e-10 1.8838244558297705 4.1e-10 1.8356263295976258 4.11e-10 1.8354153957148325 4.1199999999999997e-10 1.835860458087831 4.1299999999999997e-10 1.7461385482198315 4.1399999999999997e-10 1.8143299836175721 4.15e-10 1.7768024346431 4.16e-10 1.8363485632345298 4.17e-10 1.7991204969758987 4.18e-10 1.7840041619902052 4.19e-10 1.8406721253244793 4.2e-10 1.7982867600832322 4.21e-10 1.8510778797325091 4.22e-10 1.7285390459621608 4.23e-10 1.7226596699613645 4.24e-10 1.8760901879359762 4.25e-10 1.8851881731024351 4.26e-10 1.7287553738728014 4.2699999999999997e-10 1.7888800960150364 4.2799999999999997e-10 1.7432209638220937 4.2899999999999997e-10 1.9234426572097303 4.3e-10 1.819920651739209 4.31e-10 1.8127877576206823 4.32e-10 1.87781549424925 4.33e-10 1.8435796815488958 4.34e-10 1.901606241201804 4.35e-10 1.700960152451053 4.36e-10 1.7177385852325247 4.37e-10 1.8463234112552593 4.38e-10 1.8622843634187132 4.39e-10 1.7484774771714369 4.4e-10 1.6772642161592974 4.41e-10 1.817621391495752 4.4199999999999997e-10 1.7827212774598984 4.4299999999999997e-10 1.8280403551113702 4.4399999999999997e-10 1.8174943454569108 4.45e-10 1.7924371536282844 4.46e-10 1.801220738448344 4.47e-10 1.8013644518004035 4.48e-10 1.7860431442457476 4.49e-10 1.8661011116481365 4.5e-10 1.8508099409228644 4.51e-10 1.7476207731585311 4.52e-10 1.9131268042883363 4.53e-10 1.7522149207588655 4.54e-10 1.7638899363544887 4.55e-10 1.8257668641898122 4.56e-10 1.7486189828413752 4.5699999999999997e-10 1.785248201213846 4.5799999999999997e-10 1.7698127595602964 4.5899999999999997e-10 1.7881559838870802 4.6e-10 1.821174480421877 4.61e-10 1.8209177614485175 4.62e-10 1.8032554690869873 4.63e-10 1.9184077853973227 4.64e-10 1.8620001107636455 4.65e-10 1.7774974327053032 4.659999999999999e-10 1.7069906854888008 4.67e-10 1.7562467763764518 4.68e-10 1.8696195057111453 4.69e-10 1.7991754969113731 4.7e-10 1.7441117406583981 4.71e-10 1.8344759543588263 4.72e-10 1.7970572775524805 4.73e-10 1.8172740842526325 4.74e-10 1.7852931049232206 4.75e-10 1.711773438289105 4.76e-10 1.798600426889991 4.77e-10 1.826698473233538 4.78e-10 1.815103656867173 4.79e-10 1.761401492711581 4.8e-10 1.7222499853998448 4.81e-10 1.7209806623698154 4.82e-10 1.8688608085205876 4.83e-10 1.7669048060832429 4.84e-10 1.9225069843479328 4.85e-10 1.6567666307541196 4.86e-10 1.7976397148880867 4.87e-10 1.8038959678870687 4.88e-10 1.740273498184448 4.89e-10 1.7238357021617088 4.9e-10 1.744736730991738 4.91e-10 1.8416528027836203 4.92e-10 1.7710054873761205 4.93e-10 1.8065382938328542 4.94e-10 1.8467351699390382 4.949999999999999e-10 1.7517406236619908 4.959999999999999e-10 1.8111626523422377 4.97e-10 1.8049952466339796 4.98e-10 1.8624713381600624 4.99e-10 1.756825322968963 5e-10 1.8230215066994424 5.01e-10 1.8047596773632115 5.02e-10 1.7691582383649247 5.03e-10 1.776527388433708 5.04e-10 1.8285584408807574 5.05e-10 1.878148174638425 5.06e-10 1.8716940109079903 5.07e-10 1.7140833118525667 5.08e-10 1.8934540728222315 5.09e-10 1.787869340274448 5.1e-10 1.7816223695262674 5.11e-10 1.7398388461778926 5.12e-10 1.9208628399944885 5.13e-10 1.7578018165496037 5.14e-10 1.8201931652239416 5.15e-10 1.782399372873001 5.16e-10 1.8492265548137337 5.17e-10 1.7690080947562488 5.18e-10 1.746356156592914 5.19e-10 1.8205821427636741 5.2e-10 1.7489023505862815 5.21e-10 1.8330610400551117 5.22e-10 1.8278356840858219 5.23e-10 1.7585835665273093 5.239999999999999e-10 1.7732646235737677 5.249999999999999e-10 1.7918912504038407 5.259999999999999e-10 1.8300253539630849 5.269999999999999e-10 1.825037426044296 5.28e-10 1.7519497888750004 5.29e-10 1.658958454623725 5.3e-10 1.784827987368962 5.31e-10 1.8196502450844019 5.32e-10 1.791747838826964 5.33e-10 1.8043995484581032 5.34e-10 1.8262817743241246 5.35e-10 1.8192746564071494 5.36e-10 1.850101480759782 5.37e-10 1.7596241195400775 5.38e-10 1.8209221903764246 5.39e-10 1.7416812264188861 5.4e-10 1.7566804021632088 5.41e-10 1.800619455327467 5.42e-10 1.7316134676787422 5.43e-10 1.8133152741519496 5.44e-10 1.7595159301935286 5.45e-10 1.829640273937183 5.46e-10 1.816673657934003 5.47e-10 1.8243128459951368 5.48e-10 1.7832834675470786 5.49e-10 1.7673523550592465 5.5e-10 1.855967411042847 5.51e-10 1.842431721061815 5.52e-10 1.8535822539789917 5.53e-10 1.8002718355940042 5.539999999999999e-10 1.7736578314713216 5.549999999999999e-10 1.8581225833191455 5.559999999999999e-10 1.8863335110115251 5.569999999999999e-10 1.8292718527321283 5.58e-10 1.8504306886704316 5.59e-10 1.907204015542831 5.6e-10 1.867644825370096 5.61e-10 1.7895691710705306 5.62e-10 1.7717031063028077 5.63e-10 1.8589659870895174 5.64e-10 1.7520608193764458 5.65e-10 1.7673046374896642 5.66e-10 1.8797024714756623 5.67e-10 1.8723881451528723 5.68e-10 1.7980278488489865 5.69e-10 1.7544440709774907 5.7e-10 1.7878388951825717 5.71e-10 1.8119002192863294 5.72e-10 1.8075343186780546 5.73e-10 1.7260182035556981 5.74e-10 1.8164512970298554 5.75e-10 1.7975973806434662 5.76e-10 1.7920731871350262 5.77e-10 1.7978182283950976 5.78e-10 1.7851366070920471 5.79e-10 1.8681694571070846 5.8e-10 1.6697517709348788 5.81e-10 1.8136886629817548 5.82e-10 1.818750526834614 5.83e-10 1.7303057059281757 5.839999999999999e-10 1.7964848555488024 5.849999999999999e-10 1.8944266154007154 5.859999999999999e-10 1.8249433803845476 5.869999999999999e-10 1.794861105980307 5.88e-10 1.8542432163031826 5.89e-10 1.7698398573180225 5.9e-10 1.7193215738045626 5.91e-10 1.8484999969116152 5.92e-10 1.8263555125679232 5.93e-10 1.824811953678718 5.94e-10 1.7804789333266877 5.95e-10 1.8742613025699866 5.96e-10 1.7739090804924966 5.97e-10 1.8988071266079334 5.98e-10 1.7191181936361077 5.99e-10 1.821636471950016 6e-10 1.810605525099203 6.01e-10 1.8230289736698655 6.02e-10 1.912455582492238 6.03e-10 1.8243995402060837 6.04e-10 1.7390175106251413 6.05e-10 1.831746642753366 6.06e-10 1.7000517346861064 6.07e-10 1.8960077436199678 6.08e-10 1.73392275983703 6.09e-10 1.8386824448234094 6.1e-10 1.7974328529846102 6.11e-10 1.8874225309537278 6.12e-10 1.7879857808223683 6.13e-10 1.8252529116892917 6.139999999999999e-10 1.8423393058129136 6.149999999999999e-10 1.8265160554194215 6.159999999999999e-10 1.7566400034211151 6.169999999999999e-10 1.815756611494019 6.18e-10 1.7400944866567067 6.19e-10 1.8476483662773153 6.2e-10 1.8276249310169597 6.21e-10 1.858207096323692 6.22e-10 1.7711697331352505 6.23e-10 1.8236849819127234 6.24e-10 1.813051420383545 6.25e-10 1.82422339530917 6.26e-10 1.818728383774115 6.27e-10 1.7868399442086642 6.28e-10 1.8092576203328024 6.29e-10 1.818233442776927 6.3e-10 1.75352769083795 6.31e-10 1.7923180014004991 6.32e-10 1.7858402393270185 6.33e-10 1.8075951502652283 6.34e-10 1.7154711290647897 6.35e-10 1.8959510328864009 6.36e-10 1.793366461235506 6.37e-10 1.8134112203475095 6.38e-10 1.8439766248030367 6.39e-10 1.8231321471842703 6.4e-10 1.8429297466303034 6.41e-10 1.8119094852500677 6.42e-10 1.9533099454171206 6.43e-10 1.7773958929110782 6.439999999999999e-10 1.8162176925931017 6.449999999999999e-10 1.75217577456288 6.459999999999999e-10 1.7806488310237032 6.469999999999999e-10 1.7968078486250587 6.48e-10 1.824250046206668 6.49e-10 1.7810431101840465 6.5e-10 1.800580708604623 6.51e-10 1.8548258632565462 6.52e-10 1.821125233247144 6.53e-10 1.745311416938016 6.54e-10 1.8066166528530068 6.55e-10 1.8085981864666556 6.56e-10 1.7893678836424871 6.57e-10 1.8228367479391836 6.58e-10 1.8207967870317812 6.59e-10 1.8449281209449302 6.6e-10 1.7174613353639259 6.61e-10 1.86460271783021 6.62e-10 1.7460459959721701 6.63e-10 1.7982341858172528 6.64e-10 1.802965257523087 6.65e-10 1.7867678346313938 6.66e-10 1.7968733978233224 6.67e-10 1.8307795866537817 6.68e-10 1.8022546775632373 6.69e-10 1.862757137280307 6.7e-10 1.7739424390892082 6.71e-10 1.8188128756113326 6.72e-10 1.8174509014530535 6.73e-10 1.8007479537270499 6.739999999999999e-10 1.785063822450471 6.749999999999999e-10 1.8582879183429295 6.759999999999999e-10 1.8334257911408223 6.769999999999999e-10 1.8270179358115854 6.78e-10 1.7568333538112304 6.79e-10 1.9242127701720535 6.8e-10 1.8132323437034235 6.81e-10 1.770007361169011 6.82e-10 1.7916846783220268 6.83e-10 1.8352443153367546 6.84e-10 1.7920834028383197 6.85e-10 1.7370376385959787 6.86e-10 1.7683310464874726 6.87e-10 1.8623679149205443 6.88e-10 1.8590608004884486 6.89e-10 1.788174206927317 6.9e-10 1.8741859109219101 6.91e-10 1.8103223816545033 6.92e-10 1.8234041569382933 6.93e-10 1.8606673862276464 6.94e-10 1.786019157921935 6.95e-10 1.7661121323875908 6.96e-10 1.8400603474720265 6.97e-10 1.8000420915759696 6.98e-10 1.7719019936285225 6.99e-10 1.712073491366161 7e-10 1.8366475056838294 7.01e-10 1.7959497247569407 7.02e-10 1.8428514905576274 7.03e-10 1.872516242374966 7.039999999999999e-10 1.8605718857967617 7.049999999999999e-10 1.7948308141336535 7.059999999999999e-10 1.7661481097471858 7.069999999999999e-10 1.74365532336692 7.08e-10 1.7205625251236287 7.09e-10 1.759651547327707 7.1e-10 1.8236611046690991 7.11e-10 1.8324704191193772 7.12e-10 1.8434610077593012 7.13e-10 1.8640864757364655 7.14e-10 1.7295286419458944 7.15e-10 1.769698297998667 7.16e-10 1.8247180562692784 7.17e-10 1.8187227468522231 7.18e-10 1.8206584946712643 7.19e-10 1.8365686171273803 7.2e-10 1.8052250276263226 7.21e-10 1.7337699135041067 7.22e-10 1.8644204671611961 7.23e-10 1.7855670918743063 7.24e-10 1.749743167213522 7.25e-10 1.8335813556985625 7.26e-10 1.7984286081015863 7.27e-10 1.7931734385635292 7.28e-10 1.8760828776514678 7.29e-10 1.6839716307910235 7.3e-10 1.7360615718734576 7.31e-10 1.7946367652942796 7.32e-10 1.811867312712953 7.33e-10 1.7916360136612055 7.339999999999999e-10 1.7971393992028963 7.349999999999999e-10 1.8389979352827506 7.359999999999999e-10 1.7687920793574998 7.369999999999999e-10 1.783670100866354 7.38e-10 1.8884203457086493 7.39e-10 1.7978171815850694 7.4e-10 1.8548711645868108 7.41e-10 1.7930575129336868 7.42e-10 1.8281913323495569 7.43e-10 1.7846863802972124 7.44e-10 1.7464589178018726 7.45e-10 1.8234037831026242 7.46e-10 1.797251717825056 7.47e-10 1.7235837497885498 7.48e-10 1.7523216731660756 7.49e-10 1.8057420480752815 7.5e-10 1.846613504674974 7.51e-10 1.811860029804209 7.52e-10 1.6892734053883174 7.53e-10 1.8925185660521109 7.54e-10 1.7994583271502749 7.55e-10 1.8436887586554327 7.56e-10 1.7591101254097907 7.57e-10 1.7805637152974871 7.58e-10 1.7795657653432186 7.59e-10 1.7740374555529117 7.6e-10 1.7857571403054757 7.61e-10 1.8596668012361803 7.62e-10 1.7899490606373392 7.63e-10 1.8004902087130037 7.639999999999999e-10 1.7964105633456198 7.649999999999999e-10 1.8250007974241318 7.659999999999999e-10 1.7635483228511701 7.669999999999999e-10 1.7990850918641164 7.68e-10 1.8648654512713216 7.69e-10 1.802233893862316 7.7e-10 1.6722897402715025 7.71e-10 1.790759216893517 7.72e-10 1.8709710391443508 7.73e-10 1.8152992653394886 7.74e-10 1.833051773879549 7.75e-10 1.7403377794195354 7.76e-10 1.7259660010501063 7.77e-10 1.8346228622079699 7.78e-10 1.8493144863191515 7.79e-10 1.7927757606793253 7.8e-10 1.812907952665399 7.81e-10 1.7250011942687657 7.82e-10 1.7713184108905535 7.83e-10 1.762834707685918 7.84e-10 1.8318748395790645 7.85e-10 1.9339138683788997 7.86e-10 1.8346485609350764 7.87e-10 1.8447022800962098 7.88e-10 1.8020114600973451 7.89e-10 1.8243385368687246 7.9e-10 1.7853428614225957 7.91e-10 1.8510898260006554 7.92e-10 1.784661880930487 7.93e-10 1.82549693058064 7.939999999999999e-10 1.8723128095596708 7.949999999999999e-10 1.8221048745781152 7.959999999999999e-10 1.8620365630330349 7.969999999999999e-10 1.7833027350082733 7.979999999999999e-10 1.8118069666968888 7.99e-10 1.8587396347991365 8e-10 1.7841709936672114 8.01e-10 1.9131806144636598 8.02e-10 1.7505408712398687 8.03e-10 1.782199301346752 8.04e-10 1.850046744173317 8.05e-10 1.9181098637299647 8.06e-10 1.814784504973343 8.07e-10 1.7746263894216463 8.08e-10 1.75218104201 8.09e-10 1.7889384011906453 8.1e-10 1.8360870410662768 8.11e-10 1.7900627777368132 8.12e-10 1.8272200417613464 8.13e-10 1.7929465640711988 8.14e-10 1.7919983130975239 8.15e-10 1.752974627690929 8.16e-10 1.7594834511540691 8.17e-10 1.7597674121316627 8.18e-10 1.7596366227258455 8.19e-10 1.7795650758694423 8.2e-10 1.8109901525360426 8.21e-10 1.785978587335922 8.22e-10 1.8748426864790013 8.23e-10 1.8078894971675943 8.239999999999999e-10 1.8019546588833577 8.249999999999999e-10 1.6992430980299866 8.259999999999999e-10 1.7562782123018028 8.269999999999999e-10 1.8199732341796022 8.279999999999999e-10 1.860756901564059 8.29e-10 1.7917952435550133 8.3e-10 1.848605542992006 8.31e-10 1.7567519498814677 8.32e-10 1.8353714753319588 8.33e-10 1.8182853354159447 8.34e-10 1.8418037300048664 8.35e-10 1.7577661835041734 8.36e-10 1.7001377148108776 8.37e-10 1.7601630924638396 8.38e-10 1.8070846291783769 8.39e-10 1.7224890933540478 8.4e-10 1.784297514566162 8.41e-10 1.8767380380985081 8.42e-10 1.8150806958946841 8.43e-10 1.8011219580826732 8.44e-10 1.7203647062106653 8.45e-10 1.7418179916220722 8.46e-10 1.7433501661200221 8.47e-10 1.7432519540294225 8.48e-10 1.8591273862928763 8.49e-10 1.7700511360055853 8.5e-10 1.7703663896115938 8.51e-10 1.769125782205116 8.52e-10 1.8217211612542061 8.53e-10 1.7245347415777093 8.539999999999999e-10 1.798379891964522 8.549999999999999e-10 1.6836275550319135 8.559999999999999e-10 1.8530819789480315 8.569999999999999e-10 1.7379419804849534 8.579999999999999e-10 1.7375099159982266 8.59e-10 1.7898973491726056 8.6e-10 1.7811357943937307 8.61e-10 1.7581252092590578 8.62e-10 1.791652377738449 8.63e-10 1.8097140698120735 8.64e-10 1.8858063445069522 8.65e-10 1.8063151540077766 8.66e-10 1.830147813065551 8.67e-10 1.8057998060574816 8.68e-10 1.8418735698182511 8.69e-10 1.7544348621473154 8.7e-10 1.7823387148753738 8.71e-10 1.678175300185211 8.72e-10 1.8258348100599173 8.73e-10 1.8135190690903094 8.74e-10 1.8150146962124287 8.75e-10 1.764481559988479 8.76e-10 1.7454780247836157 8.77e-10 1.792284604867153 8.78e-10 1.7692004168703577 8.79e-10 1.851796009838188 8.8e-10 1.8187067312602472 8.81e-10 1.7641183675521557 8.82e-10 1.8631466349470955 8.83e-10 1.7776852932530751 8.839999999999999e-10 1.7901437984645716 8.849999999999999e-10 1.8399639347855168 8.859999999999999e-10 1.7908891962474605 8.869999999999999e-10 1.8010105782948063 8.879999999999999e-10 1.7918552425728702 8.89e-10 1.765447093017369 8.9e-10 1.7509180086592075 8.91e-10 1.8756888804393925 8.92e-10 1.754168020689471 8.93e-10 1.829895777662181 8.94e-10 1.811907832827598 8.95e-10 1.6726762944696978 8.96e-10 1.7457617791632007 8.97e-10 1.8258630800572744 8.98e-10 1.7921440432881328 8.99e-10 1.801590430041287 9e-10 1.8070453936926343 9.01e-10 1.7529747711153165 9.02e-10 1.8092441011412674 9.03e-10 1.7336168822487004 9.04e-10 1.8677764112567559 9.05e-10 1.7777593800456402 9.06e-10 1.893690189911193 9.07e-10 1.836376805068381 9.08e-10 1.8198774489008984 9.09e-10 1.8327731312237616 9.1e-10 1.8477232657861382 9.11e-10 1.790186774269682 9.12e-10 1.7473540131702119 9.13e-10 1.7799986076720848 9.139999999999999e-10 1.8055079183349747 9.149999999999999e-10 1.7295124054978688 9.159999999999999e-10 1.7477266284787685 9.169999999999999e-10 1.7834091218976642 9.179999999999999e-10 1.8922080608794534 9.19e-10 1.7384788128187953 9.2e-10 1.8707254109008722 9.21e-10 1.7919668283031653 9.22e-10 1.7968803876171973 9.23e-10 1.8068271538451122 9.24e-10 1.793063502124037 9.25e-10 1.7670360951473387 9.26e-10 1.8873737882129125 9.27e-10 1.7921919762515865 9.28e-10 1.8294340147593202 9.29e-10 1.850236557846241 9.3e-10 1.7632986753181912 9.31e-10 1.7472956968168327 9.319999999999999e-10 1.806390181049123 9.33e-10 1.7853187151395276 9.34e-10 1.9024772000922066 9.35e-10 1.7375303652664222 9.36e-10 1.7794732482279492 9.37e-10 1.8117073264709025 9.38e-10 1.8652355056069247 9.39e-10 1.846170735995214 9.4e-10 1.8863047168622653 9.41e-10 1.7878229085249477 9.42e-10 1.79096248162636 9.43e-10 1.8197121474978768 9.44e-10 1.8195723387891394 9.45e-10 1.8127146431083971 9.46e-10 1.6623369568141189 9.47e-10 1.900305188879959 9.48e-10 1.7976251448282183 9.49e-10 1.7562591224851525 9.5e-10 1.7742370736652362 9.51e-10 1.7750538338566546 9.52e-10 1.7875627047656126 9.53e-10 1.8619167220371267 9.54e-10 1.8047847315173406 9.55e-10 1.8263720693496142 9.56e-10 1.8040925111110278 9.57e-10 1.859819151513112 9.58e-10 1.7850153228049692 9.589999999999999e-10 1.7948334638906787 9.6e-10 1.6717160386607328 9.609999999999999e-10 1.8434850811826677 9.62e-10 1.7367087774707384 9.629999999999999e-10 1.7872332280177865 9.64e-10 1.8217623955848858 9.65e-10 1.7678940052253669 9.66e-10 1.7308484392785115 9.67e-10 1.8759407158620387 9.68e-10 1.77803358313981 9.69e-10 1.7709803104497477 9.7e-10 1.794724149276826 9.71e-10 1.761325261399729 9.72e-10 1.828053030762344 9.73e-10 1.778153855847143 9.74e-10 1.781611390736185 9.75e-10 1.7733100619094353 9.76e-10 1.798373614273015 9.77e-10 1.803669997105389 9.78e-10 1.776839879375547 9.79e-10 1.8183696344664826 9.8e-10 1.8487037887224094 9.81e-10 1.7636801047000172 9.82e-10 1.8175832541878707 9.83e-10 1.829455644904446 9.84e-10 1.7786785030182906 9.85e-10 1.7805657053754744 9.86e-10 1.825058180598205 9.87e-10 1.7731402844990618 9.88e-10 1.7531113839367622 9.89e-10 1.904470847489502 9.899999999999999e-10 1.887249892742456 9.91e-10 1.895091283144411 9.919999999999999e-10 1.789897782398459 9.93e-10 1.847641852554629 9.94e-10 1.7202389943290006 9.95e-10 1.8650321301439403 9.96e-10 1.8049151335697164 9.97e-10 1.7192417348562263 9.98e-10 1.8421787562099765 9.99e-10 1.747012443705723 1e-09 1.8307916677895917 1.001e-09 1.8732391450409176 1.002e-09 1.773605648436234 1.003e-09 1.8306974983381126 1.004e-09 1.8052731445585808 1.005e-09 1.8114284166524428 1.006e-09 1.7573035437570868 1.007e-09 1.7928436982801128 1.008e-09 1.8957763053249386 1.009e-09 1.8205497236278276 1.01e-09 1.8544019206596778 1.011e-09 1.7042502990064174 1.012e-09 1.7665641201505424 1.013e-09 1.8472377485970752 1.014e-09 1.7818840903173851 1.015e-09 1.8076864505974983 1.016e-09 1.756231484497302 1.017e-09 1.770716217356349 1.018e-09 1.7428312737560143 1.0189999999999999e-09 1.7389466162950689 1.02e-09 1.8181090968500968 1.0209999999999999e-09 1.7193420887791637 1.022e-09 1.8678941634267048 1.0229999999999999e-09 1.7202163776977981 1.024e-09 1.7380114821998365 1.025e-09 1.7652594106792674 1.026e-09 1.7785658184193145 1.027e-09 1.8421385644367119 1.028e-09 1.8953146397234306 1.029e-09 1.793209307305873 1.03e-09 1.7601217771924824 1.031e-09 1.87361853102333 1.032e-09 1.787731373622 1.033e-09 1.8607367351573707 1.034e-09 1.866299572172361 1.035e-09 1.7793260367855694 1.036e-09 1.759329524691219 1.037e-09 1.7848101621709407 1.038e-09 1.8370878831906974 1.039e-09 1.7921149526739006 1.04e-09 1.774430510090326 1.041e-09 1.8271559737885121 1.042e-09 1.7706236456445168 1.043e-09 1.774652322480455 1.044e-09 1.825010673579877 1.045e-09 1.7206610191717606 1.046e-09 1.7957731383428255 1.047e-09 1.7682468087336511 1.0479999999999999e-09 1.746790064618665 1.049e-09 1.778772733987166 1.0499999999999999e-09 1.8151265637883438 1.051e-09 1.8013537784384916 1.0519999999999999e-09 1.856313612619457 1.053e-09 1.8451474883177252 1.0539999999999999e-09 1.7806056888907302 1.055e-09 1.8039728129020947 1.056e-09 1.792626322477244 1.057e-09 1.7396442378245998 1.058e-09 1.855352660283471 1.059e-09 1.848683732279594 1.06e-09 1.8236110207704395 1.061e-09 1.8335145803470152 1.062e-09 1.7900518307637907 1.063e-09 1.7806196884728203 1.064e-09 1.7605010813778135 1.065e-09 1.730895596854859 1.066e-09 1.782853391904774 1.067e-09 1.797300553513528 1.068e-09 1.810643288537534 1.069e-09 1.8267778926449867 1.07e-09 1.8142733756248146 1.071e-09 1.77041443675756 1.072e-09 1.6163787181909715 1.073e-09 1.7987961838530422 1.074e-09 1.7726933711684798 1.075e-09 1.8109699862702884 1.076e-09 1.7012167264226257 1.077e-09 1.8493982411172174 1.078e-09 1.8006088612368427 1.0789999999999999e-09 1.808286329873655 1.08e-09 1.828556819073419 1.0809999999999999e-09 1.770387476460522 1.082e-09 1.81772703963025 1.0829999999999999e-09 1.860302404996583 1.084e-09 1.7400575961201579 1.085e-09 1.871507221626871 1.086e-09 1.7441897124758727 1.087e-09 1.8084570794540569 1.088e-09 1.7999077236417211 1.089e-09 1.8260393418920124 1.09e-09 1.7785239613769888 1.091e-09 1.8231856791663446 1.092e-09 1.7427504199236528 1.093e-09 1.905952863032093 1.094e-09 1.7771383802868401 1.095e-09 1.6775983677162927 1.096e-09 1.8003294595359596 1.097e-09 1.7539977097348958 1.098e-09 1.7459189778331325 1.099e-09 1.8125301152264142 1.1e-09 1.8350062857529095 1.101e-09 1.7226020709079726 1.102e-09 1.8420855889765186 1.103e-09 1.7006517298305193 1.104e-09 1.8061692712286752 1.105e-09 1.8408684027924378 1.106e-09 1.8093912528538099 1.107e-09 1.7487511745791433 1.1079999999999999e-09 1.752693423544563 1.109e-09 1.7822399819872747 1.1099999999999999e-09 1.846499342814817 1.111e-09 1.7043333507061296 1.1119999999999999e-09 1.7394353613609939 1.113e-09 1.894944635320011 1.1139999999999999e-09 1.8416078303245882 1.115e-09 1.81683951751422 1.116e-09 1.8426367806606443 1.117e-09 1.835256703741222 1.118e-09 1.726527422663427 1.119e-09 1.8642935290425964 1.12e-09 1.8054364089664166 1.121e-09 1.7781600386134702 1.122e-09 1.7956118154713652 1.123e-09 1.8406771423690038 1.124e-09 1.7670945925239647 1.125e-09 1.8068705909376428 1.126e-09 1.808529097222773 1.127e-09 1.814690803190746 1.128e-09 1.7955992187548717 1.129e-09 1.8639907152870945 1.13e-09 1.889226890670328 1.131e-09 1.7676986813516193 1.132e-09 1.7767428370689018 1.133e-09 1.7918661344485867 1.134e-09 1.8244366952794808 1.135e-09 1.8291183771870994 1.136e-09 1.8099615848485864 1.137e-09 1.8580861396328319 1.138e-09 1.8260994130986041 1.1389999999999999e-09 1.8138837710119475 1.14e-09 1.8512215169745698 1.1409999999999999e-09 1.8903600916238752 1.142e-09 1.754563081488777 1.1429999999999999e-09 1.7628083597381352 1.144e-09 1.8266732840414182 1.145e-09 1.8093739505874833 1.146e-09 1.7869054398133837 1.147e-09 1.8657569498533015 1.148e-09 1.805504055510069 1.149e-09 1.7309632768008525 1.15e-09 1.8002638688274069 1.151e-09 1.825407783877815 1.152e-09 1.874094638100059 1.153e-09 1.7722373497110744 1.154e-09 1.7701524905912047 1.155e-09 1.7237302241715038 1.156e-09 1.9127116894731213 1.157e-09 1.8134956215208273 1.158e-09 1.7848328623676892 1.159e-09 1.771806599980849 1.16e-09 1.801963314698213 1.161e-09 1.9302890529761851 1.162e-09 1.8787136702736111 1.163e-09 1.7889506571147427 1.164e-09 1.8510296937261987 1.165e-09 1.8445147232031411 1.166e-09 1.8079619559055204 1.167e-09 1.81912357842595 1.1679999999999999e-09 1.780158243553111 1.169e-09 1.7674330905981952 1.1699999999999999e-09 1.8545573858426745 1.171e-09 1.7794187978172162 1.1719999999999999e-09 1.8163423361846613 1.173e-09 1.831849254217131 1.1739999999999999e-09 1.869905023932512 1.175e-09 1.924306308377335 1.176e-09 1.8017218526564425 1.177e-09 1.8401142410939364 1.178e-09 1.8225194988210294 1.179e-09 1.6918884423686655 1.18e-09 1.7588780829659019 1.181e-09 1.7635219628661005 1.182e-09 1.8409439974685236 1.183e-09 1.8273795333136216 1.184e-09 1.7782928500118256 1.185e-09 1.9055368994089286 1.186e-09 1.8611336628111574 1.187e-09 1.8105285102396547 1.188e-09 1.8315517737517129 1.189e-09 1.8379038009255761 1.19e-09 1.8143143741442602 1.191e-09 1.9277951566858063 1.192e-09 1.800959907100053 1.193e-09 1.7395190054555465 1.194e-09 1.8245662182401852 1.195e-09 1.856660550324694 1.196e-09 1.796581371392587 1.197e-09 1.7592033685624031 1.198e-09 1.809804220861666 1.1989999999999999e-09 1.7575652480138817 1.2e-09 1.8047414882765604 1.2009999999999999e-09 1.7679461141864146 1.202e-09 1.800847971401337 1.2029999999999999e-09 1.7618626214906028 1.204e-09 1.7549666415104326 1.205e-09 1.7650068516329693 1.206e-09 1.711050469408307 1.207e-09 1.7757098815347383 1.208e-09 1.7885537824176347 1.209e-09 1.773410611782208 1.21e-09 1.8466566381166925 1.211e-09 1.7957744381263108 1.212e-09 1.8164730029556375 1.213e-09 1.904794255200924 1.214e-09 1.800585986717807 1.215e-09 1.7146263805300097 1.216e-09 1.8258715066388116 1.217e-09 1.8257934326118699 1.218e-09 1.786317751968894 1.219e-09 1.8598486288237048 1.22e-09 1.8074504839201115 1.221e-09 1.7966373253842893 1.222e-09 1.6833448859609463 1.223e-09 1.7568889994500125 1.224e-09 1.7875612540167818 1.225e-09 1.7777654302509929 1.226e-09 1.7885089068973967 1.227e-09 1.8237110509672816 1.2279999999999999e-09 1.805560993328292 1.229e-09 1.7931815873892052 1.2299999999999999e-09 1.811166711441565 1.231e-09 1.8278429934347404 1.2319999999999999e-09 1.848404136021536 1.233e-09 1.8401088950812043 1.2339999999999999e-09 1.754137090175088 1.235e-09 1.8569821317338004 1.236e-09 1.800873584882028 1.237e-09 1.837156744635742 1.238e-09 1.74943857433845 1.239e-09 1.845086962204781 1.24e-09 1.8501388273746693 1.241e-09 1.828171948853973 1.242e-09 1.771698325667288 1.243e-09 1.803109259961004 1.244e-09 1.7568996451752257 1.245e-09 1.7938895188296662 1.246e-09 1.7374329395524684 1.247e-09 1.8190048016454963 1.248e-09 1.8038300762395076 1.249e-09 1.8351053071855956 1.25e-09 1.9362935974763764 1.251e-09 1.8322846107303972 1.252e-09 1.851908037091428 1.253e-09 1.7518454400034997 1.254e-09 1.8396801856801337 1.255e-09 1.7853368573541657 1.256e-09 1.7994843296152447 1.257e-09 1.8355527999893855 1.258e-09 1.8173783420459846 1.2589999999999999e-09 1.7451359926731782 1.26e-09 1.7595897142935342 1.2609999999999999e-09 1.813572272773716 1.262e-09 1.7779480325190165 1.2629999999999999e-09 1.7879974159963576 1.264e-09 1.7542989075444282 1.265e-09 1.7190735354199367 1.266e-09 1.80755844633075 1.267e-09 1.8949797745682886 1.268e-09 1.850405568191556 1.269e-09 1.7350034142666702 1.27e-09 1.8172473394353643 1.271e-09 1.7449572129681628 1.272e-09 1.8345568380636275 1.273e-09 1.791685901977166 1.274e-09 1.7660989969531031 1.275e-09 1.7325653454849608 1.276e-09 1.7914119816197445 1.277e-09 1.9206918437509912 1.278e-09 1.714149614587122 1.279e-09 1.8145209378743379 1.28e-09 1.7495071000598708 1.281e-09 1.8340754698075872 1.282e-09 1.7621837499994035 1.283e-09 1.7307353555805027 1.284e-09 1.6815868194019923 1.285e-09 1.8681214500816878 1.286e-09 1.7758025225133685 1.287e-09 1.7929611692077283 1.2879999999999999e-09 1.7836909270069126 1.289e-09 1.839577492198185 1.2899999999999999e-09 1.7564033823455876 1.291e-09 1.79166049032974 1.2919999999999999e-09 1.7973135941286533 1.293e-09 1.7682449653986543 1.2939999999999999e-09 1.8339599494280396 1.295e-09 1.7597987330173 1.296e-09 1.7358033138069835 1.297e-09 1.812090848014868 1.298e-09 1.741269091432389 1.299e-09 1.7606107002845843 1.3e-09 1.787386855657799 1.301e-09 1.829499649684573 1.302e-09 1.7948194051347042 1.303e-09 1.8121732485674862 1.304e-09 1.730289554248866 1.305e-09 1.838032170385866 1.306e-09 1.7827162555962357 1.307e-09 1.8471226820648345 1.308e-09 1.8831064446672776 1.309e-09 1.7306142246456628 1.31e-09 1.8054040099980664 1.311e-09 1.7663091506490087 1.312e-09 1.8928509531586544 1.313e-09 1.8291761136491622 1.314e-09 1.7282993741749924 1.315e-09 1.7857402138824676 1.316e-09 1.7489594328960185 1.317e-09 1.7845436285090757 1.318e-09 1.7326593462406426 1.3189999999999999e-09 1.8107164013801909 1.32e-09 1.8108797574284257 1.3209999999999999e-09 1.8514336849449706 1.322e-09 1.7609327540201831 1.3229999999999999e-09 1.769177057281653 1.324e-09 1.7942815908746232 1.3249999999999999e-09 1.930642451302282 1.326e-09 1.8724336062997504 1.327e-09 1.7065058876528507 1.328e-09 1.7561741643742703 1.329e-09 1.7234817482593896 1.33e-09 1.7698621405495285 1.331e-09 1.8980453667039612 1.332e-09 1.825891641398717 1.333e-09 1.8293340953207342 1.334e-09 1.7892497392071771 1.335e-09 1.8260102527517308 1.336e-09 1.795372188639134 1.337e-09 1.809362792128254 1.338e-09 1.892679203247137 1.339e-09 1.8730787212990938 1.34e-09 1.8097481819165175 1.341e-09 1.8379120158974642 1.342e-09 1.8373954655981983 1.343e-09 1.7217437819913641 1.344e-09 1.8302526716112473 1.345e-09 1.846966539523164 1.346e-09 1.7781298979311184 1.347e-09 1.8183861011475981 1.3479999999999999e-09 1.7393233669910384 1.349e-09 1.7656424171195229 1.3499999999999999e-09 1.7110051786327078 1.351e-09 1.8506611856544586 1.3519999999999999e-09 1.7880959935381908 1.353e-09 1.8939776163986648 1.3539999999999999e-09 1.8081034897032848 1.355e-09 1.7739557537714148 1.356e-09 1.8024061668966749 1.357e-09 1.7082227149060107 1.358e-09 1.8158788762868894 1.359e-09 1.7977813209311164 1.36e-09 1.8289313398692013 1.361e-09 1.7865567057672946 1.362e-09 1.893970048569892 1.363e-09 1.8328019348662283 1.364e-09 1.7930936159891282 1.365e-09 1.7599031002030874 1.366e-09 1.7983874378195515 1.367e-09 1.7910185229182358 1.368e-09 1.8472871381097011 1.369e-09 1.7630826368795174 1.37e-09 1.7049285281049864 1.371e-09 1.8284648551815685 1.372e-09 1.8870849723632364 1.373e-09 1.7770931883903405 1.374e-09 1.750412283998057 1.375e-09 1.80637457458647 1.376e-09 1.7690535143009074 1.377e-09 1.7929206634578474 1.378e-09 1.7047232605548812 1.3789999999999999e-09 1.8232968751576575 1.38e-09 1.7887877651379833 1.3809999999999999e-09 1.8002215620873914 1.382e-09 1.84025124689582 1.3829999999999999e-09 1.767153740767128 1.384e-09 1.7766825855841029 1.3849999999999999e-09 1.77540684855075 1.386e-09 1.8050918215543084 1.387e-09 1.7298516591114876 1.388e-09 1.7470760413889899 1.389e-09 1.942664991199081 1.39e-09 1.8265563188207443 1.391e-09 1.789928617674396 1.392e-09 1.7690585610807976 1.393e-09 1.7599596431199311 1.394e-09 1.7649533003048568 1.395e-09 1.849209596069471 1.396e-09 1.8319748563596503 1.397e-09 1.8377100591741795 1.398e-09 1.740623905867218 1.399e-09 1.8174193715738012 1.4e-09 1.764942847158238 1.401e-09 1.7559057703317973 1.402e-09 1.7391526675789222 1.403e-09 1.7893303148068402 1.404e-09 1.7568744576949147 1.405e-09 1.7981883390388178 1.406e-09 1.9424229888278202 1.407e-09 1.802411190758668 1.4079999999999999e-09 1.7900511720503698 1.409e-09 1.9168387290737332 1.4099999999999999e-09 1.794411177214847 1.411e-09 1.7828647848885097 1.4119999999999999e-09 1.7809106640585222 1.413e-09 1.6819428018878253 1.4139999999999999e-09 1.7690544972186801 1.415e-09 1.8256517119833742 1.416e-09 1.8869420236317234 1.417e-09 1.718688924982191 1.418e-09 1.8309494936054826 1.419e-09 1.8387842579907676 1.42e-09 1.764196469232774 1.421e-09 1.8176800266742563 1.422e-09 1.7342051378594374 1.423e-09 1.8156456970936903 1.424e-09 1.8445432725451483 1.425e-09 1.8248351510847 1.426e-09 1.7983893447760733 1.427e-09 1.847293250371805 1.428e-09 1.8513287845916808 1.429e-09 1.6799625444008002 1.43e-09 1.8642456099791218 1.431e-09 1.8143643289392826 1.432e-09 1.8732400102789843 1.433e-09 1.8289204184641656 1.434e-09 1.8157072726784413 1.435e-09 1.7140949013820075 1.436e-09 1.8154398326414045 1.437e-09 1.8811177400945487 1.438e-09 1.7794553552666472 1.4389999999999999e-09 1.8086058808422938 1.44e-09 1.7400653564267383 1.4409999999999999e-09 1.748930182593335 1.442e-09 1.865613074242582 1.4429999999999999e-09 1.8896560882467022 1.444e-09 1.849584630139533 1.4449999999999999e-09 1.7665578374063513 1.446e-09 1.7336306986887808 1.447e-09 1.762411530937544 1.448e-09 1.795506150935001 1.449e-09 1.8119233411493063 1.45e-09 1.7058398177016176 1.451e-09 1.7648822093035321 1.452e-09 1.840929588557277 1.453e-09 1.8345034701479008 1.454e-09 1.8303257641790736 1.455e-09 1.8803813846771322 1.456e-09 1.7518542642838075 1.457e-09 1.8011014238138978 1.458e-09 1.7469382783923704 1.459e-09 1.785702384517498 1.46e-09 1.786324841507256 1.461e-09 1.7369247240908439 1.462e-09 1.7523145823206905 1.463e-09 1.7707628864539189 1.464e-09 1.7157776917217773 1.465e-09 1.7681271812198542 1.466e-09 1.8586221560234115 1.467e-09 1.800794132114973 1.4679999999999999e-09 1.8047843066455331 1.469e-09 1.7245106374920995 1.4699999999999999e-09 1.799725351696766 1.471e-09 1.8304067483751791 1.4719999999999999e-09 1.8759612331383657 1.473e-09 1.8732721187367356 1.4739999999999999e-09 1.7271599037325889 1.475e-09 1.839466896848736 1.476e-09 1.7658028902415992 1.477e-09 1.7418452896674117 1.478e-09 1.7682763977401357 1.479e-09 1.7801466000349904 1.48e-09 1.8181821462261802 1.481e-09 1.8191771560319405 1.482e-09 1.8568998291512884 1.483e-09 1.848961238339654 1.484e-09 1.8070101408726786 1.485e-09 1.820052759503086 1.486e-09 1.7868188594134535 1.487e-09 1.7667535734999869 1.488e-09 1.77544393020147 1.489e-09 1.7768092953810364 1.49e-09 1.8128313004295133 1.491e-09 1.7795800083486257 1.492e-09 1.877641908245959 1.493e-09 1.8071904483974934 1.494e-09 1.8177039279179634 1.495e-09 1.8523621106844097 1.496e-09 1.7709689918688192 1.497e-09 1.75825336271809 1.498e-09 1.8217007675290426 1.4989999999999999e-09 1.8326380061896148 1.5e-09 1.8097449263005585 1.5009999999999999e-09 1.813308096299691 1.502e-09 1.8178538072599704 1.5029999999999999e-09 1.833431699583637 1.504e-09 1.6914787066999168 1.5049999999999999e-09 1.7633822804071757 1.506e-09 1.7568340020345297 1.507e-09 1.771816477500553 1.508e-09 1.7724735843646817 1.509e-09 1.7412360197585735 1.51e-09 1.7752896837364478 1.511e-09 1.8373540633883516 1.512e-09 1.8956698157611842 1.513e-09 1.8136745465925805 1.514e-09 1.8121810826869125 1.515e-09 1.8328397878540954 1.516e-09 1.850671079385113 1.517e-09 1.8940720461873244 1.518e-09 1.7468259653525668 1.519e-09 1.7892247426947565 1.52e-09 1.7274317710169167 1.521e-09 1.8344719763637682 1.522e-09 1.8059940265259466 1.523e-09 1.7329123524297168 1.524e-09 1.8624960410491875 1.525e-09 1.7677920714173492 1.526e-09 1.7987497956242002 1.527e-09 1.8654898548099186 1.5279999999999999e-09 1.7965783129300217 1.529e-09 1.7655290826022194 1.5299999999999999e-09 1.8439177576075763 1.531e-09 1.7942557587949777 1.5319999999999999e-09 1.7619034267898686 1.533e-09 1.849453796656738 1.5339999999999999e-09 1.731159383855718 1.535e-09 1.7601915514351725 1.536e-09 1.7125321656204582 1.537e-09 1.7883061796189277 1.538e-09 1.7544650424770238 1.539e-09 1.8403429802580444 1.54e-09 1.8013854856396325 1.541e-09 1.8112544780392459 1.542e-09 1.737713422940047 1.543e-09 1.8549718045799135 1.544e-09 1.8695250431253665 1.545e-09 1.8029717246468875 1.546e-09 1.8385532670009952 1.547e-09 1.797544197031937 1.548e-09 1.7204544592458486 1.549e-09 1.8266378953892053 1.55e-09 1.7667813566542758 1.551e-09 1.7456221593975818 1.552e-09 1.7873142789098664 1.553e-09 1.8976796946400558 1.554e-09 1.8480383675899543 1.555e-09 1.8210746016958395 1.556e-09 1.7580199920763249 1.5569999999999999e-09 1.8060624681681396 1.558e-09 1.8087735593321532 1.5589999999999999e-09 1.8580861393156585 1.56e-09 1.7389176902502117 1.5609999999999999e-09 1.8675300833565356 1.562e-09 1.8400792621438828 1.5629999999999999e-09 1.7647441307017162 1.564e-09 1.6885160707159323 1.5649999999999999e-09 1.9184891009518446 1.566e-09 1.847601972305364 1.567e-09 1.826459719091489 1.568e-09 1.7259350933660742 1.569e-09 1.766577021859634 1.57e-09 1.8371504242449936 1.571e-09 1.7535809293727425 1.572e-09 1.7083470934724823 1.573e-09 1.8396604612289276 1.574e-09 1.8088998383594195 1.575e-09 1.805900995911195 1.576e-09 1.8044038662651412 1.577e-09 1.767318724132039 1.578e-09 1.81835705409212 1.579e-09 1.8781683863277547 1.58e-09 1.8348311597675244 1.581e-09 1.7994484140418014 1.582e-09 1.809738644461062 1.583e-09 1.8638426232620295 1.584e-09 1.8889270195640078 1.585e-09 1.8361261635356985 1.586e-09 1.781412837646459 1.587e-09 1.7768522613334474 1.5879999999999999e-09 1.7983747742101104 1.589e-09 1.8279562575214858 1.5899999999999999e-09 1.8418201032928312 1.591e-09 1.7647477804307588 1.5919999999999999e-09 1.7795412466277287 1.593e-09 1.799022300302217 1.5939999999999999e-09 1.810389803042104 1.595e-09 1.8896614660565503 1.5959999999999999e-09 1.876023740011681 1.597e-09 1.8234405810780123 1.598e-09 1.8006892821636744 1.599e-09 1.850044597095915 1.6e-09 1.7564348571360398 1.601e-09 1.8460182637307854 1.602e-09 1.7845181974459983 1.603e-09 1.7031275273905495 1.604e-09 1.9145887349731687 1.605e-09 1.8423155826423907 1.606e-09 1.7980971984869325 1.607e-09 1.7296646979957155 1.608e-09 1.8547199284202174 1.609e-09 1.7424282996967202 1.61e-09 1.8114842717753126 1.611e-09 1.7576655446909042 1.612e-09 1.805488540550859 1.613e-09 1.8734898518273666 1.614e-09 1.7816889027858573 1.615e-09 1.734367942742619 1.616e-09 1.898342420278017 1.6169999999999999e-09 1.785354916423978 1.618e-09 1.8114748672050494 1.6189999999999999e-09 1.7799371773388148 1.62e-09 1.6753974295813128 1.6209999999999999e-09 1.7872880139758371 1.622e-09 1.7846883914065763 1.6229999999999999e-09 1.7766070543834942 1.624e-09 1.8392280987267335 1.6249999999999999e-09 1.74998377235358 1.626e-09 1.7399183179671125 1.627e-09 1.8475426767928738 1.628e-09 1.791977756546757 1.629e-09 1.7640892607303469 1.63e-09 1.7900471918353467 1.631e-09 1.8355681283704819 1.632e-09 1.7926427053392355 1.633e-09 1.88171589739271 1.634e-09 1.7770789983617987 1.635e-09 1.8016466409789071 1.636e-09 1.8085488421477736 1.637e-09 1.849931260126366 1.638e-09 1.8067289372925426 1.639e-09 1.7238652861882964 1.64e-09 1.7981033648313909 1.641e-09 1.81143742124418 1.642e-09 1.7917616549998214 1.643e-09 1.758116340138363 1.644e-09 1.7700568524645068 1.645e-09 1.8166467252495202 1.646e-09 1.7518118223834025 1.647e-09 1.7654329443100893 1.6479999999999999e-09 1.7707758703511738 1.649e-09 1.7106719317782508 1.6499999999999999e-09 1.8079931433888017 1.651e-09 1.8112920035167326 1.6519999999999999e-09 1.782417748700467 1.653e-09 1.8747578472514177 1.6539999999999999e-09 1.8343692317810008 1.655e-09 1.771343392817841 1.6559999999999999e-09 1.7474338597283214 1.657e-09 1.8084528702878775 1.658e-09 1.8336025842390296 1.659e-09 1.8262084029798915 1.66e-09 1.7098823318280505 1.661e-09 1.7495508840877874 1.662e-09 1.8273504419571402 1.663e-09 1.8009601860429243 1.664e-09 1.7172665502115703 1.665e-09 1.892319821503463 1.666e-09 1.7832066296766436 1.667e-09 1.7708445652987006 1.668e-09 1.661204674345291 1.669e-09 1.8188701663645026 1.67e-09 1.8519622823884194 1.671e-09 1.8319032806074123 1.672e-09 1.7674893453592253 1.673e-09 1.765784612948654 1.674e-09 1.6895063306463638 1.675e-09 1.7715789660976227 1.676e-09 1.816468853459656 1.6769999999999999e-09 1.8278408783417681 1.678e-09 1.688450294801438 1.6789999999999999e-09 1.737469416282209 1.68e-09 1.7363669782686535 1.6809999999999999e-09 1.8159207357486478 1.682e-09 1.8436839903949593 1.6829999999999999e-09 1.7957750226627183 1.684e-09 1.8176049010484896 1.6849999999999999e-09 1.8368400670868623 1.686e-09 1.7251439092936964 1.687e-09 1.8499891785367606 1.688e-09 1.7870871843100045 1.689e-09 1.8725873571978409 1.69e-09 1.782433225851356 1.691e-09 1.704581251943944 1.692e-09 1.7848197145450322 1.693e-09 1.783327079719334 1.694e-09 1.8342596848733246 1.695e-09 1.764744488512242 1.696e-09 1.8258037732218053 1.697e-09 1.8004495625609962 1.698e-09 1.8561216827369516 1.699e-09 1.8265508572765154 1.7e-09 1.7865876161518606 1.701e-09 1.8445857209212193 1.702e-09 1.783675541955301 1.703e-09 1.804549698544078 1.704e-09 1.7503439035874362 1.705e-09 1.7852836554197689 1.706e-09 1.746924186528206 1.707e-09 1.8848705870382685 1.7079999999999999e-09 1.744067897043014 1.709e-09 1.7581007387137515 1.7099999999999999e-09 1.7320601978296233 1.711e-09 1.7647792189917706 1.7119999999999999e-09 1.674832987958289 1.713e-09 1.8947716412891322 1.7139999999999999e-09 1.8689648909904624 1.715e-09 1.770729993561805 1.7159999999999999e-09 1.787067465163069 1.717e-09 1.7687404106375728 1.718e-09 1.797560518942488 1.719e-09 1.8112806360280773 1.72e-09 1.822306651188418 1.721e-09 1.8256385768774597 1.722e-09 1.8114050220077798 1.723e-09 1.90643353789987 1.724e-09 1.7632817062208008 1.725e-09 1.87259206746568 1.726e-09 1.8393605451634358 1.727e-09 1.774680470287165 1.728e-09 1.850460739127548 1.729e-09 1.7836232262864917 1.73e-09 1.7994180258438124 1.731e-09 1.8413310392524191 1.732e-09 1.8032349716225073 1.733e-09 1.8486667638678878 1.734e-09 1.8215038321756847 1.735e-09 1.859414353970539 1.736e-09 1.7763148470702315 1.7369999999999999e-09 1.7776670222307156 1.738e-09 1.9098994639020765 1.7389999999999999e-09 1.7689647026779323 1.74e-09 1.740601474025087 1.7409999999999999e-09 1.847557016144837 1.742e-09 1.811941443814922 1.7429999999999999e-09 1.8319911272308305 1.744e-09 1.78767029899441 1.7449999999999999e-09 1.6984926567879413 1.746e-09 1.843105070776269 1.747e-09 1.8352413786981105 1.748e-09 1.8221452272928897 1.749e-09 1.7740895955567582 1.75e-09 1.7653775205887423 1.751e-09 1.8925885411181769 1.752e-09 1.87182212286232 1.753e-09 1.790530624921752 1.754e-09 1.777718555916723 1.755e-09 1.719069634265909 1.756e-09 1.8563662813822817 1.757e-09 1.8000602373008787 1.758e-09 1.685304004287342 1.759e-09 1.8104080050884237 1.76e-09 1.8724486918269676 1.761e-09 1.6922943685738265 1.762e-09 1.805183570758772 1.763e-09 1.7949913054305853 1.764e-09 1.8472053020444683 1.765e-09 1.7238471171003957 1.766e-09 1.734360564976084 1.767e-09 1.7031171483409737 1.7679999999999999e-09 1.8342593756481755 1.769e-09 1.7862519167905604 1.7699999999999999e-09 1.7567959754447544 1.771e-09 1.746674728310066 1.7719999999999999e-09 1.8950204307435317 1.773e-09 1.8758627341974519 1.7739999999999999e-09 1.7853115972089904 1.775e-09 1.837547335886003 1.7759999999999999e-09 1.9300308665315136 1.777e-09 1.815661990375861 1.778e-09 1.748839027824953 1.779e-09 1.7756358118650009 1.78e-09 1.9023151953081772 1.781e-09 1.7878699037795702 1.782e-09 1.7083631669237025 1.783e-09 1.8100142376096193 1.784e-09 1.769971406123004 1.785e-09 1.8086823962564058 1.786e-09 1.7344485756014008 1.787e-09 1.8106358757394212 1.788e-09 1.7098530774972531 1.789e-09 1.7924271946865633 1.79e-09 1.7620767230847099 1.791e-09 1.7962028654605413 1.792e-09 1.8393479945133908 1.793e-09 1.8568782003627207 1.794e-09 1.7515189820303296 1.795e-09 1.8007390427564218 1.796e-09 1.7772718547826543 1.7969999999999999e-09 1.747941383796009 1.798e-09 1.8360442197617133 1.7989999999999999e-09 1.7967545249287524 1.8e-09 1.6744526841431164 1.8009999999999999e-09 1.7929161254464476 1.802e-09 1.7880570503464885 1.8029999999999999e-09 1.7932958510575654 1.804e-09 1.80569519935621 1.8049999999999999e-09 1.8008942869793294 1.806e-09 1.7941696348155192 1.8069999999999999e-09 1.7649075032696229 1.808e-09 1.8073378716785493 1.809e-09 1.8473227310474298 1.81e-09 1.7503610638119074 1.811e-09 1.761437507352811 1.812e-09 1.809832132840123 1.813e-09 1.832696896072372 1.814e-09 1.857384755590635 1.815e-09 1.8334884893617969 1.816e-09 1.8551664700308061 1.817e-09 1.7079383068406355 1.818e-09 1.7731122709094942 1.819e-09 1.7494266720385045 1.82e-09 1.8294082415930653 1.821e-09 1.7640417757352294 1.822e-09 1.763503577479405 1.823e-09 1.7854450123695822 1.824e-09 1.749394784379041 1.825e-09 1.7508664152086997 1.826e-09 1.857434333208734 1.827e-09 1.7716004623261097 1.8279999999999999e-09 1.7845431727019558 1.829e-09 1.8083000196520285 1.8299999999999999e-09 1.7618943071413222 1.831e-09 1.8623688551516595 1.8319999999999999e-09 1.787677357467324 1.833e-09 1.764922325924321 1.8339999999999999e-09 1.8494479027837474 1.835e-09 1.7796351326405557 1.8359999999999999e-09 1.7469524342503973 1.837e-09 1.7341803672423188 1.838e-09 1.7765510881190525 1.839e-09 1.8317347748977357 1.84e-09 1.8088656876943057 1.841e-09 1.7857352774334585 1.842e-09 1.8085996195241087 1.843e-09 1.7754240094938443 1.844e-09 1.777323642728545 1.845e-09 1.7780715540283114 1.846e-09 1.7505300182926862 1.847e-09 1.77096138057907 1.848e-09 1.816192239654103 1.849e-09 1.6850949790553718 1.85e-09 1.8209846122520061 1.851e-09 1.7355342361239545 1.852e-09 1.7971077265258513 1.853e-09 1.8123609715662872 1.854e-09 1.767006824438773 1.855e-09 1.8109504739818114 1.856e-09 1.8291723582007333 1.8569999999999999e-09 1.8176855111890642 1.858e-09 1.8417384230290827 1.8589999999999999e-09 1.7609852488508655 1.86e-09 1.7685699288106935 1.8609999999999999e-09 1.8227503260480264 1.862e-09 1.7510591652165997 1.863e-09 1.8563774405173652 1.8639999999999998e-09 1.7420226986949112 1.865e-09 1.8524401527316459 1.866e-09 1.8452123595121384 1.867e-09 1.7963257145991034 1.868e-09 1.815912940484569 1.869e-09 1.8774144533489923 1.87e-09 1.7660022365235337 1.871e-09 1.8414335193332783 1.872e-09 1.9385007046105676 1.873e-09 1.8060811100486502 1.874e-09 1.8792795317193893 1.875e-09 1.7925507542569248 1.876e-09 1.855938302292495 1.877e-09 1.7663246537579245 1.878e-09 1.7076790874899912 1.879e-09 1.8059971290921013 1.88e-09 1.8827661663048878 1.881e-09 1.8513664620906891 1.882e-09 1.7776467974335963 1.883e-09 1.772761533421408 1.884e-09 1.9075664185201247 1.885e-09 1.792027077110943 1.886e-09 1.748410016116054 1.8869999999999998e-09 1.8172006687732811 1.888e-09 1.7383586928515373 1.889e-09 1.8425690190611332 1.89e-09 1.885877770377609 1.8909999999999998e-09 1.80533380036759 1.892e-09 1.8252008428693582 1.893e-09 1.7688119820168107 1.894e-09 1.830772448718816 1.8949999999999998e-09 1.8157240555671963 1.896e-09 1.7097223571401567 1.897e-09 1.8155167478373169 1.898e-09 1.7712324403512723 1.899e-09 1.7761857369311616 1.9e-09 1.7589937619099707 1.901e-09 1.856536476248045 1.902e-09 1.821195395783206 1.903e-09 1.6873627214796463 1.904e-09 1.7384586777855104 1.905e-09 1.8078844858831327 1.906e-09 1.8594208495621225 1.907e-09 1.8657463392528124 1.908e-09 1.8464187624862107 1.909e-09 1.7706928235205082 1.91e-09 1.8567854684442535 1.911e-09 1.9024380850087017 1.912e-09 1.7464875605762318 1.913e-09 1.8789724501786298 1.914e-09 1.8082371135655415 1.915e-09 1.8518239063730881 1.916e-09 1.8270428202012545 1.917e-09 1.7466329984455857 1.9179999999999998e-09 1.8234488792280799 1.919e-09 1.789517019844906 1.92e-09 1.8225658108889509 1.921e-09 1.8367389848028544 1.9219999999999998e-09 1.7649405257778121 1.923e-09 1.796612775616442 1.924e-09 1.7956320341160312 1.925e-09 1.7903614808211976 1.9259999999999998e-09 1.903077553634768 1.927e-09 1.8144468078353437 1.928e-09 1.7433867004255619 1.929e-09 1.7583419733304537 1.93e-09 1.869309320666432 1.931e-09 1.7466883804274582 1.932e-09 1.8155759072601518 1.933e-09 1.8154279226067727 1.934e-09 1.8120216842409609 1.935e-09 1.765672504797491 1.936e-09 1.762113080400395 1.937e-09 1.7788776266031385 1.938e-09 1.77111464636533 1.939e-09 1.794178602906243 1.94e-09 1.7774980794420867 1.941e-09 1.7393328161813901 1.942e-09 1.8370973556648458 1.943e-09 1.8759747558700104 1.944e-09 1.8542961862672318 1.945e-09 1.7697183604614237 1.946e-09 1.8562313580043068 1.947e-09 1.775875639578808 1.948e-09 1.8375003925553588 1.9489999999999998e-09 1.7754596952032236 1.95e-09 1.8453094708275983 1.951e-09 1.7794681246358004 1.952e-09 1.7442313026487801 1.9529999999999998e-09 1.826625433593038 1.954e-09 1.7983939460931095 1.955e-09 1.8459197262034208 1.956e-09 1.8864636461007807 1.9569999999999998e-09 1.8335335781623463 1.958e-09 1.7431400471608443 1.959e-09 1.8595490102109595 1.96e-09 1.7769950153687863 1.961e-09 1.8363415844384023 1.962e-09 1.7295967724679844 1.963e-09 1.8101377001346837 1.964e-09 1.8000596002341192 1.965e-09 1.722801680746021 1.966e-09 1.8572864564969234 1.967e-09 1.7851496029094789 1.968e-09 1.8178378898050371 1.969e-09 2.000555807753832 1.97e-09 1.804801198646417 1.971e-09 1.8062811711897688 1.972e-09 1.7799356499156436 1.973e-09 1.8455095103668326 1.974e-09 1.812322738091176 1.975e-09 1.800248893203056 1.976e-09 1.8912638168225488 1.977e-09 1.7919389206506324 1.978e-09 1.8699046082661388 1.979e-09 1.7511640206630492 1.9799999999999998e-09 1.7067001659344383 1.981e-09 1.8489354884183795 1.982e-09 1.8155304394278728 1.983e-09 1.8212187218419642 1.9839999999999998e-09 1.755529292446399 1.985e-09 1.765617594570193 1.986e-09 1.8064081669386318 1.987e-09 1.8299173529367887 1.988e-09 1.7858664734470897 1.989e-09 1.7884114546245287 1.99e-09 1.7615130619176749 1.991e-09 1.8127916152824974 1.992e-09 1.7956671828545911 1.993e-09 1.749794706773225 1.994e-09 1.7845271649457461 1.995e-09 1.8348027068327823 1.996e-09 1.7357819557783416 1.997e-09 1.8382385237939223 1.998e-09 1.8021084119900195 1.999e-09 1.7961246548846244 2e-09 1.7001268337191668 2.001e-09 1.814303251589181 2.002e-09 1.8080944483244952 2.003e-09 1.7411819339976264 2.004e-09 1.724784241033908 2.005e-09 1.8898862173999178 2.006e-09 1.8119947000753645 2.0069999999999998e-09 1.805523773029348 2.008e-09 1.8380434642674732 2.009e-09 1.8420406550618154 2.01e-09 1.835411697058803 2.0109999999999998e-09 1.8348798936942163 2.012e-09 1.8112376476533862 2.013e-09 1.7785418038856604 2.014e-09 1.7406910554904658 2.0149999999999998e-09 1.8514220661213245 2.016e-09 1.8811219603944467 2.017e-09 1.7361561020172513 2.018e-09 1.8018550120601775 2.019e-09 1.8416486877289806 2.02e-09 1.7688358794447898 2.021e-09 1.8049408884652194 2.022e-09 1.867176372679273 2.023e-09 1.7588464307328622 2.024e-09 1.7773372402586962 2.025e-09 1.7933724026089115 2.026e-09 1.8043467267483764 2.027e-09 1.8919207848959896 2.028e-09 1.838099182001708 2.029e-09 1.855216908371293 2.03e-09 1.8045003800264126 2.031e-09 1.7963816440344913 2.032e-09 1.6789774021073063 2.033e-09 1.7941775474334063 2.034e-09 1.7637316879145242 2.035e-09 1.75723338674449 2.036e-09 1.8411758245693728 2.037e-09 1.7598532919807721 2.0379999999999998e-09 1.813549030665099 2.039e-09 1.8704001222426045 2.04e-09 1.7751857121557824 2.041e-09 1.759997437514286 2.0419999999999998e-09 1.7935150680200553 2.043e-09 1.8135775090933373 2.044e-09 1.7783195527725535 2.045e-09 1.7573164552889249 2.0459999999999998e-09 1.8333128756907733 2.047e-09 1.83255561777123 2.048e-09 1.854333148059684 2.049e-09 1.830508112234908 2.05e-09 1.8089214210894078 2.051e-09 1.820324052086923 2.052e-09 1.8162152028412717 2.053e-09 1.721072297345987 2.054e-09 1.7609456948546738 2.055e-09 1.8228906864710963 2.056e-09 1.8163364240202418 2.057e-09 1.8255894779656814 2.058e-09 1.7878958733987713 2.059e-09 1.8391741920224516 2.06e-09 1.71521705250833 2.061e-09 1.772384494204397 2.062e-09 1.809041949017818 2.063e-09 1.9733111690195237 2.064e-09 1.8068890139043812 2.065e-09 1.797920015427204 2.066e-09 1.7636176191721629 2.067e-09 1.797830673989838 2.068e-09 1.819410627422258 2.0689999999999998e-09 1.8111989316136228 2.07e-09 1.7729810971958215 2.071e-09 1.7817567982189515 2.072e-09 1.7025738485321171 2.0729999999999998e-09 1.812749511389374 2.074e-09 1.8622974553041418 2.075e-09 1.751606707309626 2.076e-09 1.7226271371164454 2.0769999999999998e-09 1.7700309087567974 2.078e-09 1.797662524632627 2.079e-09 1.7560906389346307 2.08e-09 1.7487447984853417 2.081e-09 1.775644047007772 2.082e-09 1.882471424809917 2.083e-09 1.8183315145787367 2.084e-09 1.7996730476743215 2.085e-09 1.8566631454241789 2.086e-09 1.7995900277950618 2.087e-09 1.7973009586786062 2.088e-09 1.7561202460726502 2.089e-09 1.8317360357265429 2.09e-09 1.7442540485631552 2.091e-09 1.8596053324149804 2.092e-09 1.8046920862499314 2.093e-09 1.7685544973264884 2.094e-09 1.8527162724618214 2.095e-09 1.6965967759090925 2.0959999999999998e-09 1.8744941155190473 2.097e-09 1.7953411511861526 2.098e-09 1.7433798893517558 2.099e-09 1.8007439445975093 2.0999999999999998e-09 1.7955186192867978 2.101e-09 1.8372661127701542 2.102e-09 1.8176378622994473 2.103e-09 1.8028303261134146 2.1039999999999998e-09 1.8136774410643648 2.105e-09 1.7198589857636908 2.106e-09 1.8081139850895376 2.107e-09 1.70252754296136 2.1079999999999998e-09 1.8095864828316814 2.109e-09 1.7007455455595608 2.11e-09 1.8631080325448899 2.111e-09 1.856089875148557 2.112e-09 1.7604478844650486 2.113e-09 1.7870116115655577 2.114e-09 1.804727872600552 2.115e-09 1.8047025374046737 2.116e-09 1.8308476697614986 2.117e-09 1.8082890355323853 2.118e-09 1.7856977030442487 2.119e-09 1.8035481520739778 2.12e-09 1.728791206133946 2.121e-09 1.765423817367657 2.122e-09 1.7862489275190576 2.123e-09 1.8468793526949685 2.124e-09 1.763649778823239 2.125e-09 1.8406493111832574 2.126e-09 1.8219161386170806 2.1269999999999998e-09 1.8418866691022004 2.128e-09 1.8750389244111212 2.129e-09 1.8210254053221786 2.13e-09 1.7831692950473665 2.1309999999999998e-09 1.788413119007913 2.132e-09 1.739512956688317 2.133e-09 1.710392970843595 2.134e-09 1.788689198070775 2.1349999999999998e-09 1.7799983115232691 2.136e-09 1.713396929503704 2.137e-09 1.8612232010274468 2.138e-09 1.7970783840641231 2.139e-09 1.7895261980578208 2.14e-09 1.8201893211002536 2.141e-09 1.846523640397396 2.142e-09 1.7548841575259087 2.143e-09 1.8530727949562984 2.144e-09 1.8751825959852053 2.145e-09 1.7504073116173535 2.146e-09 1.8754313879368902 2.147e-09 1.8144947280770694 2.148e-09 1.859474707046092 2.149e-09 1.7811279145846537 2.15e-09 1.8270912457117376 2.151e-09 1.812020942558207 2.152e-09 1.84072411513405 2.153e-09 1.8794175852980566 2.154e-09 1.7672462971123497 2.155e-09 1.7882690742369727 2.156e-09 1.7960489307686762 2.157e-09 1.856698006701607 2.1579999999999998e-09 1.8223440521269834 2.159e-09 1.8519406202376094 2.16e-09 1.842387628378668 2.161e-09 1.7362397913135608 2.1619999999999998e-09 1.7264769481638265 2.163e-09 1.8366783087609782 2.164e-09 1.9339389110987868 2.165e-09 1.7836488588339654 2.1659999999999998e-09 1.803340015978087 2.167e-09 1.7827102689152667 2.168e-09 1.7330295954320543 2.169e-09 1.7225861311354593 2.17e-09 1.722081678751616 2.171e-09 1.7903277256417114 2.172e-09 1.7027288944360799 2.173e-09 1.7520016432178145 2.174e-09 1.8481313404438133 2.175e-09 1.6972251216600418 2.176e-09 1.8497485043668973 2.177e-09 1.822116523900865 2.178e-09 1.8214741497337057 2.179e-09 1.8617009778849516 2.18e-09 1.8005236356004914 2.181e-09 1.782020638129185 2.182e-09 1.8244429298552112 2.183e-09 1.8158364508957707 2.184e-09 1.7746191974972436 2.185e-09 1.797393312824731 2.186e-09 1.8492772404796936 2.187e-09 1.8166341461893434 2.188e-09 1.7696802654404276 2.1889999999999998e-09 1.7841599198039357 2.19e-09 1.792613915802171 2.191e-09 1.734601646783377 2.192e-09 1.7719067013394574 2.1929999999999998e-09 1.8701429389757551 2.194e-09 1.9037594531378925 2.195e-09 1.8503851622894847 2.196e-09 1.7593333714052561 2.1969999999999998e-09 1.7182060713397862 2.198e-09 1.8310639832340327 2.199e-09 1.850708158792943 2.2e-09 1.8752371477649115 2.201e-09 1.75018010735786 2.202e-09 1.721087024707753 2.203e-09 1.8643010621365579 2.204e-09 1.803805342620084 2.205e-09 1.7552758360486984 2.206e-09 1.841123833227943 2.207e-09 1.8246749483519933 2.208e-09 1.7837962409726336 2.209e-09 1.8585963928157705 2.21e-09 1.7683465014352895 2.211e-09 1.8180899791494574 2.212e-09 1.868086317048989 2.213e-09 1.8203054861450148 2.214e-09 1.8376103178251022 2.215e-09 1.7972968432296215 2.2159999999999998e-09 1.777309596999076 2.217e-09 1.8319064624142827 2.218e-09 1.7862483437061265 2.219e-09 1.782704889589241 2.2199999999999998e-09 1.7851535704017203 2.221e-09 1.7750154042401356 2.222e-09 1.839428702406151 2.223e-09 1.7666344621328605 2.2239999999999998e-09 1.7609180079410045 2.225e-09 1.6984284505046623 2.226e-09 1.837407700979508 2.227e-09 1.835421839736687 2.2279999999999998e-09 1.8532866636101408 2.229e-09 1.8337214377202329 2.23e-09 1.7942334898200298 2.231e-09 1.8684315509008895 2.232e-09 1.9105219454930806 2.233e-09 1.8407188251794313 2.234e-09 1.7835174479141394 2.235e-09 1.7860900131233608 2.236e-09 1.7808274745464947 2.237e-09 1.821973677268381 2.238e-09 1.7788606866306131 2.239e-09 1.7784875262545166 2.24e-09 1.7682080919848628 2.241e-09 1.8149160577523435 2.242e-09 1.781636134403415 2.243e-09 1.7584528283031011 2.244e-09 1.798609570737421 2.245e-09 1.7963634515395737 2.246e-09 1.7416355616424308 2.2469999999999998e-09 1.8372864747284994 2.248e-09 1.8264947434922953 2.249e-09 1.8346922239151782 2.25e-09 1.8814806797252177 2.2509999999999998e-09 1.7179741140099727 2.252e-09 1.736405374048076 2.253e-09 1.840897864600346 2.254e-09 1.8408946905205459 2.2549999999999998e-09 1.7402961784480964 2.256e-09 1.806007851670607 2.257e-09 1.8044650030325253 2.258e-09 1.7896164624170834 2.259e-09 1.8808968189030986 2.26e-09 1.8798266956057204 2.261e-09 1.7993321227024293 2.262e-09 1.6898257493150146 2.263e-09 1.7776138404338668 2.264e-09 1.8630757706119812 2.265e-09 1.750117842302465 2.266e-09 1.8220893665837585 2.267e-09 1.8401741024543523 2.268e-09 1.7476659930094713 2.269e-09 1.704061461068686 2.27e-09 1.8838188889715362 2.271e-09 1.7528600603527333 2.272e-09 1.7963743922897935 2.273e-09 1.7458284410897826 2.274e-09 1.8191398634580154 2.275e-09 1.8465285652631913 2.276e-09 1.7958504014107588 2.277e-09 1.7666859763784886 2.2779999999999998e-09 1.790002024554434 2.279e-09 1.8486018378684124 2.28e-09 1.8204992321807072 2.281e-09 1.7523819990054648 2.2819999999999998e-09 1.8511179835964975 2.283e-09 1.8911690852751375 2.284e-09 1.8234325885674016 2.285e-09 1.7991876450184174 2.2859999999999998e-09 1.7708031322854352 2.287e-09 1.8727229765574054 2.288e-09 1.7637543579271044 2.289e-09 1.8624788801271597 2.29e-09 1.7870154302329782 2.291e-09 1.8341666037710118 2.292e-09 1.7653531616807037 2.293e-09 1.8002563525233892 2.294e-09 1.9052973213006157 2.295e-09 1.7924835470891978 2.296e-09 1.7411411712958076 2.297e-09 1.7993118053450483 2.298e-09 1.7988941407615846 2.299e-09 1.7968315641029737 2.3e-09 1.761503157685743 2.301e-09 1.7739960742633307 2.302e-09 1.8051119262105648 2.303e-09 1.816203747072596 2.304e-09 1.7430483773288037 2.305e-09 1.8108295852237124 2.306e-09 1.7316774230397831 2.307e-09 1.817121376546284 2.308e-09 1.8319824726837715 2.3089999999999998e-09 1.8350972522558304 2.31e-09 1.8373031228344416 2.311e-09 1.8160024905102254 2.312e-09 1.792217408414541 2.3129999999999998e-09 1.8723050884197667 2.314e-09 1.778889092340378 2.315e-09 1.8540380012928757 2.316e-09 1.7983072243453506 2.3169999999999998e-09 1.7905899870849835 2.318e-09 1.8073695852952292 2.319e-09 1.7314217204188753 2.32e-09 1.7839564132874297 2.321e-09 1.7336910520994493 2.322e-09 1.9027546586489674 2.323e-09 1.7567627116425986 2.324e-09 1.8856686816584682 2.325e-09 1.8825087186402234 2.326e-09 1.8130050572187524 2.327e-09 1.7549070665689601 2.328e-09 1.7903767475223953 2.329e-09 1.8064720140962254 2.33e-09 1.8109941970135244 2.331e-09 1.8023285847223025 2.332e-09 1.8759731704578846 2.333e-09 1.744807814905188 2.334e-09 1.8649162100141956 2.335e-09 1.9585761991054529 2.3359999999999998e-09 1.786701397984945 2.337e-09 1.7589151398513188 2.338e-09 1.8773242681047553 2.339e-09 1.853544343331604 2.3399999999999998e-09 1.6596471858514743 2.341e-09 1.691251571740068 2.342e-09 1.7655037084002265 2.343e-09 1.836313873136797 2.3439999999999998e-09 1.753071746605256 2.345e-09 1.7793438275899633 2.346e-09 1.8292960679164292 2.347e-09 1.8756466404420151 2.3479999999999998e-09 1.8270677748597697 2.349e-09 1.8164660760307805 2.35e-09 1.8193143785199186 2.351e-09 1.7445263680439491 2.352e-09 1.8429622631432245 2.353e-09 1.8101561674720135 2.354e-09 1.8409345701798059 2.355e-09 1.767652888003606 2.356e-09 1.7342989465626666 2.357e-09 1.7955217998999176 2.358e-09 1.8452858915663886 2.359e-09 1.787649514603989 2.36e-09 1.8490339272550556 2.361e-09 1.7816804163447557 2.362e-09 1.7427956822596682 2.363e-09 1.8045431038006128 2.364e-09 1.8904483259650995 2.365e-09 1.8972568299955264 2.366e-09 1.7669546267154057 2.3669999999999998e-09 1.9156062259021998 2.368e-09 1.819127757248027 2.369e-09 1.8026601091144638 2.37e-09 1.7282597579932386 2.3709999999999998e-09 1.8380619301799657 2.372e-09 1.8092566230528009 2.373e-09 1.8653845188554092 2.374e-09 1.81441779841455 2.3749999999999998e-09 1.7409768020121825 2.376e-09 1.7886107040927244 2.377e-09 1.805300477919104 2.378e-09 1.7749524067359361 2.3789999999999997e-09 1.8218381828913441 2.38e-09 1.7438152611201967 2.381e-09 1.712830941714298 2.382e-09 1.819130718880955 2.383e-09 1.7911827308584503 2.384e-09 1.7633578312529814 2.385e-09 1.7697708949293323 2.386e-09 1.7008962733329973 2.387e-09 1.8029480195487997 2.388e-09 1.8094564570121563 2.389e-09 1.8415708943075102 2.39e-09 1.8509692594073093 2.391e-09 1.8177082733629257 2.392e-09 1.7248339060431626 2.393e-09 1.753452630426304 2.394e-09 1.8281104877536862 2.395e-09 1.8057999763910213 2.396e-09 1.7879826161190824 2.397e-09 1.8829993624142918 2.3979999999999998e-09 1.843242765750632 2.399e-09 1.8370607054150758 2.4e-09 1.7531349131552774 2.401e-09 1.8275426896679967 2.4019999999999998e-09 1.7415579100430247 2.403e-09 1.8582389715528147 2.404e-09 1.7666048355266182 2.405e-09 1.8381344617898523 2.4059999999999998e-09 1.7679025235806787 2.407e-09 1.8678048763870623 2.408e-09 1.7561643443117254 2.409e-09 1.7838599060131684 2.41e-09 1.805773943493171 2.411e-09 1.8597719240850956 2.412e-09 1.8080810074758522 2.413e-09 1.803639414483628 2.414e-09 1.7550354575463243 2.415e-09 1.838350903540218 2.416e-09 1.6835220533397153 2.417e-09 1.7443180259359266 2.418e-09 1.746295797788741 2.419e-09 1.7939924114793082 2.42e-09 1.8523786801755422 2.421e-09 1.7938007414806862 2.422e-09 1.8744734880144878 2.423e-09 1.7969370965086469 2.424e-09 1.8247613111809833 2.425e-09 1.813678200115674 2.426e-09 1.8349072193275229 2.427e-09 1.7626725798106668 2.428e-09 1.7395364443282184 2.4289999999999998e-09 1.7534703924828177 2.43e-09 1.844144332127861 2.431e-09 1.6880471059609377 2.432e-09 1.7872057640349874 2.4329999999999998e-09 1.8644403165041021 2.434e-09 1.7499903911511374 2.435e-09 1.7959702342497814 2.436e-09 1.79616786782511 2.4369999999999998e-09 1.7192702847943253 2.438e-09 1.8442173971687157 2.439e-09 1.7778998348489905 2.44e-09 1.801537376310534 2.441e-09 1.770262448979509 2.442e-09 1.8036822990614885 2.443e-09 1.6992899163151072 2.444e-09 1.8372703090448395 2.445e-09 1.89787844576997 2.446e-09 1.8832035361176966 2.447e-09 1.7893736514021683 2.448e-09 1.759807395116358 2.449e-09 1.8045086398599368 2.45e-09 1.778681672855529 2.451e-09 1.6807199166802118 2.452e-09 1.8036908115891004 2.453e-09 1.8297275430334479 2.454e-09 1.743249216001368 2.455e-09 1.7936729480354725 2.4559999999999998e-09 1.7414845126232354 2.457e-09 1.7638107231067504 2.458e-09 1.773646945959692 2.459e-09 1.8176340125998263 2.4599999999999998e-09 1.762846295268268 2.461e-09 1.758739995808921 2.462e-09 1.8045258545891034 2.463e-09 1.7720990546737774 2.4639999999999998e-09 1.792504947741134 2.465e-09 1.776941271366682 2.466e-09 1.9244480956953847 2.467e-09 1.8416263194922515 2.4679999999999997e-09 1.7690022192059671 2.469e-09 1.792214890035625 2.47e-09 1.7664417230375744 2.471e-09 1.7830000502941148 2.472e-09 1.812587787205229 2.473e-09 1.8222287090445564 2.474e-09 1.814793568542333 2.475e-09 1.7181481137870003 2.476e-09 1.7570664669439564 2.477e-09 1.7342511370504339 2.478e-09 1.8752200039503208 2.479e-09 1.8462105782530138 2.48e-09 1.7675510186270078 2.481e-09 1.7120815890532288 2.482e-09 1.7848512883055672 2.483e-09 1.8307452300827607 2.484e-09 1.7735383467770125 2.485e-09 1.8664706303088803 2.486e-09 1.7073431484548514 2.4869999999999998e-09 1.827873291394038 2.488e-09 1.8231259052384012 2.489e-09 1.8081588042542027 2.49e-09 1.8029471066075466 2.4909999999999998e-09 1.763357688189723 2.492e-09 1.7712008338007885 2.493e-09 1.8411482798856278 2.494e-09 1.824243360474031 2.4949999999999998e-09 1.8066785267740808 2.496e-09 1.7586663097795656 2.497e-09 1.7932471497735396 2.498e-09 1.8147625534848015 2.4989999999999997e-09 1.8711935071477708 2.5e-09 1.771279538858893 2.501e-09 1.8356642527722895 2.502e-09 1.7786836275605429 2.503e-09 1.815455048678188 2.504e-09 1.7636062193171336 2.505e-09 1.7181485795971672 2.506e-09 1.8831732432016122 2.507e-09 1.7623196806961607 2.508e-09 1.7751167798996799 2.509e-09 1.813921020306556 2.51e-09 1.754801795420725 2.511e-09 1.8178598569808193 2.512e-09 1.7944500654604716 2.513e-09 1.8071002108835885 2.514e-09 1.7575224370706928 2.515e-09 1.7068890835275228 2.516e-09 1.7425544642910993 2.517e-09 1.794528547269032 2.5179999999999998e-09 1.7679014887718496 2.519e-09 1.8039603392261174 2.52e-09 1.8583582704617578 2.521e-09 1.8793936874106023 2.5219999999999998e-09 1.7997702130575084 2.523e-09 1.7941209244539003 2.524e-09 1.6848241979144047 2.525e-09 1.7484775385576807 2.5259999999999998e-09 1.7867602334701067 2.527e-09 1.7915495319762411 2.528e-09 1.7557977117886507 2.529e-09 1.8153526793212411 2.53e-09 1.7586968267719116 2.531e-09 1.7838914302195146 2.532e-09 1.8224686296548147 2.533e-09 1.7362992939672555 2.534e-09 1.7906753863026468 2.535e-09 1.776016403460307 2.536e-09 1.8037217776998569 2.537e-09 1.7919092757583228 2.538e-09 1.7448916296373118 2.539e-09 1.8455549164001626 2.54e-09 1.8290545808081238 2.541e-09 1.8006454853024052 2.542e-09 1.814708959409782 2.543e-09 1.8660615314035964 2.544e-09 1.813631206433834 2.545e-09 1.8689036745017216 2.546e-09 1.8215736119235788 2.547e-09 1.812021467467155 2.548e-09 1.8645331123408395 2.5489999999999998e-09 1.7406739985073902 2.55e-09 1.7372627123284898 2.551e-09 1.7747422065186502 2.552e-09 1.694261668963809 2.5529999999999998e-09 1.7735710349323233 2.554e-09 1.8280683140103824 2.555e-09 1.8206389378741252 2.556e-09 1.8272892067368482 2.5569999999999998e-09 1.7985331459869662 2.558e-09 1.7887420940330199 2.559e-09 1.8284874493155676 2.56e-09 1.825891110212258 2.561e-09 1.7272751548429903 2.562e-09 1.8284707913496685 2.563e-09 1.8020714275892187 2.564e-09 1.7673035681794018 2.565e-09 1.7417155249611327 2.566e-09 1.809604306119507 2.567e-09 1.9252136696218418 2.568e-09 1.7440846811116266 2.569e-09 1.767762371406903 2.57e-09 1.812991701452817 2.571e-09 1.8239828063001278 2.572e-09 1.7507663123893895 2.573e-09 1.8071238433685528 2.574e-09 1.790302884512692 2.575e-09 1.8257126895435603 2.5759999999999998e-09 1.7967415987897468 2.577e-09 1.8016376180760398 2.578e-09 1.8685943424311402 2.579e-09 1.8758402291261191 2.5799999999999998e-09 1.7494167564132714 2.581e-09 1.828951435620468 2.582e-09 1.804352407767331 2.583e-09 1.7010505060726986 2.5839999999999998e-09 1.805453069588562 2.585e-09 1.862554529258802 2.586e-09 1.8135832187465688 2.587e-09 1.7846500610611196 2.5879999999999997e-09 1.8263366522354756 2.589e-09 1.8382604452039806 2.59e-09 1.8275180482222324 2.591e-09 1.7682923966942594 2.592e-09 1.7981721818586152 2.593e-09 1.7814130388972038 2.594e-09 1.802457515119435 2.595e-09 1.7637185818280017 2.596e-09 1.712830016559909 2.597e-09 1.8210858960785459 2.598e-09 1.6573440204866747 2.599e-09 1.7607657167460473 2.6e-09 1.8622830816197842 2.601e-09 1.8075987608074664 2.602e-09 1.7811103812610636 2.603e-09 1.8026543101112482 2.604e-09 1.7906910608160034 2.605e-09 1.7925450551712934 2.606e-09 1.7376511616500756 2.6069999999999998e-09 1.7997429361404487 2.608e-09 1.9033610433865416 2.609e-09 1.7883338959366293 2.61e-09 1.8374564537852547 2.6109999999999998e-09 1.7906704253971928 2.612e-09 1.877916209498418 2.613e-09 1.747919801105723 2.614e-09 1.7819713998459155 2.6149999999999998e-09 1.7668142907702489 2.616e-09 1.6811545818354938 2.617e-09 1.7807102106616264 2.618e-09 1.850987978964379 2.6189999999999997e-09 1.8329928651883716 2.62e-09 1.7537662346756189 2.621e-09 1.802543871097833 2.622e-09 1.8356363541845275 2.623e-09 1.7533299277931078 2.624e-09 1.8192378537834355 2.625e-09 1.7796357381833383 2.626e-09 1.7588563437843734 2.627e-09 1.802088042548117 2.628e-09 1.843095291743848 2.629e-09 1.8262123702915285 2.63e-09 1.7492635607428502 2.631e-09 1.8232768262058636 2.632e-09 1.8334897355765638 2.633e-09 1.8189124419781495 2.634e-09 1.8312739942064988 2.635e-09 1.8456003351783228 2.636e-09 1.7847124855814709 2.637e-09 1.87929910548512 2.6379999999999998e-09 1.7921251436372387 2.639e-09 1.7491817793341848 2.64e-09 1.8771166649192388 2.641e-09 1.8792341342809706 2.6419999999999998e-09 1.7963080675746115 2.643e-09 1.688886295307572 2.644e-09 1.77597515609209 2.645e-09 1.7186134053557667 2.6459999999999998e-09 1.72477796092648 2.647e-09 1.9824463836036803 2.648e-09 1.8475294868380239 2.649e-09 1.886910262038694 2.6499999999999997e-09 1.7988984081239714 2.651e-09 1.7978901063238697 2.652e-09 1.8886810367422207 2.653e-09 1.7338303531463874 2.654e-09 1.7603998494291098 2.655e-09 1.7877557228553622 2.656e-09 1.8162613757311994 2.657e-09 1.8113989108161679 2.658e-09 1.792601443749684 2.659e-09 1.817444169241283 2.66e-09 1.73791080387729 2.661e-09 1.8462673180558267 2.662e-09 1.847823988153066 2.663e-09 1.8311649993701622 2.664e-09 1.8401297409939579 2.6649999999999998e-09 1.6942181311589743 2.666e-09 1.7849593454509158 2.667e-09 1.8333572252203463 2.668e-09 1.7511852758854476 2.6689999999999998e-09 1.7868915080610792 2.67e-09 1.7968201578728418 2.671e-09 1.8609198783568581 2.672e-09 1.8530150912755206 2.6729999999999998e-09 1.8477208818697748 2.674e-09 1.7991740095382747 2.675e-09 1.7587732277316688 2.676e-09 1.7453625493938365 2.6769999999999998e-09 1.728060765938144 2.678e-09 1.8636384471425138 2.679e-09 1.763431394736861 2.68e-09 1.7762669441827215 2.681e-09 1.69349669913945 2.682e-09 1.8085704984150872 2.683e-09 1.715662960471639 2.684e-09 1.803444160386408 2.685e-09 1.809397981425202 2.686e-09 1.7486604124034884 2.687e-09 1.7139927795093195 2.688e-09 1.7948625166614738 2.689e-09 1.7739632327848103 2.69e-09 1.8179846022449397 2.691e-09 1.7913393910576894 2.692e-09 1.8082440500520527 2.693e-09 1.818110122577521 2.694e-09 1.7819003921302654 2.695e-09 1.8565276422188248 2.6959999999999998e-09 1.8005317481379006 2.697e-09 1.8525978228169622 2.698e-09 1.7648730277187823 2.699e-09 1.7899015153788136 2.6999999999999998e-09 1.7367827986678495 2.701e-09 1.7490062513535418 2.702e-09 1.6495537839320746 2.703e-09 1.7506331781883457 2.7039999999999998e-09 1.7441517625266818 2.705e-09 1.7613943934398892 2.706e-09 1.6966318392103885 2.707e-09 1.760815537106267 2.7079999999999997e-09 1.7973359009545364 2.709e-09 1.779177137885347 2.71e-09 1.7771785250423258 2.711e-09 1.7967821358053648 2.712e-09 1.8082798865351533 2.713e-09 1.8239705232079868 2.714e-09 1.7783362698325718 2.715e-09 1.7994508277104573 2.716e-09 1.8721830643438324 2.717e-09 1.9333034939980238 2.718e-09 1.840914039200379 2.719e-09 1.8184969430011766 2.72e-09 1.7880121673125056 2.721e-09 1.8296888931935613 2.722e-09 1.847212159814374 2.723e-09 1.8311320984690684 2.724e-09 1.805027412354843 2.725e-09 1.7929205827650985 2.726e-09 1.856179603216756 2.7269999999999998e-09 1.8315905068896363 2.728e-09 1.6821726008616473 2.729e-09 1.7689587659859243 2.73e-09 1.757118488455099 2.7309999999999998e-09 1.7927157808453171 2.732e-09 1.8089422402507127 2.733e-09 1.8587866343370756 2.734e-09 1.7694460977261661 2.7349999999999998e-09 1.7574819073064585 2.736e-09 1.8258493513104086 2.737e-09 1.825712094977645 2.738e-09 1.7556715379710335 2.7389999999999997e-09 1.8464178454372415 2.74e-09 1.8922887881794577 2.741e-09 1.8058805056669247 2.742e-09 1.74770653574237 2.743e-09 1.7707185105134748 2.744e-09 1.7781445026729419 2.745e-09 1.7397878947955567 2.746e-09 1.9378893943766344 2.747e-09 1.8206631648623726 2.748e-09 1.8275447710391277 2.749e-09 1.8436162894286463 2.75e-09 1.733459557621244 2.751e-09 1.8771672330410858 2.752e-09 1.7629525447800556 2.753e-09 1.9038634111678474 2.754e-09 1.6640362738708305 2.755e-09 1.7281591667876608 2.756e-09 1.844336324288649 2.757e-09 1.840992365297963 2.7579999999999998e-09 1.7444208812910669 2.759e-09 1.8773189464423965 2.76e-09 1.8425013868651525 2.761e-09 1.8830863186192244 2.7619999999999998e-09 1.8566770440806935 2.763e-09 1.8638107631134524 2.764e-09 1.7757811879249126 2.765e-09 1.7570873486776653 2.7659999999999998e-09 1.7953174533630663 2.767e-09 1.765022990188681 2.768e-09 1.830164784715833 2.769e-09 1.763067516221333 2.7699999999999997e-09 1.8842212326970031 2.771e-09 1.8390634086178634 2.772e-09 1.747873738613765 2.773e-09 1.9592527424872022 2.774e-09 1.829378780389506 2.775e-09 1.7991751434312073 2.776e-09 1.7823845338782398 2.777e-09 1.836773011130522 2.778e-09 1.742175014209424 2.779e-09 1.7991164463630778 2.78e-09 1.87987916440562 2.781e-09 1.7669283117477 2.782e-09 1.7840861260485446 2.783e-09 1.9368918814247038 2.784e-09 1.8010291068678668 2.7849999999999998e-09 1.8182553812557956 2.786e-09 1.7802402706286928 2.787e-09 1.8041711860104706 2.788e-09 1.8442204591698421 2.7889999999999998e-09 1.7709661737964009 2.79e-09 1.7210233586714094 2.791e-09 1.79085751234317 2.792e-09 1.780191141839042 2.7929999999999998e-09 1.895769231631867 2.794e-09 1.7850787309666392 2.795e-09 1.668526209646838 2.796e-09 1.8292206054335847 2.7969999999999998e-09 1.7703107757307157 2.798e-09 1.7887416132187057 2.799e-09 1.79674146976519 2.8e-09 1.8468047287722096 2.801e-09 1.7910423049191417 2.802e-09 1.7679690408541993 2.803e-09 1.738310940400254 2.804e-09 1.8175634647657177 2.805e-09 1.88761695979015 2.806e-09 1.8076748516908627 2.807e-09 1.790815385173336 2.808e-09 1.735355795793046 2.809e-09 1.8231180255566126 2.81e-09 1.8005955224409653 2.811e-09 1.8069534285480224 2.812e-09 1.8363004182577605 2.813e-09 1.7656493526850316 2.814e-09 1.7548810678418079 2.815e-09 1.762635636096989 2.8159999999999998e-09 1.809729376787982 2.817e-09 1.725003399596277 2.818e-09 1.7780673845214061 2.819e-09 1.7967062200396873 2.8199999999999998e-09 1.7371531320386822 2.821e-09 1.7343131111016452 2.822e-09 1.7968469778367888 2.823e-09 1.7907009098128293 2.8239999999999998e-09 1.798647542803194 2.825e-09 1.770213340667814 2.826e-09 1.8689375184124253 2.827e-09 1.829697347246172 2.8279999999999997e-09 1.7754590041406375 2.829e-09 1.8471542690803906 2.83e-09 1.8671268194629662 2.831e-09 1.757096930087309 2.832e-09 1.7189329850952075 2.833e-09 1.788678401803349 2.834e-09 1.806106903947638 2.835e-09 1.8089738867243264 2.836e-09 1.7054210139424997 2.837e-09 1.870887572646218 2.838e-09 1.8689559282027262 2.839e-09 1.8843191361748282 2.84e-09 1.9101539527601212 2.841e-09 1.7939525831270324 2.842e-09 1.7287993541503657 2.843e-09 1.8029583400309082 2.844e-09 1.7497019902252542 2.845e-09 1.754008767954352 2.846e-09 1.7709107327017546 2.8469999999999998e-09 1.785720691520198 2.848e-09 1.7438529733753718 2.849e-09 1.7338176575902196 2.85e-09 1.7986465402258893 2.8509999999999998e-09 1.8390209433901852 2.852e-09 1.7925695004932005 2.853e-09 1.7671259663724956 2.854e-09 1.746339152079205 2.8549999999999998e-09 1.7237479742881028 2.856e-09 1.7920967565350951 2.857e-09 1.8155878093139177 2.858e-09 1.7726464883573114 2.8589999999999997e-09 1.8937861724665186 2.86e-09 1.733371577398758 2.861e-09 1.7465395267748292 2.862e-09 1.685187428527627 2.863e-09 1.722381121722338 2.864e-09 1.7832839088425978 2.865e-09 1.7591338656208377 2.866e-09 1.8110677336683103 2.867e-09 1.7771207836941834 2.868e-09 1.884984616075706 2.869e-09 1.7593823333463208 2.87e-09 1.829071659646377 2.871e-09 1.9325558268507306 2.872e-09 1.7948866843938487 2.873e-09 1.7276102305226206 2.874e-09 1.8568990291574703 2.875e-09 1.6952747136367863 2.876e-09 1.7538090562586142 2.877e-09 1.8128308723550168 2.8779999999999998e-09 1.7935723468874663 2.879e-09 1.6795409967496737 2.88e-09 1.8509251887686515 2.881e-09 1.8025495090067911 2.8819999999999998e-09 1.7565426035486251 2.883e-09 1.6883754095868233 2.884e-09 1.7800983699596917 2.885e-09 1.8383901725722982 2.8859999999999998e-09 1.7840421513004197 2.887e-09 1.793816373945527 2.888e-09 1.8061606773557777 2.889e-09 1.6826831990776838 2.8899999999999997e-09 1.7883330465843508 2.891e-09 1.8160546793270373 2.892e-09 1.8016944616187076 2.893e-09 1.7237465438243926 2.894e-09 1.7359326165771591 2.895e-09 1.8719025096135868 2.896e-09 1.8038766432146607 2.897e-09 1.8018582723846155 2.898e-09 1.6765687683552748 2.899e-09 1.797584739910605 2.9e-09 1.8049019301248 2.901e-09 1.7541389297897847 2.902e-09 1.8513530369706301 2.903e-09 1.8114862215825958 2.904e-09 1.7839538631220124 2.9049999999999998e-09 1.745093833233442 2.906e-09 1.8031502013547094 2.907e-09 1.7889098384904973 2.908e-09 1.8126700582134956 2.9089999999999998e-09 1.7818140281547141 2.91e-09 1.7851880916945917 2.911e-09 1.7777230584039094 2.912e-09 1.8617331582813592 2.9129999999999998e-09 1.953903806374917 2.914e-09 1.8317260264225574 2.915e-09 1.7991088401646897 2.916e-09 1.7879714086905745 2.9169999999999997e-09 1.7301538862130061 2.918e-09 1.815078251241026 2.919e-09 1.7788370984707156 2.92e-09 1.8023397048128174 2.9209999999999997e-09 1.7341194085954066 2.922e-09 1.8872068620101845 2.923e-09 1.7768795311456111 2.924e-09 1.7469248209804966 2.925e-09 1.8167042519169148 2.926e-09 1.8417847594203127 2.927e-09 1.842089496287075 2.928e-09 1.8900374329234577 2.929e-09 1.694362092103613 2.93e-09 1.782036484035169 2.931e-09 1.6979851168026812 2.932e-09 1.873655364211434 2.933e-09 1.7401372068214858 2.934e-09 1.77081678194371 2.935e-09 1.8516066898568424 2.9359999999999998e-09 1.818276700876479 2.937e-09 1.8300276451444062 2.938e-09 1.7546071503418166 2.939e-09 1.7869001211766504 2.9399999999999998e-09 1.7629573695697698 2.941e-09 1.791831287547866 2.942e-09 1.8025030495878174 2.943e-09 1.8453928774385764 2.9439999999999998e-09 1.7153852683550237 2.945e-09 1.7700871458666365 2.946e-09 1.8647343892262183 2.947e-09 1.7888195944965497 2.9479999999999997e-09 1.7146990912224136 2.949e-09 1.775725770077302 2.95e-09 1.8752564893941672 2.951e-09 1.763562763221654 2.952e-09 1.809755835507349 2.953e-09 1.7519560438764743 2.954e-09 1.8106586204528325 2.955e-09 1.8339131351712337 2.956e-09 1.7097425316705166 2.957e-09 1.7949616898439715 2.958e-09 1.8247830546955492 2.959e-09 1.7230989636037066 2.96e-09 1.787122332696018 2.961e-09 1.9187397411030327 2.962e-09 1.8523032332923224 2.963e-09 1.8754029433455859 2.964e-09 1.7549725787254893 2.965e-09 1.77252324178208 2.966e-09 1.9019338449669851 2.9669999999999998e-09 1.744832842682007 2.968e-09 1.8650865806021186 2.969e-09 1.8183042113059769 2.97e-09 1.8631604774454604 2.9709999999999998e-09 1.8118337086804388 2.972e-09 1.7969086929354487 2.973e-09 1.8387387313536752 2.974e-09 1.8587123339894691 2.9749999999999998e-09 1.7808539712770695 2.976e-09 1.8431615804361163 2.977e-09 1.7062462722785916 2.978e-09 1.7694476896521367 2.9789999999999997e-09 1.7977396929480587 2.98e-09 1.7432392672842258 2.981e-09 1.7643269442262137 2.982e-09 1.8126989369775273 2.983e-09 1.6839550581367644 2.984e-09 1.6983287485307752 2.985e-09 1.768125557131666 2.986e-09 1.7115348747527936 2.987e-09 1.7416179920232189 2.988e-09 1.8323785552298257 2.989e-09 1.8267927068865764 2.99e-09 1.7064017327137677 2.991e-09 1.7941724934688847 2.992e-09 1.7493145546949915 2.993e-09 1.6808148691114357 2.994e-09 1.7535524790052488 2.995e-09 1.8051438820129435 2.996e-09 1.8356005763988343 2.997e-09 1.8495880759481236 2.9979999999999998e-09 1.7219273561906188 2.999e-09 1.8162513364189947 3e-09 1.811115815468916 3.001e-09 1.7440379232956436 3.0019999999999998e-09 1.7961708012571975 3.003e-09 1.795941472955051 3.004e-09 1.8668777717869025 3.005e-09 1.76212871447922 3.0059999999999998e-09 1.7433998561203443 3.007e-09 1.7904860767040225 3.008e-09 1.8127767984312892 3.009e-09 1.818971593611682 3.0099999999999997e-09 1.7662182340868466 3.011e-09 1.8374347992628797 3.012e-09 1.7977609693213599 3.013e-09 1.7982350813371084 3.014e-09 1.8692518973401424 3.015e-09 1.728755047652152 3.016e-09 1.760932203988584 3.017e-09 1.7165147845552666 3.018e-09 1.8285484680171578 3.019e-09 1.7923902647601244 3.02e-09 1.671460850522762 3.021e-09 1.8318220675439099 3.022e-09 1.858589652745269 3.023e-09 1.816964689481314 3.024e-09 1.8956383334998468 3.0249999999999998e-09 1.857648718760274 3.026e-09 1.7769473925974528 3.027e-09 1.8263646586601747 3.028e-09 1.7850257978938882 3.0289999999999998e-09 1.7781154645525667 3.03e-09 1.76727034046967 3.031e-09 1.7784617833997285 3.032e-09 1.7927199274989085 3.0329999999999998e-09 1.7613410818921182 3.034e-09 1.85133744850996 3.035e-09 1.7515620332602795 3.036e-09 1.7953229173833227 3.0369999999999997e-09 1.7788886854848764 3.038e-09 1.7381416414378748 3.039e-09 1.7718793671661497 3.04e-09 1.6619519773795084 3.0409999999999997e-09 1.675235707380064 3.042e-09 1.7884349072204895 3.043e-09 1.7954123577808667 3.044e-09 1.7632902794443004 3.045e-09 1.7944649962887642 3.046e-09 1.8888524319114706 3.047e-09 1.7503382774877876 3.048e-09 1.7880420615053472 3.049e-09 1.8634713380313963 3.05e-09 1.8200228285048015 3.051e-09 1.7485776850578276 3.052e-09 1.8430906417419362 3.053e-09 1.7668231670164543 3.054e-09 1.7737623582490027 3.055e-09 1.773272578477332 3.0559999999999998e-09 1.7841329131733503 3.057e-09 1.9332698052638266 3.058e-09 1.6990561729647886 3.059e-09 1.8615290119296382 3.0599999999999998e-09 1.8576336935718056 3.061e-09 1.8372243636800838 3.062e-09 1.8372067714405986 3.063e-09 1.7648797074101188 3.0639999999999998e-09 1.8552498042220975 3.065e-09 1.8029188546133157 3.066e-09 1.8093878545352802 3.067e-09 1.792264125057625 3.0679999999999997e-09 1.815704081529921 3.069e-09 1.8611497473299141 3.07e-09 1.7464860062700518 3.071e-09 1.7818175637749292 3.072e-09 1.7031488193337734 3.073e-09 1.8179145126604743 3.074e-09 1.7143464829855666 3.075e-09 1.9057534133373273 3.076e-09 1.8365284578861265 3.077e-09 1.8140005129059487 3.078e-09 1.83991062820114 3.079e-09 1.8405456856006648 3.08e-09 1.8461977965604168 3.081e-09 1.747170933209969 3.082e-09 1.8230763793473386 3.083e-09 1.7448557844824513 3.084e-09 1.8023104617066739 3.085e-09 1.8105230004127573 3.086e-09 1.7726630633073663 3.0869999999999998e-09 1.8662023510100423 3.088e-09 1.8413528630947888 3.089e-09 1.8286155284351924 3.09e-09 1.8639641776026334 3.0909999999999998e-09 1.786579249664621 3.092e-09 1.7870308985004397 3.093e-09 1.79419944371866 3.094e-09 1.932414186683717 3.0949999999999998e-09 1.7569252763920458 3.096e-09 1.7949800840758312 3.097e-09 1.840364226542119 3.098e-09 1.8635669908360386 3.0989999999999997e-09 1.8512255857098923 3.1e-09 1.7232511657018061 3.101e-09 1.8265234419036296 3.102e-09 1.7257476219956487 3.103e-09 1.8062309030649402 3.104e-09 1.772852461377987 3.105e-09 1.7669219513077234 3.106e-09 1.7773762912203688 3.107e-09 1.7416600080793456 3.108e-09 1.7665861998288326 3.109e-09 1.739307141282028 3.11e-09 1.8368292884627693 3.111e-09 1.86171389058052 3.112e-09 1.8608856959295645 3.113e-09 1.7101061788800922 3.1139999999999998e-09 1.8191522246221017 3.115e-09 1.7008932675819328 3.116e-09 1.715783041007146 3.117e-09 1.7824816886872932 3.1179999999999998e-09 1.8035219211816236 3.119e-09 1.7591210687974086 3.12e-09 1.8186295161113557 3.121e-09 1.7680902227273476 3.1219999999999998e-09 1.7859141593327157 3.123e-09 1.7852460530474932 3.124e-09 1.6773660119629112 3.125e-09 1.7895639497194828 3.1259999999999998e-09 1.8516335200538736 3.127e-09 1.8276933024069115 3.128e-09 1.7907090211449141 3.129e-09 1.8073239696363161 3.1299999999999997e-09 1.8450719989638975 3.131e-09 1.804491159073198 3.132e-09 1.8583145273312096 3.133e-09 1.8099110032287287 3.134e-09 1.7865938490989015 3.135e-09 1.794440094993333 3.136e-09 1.8615372886336068 3.137e-09 1.7457451909141277 3.138e-09 1.82455999014401 3.139e-09 1.8164538137121462 3.14e-09 1.8766911302937215 3.141e-09 1.8023884501242748 3.142e-09 1.7881782668837995 3.143e-09 1.7334160554882505 3.144e-09 1.8573419988419342 3.1449999999999998e-09 1.7638681565750842 3.146e-09 1.820028530141227 3.147e-09 1.904173895830071 3.148e-09 1.820039494325106 3.1489999999999998e-09 1.8286294999812958 3.15e-09 1.7849402124335223 3.151e-09 1.7968948741274273 3.152e-09 1.8106553727812758 3.1529999999999998e-09 1.735769489732352 3.154e-09 1.725279036716107 3.155e-09 1.8699803536595294 3.156e-09 1.8373765828557167 3.1569999999999997e-09 1.7647209842479545 3.158e-09 1.8157762481858672 3.159e-09 1.7718866558961075 3.16e-09 1.8201891467914477 3.1609999999999997e-09 1.7662633646110155 3.162e-09 1.8659760674276504 3.163e-09 1.701164396015645 3.164e-09 1.839775066535964 3.165e-09 1.8219142641608905 3.166e-09 1.7766115291230264 3.167e-09 1.7798644335406268 3.168e-09 1.6698443289009828 3.169e-09 1.8407927703465523 3.17e-09 1.7669675495441297 3.171e-09 1.799307151099093 3.172e-09 1.716933461643865 3.173e-09 1.809974910012526 3.174e-09 1.7415710980774277 3.175e-09 1.696191820174041 3.1759999999999998e-09 1.8445167962942723 3.177e-09 1.7475688298948837 3.178e-09 1.743390157196683 3.179e-09 1.8617574720981342 3.1799999999999998e-09 1.8232515010881227 3.181e-09 1.8880557578622719 3.182e-09 1.7792422987021932 3.183e-09 1.7933199087362033 3.1839999999999998e-09 1.8070552312555566 3.185e-09 1.7666758589022056 3.186e-09 1.7610758391848982 3.187e-09 1.8157716948607754 3.1879999999999997e-09 1.863434911357046 3.189e-09 1.8979179890770714 3.19e-09 1.8835420027832834 3.191e-09 1.7467260584769526 3.1919999999999997e-09 1.759597975138921 3.193e-09 1.8130791798309647 3.194e-09 1.7983495496881434 3.195e-09 1.7592332463610683 3.196e-09 1.8200731114775577 3.197e-09 1.8473438331574148 3.198e-09 1.8222077848910847 3.199e-09 1.7604584074510072 3.2e-09 1.7956273499352389 3.201e-09 1.7636231758195977 3.202e-09 1.7729651877257153 3.203e-09 1.830922242487647 3.204e-09 1.7780837945352335 3.205e-09 1.7771208773138878 3.206e-09 1.8751940864582177 3.2069999999999998e-09 1.7119568763579145 3.208e-09 1.8321126788074218 3.209e-09 1.7801427688850269 3.21e-09 1.836732392614006 3.2109999999999998e-09 1.7669690071650745 3.212e-09 1.7722827929300562 3.213e-09 1.7721569466432963 3.214e-09 1.7804960891380537 3.2149999999999998e-09 1.801551923119656 3.216e-09 1.9441644849655892 3.217e-09 1.790743733809249 3.218e-09 1.6699272753728105 3.2189999999999997e-09 1.7894719790324787 3.22e-09 1.8054996013301265 3.221e-09 1.8202628823556077 3.222e-09 1.738045531062031 3.223e-09 1.8150331570796823 3.224e-09 1.8163299967528508 3.225e-09 1.8531031010494448 3.226e-09 1.763596281097906 3.227e-09 1.7793488495099163 3.228e-09 1.7593207694081914 3.229e-09 1.809187682514002 3.23e-09 1.8952255912569318 3.231e-09 1.7392010435388325 3.232e-09 1.7611997434657172 3.233e-09 1.8804378963062731 3.2339999999999998e-09 1.845987706030885 3.235e-09 1.8350205519221996 3.236e-09 1.807009712219422 3.237e-09 1.8436731355004579 3.2379999999999998e-09 1.8083084180362496 3.239e-09 1.7792377915826454 3.24e-09 1.7408315652170099 3.241e-09 1.8632526744965707 3.2419999999999998e-09 1.8608367394391467 3.243e-09 1.797497063844761 3.244e-09 1.8154824023302376 3.245e-09 1.6989370274880309 3.2459999999999998e-09 1.8027355897898365 3.247e-09 1.8489531341632828 3.248e-09 1.751883652817323 3.249e-09 1.7550332217726228 3.2499999999999997e-09 1.7940430661105262 3.251e-09 1.7373518817927123 3.252e-09 1.8628130998570624 3.253e-09 1.8824997212853831 3.254e-09 1.7531569982072372 3.255e-09 1.8246257042336258 3.256e-09 1.7928065271401161 3.257e-09 1.8049655075366424 3.258e-09 1.82947585519907 3.259e-09 1.8027769345644007 3.26e-09 1.8043738504844387 3.261e-09 1.8120464633845226 3.262e-09 1.7583118149480477 3.263e-09 1.8173656487584042 3.264e-09 1.835952588079555 3.2649999999999998e-09 1.9287118407091193 3.266e-09 1.811592063655109 3.267e-09 1.7685414008597615 3.268e-09 1.7967951776256474 3.2689999999999998e-09 1.8177683319794886 3.27e-09 1.8158580242081135 3.271e-09 1.8911763041113083 3.272e-09 1.887124780059019 3.2729999999999998e-09 1.7945350022372666 3.274e-09 1.860182600346373 3.275e-09 1.7463000665847437 3.276e-09 1.7592938918494705 3.2769999999999997e-09 1.809177232904869 3.278e-09 1.7585004916272577 3.279e-09 1.8842302978678214 3.28e-09 1.8524495691959146 3.2809999999999997e-09 1.8025664541213966 3.282e-09 1.844756878057554 3.283e-09 1.842506122895859 3.284e-09 1.7631469887702051 3.285e-09 1.8478761769094865 3.286e-09 1.828028146957185 3.287e-09 1.8276702683818247 3.288e-09 1.7136644724933663 3.289e-09 1.8342772551701967 3.29e-09 1.8015694708114725 3.291e-09 1.7559139251222973 3.292e-09 1.758357728911282 3.293e-09 1.6936560439821433 3.294e-09 1.8594710214548105 3.295e-09 1.719825171241915 3.2959999999999998e-09 1.79873958450849 3.297e-09 1.8813987016931601 3.298e-09 1.7214678787761315 3.299e-09 1.779372234616311 3.2999999999999998e-09 1.8107049976801166 3.301e-09 1.8472284858251244 3.302e-09 1.766699006002537 3.303e-09 1.8378089117989782 3.3039999999999998e-09 1.8296959490741445 3.305e-09 1.8151931869630247 3.306e-09 1.811390083594042 3.307e-09 1.763395158066241 3.3079999999999997e-09 1.812445935190732 3.309e-09 1.7119459063808917 3.31e-09 1.7764399538794635 3.311e-09 1.9225599414758716 3.3119999999999997e-09 1.8507623915543594 3.313e-09 1.8357240272010347 3.314e-09 1.7756644226004212 3.315e-09 1.7573018079298393 3.316e-09 1.793669615330178 3.317e-09 1.7230907226711762 3.318e-09 1.8221177672540942 3.319e-09 1.7784089377306667 3.32e-09 1.859850604482811 3.321e-09 1.7824621124200803 3.322e-09 1.7636914854944046 3.323e-09 1.7793338812426225 3.324e-09 1.82765347520753 3.325e-09 1.7356985809558971 3.326e-09 1.7532304725814618 3.3269999999999998e-09 1.8286878189310154 3.328e-09 1.8244468990930536 3.329e-09 1.8231005109239449 3.33e-09 1.7938158873086674 3.3309999999999998e-09 1.8457551925040863 3.332e-09 1.786556863432691 3.333e-09 1.8123944317967824 3.334e-09 1.7805927778621047 3.3349999999999998e-09 1.7160051660510884 3.336e-09 1.7347454802166324 3.337e-09 1.8401315739479593 3.338e-09 1.77763439592071 3.3389999999999997e-09 1.7993267790850764 3.34e-09 1.7441009795205915 3.341e-09 1.7722248313476239 3.342e-09 1.8085968891924356 3.3429999999999997e-09 1.7912536228884814 3.344e-09 1.7296743708407545 3.345e-09 1.8494123716443847 3.346e-09 1.7526420737185324 3.347e-09 1.8387472064771873 3.348e-09 1.8017101894799432 3.349e-09 1.7387787930421328 3.35e-09 1.7493821560542073 3.351e-09 1.8492637435095525 3.352e-09 1.8085569816205402 3.353e-09 1.8756864080941253 3.3539999999999998e-09 1.8442214270383408 3.355e-09 1.8072547570124078 3.356e-09 1.7423311594769508 3.357e-09 1.8026862457151918 3.3579999999999998e-09 1.7200220452356407 3.359e-09 1.8199780111188564 3.36e-09 1.7699202527499835 3.361e-09 1.8007464464029102 3.3619999999999998e-09 1.8582759625850755 3.363e-09 1.735676124853503 3.364e-09 1.724729536102189 3.365e-09 1.760702236676487 3.3659999999999998e-09 1.8734331608209627 3.367e-09 1.834131200984706 3.368e-09 1.7507205210574286 3.369e-09 1.7491850815469485 3.3699999999999997e-09 1.7951863848132876 3.371e-09 1.8087583424422322 3.372e-09 1.7557303658871193 3.373e-09 1.7757577017685064 3.374e-09 1.8209430073028334 3.375e-09 1.8654287780870618 3.376e-09 1.8200905407707093 3.377e-09 1.7933256188138276 3.378e-09 1.756666391306566 3.379e-09 1.7886836198126845 3.38e-09 1.7428170673353076 3.381e-09 1.7152178833141754 3.382e-09 1.8875806471544723 3.383e-09 1.7983318080678445 3.384e-09 1.779161336197495 3.3849999999999998e-09 1.819933066405229 3.386e-09 1.773429168384406 3.387e-09 1.830438142549779 3.388e-09 1.7823587123196423 3.3889999999999998e-09 1.8159948338145289 3.39e-09 1.8600915525267363 3.391e-09 1.7468384984945917 3.392e-09 1.8258106338754911 3.3929999999999998e-09 1.853594950683208 3.394e-09 1.8406963730386037 3.395e-09 1.8160041824477597 3.396e-09 1.7985420476839726 3.3969999999999997e-09 1.758544044167784 3.398e-09 1.7927283488607613 3.399e-09 1.7942033992934705 3.4e-09 1.7873179410485707 3.4009999999999997e-09 1.7351267969586808 3.402e-09 1.7658577831431521 3.403e-09 1.7789346297289599 3.404e-09 1.788792393043495 3.405e-09 1.7667233155559527 3.406e-09 1.7292466180312187 3.407e-09 1.8020154021898622 3.408e-09 1.8153135318067224 3.409e-09 1.8268993396714537 3.41e-09 1.8144661117823297 3.411e-09 1.6657124548604012 3.412e-09 1.815429614742632 3.413e-09 1.808834891916839 3.414e-09 1.8127856424586002 3.415e-09 1.8269781188380694 3.4159999999999998e-09 1.8449693248704289 3.417e-09 1.8276179269835915 3.418e-09 1.6467161544677784 3.419e-09 1.905609764720312 3.4199999999999998e-09 1.869012345887835 3.421e-09 1.846145788484033 3.422e-09 1.8490144833189184 3.423e-09 1.7654175124108187 3.4239999999999998e-09 1.7223396903404993 3.425e-09 1.8096272824035495 3.426e-09 1.8123688108992413 3.427e-09 1.7449003204036768 3.4279999999999997e-09 1.843017800415538 3.429e-09 1.7955448584985618 3.43e-09 1.7713254339192366 3.431e-09 1.9067992471278126 3.4319999999999997e-09 1.7225539622126096 3.433e-09 1.9100861323674914 3.434e-09 1.7117159491099851 3.435e-09 1.842403469522921 3.436e-09 1.8023433345190563 3.437e-09 1.8620328448184635 3.438e-09 1.785266988449143 3.439e-09 1.8335371105615657 3.44e-09 1.8124087033550191 3.441e-09 1.8484059751751565 3.442e-09 1.7852061390538554 3.443e-09 1.8291046072233275 3.444e-09 1.72551910703472 3.445e-09 1.7383514122203676 3.446e-09 1.8341222870876006 3.4469999999999998e-09 1.7486526443343187 3.448e-09 1.809599169930952 3.449e-09 1.8092533637826453 3.45e-09 1.8275998779334726 3.4509999999999998e-09 1.8250930837937607 3.452e-09 1.8770901535541005 3.453e-09 1.732202921820394 3.454e-09 1.7223754953461077 3.4549999999999998e-09 1.789356734211426 3.456e-09 1.7951962592062645 3.457e-09 1.8025741414680243 3.458e-09 1.769329063197494 3.4589999999999997e-09 1.817165380979011 3.46e-09 1.7457012008726827 3.461e-09 1.8720726979707425 3.462e-09 1.7822503310295938 3.4629999999999997e-09 1.7898290580863814 3.464e-09 1.7081953204183393 3.465e-09 1.8065609544473649 3.466e-09 1.7238171399729694 3.467e-09 1.7972601067047578 3.468e-09 1.7951722613781944 3.469e-09 1.749858508583496 3.47e-09 1.765969749140841 3.471e-09 1.8074190661604863 3.472e-09 1.8078888467079264 3.473e-09 1.8325684982783272 3.4739999999999998e-09 1.755993038172448 3.475e-09 1.8084695425790518 3.476e-09 1.8354828746273886 3.477e-09 1.7597693349631642 3.4779999999999998e-09 1.8656123002885827 3.479e-09 1.8291502547290033 3.48e-09 1.8702170882892148 3.481e-09 1.7559803326433112 3.4819999999999998e-09 1.8072975116245336 3.483e-09 1.7859581911457683 3.484e-09 1.7078458284507223 3.485e-09 1.8810958886444415 3.4859999999999997e-09 1.7575522994971746 3.487e-09 1.6702706482953533 3.488e-09 1.815229850579632 3.489e-09 1.7975386879222541 3.4899999999999997e-09 1.6479308064650804 3.491e-09 1.8119787658253659 3.492e-09 1.792705537257539 3.493e-09 1.747343109559249 3.494e-09 1.802181929802624 3.495e-09 1.7984891604462478 3.496e-09 1.7894017772186106 3.497e-09 1.847039100055053 3.498e-09 1.7995962456131007 3.499e-09 1.8009228093525864 3.5e-09 1.7411875077507648 3.501e-09 1.8427003552239913 3.502e-09 1.8140430964496752 3.503e-09 1.7807531922694466 3.504e-09 1.7992181319714708 3.5049999999999998e-09 1.8079431795961116 3.506e-09 1.8124249515332584 3.507e-09 1.8640529757218813 3.508e-09 1.7869735008829912 3.5089999999999998e-09 1.8324500339797747 3.51e-09 1.8449564675503702 3.511e-09 1.7732474088952088 3.512e-09 1.698124733875834 3.5129999999999998e-09 1.7918416085171358 3.514e-09 1.8721881764375072 3.515e-09 1.7474458883010056 3.516e-09 1.8303849642705834 3.5169999999999997e-09 1.7797506923223603 3.518e-09 1.8348509035741893 3.519e-09 1.8290006551538482 3.52e-09 1.714079377311601 3.5209999999999997e-09 1.7762170376564628 3.522e-09 1.7098023725565326 3.523e-09 1.7089160346871113 3.524e-09 1.84773018189305 3.525e-09 1.7855442224525304 3.526e-09 1.791255727235488 3.527e-09 1.8028123401169325 3.528e-09 1.785743541634033 3.529e-09 1.7510467420312137 3.53e-09 1.8701648972075404 3.531e-09 1.7389739422311563 3.532e-09 1.7774943951308289 3.533e-09 1.8399067110610277 3.534e-09 1.7733126570983504 3.535e-09 1.7826676015153256 3.5359999999999998e-09 1.7889847485088526 3.537e-09 1.8641377329788098 3.538e-09 1.8319887567854707 3.539e-09 1.8258894730832456 3.5399999999999998e-09 1.7883661557962478 3.541e-09 1.8462703544884167 3.542e-09 1.7791082704358636 3.543e-09 1.7807805336303224 3.5439999999999998e-09 1.8171985804865816 3.545e-09 1.7110574109237537 3.546e-09 1.8167178378953193 3.547e-09 1.7374033491700016 3.5479999999999997e-09 1.8092385208718789 3.549e-09 1.823892207353997 3.55e-09 1.813062279908793 3.551e-09 1.8539100700682092 3.5519999999999997e-09 1.8709876166599186 3.553e-09 1.7798224926692734 3.554e-09 1.7830332046483814 3.555e-09 1.7698206858169827 3.556e-09 1.7815282437683015 3.557e-09 1.795671085139874 3.558e-09 1.7971971647176157 3.559e-09 1.8906127262033428 3.56e-09 1.7927411759251504 3.561e-09 1.8298951314208332 3.562e-09 1.7714153508300423 3.563e-09 1.7568016945016065 3.564e-09 1.8760302812006557 3.565e-09 1.8010296379050548 3.566e-09 1.775092769828142 3.5669999999999998e-09 1.750022240633148 3.568e-09 1.7580174299084501 3.569e-09 1.7522554551708758 3.57e-09 1.7857208106556426 3.5709999999999998e-09 1.8608147607907561 3.572e-09 1.7927128229182303 3.573e-09 1.8041201407184864 3.574e-09 1.7573137918315402 3.5749999999999998e-09 1.8032667014968196 3.576e-09 1.7572585397908256 3.577e-09 1.8216188093066885 3.578e-09 1.7993029592683354 3.5789999999999997e-09 1.7902501661729733 3.58e-09 1.884632870477362 3.581e-09 1.7487097061896297 3.582e-09 1.836157841263605 3.5829999999999997e-09 1.7732855665272036 3.584e-09 1.8598466949182995 3.585e-09 1.7592213430839927 3.586e-09 1.7651637077913551 3.587e-09 1.8205423518611539 3.588e-09 1.7461971603968485 3.589e-09 1.7620401369854162 3.59e-09 1.758928034284252 3.591e-09 1.8994060030166757 3.592e-09 1.7770414853504928 3.593e-09 1.829621360372261 3.5939999999999998e-09 1.7813587594285483 3.595e-09 1.760138404213168 3.596e-09 1.807915346257874 3.597e-09 1.6905198742116478 3.5979999999999998e-09 1.7453404057489803 3.599e-09 1.786478463721993 3.6e-09 1.7675539968807112 3.601e-09 1.8844063592710547 3.6019999999999998e-09 1.8112084090975213 3.603e-09 1.7717688346600708 3.604e-09 1.8099311858067693 3.605e-09 1.7942652503462166 3.6059999999999997e-09 1.807451734644417 3.607e-09 1.777889207591607 3.608e-09 1.829656147958262 3.609e-09 1.868464737975633 3.6099999999999997e-09 1.7929127269230622 3.611e-09 1.8326723409486618 3.612e-09 1.8439335975581528 3.613e-09 1.8809967138288801 3.6139999999999997e-09 1.7729510639280872 3.615e-09 1.7243817589399026 3.616e-09 1.7778990576021507 3.617e-09 1.8339510814562667 3.618e-09 1.7946913302328877 3.619e-09 1.834739587475157 3.62e-09 1.7466041336850942 3.621e-09 1.7810057011344713 3.622e-09 1.8187114840296914 3.623e-09 1.8074747673615186 3.624e-09 1.7151233785702744 3.6249999999999998e-09 1.7963397947904047 3.626e-09 1.8600501082389436 3.627e-09 1.7797660401538073 3.628e-09 1.8484802331869428 3.6289999999999998e-09 1.828766775497511 3.63e-09 1.8361796909898858 3.631e-09 1.7798040161138236 3.632e-09 1.6972548295124301 3.6329999999999998e-09 1.7474616369002234 3.634e-09 1.7531421367140774 3.635e-09 1.8499538636562813 3.636e-09 1.849141679277587 3.6369999999999997e-09 1.823058474008381 3.638e-09 1.6875608543128544 3.639e-09 1.779921625188006 3.64e-09 1.815378601330935 3.6409999999999997e-09 1.7538886123642248 3.642e-09 1.825158064118559 3.643e-09 1.8267655790685402 3.644e-09 1.836931170704424 3.645e-09 1.7338394090343048 3.646e-09 1.8723314437303167 3.647e-09 1.8430551736634155 3.648e-09 1.8565814954287194 3.649e-09 1.7345255925628205 3.65e-09 1.8246307216943465 3.651e-09 1.7649099288451253 3.652e-09 1.834391407020743 3.653e-09 1.7972510189659958 3.654e-09 1.8908226957041974 3.655e-09 1.776632937654221 3.6559999999999998e-09 1.724148651150006 3.657e-09 1.7476013041806564 3.658e-09 1.804879819867458 3.659e-09 1.8636008889661224 3.6599999999999998e-09 1.88266143394082 3.661e-09 1.858268287142797 3.662e-09 1.8348559978509995 3.663e-09 1.8122360656756782 3.6639999999999998e-09 1.8219511018311665 3.665e-09 1.8388895054995071 3.666e-09 1.7805087260367438 3.667e-09 1.815547997452038 3.6679999999999997e-09 1.738997477560798 3.669e-09 1.849861418302576 3.67e-09 1.873267182257988 3.671e-09 1.858059851879275 3.6719999999999997e-09 1.7958148321441365 3.673e-09 1.8000197898073416 3.674e-09 1.8620159932775406 3.675e-09 1.791283517714696 3.676e-09 1.7853642703513755 3.677e-09 1.7649609556057593 3.678e-09 1.86644355240519 3.679e-09 1.8644551639772589 3.68e-09 1.7051170954217205 3.681e-09 1.8084594947064208 3.682e-09 1.8272867732226563 3.6829999999999998e-09 1.8091164844124252 3.684e-09 1.8215687217107708 3.685e-09 1.6982443284223963 3.686e-09 1.8051654533525396 3.6869999999999998e-09 1.838095862964724 3.688e-09 1.7376522538446082 3.689e-09 1.8181111084222032 3.69e-09 1.8451174539114064 3.6909999999999998e-09 1.8404835068772765 3.692e-09 1.8843000974749253 3.693e-09 1.8206316744019282 3.694e-09 1.7403771077944636 3.6949999999999998e-09 1.7924244571531616 3.696e-09 1.8273549743793276 3.697e-09 1.8097018149552662 3.698e-09 1.801147268087807 3.6989999999999997e-09 1.8692640445602167 3.7e-09 1.7608432719236897 3.701e-09 1.9996918025227906 3.702e-09 1.704324934828937 3.7029999999999997e-09 1.816371426662195 3.704e-09 1.814654070296587 3.705e-09 1.822396218965113 3.706e-09 1.8017556058077442 3.707e-09 1.7459825131788393 3.708e-09 1.789574276325932 3.709e-09 1.7860955786663963 3.71e-09 1.8471906727114678 3.711e-09 1.6960722919530091 3.712e-09 1.7728701577563017 3.713e-09 1.8171715268659978 3.7139999999999998e-09 1.8724336791803105 3.715e-09 1.7954704172705185 3.716e-09 1.800417039532943 3.717e-09 1.7926368741986753 3.7179999999999998e-09 1.6894476491881962 3.719e-09 1.8474946038351001 3.72e-09 1.7879458445469985 3.721e-09 1.8068642690193488 3.7219999999999998e-09 1.7320668422143963 3.723e-09 1.8190414520324536 3.724e-09 1.766491467341219 3.725e-09 1.7930383075250258 3.726e-09 1.852687776663013 3.727e-09 1.8441741322130207 3.7279999999999995e-09 1.8195008843173095 3.729e-09 1.7772614288876534 3.73e-09 1.6756278512868992 3.731e-09 1.7186876579225363 3.732e-09 1.8602273668233935 3.733e-09 1.7923215632152036 3.734e-09 1.9462773732343068 3.735e-09 1.849179892751051 3.736e-09 1.7816658241578567 3.737e-09 1.7929947224414293 3.738e-09 1.7766584986673553 3.739e-09 1.7952604872690137 3.74e-09 1.7509048412441084 3.741e-09 1.7743763632722598 3.742e-09 1.8267829594391156 3.743e-09 1.863222089788688 3.744e-09 1.831632396638482 3.745e-09 1.7361704261133497 3.746e-09 1.7467734359040428 3.7469999999999996e-09 1.8054328970217268 3.748e-09 1.8522674134768218 3.749e-09 1.729003631718143 3.75e-09 1.7762559129398707 3.751e-09 1.7270582536697243 3.752e-09 1.8259870345485032 3.753e-09 1.7360166462559967 3.754e-09 1.8368438893191457 3.7549999999999995e-09 1.8792724872862057 3.756e-09 1.784341421123586 3.757e-09 1.804800226579039 3.758e-09 1.7023369119548686 3.759e-09 1.776740213871041 3.76e-09 1.8498284608961395 3.761e-09 1.7642779275794127 3.762e-09 1.8048114714307888 3.7629999999999995e-09 1.7407693603443484 3.764e-09 1.84479845730458 3.765e-09 1.8099458408948028 3.766e-09 1.818348230219536 3.767e-09 1.7660200689139929 3.768e-09 1.8170568327217727 3.769e-09 1.8505073444355933 3.77e-09 1.7450170352930066 3.771e-09 1.888237106341522 3.772e-09 1.834543588181825 3.773e-09 1.8517002428089255 3.7739999999999996e-09 1.792649556574435 3.775e-09 1.6918296680582112 3.776e-09 1.8385632632782865 3.777e-09 1.7798405463538953 3.778e-09 1.8730675285949288 3.779e-09 1.854563396820807 3.78e-09 1.7394052536039661 3.781e-09 1.7217052530207553 3.7819999999999996e-09 1.7387611299278347 3.783e-09 1.8402818420612552 3.784e-09 1.8308416153100084 3.785e-09 1.7997412843513751 3.786e-09 1.7854810263525922 3.787e-09 1.8928322760193501 3.788e-09 1.6575080580939443 3.789e-09 1.8166897851825021 3.7899999999999995e-09 1.728897370731837 3.791e-09 1.8396816237230134 3.792e-09 1.80942106847049 3.793e-09 1.7915693700354736 3.794e-09 1.8131085688991309 3.795e-09 1.6851088807329708 3.796e-09 1.8572983974236095 3.797e-09 1.8539586550234661 3.798e-09 1.765015392427326 3.799e-09 1.8201243911697216 3.8e-09 1.860245665405242 3.801e-09 1.7754514522065707 3.802e-09 1.8976017514199124 3.803e-09 1.8678889299255057 3.804e-09 1.764179665035127 3.805e-09 1.842408890671386 3.806e-09 1.81274388458848 3.807e-09 1.8498532686470983 3.808e-09 1.778649592349076 3.8089999999999996e-09 1.6847912506151907 3.81e-09 1.8021602604774023 3.811e-09 1.7507138372684787 3.812e-09 1.7982008159983698 3.813e-09 1.7630220331027966 3.814e-09 1.7158243998487717 3.815e-09 1.9029702050637076 3.816e-09 1.8065701188815775 3.8169999999999995e-09 1.8823362026641655 3.818e-09 1.7658792016918405 3.819e-09 1.8012651596853522 3.82e-09 1.7413284801021987 3.821e-09 1.887486705413694 3.822e-09 1.7235018462911718 3.823e-09 1.7788070572419434 3.824e-09 1.8097885362814587 3.825e-09 1.8876526786435361 3.826e-09 1.7750730470704768 3.827e-09 1.7601262448234696 3.828e-09 1.8105893668300834 3.829e-09 1.7785435532323546 3.83e-09 1.8142373374707688 3.831e-09 1.7122349317407721 3.832e-09 1.8220106473208197 3.833e-09 1.8707620882246208 3.834e-09 1.784077994057129 3.835e-09 1.6902308129670174 3.8359999999999996e-09 1.837996822754092 3.837e-09 1.8454597466005878 3.838e-09 1.826382955725631 3.839e-09 1.7677198078723009 3.84e-09 1.8237522287083159 3.841e-09 1.895567740717619 3.842e-09 1.8716983192233767 3.843e-09 1.6568544388746156 3.8439999999999995e-09 1.8059841143979407 3.845e-09 1.7906130177630784 3.846e-09 1.8689725923692255 3.847e-09 1.8201042071441678 3.848e-09 1.705695592545631 3.849e-09 1.6793821432231604 3.85e-09 1.7969685499633918 3.851e-09 1.737469025335948 3.8519999999999995e-09 1.7808502930262262 3.853e-09 1.8447160605054522 3.854e-09 1.8377792930183903 3.855e-09 1.7847079287390284 3.856e-09 1.7847257765482392 3.857e-09 1.7506439271081289 3.858e-09 1.8253036383500185 3.859e-09 1.725166442659885 3.86e-09 1.845201199981116 3.861e-09 1.7725804759774977 3.862e-09 1.7544900394805534 3.8629999999999996e-09 1.751988618182105 3.864e-09 1.870308063250762 3.865e-09 1.7995884569641254 3.866e-09 1.7966254893915048 3.867e-09 1.8367760003794684 3.868e-09 1.7718209792783088 3.869e-09 1.8356241327063687 3.87e-09 1.7837760616590856 3.8709999999999996e-09 1.716278789639442 3.872e-09 1.804843692519976 3.873e-09 1.877642447343656 3.874e-09 1.8273711263505845 3.875e-09 1.8482338856800764 3.876e-09 1.8914418754740425 3.877e-09 1.8414920121298544 3.878e-09 1.7894638760238597 3.8789999999999995e-09 1.8015770021350934 3.88e-09 1.7907324660923567 3.881e-09 1.771872761494127 3.882e-09 1.7784200853514314 3.883e-09 1.8255903247437655 3.884e-09 1.7792279840398046 3.885e-09 1.8291794410293813 3.886e-09 1.7378273324788496 3.887e-09 1.7859395501527036 3.888e-09 1.7988103743694257 3.889e-09 1.8102306793257734 3.89e-09 1.7940364987527055 3.891e-09 1.8365545763726383 3.892e-09 1.7802573993749908 3.893e-09 1.8055126847928658 3.894e-09 1.734830348985464 3.895e-09 1.6844302880904345 3.896e-09 1.7426513042379046 3.897e-09 1.7786747405657137 3.8979999999999996e-09 1.7452593604980335 3.899e-09 1.8304149794219733 3.9e-09 1.6985123070627481 3.901e-09 1.7976261092755998 3.902e-09 1.8271833674646838 3.903e-09 1.8019573753352633 3.904e-09 1.8697420798186377 3.905e-09 1.7828826307151378 3.9059999999999995e-09 1.8169825786453784 3.907e-09 1.7399515984035736 3.908e-09 1.8492437531310197 3.909e-09 1.7445073764332004 3.91e-09 1.8161909380775638 3.911e-09 1.735293175555252 3.912e-09 1.756598462033878 3.913e-09 1.78055936233161 3.9139999999999995e-09 1.8516509371263883 3.915e-09 1.8080540721438034 3.916e-09 1.7699155184585114 3.917e-09 1.771221925465838 3.918e-09 1.8316634466490183 3.919e-09 1.7339708682352974 3.92e-09 1.8311936942447704 3.921e-09 1.7964199295452847 3.922e-09 1.779001008627285 3.923e-09 1.836500452952153 3.924e-09 1.914367365265056 3.9249999999999996e-09 1.8142595819076197 3.926e-09 1.8172774212837415 3.927e-09 1.7488399844790998 3.928e-09 1.8952328758111223 3.929e-09 1.8201722066466892 3.93e-09 1.8657243828658623 3.931e-09 1.7437369438574615 3.932e-09 1.8193316607116996 3.9329999999999995e-09 1.750941092795846 3.934e-09 1.7937870883401292 3.935e-09 1.8099612287330844 3.936e-09 1.7759187539017074 3.937e-09 1.8450603579449016 3.938e-09 1.7924113264046717 3.939e-09 1.8665320462941835 3.94e-09 1.8718439827266666 3.9409999999999995e-09 1.81300684695517 3.942e-09 1.7818338327492744 3.943e-09 1.8098552500900413 3.944e-09 1.826017253941129 3.945e-09 1.8063981099654456 3.946e-09 1.7957706186056563 3.947e-09 1.8981171602534048 3.948e-09 1.808597997232972 3.949e-09 1.8212003730338502 3.95e-09 1.7945530638223275 3.951e-09 1.8014044335853086 3.952e-09 1.741370418243568 3.953e-09 1.8417398843775443 3.954e-09 1.804772378124726 3.955e-09 1.8299007476042581 3.956e-09 1.835434973690841 3.957e-09 1.8540308709792797 3.958e-09 1.7705311261491652 3.959e-09 1.7661491560697857 3.9599999999999996e-09 1.834479270507401 3.961e-09 1.8606142678109043 3.962e-09 1.7718186600071484 3.963e-09 1.7846693802681506 3.964e-09 1.8477623597805115 3.965e-09 1.8895803124957475 3.966e-09 1.7834194656088673 3.967e-09 1.7690634193111727 3.9679999999999995e-09 1.831879941303993 3.969e-09 1.72807206337957 3.97e-09 1.7857111896628421 3.971e-09 1.74725497935257 3.972e-09 1.792961535746662 3.973e-09 1.8505215349149826 3.974e-09 1.8245094633750831 3.975e-09 1.7766478550272273 3.976e-09 1.8223774532118497 3.977e-09 1.7341906914521947 3.978e-09 1.7059503799684277 3.979e-09 1.7475478422101502 3.98e-09 1.836428907783954 3.981e-09 1.8317411941683264 3.982e-09 1.8177231282657749 3.983e-09 1.8273734660279795 3.984e-09 1.8040971917820612 3.985e-09 1.8357441960627867 3.986e-09 1.826067171999365 3.9869999999999996e-09 1.7960729285669776 3.988e-09 1.7825652539248718 3.989e-09 1.7749203265895288 3.99e-09 1.7923845274540346 3.991e-09 1.8189301024600821 3.992e-09 1.8319214415814344 3.993e-09 1.8495099185339663 3.994e-09 1.8286723298793013 3.9949999999999995e-09 1.8799341092940114 3.996e-09 1.7231932947175712 3.997e-09 1.786594408965189 3.998e-09 1.8425007601626409 3.999e-09 1.758615616611066 4e-09 1.7867026803964632 4.001e-09 1.8207448537156905 4.002e-09 1.8188815959002196 4.0029999999999995e-09 1.8580179585184484 4.004e-09 1.8062897869587096 4.005e-09 1.762122824607041 4.006e-09 1.7570005382838716 4.007e-09 1.8204810837350651 4.008e-09 1.7410360335289767 4.009e-09 1.8287881127676602 4.01e-09 1.841351930613003 4.011e-09 1.805934931299287 4.012e-09 1.8316215991175384 4.013e-09 1.8064973764130863 4.0139999999999996e-09 1.7345171587925987 4.015e-09 1.7860375594034554 4.016e-09 1.7729025722601137 4.017e-09 1.7530156220640287 4.018e-09 1.7320025082157309 4.019e-09 1.7740811021911296 4.02e-09 1.8064716704578356 4.021e-09 1.7929552807743097 4.0219999999999996e-09 1.7600441303213612 4.023e-09 1.7966563231858959 4.024e-09 1.7856995434771061 4.025e-09 1.783550291638169 4.026e-09 1.82248256091233 4.027e-09 1.8655041290450545 4.028e-09 1.775612254213613 4.029e-09 1.7877979257087036 4.0299999999999995e-09 1.8094035543402587 4.031e-09 1.7653999751552163 4.032e-09 1.7449071477812303 4.033e-09 1.7353845944631492 4.034e-09 1.7904128065749079 4.035e-09 1.831842708790152 4.036e-09 1.7783678982201554 4.037e-09 1.7319606119913624 4.038e-09 1.7905049159942348 4.039e-09 1.7241253520171922 4.04e-09 1.8720199212759545 4.041e-09 1.7995238248860772 4.042e-09 1.7910720871977004 4.043e-09 1.8164955699327 4.044e-09 1.8232824633473912 4.045e-09 1.7703385760599042 4.046e-09 1.6948479490269717 4.047e-09 1.8234699839728998 4.048e-09 1.8497271208518558 4.0489999999999996e-09 1.7781693007884234 4.05e-09 1.8669487410334844 4.051e-09 1.815659685489198 4.052e-09 1.81894442920656 4.053e-09 1.9400630764343885 4.054e-09 1.824963922131973 4.055e-09 1.8906813340615962 4.056e-09 1.81266164367322 4.0569999999999995e-09 1.849108999327484 4.058e-09 1.856763746964268 4.059e-09 1.8344696449845197 4.06e-09 1.7221496293816667 4.061e-09 1.8254200345205334 4.062e-09 1.8296082289821591 4.063e-09 1.929044320567583 4.064e-09 1.7554242022232371 4.0649999999999995e-09 1.8752132571935203 4.066e-09 1.7966707096959105 4.067e-09 1.685233675389946 4.068e-09 1.7765304153523964 4.069e-09 1.8165267073273608 4.07e-09 1.8326024496996638 4.071e-09 1.783174550396772 4.072e-09 1.7899934960304345 4.073e-09 1.885549230619548 4.074e-09 1.8274775258439448 4.075e-09 1.812618280651234 4.0759999999999996e-09 1.7798114073116849 4.077e-09 1.793512045118782 4.078e-09 1.787534006434439 4.079e-09 1.762456822181754 4.08e-09 1.737184005015169 4.081e-09 1.8084421573806984 4.082e-09 1.858495601789877 4.083e-09 1.801843159018142 4.0839999999999995e-09 1.8008306612203702 4.085e-09 1.7869546424742853 4.086e-09 1.8040644376944224 4.087e-09 1.8041424796583627 4.088e-09 1.7540850200236702 4.089e-09 1.7831650926490406 4.09e-09 1.8420585754241312 4.091e-09 1.8372232844583651 4.0919999999999995e-09 1.7703310693823595 4.093e-09 1.8516198035359812 4.094e-09 1.814170189907066 4.095e-09 1.74286964034255 4.096e-09 1.7311509151178868 4.097e-09 1.745973757171273 4.098e-09 1.9326648115973768 4.099e-09 1.8102969401223485 4.1e-09 1.8425078237636536 4.101e-09 1.7695314924992334 4.102e-09 1.788714872501946 4.1029999999999996e-09 1.75682377553084 4.104e-09 1.8450774230570393 4.105e-09 1.7362709910543808 4.106e-09 1.8772336334103399 4.107e-09 1.7827430158884023 4.108e-09 1.8167571302470724 4.109e-09 1.691583265114207 4.11e-09 1.7867805033389634 4.1109999999999996e-09 1.7265206531552273 4.112e-09 1.8391817573695866 4.113e-09 1.8292927695529284 4.114e-09 1.8024929130122829 4.115e-09 1.7315431423465282 4.116e-09 1.8432521291573072 4.117e-09 1.8597038577718652 4.118e-09 1.754212940814042 4.1189999999999995e-09 1.8336248871081795 4.12e-09 1.8209113877137444 4.121e-09 1.846668460451014 4.122e-09 1.7340347597046255 4.123e-09 1.865432592174745 4.124e-09 1.7847310419344526 4.125e-09 1.7981883081281365 4.126e-09 1.8760812592942322 4.127e-09 1.7592520653502755 4.128e-09 1.8669657690002837 4.129e-09 1.7163836173807523 4.13e-09 1.709450293752784 4.131e-09 1.7931703612883687 4.132e-09 1.7589967983255408 4.133e-09 1.7710810695841994 4.134e-09 1.7344053071453929 4.135e-09 1.7668123636877333 4.136e-09 1.796944862325345 4.137e-09 1.7444927348096118 4.1379999999999996e-09 1.7714869194606941 4.139e-09 1.7891806023007242 4.14e-09 1.8229631515909677 4.141e-09 1.7484632774932731 4.142e-09 1.8855218036933605 4.143e-09 1.8529283359489814 4.144e-09 1.7483941891603867 4.145e-09 1.8008463249092441 4.1459999999999995e-09 1.7495057912437761 4.147e-09 1.801589647473325 4.148e-09 1.809867143418938 4.149e-09 1.7733326203652446 4.15e-09 1.7975454413130278 4.151e-09 1.8075543862021077 4.152e-09 1.7632868654845526 4.153e-09 1.8454389119305612 4.1539999999999995e-09 1.7845520566038284 4.155e-09 1.7704080040526298 4.156e-09 1.7888126776797515 4.157e-09 1.8263996613158509 4.158e-09 1.8488800304889879 4.159e-09 1.7815248662515881 4.16e-09 1.8342665798869648 4.161e-09 1.8788024765651068 4.162e-09 1.7791133765315774 4.163e-09 1.8326371458954376 4.164e-09 1.783758761618367 4.1649999999999996e-09 1.7163023809589832 4.166e-09 1.8161222490501578 4.167e-09 1.8510408751072438 4.168e-09 1.7247088223825826 4.169e-09 1.805967110437358 4.17e-09 1.8770177033552375 4.171e-09 1.7561351869051953 4.172e-09 1.7862750426249399 4.1729999999999995e-09 1.812058427319155 4.174e-09 1.7979502929436517 4.175e-09 1.8524524434233185 4.176e-09 1.818356789690822 4.177e-09 1.8684319745445124 4.178e-09 1.747090452764852 4.179e-09 1.9578269385021325 4.18e-09 1.8635909006226945 4.1809999999999995e-09 1.8079704859788102 4.182e-09 1.8509493501058056 4.183e-09 1.7595311916331804 4.184e-09 1.826267918509757 4.185e-09 1.8199007765563757 4.186e-09 1.8040337981698984 4.187e-09 1.8474784280400203 4.188e-09 1.7336013932547731 4.189e-09 1.8372143995694048 4.19e-09 1.754619657698579 4.191e-09 1.7862177157394636 4.1919999999999996e-09 1.8210203557705884 4.193e-09 1.7816994995686326 4.194e-09 1.7236565716894088 4.195e-09 1.8463395824893516 4.196e-09 1.7379604746243853 4.197e-09 1.798232817168173 4.198e-09 1.7399941856508718 4.199e-09 1.793893931640932 4.1999999999999996e-09 1.9187244972489874 4.201e-09 1.7973934020060527 4.202e-09 1.8219138180648207 4.203e-09 1.762619592973922 4.204e-09 1.8046146891240658 4.205e-09 1.836305058800699 4.206e-09 1.8578358934939236 4.207e-09 1.7565673279284195 4.2079999999999995e-09 1.7749732869972341 4.209e-09 1.775370431441236 4.21e-09 1.9643249415770072 4.211e-09 1.9153207328041058 4.212e-09 1.835275717541051 4.213e-09 1.8784387669118627 4.214e-09 1.8078787804810201 4.215e-09 1.76759675451762 4.2159999999999995e-09 1.848000037920973 4.217e-09 1.7735556961471808 4.218e-09 1.745107396240987 4.219e-09 1.869622337327942 4.22e-09 1.7496436876329096 4.221e-09 1.820116317023686 4.222e-09 1.8057332060451465 4.223e-09 1.7029540634232119 4.224e-09 1.853194212739642 4.225e-09 1.8416750309882834 4.226e-09 1.7391656066176882 4.2269999999999996e-09 1.8707049560860967 4.228e-09 1.854446484355639 4.229e-09 1.8140539331552508 4.23e-09 1.7801124411817968 4.231e-09 1.7977261630491086 4.232e-09 1.8555448676116115 4.233e-09 1.767785635029425 4.234e-09 1.8200896643411504 4.2349999999999995e-09 1.7697293700395522 4.236e-09 1.8832119322570278 4.237e-09 1.8080788111847996 4.238e-09 1.7753059612036517 4.239e-09 1.775200845548516 4.24e-09 1.7879338436952998 4.241e-09 1.8213813764194793 4.242e-09 1.794585944887738 4.2429999999999995e-09 1.7671904041993698 4.244e-09 1.7975867638229974 4.245e-09 1.8433638729339448 4.246e-09 1.7933615601573953 4.247e-09 1.796501555194579 4.248e-09 1.7313008194018267 4.249e-09 1.8237491185078947 4.25e-09 1.7384623899309621 4.251e-09 1.8010018136415356 4.252e-09 1.7853025405730083 4.253e-09 1.742688694238176 4.2539999999999996e-09 1.7909903500906739 4.255e-09 1.7681601724934852 4.256e-09 1.715420968386165 4.257e-09 1.901673254371432 4.258e-09 1.7597872446692349 4.259e-09 1.7082834597662795 4.26e-09 1.8774177783537072 4.261e-09 1.7867315483790522 4.2619999999999996e-09 1.8322112072021666 4.263e-09 1.8236292935527103 4.264e-09 1.8232973832526989 4.265e-09 1.900763538933874 4.266e-09 1.7838109327128364 4.267e-09 1.8133879762865914 4.268e-09 1.7214884166820614 4.269e-09 1.7277895695205618 4.2699999999999995e-09 1.7217510060500776 4.271e-09 1.819435907701584 4.272e-09 1.7667013701609962 4.273e-09 1.7463272036861952 4.274e-09 1.8005500638294187 4.275e-09 1.721482657121868 4.276e-09 1.7797755023146278 4.277e-09 1.787407873979768 4.278e-09 1.776638146805512 4.279e-09 1.9147675593588056 4.28e-09 1.740090769015028 4.281e-09 1.766099256765258 4.282e-09 1.8143243789743153 4.283e-09 1.7985620504668975 4.284e-09 1.7122935306096563 4.285e-09 1.8378008302903621 4.286e-09 1.7630243633789628 4.287e-09 1.799608517928063 4.288e-09 1.7838143544075646 4.2889999999999996e-09 1.7474297777073788 4.29e-09 1.8380161045208603 4.291e-09 1.7899696915832959 4.292e-09 1.863833406378181 4.293e-09 1.7387868997077576 4.294e-09 1.7661654665196056 4.295e-09 1.7849432001175067 4.296e-09 1.8611318805313102 4.2969999999999995e-09 1.7638205239878328 4.298e-09 1.8245578634500113 4.299e-09 1.8524436909628736 4.3e-09 1.7708196440927346 4.301e-09 1.6340987085993361 4.302e-09 1.7591939310010771 4.303e-09 1.7871235668312764 4.304e-09 1.816008887787486 4.3049999999999995e-09 1.9000568923131098 4.306e-09 1.7956263341704561 4.307e-09 1.7991445904052905 4.308e-09 1.782689365867961 4.309e-09 1.8117760719768812 4.31e-09 1.6858414442636775 4.311e-09 1.8482478357681709 4.312e-09 1.815794439692008 4.313e-09 1.793242977553835 4.314e-09 1.7855442085463973 4.315e-09 1.7512272756221536 4.3159999999999996e-09 1.7477898549887283 4.317e-09 1.7503558755078688 4.318e-09 1.819214149012609 4.319e-09 1.8178065963612429 4.32e-09 1.7194936009597623 4.321e-09 1.8535569143569794 4.322e-09 1.779261553041018 4.323e-09 1.825820508486345 4.3239999999999995e-09 1.8103003357405416 4.325e-09 1.7949958572262803 4.326e-09 1.7960200338018388 4.327e-09 1.799282406914187 4.328e-09 1.836421764585402 4.329e-09 1.8383618836839821 4.33e-09 1.8341086904522383 4.331e-09 1.837128110226328 4.3319999999999995e-09 1.79957859495394 4.333e-09 1.7574685739858638 4.334e-09 1.844621827822053 4.335e-09 1.6939695684288165 4.336e-09 1.7792045718790515 4.337e-09 1.7349765575845146 4.338e-09 1.8021414314559168 4.339e-09 1.795465934456453 4.34e-09 1.734892067961914 4.341e-09 1.7325305243314464 4.342e-09 1.7921700235225497 4.3429999999999996e-09 1.779591821156911 4.344e-09 1.7446293035398135 4.345e-09 1.7835918313915873 4.346e-09 1.8687022739345567 4.347e-09 1.7622439112954398 4.348e-09 1.822322452301093 4.349e-09 1.815974246417369 4.35e-09 1.7958314715515378 4.3509999999999996e-09 1.7735925108853914 4.352e-09 1.7769968126821178 4.353e-09 1.7646185858486816 4.354e-09 1.7825788079340665 4.355e-09 1.8263745433905698 4.356e-09 1.7415098633025479 4.357e-09 1.76304694706609 4.358e-09 1.8293710905026257 4.3589999999999995e-09 1.8216271967455506 4.36e-09 1.816898939094882 4.361e-09 1.811911048807893 4.362e-09 1.7384793876199107 4.363e-09 1.738571784400444 4.364e-09 1.8733187081610574 4.365e-09 1.7917496995629827 4.366e-09 1.852306280135698 4.3669999999999995e-09 1.8092044539516274 4.368e-09 1.7909994597903656 4.369e-09 1.7609061950861473 4.37e-09 1.7514858043769967 4.371e-09 1.7951923138694974 4.372e-09 1.8351813952308227 4.373e-09 1.7800372294085594 4.374e-09 1.7057586079748708 4.375e-09 1.8291926389257105 4.376e-09 1.7769905176588379 4.377e-09 1.8213916308732068 4.3779999999999996e-09 1.8100880368409198 4.379e-09 1.7143085999666976 4.38e-09 1.7226911316045783 4.381e-09 1.8278790379708136 4.382e-09 1.8762951158264891 4.383e-09 1.8832298153737175 4.384e-09 1.7675531259182904 4.385e-09 1.783743732764864 4.3859999999999995e-09 1.7848731966550144 4.387e-09 1.7966571342341968 4.388e-09 1.6666560273731892 4.389e-09 1.8235680828134357 4.39e-09 1.7292062003841997 4.391e-09 1.7238111992820493 4.392e-09 1.7555610064555343 4.393e-09 1.7927507070530757 4.3939999999999995e-09 1.7310670266101063 4.395e-09 1.7721788204867968 4.396e-09 1.896883783742216 4.397e-09 1.8601840148429827 4.398e-09 1.8179492025309876 4.399e-09 1.804931368546835 4.4e-09 1.796426946157079 4.401e-09 1.828516352581993 4.402e-09 1.7155595315699392 4.403e-09 1.7897700505265428 4.404e-09 1.8466461844315225 4.4049999999999996e-09 1.7805134488021879 4.406e-09 1.7859253901101 4.407e-09 1.7717125887125655 4.408e-09 1.87376914619857 4.409e-09 1.8100064224729309 4.41e-09 1.772270106898788 4.411e-09 1.8537048097624556 4.412e-09 1.7851002727790515 4.4129999999999995e-09 1.7365438696417164 4.414e-09 1.752513939850097 4.415e-09 1.8218846336417467 4.416e-09 1.844246208252535 4.417e-09 1.7701563339544764 4.418e-09 1.7831634428812517 4.419e-09 1.78821866458754 4.42e-09 1.835820945469855 4.4209999999999995e-09 1.8301960921470242 4.422e-09 1.8494493373742955 4.423e-09 1.7722656326236035 4.424e-09 1.7433703994687242 4.425e-09 1.7601200827926256 4.426e-09 1.8119060027400542 4.427e-09 1.8046416496766506 4.428e-09 1.70397947837902 4.429e-09 1.83787398383966 4.43e-09 1.7126093879758677 4.431e-09 1.8931883019416882 4.4319999999999996e-09 1.7674807973896103 4.433e-09 1.8663590779115733 4.434e-09 1.754470668567566 4.435e-09 1.730364506167612 4.436e-09 1.7479012715256834 4.437e-09 1.78423633792037 4.438e-09 1.7492651117794982 4.439e-09 1.8379917792714302 4.4399999999999996e-09 1.7751290235980426 4.441e-09 1.7833838209332336 4.442e-09 1.7879232418171496 4.443e-09 1.7980577809446794 4.444e-09 1.7553298900714571 4.445e-09 1.8109622136559864 4.446e-09 1.8254372397446539 4.447e-09 1.7208426991284127 4.4479999999999995e-09 1.7973732187255067 4.449e-09 1.783690576339366 4.45e-09 1.8257225546335338 4.451e-09 1.7438199681606665 4.452e-09 1.7709139620768466 4.453e-09 1.794560161957345 4.454e-09 1.7667197044910543 4.455e-09 1.780310254770077 4.4559999999999995e-09 1.7868374577028305 4.457e-09 1.8119328108184787 4.458e-09 1.8351673931383006 4.459e-09 1.778851904971721 4.46e-09 1.8093082551856607 4.461e-09 1.7491331085679205 4.462e-09 1.863516449231385 4.463e-09 1.8112186009196796 4.464e-09 1.84851688901149 4.465e-09 1.734943530826389 4.466e-09 1.787447479770971 4.4669999999999996e-09 1.808716042393092 4.468e-09 1.7749122575648717 4.469e-09 1.7347420340896706 4.47e-09 1.788342425108674 4.471e-09 1.7778266755671466 4.472e-09 1.7730226528389685 4.473e-09 1.7846664418598719 4.474e-09 1.7804704930862456 4.4749999999999995e-09 1.7452314208087172 4.476e-09 1.8327900186001724 4.477e-09 1.8471433065672158 4.478e-09 1.84047150210862 4.479e-09 1.9521010246476913 4.48e-09 1.7538790548557632 4.481e-09 1.7604665995256499 4.482e-09 1.8313487558330843 4.4829999999999995e-09 1.801573404476279 4.484e-09 1.773507930318884 4.485e-09 1.7849833893684923 4.486e-09 1.8217388384839583 4.487e-09 1.8692471456956792 4.488e-09 1.8310941653763084 4.489e-09 1.8053467458161112 4.49e-09 1.7959450136440906 4.491e-09 1.759549327827365 4.492e-09 1.6512103540480392 4.493e-09 1.8324998686621168 4.4939999999999996e-09 1.7789857164536442 4.495e-09 1.8093477460299707 4.496e-09 1.8024047112891715 4.497e-09 1.835687208237054 4.498e-09 1.7832393227594634 4.499e-09 1.850426413072855 4.5e-09 1.8122811475019582 4.501e-09 1.775981158472461 4.5019999999999995e-09 1.8172954724016974 4.503e-09 1.8989416184984291 4.504e-09 1.8110181720777738 4.505e-09 1.784916205309292 4.506e-09 1.824516453357862 4.507e-09 1.7969546109826087 4.508e-09 1.7733525599975948 4.509e-09 1.7731401798193658 4.5099999999999995e-09 1.8140846956435956 4.511e-09 1.868721314762469 4.512e-09 1.8009898538773499 4.513e-09 1.8421124492454908 4.514e-09 1.8522062034458968 4.515e-09 1.8184975220835866 4.516e-09 1.6397170738715183 4.517e-09 1.7632910627287999 4.518e-09 1.814756569895544 4.519e-09 1.8513788085487666 4.52e-09 1.7131715778373955 4.521e-09 1.7456660768043462 4.522e-09 1.7134737872762515 4.523e-09 1.86152734268761 4.524e-09 1.681540881772873 4.525e-09 1.7503499757237415 4.526e-09 1.8332824011092193 4.527e-09 1.7564903653493058 4.528e-09 1.7859278668596554 4.5289999999999996e-09 1.7653495897670892 4.53e-09 1.8251789801225682 4.531e-09 1.7160932492011562 4.532e-09 1.787027772059142 4.533e-09 1.749442036733137 4.534e-09 1.8374605330089762 4.535e-09 1.7326710177873406 4.536e-09 1.813191305223897 4.5369999999999995e-09 1.7335746672718626 4.538e-09 1.8803871921924373 4.539e-09 1.8023325751313062 4.54e-09 1.8624355637976648 4.541e-09 1.8355011998471404 4.542e-09 1.8139020616360253 4.543e-09 1.8441270902829865 4.544e-09 1.8058927561134726 4.5449999999999995e-09 1.8024627027200244 4.546e-09 1.841540283721111 4.547e-09 1.8623968136843931 4.548e-09 1.8465617460701904 4.549e-09 1.8215776809746882 4.55e-09 1.8327829452671405 4.551e-09 1.8240806648244625 4.552e-09 1.7662756459280924 4.553e-09 1.7945311853500332 4.554e-09 1.8812262248171554 4.555e-09 1.7675847922366954 4.5559999999999996e-09 1.744851754324019 4.557e-09 1.8348656125120024 4.558e-09 1.7814491829800978 4.559e-09 1.7970768833835902 4.56e-09 1.7582710519091356 4.561e-09 1.853024719074163 4.562e-09 1.7550621838915437 4.563e-09 1.8436935559850627 4.5639999999999995e-09 1.8580488152247572 4.565e-09 1.7428501219651793 4.566e-09 1.7573259044848901 4.567e-09 1.7749440853581198 4.568e-09 1.8526608186409967 4.569e-09 1.770062566928969 4.57e-09 1.7908300734152716 4.571e-09 1.7791064377808838 4.5719999999999995e-09 1.7459418619919185 4.573e-09 1.8341653900474955 4.574e-09 1.791081993058946 4.575e-09 1.8531604459488584 4.576e-09 1.731176423002348 4.577e-09 1.742321814985959 4.578e-09 1.7954952606438177 4.579e-09 1.7961194749126326 4.58e-09 1.7486232252451002 4.581e-09 1.7594039528617804 4.582e-09 1.7848836206187104 4.5829999999999996e-09 1.8590048464619275 4.584e-09 1.7987888113162196 4.585e-09 1.794237163705465 4.586e-09 1.7719964448710321 4.587e-09 1.8288075796717191 4.588e-09 1.8124072346749294 4.589e-09 1.8036964296085973 4.59e-09 1.7862780850478268 4.5909999999999996e-09 1.8307713451106689 4.592e-09 1.83977098413826 4.593e-09 1.8724395026046499 4.594e-09 1.860339670021363 4.595e-09 1.8365549541191433 4.596e-09 1.7639740908816974 4.597e-09 1.844339269126893 4.598e-09 1.7557663650283188 4.5989999999999995e-09 1.8167854525550178 4.6e-09 1.8472048904070444 4.601e-09 1.8140650085059826 4.602e-09 1.8078623502485944 4.603e-09 1.917596680353839 4.604e-09 1.8261046693456113 4.605e-09 1.7917138303867637 4.606e-09 1.8231178922006774 4.6069999999999995e-09 1.813863966289514 4.608e-09 1.8841963323619935 4.609e-09 1.8046428543085415 4.61e-09 1.7908120078785166 4.611e-09 1.774851645157821 4.612e-09 1.7530082756280079 4.613e-09 1.71968386063504 4.614e-09 1.8270349463851003 4.615e-09 1.8186691347602884 4.616e-09 1.8250817798771712 4.617e-09 1.8772799711335297 4.6179999999999996e-09 1.79827720201357 4.619e-09 1.832172755520971 4.62e-09 1.8731982926738955 4.621e-09 1.798439036151863 4.622e-09 1.8272618349367948 4.623e-09 1.7998784465081166 4.624e-09 1.8507955723565794 4.625e-09 1.8132106488270447 4.6259999999999995e-09 1.7997068179144662 4.627e-09 1.8544055447788872 4.628e-09 1.7827347602008607 4.629e-09 1.7569350062609543 4.63e-09 1.7765255967737064 4.631e-09 1.9282201230082274 4.632e-09 1.763392533622862 4.633e-09 1.7628288052602303 4.6339999999999995e-09 1.7931189691851852 4.635e-09 1.9213354749125848 4.636e-09 1.7446476039552692 4.637e-09 1.7433941827160035 4.638e-09 1.7743039965185856 4.639e-09 1.787967817998626 4.64e-09 1.8404733754194773 4.641e-09 1.7759270608229472 4.642e-09 1.8435233510004294 4.643e-09 1.7973140033336341 4.644e-09 1.760482913382882 4.6449999999999996e-09 1.76921572475008 4.646e-09 1.8039532732747818 4.647e-09 1.7250832271858563 4.648e-09 1.7600013000945371 4.649e-09 1.828642504202374 4.65e-09 1.752444932601016 4.651e-09 1.6306754459040769 4.652e-09 1.8216509549434141 4.6529999999999995e-09 1.7535071666442577 4.654e-09 1.802507170897513 4.655e-09 1.8081353962407778 4.656e-09 1.8011327224888671 4.657e-09 1.8271942779921806 4.658e-09 1.8762208356452394 4.659e-09 1.8286992625019067 4.66e-09 1.8632164975883878 4.6609999999999995e-09 1.828235342636673 4.662e-09 1.8539581640026348 4.663e-09 1.7257664892022426 4.664e-09 1.8257773654280627 4.665e-09 1.8092392307725824 4.666e-09 1.7168550549094732 4.667e-09 1.799430286118944 4.668e-09 1.7838752083752756 4.669e-09 1.8284673327237397 4.67e-09 1.8780001630290546 4.671e-09 1.8259751724372728 4.6719999999999996e-09 1.7660246888825648 4.673e-09 1.8055439294636413 4.674e-09 1.8138953151564157 4.675e-09 1.8025580633914966 4.676e-09 1.8286961998980313 4.677e-09 1.85280221906228 4.678e-09 1.7604672599731757 4.679e-09 1.7956822469046227 4.6799999999999996e-09 1.7999292806300613 4.681e-09 1.800465653022716 4.682e-09 1.8009963164410705 4.683e-09 1.8245285767541086 4.684e-09 1.872259430609179 4.685e-09 1.8405021309791179 4.686e-09 1.7232098471147732 4.687e-09 1.7754811353142552 4.6879999999999995e-09 1.8456929419967039 4.689e-09 1.7607535693866492 4.69e-09 1.7651029893880839 4.691e-09 1.8367838568488577 4.692e-09 1.824301285785193 4.693e-09 1.772910742713373 4.694e-09 1.8175989919788185 4.695e-09 1.710907119572098 4.6959999999999995e-09 1.8258028991979978 4.697e-09 1.8036675416634889 4.698e-09 1.8095544324446964 4.699e-09 1.8508629194295902 4.7e-09 1.8728623704953942 4.701e-09 1.8380941689215855 4.702e-09 1.7680666299987808 4.703e-09 1.830523650776481 4.704e-09 1.8314844501682381 4.705e-09 1.7569425424908944 4.706e-09 1.8121890458154408 4.7069999999999996e-09 1.8719726191515667 4.708e-09 1.7316344826315644 4.709e-09 1.8218741229503717 4.71e-09 1.7642305092708295 4.711e-09 1.8130559150380112 4.712e-09 1.8039541939280739 4.713e-09 1.7674908082417722 4.714e-09 1.8815889934808454 4.7149999999999995e-09 1.7708636062650014 4.716e-09 1.8558618388129653 4.717e-09 1.764129036080743 4.718e-09 1.8043154710295588 4.719e-09 1.801434695101074 4.72e-09 1.7417145744552707 4.721e-09 1.8239047153539456 4.722e-09 1.7274641064976985 4.7229999999999995e-09 1.682759974713432 4.724e-09 1.9028555866982184 4.725e-09 1.746241695259921 4.726e-09 1.7319626455159107 4.727e-09 1.7654057037130615 4.728e-09 1.7282253847891014 4.729e-09 1.8674124288629075 4.73e-09 1.7488179281338223 4.731e-09 1.887310918959741 4.732e-09 1.7692147698205833 4.733e-09 1.8201979160752608 4.7339999999999996e-09 1.8763213479997556 4.735e-09 1.8276695609902172 4.736e-09 1.8236355477226174 4.737e-09 1.827454869051527 4.738e-09 1.8665538541212674 4.739e-09 1.7651222753058184 4.74e-09 1.8032847946506312 4.741e-09 1.8502233709418894 4.7419999999999995e-09 1.7797363959350117 4.743e-09 1.7447826662580939 4.744e-09 1.8870994796029998 4.745e-09 1.8026263002354252 4.746e-09 1.7947572312272042 4.747e-09 1.8555822318660007 4.748e-09 1.8338956366885504 4.749e-09 1.7301910158881426 4.7499999999999995e-09 1.7130521484533912 4.751e-09 1.762585353254417 4.752e-09 1.7939223173473864 4.753e-09 1.842131677581162 4.754e-09 1.8221663076967027 4.755e-09 1.777398520081129 4.756e-09 1.8244765899608086 4.757e-09 1.7572254312783704 4.7579999999999995e-09 1.7258524813809017 4.759e-09 1.8016207789953755 4.76e-09 1.8189978952514838 4.7609999999999996e-09 1.8601479206265732 4.762e-09 1.801906725297832 4.763e-09 1.867851559893478 4.764e-09 1.7570656925346064 4.765e-09 1.8216540198736815 4.766e-09 1.7803364684598295 4.767e-09 1.7862405594965043 4.768e-09 1.836505738526418 4.7689999999999996e-09 1.8129481911237821 4.77e-09 1.8518747265484357 4.771e-09 1.7856480895565796 4.772e-09 1.8636790229885256 4.773e-09 1.8288663024903598 4.774e-09 1.7151537452862702 4.775e-09 1.7532460515949448 4.776e-09 1.8382829349989018 4.7769999999999995e-09 1.7747941431740455 4.778e-09 1.8441363847905405 4.779e-09 1.7910801146910071 4.78e-09 1.6873367650166227 4.781e-09 1.7700926249186917 4.782e-09 1.7241842573787542 4.783e-09 1.8743002087912093 4.784e-09 1.796957746515116 4.7849999999999995e-09 1.779666945177568 4.786e-09 1.8259740313380874 4.787e-09 1.8719553036194347 4.788e-09 1.760443362266521 4.789e-09 1.785258095108623 4.79e-09 1.8741254501869615 4.791e-09 1.8172728236832014 4.792e-09 1.8713463257948983 4.793e-09 1.7495639203170035 4.794e-09 1.7254814834637586 4.795e-09 1.705127497599709 4.7959999999999996e-09 1.7956574868272683 4.797e-09 1.7673875182863406 4.798e-09 1.7012030473203943 4.799e-09 1.8942501817353836 4.8e-09 1.7445364552655311 4.801e-09 1.7500853484984467 4.802e-09 1.74219783921639 4.803e-09 1.7788540436790863 4.8039999999999995e-09 1.8508936359863621 4.805e-09 1.7854116180577784 4.806e-09 1.7449941818501167 4.807e-09 1.8015247029063888 4.808e-09 1.8647973314551898 4.809e-09 1.781209293022014 4.81e-09 1.7764218493143156 4.811e-09 1.8481915764178152 4.8119999999999995e-09 1.8045702027396082 4.813e-09 1.8285374324190797 4.814e-09 1.811256725796657 4.815e-09 1.898994131176133 4.816e-09 1.7683497693405181 4.817e-09 1.7932536983579332 4.818e-09 1.7997585321137004 4.819e-09 1.8014589464653161 4.82e-09 1.865514052939183 4.821e-09 1.832040898678432 4.822e-09 1.8467980528232275 4.8229999999999996e-09 1.77413878560707 4.824e-09 1.7094590277932966 4.825e-09 1.8253311136320844 4.826e-09 1.8062836868783823 4.827e-09 1.8248594798654185 4.828e-09 1.837135283700965 4.829e-09 1.78178282892891 4.83e-09 1.7430085296887292 4.8309999999999996e-09 1.7295856980827127 4.832e-09 1.7625913582370898 4.833e-09 1.7507057238992312 4.834e-09 1.7893854088840975 4.835e-09 1.892345081679362 4.836e-09 1.7813022938600434 4.837e-09 1.773804774328816 4.838e-09 1.7838345198809296 4.8389999999999995e-09 1.8059878336685629 4.84e-09 1.8863851720999714 4.841e-09 1.8000224553755266 4.842e-09 1.7650419474245742 4.843e-09 1.878930035182073 4.844e-09 1.800856437563888 4.845e-09 1.7535940850812208 4.846e-09 1.8248202232812936 4.8469999999999995e-09 1.8080176272795505 4.848e-09 1.923111497343316 4.849e-09 1.8590300112748013 4.85e-09 1.723881812835053 4.851e-09 1.814422460781221 4.852e-09 1.7844040521581244 4.853e-09 1.7867015430992113 4.854e-09 1.8610023190328107 4.855e-09 1.7644563460092544 4.856e-09 1.8127975336613396 4.857e-09 1.8424649074904065 4.8579999999999996e-09 1.8053775206395632 4.859e-09 1.797773246581477 4.86e-09 1.8831762540564057 4.861e-09 1.8559229626331586 4.862e-09 1.8747842116035174 4.863e-09 1.745427887877299 4.864e-09 1.7309183084151358 4.865e-09 1.7725925516827084 4.8659999999999995e-09 1.7509570497632774 4.867e-09 1.8430606119956443 4.868e-09 1.7739697972209025 4.869e-09 1.8514488536389018 4.87e-09 1.7767438629492207 4.871e-09 1.9474334668810132 4.872e-09 1.836041655789102 4.873e-09 1.8189455937163697 4.8739999999999995e-09 1.7373546988614958 4.875e-09 1.8613385990105782 4.876e-09 1.7798118189071985 4.877e-09 1.8099325376539668 4.878e-09 1.8380942542072898 4.879e-09 1.777932644086802 4.88e-09 1.7198998256503946 4.881e-09 1.8344397497248013 4.882e-09 1.7815574865047388 4.883e-09 1.894939576188724 4.884e-09 1.7857383663828659 4.8849999999999996e-09 1.791088852061788 4.886e-09 1.7885577672889454 4.887e-09 1.7902764225410623 4.888e-09 1.7729820111079737 4.889e-09 1.7949660014394457 4.89e-09 1.828579469527729 4.891e-09 1.7659217073345768 4.892e-09 1.8448805732642268 4.8929999999999995e-09 1.8193223510918486 4.894e-09 1.8664345058988274 4.895e-09 1.7685936153135624 4.896e-09 1.7063081747829794 4.897e-09 1.8182131171555456 4.898e-09 1.7935508160807503 4.899e-09 1.7981428381574203 4.9e-09 1.7166600315505822 4.9009999999999995e-09 1.7182758792847932 4.902e-09 1.7461675225422362 4.903e-09 1.7624365181565187 4.904e-09 1.8347603791099358 4.905e-09 1.8926591078969681 4.906e-09 1.7136679042084129 4.907e-09 1.8169097637218068 4.908e-09 1.7974303030419199 4.9089999999999995e-09 1.8154085032560234 4.91e-09 1.8161278589364362 4.911e-09 1.7847088845650545 4.9119999999999996e-09 1.8791999959862267 4.913e-09 1.8057469600506606 4.914e-09 1.7267083565740193 4.915e-09 1.8848301608544378 4.916e-09 1.8206010266848176 4.917e-09 1.8133339536476087 4.918e-09 1.8220523191015148 4.919e-09 1.805315231066345 4.9199999999999996e-09 1.7558448828162823 4.921e-09 1.8314299636269664 4.922e-09 1.7195620074117612 4.923e-09 1.764611315914916 4.924e-09 1.8239925084422062 4.925e-09 1.8126177930333227 4.926e-09 1.805155180931018 4.927e-09 1.8143036744879086 4.9279999999999995e-09 1.7841963970256542 4.929e-09 1.8191232388247547 4.93e-09 1.7463798795662955 4.931e-09 1.946260585513055 4.932e-09 1.7584049685764882 4.933e-09 1.7439977212409254 4.934e-09 1.8265115047140759 4.935e-09 1.7912360845514061 4.9359999999999995e-09 1.724333238806797 4.937e-09 1.8090963677310534 4.938e-09 1.8411963961494608 4.939e-09 1.8873074614822236 4.94e-09 1.7470534141462126 4.941e-09 1.8015999108807155 4.942e-09 1.7439294747486596 4.943e-09 1.800350057791276 4.944e-09 1.7337063583275576 4.945e-09 1.801612699182223 4.946e-09 1.7234671017303436 4.9469999999999996e-09 1.6647890071341662 4.948e-09 1.8707963655258255 4.949e-09 1.850804779393036 4.95e-09 1.820778302832217 4.951e-09 1.8211701690401814 4.952e-09 1.7757951249906965 4.953e-09 1.78983407339323 4.954e-09 1.7496498263509859 4.9549999999999995e-09 1.7663985005690857 4.956e-09 1.774657012059998 4.957e-09 1.8441057518799504 4.958e-09 1.8514836034161866 4.959e-09 1.747631824073693 4.96e-09 1.9714579213135166 4.961e-09 1.7961334762244896 4.962e-09 1.8539463720893061 4.9629999999999995e-09 1.8666084836674546 4.964e-09 1.804725700382607 4.965e-09 1.7925054905614284 4.966e-09 1.8311335138117524 4.967e-09 1.8789512324726083 4.968e-09 1.8162627635639519 4.969e-09 1.9201109914919194 4.97e-09 1.822811138835936 4.971e-09 1.8513197515918591 4.972e-09 1.8010785573333594 4.973e-09 1.7821361711515853 4.9739999999999996e-09 1.8466907018356968 4.975e-09 1.8196064988649476 4.976e-09 1.794934559092169 4.977e-09 1.7247635098857372 4.978e-09 1.8449482172715739 4.979e-09 1.802807784850055 4.98e-09 1.6975163152129311 4.981e-09 1.9162688680384337 4.9819999999999995e-09 1.7190828154615714 4.983e-09 1.7492078975283383 4.984e-09 1.8594296748574473 4.985e-09 1.7831008994222763 4.986e-09 1.8132717882409546 4.987e-09 1.7429795942565738 4.988e-09 1.8850182642969415 4.989e-09 1.8779342847457707 4.9899999999999995e-09 1.7461395653607505 4.991e-09 1.8857754295583329 4.992e-09 1.748540623082337 4.993e-09 1.8024428079095174 4.994e-09 1.7998508603321084 4.995e-09 1.808853374628129 4.996e-09 1.864323760724961 4.997e-09 1.8313132401273626 4.9979999999999995e-09 1.7423663174366704 4.999e-09 1.7901767195202436 5e-09 1.859036184920056 5.0009999999999996e-09 1.7972301500821757 5.002e-09 1.7940931503135815 5.003e-09 1.7549214978959873 5.004e-09 1.787344440305178 5.005e-09 1.7787038242595052 5.006e-09 1.812575159679586 5.007e-09 1.8666005353937165 5.008e-09 1.7613276357613157 5.0089999999999996e-09 1.9243685297602242 5.01e-09 1.788417802384982 5.011e-09 1.829012956591981 5.012e-09 1.6886979984083113 5.013e-09 1.8052127536970637 5.014e-09 1.751984294283188 5.015e-09 1.8342437162254293 5.016e-09 1.702528677123809 5.0169999999999995e-09 1.8323424472939691 5.018e-09 1.8302425360489247 5.019e-09 1.7605438597467575 5.02e-09 1.9513733756278877 5.021e-09 1.8466978958041964 5.022e-09 1.838226563315847 5.023e-09 1.7864853488012749 5.024e-09 1.8135285134993187 5.0249999999999995e-09 1.7477357722252091 5.026e-09 1.766297289272508 5.027e-09 1.8068726494919727 5.028e-09 1.8294931813976147 5.029e-09 1.7796246879473876 5.03e-09 1.7617979617908963 5.031e-09 1.8528348015518235 5.032e-09 1.7896015426047112 5.033e-09 1.7433925029832407 5.034e-09 1.7529321692212292 5.035e-09 1.8322176548084808 5.0359999999999996e-09 1.815674901621624 5.037e-09 1.8091189814817001 5.038e-09 1.8987343858361732 5.039e-09 1.9104441067875308 5.04e-09 1.8197817494722994 5.041e-09 1.8383099837142445 5.042e-09 1.8562117421638944 5.043e-09 1.8719776435051463 5.0439999999999995e-09 1.8088026711072804 5.045e-09 1.8234466106093206 5.046e-09 1.780020009138736 5.047e-09 1.8131480278423877 5.048e-09 1.8228535396215706 5.049e-09 1.8555307956504543 5.05e-09 1.859945172597121 5.051e-09 1.8207742945097678 5.0519999999999995e-09 1.8689634027093411 5.053e-09 1.7917258396228442 5.054e-09 1.8290279921405543 5.055e-09 1.8545992064571335 5.056e-09 1.8864676038525834 5.057e-09 1.8426103830287772 5.058e-09 1.834909336359007 5.059e-09 1.712557191740639 5.06e-09 1.8243141068219757 5.061e-09 1.8612436112456683 5.062e-09 1.8092383399088994 5.0629999999999996e-09 1.72695434664864 5.064e-09 1.8250263282786319 5.065e-09 1.7421410255568455 5.066e-09 1.9096837359735097 5.067e-09 1.8086025440866116 5.068e-09 1.7640394102267807 5.069e-09 1.7987398832706454 5.07e-09 1.7335708435310757 5.0709999999999995e-09 1.8631448733558753 5.072e-09 1.7645144214238373 5.073e-09 1.7586960006063965 5.074e-09 1.8194079318499061 5.075e-09 1.82873053458324 5.076e-09 1.8130784203000432 5.077e-09 1.7539068016625325 5.078e-09 1.8422042916408976 5.0789999999999995e-09 1.851262480210894 5.08e-09 1.7765520214175856 5.081e-09 1.6972894346155276 5.082e-09 1.6691584333788534 5.083e-09 1.79070044885932 5.084e-09 1.800483378967493 5.085e-09 1.790454118452659 5.086e-09 1.8929081167958253 5.0869999999999995e-09 1.7917376383180728 5.088e-09 1.7994564505904365 5.089e-09 1.8621243512380576 5.09e-09 1.797515066115408 5.091e-09 1.7811875807945348 5.092e-09 1.8801473669505364 5.093e-09 1.8252266443746217 5.094e-09 1.822920867923984 5.095e-09 1.8890564881520402 5.096e-09 1.7920453847725846 5.097e-09 1.8057654050321448 5.0979999999999996e-09 1.6975360891274305 5.099e-09 1.852060645420377 5.1e-09 1.827002298794332 5.101e-09 1.7747779541205975 5.102e-09 1.7945504451177658 5.103e-09 1.7684258403430115 5.104e-09 1.787011200387376 5.105e-09 1.7681807880167777 5.1059999999999995e-09 1.8155657857878886 5.107e-09 1.7923778480295156 5.108e-09 1.7353655615892372 5.109e-09 1.8676150946914591 5.11e-09 1.9038936772403194 5.111e-09 1.7116100494492728 5.112e-09 1.860501172188971 5.113e-09 1.7479546268091162 5.1139999999999995e-09 1.7689484192776932 5.115e-09 1.8595200584433902 5.116e-09 1.7253641589815376 5.117e-09 1.8251397124180517 5.118e-09 1.7746695478567327 5.119e-09 1.8245242227854126 5.12e-09 1.7773200637009863 5.121e-09 1.8189637307748165 5.122e-09 1.7060755269999615 5.123e-09 1.7892391357614583 5.124e-09 1.9262962545959916 5.1249999999999996e-09 1.8605265852493673 5.126e-09 1.8072580384182033 5.127e-09 1.8681054723507509 5.128e-09 1.7312025075555595 5.129e-09 1.8171697351661207 5.13e-09 1.7897385185992696 5.131e-09 1.8247494995835063 5.132e-09 1.809683137209803 5.1329999999999995e-09 1.8213922682864576 5.134e-09 1.8737440773344387 5.135e-09 1.7609167601043338 5.136e-09 1.7901333266459143 5.137e-09 1.6720974673090243 5.138e-09 1.745597356174432 5.139e-09 1.7526065775652695 5.14e-09 1.7822731460025167 5.1409999999999995e-09 1.761439632399462 5.142e-09 1.7966965759007971 5.143e-09 1.7887231593797146 5.144e-09 1.7855591552120424 5.145e-09 1.8495726777711194 5.146e-09 1.784486707483284 5.147e-09 1.7682644846601845 5.148e-09 1.7620904418968997 5.1489999999999995e-09 1.7518686974175235 5.15e-09 1.803133302060264 5.151e-09 1.794427023556683 5.1519999999999996e-09 1.8762278996690371 5.153e-09 1.7799000876429192 5.154e-09 1.806095639843807 5.155e-09 1.820550973988247 5.156e-09 1.7432396901190357 5.157e-09 1.8064059356541777 5.158e-09 1.7391832472210824 5.159e-09 1.7833611586857732 5.1599999999999996e-09 1.8295005537724711 5.161e-09 1.792797553666973 5.162e-09 1.8452730654437521 5.163e-09 1.8090347982597808 5.164e-09 1.8163529393632307 5.165e-09 1.7662262746870412 5.166e-09 1.7412729423740223 5.167e-09 1.8884486269157512 5.1679999999999995e-09 1.883700209057955 5.169e-09 1.8326003931629438 5.17e-09 1.79186501682012 5.171e-09 1.7041119351054783 5.172e-09 1.8084389706505377 5.173e-09 1.7534077882623578 5.174e-09 1.8064033645618114 5.175e-09 1.7613258140372405 5.1759999999999995e-09 1.8306595688472551 5.177e-09 1.8076782273876766 5.178e-09 1.8062055521812959 5.179e-09 1.7442056014433833 5.18e-09 1.8131225441224204 5.181e-09 1.803423908806955 5.182e-09 1.8641599267820197 5.183e-09 1.816307791764157 5.184e-09 1.8568647747689784 5.185e-09 1.7919442192869388 5.186e-09 1.844138140343641 5.1869999999999996e-09 1.8372572972389682 5.188e-09 1.7551022255549018 5.189e-09 1.8124416626928481 5.19e-09 1.8193198966720894 5.191e-09 1.7005922751297982 5.192e-09 1.7811550990144498 5.193e-09 1.7920323652703605 5.194e-09 1.7865277805461055 5.1949999999999995e-09 1.7335322093329941 5.196e-09 1.8529335912771774 5.197e-09 1.8582244137501147 5.198e-09 1.7386439796731141 5.199e-09 1.7948281132393638 5.2e-09 1.754645456124719 5.201e-09 1.849850879899086 5.202e-09 1.8325277327354847 5.2029999999999995e-09 1.7741626105273594 5.204e-09 1.7883868982968267 5.205e-09 1.8542324416452596 5.206e-09 1.767443279729199 5.207e-09 1.8179328904699292 5.208e-09 1.834649503026382 5.209e-09 1.8286726350451052 5.21e-09 1.784403715302959 5.211e-09 1.8585797874957983 5.212e-09 1.8396779961224692 5.213e-09 1.853016839037002 5.2139999999999996e-09 1.808286516237374 5.215e-09 1.7772124082299716 5.216e-09 1.7834093279336898 5.217e-09 1.8747692017326838 5.218e-09 1.9019280148495559 5.219e-09 1.7988606785101908 5.22e-09 1.7805270531341997 5.221e-09 1.7095561064739055 5.2219999999999995e-09 1.864523250712416 5.223e-09 1.7937187091482378 5.224e-09 1.7697456328722365 5.225e-09 1.7072905826919604 5.226e-09 1.8282919433712674 5.227e-09 1.817076504494871 5.228e-09 1.7788182471905436 5.229e-09 1.7607090436003845 5.2299999999999995e-09 1.8667217441245643 5.231e-09 1.8152579895715497 5.232e-09 1.8167009279654458 5.233e-09 1.8492612601438332 5.234e-09 1.759526261878357 5.235e-09 1.7808606688606534 5.236e-09 1.7430947343061922 5.237e-09 1.7628144907179146 5.2379999999999995e-09 1.8245468490014058 5.239e-09 1.8152818311197803 5.24e-09 1.8611861406220682 5.2409999999999996e-09 1.8413719500550116 5.242e-09 1.797891819273289 5.243e-09 1.77147828894306 5.244e-09 1.7895106296952359 5.245e-09 1.8095461311900964 5.246e-09 1.801644741242988 5.247e-09 1.8171899999363739 5.248e-09 1.9061464627201103 5.2489999999999996e-09 1.7764080939309495 5.25e-09 1.7629953533949076 5.251e-09 1.7265731522538472 5.252e-09 1.7961145099190827 5.253e-09 1.8539555119701605 5.254e-09 1.8176492085864304 5.255e-09 1.7981015494352972 5.256e-09 1.8124503455214285 5.2569999999999995e-09 1.9416977582944819 5.258e-09 1.8381599162367628 5.259e-09 1.818924281665604 5.26e-09 1.7570756757267167 5.261e-09 1.8302349778698732 5.262e-09 1.8923579833787239 5.263e-09 1.845807450151605 5.264e-09 1.8528272014987983 5.2649999999999995e-09 1.8468012355179162 5.266e-09 1.7012871715810904 5.267e-09 1.7689022781180208 5.268e-09 1.761219935006286 5.269e-09 1.7732887126187304 5.27e-09 1.775995457624072 5.271e-09 1.781504580699847 5.272e-09 1.7742334440346552 5.273e-09 1.7917682762149072 5.274e-09 1.8278146427214934 5.275e-09 1.7548307908173937 5.2759999999999996e-09 1.9341414056694122 5.277e-09 1.8070015783455036 5.278e-09 1.8163063399388266 5.279e-09 1.855074939812392 5.28e-09 1.842747155178841 5.281e-09 1.8290264277437387 5.282e-09 1.803859254582134 5.283e-09 1.7144962508271875 5.2839999999999995e-09 1.7786320417405865 5.285e-09 1.7708978756317368 5.286e-09 1.8361696248109356 5.287e-09 1.8709459619563227 5.288e-09 1.803210086317378 5.289e-09 1.8261788156452434 5.29e-09 1.8333912636470975 5.291e-09 1.8466931789555228 5.2919999999999995e-09 1.6897883699141178 5.293e-09 1.81319187101832 5.294e-09 1.781204117593357 5.295e-09 1.787782942831556 5.296e-09 1.720378593911835 5.297e-09 1.8786671861229867 5.298e-09 1.7739132410385265 5.299e-09 1.8209311963496684 5.2999999999999995e-09 1.8410324517694483 5.301e-09 1.7599429238910065 5.302e-09 1.7943751134071722 5.3029999999999996e-09 1.745413717569587 5.304e-09 1.832111258463196 5.305e-09 1.8855177610564176 5.306e-09 1.8252066605375064 5.307e-09 1.7994830251723826 5.308e-09 1.752502925237971 5.309e-09 1.8403840713452149 5.31e-09 1.794756128612954 5.3109999999999995e-09 1.862177847793925 5.312e-09 1.8318509969802308 5.313e-09 1.7720018352787243 5.314e-09 1.831479420154026 5.315e-09 1.7606770560907767 5.316e-09 1.790174940542841 5.317e-09 1.872434054164246 5.318e-09 1.8419667798022206 5.3189999999999995e-09 1.8275755375182818 5.32e-09 1.8442804042311565 5.321e-09 1.7563765548384977 5.322e-09 1.792938557788144 5.323e-09 1.7501439517514246 5.324e-09 1.7961073719367562 5.325e-09 1.8538722909844365 5.326e-09 1.8524295414033578 5.3269999999999995e-09 1.7914953771962248 5.328e-09 1.8390665379723452 5.329e-09 1.6894072998529654 5.3299999999999996e-09 1.7924371301651816 5.331e-09 1.8637974577612024 5.332e-09 1.7919287930901378 5.333e-09 1.8329566353939548 5.334e-09 1.7773957900420423 5.335e-09 1.8736669708117446 5.336e-09 1.7093817155249431 5.337e-09 1.7608890806567625 5.3379999999999996e-09 1.7869966869572265 5.339e-09 1.7821312812794987 5.34e-09 1.7586107521096574 5.341e-09 1.8180850203399954 5.342e-09 1.8358685141891342 5.343e-09 1.8300233361610572 5.344e-09 1.7917067117606333 5.345e-09 1.8215381630475032 5.3459999999999995e-09 1.7850525898787355 5.347e-09 1.8113752839624695 5.348e-09 1.797718271233125 5.349e-09 1.8262673129017308 5.35e-09 1.7005159234858205 5.351e-09 1.7758101370112913 5.352e-09 1.7839700658604398 5.353e-09 1.8875383559618995 5.3539999999999995e-09 1.6480616149793756 5.355e-09 1.8079587931939523 5.356e-09 1.8090651002950155 5.357e-09 1.7620455224862255 5.358e-09 1.7490954063655748 5.359e-09 1.852977147698775 5.36e-09 1.757053774247912 5.361e-09 1.7028261428506672 5.362e-09 1.7877662647457784 5.363e-09 1.7752198905169891 5.364e-09 1.8158190384046817 5.3649999999999996e-09 1.7646047995899328 5.366e-09 1.8421884716319412 5.367e-09 1.846491430574288 5.368e-09 1.8258909871146183 5.369e-09 1.8221723886233538 5.37e-09 1.8262874881163866 5.371e-09 1.814569895558657 5.372e-09 1.7945345162521573 5.3729999999999995e-09 1.854744471492222 5.374e-09 1.7808802169704492 5.375e-09 1.881874221719782 5.376e-09 1.8219387000243483 5.377e-09 1.7325609385792489 5.378e-09 1.754782759933031 5.379e-09 1.752598820577176 5.38e-09 1.8346747819598481 5.3809999999999995e-09 1.751935187659675 5.382e-09 1.847293697901253 5.383e-09 1.8319922747490223 5.384e-09 1.790434330285569 5.385e-09 1.7458771766584462 5.386e-09 1.7507347828990236 5.387e-09 1.8089209818546415 5.388e-09 1.8293865135424494 5.3889999999999995e-09 1.8192889193413266 5.39e-09 1.7635487151476807 5.391e-09 1.750792431201271 5.3919999999999996e-09 1.7814215365557804 5.393e-09 1.7452982730319306 5.394e-09 1.7841005551898477 5.395e-09 1.8075440973947268 5.396e-09 1.8207376569403009 5.397e-09 1.8277252858500823 5.398e-09 1.8176001401837816 5.399e-09 1.8698276338584905 5.3999999999999996e-09 1.8444325296531643 5.401e-09 1.7845179773912005 5.402e-09 1.7731552245403148 5.403e-09 1.8287007610052213 5.404e-09 1.8646695642225681 5.405e-09 1.7988145801307205 5.406e-09 1.8729536490063363 5.407e-09 1.7945164177993314 5.4079999999999995e-09 1.6891466157271717 5.409e-09 1.820325054849917 5.41e-09 1.9143727935118855 5.411e-09 1.8267448701842406 5.412e-09 1.888994641331831 5.413e-09 1.8753507933282976 5.414e-09 1.8418043769029935 5.415e-09 1.779976460561004 5.4159999999999995e-09 1.8814824951357925 5.417e-09 1.7661742290168594 5.418e-09 1.7917843124285318 5.419e-09 1.716556534695509 5.42e-09 1.7876952445081522 5.421e-09 1.7439438380344603 5.422e-09 1.7958559004183052 5.423e-09 1.8285812276917857 5.424e-09 1.7352738885021424 5.425e-09 1.813799759960211 5.426e-09 1.8636266892056763 5.4269999999999996e-09 1.735864383167227 5.428e-09 1.7836859408928627 5.429e-09 1.748489452010407 5.43e-09 1.8053356339038913 5.431e-09 1.7875380280562374 5.432e-09 1.8167396126681794 5.433e-09 1.766091248767178 5.434e-09 1.805094808886652 5.4349999999999995e-09 1.889479080720301 5.436e-09 1.787615182304654 5.437e-09 1.797698499844002 5.438e-09 1.8341578739344433 5.439e-09 1.8073656547595383 5.44e-09 1.931754190328233 5.441e-09 1.822419626070854 5.442e-09 1.8140065223855328 5.4429999999999995e-09 1.7973357762463067 5.444e-09 1.7818870563761764 5.445e-09 1.8163142572891966 5.446e-09 1.8030639330985365 5.447e-09 1.7890162876144768 5.448e-09 1.857462055661159 5.449e-09 1.8385062048375471 5.45e-09 1.8418730160826138 5.4509999999999995e-09 1.85366323220578 5.452e-09 1.8035378103943158 5.453e-09 1.8246941458225063 5.4539999999999996e-09 1.8267549672440482 5.455e-09 1.7683249855124799 5.456e-09 1.7856149253205644 5.457e-09 1.8044467087403635 5.458e-09 1.7990624569622071 5.459e-09 1.7769936584025106 5.46e-09 1.7928084662207047 5.461e-09 1.8450338388371377 5.4619999999999995e-09 1.7877616237156129 5.463e-09 1.8110465266079825 5.464e-09 1.802736457940206 5.465e-09 1.8590646562593638 5.466e-09 1.7444470985850482 5.467e-09 1.8614953789159985 5.468e-09 1.8075050562610153 5.469e-09 1.7498428451246315 5.4699999999999995e-09 1.853149336635916 5.471e-09 1.6197105763046915 5.472e-09 1.7560306281146385 5.473e-09 1.7521567680924321 5.474e-09 1.8620664003679588 5.475e-09 1.8592899302217754 5.476e-09 1.8572012633836064 5.477e-09 1.82167064053524 5.4779999999999995e-09 1.953298516274407 5.479e-09 1.8513793420996065 5.48e-09 1.7915504475112083 5.4809999999999996e-09 1.7778568553370497 5.482e-09 1.8832566210928041 5.483e-09 1.8947336711079008 5.484e-09 1.7838655164332933 5.485e-09 1.804907362520843 5.486e-09 1.7250722443205178 5.487e-09 1.814795370731238 5.488e-09 1.7282041869005282 5.4889999999999996e-09 1.8183572529068845 5.49e-09 1.8365396076435416 5.491e-09 1.8807399262810514 5.492e-09 1.8236535000235392 5.493e-09 1.8000896723623923 5.494e-09 1.839436773616336 5.495e-09 1.8499841097946994 5.496e-09 1.7944535656017606 5.4969999999999995e-09 1.8233979242902403 5.498e-09 1.7803276474718546 5.499e-09 1.7664352376244603 5.5e-09 1.8423263350292374 5.501e-09 1.82131952150212 5.502e-09 1.796582080486544 5.503e-09 1.8084791368579718 5.504e-09 1.7785861025673095 5.5049999999999995e-09 1.8368283516174833 5.506e-09 1.7090567123283265 5.507e-09 1.7925002863243487 5.508e-09 1.8595687519344752 5.509e-09 1.7638512198146432 5.51e-09 1.7967217290797626 5.511e-09 1.819450055456787 5.512e-09 1.781942531314255 5.513e-09 1.8506574621746688 5.514e-09 1.8982829324016048 5.515e-09 1.8025295472806424 5.5159999999999996e-09 1.8218590468375964 5.517e-09 1.7583226167839392 5.518e-09 1.748101581336653 5.519e-09 1.78010274578004 5.52e-09 1.714030071795216 5.521e-09 1.8015807630505214 5.522e-09 1.794229523468764 5.523e-09 1.76512717756847 5.5239999999999995e-09 1.82683224187814 5.525e-09 1.840909260872928 5.526e-09 1.79474641072278 5.527e-09 1.7747723135960694 5.528e-09 1.804228407833914 5.529e-09 1.7782859270959772 5.53e-09 1.824565043706244 5.531e-09 1.8197944772721022 5.5319999999999995e-09 1.7986675322630783 5.533e-09 1.7695889189894018 5.534e-09 1.776291873203073 5.535e-09 1.8214946767826519 5.536e-09 1.8504287005750792 5.537e-09 1.8072955786171718 5.538e-09 1.7343030978607274 5.539e-09 1.8964448379294454 5.5399999999999995e-09 1.7051770905044823 5.541e-09 1.7635835788377212 5.542e-09 1.7934610043834578 5.5429999999999996e-09 1.8423574556923898 5.544e-09 1.773670906249908 5.545e-09 1.8540810968594845 5.546e-09 1.777776609295583 5.547e-09 1.7726681659062897 5.548e-09 1.7122659224018153 5.549e-09 1.736171008217615 5.55e-09 1.7791644232131867 5.5509999999999995e-09 1.8368967872601196 5.552e-09 1.7396076519674044 5.553e-09 1.7726990109835132 5.554e-09 1.7998236668439767 5.555e-09 1.7105791470102971 5.556e-09 1.8030671487674166 5.557e-09 1.8381598529719638 5.558e-09 1.8144745146456078 5.5589999999999995e-09 1.8474100848360762 5.56e-09 1.835891006996061 5.561e-09 1.8450056394310257 5.562e-09 1.712012630196584 5.563e-09 1.888288125399718 5.564e-09 1.7803852066115478 5.565e-09 1.7714594501491663 5.566e-09 1.7971984430222225 5.5669999999999995e-09 1.8482509026978224 5.568e-09 1.8330457414922365 5.569e-09 1.8117436559662512 5.5699999999999996e-09 1.8009336177260102 5.571e-09 1.7291205953285191 5.572e-09 1.823450923970638 5.573e-09 1.7454147282908812 5.574e-09 1.7992311621177333 5.575e-09 1.7900393966136365 5.576e-09 1.808070530977259 5.577e-09 1.8233070823356046 5.5779999999999996e-09 1.7888231812904352 5.579e-09 1.812494649111924 5.58e-09 1.8727281315646858 5.581e-09 1.8189044174794238 5.582e-09 1.7868739157439801 5.583e-09 1.8266039232531084 5.584e-09 1.8175459398687155 5.585e-09 1.8603139634686081 5.5859999999999995e-09 1.768239102014744 5.587e-09 1.9150726472754316 5.588e-09 1.8169862473825542 5.589e-09 1.7306434442496883 5.59e-09 1.805882334875709 5.591e-09 1.8087290789156414 5.592e-09 1.766042109044546 5.593e-09 1.8907316493739674 5.5939999999999995e-09 1.8412409767492197 5.595e-09 1.7664461995680476 5.596e-09 1.727977739535166 5.597e-09 1.822752048420534 5.598e-09 1.772071132710114 5.599e-09 1.8048002527307683 5.6e-09 1.8187904235013936 5.601e-09 1.7264991383358217 5.602e-09 1.8211493369470682 5.603e-09 1.7896768407769694 5.604e-09 1.7607808598162928 5.6049999999999996e-09 1.91097073362534 5.606e-09 1.7713227732792716 5.607e-09 1.8516433968110952 5.608e-09 1.790840277510007 5.609e-09 1.7710128162545438 5.61e-09 1.7827853918890306 5.611e-09 1.7178402583356267 5.612e-09 1.807913415625039 5.6129999999999995e-09 1.795076085689594 5.614e-09 1.6693184830697718 5.615e-09 1.713539822282425 5.616e-09 1.7042912411852427 5.617e-09 1.8648124001639483 5.618e-09 1.8557657641091785 5.619e-09 1.8214273561064735 5.62e-09 1.7433640019400662 5.6209999999999995e-09 1.7240249214180883 5.622e-09 1.8404071464433531 5.623e-09 1.8657875780090998 5.624e-09 1.701953932795524 5.625e-09 1.7684443547503323 5.626e-09 1.7141776038160952 5.627e-09 1.8426490813725687 5.628e-09 1.8361116671672884 5.6289999999999995e-09 1.782402144202755 5.63e-09 1.7550825353042787 5.631e-09 1.794687206356073 5.6319999999999996e-09 1.7983894888131238 5.633e-09 1.7438283861305721 5.634e-09 1.864228942339781 5.635e-09 1.759381164261481 5.636e-09 1.8747638045081738 5.637e-09 1.8830068373669855 5.638e-09 1.788967010931491 5.639e-09 1.7037612932118524 5.6399999999999995e-09 1.9006698313992163 5.641e-09 1.8807649956520804 5.642e-09 1.830606312012736 5.643e-09 1.724747267540442 5.644e-09 1.89738378586364 5.645e-09 1.8380384854669125 5.646e-09 1.7820360882165998 5.647e-09 1.682622625809929 5.6479999999999995e-09 1.8091507068533812 5.649e-09 1.810231027152283 5.65e-09 1.7840125589189026 5.651e-09 1.8053564123054722 5.652e-09 1.8529123161488124 5.653e-09 1.8141111324493397 5.654e-09 1.8519303057150929 5.655e-09 1.8833607783947093 5.6559999999999995e-09 1.8001811165137536 5.657e-09 1.777671097298369 5.658e-09 1.8055194190298425 5.659e-09 1.8208038207614876 5.66e-09 1.7110724066798104 5.661e-09 1.7810256022755395 5.662e-09 1.7458751238806691 5.663e-09 1.8718207976203705 5.664e-09 1.8012995473719045 5.665e-09 1.835018853173317 5.666e-09 1.8517042443984482 5.6669999999999996e-09 1.7421288638642498 5.668e-09 1.8110977857976802 5.669e-09 1.7600283263660943 5.67e-09 1.8322173450985075 5.671e-09 1.777210457711851 5.672e-09 1.779578524815677 5.673e-09 1.7664934924912197 5.674e-09 1.919764137405297 5.6749999999999995e-09 1.7935516068260389 5.676e-09 1.7601877875461884 5.677e-09 1.8481940774686534 5.678e-09 1.7670852026041528 5.679e-09 1.864438304397663 5.68e-09 1.8531073642680596 5.681e-09 1.833172566899354 5.682e-09 1.7397921866695982 5.6829999999999995e-09 1.7625406477633179 5.684e-09 1.8047177597090873 5.685e-09 1.8439297247332114 5.686e-09 1.7604440477454115 5.687e-09 1.8507760334725936 5.688e-09 1.846905476774041 5.689e-09 1.7757673403687027 5.69e-09 1.759023606163802 5.6909999999999995e-09 1.7468466273498422 5.692e-09 1.7972276525584359 5.693e-09 1.7843559010257415 5.6939999999999996e-09 1.8350102798297399 5.695e-09 1.837866026630433 5.696e-09 1.7379851828814277 5.697e-09 1.795559203968653 5.698e-09 1.7535086598364804 5.699e-09 1.7705562183811008 5.7e-09 1.7042260421111854 5.701e-09 1.7539437692377504 5.7019999999999995e-09 1.8428675363310236 5.703e-09 1.8739504492391394 5.704e-09 1.7521374056262646 5.705e-09 1.7523340509194505 5.706e-09 1.9083584301359198 5.707e-09 1.921395592005486 5.708e-09 1.8140082843968235 5.709e-09 1.7320139163936792 5.7099999999999995e-09 1.777290975850761 5.711e-09 1.8257149561258759 5.712e-09 1.81414264449352 5.713e-09 1.9039699967951333 5.714e-09 1.7840714994109528 5.715e-09 1.7741757359120973 5.716e-09 1.7969597242652573 5.717e-09 1.8480772527274014 5.7179999999999995e-09 1.8068247569251863 5.719e-09 1.8465369810802135 5.72e-09 1.8490467601292289 5.7209999999999996e-09 1.7810084528573005 5.722e-09 1.822862246594403 5.723e-09 1.8378120913349878 5.724e-09 1.7640054033306158 5.725e-09 1.8491531444261977 5.726e-09 1.838614978804365 5.727e-09 1.8039250518871062 5.728e-09 1.7642566087783464 5.7289999999999996e-09 1.7155807767623854 5.73e-09 1.8230582974618312 5.731e-09 1.7495863123346842 5.732e-09 1.7211592484220335 5.733e-09 1.7885236465760446 5.734e-09 1.8738230397723494 5.735e-09 1.8719794329135115 5.736e-09 1.8133973824880767 5.7369999999999995e-09 1.7071485608975954 5.738e-09 1.7226850578150632 5.739e-09 1.8497545252086098 5.74e-09 1.8508561555795788 5.741e-09 1.8058032406718558 5.742e-09 1.7659377973510912 5.743e-09 1.8618360478493545 5.744e-09 1.7510663696491313 5.7449999999999995e-09 1.7894821761390662 5.746e-09 1.7438042712406636 5.747e-09 1.7720907191409374 5.748e-09 1.7999402517408085 5.749e-09 1.8173995617239282 5.75e-09 1.7880363698475141 5.751e-09 1.9192053229638375 5.752e-09 1.8760608415476376 5.753e-09 1.821310828760214 5.754e-09 1.7994493622620427 5.755e-09 1.8311672463786923 5.7559999999999996e-09 1.7924599712470866 5.757e-09 1.7402969352533864 5.758e-09 1.7944681266740607 5.759e-09 1.8472497066432274 5.76e-09 1.8099109954885335 5.761e-09 1.7250369139602457 5.762e-09 1.8599653629171826 5.763e-09 1.8026129053785651 5.7639999999999995e-09 1.7831203878765467 5.765e-09 1.7185271393147867 5.766e-09 1.7221726779637763 5.767e-09 1.8231970188235391 5.768e-09 1.8266764723358868 5.769e-09 1.7661491258932107 5.77e-09 1.8032909091222693 5.771e-09 1.7713473615514155 5.7719999999999995e-09 1.8383320774074179 5.773e-09 1.8396965205199902 5.774e-09 1.7597005766069989 5.775e-09 1.7187331387295224 5.776e-09 1.9084109383202554 5.777e-09 1.8559915592375602 5.778e-09 1.8769219443971874 5.779e-09 1.753481249996659 5.7799999999999995e-09 1.7679761467199162 5.781e-09 1.7470801282768345 5.782e-09 1.70088076755607 5.7829999999999996e-09 1.71958046301264 5.784e-09 1.796399812014154 5.785e-09 1.7614679048809434 5.786e-09 1.7847967033132537 5.787e-09 1.7654219514522718 5.788e-09 1.8621821159164682 5.789e-09 1.7832116095822712 5.79e-09 1.7992127208167932 5.7909999999999995e-09 1.8503129904226574 5.792e-09 1.7311079016196782 5.793e-09 1.8042473246891624 5.794e-09 1.802803977100875 5.795e-09 1.7314880923510496 5.796e-09 1.8420468185629961 5.797e-09 1.8092273873167977 5.798e-09 1.7620583721468683 5.7989999999999995e-09 1.7339039299990966 5.8e-09 1.7323956341396178 5.801e-09 1.8261500794924712 5.802e-09 1.7786148137739874 5.803e-09 1.8243446885506724 5.804e-09 1.9393323967109366 5.805e-09 1.721349081674183 5.806e-09 1.8253643582354313 5.8069999999999995e-09 1.8810122197959631 5.808e-09 1.8022766050786012 5.809e-09 1.833055883194034 5.8099999999999996e-09 1.837856700294735 5.811e-09 1.7637885687580224 5.812e-09 1.8151024783196608 5.813e-09 1.846889937683227 5.814e-09 1.9375855108290236 5.815e-09 1.8287890403326157 5.816e-09 1.8194110808468054 5.817e-09 1.795501474963553 5.8179999999999996e-09 1.7465689628667111 5.819e-09 1.8101295193687963 5.82e-09 1.8212157452890803 5.821e-09 1.7823871614262674 5.822e-09 1.844902404622344 5.823e-09 1.8522355851475685 5.824e-09 1.9073896136041475 5.825e-09 1.811770148264565 5.8259999999999995e-09 1.7597367654189455 5.827e-09 1.6763878725932533 5.828e-09 1.8472022234608312 5.829e-09 1.8326151302041318 5.83e-09 1.7752290354473483 5.831e-09 1.7725190974463265 5.832e-09 1.7487765543481786 5.833e-09 1.7633898844736389 5.8339999999999995e-09 1.8238813187951115 5.835e-09 1.8244251095170954 5.836e-09 1.7996179910230574 5.837e-09 1.807067713659363 5.838e-09 1.7165754827873905 5.839e-09 1.730520946948285 5.84e-09 1.6892198084045504 5.841e-09 1.7601622215266421 5.8419999999999995e-09 1.7525784219992828 5.843e-09 1.780424528058535 5.844e-09 1.7668454741694872 5.8449999999999996e-09 1.80577757035643 5.846e-09 1.895027451056116 5.847e-09 1.8650029946031645 5.848e-09 1.8059321091167406 5.849e-09 1.8653371316696368 5.85e-09 1.9220827609953066 5.851e-09 1.7327355854839062 5.852e-09 1.6891720829747323 5.8529999999999995e-09 1.7608583889536173 5.854e-09 1.8696708997930176 5.855e-09 1.8578437292074954 5.856e-09 1.8728448614192215 5.857e-09 1.7066589629246172 5.858e-09 1.7208785395413218 5.859e-09 1.7538788101175071 5.86e-09 1.7654853585890102 5.8609999999999995e-09 1.8345428828400991 5.862e-09 1.792005023581759 5.863e-09 1.8223984423775634 5.864e-09 1.7190690671842355 5.865e-09 1.7563957551907767 5.866e-09 1.806045046429489 5.867e-09 1.7631648213949591 5.868e-09 1.7483828976945508 5.8689999999999995e-09 1.8178315371697027 5.87e-09 1.7647157911767288 5.871e-09 1.7826444201775564 5.8719999999999996e-09 1.840686570940112 5.873e-09 1.847792601110599 5.874e-09 1.7994343839748852 5.875e-09 1.7836342235930738 5.876e-09 1.7169756105584137 5.877e-09 1.7571806407644204 5.878e-09 1.9358752098825056 5.879e-09 1.807965731735837 5.8799999999999995e-09 1.78822290239858 5.881e-09 1.7319403420111374 5.882e-09 1.7467074911219322 5.883e-09 1.7631661254543352 5.884e-09 1.7940469058587303 5.885e-09 1.7105403208936125 5.886e-09 1.8411035874915782 5.887e-09 1.7629838997579999 5.8879999999999995e-09 1.7502604095060337 5.889e-09 1.781617861974563 5.89e-09 1.795911715321045 5.891e-09 1.8560044554364088 5.892e-09 1.8584776971186816 5.893e-09 1.68144889542282 5.894e-09 1.7516910185128471 5.895e-09 1.8285034729805634 5.8959999999999995e-09 1.7362349622209177 5.897e-09 1.812621869394946 5.898e-09 1.7946481048899887 5.8989999999999996e-09 1.7721975354349664 5.9e-09 1.7487173335798087 5.901e-09 1.8575881444915396 5.902e-09 1.871772319319988 5.903e-09 1.7392064765738555 5.904e-09 1.838392820166192 5.905e-09 1.7713387221566304 5.906e-09 1.8035403295381922 5.9069999999999996e-09 1.7761957230895902 5.908e-09 1.7527206663464427 5.909e-09 1.7281510717586959 5.91e-09 1.789762647823191 5.911e-09 1.8236894711667577 5.912e-09 1.9148651979011424 5.913e-09 1.8139774081276139 5.914e-09 1.8866847628860948 5.9149999999999995e-09 1.7819576029933049 5.916e-09 1.815668467351432 5.917e-09 1.8706750836079171 5.918e-09 1.8201033780170066 5.919e-09 1.842164422777861 5.92e-09 1.8286599151222558 5.921e-09 1.8050530341318116 5.922e-09 1.831064454386081 5.9229999999999995e-09 1.80275986960653 5.924e-09 1.75741736229878 5.925e-09 1.78283798357874 5.926e-09 1.829041744310928 5.927e-09 1.7376181046073034 5.928e-09 1.781343184453302 5.929e-09 1.8273442565932785 5.93e-09 1.7778223118781438 5.9309999999999995e-09 1.6891219623098612 5.932e-09 1.724876263810868 5.933e-09 1.786422082121672 5.9339999999999996e-09 1.7532174536637317 5.935e-09 1.8832398777302706 5.936e-09 1.8030377133925073 5.937e-09 1.8123192633952854 5.938e-09 1.737335215961369 5.939e-09 1.8542317949549152 5.94e-09 1.8171613288606874 5.941e-09 1.775715842570111 5.9419999999999995e-09 1.7574801928447454 5.943e-09 1.7429739746730477 5.944e-09 1.8082000839433752 5.945e-09 1.8219610054414475 5.946e-09 1.836484086930578 5.947e-09 1.8346966834152671 5.948e-09 1.7791739520743324 5.949e-09 1.8245509774477264 5.9499999999999995e-09 1.8003543529259247 5.951e-09 1.8862679686697672 5.952e-09 1.7690683927167934 5.953e-09 1.8140657277638594 5.954e-09 1.7568135641166103 5.955e-09 1.7996487250950688 5.956e-09 1.7841867162379161 5.957e-09 1.7004664511356473 5.9579999999999995e-09 1.8070927070820793 5.959e-09 1.8840191376599962 5.96e-09 1.7965101818479674 5.9609999999999996e-09 1.8440656962856712 5.962e-09 1.789393337264102 5.963e-09 1.8645049487428955 5.964e-09 1.7425023952841137 5.965e-09 1.7828843738341986 5.966e-09 1.7850751570794945 5.967e-09 1.8405974533863991 5.968e-09 1.812058784471234 5.9689999999999996e-09 1.7886137828960502 5.97e-09 1.7702407378110483 5.971e-09 1.760268709967517 5.972e-09 1.7561771579188603 5.973e-09 1.8382774890755886 5.974e-09 1.7597422552781405 5.975e-09 1.8142557443072205 5.976e-09 1.8734662772718633 5.9769999999999995e-09 1.7454055286259287 5.978e-09 1.8116283951605243 5.979e-09 1.8263171657960167 5.98e-09 1.775185261257882 5.981e-09 1.7718039379337542 5.982e-09 1.8408636152409577 5.983e-09 1.7896312215946397 5.984e-09 1.9327199898841936 5.9849999999999995e-09 1.8088417311266618 5.986e-09 1.7802924017002035 5.987e-09 1.811000712756399 5.988e-09 1.798911632929004 5.989e-09 1.7336812304990874 5.99e-09 1.8048712319480886 5.991e-09 1.8249103785910294 5.992e-09 1.7868480053189526 5.9929999999999995e-09 1.8344028066147557 5.994e-09 1.7840684411654733 5.995e-09 1.7157151050618187 5.9959999999999996e-09 1.7639914777999075 5.997e-09 1.7586689655869225 5.998e-09 1.7208668794967932 5.999e-09 1.8847446077145824 6e-09 1.7824639027205122 6.001e-09 1.7960485443815404 6.002e-09 1.8077411122236258 6.003e-09 1.8310264915748267 6.0039999999999995e-09 1.7384058310725417 6.005e-09 1.8184102871031822 6.006e-09 1.7849931080154997 6.007e-09 1.7843273299969058 6.008e-09 1.6837308143699108 6.009e-09 1.728896357091126 6.01e-09 1.7493157649064408 6.011e-09 1.7871397250569399 6.0119999999999995e-09 1.802583880148273 6.013e-09 1.8776786849763303 6.014e-09 1.8515806617124602 6.015e-09 1.8517161336383994 6.016e-09 1.7041875421975718 6.017e-09 1.7888540389492367 6.018e-09 1.7753897841146102 6.019e-09 1.7825263867070202 6.0199999999999995e-09 1.7374322501512591 6.021e-09 1.8548612323750582 6.022e-09 1.7629731793371028 6.0229999999999996e-09 1.8029619997092483 6.024e-09 1.8219410619319962 6.025e-09 1.9047543449126576 6.026e-09 1.6412651515017527 6.027e-09 1.8115106950405782 6.028e-09 1.8167906168206818 6.029e-09 1.8794650371875485 6.03e-09 1.8435724138540306 6.0309999999999995e-09 1.8435376760339584 6.032e-09 1.7625777770579396 6.033e-09 1.8486924308384876 6.034e-09 1.737595236458447 6.035e-09 1.725820974749392 6.036e-09 1.8460646369485263 6.037e-09 1.7522322609701204 6.038e-09 1.7584967184719438 6.0389999999999995e-09 1.7891929887772386 6.04e-09 1.8063571944546049 6.041e-09 1.691896763456652 6.042e-09 1.761071520480275 6.043e-09 1.7516791117347792 6.044e-09 1.7782844589598006 6.045e-09 1.8061248906184801 6.046e-09 1.7976211535187108 6.0469999999999995e-09 1.846582304841519 6.048e-09 1.7259622030449386 6.049e-09 1.7443325902908617 6.0499999999999996e-09 1.8887818083242283 6.051e-09 1.8624047418001881 6.052e-09 1.7513950573062071 6.053e-09 1.8078529337766214 6.054e-09 1.7302195470694532 6.055e-09 1.8153986556547164 6.056e-09 1.756450004514507 6.057e-09 1.7349278741504004 6.0579999999999996e-09 1.860497387362103 6.059e-09 1.8243574631468262 6.06e-09 1.7853532845963829 6.061e-09 1.806251592391252 6.062e-09 1.7990273571879154 6.063e-09 1.8619185987075695 6.064e-09 1.8331495458100275 6.065e-09 1.7638686740622684 6.0659999999999995e-09 1.8436698059466794 6.067e-09 1.7803597921418126 6.068e-09 1.8293362672560665 6.069e-09 1.8643771302999819 6.07e-09 1.8919771571087902 6.071e-09 1.7384997254715069 6.072e-09 1.7699844497257309 6.073e-09 1.6903225052343869 6.0739999999999995e-09 1.7653926215084506 6.075e-09 1.7808057034413742 6.076e-09 1.8256321722183309 6.077e-09 1.839732630632204 6.078e-09 1.7001594989301556 6.079e-09 1.8138547841109092 6.08e-09 1.8118934165109042 6.081e-09 1.782257875466488 6.0819999999999995e-09 1.7213638070263533 6.083e-09 1.756216504671035 6.084e-09 1.8276765211467216 6.0849999999999996e-09 1.8173625681459369 6.086e-09 1.8211939984493055 6.087e-09 1.843090165108741 6.088e-09 1.8098712683419127 6.089e-09 1.8243238990954107 6.09e-09 1.817493644640454 6.091e-09 1.8026284884915384 6.092e-09 1.8261621270670827 6.0929999999999995e-09 1.8406161089872548 6.094e-09 1.7735887469059726 6.095e-09 1.801165820514737 6.096e-09 1.7732979183138515 6.097e-09 1.8467892059883615 6.098e-09 1.8929158798812877 6.099e-09 1.751626645088695 6.1e-09 1.8393507469521324 6.1009999999999995e-09 1.7969227609608738 6.102e-09 1.8782044638505382 6.103e-09 1.8105315962045399 6.104e-09 1.7277044825785663 6.105e-09 1.826335082371423 6.106e-09 1.8230003704980582 6.107e-09 1.7585694045269862 6.108e-09 1.8149074815999584 6.1089999999999995e-09 1.8862743116931173 6.11e-09 1.8315133532628296 6.111e-09 1.7886522583170616 6.1119999999999996e-09 1.8604752630941404 6.113e-09 1.7507915965631953 6.114e-09 1.8117699328637267 6.115e-09 1.7980533279332012 6.116e-09 1.7954597196740736 6.117e-09 1.8079091469520387 6.118e-09 1.809718076932344 6.119e-09 1.818667279308284 6.1199999999999995e-09 1.8263391505015802 6.121e-09 1.9321315580186549 6.122e-09 1.848047434015143 6.123e-09 1.7337806957413762 6.124e-09 1.761180962653991 6.125e-09 1.8021372396908772 6.126e-09 1.822346523802485 6.127e-09 1.737324176550831 6.1279999999999995e-09 1.7491902867380855 6.129e-09 1.7910443472198627 6.13e-09 1.8934223856925665 6.131e-09 1.818743472068674 6.132e-09 1.8292124887229406 6.133e-09 1.8238719265138954 6.134e-09 1.8074014549078719 6.135e-09 1.8126903752438748 6.1359999999999995e-09 1.7720991754330035 6.137e-09 1.7849326891470063 6.138e-09 1.7902050913921044 6.1389999999999996e-09 1.8645927294787752 6.14e-09 1.769200638745107 6.141e-09 1.7977640164550681 6.142e-09 1.7790921587463924 6.143e-09 1.8343966984379583 6.144e-09 1.7947126937048126 6.145e-09 1.8713891482263483 6.146e-09 1.6770845548946356 6.1469999999999996e-09 1.7857176696109416 6.148e-09 1.8042765855476726 6.149e-09 1.8130913090191985 6.15e-09 1.7137834695519079 6.151e-09 1.7113021905101096 6.152e-09 1.7432601766115456 6.153e-09 1.7464232184222725 6.154e-09 1.793712709790415 6.1549999999999995e-09 1.766417675126457 6.156e-09 1.8644671390299759 6.157e-09 1.7702311429756667 6.158e-09 1.905038029632895 6.159e-09 1.8365449286449926 6.16e-09 1.846785666880582 6.161e-09 1.7601997641389886 6.162e-09 1.7997728722327986 6.1629999999999995e-09 1.808666314104089 6.164e-09 1.7217832498015313 6.165e-09 1.8354344947905175 6.166e-09 1.88150744181337 6.167e-09 1.797356137123217 6.168e-09 1.7761898077024398 6.169e-09 1.772381968732348 6.17e-09 1.7859054188574541 6.1709999999999995e-09 1.7697206109697738 6.172e-09 1.7692425836163248 6.173e-09 1.7585717322568863 6.1739999999999996e-09 1.8297830533031378 6.175e-09 1.7729248122970542 6.176e-09 1.7898157696494181 6.177e-09 1.867744372100297 6.178e-09 1.8563167567783896 6.179e-09 1.8145263253180486 6.18e-09 1.817211085755058 6.181e-09 1.820752777423632 6.1819999999999995e-09 1.8321743368811558 6.183e-09 1.8402991944467328 6.184e-09 1.7577594764315116 6.185e-09 1.787920155978242 6.186e-09 1.7974914794030377 6.187e-09 1.6748339798510796 6.188e-09 1.7722071443642706 6.189e-09 1.829599208960182 6.1899999999999995e-09 1.8183170461810392 6.191e-09 1.8523109315189517 6.192e-09 1.755655413462606 6.193e-09 1.8473951749011863 6.194e-09 1.81338714770946 6.195e-09 1.6303987504297746 6.196e-09 1.8643170503206985 6.197e-09 1.7582428703529416 6.1979999999999995e-09 1.7933778187052594 6.199e-09 1.7047311659519948 6.2e-09 1.818050832076376 6.2009999999999996e-09 1.7986886170541514 6.202e-09 1.740758749631812 6.203e-09 1.8665675432649667 6.204e-09 1.7677197268619003 6.205e-09 1.7611667057453375 6.206e-09 1.8609870628501273 6.207e-09 1.8404710520446759 6.208e-09 1.8351733997064124 6.2089999999999995e-09 1.8107803810496546 6.21e-09 1.837222097995097 6.211e-09 1.7641370371542289 6.212e-09 1.7543757227821632 6.213e-09 1.8208495196776016 6.214e-09 1.7351510572960702 6.215e-09 1.753163275089296 6.216e-09 1.7924708701077021 6.2169999999999995e-09 1.7482753110079603 6.218e-09 1.861029385103163 6.219e-09 1.8600346479220455 6.22e-09 1.7812991979186021 6.221e-09 1.7989040682528705 6.222e-09 1.8910987189771147 6.223e-09 1.7667467484779376 6.224e-09 1.8637761363873773 6.2249999999999995e-09 1.8609300421515964 6.226e-09 1.7740947563525717 6.227e-09 1.8071813502696776 6.2279999999999996e-09 1.7350369815773745 6.229e-09 1.801630738388885 6.23e-09 1.791881064590499 6.231e-09 1.812445888586583 6.232e-09 1.7417130187236536 6.2329999999999995e-09 1.7722235201650798 6.234e-09 1.8086542201841171 6.235e-09 1.8463143463561207 6.2359999999999996e-09 1.7713275895535898 6.237e-09 1.7313284393950832 6.238e-09 1.8365630557151265 6.239e-09 1.819159703892867 6.24e-09 1.7451209400698076 6.241e-09 1.91706902203636 6.242e-09 1.7542788026759086 6.243e-09 1.754755331594661 6.2439999999999995e-09 1.887406592764994 6.245e-09 1.808382694368498 6.246e-09 1.7883637834116217 6.247e-09 1.8151733079498822 6.248e-09 1.8085297825471214 6.249e-09 1.7679230935813948 6.25e-09 1.8671086267873582 6.251e-09 1.81478555901455 6.2519999999999995e-09 1.8139878136964762 6.253e-09 1.8304658562982528 6.254e-09 1.8240886631095627 6.255e-09 1.761846852013103 6.256e-09 1.8529832890667637 6.257e-09 1.7582837923016923 6.258e-09 1.7480205234962307 6.259e-09 1.7701768111804748 6.2599999999999995e-09 1.8745860582907732 6.261e-09 1.7347488080091793 6.262e-09 1.7521405111255015 6.2629999999999996e-09 1.7733563971040291 6.264e-09 1.723162279949302 6.265e-09 1.8395906349588669 6.266e-09 1.687153206975914 6.267e-09 1.8297739632699022 6.268e-09 1.8390299240611057 6.269e-09 1.6750505649969276 6.27e-09 1.832208960617958 6.2709999999999995e-09 1.786294653192085 6.272e-09 1.8740541499077772 6.273e-09 1.8840381350187483 6.274e-09 1.8090565479984244 6.275e-09 1.8191057674310076 6.276e-09 1.8689071238322996 6.277e-09 1.7455021256012029 6.278e-09 1.68881269430246 6.2789999999999995e-09 1.8176668290431124 6.28e-09 1.7976520670587028 6.281e-09 1.8071213772072794 6.282e-09 1.8466952896991045 6.283e-09 1.7744770770617773 6.284e-09 1.865742797827867 6.285e-09 1.841138128677556 6.286e-09 1.7925362373253828 6.2869999999999995e-09 1.7846666458764522 6.288e-09 1.760369896919397 6.289e-09 1.8703287786877334 6.2899999999999996e-09 1.754073387163817 6.291e-09 1.891606832070809 6.292e-09 1.8475034863243085 6.293e-09 1.8256454690505806 6.294e-09 1.8272237402476352 6.295e-09 1.797589649251576 6.296e-09 1.7283773260358994 6.297e-09 1.8101816257966101 6.2979999999999996e-09 1.8092352575156199 6.299e-09 1.84126301264458 6.3e-09 1.7899445426544298 6.301e-09 1.825716846076356 6.302e-09 1.6914109553488719 6.303e-09 1.709816730782065 6.304e-09 1.8083471657110477 6.305e-09 1.8056806765736122 6.3059999999999995e-09 1.7361309576193915 6.307e-09 1.8357529970655684 6.308e-09 1.830671320767674 6.309e-09 1.7936609035943507 6.31e-09 1.83828183571003 6.311e-09 1.906800141808463 6.312e-09 1.8000116753700235 6.313e-09 1.7225941087315104 6.3139999999999995e-09 1.7227515062610093 6.315e-09 1.857741407325504 6.316e-09 1.798337319712169 6.317e-09 1.7932105760132784 6.318e-09 1.756400754102746 6.319e-09 1.890299828470594 6.32e-09 1.8201196055639204 6.321e-09 1.6936731186833063 6.3219999999999995e-09 1.8147259380534757 6.323e-09 1.7971357024927554 6.324e-09 1.831454390693738 6.3249999999999996e-09 1.8825577587208733 6.326e-09 1.7941069684017383 6.327e-09 1.780819971786566 6.328e-09 1.8234109814757722 6.329e-09 1.7548322669285439 6.33e-09 1.7263199518705918 6.331e-09 1.8472876243876657 6.332e-09 1.7470513938481684 6.3329999999999995e-09 1.862608679390951 6.334e-09 1.7723112590943195 6.335e-09 1.7048799974684132 6.336e-09 1.8273191954691925 6.337e-09 1.8041386307815896 6.338e-09 1.8069774053341414 6.339e-09 1.7717059819976766 6.34e-09 1.8244144311744062 6.3409999999999995e-09 1.7765046106214997 6.342e-09 1.8298860673962523 6.343e-09 1.778745148836656 6.344e-09 1.807657446309042 6.345e-09 1.7625244138487635 6.346e-09 1.7429916542072281 6.347e-09 1.842534259611778 6.348e-09 1.8412320904687018 6.3489999999999995e-09 1.8877597591239392 6.35e-09 1.7828984170769577 6.351e-09 1.7592106182423972 6.3519999999999996e-09 1.7779769806082344 6.353e-09 1.7460932899459423 6.354e-09 1.7683145373730915 6.355e-09 1.8064443787485174 6.356e-09 1.8577507654125005 6.357e-09 1.7734889730449601 6.358e-09 1.7601575058590715 6.359e-09 1.8752250365977639 6.3599999999999995e-09 1.7789925257307106 6.361e-09 1.8626067826804165 6.362e-09 1.8161313263218863 6.363e-09 1.8478852307569342 6.364e-09 1.8281738993863026 6.365e-09 1.8065163494683814 6.366e-09 1.8038569141952692 6.367e-09 1.8361688461413312 6.3679999999999995e-09 1.7614122285257399 6.369e-09 1.7866802614248742 6.37e-09 1.822790170353462 6.371e-09 1.8065745729091698 6.372e-09 1.80553644014024 6.373e-09 1.8155419461439044 6.374e-09 1.8426145581777909 6.375e-09 1.7592802482193872 6.3759999999999995e-09 1.7810079805521681 6.377e-09 1.810626345213337 6.378e-09 1.846272741083408 6.3789999999999996e-09 1.8426083872493324 6.38e-09 1.8885484022144108 6.381e-09 1.73292813463111 6.382e-09 1.8211413011129445 6.383e-09 1.72184079425274 6.3839999999999995e-09 1.731920437127652 6.385e-09 1.7841333253981804 6.386e-09 1.786675635442897 6.3869999999999996e-09 1.7239614692932401 6.388e-09 1.7458099746235272 6.389e-09 1.7617945364283238 6.39e-09 1.9247874401889589 6.391e-09 1.762945303401766 6.392e-09 1.8667836093766244 6.393e-09 1.8607187166296946 6.394e-09 1.8159873277973908 6.3949999999999995e-09 1.8692303449354706 6.396e-09 1.8678621702431522 6.397e-09 1.801561166086476 6.398e-09 1.7806580430513415 6.399e-09 1.7172200997963938 6.4e-09 1.6758436160312156 6.401e-09 1.8147168438771424 6.402e-09 1.7792840246437818 6.4029999999999995e-09 1.771629926316711 6.404e-09 1.781025386063038 6.405e-09 1.890643103222357 6.406e-09 1.808979183179443 6.407e-09 1.6875810904300508 6.408e-09 1.8472851000610802 6.409e-09 1.767906400884727 6.41e-09 1.792478833702227 6.4109999999999995e-09 1.8696618678204522 6.412e-09 1.8077865738432026 6.413e-09 1.782924275974879 6.4139999999999996e-09 1.7403231524924963 6.415e-09 1.8060418786505217 6.416e-09 1.774241801850596 6.417e-09 1.8379800875109331 6.418e-09 1.7164138432336544 6.419e-09 1.7027294272247033 6.42e-09 1.829135081021152 6.421e-09 1.7494444828477116 6.4219999999999995e-09 1.8059346792959776 6.423e-09 1.8610238429003918 6.424e-09 1.7368445868368376 6.425e-09 1.8066126187787102 6.426e-09 1.7415025289880828 6.427e-09 1.8754060672229675 6.428e-09 1.8338431937469184 6.429e-09 1.9092341040800984 6.4299999999999995e-09 1.8227117727048983 6.431e-09 1.9647825508128156 6.432e-09 1.8169582104121216 6.433e-09 1.8422281691599993 6.434e-09 1.7957212928805335 6.435e-09 1.8510037599845284 6.436e-09 1.7847162511213426 6.437e-09 1.782121620437992 6.4379999999999995e-09 1.85646760185046 6.439e-09 1.7507763860241985 6.44e-09 1.8539339482920356 6.4409999999999996e-09 1.7764808137615369 6.442e-09 1.7538015507163764 6.443e-09 1.6656405802847074 6.444e-09 1.738086055617792 6.445e-09 1.8437162014361834 6.446e-09 1.7696717328782614 6.447e-09 1.7791116532063407 6.448e-09 1.7913546622673189 6.4489999999999995e-09 1.789837959596101 6.45e-09 1.7662832331426965 6.451e-09 1.7996223197573507 6.452e-09 1.899066924131991 6.453e-09 1.7440597367526738 6.454e-09 1.7412980181041107 6.455e-09 1.7565360782868116 6.456e-09 1.8219120170583478 6.4569999999999995e-09 1.8429140144953464 6.458e-09 1.7673314649162248 6.459e-09 1.8121111985058265 6.46e-09 1.8318778002248655 6.461e-09 1.7923147341217573 6.462e-09 1.8077188597300082 6.463e-09 1.8507536834356908 6.464e-09 1.8176272419100308 6.4649999999999995e-09 1.819123195320744 6.466e-09 1.8003316761002077 6.467e-09 1.8360422653720276 6.4679999999999996e-09 1.824633266569243 6.469e-09 1.7192756030093426 6.47e-09 1.8885821914556724 6.471e-09 1.7317941836390256 6.472e-09 1.7977258071919833 6.4729999999999995e-09 1.8440822413944142 6.474e-09 1.8074384451563579 6.475e-09 1.8345546590734356 6.4759999999999996e-09 1.8061613861163954 6.477e-09 1.8456391319438177 6.478e-09 1.7532014328013747 6.479e-09 1.762830634487874 6.48e-09 1.8019917093686486 6.481e-09 1.762883293098517 6.482e-09 1.7980719414388764 6.483e-09 1.7370474932623727 6.4839999999999995e-09 1.910354763923921 6.485e-09 1.87855432571142 6.486e-09 1.8543024469792928 6.487e-09 1.7575098358232493 6.488e-09 1.9337390266035692 6.489e-09 1.8625047768203329 6.49e-09 1.7900336818337825 6.491e-09 1.7564826749113656 6.4919999999999995e-09 1.743747952473374 6.493e-09 1.9040139073989772 6.494e-09 1.8199320549518911 6.495e-09 1.6971256508410364 6.496e-09 1.8100189257329125 6.497e-09 1.7608231989614662 6.498e-09 1.7574291313903876 6.499e-09 1.8064503514783252 6.4999999999999995e-09 1.804742980277684 6.501e-09 1.710747718285092 6.502e-09 1.8251430406117168 6.5029999999999996e-09 1.7957886295564673 6.504e-09 1.795920890382956 6.505e-09 1.7364159087976359 6.506e-09 1.8567988400685833 6.507e-09 1.772635425564645 6.508e-09 1.8050854616055347 6.509e-09 1.7725263333088823 6.51e-09 1.7480302330449677 6.5109999999999995e-09 1.7918096227889226 6.512e-09 1.7696729029345248 6.513e-09 1.7890299254114221 6.514e-09 1.8580095720658212 6.515e-09 1.770808402145008 6.516e-09 1.7868334043690393 6.517e-09 1.7631772034899613 6.518e-09 1.8370558687007037 6.5189999999999995e-09 1.6912262205718958 6.52e-09 1.8912482478258104 6.521e-09 1.7887937319371012 6.522e-09 1.846374944410294 6.523e-09 1.8251785934389004 6.524e-09 1.7409550985147397 6.525e-09 1.8578367209815816 6.526e-09 1.7536408562722003 6.5269999999999995e-09 1.7867673169745393 6.528e-09 1.7376416627031277 6.529e-09 1.7965804506218246 6.5299999999999996e-09 1.8387863434371765 6.531e-09 1.7734821795012405 6.532e-09 1.8570265885424002 6.533e-09 1.7527224195687674 6.534e-09 1.8189352836717692 6.5349999999999995e-09 1.7844122055286873 6.536e-09 1.7696077833611248 6.537e-09 1.7961629010641769 6.5379999999999995e-09 1.8086419947328576 6.539e-09 1.7525392733904972 6.54e-09 1.8192391514848094 6.541e-09 1.8501225027745065 6.542e-09 1.695297044792578 6.543e-09 1.8429918469293245 6.544e-09 1.745643229191762 6.545e-09 1.700738150044179 6.5459999999999995e-09 1.84278132166212 6.547e-09 1.8458653776458251 6.548e-09 1.832924156991254 6.549e-09 1.838855076322118 6.55e-09 1.749655760464879 6.551e-09 1.7434895580411163 6.552e-09 1.8720238259607282 6.553e-09 1.7763282354521925 6.5539999999999995e-09 1.8577625650906744 6.555e-09 1.7267702690265263 6.556e-09 1.7916084251699522 6.557e-09 1.6952317993335793 6.558e-09 1.7941188390597456 6.559e-09 1.7288163289857152 6.56e-09 1.8221170782726188 6.561e-09 1.7904588361044347 6.5619999999999995e-09 1.750544746274496 6.563e-09 1.7921543887420577 6.564e-09 1.769543433747776 6.5649999999999996e-09 1.7366434565315672 6.566e-09 1.7946105947122883 6.567e-09 1.841074759871959 6.568e-09 1.9030200994462132 6.569e-09 1.7322188650671304 6.57e-09 1.8340446451211372 6.571e-09 1.774494414010541 6.572e-09 1.8046768836247244 6.5729999999999995e-09 1.8544768047063247 6.574e-09 1.8026419367103652 6.575e-09 1.7620044759599316 6.576e-09 1.7197458809088524 6.577e-09 1.7516931528156094 6.578e-09 1.8644578904812699 6.579e-09 1.7451846239213578 6.58e-09 1.794791233592903 6.5809999999999995e-09 1.8787768072506905 6.582e-09 1.8398055041303971 6.583e-09 1.7720201101223831 6.584e-09 1.7578014669167352 6.585e-09 1.8322781539468698 6.586e-09 1.824097705694769 6.587e-09 1.845099666465297 6.588e-09 1.8251702423878036 6.5889999999999995e-09 1.8611365392767747 6.59e-09 1.9158998198985446 6.591e-09 1.8312412646881429 6.5919999999999996e-09 1.7890937671946703 6.593e-09 1.8342731731947564 6.594e-09 1.9179634071085514 6.595e-09 1.758507006656465 6.596e-09 1.9132273733282443 6.597e-09 1.8208633572709303 6.598e-09 1.7818332810246724 6.599e-09 1.7204862605993743 6.5999999999999995e-09 1.7716293266779617 6.601e-09 1.791913917440645 6.602e-09 1.724254097012992 6.603e-09 1.8527499379246382 6.604e-09 1.750281825971871 6.605e-09 1.72679130427189 6.606e-09 1.802311677049972 6.607e-09 1.7751796599533185 6.6079999999999995e-09 1.746202439275145 6.609e-09 1.7511154400331228 6.61e-09 1.7793128593112446 6.611e-09 1.8313063674439636 6.612e-09 1.838429773952155 6.613e-09 1.7987635578443006 6.614e-09 1.8596372768623324 6.615e-09 1.7475667646692858 6.6159999999999995e-09 1.8367278018773172 6.617e-09 1.8091723627199199 6.618e-09 1.7218686952165176 6.6189999999999996e-09 1.9050227017304229 6.62e-09 1.8641870905387137 6.621e-09 1.7869710012375926 6.622e-09 1.8795814946624447 6.623e-09 1.767181289840411 6.6239999999999995e-09 1.8635512069320395 6.625e-09 1.7354764687506772 6.626e-09 1.8394134959840465 6.6269999999999996e-09 1.7219387824767198 6.628e-09 1.7741849688580433 6.629e-09 1.6937496718161267 6.63e-09 1.78883234900511 6.631e-09 1.8124786037463554 6.632e-09 1.7392999308825443 6.633e-09 1.79975781199548 6.634e-09 1.818517334218692 6.6349999999999995e-09 1.7873266048317338 6.636e-09 1.7562098593474753 6.637e-09 1.8507381561373726 6.638e-09 1.7799768985828976 6.639e-09 1.8059738521462765 6.64e-09 1.7890015122078746 6.641e-09 1.7091472818457234 6.642e-09 1.791401154398458 6.6429999999999995e-09 1.7668179783811042 6.644e-09 1.736627852507552 6.645e-09 1.8184549970299424 6.646e-09 1.8093302109854743 6.647e-09 1.7732330504305038 6.648e-09 1.7804110781601006 6.649e-09 1.8168602835147203 6.65e-09 1.8991369827507045 6.6509999999999995e-09 1.7668444733317232 6.652e-09 1.7337542509788384 6.653e-09 1.7517069884498702 6.6539999999999996e-09 1.7882887973801562 6.655e-09 1.8281704870625357 6.656e-09 1.7672568268721343 6.657e-09 1.796111209077217 6.658e-09 1.722045928888525 6.659e-09 1.8227871100391924 6.66e-09 1.794001570954898 6.661e-09 1.8598608001685235 6.6619999999999995e-09 1.8075326777207894 6.663e-09 1.7952913777778254 6.664e-09 1.8266211760704838 6.665e-09 1.7516809835502258 6.666e-09 1.7316132198726533 6.667e-09 1.8268073878635644 6.668e-09 1.7866056853847254 6.669e-09 1.8011883874120096 6.6699999999999995e-09 1.7769518017564494 6.671e-09 1.8128189250185125 6.672e-09 1.8441433655625992 6.673e-09 1.731504504481756 6.674e-09 1.7748115144334708 6.675e-09 1.8671595478564402 6.676e-09 1.771866951896934 6.677e-09 1.826440226770238 6.6779999999999995e-09 1.747438376234554 6.679e-09 1.82885817111718 6.68e-09 1.8196109401824216 6.6809999999999996e-09 1.7899393202269822 6.682e-09 1.8464886136485403 6.683e-09 1.8149900718585739 6.684e-09 1.7034812809717181 6.685e-09 1.7622691023297201 6.6859999999999995e-09 1.8014683579228479 6.687e-09 1.8759481765922608 6.688e-09 1.8403825121906534 6.6889999999999995e-09 1.7852477663644795 6.69e-09 1.8539738010005709 6.691e-09 1.7234129922370924 6.692e-09 1.7845616483341917 6.693e-09 1.7667058777203302 6.694e-09 1.8302273874150752 6.695e-09 1.726435925516232 6.696e-09 1.7934710714542301 6.6969999999999995e-09 1.8164200832925514 6.698e-09 1.6987127618369025 6.699e-09 1.7989677344000905 6.7e-09 1.8506273191345284 6.701e-09 1.754121046598526 6.702e-09 1.7744973983502828 6.703e-09 1.747680462313103 6.704e-09 1.8877967007112442 6.7049999999999995e-09 1.8410288387855447 6.706e-09 1.7596794547508088 6.707e-09 1.754297240223952 6.7079999999999996e-09 1.857541021469727 6.709e-09 1.8655667414155894 6.71e-09 1.7249571304554618 6.711e-09 1.7894646111454464 6.712e-09 1.8577449521221405 6.7129999999999995e-09 1.853464330652295 6.714e-09 1.8154245524391097 6.715e-09 1.8590121840561067 6.7159999999999996e-09 1.6948105664259523 6.717e-09 1.8037865677120637 6.718e-09 1.8303267584026919 6.719e-09 1.685916317403167 6.72e-09 1.8197741218964363 6.721e-09 1.8234416512182043 6.722e-09 1.8127991734091429 6.723e-09 1.752043642858096 6.7239999999999995e-09 1.82272330345026 6.725e-09 1.7859411061271566 6.726e-09 1.7504673172825334 6.727e-09 1.8205574410923593 6.728e-09 1.7935682266251936 6.729e-09 1.8536817535125938 6.73e-09 1.8375442523551766 6.731e-09 1.7448998337471253 6.7319999999999995e-09 1.7979060384657468 6.733e-09 1.7785253282179547 6.734e-09 1.7971408896892243 6.735e-09 1.8909365277724455 6.736e-09 1.7852226798450952 6.737e-09 1.8044192085725763 6.738e-09 1.7810333482235217 6.739e-09 1.8536411798331698 6.7399999999999995e-09 1.8162713674430337 6.741e-09 1.9215918353319934 6.742e-09 1.8415366862901899 6.7429999999999996e-09 1.722560508203709 6.744e-09 1.7995585740693876 6.745e-09 1.802869446788294 6.746e-09 1.864894408321543 6.747e-09 1.763392947118135 6.748e-09 1.8550088291194013 6.749e-09 1.7437080623285655 6.75e-09 1.839952028182226 6.7509999999999995e-09 1.7054952019086254 6.752e-09 1.7438344931084706 6.753e-09 1.8075067115246508 6.754e-09 1.6791588165440237 6.755e-09 1.8744801342838577 6.756e-09 1.7594671003056712 6.757e-09 1.8596058255456258 6.758e-09 1.8904047280134717 6.7589999999999995e-09 1.7500520549796075 6.76e-09 1.7858286353469517 6.761e-09 1.7162531888315327 6.762e-09 1.8460706282122996 6.763e-09 1.8496708976819964 6.764e-09 1.778109623853342 6.765e-09 1.8654981454312674 6.766e-09 1.7935028874792334 6.7669999999999995e-09 1.7850348311979336 6.768e-09 1.8219993335024705 6.769e-09 1.7638984445784067 6.7699999999999996e-09 1.8067420660887896 6.771e-09 1.7474765088602668 6.772e-09 1.7183429009826827 6.773e-09 1.7633683140340108 6.774e-09 1.8853939834129867 6.7749999999999995e-09 1.8458100829012631 6.776e-09 1.7697697369861143 6.777e-09 1.814218911341093 6.7779999999999995e-09 1.843961750056626 6.779e-09 1.874746634745973 6.78e-09 1.7789316906251305 6.781e-09 1.7368520479218637 6.782e-09 1.8767240548134678 6.783e-09 1.8386870738559555 6.784e-09 1.8016308488132171 6.785e-09 1.8453699860625798 6.7859999999999995e-09 1.8247572707657775 6.787e-09 1.8345472696176197 6.788e-09 1.8478994435196154 6.789e-09 1.7744677325628664 6.79e-09 1.8500958883440177 6.791e-09 1.894673118081011 6.792e-09 1.8520620641127568 6.793e-09 1.7768004258749395 6.7939999999999995e-09 1.8479540468943392 6.795e-09 1.8225353536404858 6.796e-09 1.7865855298912887 6.7969999999999996e-09 1.871146844830438 6.798e-09 1.8312474383347332 6.799e-09 1.746583876632991 6.8e-09 1.7972718793650113 6.801e-09 1.7434225334673379 6.8019999999999995e-09 1.7224161063064007 6.803e-09 1.846610559836771 6.804e-09 1.7386936075169759 6.8049999999999996e-09 1.8848516478091129 6.806e-09 1.8214274834596111 6.807e-09 1.8387129519566614 6.808e-09 1.8237233439830416 6.809e-09 1.799791568531915 6.81e-09 1.826044276469132 6.811e-09 1.7595651019718663 6.812e-09 1.8565024900446616 6.8129999999999995e-09 1.8408376272950098 6.814e-09 1.7613441087761872 6.815e-09 1.828157376786556 6.816e-09 1.8053994110483393 6.817e-09 1.8507499795450948 6.818e-09 1.8191332690095008 6.819e-09 1.7373935299594216 6.82e-09 1.6960145546617122 6.8209999999999995e-09 1.8328674323335714 6.822e-09 1.811762259403936 6.823e-09 1.7905794594387328 6.824e-09 1.7159912645085982 6.825e-09 1.7798240811337984 6.826e-09 1.781124049395971 6.827e-09 1.7949615779723842 6.828e-09 1.8045092955422906 6.8289999999999995e-09 1.7955032806526967 6.83e-09 1.8110558478224181 6.831e-09 1.822159826608635 6.8319999999999996e-09 1.9180567983962769 6.833e-09 1.762465443199611 6.834e-09 1.7275641838431053 6.835e-09 1.7137584415843272 6.836e-09 1.8027025880187544 6.837e-09 1.7782112434005752 6.838e-09 1.7471518159788422 6.839e-09 1.8606376891396654 6.8399999999999995e-09 1.8597263169400615 6.841e-09 1.7769551510559851 6.842e-09 1.8000884653446767 6.843e-09 1.8266016054493794 6.844e-09 1.8171918941713179 6.845e-09 1.8160141159523202 6.846e-09 1.801545675204457 6.847e-09 1.8121273126524362 6.8479999999999995e-09 1.8608362739312443 6.849e-09 1.8143161757851078 6.85e-09 1.755082538714645 6.851e-09 1.7662977161806164 6.852e-09 1.8293661270045833 6.853e-09 1.7823235781057964 6.854e-09 1.8339747998740126 6.855e-09 1.8337685033028637 6.8559999999999995e-09 1.8221837320545222 6.857e-09 1.713722518038268 6.858e-09 1.8156466863593554 6.8589999999999996e-09 1.7856410714580573 6.86e-09 1.7823885390392824 6.861e-09 1.7657606890280872 6.862e-09 1.800466418594407 6.863e-09 1.758013747337024 6.8639999999999995e-09 1.784607281383986 6.865e-09 1.8386291938209276 6.866e-09 1.8171998983472715 6.8669999999999996e-09 1.8448466015184792 6.868e-09 1.7766769435481748 6.869e-09 1.8225317317433298 6.87e-09 1.7597674944319448 6.871e-09 1.7674479557489113 6.872e-09 1.7559416874979215 6.873e-09 1.734270754642664 6.874e-09 1.836930531632278 6.8749999999999995e-09 1.759599798837219 6.876e-09 1.7740272480304493 6.877e-09 1.8216047061807612 6.878e-09 1.8403206312335212 6.879e-09 1.8005149956166588 6.88e-09 1.7746594470948847 6.881e-09 1.8057855563006056 6.882e-09 1.9319492539068248 6.8829999999999995e-09 1.7817841348282053 6.884e-09 1.8315923423123317 6.885e-09 1.8027056062213573 6.886e-09 1.7915010840798418 6.887e-09 1.7058175745427369 6.888e-09 1.754541859300802 6.889e-09 1.848677467417617 6.89e-09 1.7996107786835582 6.8909999999999995e-09 1.7294793152993897 6.892e-09 1.7301217631740737 6.893e-09 1.9062083950797852 6.8939999999999996e-09 1.8238499252055687 6.895e-09 1.783306067547956 6.896e-09 1.825727500908818 6.897e-09 1.7625175177948635 6.898e-09 1.7934540903702918 6.899e-09 1.800163253725328 6.9e-09 1.8178591579239312 6.901e-09 1.8236474838142003 6.9019999999999995e-09 1.773366352929609 6.903e-09 1.8336420617728917 6.904e-09 1.7724152439464607 6.905e-09 1.8180471247178172 6.906e-09 1.818702842738627 6.907e-09 1.7901655110402555 6.908e-09 1.8047020192897583 6.909e-09 1.7693597186484264 6.9099999999999995e-09 1.8255460559580734 6.911e-09 1.8726322002356302 6.912e-09 1.7912393026636129 6.913e-09 1.8263067883352737 6.914e-09 1.8403621658975833 6.915e-09 1.8443595585472001 6.916e-09 1.8935671537748116 6.917e-09 1.7881563944987078 6.9179999999999995e-09 1.8356817384455921 6.919e-09 1.772859209481068 6.92e-09 1.8949191004802897 6.9209999999999996e-09 1.8768216643181115 6.922e-09 1.806752621669076 6.923e-09 1.813703298801809 6.924e-09 1.7727425801190762 6.925e-09 1.8933954920797778 6.9259999999999995e-09 1.7662783171338112 6.927e-09 1.7514915334812287 6.928e-09 1.7872490936113792 6.9289999999999995e-09 1.8601928251248205 6.93e-09 1.7851928652300373 6.931e-09 1.8186561029644424 6.932e-09 1.81557980290765 6.933e-09 1.7565104234227045 6.934e-09 1.7250136800184959 6.935e-09 1.8689418719832769 6.936e-09 1.7867964381435493 6.9369999999999995e-09 1.7546482199343867 6.938e-09 1.832272101321742 6.939e-09 1.8085830695926814 6.94e-09 1.6959632868551573 6.941e-09 1.696687355238965 6.942e-09 1.8163648076386543 6.943e-09 1.8128578027556854 6.944e-09 1.8240498386794552 6.9449999999999995e-09 1.8384063545556444 6.946e-09 1.791885667836203 6.947e-09 1.7468304352709934 6.9479999999999996e-09 1.8455628236319697 6.949e-09 1.896425883075482 6.95e-09 1.8456719206908698 6.951e-09 1.8163438765296318 6.952e-09 1.688119167957789 6.9529999999999995e-09 1.8293635217089055 6.954e-09 1.7175369692953448 6.955e-09 1.807332629732435 6.9559999999999996e-09 1.7668696810295585 6.957e-09 1.7317344561788848 6.958e-09 1.77844335973915 6.959e-09 1.8553305140430227 6.96e-09 1.7008912937572178 6.961e-09 1.7951746470257797 6.962e-09 1.7826284225664466 6.963e-09 1.8357897984296112 6.9639999999999995e-09 1.8807480522465099 6.965e-09 1.7821910546499604 6.966e-09 1.743495800735784 6.967e-09 1.8442118330057597 6.968e-09 1.727115239723998 6.969e-09 1.8230062771759072 6.97e-09 1.7643311249260158 6.971e-09 1.767472958654907 6.9719999999999995e-09 1.7560400770456515 6.973e-09 1.839560725332686 6.974e-09 1.8380833703177923 6.975e-09 1.7252971234148586 6.976e-09 1.848801180090743 6.977e-09 1.8061467019887147 6.978e-09 1.748083613768821 6.979e-09 1.7823365054625793 6.9799999999999995e-09 1.8069445727072144 6.981e-09 1.8001173354978666 6.982e-09 1.8312462808245762 6.9829999999999996e-09 1.8103602182222902 6.984e-09 1.7957542912652564 6.985e-09 1.8708428065459946 6.986e-09 1.8633612779156241 6.987e-09 1.7759783597341985 6.988e-09 1.7287034288460077 6.989e-09 1.788268230852207 6.99e-09 1.8069803202447325 6.9909999999999995e-09 1.7597652789299545 6.992e-09 1.7234404687027298 6.993e-09 1.7919502554580526 6.994e-09 1.8972935452178217 6.995e-09 1.8416494378665 6.996e-09 1.7869794646119794 6.997e-09 1.8189474698791217 6.998e-09 1.8649071223187688 6.9989999999999995e-09 1.9047573664763158 7e-09 1.880911370433891 7.001e-09 1.8246115794626176 7.002e-09 1.7044359915725626 7.003e-09 1.7436277545015484 7.004e-09 1.7524127510596434 7.005e-09 1.86911666217543 7.006e-09 1.8632470913060193 7.0069999999999995e-09 1.7682553643290986 7.008e-09 1.7988166760620214 7.009e-09 1.7280929280119317 7.0099999999999996e-09 1.799634981088832 7.011e-09 1.828811792480259 7.012e-09 1.8405462718697725 7.013e-09 1.7541812675679682 7.014e-09 1.7334610911502146 7.0149999999999995e-09 1.8647197760216205 7.016e-09 1.816309980786469 7.017e-09 1.7921129470210153 7.0179999999999995e-09 1.8158437912414023 7.019e-09 1.6537601791664231 7.02e-09 1.7023069324177167 7.021e-09 1.8188881249812252 7.022e-09 1.797945225601029 7.023e-09 1.7967051162236667 7.024e-09 1.8384078204375736 7.025e-09 1.7195771214829647 7.0259999999999995e-09 1.8171534294505092 7.027e-09 1.8954326872116418 7.028e-09 1.8111652970566834 7.029e-09 1.7748988123031002 7.03e-09 1.8372768273839324 7.031e-09 1.801960672094917 7.032e-09 1.8974738670158948 7.033e-09 1.84477454033289 7.0339999999999995e-09 1.7902858940215751 7.035e-09 1.7912396599795732 7.036e-09 1.7360691439247777 7.0369999999999996e-09 1.7717613695846155 7.038e-09 1.8179573959397073 7.039e-09 1.8146332706090087 7.04e-09 1.8858727658917607 7.041e-09 1.796041265659535 7.0419999999999995e-09 1.8935078648660144 7.043e-09 1.8370043386285173 7.044e-09 1.8161620734100714 7.0449999999999996e-09 1.8613954461345392 7.046e-09 1.8017829935952727 7.047e-09 1.882175233753247 7.048e-09 1.8395601677949278 7.049e-09 1.775413966996621 7.05e-09 1.829418774243068 7.051e-09 1.8246208801811146 7.052e-09 1.7859421155741797 7.0529999999999995e-09 1.846512159306838 7.054e-09 1.880343260844972 7.055e-09 1.824759803963779 7.056e-09 1.836837764093394 7.057e-09 1.8772962576198728 7.058e-09 1.8028691542306958 7.059e-09 1.8272746832082754 7.06e-09 1.7527646691127015 7.0609999999999995e-09 1.801205788277726 7.062e-09 1.889242537774825 7.063e-09 1.7974048845726556 7.064e-09 1.7547353721012309 7.065e-09 1.7349505471584667 7.066e-09 1.8485891708293285 7.067e-09 1.9025675637759358 7.068e-09 1.8582988585214602 7.0689999999999995e-09 1.8071720702878464 7.07e-09 1.777110757017752 7.071e-09 1.843221921399397 7.0719999999999996e-09 1.9067800170528946 7.073e-09 1.8581033468137356 7.074e-09 1.826433249221936 7.075e-09 1.8216215663897408 7.076e-09 1.7964128741983059 7.0769999999999994e-09 1.7927676742883083 7.078e-09 1.8387628985565816 7.079e-09 1.7501089441013737 7.0799999999999995e-09 1.8239958417486437 7.081e-09 1.702389726359053 7.082e-09 1.7991321345789097 7.083e-09 1.8673517630946392 7.084e-09 1.8337832635137632 7.085e-09 1.8036721924423436 7.086e-09 1.794839376177355 7.087e-09 1.78674784618185 7.0879999999999995e-09 1.7870380076961028 7.089e-09 1.8444895217741542 7.09e-09 1.755347319531979 7.091e-09 1.8038161577180976 7.092e-09 1.782505481616181 7.093e-09 1.7321286893866463 7.094e-09 1.805947042815898 7.095e-09 1.8439885278677535 7.0959999999999995e-09 1.8121455720036435 7.097e-09 1.7338775864344802 7.098e-09 1.7246169275945027 7.0989999999999996e-09 1.8110438012317571 7.1e-09 1.803071974593736 7.101e-09 1.7231497023489883 7.102e-09 1.8567763539699151 7.103e-09 1.8332368175712341 7.1039999999999995e-09 1.7920423474627125 7.105e-09 1.7506721038862079 7.106e-09 1.799630789776306 7.1069999999999995e-09 1.826959175750826 7.108e-09 1.857545887152493 7.109e-09 1.8313269477342018 7.11e-09 1.719070734361555 7.111e-09 1.801552281957418 7.112e-09 1.7235498641943872 7.113e-09 1.690045278499742 7.114e-09 1.9135134689749171 7.1149999999999995e-09 1.7321669991021846 7.116e-09 1.7935054684828746 7.117e-09 1.793859229766056 7.118e-09 1.879646704723535 7.119e-09 1.8121216382659695 7.12e-09 1.8097522832227333 7.121e-09 1.7836339449370129 7.122e-09 1.7999437735511647 7.1229999999999995e-09 1.815538877987991 7.124e-09 1.7473735575092018 7.125e-09 1.7920996379617282 7.126e-09 1.8576438617737967 7.127e-09 1.7665056944674584 7.128e-09 1.7734404072317351 7.129e-09 1.8230297502233765 7.13e-09 1.7636596662079915 7.1309999999999995e-09 1.7549413824393252 7.132e-09 1.799211599303245 7.133e-09 1.8586870712287034 7.1339999999999996e-09 1.7559755244469804 7.135e-09 1.7968463426571353 7.136e-09 1.7761737444704997 7.137e-09 1.9045923245966792 7.138e-09 1.8429758222862587 7.139e-09 1.7091810386176638 7.14e-09 1.7844709574578341 7.141e-09 1.7646970930002939 7.1419999999999995e-09 1.8915018076790144 7.143e-09 1.807760647730318 7.144e-09 1.808974410238496 7.145e-09 1.8390651717864337 7.146e-09 1.7251280602527077 7.147e-09 1.8026780926957076 7.148e-09 1.7480318984418783 7.149e-09 1.853299197669419 7.1499999999999995e-09 1.7700262581304052 7.151e-09 1.7985303225194627 7.152e-09 1.816644128724226 7.153e-09 1.7574797527397643 7.154e-09 1.8973027673165674 7.155e-09 1.8899218198078842 7.156e-09 1.8011056903514007 7.157e-09 1.8062734025850986 7.1579999999999995e-09 1.874135202991468 7.159e-09 1.8192809481688097 7.16e-09 1.7958073029841894 7.1609999999999996e-09 1.7421388041553172 7.162e-09 1.7631955472353515 7.163e-09 1.7945908766121499 7.164e-09 1.754024993966521 7.165e-09 1.7580865147679356 7.1659999999999994e-09 1.827963335865355 7.167e-09 1.7539042588213376 7.168e-09 1.8187145447319086 7.1689999999999995e-09 1.6910019215650436 7.17e-09 1.839039097947738 7.171e-09 1.7824998912434806 7.172e-09 1.7845791593272269 7.173e-09 1.8017895750575086 7.174e-09 1.8476850325212923 7.175e-09 1.8321851263135154 7.176e-09 1.7427843866604606 7.1769999999999995e-09 1.8395195424567696 7.178e-09 1.8465521865427623 7.179e-09 1.8915864462279468 7.18e-09 1.905937669877336 7.181e-09 1.8577792068946406 7.182e-09 1.806246696378458 7.183e-09 1.8014807718410657 7.184e-09 1.7968772977024468 7.1849999999999995e-09 1.8835449623255531 7.186e-09 1.7760395646879794 7.187e-09 1.765332683458465 7.1879999999999996e-09 1.753495092138163 7.189e-09 1.7889850187831378 7.19e-09 1.843584742109332 7.191e-09 1.8095522996551476 7.192e-09 1.811111436824813 7.1929999999999995e-09 1.7485101539585661 7.194e-09 1.9297858104582781 7.195e-09 1.7733301851890324 7.1959999999999996e-09 1.7913872756194218 7.197e-09 1.7251073934234944 7.198e-09 1.9124015055184966 7.199e-09 1.7698120903396828 7.2e-09 1.7892215764385075 7.201e-09 1.797056673035611 7.202e-09 1.7932656055085674 7.203e-09 1.7539429126029686 7.2039999999999995e-09 1.8838145158113433 7.205e-09 1.7783774681569542 7.206e-09 1.8157096677101616 7.207e-09 1.8088086821575593 7.208e-09 1.876587798024508 7.209e-09 1.7385507104220441 7.21e-09 1.832412350033287 7.211e-09 1.780706139971161 7.2119999999999995e-09 1.7815944860158877 7.213e-09 1.7813506416607081 7.214e-09 1.804397091585793 7.215e-09 1.7639300141574572 7.216e-09 1.8286535410548415 7.217e-09 1.7338685208712272 7.218e-09 1.8500677804565915 7.219e-09 1.834971668383528 7.2199999999999995e-09 1.8134722204521556 7.221e-09 1.8369673663844703 7.222e-09 1.8671985817031735 7.2229999999999996e-09 1.8449832774619273 7.224e-09 1.8241055160069535 7.225e-09 1.731313123801597 7.226e-09 1.8238937916330782 7.227e-09 1.8070658952345853 7.2279999999999994e-09 1.7947631356831537 7.229e-09 1.7070978740059 7.23e-09 1.779436449009707 7.2309999999999995e-09 1.774516830772555 7.232e-09 1.8459298922555558 7.233e-09 1.8600207052797824 7.234e-09 1.782123432864885 7.235e-09 1.7641812891909732 7.236e-09 1.8658886537123955 7.237e-09 1.8998616988829757 7.238e-09 1.8336389495823069 7.2389999999999995e-09 1.7691966812641653 7.24e-09 1.815951050850683 7.241e-09 1.7331802861948233 7.242e-09 1.802220263715723 7.243e-09 1.777364229145064 7.244e-09 1.7849544813423193 7.245e-09 1.8965228282324946 7.246e-09 1.768233013320413 7.2469999999999995e-09 1.769564032790303 7.248e-09 1.8123381343342122 7.249e-09 1.792134425890212 7.2499999999999996e-09 1.8771796565225243 7.251e-09 1.790363298840676 7.252e-09 1.802588160968555 7.253e-09 1.80755785947227 7.254e-09 1.7666765054528402 7.2549999999999995e-09 1.7213262902145603 7.256e-09 1.8378018022534899 7.257e-09 1.731101454147555 7.2579999999999995e-09 1.714134077953684 7.259e-09 1.757611900870862 7.26e-09 1.8292213459952167 7.261e-09 1.7493616784222676 7.262e-09 1.8176674008681268 7.263e-09 1.8757996887228359 7.264e-09 1.8435286068176309 7.265e-09 1.7630587200887542 7.2659999999999995e-09 1.771853647250738 7.267e-09 1.8634740767010551 7.268e-09 1.8572699773787624 7.269e-09 1.8076193050411093 7.27e-09 1.828857520356011 7.271e-09 1.8254860637351544 7.272e-09 1.826426257234025 7.273e-09 1.7665552825454767 7.2739999999999995e-09 1.804607841186233 7.275e-09 1.8169328338191655 7.276e-09 1.7274194692637617 7.2769999999999996e-09 1.8703637244220832 7.278e-09 1.7639856272993923 7.279e-09 1.8457198998510198 7.28e-09 1.7915760192803785 7.281e-09 1.8091523700796792 7.2819999999999995e-09 1.7825924900868133 7.283e-09 1.7765356903459617 7.284e-09 1.839364917266293 7.2849999999999996e-09 1.842467317089751 7.286e-09 1.7133535096802064 7.287e-09 1.880021474623015 7.288e-09 1.768901528080318 7.289e-09 1.8396894689194259 7.29e-09 1.829846036906399 7.291e-09 1.8462385695037788 7.292e-09 1.8232958087191729 7.2929999999999995e-09 1.8664189980918757 7.294e-09 1.7932187650459976 7.295e-09 1.896411465519972 7.296e-09 1.7445449491546594 7.297e-09 1.816399992195796 7.298e-09 1.8264764074852982 7.299e-09 1.7991781563944593 7.3e-09 1.776855228622538 7.3009999999999995e-09 1.7696652334752667 7.302e-09 1.819728848829338 7.303e-09 1.8946814082985606 7.304e-09 1.9462169626389068 7.305e-09 1.7792374146869132 7.306e-09 1.8081292616369717 7.307e-09 1.8176685143638402 7.308e-09 1.739389694820677 7.3089999999999995e-09 1.7661214449281049 7.31e-09 1.8315083319743057 7.311e-09 1.7690581715391878 7.3119999999999996e-09 1.714270612948033 7.313e-09 1.740859443895641 7.314e-09 1.7399311741201056 7.315e-09 1.8173744580669087 7.316e-09 1.8847126798232297 7.3169999999999994e-09 1.7593109649437237 7.318e-09 1.7254591689797127 7.319e-09 1.8691956393139164 7.3199999999999995e-09 1.8202898867987098 7.321e-09 1.7522694393609668 7.322e-09 1.9022463479601823 7.323e-09 1.8119387787848127 7.324e-09 1.774178868351197 7.325e-09 1.680402888183156 7.326e-09 1.7281019788297391 7.327e-09 1.7737165268892763 7.3279999999999995e-09 1.7752110292464034 7.329e-09 1.8396872923115852 7.33e-09 1.8497878704089912 7.331e-09 1.7776882215171805 7.332e-09 1.7248905985330127 7.333e-09 1.7915574383501114 7.334e-09 1.70278618446798 7.335e-09 1.8871768969600955 7.3359999999999995e-09 1.7874908232860796 7.337e-09 1.8347218580267501 7.338e-09 1.8019550646412859 7.3389999999999996e-09 1.7627796799251985 7.34e-09 1.6956975859830326 7.341e-09 1.7193162455074211 7.342e-09 1.7872880968727505 7.343e-09 1.7421614109610697 7.3439999999999995e-09 1.806149274033464 7.345e-09 1.8342894115509762 7.346e-09 1.7300096977441497 7.3469999999999995e-09 1.755119568174147 7.348e-09 1.815774603048333 7.349e-09 1.79261026243444 7.35e-09 1.766949767967831 7.351e-09 1.8232215633421174 7.352e-09 1.6976719415651247 7.353e-09 1.7519762152056475 7.354e-09 1.7106308248289723 7.3549999999999995e-09 1.852078221563232 7.356e-09 1.8083604569258673 7.357e-09 1.8016093479203215 7.358e-09 1.8127754801380311 7.359e-09 1.8346935631577537 7.36e-09 1.8893141142044854 7.361e-09 1.813960548664534 7.362e-09 1.8092551975903284 7.3629999999999995e-09 1.8440459152170685 7.364e-09 1.7641060182563377 7.365e-09 1.7768259447093502 7.3659999999999996e-09 1.7239624959536388 7.367e-09 1.7838773104636747 7.368e-09 1.8397919119117212 7.369e-09 1.757918983238431 7.37e-09 1.7009823162681799 7.3709999999999995e-09 1.9491814783597343 7.372e-09 1.738737201168791 7.373e-09 1.8066646884576851 7.3739999999999996e-09 1.8157057095013647 7.375e-09 1.9174166289121721 7.376e-09 1.7941741438864283 7.377e-09 1.8151740595341213 7.378e-09 1.7693022652863863 7.379e-09 1.7901730455059657 7.38e-09 1.802110817655073 7.381e-09 1.8359658929231248 7.3819999999999995e-09 1.844562697635894 7.383e-09 1.792065549644502 7.384e-09 1.784684949290568 7.385e-09 1.8259472865142046 7.386e-09 1.779605845029761 7.387e-09 1.799949048781265 7.388e-09 1.8127944649780274 7.389e-09 1.7576531597176859 7.3899999999999995e-09 1.7297801479367132 7.391e-09 1.7290158706264271 7.392e-09 1.814219268030438 7.393e-09 1.8438503395776493 7.394e-09 1.8704035955510085 7.395e-09 1.7558458698203343 7.396e-09 1.8361426961762266 7.397e-09 1.7664127530931824 7.3979999999999995e-09 1.8945981690117182 7.399e-09 1.8083786627108562 7.4e-09 1.7496420386020437 7.4009999999999996e-09 1.8241507023068506 7.402e-09 1.783211941825605 7.403e-09 1.8444570140477168 7.404e-09 1.83049140044489 7.405e-09 1.906402854688558 7.4059999999999994e-09 1.7723581656012812 7.407e-09 1.7463725586497223 7.408e-09 1.8302288747729727 7.4089999999999995e-09 1.7900704629717277 7.41e-09 1.7938362057201074 7.411e-09 1.819107614793546 7.412e-09 1.8130256255625905 7.413e-09 1.8213276236053788 7.414e-09 1.6847278158091665 7.415e-09 1.7866360742428538 7.416e-09 1.812451051135377 7.4169999999999995e-09 1.7616795481185152 7.418e-09 1.8281651503662752 7.419e-09 1.8404180983619165 7.42e-09 1.765642001256942 7.421e-09 1.7558741959138082 7.422e-09 1.8358398098837385 7.423e-09 1.811295674236607 7.424e-09 1.7956913087350248 7.4249999999999995e-09 1.7500253286313328 7.426e-09 1.838141403040565 7.427e-09 1.7509303985634366 7.4279999999999996e-09 1.6809910070042877 7.429e-09 1.8099138204944327 7.43e-09 1.7151093244781614 7.431e-09 1.8234940653748757 7.432e-09 1.791068014319864 7.4329999999999995e-09 1.829237525607154 7.434e-09 1.820796976846225 7.435e-09 1.8145019551366315 7.4359999999999996e-09 1.802154740501383 7.437e-09 1.8385688704076353 7.438e-09 1.8120132867399341 7.439e-09 1.7687564425358706 7.44e-09 1.8602104037638354 7.441e-09 1.8335526289258484 7.442e-09 1.7510443888973855 7.443e-09 1.8481402589557923 7.4439999999999995e-09 1.8219981922261508 7.445e-09 1.7348722948296103 7.446e-09 1.7593628772484793 7.447e-09 1.7999691316648223 7.448e-09 1.812481254815476 7.449e-09 1.830980625434848 7.45e-09 1.8733601952217211 7.451e-09 1.7003152788290556 7.452e-09 1.8610403599611995 7.453e-09 1.8359945353581357 7.454e-09 1.7830507550775796 7.455e-09 1.831411934203659 7.455999999999999e-09 1.8623010451788635 7.457e-09 1.8238337710708554 7.458e-09 1.8034719699687314 7.458999999999999e-09 1.7985796810821455 7.46e-09 1.7421992285396675 7.461e-09 1.8967327283725604 7.462e-09 1.8557895847655588 7.463e-09 1.8265854276346785 7.464e-09 1.8326079555667967 7.465e-09 1.8190184545665025 7.466e-09 1.7385086793744902 7.467e-09 1.8623081673182882 7.468e-09 1.795534302699932 7.469e-09 1.800476185520678 7.47e-09 1.73343072243091 7.471e-09 1.8061813866122545 7.472e-09 1.8163497081432984 7.473e-09 1.7298163590229338 7.474e-09 1.816463280710569 7.474999999999999e-09 1.867480748569857 7.476e-09 1.8778642087406887 7.477e-09 1.7425752896737465 7.478e-09 1.7337252966030121 7.479e-09 1.7671897782147152 7.48e-09 1.790180513255834 7.481e-09 1.7154869215536392 7.482e-09 1.7473209516419328 7.483e-09 1.795342615942716 7.484e-09 1.8437265410785946 7.485e-09 1.8265499709277007 7.486e-09 1.7472404089784215 7.487e-09 1.8284331268510252 7.488e-09 1.8312794763672229 7.489e-09 1.8175487442206415 7.49e-09 1.829612638086651 7.490999999999999e-09 1.8254739045719737 7.492e-09 1.761163735212581 7.493e-09 1.8804855660205284 7.493999999999999e-09 1.8153588163276047 7.495e-09 1.8274105450203604 7.496e-09 1.7656391702753438 7.497e-09 1.81996434907379 7.498e-09 1.7589826277072604 7.499e-09 1.7848315265301822 7.5e-09 1.795729017005273 7.501e-09 1.7605367342300735 7.502e-09 1.7565231659144722 7.503e-09 1.7879565830726833 7.504e-09 1.8191351300461613 7.505e-09 1.8592671744026734 7.506e-09 1.755919366146284 7.507e-09 1.8087296176692285 7.508e-09 1.7623535305531028 7.509e-09 1.7554602171601927 7.509999999999999e-09 1.695995333670105 7.511e-09 1.9054601444253096 7.512e-09 1.8399521807360804 7.513e-09 1.727854075083149 7.514e-09 1.8242023710250344 7.515e-09 1.7328000726389754 7.516e-09 1.921640744840237 7.517e-09 1.8204167434073364 7.518e-09 1.88297272554533 7.519e-09 1.7261587482537335 7.52e-09 1.7884602053101666 7.521e-09 1.80756130255344 7.522e-09 1.795128379994801 7.523e-09 1.801191775264786 7.524e-09 1.8360798193288164 7.525e-09 1.751484316959374 7.525999999999999e-09 1.874751142646816 7.527e-09 1.8237349790578343 7.528e-09 1.8731659871297044 7.528999999999999e-09 1.8081112902810554 7.53e-09 1.7853356185315659 7.531e-09 1.9276972674696402 7.532e-09 1.7594068747122333 7.533e-09 1.8035312118643319 7.534e-09 1.753661154135134 7.535e-09 1.8535481569782224 7.536e-09 1.7213465961216161 7.537e-09 1.841003893900332 7.538e-09 1.7591588916089433 7.539e-09 1.7425270979281804 7.54e-09 1.813978511383597 7.541e-09 1.8300382174869552 7.542e-09 1.8287240462458565 7.543e-09 1.872438811370869 7.544e-09 1.862398806096272 7.544999999999999e-09 1.802807067606119 7.546e-09 1.8220852211153749 7.547e-09 1.8316880561832327 7.547999999999999e-09 1.793291571578375 7.549e-09 1.811302819756189 7.55e-09 1.8521099523981963 7.551e-09 1.8509649873254326 7.552e-09 1.796058346191295 7.553e-09 1.9091005540366868 7.554e-09 1.8336315258525648 7.555e-09 1.8142793152290293 7.556e-09 1.7750563290879513 7.557e-09 1.7586662862827969 7.558e-09 1.9019653866280923 7.559e-09 1.7581613867734551 7.56e-09 1.7976879760278608 7.561e-09 1.7429031842838985 7.562e-09 1.7345998898321628 7.563e-09 1.8219589083148875 7.563999999999999e-09 1.8492995071154263 7.565e-09 1.8184822388127928 7.566e-09 1.7844982881558829 7.567e-09 1.893215257104146 7.568e-09 1.7399174044515773 7.569e-09 1.7869107940376348 7.57e-09 1.7759643262547502 7.571e-09 1.8114072495359452 7.572e-09 1.8179860681953601 7.573e-09 1.7440931406208946 7.574e-09 1.6910380808174277 7.575e-09 1.8490314676744437 7.576e-09 1.8399688601680069 7.577e-09 1.82463282333309 7.578e-09 1.8787894530842608 7.579e-09 1.7634311992444727 7.579999999999999e-09 1.836815386387035 7.581e-09 1.7825635813056089 7.582e-09 1.7764680671768047 7.582999999999999e-09 1.8200313010496656 7.584e-09 1.7947656754975694 7.585e-09 1.7647477913949552 7.586e-09 1.7540487764627488 7.587e-09 1.8215789772014093 7.588e-09 1.7538562682586603 7.589e-09 1.742242777596183 7.59e-09 1.8013705208702933 7.591e-09 1.814261606276871 7.592e-09 1.6837319159733264 7.593e-09 1.7288510372659434 7.594e-09 1.803518144643821 7.595e-09 1.76449350598248 7.596e-09 1.839604575803766 7.597e-09 1.7272799612464982 7.598e-09 1.8042866301106535 7.598999999999999e-09 1.650520233075051 7.6e-09 1.8217001685958523 7.601e-09 1.7848787991661952 7.602e-09 1.7770354511787667 7.603e-09 1.908436776926453 7.604e-09 1.7500202224332468 7.605e-09 1.8694149046798303 7.606e-09 1.731898921404304 7.607e-09 1.749365479446021 7.608e-09 1.7143492321497684 7.609e-09 1.8068444240421755 7.61e-09 1.860959361532387 7.611e-09 1.834619281223419 7.612e-09 1.7800037988636963 7.613e-09 1.7309496956687191 7.614e-09 1.763573784307089 7.614999999999999e-09 1.8049253098906066 7.616e-09 1.7429654960110896 7.617e-09 1.7448049406186583 7.617999999999999e-09 1.791589961029908 7.619e-09 1.7984395548605965 7.62e-09 1.849689106459371 7.621e-09 1.8250510203945545 7.622e-09 1.85039151187437 7.623e-09 1.7841058631408322 7.624e-09 1.6970652053397977 7.625e-09 1.8286227902064893 7.626e-09 1.7873440793415059 7.627e-09 1.7843667124992793 7.628e-09 1.8497929825533013 7.629e-09 1.737352405736411 7.63e-09 1.7785341226203102 7.631e-09 1.7989521180132604 7.632e-09 1.8076026578020994 7.633e-09 1.7735430450251402 7.633999999999999e-09 1.7695686446794856 7.635e-09 1.8649356307602798 7.636e-09 1.834197430550742 7.636999999999999e-09 1.7411412028843736 7.638e-09 1.8408539455409512 7.639e-09 1.817248458857715 7.64e-09 1.780813078637577 7.641e-09 1.7808593026446706 7.642e-09 1.866424345205869 7.643e-09 1.7663684408354285 7.644e-09 1.7861217155663849 7.645e-09 1.727586030283444 7.646e-09 1.8635351092470567 7.647e-09 1.8204286970735686 7.648e-09 1.847617965957422 7.649e-09 1.728264141095119 7.65e-09 1.7817712709585714 7.651e-09 1.7996004085995443 7.652e-09 1.7408923965699827 7.652999999999999e-09 1.7854826869511127 7.654e-09 1.8676667699931038 7.655e-09 1.8412949010901556 7.656e-09 1.801380144945576 7.657e-09 1.857881741214122 7.658e-09 1.8690142155513148 7.659e-09 1.8264109662086034 7.66e-09 1.8097384742380997 7.661e-09 1.8884925818610219 7.662e-09 1.773760563644661 7.663e-09 1.724878977579578 7.664e-09 1.7997155856578506 7.665e-09 1.7841137408462813 7.666e-09 1.7711172775806938 7.667e-09 1.8191413885245482 7.668e-09 1.873519428390104 7.668999999999999e-09 1.8369029935758039 7.67e-09 1.8586238252980085 7.671e-09 1.8430619338173944 7.671999999999999e-09 1.759919042439172 7.673e-09 1.8042652470476275 7.674e-09 1.770902791900087 7.675e-09 1.7615402577363157 7.676e-09 1.8508129900437393 7.677e-09 1.7897031109161268 7.678e-09 1.7934277401387693 7.679e-09 1.9337867082996565 7.68e-09 1.7309657299070422 7.681e-09 1.856048300972207 7.682e-09 1.8472710237400283 7.683e-09 1.7632527002767808 7.684e-09 1.9125921347122994 7.685e-09 1.8099225981675355 7.686e-09 1.8117504176131893 7.687e-09 1.7723159539368032 7.687999999999999e-09 1.761363791831793 7.689e-09 1.760172376037192 7.69e-09 1.7699871682832493 7.691e-09 1.88775743256442 7.692e-09 1.8211929496996757 7.693e-09 1.8232562474994818 7.694e-09 1.861861666594211 7.695e-09 1.7911594640466448 7.696e-09 1.7832835847029662 7.697e-09 1.8135032600775234 7.698e-09 1.7657563012860433 7.699e-09 1.8449583830033423 7.7e-09 1.9511102668054354 7.701e-09 1.7926611471352347 7.702e-09 1.753675996638061 7.703e-09 1.7440155976822516 7.703999999999999e-09 1.7923449204682371 7.705e-09 1.7910103885083517 7.706e-09 1.7778178301586998 7.706999999999999e-09 1.7375242108341062 7.708e-09 1.817148550963095 7.709e-09 1.809566140013775 7.71e-09 1.7957140558237428 7.711e-09 1.7915112060404668 7.712e-09 1.7873135745349868 7.713e-09 1.797745650235507 7.714e-09 1.8403653136869151 7.715e-09 1.8311677279593481 7.716e-09 1.6942833714742325 7.717e-09 1.8553123623273644 7.718e-09 1.768901971818714 7.719e-09 1.808493377987871 7.72e-09 1.80170428321992 7.721e-09 1.768448623841926 7.722e-09 1.6779372946277127 7.722999999999999e-09 1.7882737193825058 7.724e-09 1.8149082761378048 7.725e-09 1.7920932710470143 7.725999999999999e-09 1.773419270787524 7.727e-09 1.9089348990093382 7.728e-09 1.7874321906308566 7.729e-09 1.7031808904267691 7.73e-09 1.7999335241627272 7.731e-09 1.7891125767865328 7.732e-09 1.7008020558393102 7.733e-09 1.7333297832894883 7.734e-09 1.8503647736664597 7.735e-09 1.8404394614996993 7.736e-09 1.9066234661273882 7.737e-09 1.8476890168309612 7.738e-09 1.7308440136350203 7.738999999999999e-09 1.8236654369037897 7.74e-09 1.7466821677914746 7.741e-09 1.8188079833825141 7.741999999999999e-09 1.7653737620948244 7.743e-09 1.751857550534386 7.744e-09 1.779050900183468 7.745e-09 1.8203050970665324 7.746e-09 1.8077583040457987 7.747e-09 1.7433890105736547 7.748e-09 1.822464469628285 7.749e-09 1.8598378444057246 7.75e-09 1.772974126342533 7.751e-09 1.8613186839173397 7.752e-09 1.7638218941621668 7.753e-09 1.80419257586195 7.754e-09 1.730058915487154 7.755e-09 1.7214732092661942 7.756e-09 1.7719509872290877 7.757e-09 1.7770607401081715 7.757999999999999e-09 1.784990873281522 7.759e-09 1.77647309969713 7.76e-09 1.8212789507848282 7.760999999999999e-09 1.8396441435489561 7.762e-09 1.8836938925088258 7.763e-09 1.7542175559093287 7.764e-09 1.7879156797710902 7.765e-09 1.786429242759973 7.766e-09 1.8204508288454306 7.767e-09 1.768253382535846 7.768e-09 1.7991824296345171 7.769e-09 1.7980006508122128 7.77e-09 1.8647979464298776 7.771e-09 1.8088635348167068 7.772e-09 1.7311104697087105 7.773e-09 1.8282372538035876 7.774e-09 1.818612259078853 7.775e-09 1.7883521206399675 7.776e-09 1.7952805476325886 7.776999999999999e-09 1.8801399586669076 7.778e-09 1.7932572842771128 7.779e-09 1.7565256275833907 7.78e-09 1.784998015346147 7.781e-09 1.7543875373597881 7.782e-09 1.8086503241626128 7.783e-09 1.759335575340566 7.784e-09 1.758106631055548 7.785e-09 1.794436840004581 7.786e-09 1.7933052108468222 7.787e-09 1.8020277409485657 7.788e-09 1.7956145014657323 7.789e-09 1.8110645190803398 7.79e-09 1.762661306041783 7.791e-09 1.8472649154771588 7.792e-09 1.7748683227821478 7.792999999999999e-09 1.7685093508096852 7.794e-09 1.7428645828019231 7.795e-09 1.7601108363269322 7.795999999999999e-09 1.7723656029175938 7.797e-09 1.8542384994227983 7.798e-09 1.802218937594359 7.799e-09 1.8403462433642073 7.8e-09 1.8063854606539622 7.801e-09 1.8607137803000944 7.802e-09 1.7877127597391436 7.803e-09 1.8809167841778596 7.804e-09 1.760411851881249 7.805e-09 1.806972504353936 7.806e-09 1.8196838422217636 7.807e-09 1.8536693906155477 7.808e-09 1.716832769466838 7.809e-09 1.7453144379256698 7.81e-09 1.8398421641303253 7.811e-09 1.7948647048631543 7.811999999999999e-09 1.7676096298930646 7.813e-09 1.8557698757820786 7.814e-09 1.845318210094298 7.814999999999999e-09 1.819891958205315 7.816e-09 1.8330261119102345 7.817e-09 1.9177441085166138 7.818e-09 1.8512604962530796 7.819e-09 1.7613813224129986 7.82e-09 1.7715482359477321 7.821e-09 1.9013000577781045 7.822e-09 1.7758880737115161 7.823e-09 1.7946830047020073 7.824e-09 1.7740575917859998 7.825e-09 1.7629660975214092 7.826e-09 1.8036477233396397 7.827e-09 1.8898895125104045 7.827999999999999e-09 1.7721370834317758 7.829e-09 1.8145781012116793 7.83e-09 1.842195270949715 7.830999999999999e-09 1.7736042826453648 7.832e-09 1.7430172194611322 7.833e-09 1.8237801855385694 7.834e-09 1.7458607319030404 7.835e-09 1.7761367385543683 7.836e-09 1.6338982068144952 7.837e-09 1.774899965905029 7.838e-09 1.8363888342835621 7.839e-09 1.797223933784632 7.84e-09 1.7785109504638283 7.841e-09 1.8508313566660584 7.842e-09 1.7459690433469046 7.843e-09 1.845628836737712 7.844e-09 1.7905938077782615 7.845e-09 1.7818418812954508 7.846e-09 1.804326370945349 7.846999999999999e-09 1.832237412865356 7.848e-09 1.8189853915996237 7.849e-09 1.883199656251732 7.849999999999999e-09 1.7894745325826142 7.851e-09 1.8706787617702925 7.852e-09 1.790103808224093 7.853e-09 1.8091942481660301 7.854e-09 1.7768803924143193 7.855e-09 1.8631913436978713 7.856e-09 1.744911837764903 7.857e-09 1.8321966963264227 7.858e-09 1.6938109270442712 7.859e-09 1.821047339826913 7.86e-09 1.7570630109713836 7.861e-09 1.8348454053670724 7.862e-09 1.7946568265812366 7.863e-09 1.809201286494231 7.864e-09 1.8606745176120527 7.865e-09 1.8246843527143166 7.865999999999999e-09 1.76972217600354 7.867e-09 1.8110215363871225 7.868e-09 1.849849922242703 7.869e-09 1.6954510024202 7.87e-09 1.7301729639775152 7.871e-09 1.7925094716603485 7.872e-09 1.8464396879646974 7.873e-09 1.723855212763242 7.874e-09 1.8107230692712082 7.875e-09 1.7183949237726606 7.876e-09 1.7203917857011648 7.877e-09 1.769514418399699 7.878e-09 1.6552751293431232 7.879e-09 1.691945832956916 7.88e-09 1.8273332334120294 7.881e-09 1.7767552886483169 7.881999999999999e-09 1.7979427241608954 7.883e-09 1.7701233239130323 7.884e-09 1.7161473952649646 7.884999999999999e-09 1.8012842575823156 7.886e-09 1.7904003834235542 7.887e-09 1.756089243455243 7.888e-09 1.7744438332274513 7.889e-09 1.6919346924190832 7.89e-09 1.7562431604382434 7.891e-09 1.7439268554300345 7.892e-09 1.9032716299996053 7.893e-09 1.841461188744818 7.894e-09 1.7324652254557398 7.895e-09 1.891783940973871 7.896e-09 1.8488588191586994 7.897e-09 1.807682873077094 7.898e-09 1.7125831019260211 7.899e-09 1.7247931290062182 7.9e-09 1.7621049720264308 7.900999999999999e-09 1.7466895636029451 7.902e-09 1.8348665698689888 7.903e-09 1.8352832034648585 7.904e-09 1.7888896583122726 7.905e-09 1.858587063857991 7.906e-09 1.8759218515936378 7.907e-09 1.8273766038928883 7.908e-09 1.848352093826026 7.909e-09 1.8302437571693044 7.91e-09 1.8536698194375887 7.911e-09 1.7572582245015849 7.912e-09 1.7759204414212382 7.913e-09 1.7049239968930354 7.914e-09 1.808787260520516 7.915e-09 1.787599806552955 7.916e-09 1.7029375475263477 7.916999999999999e-09 1.7543379804328691 7.918e-09 1.846145950143851 7.919e-09 1.8221495652440018 7.919999999999999e-09 1.7985003942139794 7.921e-09 1.7812099405881785 7.922e-09 1.7965922526792533 7.923e-09 1.7627723619895888 7.924e-09 1.7140046085483402 7.925e-09 1.823285173979401 7.926e-09 1.8100281515704613 7.927e-09 1.7737398745647226 7.928e-09 1.758243073574788 7.929e-09 1.8350571460399965 7.93e-09 1.8293061436613332 7.931e-09 1.8151701237237972 7.932e-09 1.7597379323104283 7.933e-09 1.8193950816944047 7.934e-09 1.8379296144212298 7.935e-09 1.78073675836428 7.935999999999999e-09 1.7779934665239545 7.937e-09 1.8076330066316093 7.938e-09 1.835594871059296 7.938999999999999e-09 1.8141848373550284 7.94e-09 1.7578571591282428 7.941e-09 1.774101060575272 7.942e-09 1.7960904904175248 7.943e-09 1.8330198427256685 7.944e-09 1.7899303836014193 7.945e-09 1.788045424907063 7.946e-09 1.8791302009398438 7.947e-09 1.7627519312745772 7.948e-09 1.7632931552814974 7.949e-09 1.828155280849374 7.95e-09 1.8410477804828698 7.951e-09 1.928240828367068 7.952e-09 1.6437136548822937 7.953e-09 1.8310110427282649 7.954e-09 1.8783134541193391 7.954999999999999e-09 1.8788008033168382 7.956e-09 1.838915313262065 7.957e-09 1.8856713013252873 7.958e-09 1.7546357941859116 7.959e-09 1.7949308823504593 7.96e-09 1.860700989879145 7.961e-09 1.8259902714765768 7.962e-09 1.8401482431020553 7.963e-09 1.8971639446268311 7.964e-09 1.7919931495157317 7.965e-09 1.8178463769924058 7.966e-09 1.8605017942517863 7.967e-09 1.931253397567514 7.968e-09 1.8677986155193902 7.969e-09 1.8144681002808438 7.97e-09 1.8389328044434852 7.970999999999999e-09 1.803911162918552 7.972e-09 1.8532545879837399 7.973e-09 1.8230624450720696 7.973999999999999e-09 1.8443763133297348 7.975e-09 1.873744356787674 7.976e-09 1.7650562317471123 7.977e-09 1.866691311709665 7.978e-09 1.7195512959797266 7.979e-09 1.820504401896216 7.98e-09 1.8397907048847344 7.981e-09 1.806788977045568 7.982e-09 1.741639746515015 7.983e-09 1.8089024222768277 7.984e-09 1.781611114863281 7.985e-09 1.7378761235596836 7.986e-09 1.6579636520839502 7.987e-09 1.6725009950826444 7.988e-09 1.8208533625302876 7.989e-09 1.793634990065249 7.989999999999999e-09 1.7797760665708613 7.991e-09 1.8314323961762127 7.992e-09 1.8578684507416885 7.993e-09 1.7403326777081016 7.994e-09 1.7858350935178984 7.995e-09 1.6534065870758987 7.996e-09 1.83762805097618 7.997e-09 1.7937879531365963 7.998e-09 1.8604662588580416 7.999e-09 1.802496727760308 8e-09 1.7142256197611263 8.001e-09 1.811974590095675 8.002e-09 1.7607066077526672 8.003e-09 1.8322605011015616 8.004e-09 1.830460990832906 8.005e-09 1.7638392980771487 8.005999999999999e-09 1.7298063876406058 8.007e-09 1.8425883967919943 8.008e-09 1.8163446548074622 8.008999999999999e-09 1.8021857404787722 8.01e-09 1.8108682172002952 8.011e-09 1.7743180732404567 8.012e-09 1.7427252078408666 8.013e-09 1.9145219666686542 8.014e-09 1.791963662483676 8.015e-09 1.869043956242265 8.016e-09 1.7957383656885149 8.017e-09 1.7641547881586843 8.018e-09 1.7557860505933716 8.019e-09 1.852035752639556 8.02e-09 1.7847487574381353 8.021e-09 1.7781294814738817 8.022e-09 1.7924525370584345 8.023e-09 1.855781915988221 8.024e-09 1.6860064313131238 8.024999999999999e-09 1.7925815438160602 8.026e-09 1.8155615589573357 8.027e-09 1.7577786794145196 8.027999999999999e-09 1.7152285012565658 8.029e-09 1.839906631932876 8.03e-09 1.790661437537706 8.031e-09 1.7658531657834216 8.032e-09 1.7360905871721521 8.033e-09 1.7857354677696253 8.034e-09 1.7012889920252166 8.035e-09 1.7761165760313702 8.036e-09 1.7732800979595165 8.037e-09 1.934998735694208 8.038e-09 1.8624238602092982 8.039e-09 1.901611124452374 8.04e-09 1.8275463474114697 8.040999999999999e-09 1.8911578045740394 8.042e-09 1.7882608747553463 8.043e-09 1.7781251235203475 8.043999999999999e-09 1.7845381009088328 8.045e-09 1.7522331525857557 8.046e-09 1.7909062796837092 8.047e-09 1.8094784696336124 8.048e-09 1.7180141252549452 8.049e-09 1.8243017026570216 8.05e-09 1.78654289672021 8.051e-09 1.8510043266034917 8.052e-09 1.7882680399337785 8.053e-09 1.8647409840011955 8.054e-09 1.8191271869667596 8.055e-09 1.8018482768592154 8.056e-09 1.9494906342031777 8.057e-09 1.7948744053387202 8.058e-09 1.7211864600131481 8.059e-09 1.7529413736361672 8.059999999999999e-09 1.7972809565837142 8.061e-09 1.800688123266939 8.062e-09 1.7802186327784923 8.062999999999999e-09 1.8332254167800284 8.064e-09 1.850164766855076 8.065e-09 1.8439329620336753 8.066e-09 1.8006159036179614 8.067e-09 1.7643186158911808 8.068e-09 1.7815147953570774 8.069e-09 1.765695942048241 8.07e-09 1.8308706241787034 8.071e-09 1.7665335172307208 8.072e-09 1.7122404336301338 8.073e-09 1.8478966855959982 8.074e-09 1.720722757386393 8.075e-09 1.8020423201585911 8.076e-09 1.7661627791648014 8.077e-09 1.8106402918675117 8.078e-09 1.8310210863825356 8.078999999999999e-09 1.814290088493494 8.08e-09 1.767874446665708 8.081e-09 1.7930259085725773 8.082e-09 1.8170618327883248 8.083e-09 1.8294250894901245 8.084e-09 1.884150522222608 8.085e-09 1.83503524601864 8.086e-09 1.7452954666247784 8.087e-09 1.7864643177052986 8.088e-09 1.695115572233885 8.089e-09 1.7675504277519911 8.09e-09 1.815076414059441 8.091e-09 1.8785319939916387 8.092e-09 1.8164739628344466 8.093e-09 1.7790934010426356 8.094e-09 1.7774314526409947 8.094999999999999e-09 1.8366111837520245 8.096e-09 1.8499201471438533 8.097e-09 1.689660774858201 8.097999999999999e-09 1.801776348123856 8.099e-09 1.7613407060229584 8.1e-09 1.7817252609330043 8.101e-09 1.790390007872107 8.102e-09 1.833059109170925 8.103e-09 1.8182401372178492 8.104e-09 1.7856950365005475 8.105e-09 1.7949764184414676 8.106e-09 1.805105117914483 8.107e-09 1.688516621620395 8.108e-09 1.7195455926977412 8.109e-09 1.8282262657079864 8.11e-09 1.77928179203214 8.111e-09 1.7644958201154899 8.112e-09 1.8079972182418547 8.113e-09 1.760172075975644 8.113999999999999e-09 1.8256124309297892 8.115e-09 1.7440424582227254 8.116e-09 1.8811344217859742 8.116999999999999e-09 1.7621730027133977 8.118e-09 1.6925827957244861 8.119e-09 1.7772883736636371 8.12e-09 1.7909055806363832 8.121e-09 1.7869871469318885 8.122e-09 1.7414024805441215 8.123e-09 1.7451874554213567 8.124e-09 1.807762493696635 8.125e-09 1.9044787347248686 8.126e-09 1.8644888345246442 8.127e-09 1.8716544840987936 8.128e-09 1.8347734463859264 8.129e-09 1.8136992278077357 8.129999999999999e-09 1.7913492317735813 8.131e-09 1.9289314750641195 8.132e-09 1.8075502066084608 8.132999999999999e-09 1.8165819497331004 8.134e-09 1.7240536839703935 8.135e-09 1.801364125367686 8.136e-09 1.7621623416228336 8.137e-09 1.6742786493992285 8.138e-09 1.8238941667937123 8.139e-09 1.737450170587807 8.14e-09 1.857039757343263 8.141e-09 1.8466581645232305 8.142e-09 1.6900259639999962 8.143e-09 1.8673150089997723 8.144e-09 1.773936448036497 8.145e-09 1.763035330393291 8.146e-09 1.7484391364503034 8.147e-09 1.8267752602846201 8.148e-09 1.6926229478384183 8.148999999999999e-09 1.7665935918422033 8.15e-09 1.818527801666245 8.151e-09 1.7249549666660289 8.151999999999999e-09 1.802688809826555 8.153e-09 1.772720282577931 8.154e-09 1.7425211183706295 8.155e-09 1.7763604819010421 8.156e-09 1.7940772100228317 8.157e-09 1.7409803736473266 8.158e-09 1.784354604170304 8.159e-09 1.7980865255906135 8.16e-09 1.729441930846995 8.161e-09 1.7682447542243285 8.162e-09 1.7474449935962373 8.163e-09 1.8158789554754273 8.164e-09 1.8111862801090854 8.165e-09 1.7776329362620127 8.166e-09 1.903923646232545 8.167e-09 1.8204948108255714 8.167999999999999e-09 1.800028248645639 8.169e-09 1.7798543827293174 8.17e-09 1.7787760956089094 8.171e-09 1.7804546382738895 8.172e-09 1.9024532047671505 8.173e-09 1.8313110978538725 8.174e-09 1.819485367629147 8.175e-09 1.7427787656195042 8.176e-09 1.8588534580279736 8.177e-09 1.8392240097669499 8.178e-09 1.9110095610222142 8.179e-09 1.8167160373360778 8.18e-09 1.815167833087069 8.181e-09 1.7700768062145296 8.182e-09 1.8133545989938806 8.183e-09 1.7681508417460163 8.183999999999999e-09 1.7503171431219906 8.185e-09 1.8124725967143045 8.186e-09 1.8088034464329195 8.186999999999999e-09 1.8081526588966907 8.188e-09 1.7723311611416095 8.189e-09 1.754585457902432 8.19e-09 1.8326955733593282 8.191e-09 1.8466258008945178 8.192e-09 1.8572303095958604 8.193e-09 1.7887182574559546 8.194e-09 1.7829385317619857 8.195e-09 1.745348652149233 8.196e-09 1.8038759079812885 8.197e-09 1.879552058561205 8.198e-09 1.9001419612503234 8.199e-09 1.8491324375326759 8.2e-09 1.8890607973853606 8.201e-09 1.81758361187943 8.202e-09 1.7563969029663247 8.202999999999999e-09 1.759987858746441 8.204e-09 1.8394841819130416 8.205e-09 1.8010578694220325 8.205999999999999e-09 1.8517483755829423 8.207e-09 1.8280874080978158 8.208e-09 1.6788814974528246 8.209e-09 1.835433746982008 8.21e-09 1.8142081276117041 8.211e-09 1.8323384647500762 8.212e-09 1.744558188836076 8.213e-09 1.7221658754239582 8.214e-09 1.8538604897439896 8.215e-09 1.8355573475070688 8.216e-09 1.792781667376698 8.217e-09 1.7893964117763046 8.218e-09 1.7937809907065165 8.218999999999999e-09 1.858620512962886 8.22e-09 1.802611178910123 8.221e-09 1.6898929826812694 8.221999999999999e-09 1.7570651072067978 8.223e-09 1.8202265236365058 8.224e-09 1.7878954699849623 8.225e-09 1.7774632625259557 8.226e-09 1.8173417478147573 8.227e-09 1.7525633947471693 8.228e-09 1.8568916350301639 8.229e-09 1.870213943361815 8.23e-09 1.8854653214752806 8.231e-09 1.7810940811418536 8.232e-09 1.7391333327133243 8.233e-09 1.7330744013285198 8.234e-09 1.9068008293252472 8.235e-09 1.783081634747886 8.236e-09 1.8156622176796098 8.237e-09 1.7654617306808673 8.237999999999999e-09 1.7888835976557262 8.239e-09 1.8202059255637164 8.24e-09 1.796796147774205 8.240999999999999e-09 1.805987034632297 8.242e-09 1.8185427377610717 8.243e-09 1.7298170197838458 8.244e-09 1.778756284163341 8.245e-09 1.7342302703776424 8.246e-09 1.795000388217376 8.247e-09 1.8139485491649918 8.248e-09 1.8541270405822847 8.249e-09 1.7937996687266908 8.25e-09 1.8075514427725576 8.251e-09 1.8406817005436484 8.252e-09 1.763946794230949 8.253e-09 1.7952342281705447 8.254e-09 1.7935236525580216 8.255e-09 1.8860724280011973 8.256e-09 1.7841474465661125 8.256999999999999e-09 1.8534119778033864 8.258e-09 1.7621683750980044 8.259e-09 1.8894505565141488 8.26e-09 1.6849713484501851 8.261e-09 1.7683035084718968 8.262e-09 1.793718241246407 8.263e-09 1.7525003412772544 8.264e-09 1.838317185427782 8.265e-09 1.7961417040248442 8.266e-09 1.8368859660753964 8.267e-09 1.7780006641165507 8.268e-09 1.870977092395936 8.269e-09 1.7709922490812997 8.27e-09 1.7671199830971054 8.271e-09 1.8079218432748119 8.272e-09 1.8012721675035048 8.272999999999999e-09 1.8445148545785204 8.274e-09 1.742950080970311 8.275e-09 1.8084796244057562 8.275999999999999e-09 1.7834301202400993 8.277e-09 1.70909652257173 8.278e-09 1.7605848684089214 8.279e-09 1.7551896323866627 8.28e-09 1.798253849620597 8.281e-09 1.8767885740603045 8.282e-09 1.8498338980274818 8.283e-09 1.8211931153215664 8.284e-09 1.7644889257974883 8.285e-09 1.7985312129425002 8.286e-09 1.7975286459573907 8.287e-09 1.7893816342718842 8.288e-09 1.8057228252664475 8.289e-09 1.8258411952798388 8.29e-09 1.8213847394680853 8.291e-09 1.7870977599165498 8.291999999999999e-09 1.7601521382693233 8.293e-09 1.7850047141952752 8.294e-09 1.7594163982395932 8.294999999999999e-09 1.8069369194969045 8.296e-09 1.8104851595159848 8.297e-09 1.8247970524822337 8.298e-09 1.8081180940911634 8.299e-09 1.836130883045569 8.3e-09 1.8402663110829756 8.301e-09 1.8424687334302503 8.302e-09 1.8015215090018168 8.303e-09 1.7715639651682804 8.304e-09 1.9054942457850128 8.305e-09 1.7767606172523556 8.306e-09 1.7501693310877766 8.307e-09 1.762300108164558 8.307999999999999e-09 1.827216494553979 8.309e-09 1.789819189421142 8.31e-09 1.8349819522828095 8.310999999999999e-09 1.8398445643638233 8.312e-09 1.766101623814545 8.313e-09 1.831998223085153 8.314e-09 1.701100875998923 8.315e-09 1.8432931666296388 8.316e-09 1.7849655954266264 8.317e-09 1.7227160959479786 8.318e-09 1.712883610807378 8.319e-09 1.9053838974797888 8.32e-09 1.7861934912028137 8.321e-09 1.8258584951587924 8.322e-09 1.850029119795065 8.323e-09 1.795439720313226 8.324e-09 1.7651596528999407 8.325e-09 1.8470542269948724 8.326e-09 1.7828089573685533 8.326999999999999e-09 1.852022619771876 8.328e-09 1.7375353510559837 8.329e-09 1.803930602204362 8.329999999999999e-09 1.6712586505666516 8.331e-09 1.775624261162674 8.332e-09 1.7781728024223944 8.333e-09 1.6404591124746246 8.334e-09 1.8082467673861757 8.335e-09 1.8316515016692996 8.336e-09 1.7950632255344443 8.337e-09 1.7101779382941096 8.338e-09 1.7398588415711347 8.339e-09 1.7927612861257645 8.34e-09 1.8262674444826954 8.341e-09 1.8274001285912818 8.342e-09 1.7694253274409535 8.343e-09 1.774321377741003 8.344e-09 1.8414972717915072 8.345e-09 1.7476146096145224 8.345999999999999e-09 1.7720832658214805 8.347e-09 1.8972318368089736 8.348e-09 1.80875471637749 8.349e-09 1.8554378102446012 8.35e-09 1.8400481473775432 8.351e-09 1.7399473417106188 8.352e-09 1.762837283206482 8.353e-09 1.8623609778854877 8.354e-09 1.8352977303162534 8.355e-09 1.7614390218435099 8.356e-09 1.8051247637608387 8.357e-09 1.756223207718421 8.358e-09 1.7647944555438295 8.359e-09 1.8872406227200276 8.36e-09 1.761606117589668 8.361e-09 1.7877705625586826 8.361999999999999e-09 1.787965469972172 8.363e-09 1.8659764459256638 8.364e-09 1.7539185114476232 8.364999999999999e-09 1.776041411323852 8.366e-09 1.787265080343271 8.367e-09 1.785087959105819 8.368e-09 1.8080766769852537 8.369e-09 1.8640381912808413 8.37e-09 1.7873965435360388 8.371e-09 1.847593299192147 8.372e-09 1.8395250004814798 8.373e-09 1.878868352145798 8.374e-09 1.7910637520596158 8.375e-09 1.823684549573776 8.376e-09 1.7513352778545848 8.377e-09 1.803135540670822 8.378e-09 1.8109708737529553 8.379e-09 1.7941698458524833 8.38e-09 1.8131406139483195 8.380999999999999e-09 1.826922983190269 8.382e-09 1.8413994251539643 8.383e-09 1.7521964707981397 8.383999999999999e-09 1.8093198756586504 8.385e-09 1.8136866757223302 8.386e-09 1.8443838445007645 8.387e-09 1.7556544749037308 8.388e-09 1.8362531851496509 8.389e-09 1.7491292202259234 8.39e-09 1.7387714509331125 8.391e-09 1.8439588496266355 8.392e-09 1.7262971781392469 8.393e-09 1.8897574423065644 8.394e-09 1.775205001244436 8.395e-09 1.7739359286870966 8.396e-09 1.7905376407363804 8.396999999999999e-09 1.779361399967393 8.398e-09 1.8266728127438754 8.399e-09 1.8470028961054532 8.399999999999999e-09 1.8126859911107764 8.401e-09 1.711431506062177 8.402e-09 1.8179472275942987 8.403e-09 1.8035799250053082 8.404e-09 1.8335414491557647 8.405e-09 1.727779664793173 8.406e-09 1.7835071610575481 8.407e-09 1.8290838474102395 8.408e-09 1.8632714134896062 8.409e-09 1.7777508383044416 8.41e-09 1.8046830676890933 8.411e-09 1.813998509422242 8.412e-09 1.9629057701715973 8.413e-09 1.7623503827391522 8.414e-09 1.7368210741149959 8.415e-09 1.8956311675114368 8.415999999999999e-09 1.8163212167360747 8.417e-09 1.889969051601682 8.418e-09 1.7901070054799695 8.418999999999999e-09 1.7474539725473175 8.42e-09 1.7861276238851878 8.421e-09 1.6657132038672988 8.422e-09 1.8401251108116259 8.423e-09 1.7271686818706744 8.424e-09 1.9184627223129966 8.425e-09 1.7970793386897979 8.426e-09 1.741339776530953 8.427e-09 1.842549959812395 8.428e-09 1.805041998837929 8.429e-09 1.830207631033703 8.43e-09 1.7493469299845126 8.431e-09 1.7858083827322417 8.431999999999999e-09 1.7886586316204678 8.433e-09 1.7759095396018365 8.434e-09 1.8141060997647618 8.434999999999999e-09 1.7921354532157108 8.436e-09 1.8409885854660029 8.437e-09 1.7955395165062935 8.438e-09 1.8744034956658933 8.439e-09 1.7879710238795743 8.44e-09 1.7343797129129512 8.441e-09 1.824342326634583 8.442e-09 1.766638340443513 8.443e-09 1.8399461664633656 8.444e-09 1.816833516108194 8.445e-09 1.7469262067119535 8.446e-09 1.7888710564247454 8.447e-09 1.7611723812426023 8.448e-09 1.7544654324253308 8.449e-09 1.7853457172692981 8.45e-09 1.810414540431153 8.450999999999999e-09 1.736881961889966 8.452e-09 1.8716170362609048 8.453e-09 1.6453053434567568 8.453999999999999e-09 1.833868280293712 8.455e-09 1.711236776925016 8.456e-09 1.8420881508856515 8.457e-09 1.7084850306323458 8.458e-09 1.7899732457955169 8.459e-09 1.8343433545760497 8.46e-09 1.7994817066270252 8.461e-09 1.7705609818097863 8.462e-09 1.804705692398344 8.463e-09 1.7950797326992798 8.464e-09 1.787556631384267 8.465e-09 1.7679167104434705 8.466e-09 1.8294205479375647 8.467e-09 1.6885279073031534 8.468e-09 1.8464210493060582 8.469e-09 1.8339241235340071 8.469999999999999e-09 1.752673878403395 8.471e-09 1.7545351889223946 8.472e-09 1.8357528210314986 8.473e-09 1.7750085676867176 8.474e-09 1.7427328662427537 8.475e-09 1.86986514623464 8.476e-09 1.838236579646003 8.477e-09 1.8023934929085208 8.478e-09 1.7618527842638518 8.479e-09 1.7756144958950564 8.48e-09 1.828406036626471 8.481e-09 1.8165910334193585 8.482e-09 1.868097639281304 8.483e-09 1.77624787640604 8.484e-09 1.7071110897259403 8.485e-09 1.805716556317729 8.485999999999999e-09 1.8393295671416905 8.487e-09 1.7745774957771514 8.488e-09 1.8748289954302668 8.488999999999999e-09 1.8355829239837518 8.49e-09 1.7841365806890777 8.491e-09 1.86576258367803 8.492e-09 1.8141329229230658 8.493e-09 1.747228679386439 8.494e-09 1.793003462356038 8.495e-09 1.7897298704971558 8.496e-09 1.8581921330912268 8.497e-09 1.8135059427952214 8.498e-09 1.869695663791736 8.499e-09 1.8235515843922976 8.5e-09 1.7930610840108554 8.501e-09 1.8627247315107605 8.502e-09 1.781034237888221 8.503e-09 1.8518510308774037 8.504e-09 1.735394538920977 8.504999999999999e-09 1.7935409847919566 8.506e-09 1.7973595905438327 8.507e-09 1.82800139360871 8.507999999999999e-09 1.8396363907719173 8.509e-09 1.7878733892077945 8.51e-09 1.8023088302716155 8.511e-09 1.7522618491782715 8.512e-09 1.7869099742996366 8.513e-09 1.80485445928988 8.514e-09 1.7868466755768921 8.515e-09 1.785937204226668 8.516e-09 1.7653092250593037 8.517e-09 1.7419966890575682 8.518e-09 1.8196884098716313 8.519e-09 1.727180934507043 8.52e-09 1.7627463674497879 8.520999999999999e-09 1.7813717789372123 8.522e-09 1.7633873320371554 8.523e-09 1.8000963900913083 8.523999999999999e-09 1.8203442601888686 8.525e-09 1.8520508589875209 8.526e-09 1.7603866970343442 8.527e-09 1.865053217204037 8.528e-09 1.846776623563763 8.529e-09 1.7381739580777409 8.53e-09 1.8583727887772696 8.531e-09 1.7805417308402323 8.532e-09 1.853695918340601 8.533e-09 1.8494133611896633 8.534e-09 1.7378368798448558 8.535e-09 1.80689378180732 8.536e-09 1.8045414503767345 8.537e-09 1.7678299525308627 8.538e-09 1.82905558240111 8.539e-09 1.9573677939027798 8.539999999999999e-09 1.734469287015123 8.541e-09 1.760077778723669 8.542e-09 1.7589328707038552 8.542999999999999e-09 1.856723363851323 8.544e-09 1.9017018755972106 8.545e-09 1.841021705291257 8.546e-09 1.7433994933031025 8.547e-09 1.8189895075745615 8.548e-09 1.7172354492043156 8.549e-09 1.7961112075576213 8.55e-09 1.8055607661833675 8.551e-09 1.7471823197538434 8.552e-09 1.7061489114712427 8.553e-09 1.900104914762571 8.554e-09 1.8491562558548598 8.555e-09 1.8904323300187014 8.556e-09 1.7618453309320117 8.557e-09 1.8047307789481417 8.558e-09 1.8703363334980017 8.558999999999999e-09 1.7542731833765914 8.56e-09 1.717597052692021 8.561e-09 1.7587824235092437 8.562e-09 1.900625696459675 8.563e-09 1.8095259277240299 8.564e-09 1.818828057583585 8.565e-09 1.902915511545372 8.566e-09 1.8861477382821552 8.567e-09 1.8054918261165211 8.568e-09 1.8645382239560966 8.569e-09 1.760540880436139 8.57e-09 1.839561627983849 8.571e-09 1.7405338308046276 8.572e-09 1.8214370210390032 8.573e-09 1.8558873522462014 8.574e-09 1.890096382031215 8.574999999999999e-09 1.7834873795995618 8.576e-09 1.8097309590586315 8.577e-09 1.8640180241195932 8.577999999999999e-09 1.857077223422691 8.579e-09 1.728558282426223 8.58e-09 1.8181748025599223 8.581e-09 1.894348762149526 8.582e-09 1.852252875035359 8.583e-09 1.9113442097965758 8.584e-09 1.896814723844879 8.585e-09 1.7742777335043716 8.586e-09 1.7678017384712796 8.587e-09 1.9090842518574853 8.588e-09 1.7726756985089482 8.589e-09 1.7525368588107628 8.59e-09 1.8244622770184753 8.591e-09 1.8825868728783268 8.592e-09 1.7757621565083117 8.593e-09 1.7734287902341381 8.593999999999999e-09 1.78846852296442 8.595e-09 1.796731845366774 8.596e-09 1.7879821858732932 8.596999999999999e-09 1.7889592930051046 8.598e-09 1.84719951535216 8.599e-09 1.770855266527656 8.6e-09 1.7637028500056742 8.601e-09 1.798929878087515 8.602e-09 1.8139016933738028 8.603e-09 1.79496265235408 8.604e-09 1.7520456506150546 8.605e-09 1.777598418013374 8.606e-09 1.8827322569815759 8.607e-09 1.8201555186668574 8.608e-09 1.8061060484105647 8.609e-09 1.7826813097011152 8.609999999999999e-09 1.6728693185501404 8.611e-09 1.9006218317879842 8.612e-09 1.8518653175467086 8.612999999999999e-09 1.7585436970601276 8.614e-09 1.8478691904721893 8.615e-09 1.7902859852663744 8.616e-09 1.8319269963103932 8.617e-09 1.7761489196737679 8.618e-09 1.8972489184251744 8.619e-09 1.7971729099585176 8.62e-09 1.8475757348230946 8.621e-09 1.7718879626498958 8.622e-09 1.8496906688226036 8.623e-09 1.7047670150427172 8.624e-09 1.8526505637176474 8.625e-09 1.798808000813268 8.626e-09 1.7583340768137155 8.627e-09 1.7263255946089935 8.628e-09 1.7905432517703874 8.628999999999999e-09 1.7579118234230016 8.63e-09 1.7928458979428008 8.631e-09 1.8168362264748976 8.631999999999999e-09 1.7569778589910716 8.633e-09 1.7515555677459644 8.634e-09 1.8002675718655383 8.635e-09 1.839095470385112 8.636e-09 1.8304439340180878 8.637e-09 1.8116560847417431 8.638e-09 1.8021574498047557 8.639e-09 1.739431051306906 8.64e-09 1.762883870709073 8.641e-09 1.8141637632904022 8.642e-09 1.8101003079261757 8.643e-09 1.8066272921887383 8.644e-09 1.7659808300201396 8.645e-09 1.8438409006302958 8.646e-09 1.8003622477530168 8.647e-09 1.8665196913683137 8.647999999999999e-09 1.7780628301006045 8.649e-09 1.8503237913302795 8.65e-09 1.852039840650609 8.651e-09 1.8624682124750245 8.652e-09 1.8676176424509354 8.653e-09 1.8595715897193226 8.654e-09 1.7077493520692621 8.655e-09 1.7788229831363536 8.656e-09 1.8082827771835728 8.657e-09 1.7813463462712915 8.658e-09 1.8424994220728592 8.659e-09 1.7994955371160473 8.66e-09 1.8228429036257414 8.661e-09 1.8075112591082585 8.662e-09 1.7933574926251112 8.663e-09 1.8543346824209281 8.663999999999999e-09 1.753506703675647 8.665e-09 1.8188096969649092 8.666e-09 1.8294340281316432 8.666999999999999e-09 1.8249825419449126 8.668e-09 1.7641256409554142 8.669e-09 1.8370179872126102 8.67e-09 1.8572500987650227 8.671e-09 1.8346040638000434 8.672e-09 1.7833971067026775 8.673e-09 1.7915714774697011 8.674e-09 1.8466089499988116 8.675e-09 1.8493551432743585 8.676e-09 1.7952685630581218 8.677e-09 1.7648246936169827 8.678e-09 1.8260679696836228 8.679e-09 1.8170347865503618 8.68e-09 1.747683682711722 8.681e-09 1.7750172433660751 8.682e-09 1.7326043649961966 8.682999999999999e-09 1.8088674252951102 8.684e-09 1.725804471061465 8.685e-09 1.7577721821602932 8.685999999999999e-09 1.827652280712917 8.687e-09 1.7538763486801703 8.688e-09 1.7710317071983563 8.689e-09 1.8626905083636478 8.69e-09 1.8015126341885397 8.691e-09 1.7782094570905673 8.692e-09 1.769871485708178 8.693e-09 1.7776838787312288 8.694e-09 1.7813850663514235 8.695e-09 1.7950054345222588 8.696e-09 1.8106549021686695 8.697e-09 1.7905437334040875 8.698e-09 1.8215948046523853 8.698999999999999e-09 1.7554591355072393 8.7e-09 1.8123959017469495 8.701e-09 1.8145100922293522 8.701999999999999e-09 1.840812598175894 8.703e-09 1.7881683607336225 8.704e-09 1.777129579126882 8.705e-09 1.7837812952373762 8.706e-09 1.8579099986302707 8.707e-09 1.7504426696904518 8.708e-09 1.7389373479857118 8.709e-09 1.8380855599305843 8.71e-09 1.7838584847743968 8.711e-09 1.8588843329770008 8.712e-09 1.8621875293622798 8.713e-09 1.7051886547352302 8.714e-09 1.738044174183628 8.715e-09 1.8168427939393765 8.716e-09 1.7861251790767454 8.717e-09 1.9344369814366242 8.717999999999999e-09 1.8555140633800453 8.719e-09 1.8278082521451655 8.72e-09 1.8491215432408685 8.720999999999999e-09 1.7342065756525424 8.722e-09 1.8366589737113899 8.723e-09 1.7734916371588063 8.724e-09 1.7505005617199803 8.725e-09 1.7762916057586364 8.726e-09 1.8171346336965186 8.727e-09 1.7835965214416387 8.728e-09 1.778189344272572 8.729e-09 1.8523613522849443 8.73e-09 1.7699341821897574 8.731e-09 1.8206830340103874 8.732e-09 1.8561059553728902 8.733e-09 1.8280746951220155 8.733999999999999e-09 1.7185005028821547 8.735e-09 1.7885423811305141 8.736e-09 1.7164048003808976 8.736999999999999e-09 1.776026179691345 8.738e-09 1.79898019523107 8.739e-09 1.779130067612888 8.74e-09 1.7730783211117676 8.741e-09 1.8485200645953506 8.742e-09 1.7625902385691852 8.743e-09 1.8422549577323744 8.744e-09 1.7410006305336667 8.745e-09 1.8906858517667204 8.746e-09 1.7899521506247535 8.747e-09 1.7661966268079015 8.748e-09 1.859462541185334 8.749e-09 1.8423810680736232 8.75e-09 1.8657638533304362 8.751e-09 1.815402858627053 8.752e-09 1.8805893386659462 8.752999999999999e-09 1.8611533774791056 8.754e-09 1.8049462379007042 8.755e-09 1.8732640526809734 8.755999999999999e-09 1.7572624699640529 8.757e-09 1.7778711921192585 8.758e-09 1.8771841575381318 8.759e-09 1.7489277089205235 8.76e-09 1.8090029533314875 8.761e-09 1.8062285389313226 8.762e-09 1.8003307711581986 8.763e-09 1.83463686703416 8.764e-09 1.8533377055737825 8.765e-09 1.8114211222645635 8.766e-09 1.8927360857324014 8.767e-09 1.8162795458795256 8.768e-09 1.8341370284195966 8.769e-09 1.6613154534501766 8.77e-09 1.7125992954639755 8.771e-09 1.8302476757504282 8.771999999999999e-09 1.8048400537356364 8.773e-09 1.8057115722309305 8.774e-09 1.813349898553533 8.774999999999999e-09 1.7048838317797765 8.776e-09 1.7642024951595474 8.777e-09 1.856905303380747 8.778e-09 1.8098088713118023 8.779e-09 1.7781758113868869 8.78e-09 1.7688633403477165 8.781e-09 1.7407065794522838 8.782e-09 1.8019777446490186 8.783e-09 1.845188656214756 8.784e-09 1.7737668926868935 8.785e-09 1.903317035829325 8.786e-09 1.8455781375661078 8.787e-09 1.772249258634123 8.787999999999999e-09 1.8401825228828104 8.789e-09 1.884175715762821 8.79e-09 1.8530916001819482 8.790999999999999e-09 1.7090207991310193 8.792e-09 1.796306845163494 8.793e-09 1.7869749898152307 8.794e-09 1.807310714773045 8.795e-09 1.7192259614329952 8.796e-09 1.7947773329630339 8.797e-09 1.7978965998025247 8.798e-09 1.678579850017567 8.799e-09 1.8216585978027044 8.8e-09 1.8139617946822404 8.801e-09 1.8966209784743138 8.802e-09 1.7247663388611207 8.803e-09 1.8000850889225675 8.804e-09 1.7262755744709786 8.805e-09 1.8197977320250387 8.806e-09 1.7571383476866413 8.806999999999999e-09 1.8851729917273206 8.808e-09 1.8401266982951885 8.809e-09 1.6734304847751347 8.809999999999999e-09 1.7835508485949958 8.811e-09 1.827097900749582 8.812e-09 1.824556721551488 8.813e-09 1.8205879468542323 8.814e-09 1.8639527063886443 8.815e-09 1.6922777981058672 8.816e-09 1.7301844344365398 8.817e-09 1.7828925221778704 8.818e-09 1.8311698122791467 8.819e-09 1.817004339386261 8.82e-09 1.8344798823737574 8.821e-09 1.77193212631504 8.822e-09 1.8235410662728748 8.822999999999999e-09 1.8198687165149936 8.824e-09 1.7685514999705827 8.825e-09 1.7598670394422629 8.825999999999999e-09 1.830216347220267 8.827e-09 1.7950799644784539 8.828e-09 1.7720056187705144 8.829e-09 1.8117559844279016 8.83e-09 1.8776700815644056 8.831e-09 1.743628989100848 8.832e-09 1.8432672256100089 8.833e-09 1.8663675368207517 8.834e-09 1.8056298419869503 8.835e-09 1.7900024638520737 8.836e-09 1.8526819966672328 8.837e-09 1.7284142376516574 8.838e-09 1.8007798886427033 8.839e-09 1.8049148424877954 8.84e-09 1.7454428956114854 8.841e-09 1.7262766548329997 8.841999999999999e-09 1.823352336225432 8.843e-09 1.8256803629951228 8.844e-09 1.739628541784846 8.844999999999999e-09 1.8119896599093048 8.846e-09 1.7597736430704776 8.847e-09 1.900095178244731 8.848e-09 1.9044054030760058 8.849e-09 1.8270232263731596 8.85e-09 1.8703248426097299 8.851e-09 1.8667710007846097 8.852e-09 1.8473108931430928 8.853e-09 1.887916181835258 8.854e-09 1.785060533746779 8.855e-09 1.7426455517598973 8.856e-09 1.8075057745173682 8.857e-09 1.8467597930915856 8.858e-09 1.8214969576444273 8.859e-09 1.7854244669849522 8.86e-09 1.8063741739821735 8.860999999999999e-09 1.7122669864995053 8.862e-09 1.8837243550425404 8.863e-09 1.8207903497019429 8.863999999999999e-09 1.8155332616216 8.865e-09 1.7302653006575062 8.866e-09 1.9017572045350815 8.867e-09 1.7693838282796743 8.868e-09 1.8294644141890415 8.869e-09 1.6847334181353766 8.87e-09 1.6876571873306894 8.871e-09 1.8445016106310936 8.872e-09 1.8367280006631037 8.873e-09 1.8152529989105908 8.874e-09 1.7313700981368898 8.875e-09 1.806322411506412 8.876e-09 1.7767297689593353 8.876999999999999e-09 1.8258290334398355 8.878e-09 1.826389170510413 8.879e-09 1.854239685062546 8.879999999999999e-09 1.7694455974184338 8.881e-09 1.7481809858409274 8.882e-09 1.82552931466469 8.883e-09 1.7885897318046438 8.884e-09 1.7902336285561005 8.885e-09 1.8249675557240663 8.886e-09 1.76859724709115 8.887e-09 1.7987486581781205 8.888e-09 1.8841037709851036 8.889e-09 1.7881281195234613 8.89e-09 1.8425198502072093 8.891e-09 1.8223319053323022 8.892e-09 1.8716843786986888 8.893e-09 1.8483367835606237 8.894e-09 1.8707929404836434 8.895e-09 1.7707759407831118 8.895999999999999e-09 1.8459524866924968 8.897e-09 1.7263162021204703 8.898e-09 1.8238166551242359 8.898999999999999e-09 1.7886063249175255 8.9e-09 1.7799719042145032 8.901e-09 1.7671041821768763 8.902e-09 1.7900842659100926 8.903e-09 1.8053122619964934 8.904e-09 1.8232663173052466 8.905e-09 1.7770945923746604 8.906e-09 1.7867536359490495 8.907e-09 1.824397678811402 8.908e-09 1.8293674172293688 8.909e-09 1.7705639199172487 8.91e-09 1.7297929289513894 8.911e-09 1.7470012684617124 8.911999999999999e-09 1.7888408374321119 8.913e-09 1.7739800515609845 8.914e-09 1.8097252835608741 8.914999999999999e-09 1.8074016553802719 8.916e-09 1.7967089343676006 8.917e-09 1.7391532414715178 8.918e-09 1.7883989318437346 8.919e-09 1.7915819582201904 8.92e-09 1.8542128303471925 8.921e-09 1.7207708374530446 8.922e-09 1.791621757528347 8.923e-09 1.7041078524014897 8.924e-09 1.7687545524466262 8.925e-09 1.7438226010431008 8.926e-09 1.7695331131923477 8.927e-09 1.8110585632810627 8.928e-09 1.7594569646084213 8.929e-09 1.7564189622727497 8.93e-09 1.8800727472350396 8.930999999999999e-09 1.798203124988435 8.932e-09 1.7404105692882406 8.933e-09 1.886490198779438 8.933999999999999e-09 1.7635368580746547 8.935e-09 1.7831964241192932 8.936e-09 1.8263769596844373 8.937e-09 1.7677251465956927 8.938e-09 1.9079674213702136 8.939e-09 1.8492694907562106 8.94e-09 1.8474591960973132 8.941e-09 1.8556706591461645 8.942e-09 1.7782563037623706 8.943e-09 1.7745451088662265 8.944e-09 1.7805804205362785 8.945e-09 1.7260099123478643 8.946e-09 1.8365496653304882 8.947e-09 1.7619913984107731 8.948e-09 1.8015281463995185 8.949e-09 1.841393679622842 8.949999999999999e-09 1.709130257160823 8.951e-09 1.7767856026492177 8.952e-09 1.750112501541437 8.952999999999999e-09 1.8429691700760598 8.954e-09 1.7829934800815586 8.955e-09 1.7901806864755119 8.956e-09 1.7806014975095692 8.957e-09 1.7480871474036281 8.958e-09 1.7818512088594627 8.959e-09 1.7912734908055354 8.96e-09 1.8082523551963077 8.961e-09 1.780095772548912 8.962e-09 1.8226352098882346 8.963e-09 1.8211659311085764 8.964e-09 1.7886353302124305 8.965e-09 1.730822005533537 8.965999999999999e-09 1.7870503452005657 8.967e-09 1.7910518262617006 8.968e-09 1.732127650438082 8.968999999999999e-09 1.729033958324276 8.97e-09 1.705915700832831 8.971e-09 1.8770193114731542 8.972e-09 1.758118543028292 8.973e-09 1.807724977003028 8.974e-09 1.7771166999320998 8.975e-09 1.8464258652620003 8.976e-09 1.811166079572367 8.977e-09 1.7892942009180084 8.978e-09 1.757338630831547 8.979e-09 1.8452816514100419 8.98e-09 1.7498264467683595 8.981e-09 1.857904187995574 8.982e-09 1.8286271920528863 8.983e-09 1.799581439805413 8.984e-09 1.8151532524574687 8.984999999999999e-09 1.7540419354964079 8.986e-09 1.8255059229982216 8.987e-09 1.8149838090380603 8.987999999999999e-09 1.6727659803493615 8.989e-09 1.8196552487040651 8.99e-09 1.7441219586056078 8.991e-09 1.789277500270405 8.992e-09 1.7622276451913221 8.993e-09 1.8306659583945695 8.994e-09 1.7952263698635569 8.995e-09 1.7887368601022118 8.996e-09 1.8674814994451416 8.997e-09 1.7637018917107277 8.998e-09 1.884936553425829 8.999e-09 1.7322410266699435 9e-09 1.862161542130674 9.000999999999999e-09 1.820595916021147 9.002e-09 1.85436586119922 9.003e-09 1.8355786204581344 9.003999999999999e-09 1.7423805940183033 9.005e-09 1.78399736340524 9.006e-09 1.813376715913107 9.007e-09 1.8184686456944237 9.008e-09 1.7372307529351951 9.009e-09 1.8109884968783994 9.01e-09 1.731917784531747 9.011e-09 1.8498279158734854 9.012e-09 1.8272505639199208 9.013e-09 1.8532763040029208 9.014e-09 1.7168921334540577 9.015e-09 1.7463348485897523 9.016e-09 1.8007610296273526 9.017e-09 1.8246462750674772 9.018e-09 1.7535543786527334 9.019e-09 1.8176442709236202 9.019999999999999e-09 1.8450567244742437 9.021e-09 1.7762574473914936 9.022e-09 1.7821601122852406 9.022999999999999e-09 1.7676741488895094 9.024e-09 1.7399454160776344 9.025e-09 1.8151989848112668 9.026e-09 1.881787945860063 9.027e-09 1.7945409867796795 9.028e-09 1.855071366968451 9.029e-09 1.8527387501112964 9.03e-09 1.8470676684767031 9.031e-09 1.824856282232583 9.032e-09 1.8185803145425954 9.033e-09 1.8444195223026845 9.034e-09 1.6467798144060914 9.035e-09 1.8563621053811534 9.036e-09 1.8442273814227972 9.037e-09 1.7436197684040495 9.038e-09 1.7991886512584498 9.038999999999999e-09 1.8951793144932556 9.04e-09 1.7988302009787462 9.041e-09 1.7393697282875842 9.042e-09 1.8224297392727626 9.043e-09 1.7879805205537553 9.044e-09 1.7708067826559204 9.045e-09 1.8367431849109248 9.046e-09 1.720001187102774 9.047e-09 1.7833034521708813 9.048e-09 1.8548289837675629 9.049e-09 1.826137352964801 9.05e-09 1.7756098647173915 9.051e-09 1.7512349723645557 9.052e-09 1.8098030700839607 9.053e-09 1.8723829457251804 9.054e-09 1.805541502665424 9.054999999999999e-09 1.7565630735360196 9.056e-09 1.7613509826411442 9.057e-09 1.77524115560868 9.057999999999999e-09 1.783895486364895 9.059e-09 1.7771602574389473 9.06e-09 1.7606228426277797 9.061e-09 1.809912478533814 9.062e-09 1.775524459744578 9.063e-09 1.8400416715060623 9.064e-09 1.7851027440942828 9.065e-09 1.872062300746827 9.066e-09 1.7400587327446388 9.067e-09 1.7607387869122215 9.068e-09 1.7463918151138154 9.069e-09 1.8291041392013816 9.07e-09 1.7369110764949878 9.071e-09 1.7991058174700685 9.072e-09 1.76305339603298 9.073e-09 1.821143725506007 9.073999999999999e-09 1.8767989547262618 9.075e-09 1.7859781144119942 9.076e-09 1.6956983941888555 9.076999999999999e-09 1.807376569077362 9.078e-09 1.7661636637844058 9.079e-09 1.8396782293363494 9.08e-09 1.8027530030042727 9.081e-09 1.7708691546187563 9.082e-09 1.8602782472258246 9.083e-09 1.7988135161254841 9.084e-09 1.8988972412910927 9.085e-09 1.8791051702960537 9.086e-09 1.7961840523477737 9.087e-09 1.8404098102031596 9.088e-09 1.7664586352842562 9.089e-09 1.8113986493533019 9.089999999999999e-09 1.815425494097421 9.091e-09 1.765299191774051 9.092e-09 1.7938280118242533 9.092999999999999e-09 1.899814038178129 9.094e-09 1.7882326422261527 9.095e-09 1.7957755975826302 9.096e-09 1.8274718396170893 9.097e-09 1.7874439486531555 9.098e-09 1.744795013241747 9.099e-09 1.7140740844088689 9.1e-09 1.7964164770567506 9.101e-09 1.7758058154382874 9.102e-09 1.7905812333381135 9.103e-09 1.811694729436099 9.104e-09 1.802569878947093 9.105e-09 1.8961644526684474 9.106e-09 1.8192730616227935 9.107e-09 1.7573836194451473 9.108e-09 1.751195016113559 9.108999999999999e-09 1.8203951047844382 9.11e-09 1.8146715980065447 9.111e-09 1.8258127386011795 9.111999999999999e-09 1.7435724393458782 9.113e-09 1.8091096144579966 9.114e-09 1.8143015677458683 9.115e-09 1.8452423584073543 9.116e-09 1.7759960663378296 9.117e-09 1.7708126684343015 9.118e-09 1.8617162582137192 9.119e-09 1.8155723775904546 9.12e-09 1.7387699664160219 9.121e-09 1.7692569776569675 9.122e-09 1.8005215712849771 9.123e-09 1.8754241786916785 9.124e-09 1.849194603019571 9.124999999999999e-09 1.83848896215432 9.126e-09 1.7680409932922831 9.127e-09 1.8316543691295382 9.127999999999999e-09 1.7419564869240116 9.129e-09 1.8265469263308896 9.13e-09 1.7841182054557492 9.131e-09 1.808997070327346 9.132e-09 1.7340903874084204 9.133e-09 1.8194295579436324 9.134e-09 1.889226385633703 9.135e-09 1.7518027608461133 9.136e-09 1.8470968917803452 9.137e-09 1.8143063517951843 9.138e-09 1.7769655637769224 9.139e-09 1.8552577798649017 9.14e-09 1.7695351568013473 9.141e-09 1.767874152229515 9.142e-09 1.7461875945517653 9.143e-09 1.800575820486268 9.143999999999999e-09 1.8300942714070676 9.145e-09 1.9224038560597048 9.146e-09 1.8312989710881806 9.146999999999999e-09 1.8431072167376799 9.148e-09 1.8021897923823822 9.149e-09 1.7282530407521741 9.15e-09 1.7906892493908124 9.151e-09 1.732392025359514 9.152e-09 1.801987925727516 9.153e-09 1.753377592177459 9.154e-09 1.810131414723837 9.155e-09 1.789813355318692 9.156e-09 1.789752905366089 9.157e-09 1.806107272993216 9.158e-09 1.7519473565612356 9.159e-09 1.7503714175684162 9.16e-09 1.737850393385416 9.161e-09 1.7532599072996455 9.162e-09 1.833529534026531 9.162999999999999e-09 1.8589485035117377 9.164e-09 1.7971906370912705 9.165e-09 1.8585403971845713 9.165999999999999e-09 1.7816673074751734 9.167e-09 1.7756730291798 9.168e-09 1.7856036644648756 9.169e-09 1.8041801828374993 9.17e-09 1.7495089919484341 9.171e-09 1.8422047753888513 9.172e-09 1.8088795016354453 9.173e-09 1.7776264173497787 9.174e-09 1.8007179975444387 9.175e-09 1.8351905135648887 9.176e-09 1.7993926825270385 9.177e-09 1.7675575070007647 9.178e-09 1.7895049780067738 9.178999999999999e-09 1.7784187351569527 9.18e-09 1.847071621066369 9.181e-09 1.7978850922567882 9.181999999999999e-09 1.8021583273492814 9.183e-09 1.8144990404827177 9.184e-09 1.835530534287422 9.185e-09 1.8162591981477538 9.186e-09 1.8044985379315974 9.187e-09 1.7892826300847824 9.188e-09 1.8278076535789132 9.189e-09 1.7833318912462404 9.19e-09 1.7984198988604012 9.191e-09 1.6916090318176373 9.192e-09 1.8122946292799293 9.193e-09 1.8731054441252497 9.194e-09 1.8202594094519053 9.195e-09 1.8434586313196533 9.196e-09 1.8104349221512959 9.197e-09 1.7004374091213932 9.197999999999999e-09 1.8168673258529782 9.199e-09 1.7314278981992715 9.2e-09 1.8280388641212406 9.200999999999999e-09 1.9041313254716288 9.202e-09 1.8009330167543653 9.203e-09 1.8014992480237746 9.204e-09 1.7619956949768876 9.205e-09 1.6684892706721448 9.206e-09 1.878473539494817 9.207e-09 1.8432606724664762 9.208e-09 1.907756642405081 9.209e-09 1.7918135830474218 9.21e-09 1.7746820548169686 9.211e-09 1.7816472316598695 9.212e-09 1.691297612135509 9.213e-09 1.7432986231687324 9.213999999999999e-09 1.8017301643391235 9.215e-09 1.8049967642894313 9.216e-09 1.8108845427474705 9.216999999999999e-09 1.7809967308857777 9.218e-09 1.8220818553551352 9.219e-09 1.8030210533155686 9.22e-09 1.8614500002286667 9.221e-09 1.8189258438168747 9.222e-09 1.8158515088156568 9.223e-09 1.8339388592115802 9.224e-09 1.7716721453633373 9.225e-09 1.8486527177778405 9.226e-09 1.823909671385163 9.227e-09 1.8260456427118623 9.228e-09 1.8372092779617335 9.229e-09 1.7371325429250202 9.23e-09 1.6837614488573878 9.231e-09 1.8294499182563384 9.232e-09 1.760392655245896 9.232999999999999e-09 1.8224263855719807 9.234e-09 1.6942336476525548 9.235e-09 1.7668022278956204 9.235999999999999e-09 1.822999890358145 9.237e-09 1.8532452374982367 9.238e-09 1.7787812197135806 9.239e-09 1.7433145741383562 9.24e-09 1.8045260464418684 9.241e-09 1.8028672442183362 9.242e-09 1.7614773792837901 9.243e-09 1.8499551311183506 9.244e-09 1.8223023124785778 9.245e-09 1.7741058106797964 9.246e-09 1.7714013729816804 9.247e-09 1.7189656721460032 9.248e-09 1.8119263786365714 9.249e-09 1.7758434193528403 9.25e-09 1.757625471753435 9.251e-09 1.8160005731978566 9.251999999999999e-09 1.8289406948629854 9.253e-09 1.8340751934668091 9.254e-09 1.8755773256165444 9.254999999999999e-09 1.8017552615919867 9.256e-09 1.8094130953648124 9.257e-09 1.787114413228938 9.258e-09 1.8336341271043028 9.259e-09 1.859116703998913 9.26e-09 1.8049925913144516 9.261e-09 1.782431376837881 9.262e-09 1.7718526182594887 9.263e-09 1.8334995090920445 9.264e-09 1.7575235339638788 9.265e-09 1.8196329575328956 9.266e-09 1.8624588128984731 9.267e-09 1.7736401115670737 9.267999999999999e-09 1.7758837260367824 9.269e-09 1.8913421652583908 9.27e-09 1.7543244736767376 9.270999999999999e-09 1.8530682339751652 9.272e-09 1.7397586655171178 9.273e-09 1.7286261822207065 9.274e-09 1.798103923401957 9.275e-09 1.8087327886951527 9.276e-09 1.7048649415330854 9.277e-09 1.8364375743632793 9.278e-09 1.7500867641912694 9.279e-09 1.78118393699999 9.28e-09 1.7904385110414323 9.281e-09 1.7612264204855197 9.282e-09 1.7436745707504195 9.283e-09 1.7172110527011781 9.284e-09 1.8276254024591956 9.285e-09 1.8465835564749196 9.286e-09 1.852350115918375 9.286999999999999e-09 1.7789735221171559 9.288e-09 1.810091814643922 9.289e-09 1.799268473846473 9.289999999999999e-09 1.8733235170831395 9.291e-09 1.8054001191549043 9.292e-09 1.8249061290732 9.293e-09 1.8005501614944877 9.294e-09 1.8379200178743853 9.295e-09 1.8583944859892885 9.296e-09 1.7089390715403354 9.297e-09 1.7889513050912262 9.298e-09 1.7626140732378137 9.299e-09 1.869880119352345 9.3e-09 1.7740059016089589 9.301e-09 1.7499187262691498 9.302e-09 1.8296378879681632 9.302999999999999e-09 1.76638450714189 9.304e-09 1.8326701063587452 9.305e-09 1.7534779508246836 9.305999999999999e-09 1.7948641014583648 9.307e-09 1.8334797274919565 9.308e-09 1.7617526963092278 9.309e-09 1.9187001367581842 9.31e-09 1.7909194041211025 9.311e-09 1.8851002615632517 9.312e-09 1.8167198071198962 9.313e-09 1.8123422556871334 9.314e-09 1.7954311292529244 9.315e-09 1.7723445543116745 9.316e-09 1.8116839779613705 9.317e-09 1.6842573055261636 9.318e-09 1.859802658193608 9.319e-09 1.9540023183536452 9.32e-09 1.7304806429075121 9.321e-09 1.8429338542410965 9.321999999999999e-09 1.8312364995703558 9.323e-09 1.7779099729849852 9.324e-09 1.7668470712223145 9.324999999999999e-09 1.808968849064209 9.326e-09 1.7576749409638912 9.327e-09 1.7911887745319164 9.328e-09 1.7955370936147226 9.329e-09 1.8235421368914033 9.33e-09 1.7662264678318988 9.331e-09 1.8023908956354509 9.332e-09 1.789944737989632 9.333e-09 1.7919603309499084 9.334e-09 1.820839802694583 9.335e-09 1.8386288053803768 9.336e-09 1.820064890010928 9.337e-09 1.8186109402425514 9.338e-09 1.8180665219640582 9.339e-09 1.8119447564407967 9.34e-09 1.9112693945360717 9.340999999999999e-09 1.775858731919242 9.342e-09 1.7290665257916502 9.343e-09 1.7511280388253163 9.343999999999999e-09 1.8185767882071244 9.345e-09 1.9085430241989827 9.346e-09 1.8243230790906355 9.347e-09 1.8008558941264166 9.348e-09 1.8388394762111324 9.349e-09 1.677311917333038 9.35e-09 1.786104476022237 9.351e-09 1.7928072048823371 9.352e-09 1.7566635237661063 9.353e-09 1.7545394555287843 9.354e-09 1.7614088019672012 9.355e-09 1.8532243190251625 9.356e-09 1.842387013168047 9.356999999999999e-09 1.7747530929883406 9.358e-09 1.7870498940062052 9.359e-09 1.8028502094114147 9.359999999999999e-09 1.8254464471051193 9.361e-09 1.793447408750225 9.362e-09 1.8680542089054901 9.363e-09 1.8658558548465534 9.364e-09 1.8544144339121191 9.365e-09 1.7546747594129668 9.366e-09 1.8484323780082415 9.367e-09 1.8081671382395843 9.368e-09 1.8074762421834614 9.369e-09 1.7993610838374452 9.37e-09 1.7383702267185754 9.371e-09 1.8360617268000596 9.372e-09 1.8276607872368713 9.373e-09 1.8814823951515929 9.374e-09 1.74042993945736 9.375e-09 1.841273072094929 9.375999999999999e-09 1.7244676413689133 9.377e-09 1.8348542797675296 9.378e-09 1.8176787740566105 9.378999999999999e-09 1.8990657850362624 9.38e-09 1.8605916670832607 9.381e-09 1.770823290340351 9.382e-09 1.7664746650389616 9.383e-09 1.7852088467786127 9.384e-09 1.788078322992566 9.385e-09 1.8123847740589532 9.386e-09 1.8335965101197809 9.387e-09 1.8571137045215378 9.388e-09 1.8595602954083037 9.389e-09 1.7907474789481759 9.39e-09 1.7091227368678543 9.391e-09 1.7434553235871166 9.391999999999999e-09 1.747165213788354 9.393e-09 1.7687589427058807 9.394e-09 1.852784654033671 9.394999999999999e-09 1.7687593394674042 9.396e-09 1.809015390718217 9.397e-09 1.855023927072748 9.398e-09 1.7034212991466524 9.399e-09 1.817517493542678 9.4e-09 1.7200861221613475 9.401e-09 1.9231495736045185 9.402e-09 1.8911158175648837 9.403e-09 1.8388732923977296 9.404e-09 1.7820468953006579 9.405e-09 1.7970062028248706 9.406e-09 1.8502539469350026 9.407e-09 1.774896622426956 9.408e-09 1.8303171543229244 9.409e-09 1.807192091286008 9.41e-09 1.7529849137829905 9.410999999999999e-09 1.723742380377981 9.412e-09 1.791171921388248 9.413e-09 1.8182392776130796 9.413999999999999e-09 1.7690000352807642 9.415e-09 1.78847794181849 9.416e-09 1.8552512048467555 9.417e-09 1.8113492135640021 9.418e-09 1.7934099982112357 9.419e-09 1.7645227754093147 9.42e-09 1.819058126235412 9.421e-09 1.7285890078668669 9.422e-09 1.8598133873281215 9.423e-09 1.7520949145571472 9.424e-09 1.8647071921831488 9.425e-09 1.8223617671079229 9.426e-09 1.8971920886536868 9.427e-09 1.7782007151813763 9.428e-09 1.7282672283516032 9.429e-09 1.8062415416006716 9.429999999999999e-09 1.853993359281559 9.431e-09 1.8553501581726686 9.432e-09 1.7394955334437585 9.432999999999999e-09 1.7701194619103484 9.434e-09 1.7841622282772962 9.435e-09 1.7573216816477024 9.436e-09 1.7763186456309201 9.437e-09 1.835827054494171 9.438e-09 1.7506629422599254 9.439e-09 1.8065431600491177 9.44e-09 1.8331982372651838 9.441e-09 1.7918829488935701 9.442e-09 1.8815139199165085 9.443e-09 1.7865536135420939 9.444e-09 1.807544876796569 9.445e-09 1.8109971561342384 9.445999999999999e-09 1.8770707331625216 9.447e-09 1.7567505398349677 9.448e-09 1.7917280243582792 9.448999999999999e-09 1.8524128760826073 9.45e-09 1.7746078556526805 9.451e-09 1.8389608511603057 9.452e-09 1.8127819836544332 9.453e-09 1.8059766075943857 9.454e-09 1.8690171587098017 9.455e-09 1.7815993493762823 9.456e-09 1.7447574226825238 9.457e-09 1.7983176134466208 9.458e-09 1.8585004350827374 9.459e-09 1.8211668071839893 9.46e-09 1.8093904808646801 9.461e-09 1.8152783904894307 9.462e-09 1.7708537197387497 9.463e-09 1.7011129389914752 9.464e-09 1.8659523288174993 9.464999999999999e-09 1.7590510575115401 9.466e-09 1.796387760068633 9.467e-09 1.8078259974826776 9.467999999999999e-09 1.8139803360492621 9.469e-09 1.7499383770973147 9.47e-09 1.8598538443110426 9.471e-09 1.8155392394610497 9.472e-09 1.814546827743396 9.473e-09 1.7568306385339876 9.474e-09 1.6919992470561374 9.475e-09 1.7215526727910782 9.476e-09 1.7717680385274306 9.477e-09 1.8407780455415066 9.478e-09 1.8049275236189124 9.479e-09 1.8053585475006717 9.48e-09 1.773572665796351 9.480999999999999e-09 1.8107835688544087 9.482e-09 1.8505279454705315 9.483e-09 1.835009367404982 9.483999999999999e-09 1.8015430854732408 9.485e-09 1.8067702436523896 9.486e-09 1.8624767919353225 9.487e-09 1.7478232328213104 9.488e-09 1.7717252991068646 9.489e-09 1.813699407274841 9.49e-09 1.7571241495244652 9.491e-09 1.8002500846549798 9.492e-09 1.807797205929702 9.493e-09 1.7771182220279604 9.494e-09 1.7252856600965272 9.495e-09 1.7628246317253424 9.496e-09 1.8049658289061665 9.497e-09 1.702496455152845 9.498e-09 1.7985230060250048 9.499e-09 1.883088940572621 9.499999999999999e-09 1.793558690776274 9.501e-09 1.6582295886924459 9.502e-09 1.8073874474659881 9.502999999999999e-09 1.7463447001357764 9.504e-09 1.916558330497221 9.505e-09 1.8375542404859784 9.506e-09 1.8249493766773546 9.507e-09 1.8297922278225358 9.508e-09 1.827714230623757 9.509e-09 1.6954869220023363 9.51e-09 1.859257964802922 9.511e-09 1.8234538929816182 9.512e-09 1.8047871912723408 9.513e-09 1.716121538791011 9.514e-09 1.834817751598214 9.515e-09 1.8199325880852808 9.515999999999999e-09 1.71550614824781 9.517e-09 1.7272982278078648 9.518e-09 1.75605166508996 9.518999999999999e-09 1.8405213038489863 9.52e-09 1.8982254321879635 9.521e-09 1.8311479787192233 9.521999999999999e-09 1.838773746895227 9.523e-09 1.8496851886372707 9.524e-09 1.8459084491947273 9.525e-09 1.8444782572566918 9.526e-09 1.8222158781280455 9.527e-09 1.7431570271337555 9.528e-09 1.77104164641388 9.529e-09 1.760217474705547 9.53e-09 1.7154959682349613 9.531e-09 1.8572022786403546 9.532e-09 1.8313907216687457 9.533e-09 1.783392791333575 9.534e-09 1.8364996047237432 9.534999999999999e-09 1.7707126986685242 9.536e-09 1.7742016874264126 9.537e-09 1.8853279453925418 9.537999999999999e-09 1.9214205314684585 9.539e-09 1.7940209455889025 9.54e-09 1.7456596532856588 9.541e-09 1.8582384326559804 9.542e-09 1.7370365502117182 9.543e-09 1.775317059630999 9.544e-09 1.674455244627234 9.545e-09 1.8492786677568132 9.546e-09 1.7378400604414184 9.547e-09 1.7709666219452191 9.548e-09 1.7473792324511688 9.549e-09 1.8135833964771408 9.55e-09 1.7874478494417507 9.551e-09 1.711874314061855 9.552e-09 1.7999655643443078 9.553e-09 1.8294329344548506 9.553999999999999e-09 1.8058859078676797 9.555e-09 1.8161361271523786 9.556e-09 1.7889731159152442 9.556999999999999e-09 1.765252680206729 9.558e-09 1.792095031745102 9.559e-09 1.75307246999526 9.56e-09 1.8958120531908569 9.561e-09 1.811527529160115 9.562e-09 1.782765449310952 9.563e-09 1.76647646754831 9.564e-09 1.7220442371426607 9.565e-09 1.8237784097138072 9.566e-09 1.7793632222926752 9.567e-09 1.8463631264609504 9.568e-09 1.7963367825575383 9.569e-09 1.790734031649771 9.569999999999999e-09 1.7978138404731432 9.571e-09 1.7975806324635597 9.572e-09 1.8156124021920446 9.572999999999999e-09 1.7855503167646727 9.574e-09 1.8130594590551294 9.575e-09 1.8168962597251601 9.576e-09 1.804578070389767 9.577e-09 1.8426002215037414 9.578e-09 1.7981034234987516 9.579e-09 1.7688162266214689 9.58e-09 1.812249259091485 9.581e-09 1.834228208412468 9.582e-09 1.8329121972423126 9.583e-09 1.7893104698334021 9.584e-09 1.8124995831637585 9.585e-09 1.7921814880710865 9.586e-09 1.7588907472448307 9.587e-09 1.7741614802567682 9.588e-09 1.750129954847077 9.588999999999999e-09 1.7973273706639212 9.59e-09 1.865018517207779 9.591e-09 1.845655493466223 9.591999999999999e-09 1.7339365706218959 9.593e-09 1.7745956381736299 9.594e-09 1.8524941853999468 9.595e-09 1.7923925154313913 9.596e-09 1.8643389693883878 9.597e-09 1.766898008184657 9.598e-09 1.8485316164348895 9.599e-09 1.82412923970912 9.6e-09 1.7941473001032722 9.601e-09 1.8141427763754776 9.602e-09 1.7843813342114538 9.603e-09 1.8656643866388758 9.604e-09 1.797252271594295 9.604999999999999e-09 1.7855071834700305 9.606e-09 1.8910070397541692 9.607e-09 1.8565806505625497 9.607999999999999e-09 1.8621833191835728 9.609e-09 1.858798435064562 9.61e-09 1.7858797805044806 9.611e-09 1.81754218643839 9.612e-09 1.8136059872275327 9.613e-09 1.823240820278523 9.614e-09 1.8669239154380644 9.615e-09 1.8157591827105724 9.616e-09 1.828461218338658 9.617e-09 1.7287045009016484 9.618e-09 1.891128304793121 9.619e-09 1.8713434856762639 9.62e-09 1.7233213300883656 9.621e-09 1.7902113797768728 9.622e-09 1.8330024486392122 9.623e-09 1.8455223174908253 9.623999999999999e-09 1.7185853326799265 9.625e-09 1.8095124784774357 9.626e-09 1.7983426886149638 9.626999999999999e-09 1.8995147553469898 9.628e-09 1.8237491699066501 9.629e-09 1.8664942189072116 9.63e-09 1.8311889055762987 9.631e-09 1.759756930874704 9.632e-09 1.7807355011485317 9.633e-09 1.835055324632201 9.634e-09 1.8208038628677587 9.635e-09 1.8364145337157451 9.636e-09 1.7956510035851077 9.637e-09 1.774842551089638 9.638e-09 1.815457281078414 9.639e-09 1.774958253403978 9.64e-09 1.7919681979560818 9.641e-09 1.8628090834299902 9.642e-09 1.695217039785049 9.642999999999999e-09 1.742595410683775 9.644e-09 1.7723645439730313 9.645e-09 1.7713853633525563 9.645999999999999e-09 1.7544461452872802 9.647e-09 1.886595019563667 9.648e-09 1.801217366478721 9.649e-09 1.8012930678658903 9.65e-09 1.727499749317477 9.651e-09 1.8152175294812618 9.652e-09 1.8542230811689269 9.653e-09 1.7923659317252514 9.654e-09 1.8844691471319641 9.655e-09 1.8087547796927959 9.656e-09 1.7451308097742286 9.657e-09 1.67558782432368 9.658e-09 1.8242584485446185 9.658999999999999e-09 1.7571688532905925 9.66e-09 1.7658211160282171 9.661e-09 1.711031407321687 9.661999999999999e-09 1.7382777546485082 9.663e-09 1.8221472536341552 9.664e-09 1.8124157294801397 9.665e-09 1.8031450553117052 9.666e-09 1.698527914892391 9.667e-09 1.7613576571315046 9.668e-09 1.8103704348242289 9.669e-09 1.824072830167154 9.67e-09 1.8274122566015183 9.671e-09 1.83343874732164 9.672e-09 1.744659087644478 9.673e-09 1.776098662337858 9.674e-09 1.7716071001479219 9.675e-09 1.7236513478633222 9.676e-09 1.8519681009282383 9.677e-09 1.7668835348320264 9.677999999999999e-09 1.7988782285395089 9.679e-09 1.8479575039416434 9.68e-09 1.8221976884495699 9.680999999999999e-09 1.7991220255576057 9.682e-09 1.7935342257662263 9.683e-09 1.7682593825133142 9.684e-09 1.7485192780272263 9.685e-09 1.7739248501237659 9.686e-09 1.799310982361873 9.687e-09 1.8594875708947929 9.688e-09 1.8168964655308528 9.689e-09 1.805081231106402 9.69e-09 1.954534722199731 9.691e-09 1.8050343375802804 9.692e-09 1.7425751023066145 9.693e-09 1.708494905784688 9.693999999999999e-09 1.7649344423307087 9.695e-09 1.7606137221195572 9.696e-09 1.7548199822804706 9.696999999999999e-09 1.8955326050199934 9.698e-09 1.9107767077724802 9.699e-09 1.7942583100945872 9.7e-09 1.8561490151258324 9.701e-09 1.7676723529750298 9.702e-09 1.7046670882448893 9.703e-09 1.7919865972141276 9.704e-09 1.7119258614453392 9.705e-09 1.7588001510045437 9.706e-09 1.8360465705327558 9.707e-09 1.8244827991782526 9.708e-09 1.7322459899709641 9.709e-09 1.7852460045489087 9.71e-09 1.8427054527998927 9.711e-09 1.704872926568834 9.712e-09 1.7469762871036607 9.712999999999999e-09 1.8591860010594827 9.714e-09 1.7691276923758572 9.715e-09 1.8416378926895909 9.715999999999999e-09 1.7326842776018345 9.717e-09 1.7853977646893016 9.718e-09 1.8011285526845389 9.719e-09 1.880008177854214 9.72e-09 1.788663649500878 9.721e-09 1.7880890148155255 9.722e-09 1.7855201334467017 9.723e-09 1.8208134874853812 9.724e-09 1.7231510740591724 9.725e-09 1.8730474182762182 9.726e-09 1.8545650061880172 9.727e-09 1.8046469985923688 9.728e-09 1.8222437145495967 9.729e-09 1.8075806465323216 9.73e-09 1.7742065182319136 9.731e-09 1.7551371147456687 9.731999999999999e-09 1.8404213847441702 9.733e-09 1.7962268472692378 9.734e-09 1.779735305688551 9.734999999999999e-09 1.7640630765988146 9.736e-09 1.7494691485833 9.737e-09 1.8441419718878267 9.738e-09 1.8576703870544968 9.739e-09 1.8089311135057113 9.74e-09 1.8072789848364565 9.741e-09 1.8201074203834469 9.742e-09 1.8574024632579542 9.743e-09 1.8949978667290177 9.744e-09 1.8398585130367775 9.745e-09 1.8783502738538698 9.746e-09 1.8071838830519809 9.747e-09 1.8652209975699339 9.747999999999999e-09 1.8388147004388293 9.749e-09 1.7972021687892044 9.75e-09 1.7486037826140906 9.750999999999999e-09 1.75801457313596 9.752e-09 1.8145893707163505 9.753e-09 1.906354372539734 9.754e-09 1.7567846565386198 9.755e-09 1.8446888907562815 9.756e-09 1.6501516460631065 9.757e-09 1.8530708001010507 9.758e-09 1.8469113121014111 9.759e-09 1.8137823529193806 9.76e-09 1.7500124299596194 9.761e-09 1.7806165409645633 9.762e-09 1.86292678261639 9.763e-09 1.7647209612318293 9.764e-09 1.8112534569961851 9.765e-09 1.7799319879995616 9.766e-09 1.7684290059008116 9.766999999999999e-09 1.816088538957542 9.768e-09 1.8226063285151344 9.769e-09 1.840612209405187 9.769999999999999e-09 1.7755308212309056 9.771e-09 1.8080057095589148 9.772e-09 1.7837396743263554 9.773e-09 1.8739021074270334 9.774e-09 1.8849129617967144 9.775e-09 1.7885966955216441 9.776e-09 1.8381862842066234 9.777e-09 1.7362429584134018 9.778e-09 1.8075122683098945 9.779e-09 1.7903482980104772 9.78e-09 1.7416600370310062 9.781e-09 1.806538314572417 9.782e-09 1.829734994452057 9.782999999999999e-09 1.7838120049539228 9.784e-09 1.7666892349819392 9.785e-09 1.8564636835003627 9.785999999999999e-09 1.9223497865424959 9.787e-09 1.8045560950053054 9.788e-09 1.762353135643425 9.789e-09 1.7693134964478239 9.79e-09 1.8129213158305562 9.791e-09 1.7826304341821997 9.792e-09 1.823469820505325 9.793e-09 1.7701020183942342 9.794e-09 1.6806795309200118 9.795e-09 1.8334953504632634 9.796e-09 1.743366858573195 9.797e-09 1.7551489501075972 9.798e-09 1.912422087429374 9.799e-09 1.845266551405535 9.8e-09 1.8168983907568246 9.801e-09 1.757899967476264 9.801999999999999e-09 1.7386212895692388 9.803e-09 1.8776634613775816 9.804e-09 1.8690702429280739 9.804999999999999e-09 1.7788020603112495 9.806e-09 1.823384224417807 9.807e-09 1.7856858841130205 9.808e-09 1.7859413236841544 9.809e-09 1.808191219367114 9.81e-09 1.8413020013970982 9.811e-09 1.7495569726505862 9.812e-09 1.7907488863232155 9.813e-09 1.8097524039650439 9.814e-09 1.7956574409061754 9.815e-09 1.747979759417759 9.816e-09 1.7494476095198759 9.817e-09 1.7676204038265801 9.817999999999999e-09 1.8434419696316944 9.819e-09 1.8173648786006082 9.82e-09 1.7822011159127589 9.820999999999999e-09 1.7621531920678912 9.822e-09 1.7939860518051802 9.823e-09 1.7626924353512385 9.823999999999999e-09 1.8097421580473114 9.825e-09 1.8347855707145646 9.826e-09 1.756117972990516 9.827e-09 1.7701748133991986 9.828e-09 1.9052180768010354 9.829e-09 1.8067411221506682 9.83e-09 1.7635550246338807 9.831e-09 1.8046697972479588 9.832e-09 1.7743211032414825 9.833e-09 1.8139527783621592 9.834e-09 1.827836404803093 9.835e-09 1.8217604894681911 9.836e-09 1.851878746096413 9.836999999999999e-09 1.8283695064458663 9.838e-09 1.869727728061772 9.839e-09 1.8205298956943539 9.839999999999999e-09 1.797774331649686 9.841e-09 1.7425393571379841 9.842e-09 1.8247927461951396 9.843e-09 1.7645327296155042 9.844e-09 1.7864230264324807 9.845e-09 1.8341638054466647 9.846e-09 1.6819875113952225 9.847e-09 1.7776426750893795 9.848e-09 1.8093722584612888 9.849e-09 1.738269593417968 9.85e-09 1.8116816365062638 9.851e-09 1.8671120057070223 9.852e-09 1.809089711540562 9.853e-09 1.8576455539678165 9.854e-09 1.860684360486487 9.855e-09 1.7879761559901446 9.855999999999999e-09 1.7853710462199504 9.857e-09 1.8040307403136309 9.858e-09 1.8168588944542265 9.858999999999999e-09 1.8099096559725776 9.86e-09 1.7739682453378827 9.861e-09 1.833501126776031 9.862e-09 1.7541646851486878 9.863e-09 1.7497756895530856 9.864e-09 1.7098599479152283 9.865e-09 1.7352864210686358 9.866e-09 1.8416359879125896 9.867e-09 1.763117285873737 9.868e-09 1.8289764078088364 9.869e-09 1.747697604900625 9.87e-09 1.7986542513559738 9.871e-09 1.8336853487767553 9.871999999999999e-09 1.8285264087027853 9.873e-09 1.852808917754929 9.874e-09 1.7672194293176626 9.874999999999999e-09 1.8257064193606674 9.876e-09 1.8346560819692137 9.877e-09 1.7880866323324434 9.878e-09 1.662357861822071 9.879e-09 1.8698950858734769 9.88e-09 1.861458065001701 9.881e-09 1.858674503674052 9.882e-09 1.8373049509770505 9.883e-09 1.8386000192757892 9.884e-09 1.7514263574961686 9.885e-09 1.8206867719898954 9.886e-09 1.8584038607166664 9.887e-09 1.847194485657294 9.888e-09 1.847938501415939 9.889e-09 1.9479502804503253 9.89e-09 1.9012843630760796 9.890999999999999e-09 1.7358601990802018 9.892e-09 1.8593166386090825 9.893e-09 1.7823915327064066 9.893999999999999e-09 1.7520643523783053 9.895e-09 1.8740215639010096 9.896e-09 1.7559113215879238 9.897e-09 1.7682204168238635 9.898e-09 1.878320553907194 9.899e-09 1.8939121460741464 9.9e-09 1.7891616687673018 9.901e-09 1.7832535821917177 9.902e-09 1.824841538465414 9.903e-09 1.783236246173428 9.904e-09 1.9397303377119566 9.905e-09 1.82150716150913 9.906e-09 1.7256842615016368 9.906999999999999e-09 1.832737836126842 9.908e-09 1.7553233327716977 9.909e-09 1.773010271704996 9.909999999999999e-09 1.8545606737616835 9.911e-09 1.8174794636721607 9.912e-09 1.8242852071093192 9.912999999999999e-09 1.7460005307451114 9.914e-09 1.7672195696798767 9.915e-09 1.7303507874019084 9.916e-09 1.7336594163277017 9.917e-09 1.8083318717181467 9.918e-09 1.7520576139690145 9.919e-09 1.7668184454251348 9.92e-09 1.867067756497684 9.921e-09 1.7965869651490896 9.922e-09 1.783682487944142 9.923e-09 1.8387176844140236 9.924e-09 1.8895278305316987 9.925e-09 1.7894771291836957 9.925999999999999e-09 1.8334917379238713 9.927e-09 1.8242797491488663 9.928e-09 1.8621933205422097 9.928999999999999e-09 1.8402573839602139 9.93e-09 1.8083348275475262 9.931e-09 1.7939146840729387 9.932e-09 1.788308733535624 9.933e-09 1.7714990769651382 9.934e-09 1.728776535577953 9.935e-09 1.8486264663052963 9.936e-09 1.784592901298587 9.937e-09 1.772413346041693 9.938e-09 1.8611168465211199 9.939e-09 1.789663063326889 9.94e-09 1.827916337257925 9.941e-09 1.8651183144542938 9.942e-09 1.8240362860606314 9.943e-09 1.7773781548214609 9.944e-09 1.7755162659630688 9.944999999999999e-09 1.802243682459739 9.946e-09 1.849293760979562 9.947e-09 1.8357294485285844 9.947999999999999e-09 1.7700424086992992 9.949e-09 1.7897623296451923 9.95e-09 1.7986092383106504 9.951e-09 1.7526872212274398 9.952e-09 1.7364103655288836 9.953e-09 1.7920804391057568 9.954e-09 1.783541932568415 9.955e-09 1.7821697439519504 9.956e-09 1.7499606304228768 9.957e-09 1.8230484219390026 9.958e-09 1.8559652984359587 9.959e-09 1.8491069516226903 9.96e-09 1.7701435105641479 9.960999999999999e-09 1.7772110641952261 9.962e-09 1.7513263038751439 9.963e-09 1.7443874200449212 9.963999999999999e-09 1.7765706684520202 9.965e-09 1.7766190177870045 9.966e-09 1.7523982720725149 9.967e-09 1.7864605250327403 9.968e-09 1.7226914216030333 9.969e-09 1.7906761055747225 9.97e-09 1.8714950937576482 9.971e-09 1.9565265759183825 9.972e-09 1.7437627577298582 9.973e-09 1.691578097694377 9.974e-09 1.8147445991100655 9.975e-09 1.8335352987964153 9.976e-09 1.7334740557569304 9.977e-09 1.6928785787935854 9.978e-09 1.8097177199667862 9.979e-09 1.7959155626241003 9.979999999999999e-09 1.848495140629572 9.981e-09 1.806247775159348 9.982e-09 1.7747758162024014 9.982999999999999e-09 1.763617918014475 9.984e-09 1.8221672340287913 9.985e-09 1.8615900712372757 9.986e-09 1.7925317046241973 9.987e-09 1.8268960437352921 9.988e-09 1.7791013509120228 9.989e-09 1.7518636886063266 9.99e-09 1.7693966324318113 9.991e-09 1.7793820211199705 9.992e-09 1.8423811626481532 9.993e-09 1.766803015979411 9.994e-09 1.8129770522173967 9.995e-09 1.850865256869365 9.995999999999999e-09 1.6941336018697046 9.997e-09 1.7845603715917224 9.998e-09 1.837051856791997 9.998999999999999e-09 1.8430334367892482 1e-08 1.702563724331057 1.0001e-08 1.8187348970826613 1.0001999999999999e-08 1.8014934419928401 1.0003e-08 1.801568112833238 1.0004e-08 1.8568826213902299 1.0005e-08 1.7452303537282525 1.0006e-08 1.7594261764903774 1.0007e-08 1.8508153693036185 1.0008e-08 1.9002875704097566 1.0009e-08 1.7894090501452684 1.001e-08 1.7722611958730843 1.0011e-08 1.793396579857166 1.0012e-08 1.8050524943073987 1.0013e-08 1.853802064303281 1.0014e-08 1.8463030612358717 1.0014999999999999e-08 1.7795706509073592 1.0016e-08 1.8372407268059536 1.0017e-08 1.7613571987607948 1.0017999999999999e-08 1.8015519696484659 1.0019e-08 1.7837363194509173 1.002e-08 1.8024957819861733 1.0021e-08 1.7387881186628207 1.0022e-08 1.7842352255220273 1.0023e-08 1.7434824825838642 1.0024e-08 1.7677554722487487 1.0025e-08 1.7940765560783123 1.0026e-08 1.712952070844183 1.0027e-08 1.8680719565975685 1.0028e-08 1.7249687321487082 1.0029e-08 1.8773597298122722 1.003e-08 1.8336881239596803 1.0031e-08 1.7840212449856483 1.0032e-08 1.834342734931885 1.0033e-08 1.807885062082642 1.0033999999999999e-08 1.7487497248351 1.0035e-08 1.7000071726721535 1.0036e-08 1.7625157277249228 1.0036999999999999e-08 1.765322318689418 1.0038e-08 1.7292184736756302 1.0039e-08 1.7709074021176705 1.004e-08 1.7655966792098934 1.0041e-08 1.7753323058700339 1.0042e-08 1.8881881510890848 1.0043e-08 1.819061423910043 1.0044e-08 1.753588185201602 1.0045e-08 1.7602589719931137 1.0046e-08 1.7685934400018894 1.0047e-08 1.8207728862939352 1.0048e-08 1.8029274868077032 1.0049e-08 1.7753093621505682 1.0049999999999999e-08 1.731514750544388 1.0051e-08 1.8840051230760078 1.0052e-08 1.7901020369380964 1.0052999999999999e-08 1.7022995620111099 1.0054e-08 1.7284771827126564 1.0055e-08 1.735036142628986 1.0056e-08 1.8788729423660435 1.0057e-08 1.7029748646411718 1.0058e-08 1.762399839794326 1.0059e-08 1.7436587605109397 1.006e-08 1.8019880089907343 1.0061e-08 1.8326810128145656 1.0062e-08 1.7798362007796318 1.0063e-08 1.7576351185969432 1.0064e-08 1.8386027404669418 1.0065e-08 1.7741879726801344 1.0066e-08 1.7778846445429928 1.0067e-08 1.8196514540801285 1.0068e-08 1.8230171844421934 1.0068999999999999e-08 1.8051556606817811 1.007e-08 1.8749795013659347 1.0071e-08 1.8615322031449968 1.0071999999999999e-08 1.7840280354626914 1.0073e-08 1.777189168111677 1.0074e-08 1.7079561488511055 1.0075e-08 1.784701920403324 1.0076e-08 1.786144668094694 1.0077e-08 1.7080531419672655 1.0078e-08 1.7577843746054278 1.0079e-08 1.8073205262228227 1.008e-08 1.8640866080223597 1.0081e-08 1.8157256331009424 1.0082e-08 1.7886508286701552 1.0083e-08 1.8292137425297559 1.0084e-08 1.8695971341025237 1.0084999999999999e-08 1.9175918024486935 1.0086e-08 1.785289694919058 1.0087e-08 1.7590405799237134 1.0087999999999999e-08 1.7370071127966378 1.0089e-08 1.7722942148408516 1.009e-08 1.7197137528928865 1.0090999999999999e-08 1.7138516985611005 1.0092e-08 1.8735644053100013 1.0093e-08 1.798967834262516 1.0094e-08 1.8115357860602321 1.0095e-08 1.7718089951209497 1.0096e-08 1.8277571714944176 1.0097e-08 1.84209063542377 1.0098e-08 1.7342845869493604 1.0099e-08 1.7666709362182964 1.01e-08 1.855063639023712 1.0101e-08 1.7784761015959798 1.0102e-08 1.77165816622535 1.0103e-08 1.770524482323082 1.0103999999999999e-08 1.7874991562333007 1.0105e-08 1.847814759310481 1.0106e-08 1.8135925824621355 1.0106999999999999e-08 1.8463260709580984 1.0108e-08 1.7354753890964496 1.0109e-08 1.81854135725558 1.011e-08 1.8218839184648077 1.0111e-08 1.831558503785355 1.0112e-08 1.7957176887841815 1.0113e-08 1.8024046728847842 1.0114e-08 1.6965098626368051 1.0115e-08 1.7789437572584532 1.0116e-08 1.8056363833533953 1.0117e-08 1.7779176799958407 1.0118e-08 1.8295411782824538 1.0119e-08 1.7305974631743553 1.012e-08 1.8850839092920175 1.0121e-08 1.7599829272717944 1.0122e-08 1.8552285666775872 1.0122999999999999e-08 1.8736287733498582 1.0124e-08 1.7077634195404914 1.0125e-08 1.8370446998897918 1.0125999999999999e-08 1.7091030292432947 1.0127e-08 1.7894215446668043 1.0128e-08 1.7243503516145129 1.0129e-08 1.6367545708260902 1.013e-08 1.7791202665661856 1.0131e-08 1.8668963065349804 1.0132e-08 1.7878821287813167 1.0133e-08 1.7771154472363062 1.0134e-08 1.824193580193291 1.0135e-08 1.804737155495724 1.0136e-08 1.843281511384899 1.0137e-08 1.8360759724551285 1.0138e-08 1.7801186002349234 1.0138999999999999e-08 1.7942914749747318 1.014e-08 1.6819128772118896 1.0141e-08 1.7792563626182738 1.0141999999999999e-08 1.7349249309550723 1.0143e-08 1.7414027875277538 1.0144e-08 1.7367872343275617 1.0145e-08 1.8104890388321564 1.0146e-08 1.7032786586669086 1.0147e-08 1.8263169028550685 1.0148e-08 1.831186464470756 1.0149e-08 1.9385436486313359 1.015e-08 1.8716662159612287 1.0151e-08 1.795855683605004 1.0152e-08 1.7942642645410518 1.0153e-08 1.7968570730488282 1.0154e-08 1.8461528216585903 1.0155e-08 1.7820830126490315 1.0156e-08 1.7782232647496794 1.0157e-08 1.7937124332860395 1.0157999999999999e-08 1.731665253290354 1.0159e-08 1.7453263568497785 1.016e-08 1.8564076370482943 1.0160999999999999e-08 1.881956962002043 1.0162e-08 1.7981736099702463 1.0163e-08 1.7222446717387276 1.0164e-08 1.8508624301311714 1.0165e-08 1.7023464596990958 1.0166e-08 1.8293470025808147 1.0167e-08 1.7642936449433022 1.0168e-08 1.781387017973527 1.0169e-08 1.764406659280864 1.017e-08 1.881686502564673 1.0171e-08 1.843601322694163 1.0172e-08 1.8280009366974295 1.0173e-08 1.8095446786144587 1.0173999999999999e-08 1.8226643567292429 1.0175e-08 1.8132547195158417 1.0176e-08 1.7370910913847646 1.0176999999999999e-08 1.7899997683765951 1.0178e-08 1.718233492262132 1.0179e-08 1.7462214767326303 1.018e-08 1.7862785506348446 1.0181e-08 1.7873665782249533 1.0182e-08 1.8811666879570692 1.0183e-08 1.8423556343429237 1.0184e-08 1.7857358682513211 1.0185e-08 1.799299032303707 1.0186e-08 1.8210392985858255 1.0187e-08 1.8040361155557316 1.0188e-08 1.7332112331419687 1.0189e-08 1.8253948025742115 1.019e-08 1.76223448874775 1.0191e-08 1.7730103916697364 1.0192e-08 1.8046205148960517 1.0192999999999999e-08 1.8319963993669992 1.0194e-08 1.819373719410766 1.0195e-08 1.7800596508117694 1.0195999999999999e-08 1.8951245477294467 1.0197e-08 1.865918273174773 1.0198e-08 1.7679668830018935 1.0199e-08 1.7821840912751503 1.02e-08 1.7492179847415874 1.0201e-08 1.7603650137497893 1.0202e-08 1.7737805941971685 1.0203e-08 1.803311132920548 1.0204e-08 1.7925212173717004 1.0205e-08 1.779207087304916 1.0206e-08 1.7125027453725215 1.0207e-08 1.7148136070814755 1.0208e-08 1.7966827600052249 1.0208999999999999e-08 1.8598909104306438 1.021e-08 1.771400959863619 1.0211e-08 1.7347443550393906 1.0211999999999999e-08 1.8354068415771465 1.0213e-08 1.7220114005782667 1.0214e-08 1.7523626797303702 1.0214999999999999e-08 1.8077732875703116 1.0216e-08 1.7804545530477613 1.0217e-08 1.8117039346416268 1.0218e-08 1.8582751615669446 1.0219e-08 1.6970787910942462 1.022e-08 1.8482905883611804 1.0221e-08 1.7467728726153615 1.0222e-08 1.8683277694361007 1.0223e-08 1.817311300157517 1.0224e-08 1.8292918574580495 1.0225e-08 1.7701488424323744 1.0226e-08 1.6882738833669007 1.0227e-08 1.8066181008461875 1.0227999999999999e-08 1.7638841175726032 1.0229e-08 1.7843502710516164 1.023e-08 1.7308114089305562 1.0230999999999999e-08 1.8114148501718763 1.0232e-08 1.826686304098275 1.0233e-08 1.7726998317106273 1.0234e-08 1.7273093793103391 1.0235e-08 1.7302678043058526 1.0236e-08 1.8713096376242762 1.0237e-08 1.7714949009397047 1.0238e-08 1.8335465437057739 1.0239e-08 1.7418264296977146 1.024e-08 1.7592635916270634 1.0241e-08 1.8122903431123336 1.0242e-08 1.758988596637496 1.0243e-08 1.8438800028228535 1.0244e-08 1.7754829888048866 1.0245e-08 1.8851711713198909 1.0246e-08 1.8592505294837398 1.0246999999999999e-08 1.823774969689359 1.0248e-08 1.8141249355825744 1.0249e-08 1.7629789325950649 1.0249999999999999e-08 1.762704844999267 1.0251e-08 1.8449523576333606 1.0252e-08 1.9052705990345364 1.0253e-08 1.773744879237195 1.0254e-08 1.7707609535902256 1.0255e-08 1.8295302739675292 1.0256e-08 1.7792080340613066 1.0257e-08 1.8286371403162798 1.0258e-08 1.805667893424493 1.0259e-08 1.8099646124827393 1.026e-08 1.806161997226427 1.0261e-08 1.739156430205736 1.0262e-08 1.793285049304012 1.0262999999999999e-08 1.8481781954344263 1.0264e-08 1.7916861225311453 1.0265e-08 1.787435811843705 1.0265999999999999e-08 1.7540374848301152 1.0267e-08 1.7565537239338251 1.0268e-08 1.7929475373717239 1.0269e-08 1.8784901868912844 1.027e-08 1.8400728964214625 1.0271e-08 1.768791824025069 1.0272e-08 1.7996911817513814 1.0273e-08 1.8172165229281383 1.0274e-08 1.7391358181026488 1.0275e-08 1.8355826932958492 1.0276e-08 1.7435665336076602 1.0277e-08 1.7715354570988047 1.0278e-08 1.8685544337994282 1.0279e-08 1.7233340106166064 1.028e-08 1.7823569833995159 1.0281e-08 1.789624111131632 1.0281999999999999e-08 1.7366163813317208 1.0283e-08 1.8588878689300157 1.0284e-08 1.857173877596601 1.0284999999999999e-08 1.834599923040388 1.0286e-08 1.6631107617393974 1.0287e-08 1.794952567343602 1.0288e-08 1.7909106843599578 1.0289e-08 1.7881119717582383 1.029e-08 1.7647025714433713 1.0291e-08 1.7841590303918762 1.0292e-08 1.807461457499309 1.0293e-08 1.8567347499460165 1.0294e-08 1.780049284677635 1.0295e-08 1.7693863957335143 1.0296e-08 1.7761165496139788 1.0297e-08 1.7603756560180095 1.0297999999999999e-08 1.8718853994940354 1.0299e-08 1.7722162562723354 1.03e-08 1.7382122544843446 1.0300999999999999e-08 1.7481011948414409 1.0302e-08 1.8803449387488875 1.0303e-08 1.9041623555975882 1.0303999999999999e-08 1.932952310712835 1.0305e-08 1.8546093368353345 1.0306e-08 1.7698625827288812 1.0307e-08 1.8143347495685829 1.0308e-08 1.7424965113537647 1.0309e-08 1.6798791248927583 1.031e-08 1.8534788376557145 1.0311e-08 1.7841654082553544 1.0312e-08 1.8623724863575213 1.0313e-08 1.8886335974651887 1.0314e-08 1.828068263514266 1.0315e-08 1.7714276281660413 1.0316e-08 1.897613698513493 1.0316999999999999e-08 1.6781708180853685 1.0318e-08 1.8177358890593593 1.0319e-08 1.781623216411424 1.0319999999999999e-08 1.793997601367785 1.0321e-08 1.8236366200134824 1.0322e-08 1.8186223676097577 1.0323e-08 1.7998242157283342 1.0324e-08 1.877089528775951 1.0325e-08 1.8201965933075668 1.0326e-08 1.7676915621050961 1.0327e-08 1.797873965769762 1.0328e-08 1.8459597692976404 1.0329e-08 1.7741563951644632 1.033e-08 1.8790139458260937 1.0331e-08 1.807881571134759 1.0332e-08 1.7840298618449986 1.0333e-08 1.8271239449202494 1.0334e-08 1.7890173672674585 1.0335e-08 1.8212268817742205 1.0335999999999999e-08 1.8069079578202214 1.0337e-08 1.7854449414395157 1.0338e-08 1.8918753705987423 1.0338999999999999e-08 1.9183625849493446 1.034e-08 1.8214906190095264 1.0341e-08 1.7999685658911253 1.0342e-08 1.7701930144323101 1.0343e-08 1.8569130765291708 1.0344e-08 1.7897644106760693 1.0345e-08 1.7981675943724567 1.0346e-08 1.8084804185773922 1.0347e-08 1.8071340207314728 1.0348e-08 1.7714384693372207 1.0349e-08 1.8224065562769778 1.035e-08 1.7444386333831976 1.0351e-08 1.7808264356567376 1.0351999999999999e-08 1.7817792736882205 1.0353e-08 1.8365293249471994 1.0354e-08 1.7823622012793439 1.0354999999999999e-08 1.724731648023245 1.0356e-08 1.804464171875627 1.0357e-08 1.7928409823218363 1.0358e-08 1.8317860364326521 1.0359e-08 1.7395888291890143 1.036e-08 1.8509118341544988 1.0361e-08 1.8411235210679426 1.0362e-08 1.809244904093393 1.0363e-08 1.860131987079171 1.0364e-08 1.8134342387084945 1.0365e-08 1.754757401177457 1.0366e-08 1.7393054932761964 1.0367e-08 1.8650856899048944 1.0368e-08 1.8122749917313332 1.0369e-08 1.7990817577651128 1.037e-08 1.8061287251278775 1.0370999999999999e-08 1.710227684073683 1.0372e-08 1.8104275746182323 1.0373e-08 1.76890001399134 1.0373999999999999e-08 1.795956039257026 1.0375e-08 1.8182749938174445 1.0376e-08 1.8081567020897147 1.0377e-08 1.6852019392820066 1.0378e-08 1.8349804709875237 1.0379e-08 1.8940875512097133 1.038e-08 1.8551099230579353 1.0381e-08 1.7984918124927094 1.0382e-08 1.8697344541370486 1.0383e-08 1.7979295134533673 1.0384e-08 1.7252719865025616 1.0385e-08 1.7044301916721336 1.0386e-08 1.7944175605961665 1.0386999999999999e-08 1.7697458236936179 1.0388e-08 1.688560148849556 1.0389e-08 1.8036567779593617 1.0389999999999999e-08 1.8332952092204353 1.0391e-08 1.8014388768204022 1.0392e-08 1.835145018436883 1.0392999999999999e-08 1.6880686555657634 1.0394e-08 1.9211334642243736 1.0395e-08 1.7770124929943125 1.0396e-08 1.792550133974717 1.0397e-08 1.9520757321804845 1.0398e-08 1.7630889807198937 1.0399e-08 1.8429865077106093 1.04e-08 1.7180002048518968 1.0401e-08 1.8044983371266525 1.0402e-08 1.7960991700867248 1.0403e-08 1.8558622424319053 1.0404e-08 1.7679558019913861 1.0405e-08 1.7254059809275206 1.0405999999999999e-08 1.8230399107710926 1.0407e-08 1.7536073481693708 1.0408e-08 1.8523011883373497 1.0408999999999999e-08 1.797702198601641 1.041e-08 1.8460995615836753 1.0411e-08 1.8289357544304938 1.0412e-08 1.8771687295515889 1.0413e-08 1.8193137727081803 1.0414e-08 1.8805559145669741 1.0415e-08 1.7591228452123622 1.0416e-08 1.8139792065495515 1.0417e-08 1.7595583176427425 1.0418e-08 1.7464756207270822 1.0419e-08 1.7617668518433196 1.042e-08 1.8201779890019294 1.0421e-08 1.7712470135398 1.0422e-08 1.7261812465402717 1.0423e-08 1.7885533495530084 1.0424e-08 1.7513695584768691 1.0424999999999999e-08 1.8468947567164373 1.0426e-08 1.807129648946841 1.0427e-08 1.8061448984291961 1.0427999999999999e-08 1.7250623402641438 1.0429e-08 1.7617793705531537 1.043e-08 1.7429172676635638 1.0431e-08 1.74299621050939 1.0432e-08 1.8611505332531517 1.0433e-08 1.929395204974097 1.0434e-08 1.867088266732249 1.0435e-08 1.7709146264260431 1.0436e-08 1.8035912513639512 1.0437e-08 1.87214783910005 1.0438e-08 1.8150478061057091 1.0439e-08 1.7539685726208338 1.044e-08 1.7747129441537088 1.0440999999999999e-08 1.8275164697135369 1.0442e-08 1.8220473237524013 1.0443e-08 1.7662776092115375 1.0443999999999999e-08 1.7518288325975353 1.0445e-08 1.7026656874263222 1.0446e-08 1.7850724530342958 1.0447e-08 1.7857820754756242 1.0448e-08 1.8014428207651432 1.0449e-08 1.8519342957663267 1.045e-08 1.8572634282318041 1.0451e-08 1.8022517072405546 1.0452e-08 1.8202175154766393 1.0453e-08 1.716956511130779 1.0454e-08 1.7823729131715924 1.0455e-08 1.7701331337655417 1.0456e-08 1.7566586526515935 1.0457e-08 1.8566996723559586 1.0458e-08 1.7420391334348848 1.0459e-08 1.789120603848043 1.0459999999999999e-08 1.8802511002032036 1.0461e-08 1.798812181783335 1.0462e-08 1.7308640171046386 1.0462999999999999e-08 1.8180812694220485 1.0464e-08 1.8664338160349605 1.0465e-08 1.696077884832426 1.0466e-08 1.874236175854715 1.0467e-08 1.8141950673306435 1.0468e-08 1.6680109717096538 1.0469e-08 1.792850299785569 1.047e-08 1.7953794914116015 1.0471e-08 1.8914639003983629 1.0472e-08 1.7273450596528628 1.0473e-08 1.883480611651156 1.0474e-08 1.7456054952064501 1.0475e-08 1.7881267742982445 1.0475999999999999e-08 1.7569975541456757 1.0477e-08 1.809597305509426 1.0478e-08 1.793124402480136 1.0478999999999999e-08 1.9209542504110226 1.048e-08 1.864790740754433 1.0481e-08 1.8063555692505833 1.0481999999999999e-08 1.836478624454562 1.0483e-08 1.8824480839662905 1.0484e-08 1.851287205435065 1.0485e-08 1.8749362969774896 1.0486e-08 1.8365839948850273 1.0487e-08 1.7930011040154787 1.0488e-08 1.7726069277940903 1.0489e-08 1.7530385306506158 1.049e-08 1.8341130048263463 1.0491e-08 1.76478429224506 1.0492e-08 1.8182690495156257 1.0493e-08 1.8634662799279753 1.0494e-08 1.81689394481513 1.0494999999999999e-08 1.728384595150553 1.0496e-08 1.8727847530106352 1.0497e-08 1.8369167754634081 1.0497999999999999e-08 1.8761781812790086 1.0499e-08 1.8102005653163182 1.05e-08 1.7588218233826551 1.0501e-08 1.7710522475950967 1.0502e-08 1.7480786791022476 1.0503e-08 1.8703492877702694 1.0504e-08 1.835565040341024 1.0505e-08 1.7756155076827818 1.0506e-08 1.7754803590322585 1.0507e-08 1.7885143538920116 1.0508e-08 1.7571396600070084 1.0509e-08 1.6914640476026226 1.051e-08 1.8583282400832535 1.0510999999999999e-08 1.8194808267535652 1.0512e-08 1.7651446931997476 1.0513e-08 1.7545209896049816 1.0513999999999999e-08 1.7201481843979498 1.0515e-08 1.7929350706678455 1.0516e-08 1.790570034895285 1.0516999999999999e-08 1.8683629119467917 1.0518e-08 1.8035705616166644 1.0519e-08 1.896246399864928 1.052e-08 1.8390801622974016 1.0521e-08 1.6907684950866193 1.0522e-08 1.8554454877947086 1.0523e-08 1.9132765050951077 1.0524e-08 1.7731909895540763 1.0525e-08 1.845499867009042 1.0526e-08 1.8423006980098622 1.0527e-08 1.7510525181124685 1.0528e-08 1.7873991005302632 1.0529e-08 1.7870656844386712 1.0529999999999999e-08 1.8156215594689185 1.0531e-08 1.8138720081387691 1.0532e-08 1.7692929193116844 1.0532999999999999e-08 1.659558135849146 1.0534e-08 1.884908503766503 1.0535e-08 1.9554739138247414 1.0536e-08 1.7684071804793084 1.0537e-08 1.79006456914831 1.0538e-08 1.811270349928164 1.0539e-08 1.8244897611822986 1.054e-08 1.8601070499958308 1.0541e-08 1.8077114364680782 1.0542e-08 1.7469583967961937 1.0543e-08 1.7802091375253575 1.0544e-08 1.9234067265979824 1.0545e-08 1.8575021612697091 1.0546e-08 1.8948498796378208 1.0547e-08 1.7430875978014118 1.0548e-08 1.7905560937648424 1.0548999999999999e-08 1.8637956294194225 1.055e-08 1.9221581026952415 1.0551e-08 1.8557259736369822 1.0551999999999999e-08 1.7685890565463236 1.0553e-08 1.8510030338453358 1.0554e-08 1.8395477479070708 1.0555e-08 1.8100049518659294 1.0556e-08 1.79609471111501 1.0557e-08 1.7632353756988346 1.0558e-08 1.7906740984276732 1.0559e-08 1.7757929214781467 1.056e-08 1.8206815955313798 1.0561e-08 1.8375599433586245 1.0562e-08 1.7473787285116078 1.0563e-08 1.7857895044879302 1.0564e-08 1.7410748242010625 1.0564999999999999e-08 1.7371422236086849 1.0566e-08 1.8721810624530029 1.0567e-08 1.844310656614871 1.0567999999999999e-08 1.7904952112518129 1.0569e-08 1.6983355498208101 1.057e-08 1.6992412462819935 1.0570999999999999e-08 1.7441870420704517 1.0572e-08 1.7380164864171923 1.0573e-08 1.7708215143762858 1.0574e-08 1.7995937317851882 1.0575e-08 1.7986678443930009 1.0576e-08 1.8607467283762553 1.0577e-08 1.798153348726951 1.0578e-08 1.8112095137757098 1.0579e-08 1.7564895036390658 1.058e-08 1.7302015558677544 1.0581e-08 1.7949698466404076 1.0582e-08 1.786873976841733 1.0583e-08 1.8031823816079346 1.0583999999999999e-08 1.7339510890590173 1.0585e-08 1.8086832444506247 1.0586e-08 1.810752980272205 1.0586999999999999e-08 1.821670964656974 1.0588e-08 1.7209786703709995 1.0589e-08 1.8626392068264945 1.059e-08 1.765870908703166 1.0591e-08 1.7907434689056207 1.0592e-08 1.7909255231398198 1.0593e-08 1.768014178192304 1.0594e-08 1.8468950608562873 1.0595e-08 1.844738614496056 1.0596e-08 1.8595208391241662 1.0597e-08 1.7999393666624124 1.0598e-08 1.7926712914656047 1.0599e-08 1.7743764734846115 1.0599999999999999e-08 1.8798076253716545 1.0601e-08 1.7628082122005468 1.0602e-08 1.7649906771747905 1.0602999999999999e-08 1.9160584014726822 1.0604e-08 1.8036691894619652 1.0605e-08 1.883921808205743 1.0605999999999999e-08 1.7932491923080016 1.0607e-08 1.8214810050696242 1.0608e-08 1.845851317035023 1.0609e-08 1.8949926430688848 1.061e-08 1.8332597110591862 1.0611e-08 1.7123773497975592 1.0612e-08 1.7823141677065375 1.0613e-08 1.8673755285729436 1.0614e-08 1.7696249188259203 1.0615e-08 1.7864127682965099 1.0616e-08 1.7910263934021133 1.0617e-08 1.794933627707714 1.0618e-08 1.7744226508748062 1.0618999999999999e-08 1.7875151181501499 1.062e-08 1.888754968057615 1.0621e-08 1.8390898798172892 1.0621999999999999e-08 1.8371385622509349 1.0623e-08 1.827726219832356 1.0624e-08 1.685774651333226 1.0625e-08 1.7935143664401751 1.0626e-08 1.7923862027379591 1.0627e-08 1.7490612298000618 1.0628e-08 1.771223772755807 1.0629e-08 1.840645576046822 1.063e-08 1.8021320234249951 1.0631e-08 1.7748449678047544 1.0632e-08 1.8149771012124836 1.0633e-08 1.8276501684662279 1.0634e-08 1.7886536534581217 1.0635e-08 1.8430335339116533 1.0636e-08 1.840725851870657 1.0637e-08 1.689027411212292 1.0637999999999999e-08 1.732300406624331 1.0639e-08 1.7963950232478876 1.064e-08 1.8047801632405969 1.0640999999999999e-08 1.818976727310065 1.0642e-08 1.801744960349253 1.0643e-08 1.780788523065437 1.0644e-08 1.8123264920496454 1.0645e-08 1.8837377856224047 1.0646e-08 1.8292020546777106 1.0647e-08 1.6313648357722201 1.0648e-08 1.8131173516187162 1.0649e-08 1.881616686107524 1.065e-08 1.6974937073208238 1.0651e-08 1.842590661344279 1.0652e-08 1.7946279634099593 1.0653e-08 1.7720631451980509 1.0653999999999999e-08 1.8177372739559625 1.0655e-08 1.7617860739738016 1.0656e-08 1.8450063810858781 1.0656999999999999e-08 1.7168564964036288 1.0658e-08 1.8331104997756047 1.0659e-08 1.915215349463136 1.0659999999999999e-08 1.7946029542939197 1.0661e-08 1.8907635330704264 1.0662e-08 1.743540757467168 1.0663e-08 1.7025025511100622 1.0664e-08 1.802659301948027 1.0665e-08 1.7970846635202349 1.0666e-08 1.7845784380573269 1.0667e-08 1.828043894362415 1.0668e-08 1.7891713677158727 1.0669e-08 1.7496930741115972 1.067e-08 1.8215073126323562 1.0671e-08 1.814823346344592 1.0672e-08 1.848097169285041 1.0672999999999999e-08 1.8175913164706452 1.0674e-08 1.743578676552058 1.0675e-08 1.761408496836168 1.0675999999999999e-08 1.7139974087616774 1.0677e-08 1.9001571203464491 1.0678e-08 1.8174092582771055 1.0679e-08 1.8932777333625617 1.068e-08 1.770073499923105 1.0681e-08 1.777312308123524 1.0682e-08 1.7421445726514821 1.0683e-08 1.8916762219630003 1.0684e-08 1.819621421288677 1.0685e-08 1.8010988865896576 1.0686e-08 1.7210263672689952 1.0687e-08 1.8635420360685533 1.0688e-08 1.8242852221789554 1.0688999999999999e-08 1.8332317709038475 1.069e-08 1.7278623080161357 1.0691e-08 1.8304645981063428 1.0691999999999999e-08 1.8121204448825916 1.0693e-08 1.791482005268709 1.0694e-08 1.895698187025316 1.0694999999999999e-08 1.7492890364511344 1.0696e-08 1.803891533944238 1.0697e-08 1.7561883256537736 1.0698e-08 1.76391730125245 1.0699e-08 1.7838260962945245 1.07e-08 1.7515343477985672 1.0701e-08 1.7820167540018907 1.0702e-08 1.786966976378495 1.0703e-08 1.7979022564706764 1.0704e-08 1.7888486824362275 1.0705e-08 1.8061685931827636 1.0706e-08 1.7334138068992944 1.0707e-08 1.8264073535060328 1.0707999999999999e-08 1.816462499474552 1.0709e-08 1.8405625322259929 1.071e-08 1.761594958117171 1.0710999999999999e-08 1.853440431058471 1.0712e-08 1.8256839008812622 1.0713e-08 1.872205816835688 1.0714e-08 1.7949724563238687 1.0715e-08 1.7169411643608528 1.0716e-08 1.8195042338154273 1.0717e-08 1.7721054801681817 1.0718e-08 1.6912797655725145 1.0719e-08 1.8839510791364351 1.072e-08 1.7939447033791893 1.0721e-08 1.8023766209737053 1.0722e-08 1.8291510058316955 1.0723e-08 1.791512600975553 1.0724e-08 1.7860604803061282 1.0725e-08 1.8284810452273317 1.0726e-08 1.7109428702725478 1.0726999999999999e-08 1.7869954125055154 1.0728e-08 1.7523238532133272 1.0729e-08 1.9040889122182838 1.0729999999999999e-08 1.8566959645964156 1.0731e-08 1.7375610487888105 1.0732e-08 1.7835093306931002 1.0733e-08 1.8512319090069855 1.0734e-08 1.8102032202757687 1.0735e-08 1.869826409991383 1.0736e-08 1.8137324833116488 1.0737e-08 1.806843411341406 1.0738e-08 1.8508360658519836 1.0739e-08 1.868965596033485 1.074e-08 1.795093914208869 1.0741e-08 1.7940857027696269 1.0742e-08 1.85247149716367 1.0742999999999999e-08 1.8308717598267457 1.0744e-08 1.773341764014584 1.0745e-08 1.8792310059314201 1.0745999999999999e-08 1.7019892185676704 1.0747e-08 1.8812227168019477 1.0748e-08 1.826284078030619 1.0749e-08 1.7755939002040766 1.075e-08 1.8102667306266689 1.0751e-08 1.78537973092561 1.0752e-08 1.7292827806020852 1.0753e-08 1.9386641864651466 1.0754e-08 1.8160562621607585 1.0755e-08 1.7965477448174514 1.0756e-08 1.8054807514896387 1.0757e-08 1.8518249635784203 1.0758e-08 1.7752516908269131 1.0759e-08 1.7763275507206526 1.076e-08 1.7737185414658696 1.0761e-08 1.7314175685089876 1.0761999999999999e-08 1.7662281469931536 1.0763e-08 1.7847761256133596 1.0764e-08 1.6608092489721842 1.0764999999999999e-08 1.8690190832434885 1.0766e-08 1.758106176652655 1.0767e-08 1.81149706331498 1.0768e-08 1.762116640450551 1.0769e-08 1.7531371336812485 1.077e-08 1.8238261988501685 1.0771e-08 1.764446562198836 1.0772e-08 1.7803025541879365 1.0773e-08 1.7790198802956274 1.0774e-08 1.7979462570970575 1.0775e-08 1.6870444975929757 1.0776e-08 1.8020396697606698 1.0777e-08 1.756902164504412 1.0777999999999999e-08 1.8577173116751444 1.0779e-08 1.8171610192935592 1.078e-08 1.8004263645366727 1.0780999999999999e-08 1.80009945776348 1.0782e-08 1.8130602873448391 1.0783e-08 1.8211116700756642 1.0783999999999999e-08 1.7211539454262827 1.0785e-08 1.7696130885145032 1.0786e-08 1.765260214299246 1.0787e-08 1.7979345960102915 1.0788e-08 1.9160117623501896 1.0789e-08 1.7301913099514283 1.079e-08 1.836723926696087 1.0791e-08 1.846634909330983 1.0792e-08 1.8620300574630333 1.0793e-08 1.828773680843584 1.0794e-08 1.8489153723119276 1.0795e-08 1.751596469542172 1.0796e-08 1.7804170972542919 1.0796999999999999e-08 1.8634833493621745 1.0798e-08 1.7881580495674925 1.0799e-08 1.8011757870672795 1.0799999999999999e-08 1.7379127487491186 1.0801e-08 1.858259852722742 1.0802e-08 1.6437790112343083 1.0803e-08 1.8665100163652533 1.0804e-08 1.83304452961211 1.0805e-08 1.842006985259728 1.0806e-08 1.8159952989956851 1.0807e-08 1.768969894424302 1.0808e-08 1.8527548215638936 1.0809e-08 1.8532085371745946 1.081e-08 1.7606290076112552 1.0811e-08 1.7759125578151629 1.0812e-08 1.7984743029275292 1.0813e-08 1.8301332016550043 1.0814e-08 1.7840889903950221 1.0815e-08 1.7923285645404807 1.0815999999999999e-08 1.7978844325428227 1.0817e-08 1.8121643677495258 1.0818e-08 1.8063814477051134 1.0818999999999999e-08 1.8165805189313373 1.082e-08 1.7836972079691975 1.0821e-08 1.6171823257243636 1.0822e-08 1.7912993868048401 1.0823e-08 1.8206229111321781 1.0824e-08 1.799002568270527 1.0825e-08 1.7923723195519095 1.0826e-08 1.728615831948201 1.0827e-08 1.8514632406649623 1.0828e-08 1.828461361676545 1.0829e-08 1.760656668383707 1.083e-08 1.8349416136410257 1.0831e-08 1.814815045750584 1.0831999999999999e-08 1.7673894362788962 1.0833e-08 1.7833801579012072 1.0834e-08 1.8287125784911091 1.0834999999999999e-08 1.7882693940014607 1.0836e-08 1.7457486997682965 1.0837e-08 1.8562614773528354 1.0838e-08 1.8194674854368988 1.0839e-08 1.8242127739047282 1.084e-08 1.751131378431038 1.0841e-08 1.8618258000504149 1.0842e-08 1.7358713556334957 1.0843e-08 1.7688158779824237 1.0844e-08 1.8401563051318264 1.0845e-08 1.8054916329713055 1.0846e-08 1.7257484022252632 1.0847e-08 1.744492102896096 1.0848e-08 1.752348740535673 1.0849e-08 1.7705017608362654 1.085e-08 1.856069728761761 1.0850999999999999e-08 1.8603770853686326 1.0852e-08 1.7748146808426941 1.0853e-08 1.776520117478706 1.0853999999999999e-08 1.7963234021202297 1.0855e-08 1.752905820630863 1.0856e-08 1.7539857072519045 1.0857e-08 1.8062930521836522 1.0858e-08 1.75453804705189 1.0859e-08 1.712530897667509 1.086e-08 1.8630090743909178 1.0861e-08 1.8481606415805236 1.0862e-08 1.8034247742199274 1.0863e-08 1.7773826744577064 1.0864e-08 1.7870115265659898 1.0865e-08 1.7376155068150498 1.0866e-08 1.794945933698082 1.0866999999999999e-08 1.7968019650638296 1.0868e-08 1.8930011161432767 1.0869e-08 1.8049828226860278 1.0869999999999999e-08 1.8000192180210601 1.0871e-08 1.8795623782274296 1.0872e-08 1.775689032119128 1.0872999999999999e-08 1.7457115826563658 1.0874e-08 1.784746989835775 1.0875e-08 1.8516417588175758 1.0876e-08 1.8632704496427681 1.0877e-08 1.757367393587013 1.0878e-08 1.8092636917377776 1.0879e-08 1.7679441192768397 1.088e-08 1.8169419918050673 1.0881e-08 1.7895709390672485 1.0882e-08 1.6884578494151894 1.0883e-08 1.7949552210886026 1.0884e-08 1.7763801460366377 1.0885e-08 1.6994408357071358 1.0885999999999999e-08 1.822292154845031 1.0887e-08 1.8711184152768305 1.0888e-08 1.7837256729877802 1.0888999999999999e-08 1.8423634476925979 1.089e-08 1.8332000910914137 1.0891e-08 1.8770125923332657 1.0892e-08 1.80869513719896 1.0893e-08 1.7643666846475041 1.0894e-08 1.82057937312807 1.0895e-08 1.7693805214615022 1.0896e-08 1.7078581483636561 1.0897e-08 1.9084095018868237 1.0898e-08 1.875667468251025 1.0899e-08 1.7560667921248805 1.09e-08 1.7584015074596264 1.0901e-08 1.7983098182868809 1.0901999999999999e-08 1.7221578779882045 1.0903e-08 1.7877913087816255 1.0904e-08 1.725700505364434 1.0904999999999999e-08 1.7930167234486132 1.0906e-08 1.706350324731635 1.0907e-08 1.7191823239673414 1.0907999999999999e-08 1.796874003503382 1.0909e-08 1.73077960187708 1.091e-08 1.7709004557088712 1.0911e-08 1.8541061880126655 1.0912e-08 1.8147405000062946 1.0913e-08 1.990990332023935 1.0914e-08 1.7725310871015938 1.0915e-08 1.834926179842021 1.0916e-08 1.780255200316097 1.0917e-08 1.8043476376909795 1.0918e-08 1.8292529847237669 1.0919e-08 1.7701265157377517 1.092e-08 1.7557420084775641 1.0920999999999999e-08 1.6758829391235457 1.0922e-08 1.8248164087659609 1.0923e-08 1.8183415021486788 1.0923999999999999e-08 1.84800276146826 1.0925e-08 1.7481555200740428 1.0926e-08 1.8042271781680734 1.0927e-08 1.7876283639277353 1.0928e-08 1.8228621917381285 1.0929e-08 1.7622061955233386 1.093e-08 1.7940504324889281 1.0931e-08 1.8590169626967994 1.0932e-08 1.8121438580703104 1.0933e-08 1.655124003328768 1.0934e-08 1.7681513750829574 1.0935e-08 1.7185561379013137 1.0936e-08 1.866581578607526 1.0937e-08 1.780151434571694 1.0938e-08 1.7145422689584744 1.0939e-08 1.7574132329947088 1.0939999999999999e-08 1.8112237850745938 1.0941e-08 1.8268909005272933 1.0942e-08 1.9380717526502886 1.0942999999999999e-08 1.8835595473945665 1.0944e-08 1.7544823434487462 1.0945e-08 1.7892651541571294 1.0946e-08 1.8087402700696236 1.0947e-08 1.8494521961502068 1.0948e-08 1.802027649145617 1.0949e-08 1.765137862097608 1.095e-08 1.7565379972829591 1.0951e-08 1.8037022394393774 1.0952e-08 1.825111301904003 1.0953e-08 1.8059906965278025 1.0954e-08 1.7859310594638884 1.0955e-08 1.8516180485521567 1.0955999999999999e-08 1.8602632396200216 1.0957e-08 1.7772970863043718 1.0958e-08 1.8724463210619942 1.0958999999999999e-08 1.7963909090395596 1.096e-08 1.7240571115564176 1.0961e-08 1.714145515661337 1.0961999999999999e-08 1.9149516774295474 1.0963e-08 1.7340583253377526 1.0964e-08 1.85684865706767 1.0965e-08 1.7644790305262745 1.0966e-08 1.8065296699987947 1.0967e-08 1.702608238066981 1.0968e-08 1.8629544847188835 1.0969e-08 1.7825732427385808 1.097e-08 1.7608549017135613 1.0971e-08 1.8258454892234062 1.0972e-08 1.827863971294465 1.0973e-08 1.7614165896882366 1.0974e-08 1.7777912784631724 1.0974999999999999e-08 1.7627411699771034 1.0976e-08 1.8075956936289543 1.0977e-08 1.6003697236546297 1.0977999999999999e-08 1.830488031260288 1.0979e-08 1.7025111595980111 1.098e-08 1.8786544071640685 1.0981e-08 1.8504916486389464 1.0982e-08 1.899926261727897 1.0983e-08 1.810035576416078 1.0984e-08 1.7671316667364927 1.0985e-08 1.7941040666921562 1.0986e-08 1.8911082125584233 1.0987e-08 1.7714795773376903 1.0988e-08 1.7458884692242707 1.0989e-08 1.7649592512700234 1.099e-08 1.7103212633612008 1.0990999999999999e-08 1.8366103919484453 1.0992e-08 1.8379103649414128 1.0993e-08 1.8058296719686795 1.0993999999999999e-08 1.7857576077700352 1.0995e-08 1.7469843704528243 1.0996e-08 1.7944368290960577 1.0996999999999999e-08 1.8585568048443255 1.0998e-08 1.799492806103594 1.0999e-08 1.87088240560064 1.1e-08 1.6894703520206507 1.1001e-08 1.7768185218291699 1.1002e-08 1.8291692760540597 1.1003e-08 1.7983456387374483 1.1004e-08 1.8590737604635779 1.1005e-08 1.8581498404365235 1.1006e-08 1.7675213766913869 1.1007e-08 1.7869575143960614 1.1008e-08 1.7813902021320243 1.1009e-08 1.7218835561033603 1.1009999999999999e-08 1.8547687215980138 1.1011e-08 1.8329706535542793 1.1012e-08 1.8922240864878042 1.1012999999999999e-08 1.7327410040343993 1.1014e-08 1.8334587966835558 1.1015e-08 1.747489869974814 1.1016e-08 1.7798059192781066 1.1017e-08 1.7890280440424833 1.1018e-08 1.79405693258972 1.1019e-08 1.908720985986202 1.102e-08 1.8716838955491377 1.1021e-08 1.8466798089618517 1.1022e-08 1.8335265242329273 1.1023e-08 1.7852773396609685 1.1024e-08 1.7385996103022072 1.1025e-08 1.7816930874922488 1.1026e-08 1.7594700312115057 1.1027e-08 1.811268627696557 1.1028e-08 1.799947207102361 1.1028999999999999e-08 1.8467756423867145 1.103e-08 1.8982997039079932 1.1031e-08 1.85440112030669 1.1031999999999999e-08 1.8301520617303348 1.1033e-08 1.8253174210580423 1.1034e-08 1.7466552330703795 1.1035e-08 1.712396219931362 1.1036e-08 1.764524327375644 1.1037e-08 1.7696244271876493 1.1038e-08 1.7333812706517602 1.1039e-08 1.771296285235275 1.104e-08 1.8976222006218577 1.1041e-08 1.7419925663488451 1.1042e-08 1.8346030844995016 1.1043e-08 1.8488855666005026 1.1044e-08 1.776171821723931 1.1044999999999999e-08 1.7258902905324052 1.1046e-08 1.7952357978623839 1.1047e-08 1.7636078554508352 1.1047999999999999e-08 1.7625195870284696 1.1049e-08 1.8275513480994774 1.105e-08 1.8130574730071796 1.1050999999999999e-08 1.7690192913880436 1.1052e-08 1.8002620315806026 1.1053e-08 1.851998991898205 1.1054e-08 1.7669960889533078 1.1055e-08 1.7810037300770707 1.1056e-08 1.8261244619856385 1.1057e-08 1.8192091974215265 1.1058e-08 1.744225360214286 1.1059e-08 1.908980340213487 1.106e-08 1.837445699781906 1.1061e-08 1.851364091225863 1.1062e-08 1.765509422541835 1.1063e-08 1.8252400234488206 1.1063999999999999e-08 1.8229860106773041 1.1065e-08 1.7669692296846264 1.1066e-08 1.795656234957102 1.1066999999999999e-08 1.8674690848192823 1.1068e-08 1.8221858423272856 1.1069e-08 1.7958814533600895 1.107e-08 1.8222434877342026 1.1071e-08 1.8020661484456386 1.1072e-08 1.800144062879231 1.1073e-08 1.7779282488969679 1.1074e-08 1.821446542407379 1.1075e-08 1.832799766344057 1.1076e-08 1.7725750665225557 1.1077e-08 1.8330157245388048 1.1078e-08 1.9195071224119866 1.1079e-08 1.821704814395313 1.1079999999999999e-08 1.786744924403858 1.1081e-08 1.854103154395474 1.1082e-08 1.8203537037199693 1.1082999999999999e-08 1.9184306430561158 1.1084e-08 1.8182989414070778 1.1085e-08 1.8354146870329033 1.1085999999999999e-08 1.770470066509263 1.1087e-08 1.802804855200735 1.1088e-08 1.8503912481998628 1.1089e-08 1.8295255941646063 1.109e-08 1.7419168055183452 1.1091e-08 1.781998473565828 1.1092e-08 1.7879580178112282 1.1093e-08 1.784080563494114 1.1094e-08 1.880458757395414 1.1095e-08 1.6781751558075193 1.1096e-08 1.7815596163693066 1.1097e-08 1.7152082118983232 1.1098e-08 1.870094078170247 1.1098999999999999e-08 1.7847035826193536 1.11e-08 1.7929995205443652 1.1101e-08 1.8220214465976985 1.1101999999999999e-08 1.8655989187535489 1.1103e-08 1.7208727152371492 1.1104e-08 1.7847742563118285 1.1105e-08 1.854038279704605 1.1106e-08 1.785255524650158 1.1107e-08 1.806487581402948 1.1108e-08 1.647311172035894 1.1109e-08 1.8255755107340645 1.111e-08 1.6810909076135632 1.1111e-08 1.8669501007361842 1.1112e-08 1.7969881141384103 1.1113e-08 1.7207976069325897 1.1114e-08 1.8451072881040438 1.1115e-08 1.7859254299927234 1.1116e-08 1.8317813409458485 1.1117e-08 1.7845434956417907 1.1117999999999999e-08 1.8250520964210772 1.1119e-08 1.7993001999304687 1.112e-08 1.8377072482764996 1.1120999999999999e-08 1.78016007787975 1.1122e-08 1.8038616213774672 1.1123e-08 1.7546794814061242 1.1124e-08 1.754652777002696 1.1125e-08 1.7797685465354505 1.1126e-08 1.807609702402933 1.1127e-08 1.7997533904485634 1.1128e-08 1.7847492935163205 1.1129e-08 1.8714490941642261 1.113e-08 1.741692093673294 1.1131e-08 1.7830938437763268 1.1132e-08 1.7918100074517676 1.1133e-08 1.804763792413808 1.1133999999999999e-08 1.8184283512056518 1.1135e-08 1.8122126856407643 1.1136e-08 1.720918871841962 1.1136999999999999e-08 1.7336184067404394 1.1138e-08 1.732177431014606 1.1139e-08 1.7918794439485104 1.1139999999999999e-08 1.7687794807794956 1.1141e-08 1.7149508351744571 1.1142e-08 1.8156084940942707 1.1143e-08 1.839336158070743 1.1144e-08 1.7873036315525668 1.1145e-08 1.908051593538677 1.1146e-08 1.9092405634921796 1.1147e-08 1.7860576454370634 1.1148e-08 1.8380718575550912 1.1149e-08 1.786311914100863 1.115e-08 1.8414291101995077 1.1151e-08 1.8591298636763578 1.1152e-08 1.8031166340026108 1.1152999999999999e-08 1.7673534218605862 1.1154e-08 1.852382159472158 1.1155e-08 1.804578065074582 1.1155999999999999e-08 1.7887862636631402 1.1157e-08 1.809100410721053 1.1158e-08 1.9425806813835873 1.1159e-08 1.789521149330583 1.116e-08 1.8606354235643665 1.1161e-08 1.8011706797672635 1.1162e-08 1.7602316686421071 1.1163e-08 1.7920627144878032 1.1164e-08 1.719156222368858 1.1165e-08 1.8395938037119122 1.1166e-08 1.8688088078472918 1.1167e-08 1.834019596172015 1.1168e-08 1.8475329089471573 1.1168999999999999e-08 1.8018987697011453 1.117e-08 1.753398909110327 1.1171e-08 1.7079315066427403 1.1171999999999999e-08 1.8031024872288752 1.1173e-08 1.7609900097362055 1.1174e-08 1.7637742707676731 1.1174999999999999e-08 1.7576607955746781 1.1176e-08 1.7821454716273484 1.1177e-08 1.8256383700627539 1.1178e-08 1.7675381195088768 1.1179e-08 1.7327778666481986 1.118e-08 1.7925451577186349 1.1181e-08 1.885268189172339 1.1182e-08 1.808651975254938 1.1183e-08 1.7666886736863383 1.1184e-08 1.774792783603405 1.1185e-08 1.906324798854753 1.1186e-08 1.8425870344026083 1.1187e-08 1.6834774047396426 1.1187999999999999e-08 1.7703625849924165 1.1189e-08 1.8503965909492432 1.119e-08 1.8067860499119033 1.1190999999999999e-08 1.8366939526596244 1.1192e-08 1.784841133895639 1.1193e-08 1.8110740605374225 1.1194e-08 1.733062710687507 1.1195e-08 1.7742447552552145 1.1196e-08 1.7289295694846127 1.1197e-08 1.8282577079951314 1.1198e-08 1.712993006596175 1.1199e-08 1.7971553709242565 1.12e-08 1.8805896531808992 1.1201e-08 1.8407607237043373 1.1202e-08 1.7869658112052893 1.1203e-08 1.7684528019962098 1.1204e-08 1.7684989544884036 1.1205e-08 1.8224934105433632 1.1206e-08 1.6714846158925096 1.1206999999999999e-08 1.7599540267170493 1.1208e-08 1.7206996084485662 1.1209e-08 1.8706119555949379 1.1209999999999999e-08 1.8537366228509562 1.1211e-08 1.7360925795899407 1.1212e-08 1.846492678684048 1.1213e-08 1.7590743781504627 1.1214e-08 1.7895239718460567 1.1215e-08 1.892684449519886 1.1216e-08 1.8678064238089325 1.1217e-08 1.7578944816902746 1.1218e-08 1.7344658380862177 1.1219e-08 1.810505942928418 1.122e-08 1.7969357043572136 1.1221e-08 1.8112421460480732 1.1222e-08 1.703520372946843 1.1222999999999999e-08 1.7146642678232749 1.1224e-08 1.8219983459722762 1.1225e-08 1.738642079034534 1.1225999999999999e-08 1.7285581190774488 1.1227e-08 1.8796756440772573 1.1228e-08 1.7893756115943202 1.1228999999999999e-08 1.782874091232446 1.123e-08 1.7482052709724607 1.1231e-08 1.7863263592229968 1.1232e-08 1.771051587725348 1.1233e-08 1.7984410395096728 1.1234e-08 1.8542237484235378 1.1235e-08 1.7259960279802629 1.1236e-08 1.7101248742255413 1.1237e-08 1.8584375977081662 1.1238e-08 1.8497595211176148 1.1239e-08 1.867824829816132 1.124e-08 1.677387886644313 1.1241e-08 1.7587705514082355 1.1241999999999999e-08 1.7761737747131674 1.1243e-08 1.874736791746312 1.1244e-08 1.7941604729408553 1.1244999999999999e-08 1.8124016560602214 1.1246e-08 1.787923503227634 1.1247e-08 1.7084539449065306 1.1248e-08 1.7449428634546622 1.1249e-08 1.818260053253555 1.125e-08 1.7538461128427976 1.1251e-08 1.822473181275487 1.1252e-08 1.7311404314424204 1.1253e-08 1.7871895056122766 1.1254e-08 1.798348929015756 1.1255e-08 1.762267127216387 1.1256e-08 1.7629481887653047 1.1257e-08 1.7914608964442045 1.1257999999999999e-08 1.8552770912338967 1.1259e-08 1.8069805131026024 1.126e-08 1.725643553537869 1.1260999999999999e-08 1.7669914668388995 1.1262e-08 1.8020418749926637 1.1263e-08 1.7397393336133622 1.1263999999999999e-08 1.81209767300048 1.1265e-08 1.793830334982496 1.1266e-08 1.8247888283958966 1.1267e-08 1.8599736935874063 1.1268e-08 1.9003781256058778 1.1269e-08 1.8366953319907904 1.127e-08 1.7649737803146976 1.1271e-08 1.7425373473554355 1.1272e-08 1.8031773017303427 1.1273e-08 1.6734048312832774 1.1274e-08 1.8148992780804285 1.1275e-08 1.7329413050376052 1.1276e-08 1.8020742575335627 1.1276999999999999e-08 1.8711765906886906 1.1278e-08 1.7907928008153329 1.1279e-08 1.7673754334125436 1.1279999999999999e-08 1.777508236850341 1.1281e-08 1.747120850484974 1.1282e-08 1.8022856734268144 1.1283e-08 1.8424195818487952 1.1284e-08 1.8930479493347134 1.1285e-08 1.7619252785137776 1.1286e-08 1.8091716688473316 1.1287e-08 1.8313111495282421 1.1288e-08 1.866191126002962 1.1289e-08 1.86523414642576 1.129e-08 1.8414525824722299 1.1291e-08 1.8151188441890487 1.1292e-08 1.7478582463630083 1.1292999999999999e-08 1.863079682478486 1.1294e-08 1.7849655039270593 1.1295e-08 1.8176599470213377 1.1295999999999999e-08 1.9055245465035138 1.1297e-08 1.8538231251344701 1.1298e-08 1.8795916538068236 1.1298999999999999e-08 1.9034194800706234 1.13e-08 1.7986839152480028 1.1301e-08 1.758904677584429 1.1302e-08 1.8128875269827662 1.1303e-08 1.7813244670328758 1.1304e-08 1.7111521947262862 1.1305e-08 1.8207447778867736 1.1306e-08 1.7847869266994627 1.1307e-08 1.7741467832396398 1.1308e-08 1.8403937749356265 1.1309e-08 1.7329662277775444 1.131e-08 1.7840688727163676 1.1311e-08 1.8713414374863644 1.1311999999999999e-08 1.8717111371698314 1.1313e-08 1.8224747418874376 1.1314e-08 1.739635422589434 1.1314999999999999e-08 1.8173236662973355 1.1316e-08 1.868320169431667 1.1317e-08 1.7910869417674458 1.1318e-08 1.7950092064466858 1.1319e-08 1.713200128134391 1.132e-08 1.700440840659751 1.1321e-08 1.7199424347267178 1.1322e-08 1.7295640612536156 1.1323e-08 1.7168826763458025 1.1324e-08 1.8493824055335042 1.1325e-08 1.7767301949056014 1.1326e-08 1.7812564895439513 1.1327e-08 1.8460074344379778 1.1328e-08 1.7326966273268491 1.1329e-08 1.7694582742685396 1.133e-08 1.9401592740389868 1.1330999999999999e-08 1.7530651573581455 1.1332e-08 1.8096381277418876 1.1333e-08 1.792961285540453 1.1333999999999999e-08 1.7700034855656173 1.1335e-08 1.8290309053558134 1.1336e-08 1.7312365658629485 1.1337e-08 1.7639557161717545 1.1338e-08 1.7464402165850557 1.1339e-08 1.9167771737580876 1.134e-08 1.7944905521426953 1.1341e-08 1.832674852588009 1.1342e-08 1.8088021267093566 1.1343e-08 1.820217286996428 1.1344e-08 1.7265303851576252 1.1345e-08 1.715620497961188 1.1346e-08 1.7786284019570624 1.1346999999999999e-08 1.8332254303117432 1.1348e-08 1.7602539427745163 1.1349e-08 1.8073983651247123 1.1349999999999999e-08 1.8591326114751408 1.1351e-08 1.9350264243494533 1.1352e-08 1.8224260693970105 1.1352999999999999e-08 1.7919963076778695 1.1354e-08 1.8052297814747846 1.1355e-08 1.7747002414787705 1.1356e-08 1.8489447506047187 1.1357e-08 1.845778313331421 1.1358e-08 1.8015258247212826 1.1359e-08 1.7219682051226792 1.136e-08 1.742860359986857 1.1361e-08 1.7830596887920245 1.1362e-08 1.7787256820285022 1.1363e-08 1.7749716534079378 1.1364e-08 1.795463744263158 1.1365e-08 1.7876143772470683 1.1365999999999999e-08 1.8742643507563677 1.1367e-08 1.8212911061285884 1.1368e-08 1.8016086910495739 1.1368999999999999e-08 1.7508009322883382 1.137e-08 1.8320828654053019 1.1371e-08 1.7331289326931991 1.1372e-08 1.758740127951533 1.1373e-08 1.850409455099444 1.1374e-08 1.8463384901887685 1.1375e-08 1.8832260783468027 1.1376e-08 1.8361148495569666 1.1377e-08 1.8517519260362685 1.1378e-08 1.7992094991660181 1.1379e-08 1.8406807459886079 1.138e-08 1.790678851807173 1.1381e-08 1.7367695579065097 1.1381999999999999e-08 1.7071467497385397 1.1383e-08 1.8515482810148436 1.1384e-08 1.8033406887738674 1.1384999999999999e-08 1.768335742501122 1.1386e-08 1.8601810406237724 1.1387e-08 1.8317810838902606 1.1387999999999999e-08 1.7873040998645955 1.1389e-08 1.7878515074926287 1.139e-08 1.8158545934679566 1.1391e-08 1.8844356092954495 1.1392e-08 1.8336839519362473 1.1393e-08 1.7919271738448372 1.1394e-08 1.7914326664278173 1.1395e-08 1.8176854797661788 1.1396e-08 1.8601541155261814 1.1397e-08 1.7727069470055605 1.1398e-08 1.7697644336596892 1.1399e-08 1.804155165539969 1.14e-08 1.861936912833375 1.1400999999999999e-08 1.7480820803843844 1.1402e-08 1.7808758015018828 1.1403e-08 1.884475947210933 1.1403999999999999e-08 1.7317583629866315 1.1405e-08 1.753206553048044 1.1406e-08 1.7801273270749407 1.1407e-08 1.734121510459921 1.1408e-08 1.7664164959174642 1.1409e-08 1.8332482455732346 1.141e-08 1.7976600572468096 1.1411e-08 1.8031342641751869 1.1412e-08 1.7333438468801994 1.1413e-08 1.775549457840615 1.1414e-08 1.8100987013682825 1.1415e-08 1.824015820174123 1.1416e-08 1.8277667111340512 1.1417e-08 1.8551409316521024 1.1418e-08 1.840027427010904 1.1419e-08 1.7961427246508437 1.1419999999999999e-08 1.792105860450081 1.1421e-08 1.8139623858768659 1.1422e-08 1.836399431060296 1.1422999999999999e-08 1.7788390057946866 1.1424e-08 1.8584195790852893 1.1425e-08 1.7323689648757845 1.1426e-08 1.8174443889903311 1.1427e-08 1.795429488369979 1.1428e-08 1.783539959554008 1.1429e-08 1.737834960068688 1.143e-08 1.7715645633931716 1.1431e-08 1.837464537825074 1.1432e-08 1.7888303729695922 1.1433e-08 1.8449129859943494 1.1434e-08 1.8521514668569172 1.1435e-08 1.8208871180217765 1.1435999999999999e-08 1.7975501264282003 1.1437e-08 1.8136491093173137 1.1438e-08 1.8346437996028453 1.1438999999999999e-08 1.7316477685909453 1.144e-08 1.852971535162595 1.1441e-08 1.7601091414373031 1.1441999999999999e-08 1.8674351189399598 1.1443e-08 1.7722733869719878 1.1444e-08 1.8171981511026292 1.1445e-08 1.804287846218863 1.1446e-08 1.827051441051806 1.1447e-08 1.852943197907288 1.1448e-08 1.7935201355293493 1.1449e-08 1.816428061224641 1.145e-08 1.790885273690154 1.1451e-08 1.865699876903077 1.1452e-08 1.8618031863516329 1.1453e-08 1.8539727978547045 1.1454e-08 1.746882295189108 1.1454999999999999e-08 1.8594625618943672 1.1456e-08 1.7712222336631729 1.1457e-08 1.842949299454489 1.1457999999999999e-08 1.8152693151101433 1.1459e-08 1.8392393030965881 1.146e-08 1.7739489199266496 1.1461e-08 1.864803194420394 1.1462e-08 1.7781510803098595 1.1463e-08 1.8386002891462938 1.1464e-08 1.787117390731341 1.1465e-08 1.766128059194748 1.1466e-08 1.786221898469831 1.1467e-08 1.8570430804132099 1.1468e-08 1.8515420058109173 1.1469e-08 1.7401180788286932 1.147e-08 1.7653911378087688 1.1470999999999999e-08 1.8407718951842154 1.1472e-08 1.7263218841317436 1.1473e-08 1.8088278414593035 1.1473999999999999e-08 1.8477811209670623 1.1475e-08 1.7992122467167047 1.1476e-08 1.7900477092084917 1.1476999999999999e-08 1.7223761996702631 1.1478e-08 1.8400073355679407 1.1479e-08 1.7948986009841579 1.148e-08 1.8034392247670636 1.1481e-08 1.773945112521476 1.1482e-08 1.8240455771179553 1.1483e-08 1.7452511080185198 1.1484e-08 1.8423526540253758 1.1485e-08 1.8356319818071325 1.1486e-08 1.792801481080899 1.1487e-08 1.81714736131813 1.1488e-08 1.8658720964641091 1.1489e-08 1.8028823340177889 1.1489999999999999e-08 1.7913266202385278 1.1491e-08 1.7020329961203167 1.1492e-08 1.8293935388965599 1.1492999999999999e-08 1.8273582299323596 1.1494e-08 1.7625689216220457 1.1495e-08 1.8624922996155053 1.1496e-08 1.873398966532854 1.1497e-08 1.7942035179742626 1.1498e-08 1.7709456992386763 1.1499e-08 1.8183680795145727 1.15e-08 1.8406009296518362 1.1501e-08 1.8261779144887444 1.1502e-08 1.7849392801666704 1.1503e-08 1.8500909515302324 1.1504e-08 1.8187010095456582 1.1505e-08 1.8220393893610112 1.1506e-08 1.7817138133099253 1.1507e-08 1.7172440500234853 1.1508e-08 1.8218789665331834 1.1508999999999999e-08 1.7918603594076237 1.151e-08 1.8274898328424203 1.1511e-08 1.8493996029330282 1.1511999999999999e-08 1.8016088417936151 1.1513e-08 1.7878203088480267 1.1514e-08 1.8283641663978039 1.1515e-08 1.73036022850371 1.1516e-08 1.724611365035749 1.1517e-08 1.796831110512532 1.1518e-08 1.7749436064641329 1.1519e-08 1.8281720561349057 1.152e-08 1.831794743289961 1.1521e-08 1.7677830016678082 1.1522e-08 1.6449466866737763 1.1523e-08 1.7919050719255496 1.1524e-08 1.796012794806501 1.1524999999999999e-08 1.873841656122228 1.1526e-08 1.9256402236273615 1.1527e-08 1.8898487681080505 1.1527999999999999e-08 1.8574408027399427 1.1529e-08 1.6857451932178813 1.153e-08 1.7838895775395507 1.1530999999999999e-08 1.8927748592516096 1.1532e-08 1.7406731508306863 1.1533e-08 1.8883650276074007 1.1534e-08 1.8142021945543383 1.1535e-08 1.7060520922614173 1.1536e-08 1.7897174427816753 1.1537e-08 1.7617115637736689 1.1538e-08 1.7431511779939886 1.1539e-08 1.863193390368165 1.154e-08 1.7518550529001433 1.1541e-08 1.8641722645158214 1.1542e-08 1.8118403886973744 1.1543e-08 1.7751185450871867 1.1543999999999999e-08 1.7671045662277882 1.1545e-08 1.7297372584542536 1.1546e-08 1.8758835522415769 1.1546999999999999e-08 1.8493592330262707 1.1548e-08 1.7645369016212304 1.1549e-08 1.7428326293692158 1.155e-08 1.8432950527486172 1.1551e-08 1.9768988686993516 1.1552e-08 1.8329463773708732 1.1553e-08 1.7513752241145404 1.1554e-08 1.8180964356856573 1.1555e-08 1.7874393884762523 1.1556e-08 1.7830448941157067 1.1557e-08 1.7310556139081181 1.1558e-08 1.7613869665739585 1.1559e-08 1.8521811366801089 1.1559999999999999e-08 1.802629395143196 1.1561e-08 1.813747663422957 1.1562e-08 1.846235994753147 1.1562999999999999e-08 1.6927479464667226 1.1564e-08 1.7698544883132683 1.1565e-08 1.8021234692704613 1.1565999999999999e-08 1.8288795819783377 1.1567e-08 1.832908480744604 1.1568e-08 1.832081253845427 1.1569e-08 1.6924191023233908 1.157e-08 1.8721284834722538 1.1571e-08 1.9119310968558139 1.1572e-08 1.7466964647063392 1.1573e-08 1.7900459115960283 1.1574e-08 1.8588498298506713 1.1575e-08 1.8153242330522303 1.1576e-08 1.793518888718589 1.1577e-08 1.8284566875103632 1.1578e-08 1.7793318851851476 1.1578999999999999e-08 1.788194190316844 1.158e-08 1.7652523408793594 1.1581e-08 1.8332565961325935 1.1581999999999999e-08 1.8541832024119436 1.1583e-08 1.7639298554029128 1.1584e-08 1.8042471261611301 1.1585e-08 1.8398945252840935 1.1586e-08 1.8145230406839088 1.1587e-08 1.9289991664323678 1.1588e-08 1.8451644191502474 1.1589e-08 1.8169593075443329 1.159e-08 1.7536101477030361 1.1591e-08 1.7153888422341168 1.1592e-08 1.7517516509840905 1.1593e-08 1.8257290928683632 1.1594e-08 1.8495771626779205 1.1594999999999999e-08 1.7605383420140748 1.1596e-08 1.7588466612300404 1.1597e-08 1.834027706021359 1.1597999999999999e-08 1.7991136847124298 1.1599e-08 1.8153677519887854 1.16e-08 1.8124242754772604 1.1600999999999999e-08 1.7835896933282072 1.1602e-08 1.8870685458186098 1.1603e-08 1.801817467221314 1.1604e-08 1.827511104281367 1.1605e-08 1.860376518839834 1.1606e-08 1.759000110307833 1.1607e-08 1.7409327744256107 1.1608e-08 1.7845504679739117 1.1609e-08 1.7750418945324582 1.161e-08 1.8438193617903997 1.1611e-08 1.761407874833141 1.1612e-08 1.803525210816205 1.1613e-08 1.8353075951144697 1.1613999999999999e-08 1.9120809178984863 1.1615e-08 1.8062177753061892 1.1616e-08 1.847416900053328 1.1616999999999999e-08 1.8155303770357922 1.1618e-08 1.8212763952826794 1.1619e-08 1.8137102066982096 1.1619999999999999e-08 1.7703064646044333 1.1621e-08 1.8136995642149711 1.1622e-08 1.8751894122349038 1.1623e-08 1.8283457583882705 1.1624e-08 1.780102325717282 1.1625e-08 1.8526846357186193 1.1626e-08 1.8176676458654688 1.1627e-08 1.700485220147818 1.1628e-08 1.891314367831003 1.1629e-08 1.7845221774870828 1.163e-08 1.8004572530403178 1.1631e-08 1.7591869593460796 1.1632e-08 1.8207446684426551 1.1632999999999999e-08 1.851685595736578 1.1634e-08 1.775383474827302 1.1635e-08 1.7508845761176248 1.1635999999999999e-08 1.8190336956684057 1.1637e-08 1.8040158893907323 1.1638e-08 1.8055398928838382 1.1639e-08 1.780523554872576 1.164e-08 1.7883400256289173 1.1641e-08 1.7718809605858274 1.1642e-08 1.8140103748949319 1.1643e-08 1.771974408904961 1.1644e-08 1.7782340018994138 1.1645e-08 1.784212455810614 1.1646e-08 1.8145552156442195 1.1647e-08 1.7648571358898275 1.1648e-08 1.8795298412988704 1.1648999999999999e-08 1.7156859618319287 1.165e-08 1.768451362784043 1.1651e-08 1.8142607187780753 1.1651999999999999e-08 1.8084438010883404 1.1653e-08 1.6892115419089677 1.1654e-08 1.6844034228655334 1.1654999999999999e-08 1.836081169265568 1.1656e-08 1.7911466438821464 1.1657e-08 1.8410091025721715 1.1658e-08 1.7811216436832995 1.1659e-08 1.856945517400887 1.166e-08 1.7426865046719973 1.1661e-08 1.7624745733381806 1.1662e-08 1.7361058402670553 1.1663e-08 1.8045182822845411 1.1664e-08 1.8116095692287484 1.1665e-08 1.7499849039896276 1.1666e-08 1.7666946335913336 1.1667e-08 1.8304293085284478 1.1667999999999999e-08 1.8756943605922438 1.1669e-08 1.8613929123795374 1.167e-08 1.8336620868205318 1.1670999999999999e-08 1.8656148582710796 1.1672e-08 1.8566274851024562 1.1673e-08 1.6983830968418792 1.1674e-08 1.7982464709542783 1.1675e-08 1.7864747026257703 1.1676e-08 1.743685898081209 1.1677e-08 1.8560463015224902 1.1678e-08 1.7597056233568458 1.1679e-08 1.8027707248407228 1.168e-08 1.7950462309776456 1.1681e-08 1.7661812804213957 1.1682e-08 1.6414261809039254 1.1683e-08 1.7490295458753635 1.1683999999999999e-08 1.7654513094998687 1.1685e-08 1.8356494764201918 1.1686e-08 1.880266543894631 1.1686999999999999e-08 1.838334503382105 1.1688e-08 1.8476202136672477 1.1689e-08 1.7616868495365 1.1689999999999999e-08 1.74336640458928 1.1691e-08 1.7988160963491127 1.1692e-08 1.7123484178155954 1.1693e-08 1.779393104515745 1.1694e-08 1.833202803138733 1.1695e-08 1.7430905833976384 1.1696e-08 1.8408648788737172 1.1697e-08 1.7966905187754534 1.1698e-08 1.7822154797914427 1.1699e-08 1.806199483397283 1.17e-08 1.7086563246931026 1.1701e-08 1.7909644371021425 1.1702e-08 1.7229206059688922 1.1702999999999999e-08 1.7941647017502782 1.1704e-08 1.6895448228311487 1.1705e-08 1.6867767387315409 1.1705999999999999e-08 1.9234311307375356 1.1707e-08 1.786767126068457 1.1708e-08 1.7951146310616453 1.1708999999999999e-08 1.8041578490401404 1.171e-08 1.8470219180017267 1.1711e-08 1.8122621438362783 1.1712e-08 1.693913693271652 1.1713e-08 1.8075954276698056 1.1714e-08 1.7778991424936383 1.1715e-08 1.7999638649463119 1.1716e-08 1.7271232750545977 1.1717e-08 1.8074576885950067 1.1718e-08 1.812953412247093 1.1719e-08 1.706422375425296 1.172e-08 1.7441868459707455 1.1721e-08 1.8114856570267517 1.1721999999999999e-08 1.7374731494614861 1.1723e-08 1.835221125925938 1.1724e-08 1.8122617713057279 1.1724999999999999e-08 1.7877946669936864 1.1726e-08 1.7777281659408637 1.1727e-08 1.82375370021647 1.1728e-08 1.8286783094636625 1.1729e-08 1.8599795062987374 1.173e-08 1.9170037318199038 1.1731e-08 1.8590483578228005 1.1732e-08 1.7984915280494964 1.1733e-08 1.7709546980554984 1.1734e-08 1.7264429357668862 1.1735e-08 1.7412317114170692 1.1736e-08 1.8007894599538168 1.1737e-08 1.7508999225083457 1.1737999999999999e-08 1.7912003200756776 1.1739e-08 1.7448849600352858 1.174e-08 1.7975523918302374 1.1740999999999999e-08 1.8341412030531374 1.1742e-08 1.6899843599271167 1.1743e-08 1.8063323430717708 1.1743999999999999e-08 1.823569037255806 1.1745e-08 1.8584723441736883 1.1746e-08 1.8444723066944262 1.1747e-08 1.829529114119882 1.1748e-08 1.7512019916440482 1.1749e-08 1.8462915392854944 1.175e-08 1.8086593181907265 1.1751e-08 1.7920718158912503 1.1752e-08 1.8031616856391057 1.1753e-08 1.8149850949146538 1.1754e-08 1.8099948805472126 1.1755e-08 1.8506024552176843 1.1756e-08 1.8374383071469835 1.1756999999999999e-08 1.8306022290733643 1.1758e-08 1.8461750808097037 1.1759e-08 1.8031394812947406 1.1759999999999999e-08 1.8391523633115634 1.1761e-08 1.7934369983648528 1.1762e-08 1.7526916369992844 1.1763e-08 1.8690071970278457 1.1764e-08 1.882691052538777 1.1765e-08 1.810183043080507 1.1766e-08 1.804238908222226 1.1767e-08 1.7674124751797626 1.1768e-08 1.7824212135342676 1.1769e-08 1.9463195133850244 1.177e-08 1.8075936490822397 1.1771e-08 1.7191366548673053 1.1772e-08 1.8739367200698844 1.1772999999999999e-08 1.7911294115880525 1.1774e-08 1.8210519139462185 1.1775e-08 1.8664484939503796 1.1775999999999999e-08 1.893639994167286 1.1777e-08 1.7862612661605788 1.1778e-08 1.78803226874889 1.1778999999999999e-08 1.7188094054934187 1.178e-08 1.7968834296001452 1.1781e-08 1.824183464175248 1.1782e-08 1.7109112659152328 1.1783e-08 1.8210255988545818 1.1784e-08 1.7691511681630114 1.1785e-08 1.7248489818732984 1.1786e-08 1.7512105497956956 1.1787e-08 1.7664388311343286 1.1788e-08 1.8460862592143235 1.1789e-08 1.805065348476004 1.179e-08 1.751906082011584 1.1791e-08 1.7630826018320385 1.1791999999999999e-08 1.6486951477714413 1.1793e-08 1.7832610606104942 1.1794e-08 1.8191942965604126 1.1794999999999999e-08 1.8043137406668943 1.1796e-08 1.7466373739503431 1.1797e-08 1.8623072744367157 1.1797999999999999e-08 1.7417141293321434 1.1799e-08 1.7994026651869968 1.18e-08 1.768147228113954 1.1801e-08 1.7922271523831759 1.1802e-08 1.776577193375312 1.1803e-08 1.850571178294113 1.1804e-08 1.8986440193906648 1.1805e-08 1.7623625178627191 1.1806e-08 1.7711240129506947 1.1807e-08 1.7966034249794358 1.1808e-08 1.8385194721274938 1.1809e-08 1.8137546609654203 1.181e-08 1.8004467265503685 1.1810999999999999e-08 1.790118915249648 1.1812e-08 1.8280106559549547 1.1813e-08 1.7871105752312195 1.1813999999999999e-08 1.8200917674252526 1.1815e-08 1.823262539535303 1.1816e-08 1.752768019490171 1.1817e-08 1.9425154312690887 1.1818e-08 1.886082600979732 1.1819e-08 1.7926759376925132 1.182e-08 1.8242916038790882 1.1821e-08 1.7787193810202464 1.1822e-08 1.7961264480910257 1.1823e-08 1.8179417724606308 1.1824e-08 1.8031924511094362 1.1825e-08 1.793071793464864 1.1826e-08 1.7791383896461475 1.1826999999999999e-08 1.8395505327580428 1.1828e-08 1.792531848538641 1.1829e-08 1.7558555325200562 1.1829999999999999e-08 1.8115229394826389 1.1831e-08 1.7981147118403815 1.1832e-08 1.8376593702363708 1.1832999999999999e-08 1.792259553336697 1.1834e-08 1.7928573511242998 1.1835e-08 1.805754411072815 1.1836e-08 1.7394618954126133 1.1837e-08 1.8105271889482148 1.1838e-08 1.769975556890894 1.1839e-08 1.8579293903225897 1.184e-08 1.8513180281335935 1.1841e-08 1.8977444812359783 1.1842e-08 1.7824455905928311 1.1843e-08 1.8186800384188972 1.1844e-08 1.8392453911401188 1.1845e-08 1.8042637246213795 1.1845999999999999e-08 1.7758478199926944 1.1847e-08 1.722817606703421 1.1848e-08 1.8320301727766535 1.1848999999999999e-08 1.8068415488163785 1.185e-08 1.8076836758438541 1.1851e-08 1.7895464130925005 1.1852e-08 1.7405252871450911 1.1853e-08 1.8520717059305027 1.1854e-08 1.8395546378204914 1.1855e-08 1.8153255002339581 1.1856e-08 1.8907934405518945 1.1857e-08 1.8869755187422415 1.1858e-08 1.7190452381964605 1.1859e-08 1.8482867712811388 1.186e-08 1.7662027393015753 1.1861e-08 1.8033501977924562 1.1861999999999999e-08 1.7513898932714005 1.1863e-08 1.9041917166819997 1.1864e-08 1.9349758449650176 1.1864999999999999e-08 1.802256416892746 1.1866e-08 1.8007187308069237 1.1867e-08 1.741139793937838 1.1867999999999999e-08 1.8508715422746282 1.1869e-08 1.8200113269109006 1.187e-08 1.844597165306006 1.1871e-08 1.7664335379233802 1.1872e-08 1.855572023553445 1.1873e-08 1.7873806796033254 1.1874e-08 1.90282408423605 1.1875e-08 1.8200963055060138 1.1876e-08 1.8161175697989267 1.1877e-08 1.7393159488421306 1.1878e-08 1.8291084031094218 1.1879e-08 1.6917577833124695 1.188e-08 1.8629099356630547 1.1880999999999999e-08 1.7933154366825435 1.1882e-08 1.7343859557574843 1.1883e-08 1.7917573346151079 1.1883999999999999e-08 1.7485593637254384 1.1885e-08 1.7986878460851101 1.1886e-08 1.7271554589530689 1.1887e-08 1.8328019282112693 1.1888e-08 1.7340767394447285 1.1889e-08 1.7594408587470827 1.189e-08 1.8175071757863035 1.1891e-08 1.7650176284421162 1.1892e-08 1.7768686577767399 1.1893e-08 1.8355692492916214 1.1894e-08 1.820120048589921 1.1895e-08 1.763253028452455 1.1896e-08 1.7534186875335747 1.1897e-08 1.8038231223157424 1.1898e-08 1.859711803215497 1.1899e-08 1.737902970684456 1.1899999999999999e-08 1.8092520862447328 1.1901e-08 1.8719238233018611 1.1902e-08 1.7818420564475868 1.1902999999999999e-08 1.7962548260749802 1.1904e-08 1.82099756372651 1.1905e-08 1.8601251734116622 1.1906e-08 1.7842861882299865 1.1907e-08 1.7054347013302884 1.1908e-08 1.802403632359815 1.1909e-08 1.8150693616971003 1.191e-08 1.720136335758256 1.1911e-08 1.7959509459844765 1.1912e-08 1.7570962186600072 1.1913e-08 1.8693187496880035 1.1914e-08 1.8412345696775638 1.1915e-08 1.8128262744210506 1.1915999999999999e-08 1.7969144918913502 1.1917e-08 1.7914404154945525 1.1918e-08 1.8986376752807086 1.1918999999999999e-08 1.77180502958172 1.192e-08 1.812589999789318 1.1921e-08 1.8284820011323046 1.1921999999999999e-08 1.8138084283285507 1.1923e-08 1.8218276514546718 1.1924e-08 1.8371369876016448 1.1925e-08 1.6990319517045256 1.1926e-08 1.8448849529644762 1.1927e-08 1.8542403217034018 1.1928e-08 1.7501582433332499 1.1929e-08 1.8690074021862715 1.193e-08 1.7492316350136923 1.1931e-08 1.8645669344712996 1.1932e-08 1.8118013054509676 1.1933e-08 1.8595244235422344 1.1934e-08 1.8383204433435252 1.1934999999999999e-08 1.853525021509125 1.1936e-08 1.7461289980243724 1.1937e-08 1.825932451493058 1.1937999999999999e-08 1.703169998098544 1.1939e-08 1.8065833558775077 1.194e-08 1.822246061999306 1.1941e-08 1.807260013360111 1.1942e-08 1.852718170939771 1.1943e-08 1.7395625535303887 1.1944e-08 1.7844292036251064 1.1945e-08 1.846228189203948 1.1946e-08 1.7785296481979038 1.1947e-08 1.80147690096615 1.1948e-08 1.8286599843808053 1.1949e-08 1.7819546974171705 1.195e-08 1.787860176493564 1.1950999999999999e-08 1.8904221375035375 1.1952e-08 1.8004529947194279 1.1953e-08 1.7892806800761254 1.1953999999999999e-08 1.6543585835905432 1.1955e-08 1.7298565756113145 1.1956e-08 1.8013431516045646 1.1956999999999999e-08 1.7885314159413626 1.1958e-08 1.8805924082556404 1.1959e-08 1.8483639142091224 1.196e-08 1.8438521407100263 1.1961e-08 1.8016163456113297 1.1962e-08 1.807237213749532 1.1963e-08 1.7551575505510129 1.1964e-08 1.8266573733064468 1.1965e-08 1.7177970309554735 1.1966e-08 1.8574290888695593 1.1967e-08 1.817761297207489 1.1968e-08 1.8165736151454643 1.1969e-08 1.8215529266794563 1.1969999999999999e-08 1.787573480097265 1.1971e-08 1.8350227242797956 1.1972e-08 1.767325936066652 1.1972999999999999e-08 1.8470852458144478 1.1974e-08 1.8332163898357536 1.1975e-08 1.7818841837865134 1.1976e-08 1.7167444926092452 1.1977e-08 1.8702241028168238 1.1978e-08 1.8487155223231635 1.1979e-08 1.8385651866283266 1.198e-08 1.7318305834130656 1.1981e-08 1.7951538646032792 1.1982e-08 1.80552736315284 1.1983e-08 1.8326913394419626 1.1984e-08 1.7925962267615425 1.1985e-08 1.8324912190537066 1.1985999999999999e-08 1.7951177695722105 1.1987e-08 1.8329068695824393 1.1988e-08 1.731786651570549 1.1988999999999999e-08 1.772412675133909 1.199e-08 1.8274531727212853 1.1991e-08 1.8630483183593927 1.1991999999999999e-08 1.821961532490824 1.1993e-08 1.8002338156518505 1.1994e-08 1.820110583524409 1.1995e-08 1.826756476988337 1.1996e-08 1.8076869998345717 1.1997e-08 1.772157187390528 1.1998e-08 1.8882307120030302 1.1999e-08 1.7979905546267625 1.2e-08 1.7637868567107478 1.2001e-08 1.8650657849446026 1.2002e-08 1.8195419796162249 1.2003e-08 1.7915950987293696 1.2004e-08 1.870216055384468 1.2004999999999999e-08 1.7964342703121112 1.2006e-08 1.7621573312965209 1.2007e-08 1.7416833760836503 1.2007999999999999e-08 1.7680383578433798 1.2009e-08 1.7245248064185836 1.201e-08 1.782906285524856 1.2010999999999999e-08 1.8285620310278858 1.2012e-08 1.8077635605364981 1.2013e-08 1.8660960973615952 1.2014e-08 1.8251563249144929 1.2015e-08 1.800924779975803 1.2016e-08 1.8041721300998086 1.2017e-08 1.7797936327702024 1.2018e-08 1.8791879245746572 1.2019e-08 1.703955466880328 1.202e-08 1.7873290750662902 1.2021e-08 1.8894979936719203 1.2022e-08 1.8271279014803783 1.2023e-08 1.779192888609906 1.2023999999999999e-08 1.787650580738134 1.2025e-08 1.7809438789439587 1.2026e-08 1.8549734244352134 1.2026999999999999e-08 1.8407294677999428 1.2028e-08 1.8271124568557744 1.2029e-08 1.7477697038539832 1.203e-08 1.6977094102436645 1.2031e-08 1.8530739674487406 1.2032e-08 1.7975560230196916 1.2033e-08 1.790275132118386 1.2034e-08 1.763707009634428 1.2035e-08 1.8654263457553963 1.2036e-08 1.851823602705475 1.2037e-08 1.8061771342233324 1.2038e-08 1.7714134588094093 1.2039e-08 1.7392901373127823 1.2039999999999999e-08 1.8399331795243727 1.2041e-08 1.9194354907591684 1.2042e-08 1.8393408555898292 1.2042999999999999e-08 1.8282246779246223 1.2044e-08 1.8263516587973012 1.2045e-08 1.828370533147889 1.2045999999999999e-08 1.913696794486556 1.2047e-08 1.8682400724349082 1.2048e-08 1.8145384599288672 1.2049e-08 1.7626588163116916 1.205e-08 1.8294553661486217 1.2051e-08 1.7971041271458696 1.2052e-08 1.8180319788535264 1.2053e-08 1.9039146986816056 1.2054e-08 1.7524303512584707 1.2055e-08 1.8185424805787636 1.2056e-08 1.7931428884240586 1.2057e-08 1.8319034030199095 1.2058e-08 1.7612826596677758 1.2058999999999999e-08 1.7711032801021953 1.206e-08 1.8230658950915453 1.2061e-08 1.7555856908988319 1.2061999999999999e-08 1.8088843661227498 1.2063e-08 1.849109751513982 1.2064e-08 1.8122205977144477 1.2065e-08 1.833933986365346 1.2066e-08 1.7913309430249489 1.2067e-08 1.8797985594050697 1.2068e-08 1.779096386254474 1.2069e-08 1.8765928784954808 1.207e-08 1.716807834541822 1.2071e-08 1.7650390595472634 1.2072e-08 1.7534376282289494 1.2073e-08 1.7750815535529763 1.2074e-08 1.8006667171205466 1.2074999999999999e-08 1.8345150170596227 1.2076e-08 1.832876300079984 1.2077e-08 1.712350869969282 1.2077999999999999e-08 1.860678729976092 1.2079e-08 1.7602115855872913 1.208e-08 1.8429228145733694 1.2080999999999999e-08 1.8534378365449533 1.2082e-08 1.8710121123424415 1.2083e-08 1.8644516310712262 1.2084e-08 1.7820236040896051 1.2085e-08 1.7693579015490852 1.2086e-08 1.818188752586437 1.2087e-08 1.8863352384741854 1.2088e-08 1.8789347970028638 1.2089e-08 1.7738808927648095 1.209e-08 1.8143784764595732 1.2091e-08 1.8744325984411883 1.2092e-08 1.7977581799663251 1.2093e-08 1.706687810628091 1.2093999999999999e-08 1.7505440465372821 1.2095e-08 1.8089928450074106 1.2096e-08 1.779685137385083 1.2096999999999999e-08 1.7415098593433709 1.2098e-08 1.7419938841569622 1.2099e-08 1.8129153130135656 1.2099999999999999e-08 1.7998896478939268 1.2101e-08 1.8237818875256904 1.2102e-08 1.7575482061811376 1.2103e-08 1.8127970077389493 1.2104e-08 1.7637742889545416 1.2105e-08 1.8494316614481923 1.2106e-08 1.9140473369097852 1.2107e-08 1.792788980947409 1.2108e-08 1.8232645796511167 1.2109e-08 1.848430255281203 1.211e-08 1.8680295576274286 1.2111e-08 1.7644434231578527 1.2112e-08 1.8009896970678523 1.2112999999999999e-08 1.818268341079336 1.2114e-08 1.685755443782235 1.2115e-08 1.7453224089064703 1.2115999999999999e-08 1.7711361110572716 1.2117e-08 1.8489111119396877 1.2118e-08 1.7759869792225662 1.2119e-08 1.820681546390217 1.212e-08 1.8078646769255882 1.2121e-08 1.7684406870261409 1.2122e-08 1.8055186536096068 1.2123e-08 1.7539218741823426 1.2124e-08 1.8027304848469097 1.2125e-08 1.914022266688929 1.2126e-08 1.7373748943666318 1.2127e-08 1.7140221740096675 1.2128e-08 1.7787676279521145 1.2128999999999999e-08 1.7652135438031051 1.213e-08 1.8024550248351736 1.2131e-08 1.8763512639778757 1.2131999999999999e-08 1.8335783340234082 1.2133e-08 1.8177772614913252 1.2134e-08 1.8095603525812947 1.2134999999999999e-08 1.894420067944878 1.2136e-08 1.7977434439294835 1.2137e-08 1.7482980632538505 1.2138e-08 1.819832341443482 1.2139e-08 1.8777567374007127 1.214e-08 1.832729845925518 1.2141e-08 1.8063248363699755 1.2142e-08 1.7315638232974129 1.2143e-08 1.7474667207688412 1.2144e-08 1.8314780834973583 1.2145e-08 1.807087573746924 1.2146e-08 1.8799181511955052 1.2147e-08 1.8106836747228399 1.2147999999999999e-08 1.8262127441685232 1.2149e-08 1.817420610699417 1.215e-08 1.7559367270229955 1.2150999999999999e-08 1.8327442134415741 1.2152e-08 1.8321992295256748 1.2153e-08 1.8400915662574557 1.2154e-08 1.7466939998091142 1.2155e-08 1.8623158773933457 1.2156e-08 1.7922954823569794 1.2157e-08 1.8088353400327664 1.2158e-08 1.8289006573178157 1.2159e-08 1.7957527143227479 1.216e-08 1.6946828517187285 1.2161e-08 1.7266911980178974 1.2162e-08 1.8272361122266358 1.2163e-08 1.8082748972936873 1.2163999999999999e-08 1.8949468000134506 1.2165e-08 1.7625551804146846 1.2166e-08 1.7774657382346473 1.2166999999999999e-08 1.8743698788889538 1.2168e-08 1.778575531080537 1.2169e-08 1.8390909254882957 1.2169999999999999e-08 1.8062012617654708 1.2171e-08 1.7471081924946374 1.2172e-08 1.7647163351800763 1.2173e-08 1.8218903919032463 1.2174e-08 1.8233832970876351 1.2175e-08 1.8367611492210312 1.2176e-08 1.7978082440263419 1.2177e-08 1.7908663622769192 1.2178e-08 1.7137002828479444 1.2179e-08 1.7925118200874808 1.218e-08 1.8724076477910458 1.2181e-08 1.774772958208555 1.2182e-08 1.8213391443539995 1.2182999999999999e-08 1.8619771469820203 1.2184e-08 1.884578236641725 1.2185e-08 1.7426440580470552 1.2185999999999999e-08 1.7334311404212586 1.2187e-08 1.7561169226844964 1.2188e-08 1.7768440594088568 1.2188999999999999e-08 1.786473353870458 1.219e-08 1.7516547155542757 1.2191e-08 1.673617157589251 1.2192e-08 1.7647748917234032 1.2193e-08 1.8538249131296278 1.2194e-08 1.733712757197112 1.2195e-08 1.7399929364978481 1.2196e-08 1.7605902737205164 1.2197e-08 1.7308679398740823 1.2198e-08 1.774738790197676 1.2199e-08 1.8089141457106608 1.22e-08 1.7669009948525414 1.2201e-08 1.7787012763576415 1.2201999999999999e-08 1.761094886597017 1.2203e-08 1.786951755002384 1.2204e-08 1.7525165055195557 1.2204999999999999e-08 1.7779373437420618 1.2206e-08 1.7818666262123635 1.2207e-08 1.7927668227437028 1.2208e-08 1.7716242031796148 1.2209e-08 1.8388319640331843 1.221e-08 1.8689539237494883 1.2211e-08 1.8572053620377538 1.2212e-08 1.8872224224315164 1.2213e-08 1.7622718115093519 1.2214e-08 1.769317783642454 1.2215e-08 1.789983955844229 1.2216e-08 1.837667119618435 1.2217e-08 1.7731511878630566 1.2217999999999999e-08 1.7759117635407695 1.2219e-08 1.8249089403186065 1.222e-08 1.8715646238655208 1.2220999999999999e-08 1.7821499444572888 1.2222e-08 1.8157705415968448 1.2223e-08 1.8897306778623695 1.2223999999999999e-08 1.7721125350246787 1.2225e-08 1.7607863330257898 1.2226e-08 1.8254780155252277 1.2227e-08 1.6682342067748746 1.2228e-08 1.8964023825371004 1.2229e-08 1.8148559187092836 1.223e-08 1.7963820419407615 1.2231e-08 1.8108067748377712 1.2232e-08 1.7425396903815185 1.2233e-08 1.7962436871102476 1.2234e-08 1.7633052541031538 1.2235e-08 1.9057584452380592 1.2236e-08 1.8134233491015104 1.2236999999999999e-08 1.8287940208463136 1.2238e-08 1.7429362194024525 1.2239e-08 1.837081800144356 1.2239999999999999e-08 1.7356183249365726 1.2241e-08 1.715444490205092 1.2242e-08 1.8134416880884818 1.2243e-08 1.7590551150552074 1.2244e-08 1.8888706960782198 1.2245e-08 1.8286964073021443 1.2246e-08 1.8288307050098473 1.2247e-08 1.7898962188967653 1.2248e-08 1.7665885343043415 1.2249e-08 1.768204032165394 1.225e-08 1.796257703558406 1.2251e-08 1.8701670189086483 1.2252e-08 1.808121864072557 1.2252999999999999e-08 1.8089118895640122 1.2254e-08 1.7942851919477105 1.2255e-08 1.816118545287038 1.2255999999999999e-08 1.8512837995826568 1.2257e-08 1.8387723338751583 1.2258e-08 1.8176765681251275 1.2258999999999999e-08 1.830711117697545 1.226e-08 1.7803142274066746 1.2261e-08 1.69652628430492 1.2262e-08 1.7549249192760328 1.2263e-08 1.775243877567384 1.2264e-08 1.8246631056642557 1.2265e-08 1.732999184420145 1.2266e-08 1.8102522281826467 1.2267e-08 1.8215510113017948 1.2268e-08 1.7694309102399977 1.2269e-08 1.7998921217319341 1.227e-08 1.7722225986828617 1.2271e-08 1.7902308864201393 1.2271999999999999e-08 1.8308327979398829 1.2273e-08 1.826936781393953 1.2274e-08 1.8223640923585893 1.2274999999999999e-08 1.8209430535182052 1.2276e-08 1.678281892555793 1.2277e-08 1.7960723070186897 1.2277999999999999e-08 1.8073540353847282 1.2279e-08 1.8383913785559993 1.228e-08 1.834772245728567 1.2281e-08 1.7820786064816327 1.2282e-08 1.8596687300127506 1.2283e-08 1.8527817925840935 1.2284e-08 1.7625455965296648 1.2285e-08 1.814107678543157 1.2286e-08 1.8343807672289818 1.2287e-08 1.7380657586480537 1.2288e-08 1.718893711147131 1.2289e-08 1.8833931715071657 1.229e-08 1.748387094139412 1.2290999999999999e-08 1.877483163339027 1.2292e-08 1.8235792116267031 1.2293e-08 1.8409106343464052 1.2293999999999999e-08 1.7698930028676623 1.2295e-08 1.7958013922241143 1.2296e-08 1.6986953205671194 1.2297e-08 1.7957091984035867 1.2298e-08 1.8335329661479383 1.2299e-08 1.8748255408837966 1.23e-08 1.783108899773301 1.2301e-08 1.8319399663753988 1.2302e-08 1.754085718820702 1.2303e-08 1.8066189913298512 1.2304e-08 1.7731287978930423 1.2305e-08 1.8534422617825166 1.2306e-08 1.8641008327793214 1.2306999999999999e-08 1.767043415945501 1.2308e-08 1.7510908028215584 1.2309e-08 1.7444341184042245 1.2309999999999999e-08 1.8515408769927304 1.2311e-08 1.8379217758297979 1.2312e-08 1.7561190797229143 1.2312999999999999e-08 1.8804242579130253 1.2314e-08 1.7929192153243556 1.2315e-08 1.8429559034615197 1.2316e-08 1.7897827752441844 1.2317e-08 1.8157798617208896 1.2318e-08 1.7354030865006123 1.2319e-08 1.8692077138588965 1.232e-08 1.802770199337027 1.2321e-08 1.9201791026721833 1.2322e-08 1.8828504959641272 1.2323e-08 1.782684241565637 1.2324e-08 1.838687424030125 1.2325e-08 1.7848254204028384 1.2325999999999999e-08 1.7464552992759423 1.2327e-08 1.7819106670660663 1.2328e-08 1.7740837428578953 1.2328999999999999e-08 1.7934253598514127 1.233e-08 1.828951101655296 1.2331e-08 1.7505048116707707 1.2332e-08 1.7259764574270355 1.2333e-08 1.778280798220488 1.2334e-08 1.9014653196896831 1.2335e-08 1.7331763104802065 1.2336e-08 1.791042380347207 1.2337e-08 1.7505852154293904 1.2338e-08 1.7279321694818368 1.2339e-08 1.7910172934181652 1.234e-08 1.7927776747340056 1.2341e-08 1.8532541510805933 1.2341999999999999e-08 1.7569787980009233 1.2343e-08 1.8190419129222173 1.2344e-08 1.7532988768388165 1.2344999999999999e-08 1.8121954063200159 1.2346e-08 1.8008964983687832 1.2347e-08 1.8245471643456692 1.2347999999999999e-08 1.8174246381817087 1.2349e-08 1.6862819751646507 1.235e-08 1.8081370624527526 1.2351e-08 1.7658695351791893 1.2352e-08 1.7029467742942879 1.2353e-08 1.8816444904759488 1.2354e-08 1.837589458260854 1.2355e-08 1.8657862515240304 1.2356e-08 1.7967412931580597 1.2357e-08 1.7835460871213198 1.2358e-08 1.8833486332350495 1.2359e-08 1.830188157433419 1.236e-08 1.8873013170327486 1.2360999999999999e-08 1.7665733001521349 1.2362e-08 1.821219457514062 1.2363e-08 1.768226818781608 1.2363999999999999e-08 1.832348259795637 1.2365e-08 1.7751028584201771 1.2366e-08 1.8048450114580816 1.2366999999999999e-08 1.8313494072159693 1.2368e-08 1.740111853199438 1.2369e-08 1.760447251224976 1.237e-08 1.8439035888186803 1.2371e-08 1.858526405338785 1.2372e-08 1.808133933997143 1.2373e-08 1.7624586619052995 1.2374e-08 1.747404890905262 1.2375e-08 1.8456313375165312 1.2376e-08 1.903597629169524 1.2376999999999999e-08 1.798710854760916 1.2378e-08 1.7387391442875026 1.2379e-08 1.7209925973880367 1.2379999999999999e-08 1.8318269388801858 1.2381e-08 1.7852204552582809 1.2382e-08 1.7594363569600948 1.2382999999999999e-08 1.7970367156737959 1.2384e-08 1.7147213703676436 1.2385e-08 1.8405316260524964 1.2386e-08 1.7571721336462405 1.2387e-08 1.858022208771531 1.2388e-08 1.8234105055177283 1.2389e-08 1.819561731994981 1.239e-08 1.8268299554208964 1.2391e-08 1.8481967166625375 1.2392e-08 1.7847813566024255 1.2393e-08 1.8433502767262728 1.2394e-08 1.7967698842161504 1.2395e-08 1.8076301269894202 1.2395999999999999e-08 1.7984953751335007 1.2397e-08 1.835084680263215 1.2398e-08 1.8174544449769383 1.2398999999999999e-08 1.8652510246442073 1.24e-08 1.7980420092986815 1.2401e-08 1.8287444061511235 1.2401999999999999e-08 1.7766768455214312 1.2403e-08 1.7788875120830487 1.2404e-08 1.8201879252415478 1.2405e-08 1.8321944980401257 1.2406e-08 1.760883097751964 1.2407e-08 1.883258741463872 1.2408e-08 1.684789075547232 1.2409e-08 1.8430493742818546 1.241e-08 1.807126996036781 1.2411e-08 1.7516299182383939 1.2412e-08 1.775321785743656 1.2413e-08 1.7663304969668272 1.2414e-08 1.8366601924165937 1.2414999999999999e-08 1.810293660318603 1.2416e-08 1.8767581205376018 1.2417e-08 1.7488356714747468 1.2417999999999999e-08 1.8612504384305666 1.2419e-08 1.7576766075417813 1.242e-08 1.7016814430676217 1.2421e-08 1.894254759924193 1.2422e-08 1.7906950437507405 1.2423e-08 1.787327423309985 1.2424e-08 1.7533117970838135 1.2425e-08 1.7957424698717723 1.2426e-08 1.8085418557095876 1.2427e-08 1.8432070585990195 1.2428e-08 1.7493324153240297 1.2429e-08 1.7225269767272389 1.243e-08 1.8035104565449505 1.2430999999999999e-08 1.8432558655834121 1.2432e-08 1.742453990230488 1.2433e-08 1.8079053527027515 1.2433999999999999e-08 1.7505941286157467 1.2435e-08 1.829840942181968 1.2436e-08 1.8396072517806161 1.2436999999999999e-08 1.7763034305219956 1.2438e-08 1.8846137085804102 1.2439e-08 1.8030310537963135 1.244e-08 1.8451798872464062 1.2441e-08 1.914667080251441 1.2442e-08 1.7685863266031217 1.2443e-08 1.8099783728777559 1.2444e-08 1.8464690335583611 1.2445e-08 1.8349444607491783 1.2446e-08 1.7964035638494615 1.2447e-08 1.8648326075637567 1.2448e-08 1.7905725830816261 1.2449e-08 1.8184363107204395 1.2449999999999999e-08 1.830346854030122 1.2451e-08 1.8170908207259229 1.2452e-08 1.7849112926288349 1.2452999999999999e-08 1.7596469185300245 1.2454e-08 1.8480431880453054 1.2455e-08 1.8098114965414933 1.2455999999999999e-08 1.8398372477144522 1.2457e-08 1.8065246190217394 1.2458e-08 1.7489738171646192 1.2459e-08 1.7238705486046682 1.246e-08 1.805896185699643 1.2461e-08 1.8487471018994315 1.2462e-08 1.8260139108566253 1.2463e-08 1.8592586505334023 1.2464e-08 1.8851948562828886 1.2465e-08 1.6996695047337451 1.2465999999999999e-08 1.7930610305442738 1.2467e-08 1.8534244598555807 1.2468e-08 1.7165695939358259 1.2468999999999999e-08 1.7912156427528358 1.247e-08 1.7719585091489463 1.2471e-08 1.894917783778049 1.2471999999999999e-08 1.7861620847291635 1.2473e-08 1.8531443488484471 1.2474e-08 1.811895757508094 1.2475e-08 1.8209088665711914 1.2476e-08 1.7807663810495664 1.2477e-08 1.823246587774358 1.2478e-08 1.6681532749288512 1.2479e-08 1.7922019238532148 1.248e-08 1.8791681170708858 1.2481e-08 1.777140971860185 1.2482e-08 1.7626692683720895 1.2483e-08 1.7584995180312988 1.2484e-08 1.7910174192334805 1.2484999999999999e-08 1.7776314617048445 1.2486e-08 1.7208494297287997 1.2487e-08 1.7795209574336672 1.2487999999999999e-08 1.807437353106175 1.2489e-08 1.839641736470896 1.249e-08 1.8369025487406225 1.2490999999999999e-08 1.802256592651405 1.2492e-08 1.8100658996293453 1.2493e-08 1.7612447459899272 1.2494e-08 1.8057341108002931 1.2495e-08 1.7597594500882394 1.2496e-08 1.7473685322535826 1.2497e-08 1.7882075382365021 1.2498e-08 1.7993745832548562 1.2499e-08 1.7577686966684396 1.25e-08 1.7774549890981115 1.2501e-08 1.7279942076356172 1.2502e-08 1.781359233216506 1.2503e-08 1.8510155247251046 1.2503999999999999e-08 1.7695158039995056 1.2505e-08 1.8355623726772177 1.2506e-08 1.7823820922463272 1.2506999999999999e-08 1.7872023867157705 1.2508e-08 1.8142455656148462 1.2509e-08 1.7579918003265054 1.251e-08 1.862523044989111 1.2511e-08 1.7959060454743045 1.2512e-08 1.9042250420288913 1.2513e-08 1.8210188330583765 1.2514e-08 1.798008274681384 1.2515e-08 1.8221515132590316 1.2516e-08 1.7967493989716814 1.2517e-08 1.712743023704278 1.2518e-08 1.6819469777228369 1.2519e-08 1.8040170698918512 1.2519999999999999e-08 1.785610258619256 1.2521e-08 1.8473594799964825 1.2522e-08 1.8251042840201226 1.2522999999999999e-08 1.8263802994971507 1.2524e-08 1.8161963860907833 1.2525e-08 1.8198064601920614 1.2525999999999999e-08 1.820625863785098 1.2527e-08 1.7709617986499628 1.2528e-08 1.7755258901931683 1.2529e-08 1.8190253732460147 1.253e-08 1.8301993422574114 1.2531e-08 1.79060635054318 1.2532e-08 1.7565308080596087 1.2533e-08 1.7153127864020543 1.2534e-08 1.8469953584322538 1.2535e-08 1.8089925959792448 1.2536e-08 1.7986664499719107 1.2537e-08 1.7351359109010758 1.2538e-08 1.829864971404192 1.2538999999999999e-08 1.7859139656676146 1.254e-08 1.8608123108459669 1.2541e-08 1.8195003242385246 1.2541999999999999e-08 1.815669499256853 1.2543e-08 1.780887426777325 1.2544e-08 1.7651877329365044 1.2545e-08 1.804897863733788 1.2546e-08 1.8277959133855102 1.2547e-08 1.8537779482139753 1.2548e-08 1.7867928573761804 1.2549e-08 1.7231189104864584 1.255e-08 1.8029363431903738 1.2551e-08 1.7834745779561365 1.2552e-08 1.80964590903075 1.2553e-08 1.7849314796553408 1.2554e-08 1.8133427927965795 1.2554999999999999e-08 1.8922432280357038 1.2556e-08 1.781180681547717 1.2557e-08 1.8474715410681244 1.2557999999999999e-08 1.8211606792915727 1.2559e-08 1.9251971692834147 1.256e-08 1.7910405047988593 1.2560999999999999e-08 1.7964596423897667 1.2562e-08 1.7233951746041665 1.2563e-08 1.8251564908288849 1.2564e-08 1.7491564009540042 1.2565e-08 1.8431275784770063 1.2566e-08 1.8537950606535807 1.2567e-08 1.8725603072074675 1.2568e-08 1.731498313742033 1.2569e-08 1.7680220490977008 1.257e-08 1.8615764513243545 1.2571e-08 1.7934013090793604 1.2572e-08 1.8180537482990582 1.2573e-08 1.7977211461426306 1.2573999999999999e-08 1.8278072965257033 1.2575e-08 1.8380524857149774 1.2576e-08 1.8811733377881434 1.2576999999999999e-08 1.840873467640886 1.2578e-08 1.8738034032619606 1.2579e-08 1.806525696796177 1.2579999999999999e-08 1.7539066501382776 1.2581e-08 1.8671705664577825 1.2582e-08 1.7399656083948098 1.2583e-08 1.840511814565177 1.2584e-08 1.7651738627455977 1.2585e-08 1.8116825697283514 1.2586e-08 1.8328841739618207 1.2587e-08 1.8221846356513731 1.2588e-08 1.707906939453778 1.2589e-08 1.7927918990036522 1.259e-08 1.756763626563361 1.2591e-08 1.8571339246219174 1.2592e-08 1.8570662294195317 1.2592999999999999e-08 1.7240932441638048 1.2594e-08 1.8106712362586022 1.2595e-08 1.7263148241692257 1.2595999999999999e-08 1.7206532619900503 1.2597e-08 1.80980785179644 1.2598e-08 1.8032171634299412 1.2599e-08 1.764933326787139 1.26e-08 1.753324962723993 1.2601e-08 1.8189297805222264 1.2602e-08 1.775227992027527 1.2603e-08 1.8862578355503972 1.2604e-08 1.750514955307143 1.2605e-08 1.7498090083678346 1.2606e-08 1.818534455919414 1.2607e-08 1.7411429622934658 1.2608e-08 1.7885372232041534 1.2608999999999999e-08 1.8327595991565684 1.261e-08 1.7784221800539395 1.2611e-08 1.8510097691872742 1.2611999999999999e-08 1.764745992140869 1.2613e-08 1.8592226396198972 1.2614e-08 1.78898846319585 1.2614999999999999e-08 1.8326347793255084 1.2616e-08 1.8235221607625973 1.2617e-08 1.779233526840224 1.2618e-08 1.8288897317156685 1.2619e-08 1.9220315134892927 1.262e-08 1.8384926814976874 1.2621e-08 1.8112482464806499 1.2622e-08 1.8406286044329494 1.2623e-08 1.7276628252349915 1.2624e-08 1.8409668615938268 1.2625e-08 1.7744811711669466 1.2626e-08 1.7987852686167434 1.2627e-08 1.8275710729299341 1.2627999999999999e-08 1.7431957350348635 1.2629e-08 1.7105864030501328 1.263e-08 1.7769928250854896 1.2630999999999999e-08 1.8497927132571987 1.2632e-08 1.8443586792477096 1.2633e-08 1.754683132224925 1.2634e-08 1.8061280873037973 1.2635e-08 1.9185249211088224 1.2636e-08 1.7474435209995016 1.2637e-08 1.7874421436865375 1.2638e-08 1.7459174895120753 1.2639e-08 1.7839769403071282 1.264e-08 1.715947939201304 1.2641e-08 1.7816578971857588 1.2642e-08 1.879614977658823 1.2643e-08 1.7934883927721081 1.2643999999999999e-08 1.7271283701463018 1.2645e-08 1.8451995567598658 1.2646e-08 1.8122743632213336 1.2646999999999999e-08 1.8117530019295358 1.2648e-08 1.7891852822701841 1.2649e-08 1.7808696165220652 1.2649999999999999e-08 1.8055193164104297 1.2651e-08 1.7950809942115333 1.2652e-08 1.874950026707005 1.2653e-08 1.828358753119268 1.2654e-08 1.795565252929627 1.2655e-08 1.7742444616217454 1.2656e-08 1.8305799687693864 1.2657e-08 1.722032764838806 1.2658e-08 1.8161924496614952 1.2659e-08 1.8487591752446777 1.266e-08 1.734549472289322 1.2661e-08 1.8246367968922745 1.2662e-08 1.8127885778681017 1.2662999999999999e-08 1.8450000481270223 1.2664e-08 1.793521483531294 1.2665e-08 1.7260688556838133 1.2665999999999999e-08 1.852885944582526 1.2667e-08 1.8559417543558672 1.2668e-08 1.8246879721955567 1.2668999999999999e-08 1.7867381512778044 1.267e-08 1.8078211879537822 1.2671e-08 1.81127610484904 1.2672e-08 1.8337746495032858 1.2673e-08 1.8573588838717 1.2674e-08 1.8119813340972906 1.2675e-08 1.8292035211600726 1.2676e-08 1.7650336431016194 1.2677e-08 1.7821496173861007 1.2678e-08 1.7668651307700187 1.2678999999999999e-08 1.6971324726306376 1.268e-08 1.7986524620749542 1.2681e-08 1.9097128601872746 1.2681999999999999e-08 1.8777635827156356 1.2683e-08 1.8415899929377566 1.2684e-08 1.7482651464872652 1.2684999999999999e-08 1.7786870183067423 1.2686e-08 1.8825502556335185 1.2687e-08 1.867730913677615 1.2688e-08 1.7980259341950415 1.2689e-08 1.776999141465409 1.269e-08 1.7760779768918655 1.2691e-08 1.8238933694663122 1.2692e-08 1.8696207188156186 1.2693e-08 1.772785135860987 1.2694e-08 1.8340925005288478 1.2695e-08 1.7373695614699898 1.2696e-08 1.7618644489064084 1.2697e-08 1.7927742705741243 1.2697999999999999e-08 1.7613906089713247 1.2699e-08 1.8420714082452454 1.27e-08 1.7173078656356948 1.2700999999999999e-08 1.874266571342135 1.2702e-08 1.762219463919732 1.2703e-08 1.9168402655960668 1.2703999999999999e-08 1.7978311403654992 1.2705e-08 1.8136337130880187 1.2706e-08 1.7772106044649165 1.2707e-08 1.78959171673239 1.2708e-08 1.7227010879710665 1.2709e-08 1.797551394960363 1.271e-08 1.7527434906890829 1.2711e-08 1.7484086819965998 1.2712e-08 1.7585529810067904 1.2713e-08 1.8251196435039334 1.2714e-08 1.7776764860065748 1.2715e-08 1.7901053393971154 1.2716e-08 1.8365450756445556 1.2716999999999999e-08 1.8255403339351983 1.2718e-08 1.8060872632959546 1.2719e-08 1.8631514478083342 1.2719999999999999e-08 1.7823882932337638 1.2721e-08 1.795294349929571 1.2722e-08 1.7976944169806595 1.2723e-08 1.7993204313497708 1.2724e-08 1.8542772750081757 1.2725e-08 1.8425794567187883 1.2726e-08 1.78277478883694 1.2727e-08 1.7449694919230874 1.2728e-08 1.8385120425053187 1.2729e-08 1.818494135924974 1.273e-08 1.733241697718485 1.2731e-08 1.8702317470488448 1.2732e-08 1.827886034208202 1.2732999999999999e-08 1.8472993202648313 1.2734e-08 1.7407825253487106 1.2735e-08 1.7696208634198614 1.2735999999999999e-08 1.7634603745887376 1.2737e-08 1.7910830561648972 1.2738e-08 1.7928974841456964 1.2738999999999999e-08 1.8613863087985996 1.274e-08 1.7793413310573738 1.2741e-08 1.7531266607970672 1.2742e-08 1.8140789596221074 1.2743e-08 1.847931464571052 1.2744e-08 1.8514491781169502 1.2745e-08 1.7686149061452852 1.2746e-08 1.8104630971116273 1.2747e-08 1.7920396270376036 1.2748e-08 1.7929049346264878 1.2749e-08 1.8628442568500736 1.275e-08 1.8264776971359347 1.2751e-08 1.8067907831936991 1.2751999999999999e-08 1.759568656579655 1.2753e-08 1.8340764593543806 1.2754e-08 1.7054818211515708 1.2754999999999999e-08 1.7890324350189073 1.2756e-08 1.8603149361953857 1.2757e-08 1.7762534396598868 1.2757999999999999e-08 1.7848342044790568 1.2759e-08 1.8435102856708605 1.276e-08 1.7755990481943027 1.2761e-08 1.8415276707895283 1.2762e-08 1.7918289023107947 1.2763e-08 1.7886752575628118 1.2764e-08 1.8332626359777442 1.2765e-08 1.7856873972023255 1.2766e-08 1.7381235858860347 1.2767e-08 1.7973667867621692 1.2767999999999999e-08 1.7981806459196925 1.2769e-08 1.8740579740626437 1.277e-08 1.8552325515952806 1.2770999999999999e-08 1.693551558835756 1.2772e-08 1.8530842047740643 1.2773e-08 1.7864319118941467 1.2773999999999999e-08 1.757726001206814 1.2775e-08 1.8382750105368793 1.2776e-08 1.7910639741353005 1.2777e-08 1.770716792246982 1.2778e-08 1.7789739126144815 1.2779e-08 1.7882211653193687 1.278e-08 1.796872658980904 1.2781e-08 1.8243732985505243 1.2782e-08 1.879363235920285 1.2783e-08 1.9089597972308083 1.2784e-08 1.7610326364426525 1.2785e-08 1.804806370230468 1.2786e-08 1.8194729496467845 1.2786999999999999e-08 1.8163116946847688 1.2788e-08 1.8426578638671163 1.2789e-08 1.8188087826693244 1.2789999999999999e-08 1.8277534078355182 1.2791e-08 1.8272679745654286 1.2792e-08 1.8195617812811953 1.2792999999999999e-08 1.7611713406720928 1.2794e-08 1.8545685848626932 1.2795e-08 1.798995259181826 1.2796e-08 1.8499325120832972 1.2797e-08 1.9308620562085408 1.2798e-08 1.7730591806039617 1.2799e-08 1.774753745413298 1.28e-08 1.75477294148203 1.2801e-08 1.7619944680921409 1.2802e-08 1.7858802339137136 1.2803e-08 1.859307762602382 1.2804e-08 1.8077502732952488 1.2805e-08 1.7232083771907962 1.2805999999999999e-08 1.7650014343105451 1.2807e-08 1.8391870535662556 1.2808e-08 1.7698581124384174 1.2808999999999999e-08 1.8565835682155445 1.281e-08 1.809312123916396 1.2811e-08 1.794545934369545 1.2812e-08 1.831708843240767 1.2813e-08 1.756557485249244 1.2814e-08 1.7888762331029557 1.2815e-08 1.7058657773083516 1.2816e-08 1.8587571185107625 1.2817e-08 1.8661585798730678 1.2818e-08 1.8115343549021414 1.2819e-08 1.853622839345904 1.282e-08 1.868533462980748 1.2821e-08 1.76446937563076 1.2821999999999999e-08 1.818599413800566 1.2823e-08 1.7607471081082917 1.2824e-08 1.695672990291071 1.2824999999999999e-08 1.8527538585476635 1.2826e-08 1.754732354425252 1.2827e-08 1.9442427063515986 1.2827999999999999e-08 1.9372364526633894 1.2829e-08 1.7704641150362832 1.283e-08 1.7952508763775865 1.2831e-08 1.8638519503547473 1.2832e-08 1.7954147182801283 1.2833e-08 1.7722163491617022 1.2834e-08 1.80336219128846 1.2835e-08 1.8227578550512678 1.2836e-08 1.8422119280998797 1.2837e-08 1.868665453111574 1.2838e-08 1.7874124207078284 1.2839e-08 1.7456222466593183 1.284e-08 1.8483087418234743 1.2840999999999999e-08 1.8262597917447616 1.2842e-08 1.7837075670242866 1.2843e-08 1.7167590164541653 1.2843999999999999e-08 1.786508785061694 1.2845e-08 1.7464310521299327 1.2846e-08 1.8607316111624974 1.2846999999999999e-08 1.772331044923959 1.2848e-08 1.812061660561757 1.2849e-08 1.7149923179699176 1.285e-08 1.7917446393264205 1.2851e-08 1.7012482866994227 1.2852e-08 1.6857810514506717 1.2853e-08 1.9061771552962625 1.2854e-08 1.7388608828350336 1.2855e-08 1.8131864808399865 1.2856e-08 1.8008542320076935 1.2856999999999999e-08 1.714227100447874 1.2858e-08 1.7845513552928063 1.2859e-08 1.7958033266667877 1.2859999999999999e-08 1.8446814586123574 1.2861e-08 1.8083355340313974 1.2862e-08 1.7832807368450472 1.2862999999999999e-08 1.7779023585648055 1.2864e-08 1.8054882701252246 1.2865e-08 1.7678460294720146 1.2866e-08 1.810510845422044 1.2867e-08 1.782587635491468 1.2868e-08 1.7873166342698166 1.2869e-08 1.8213633504569766 1.287e-08 1.808997646219019 1.2871e-08 1.9174647965004281 1.2872e-08 1.8439335941728527 1.2873e-08 1.8350242283950728 1.2874e-08 1.7688923240011571 1.2875e-08 1.81889915403598 1.2875999999999999e-08 1.7615088637365548 1.2877e-08 1.8070756839976418 1.2878e-08 1.7663625549066606 1.2878999999999999e-08 1.7967423055635865 1.288e-08 1.8394927166830992 1.2881e-08 1.8974649407513826 1.2881999999999999e-08 1.8307232565780984 1.2883e-08 1.8099165307944134 1.2884e-08 1.8748574958643898 1.2885e-08 1.7985476759601375 1.2886e-08 1.7656017793257635 1.2887e-08 1.8237268647438805 1.2888e-08 1.8704716827653987 1.2889e-08 1.803422431727209 1.289e-08 1.780824739576778 1.2891e-08 1.8669465460436059 1.2892e-08 1.8698585724342995 1.2893e-08 1.8982226905991901 1.2894e-08 1.8428305966704113 1.2894999999999999e-08 1.7608316308208363 1.2896e-08 1.842216436485518 1.2897e-08 1.7415054989164396 1.2897999999999999e-08 1.8525556698261882 1.2899e-08 1.8094599257384467 1.29e-08 1.7675025075349708 1.2901e-08 1.8341979423978378 1.2902e-08 1.7857888799683153 1.2903e-08 1.7601809242880138 1.2904e-08 1.7178651512767695 1.2905e-08 1.8088462645000993 1.2906e-08 1.9111121467858578 1.2907e-08 1.8628980933791566 1.2908e-08 1.8525927765079255 1.2909e-08 1.7584866057991697 1.291e-08 1.8058192516041545 1.2910999999999999e-08 1.8451332627963062 1.2912e-08 1.8280680369176847 1.2913e-08 1.8168800796503466 1.2913999999999999e-08 1.8767532221971723 1.2915e-08 1.747563999602758 1.2916e-08 1.8174840665443113 1.2916999999999999e-08 1.752343331882369 1.2918e-08 1.8385437255592927 1.2919e-08 1.8344006169305285 1.292e-08 1.7909087038949953 1.2921e-08 1.8268911764685887 1.2922e-08 1.840302027603918 1.2923e-08 1.7555292357695285 1.2924e-08 1.837925998900033 1.2925e-08 1.757930789697178 1.2926e-08 1.7511960419780872 1.2927e-08 1.8020807338158793 1.2928e-08 1.8005357601018468 1.2929e-08 1.773470973217422 1.2929999999999999e-08 1.7949133119240201 1.2931e-08 1.816898248198227 1.2932e-08 1.8002441398707996 1.2932999999999999e-08 1.835330345712723 1.2934e-08 1.7615857246698643 1.2935e-08 1.8112439572028256 1.2935999999999999e-08 1.840538276927348 1.2937e-08 1.8265355121293807 1.2938e-08 1.8191799111407454 1.2939e-08 1.793823931195873 1.294e-08 1.7442797636240015 1.2941e-08 1.7919634234655049 1.2942e-08 1.739922734891049 1.2943e-08 1.8274268315689153 1.2944e-08 1.832258198291665 1.2945e-08 1.7247267874304701 1.2945999999999999e-08 1.7168927161400798 1.2947e-08 1.915965494608738 1.2948e-08 1.790817094677574 1.2948999999999999e-08 1.796335972690849 1.295e-08 1.7668040816498876 1.2951e-08 1.7676154653511296 1.2951999999999999e-08 1.7814414636778724 1.2953e-08 1.8238547401544045 1.2954e-08 1.8719513302032782 1.2955e-08 1.8746046205712414 1.2956e-08 1.7184331933557146 1.2957e-08 1.849367396005384 1.2958e-08 1.8179636581098633 1.2959e-08 1.7939600033643395 1.296e-08 1.8788271780347896 1.2961e-08 1.7804196462097919 1.2962e-08 1.7390377503706422 1.2963e-08 1.7353661417012447 1.2964e-08 1.8049080651373468 1.2964999999999999e-08 1.7160475634515668 1.2966e-08 1.7712977918878832 1.2967e-08 1.7003048298544545 1.2967999999999999e-08 1.8544049818827009 1.2969e-08 1.811977456611304 1.297e-08 1.7422598586011118 1.2970999999999999e-08 1.7820468152552396 1.2972e-08 1.776985396663119 1.2973e-08 1.8514633589262037 1.2974e-08 1.8762904338837252 1.2975e-08 1.7697691879936308 1.2976e-08 1.7995613539340596 1.2977e-08 1.757905422215615 1.2978e-08 1.7963174426248947 1.2979e-08 1.7745363909570218 1.298e-08 1.7231960177082346 1.2981e-08 1.8332430135022661 1.2982e-08 1.6984878149671823 1.2983e-08 1.8187819578253321 1.2983999999999999e-08 1.842092795513425 1.2985e-08 1.8067202093098707 1.2986e-08 1.8589313768201419 1.2986999999999999e-08 1.7440070666329912 1.2988e-08 1.7866173392341782 1.2989e-08 1.8032488345725326 1.299e-08 1.8456097999535075 1.2991e-08 1.7763387784466893 1.2992e-08 1.7846239970226523 1.2993e-08 1.817567168480788 1.2994e-08 1.8404427530303504 1.2995e-08 1.77434080066519 1.2996e-08 1.8217240798170202 1.2997e-08 1.8170552528231834 1.2998e-08 1.7496658072663334 1.2999e-08 1.7880132961596487 1.2999999999999999e-08 1.7703779302126328 1.3001e-08 1.7721813706383331 1.3002e-08 1.7446463584949392 1.3002999999999999e-08 1.7875940518630997 1.3004e-08 1.8589065862100647 1.3005e-08 1.849034048855025 1.3005999999999999e-08 1.8384463893354457 1.3007e-08 1.9004856279353475 1.3008e-08 1.8215819250734457 1.3009e-08 1.78341950599004 1.301e-08 1.7704657357701108 1.3011e-08 1.714429866260383 1.3012e-08 1.7965562909698816 1.3013e-08 1.8149357688942616 1.3014e-08 1.7710480020131754 1.3015e-08 1.7817123874623066 1.3016e-08 1.8457225911400932 1.3017e-08 1.7864773027357332 1.3018e-08 1.7925912885327189 1.3018999999999999e-08 1.7759596950293495 1.302e-08 1.765873946444749 1.3021e-08 1.7645148888805309 1.3021999999999999e-08 1.8503606452096526 1.3023e-08 1.6930519806825473 1.3024e-08 1.7823780084054504 1.3024999999999999e-08 1.819166635759367 1.3026e-08 1.7767580438014543 1.3027e-08 1.7760568652227375 1.3028e-08 1.79517589312762 1.3029e-08 1.796227491892574 1.303e-08 1.789837737155545 1.3031e-08 1.800738020500519 1.3032e-08 1.820481631751322 1.3033e-08 1.8903933905519148 1.3034e-08 1.7772316153209367 1.3034999999999999e-08 1.93134427519547 1.3036e-08 1.910798411589004 1.3037e-08 1.739732424144781 1.3037999999999999e-08 1.8879520533831384 1.3039e-08 1.8677890334118752 1.304e-08 1.7337600073449484 1.3040999999999999e-08 1.823375576447315 1.3042e-08 1.8306055027558799 1.3043e-08 1.8134765233005938 1.3044e-08 1.656770253075221 1.3045e-08 1.8497309669674777 1.3046e-08 1.7805907812101913 1.3047e-08 1.8858957330042652 1.3048e-08 1.7773513632689937 1.3049e-08 1.8556684864937776 1.305e-08 1.7411020827271388 1.3051e-08 1.7498268381114035 1.3052e-08 1.8061241675879478 1.3053e-08 1.7274744037032264 1.3053999999999999e-08 1.7371367301179654 1.3055e-08 1.8015582582594192 1.3056e-08 1.7773202625083115 1.3056999999999999e-08 1.8339068941329086 1.3058e-08 1.776927013586502 1.3059e-08 1.7928256441544477 1.3059999999999999e-08 1.8352384467210558 1.3061e-08 1.8160494140331476 1.3062e-08 1.7971907229913702 1.3063e-08 1.823756085183936 1.3064e-08 1.7872096786208427 1.3065e-08 1.8109092865766772 1.3066e-08 1.7851925497616667 1.3067e-08 1.7427453469455914 1.3068e-08 1.8053507395619757 1.3069e-08 1.744439421778018 1.3069999999999999e-08 1.821421610149605 1.3071e-08 1.8127125857126236 1.3072e-08 1.8204692268526956 1.3072999999999999e-08 1.8266002180006493 1.3074e-08 1.7459322629870402 1.3075e-08 1.7807747639247362 1.3075999999999999e-08 1.7059474306823743 1.3077e-08 1.754555380754832 1.3078e-08 1.7910568916015301 1.3079e-08 1.8449133814187633 1.308e-08 1.753794667337766 1.3081e-08 1.8274589324432422 1.3082e-08 1.831930929778575 1.3083e-08 1.904385452692315 1.3084e-08 1.8182658681169315 1.3085e-08 1.8344222547406321 1.3086e-08 1.8543868843193987 1.3087e-08 1.7637727100743057 1.3088e-08 1.8193732484112983 1.3088999999999999e-08 1.76715950027841 1.309e-08 1.862116979617571 1.3091e-08 1.78229831238673 1.3091999999999999e-08 1.7614056081013705 1.3093e-08 1.8119304802321334 1.3094e-08 1.7832427331655014 1.3094999999999999e-08 1.8824232458704155 1.3096e-08 1.8302891551392175 1.3097e-08 1.759504157598024 1.3098e-08 1.799077755025812 1.3099e-08 1.8329440345725148 1.31e-08 1.8257180479855692 1.3101e-08 1.9008986018260698 1.3102e-08 1.819862891546592 1.3103e-08 1.7569704265089814 1.3104e-08 1.8313304129490475 1.3105e-08 1.7676129942302994 1.3106e-08 1.7579756753315012 1.3107e-08 1.8023112774529348 1.3107999999999999e-08 1.7182776961385833 1.3109e-08 1.8228511547321429 1.311e-08 1.8469590221495347 1.3110999999999999e-08 1.8196535273665864 1.3112e-08 1.826563372487162 1.3113e-08 1.8195443461637686 1.3114e-08 1.8584433493172745 1.3115e-08 1.7448110497763683 1.3116e-08 1.8180413959437198 1.3117e-08 1.7737576492816014 1.3118e-08 1.813385170994434 1.3119e-08 1.8365342713284911 1.312e-08 1.871405034102578 1.3121e-08 1.8048347407241807 1.3122e-08 1.7537143260943417 1.3123e-08 1.7921466546630571 1.3123999999999999e-08 1.7825904671138564 1.3125e-08 1.8410295291525454 1.3126e-08 1.7781703459039566 1.3126999999999999e-08 1.8608372730275717 1.3128e-08 1.7179393866820358 1.3129e-08 1.8251706516442554 1.3129999999999999e-08 1.804087176260268 1.3131e-08 1.9212092167774533 1.3132e-08 1.80896181842452 1.3133e-08 1.768267407697422 1.3134e-08 1.7669553087317806 1.3135e-08 1.7457079797403816 1.3136e-08 1.717065796655438 1.3137e-08 1.804444212243809 1.3138e-08 1.7920229488014563 1.3139e-08 1.8108155018374046 1.314e-08 1.8070827228183608 1.3141e-08 1.7303986579499504 1.3142e-08 1.794737365534823 1.3142999999999999e-08 1.8296023154746663 1.3144e-08 1.8359431003991318 1.3145e-08 1.7720285093947232 1.3145999999999999e-08 1.7039378176241158 1.3147e-08 1.7782435204021216 1.3148e-08 1.877061226043153 1.3148999999999999e-08 1.8254346647002004 1.315e-08 1.7895207765542098 1.3151e-08 1.768676239864418 1.3152e-08 1.7438336923665645 1.3153e-08 1.7067238175427215 1.3154e-08 1.7785446274922592 1.3155e-08 1.8170816797203138 1.3156e-08 1.8742170308862978 1.3157e-08 1.7462457577335557 1.3158e-08 1.8838143928571758 1.3158999999999999e-08 1.785744370971029 1.316e-08 1.7539196670666435 1.3161e-08 1.804279529886376 1.3161999999999999e-08 1.8442199588631882 1.3163e-08 1.7947663784368582 1.3164e-08 1.8618122290816903 1.3164999999999999e-08 1.7475541936521228 1.3166e-08 1.8609159165447482 1.3167e-08 1.7492709918930711 1.3168e-08 1.8600833836305608 1.3169e-08 1.9279598596313516 1.317e-08 1.7779832267584044 1.3171e-08 1.8869091576352055 1.3172e-08 1.8124766882727865 1.3173e-08 1.7260477822596931 1.3174e-08 1.7990225429167195 1.3175e-08 1.8207319176883798 1.3176e-08 1.7938623356154448 1.3177e-08 1.8427114605696329 1.3177999999999999e-08 1.900294971791395 1.3179e-08 1.8265492984481932 1.318e-08 1.874420374159253 1.3180999999999999e-08 1.7739035403595964 1.3182e-08 1.7455892774422666 1.3183e-08 1.7783332792910884 1.3183999999999999e-08 1.7923106231821733 1.3185e-08 1.8414742400886814 1.3186e-08 1.8016618041235 1.3187e-08 1.78201152820153 1.3188e-08 1.7643495098093671 1.3189e-08 1.8869018547061243 1.319e-08 1.7484866295055945 1.3191e-08 1.7833106824053226 1.3192e-08 1.7932204441853814 1.3193e-08 1.8516014584938418 1.3194e-08 1.7817611638720674 1.3195e-08 1.8275750594875273 1.3196e-08 1.869274295687055 1.3196999999999999e-08 1.7483143861541028 1.3198e-08 1.6905836786369781 1.3199e-08 1.8053919723544936 1.3199999999999999e-08 1.8542285715012499 1.3201e-08 1.7828594821823855 1.3202e-08 1.7352397634264187 1.3203e-08 1.7552537082003972 1.3204e-08 1.8698595871182773 1.3205e-08 1.7926208097312342 1.3206e-08 1.7758494042576325 1.3207e-08 1.8498732354879204 1.3208e-08 1.7849078085115366 1.3209e-08 1.773508487178813 1.321e-08 1.7605719422214117 1.3211e-08 1.8454269385897668 1.3212e-08 1.9527972415675603 1.3212999999999999e-08 1.7628812183419829 1.3214e-08 1.8396916845621347 1.3215e-08 1.7525027083125038 1.3215999999999999e-08 1.7827821438274982 1.3217e-08 1.8244788337171345 1.3218e-08 1.8408900977504223 1.3218999999999999e-08 1.7226311965485213 1.322e-08 1.8271740000303685 1.3221e-08 1.8333590395985975 1.3222e-08 1.7519936374114113 1.3223e-08 1.878847399606351 1.3224e-08 1.8427077255452506 1.3225e-08 1.7315315497144668 1.3226e-08 1.7994817701045471 1.3227e-08 1.7790388628872942 1.3228e-08 1.7922677211987297 1.3229e-08 1.7414107224268183 1.323e-08 1.8631984964075323 1.3231e-08 1.7755948835777113 1.3231999999999999e-08 1.8474231739695075 1.3233e-08 1.767963020872645 1.3234e-08 1.8563674612510868 1.3234999999999999e-08 1.788696014964959 1.3236e-08 1.7764982132064961 1.3237e-08 1.8610040243761479 1.3237999999999999e-08 1.7232147251397312 1.3239e-08 1.8253169459812024 1.324e-08 1.739135797345794 1.3241e-08 1.8039906040775506 1.3242e-08 1.7873673254768263 1.3243e-08 1.861775860054131 1.3244e-08 1.849558825419973 1.3245e-08 1.8744682291344663 1.3246e-08 1.8405005172064937 1.3247e-08 1.7869225160211815 1.3247999999999999e-08 1.8785586751493493 1.3249e-08 1.7369308643550385 1.325e-08 1.7649462335632289 1.3250999999999999e-08 1.851547144989671 1.3252e-08 1.771938682175235 1.3253e-08 1.7846790316955348 1.3253999999999999e-08 1.7198337112688582 1.3255e-08 1.8346656637515533 1.3256e-08 1.845494603128821 1.3257e-08 1.7992371942627106 1.3258e-08 1.6937709102047513 1.3259e-08 1.7962906740641376 1.326e-08 1.7642712427990157 1.3261e-08 1.7589710226455102 1.3262e-08 1.7853590171124274 1.3263e-08 1.7823363354666322 1.3264e-08 1.8176453151877254 1.3265e-08 1.6807327413509459 1.3266e-08 1.8919064155531504 1.3266999999999999e-08 1.71676404115577 1.3268e-08 1.8270003495844003 1.3269e-08 1.8009827750348535 1.3269999999999999e-08 1.7637958195360404 1.3271e-08 1.7825218956589983 1.3272e-08 1.7998934194805998 1.3272999999999999e-08 1.795509551032406 1.3274e-08 1.850940368158755 1.3275e-08 1.7658732101594021 1.3276e-08 1.7392238662905264 1.3277e-08 1.829919812049234 1.3278e-08 1.7122662571629823 1.3279e-08 1.7826262730897389 1.328e-08 1.8127523580742169 1.3281e-08 1.8505320830556136 1.3282e-08 1.7788186784985678 1.3283e-08 1.7419916313318151 1.3284e-08 1.7035050823599474 1.3285e-08 1.7986170854627266 1.3285999999999999e-08 1.7540559702498137 1.3287e-08 1.7514368079673297 1.3288e-08 1.7536706332725704 1.3288999999999999e-08 1.7980151317739903 1.329e-08 1.8074163821418532 1.3291e-08 1.7447528088854196 1.3292e-08 1.8381557608375194 1.3293e-08 1.8439676622871817 1.3294e-08 1.7623571001699518 1.3295e-08 1.7749033599628157 1.3296e-08 1.7077025904557523 1.3297e-08 1.8620916637888802 1.3298e-08 1.7353187770981606 1.3299e-08 1.8089385554417747 1.33e-08 1.7873724690820085 1.3301e-08 1.7676742116639097 1.3301999999999999e-08 1.7834143312575153 1.3303e-08 1.7929680533319463 1.3304e-08 1.8772150805657435 1.3304999999999999e-08 1.7671753470209217 1.3306e-08 1.8327971143966693 1.3307e-08 1.9080952789616765 1.3307999999999999e-08 1.8225338789841268 1.3309e-08 1.78994580182697 1.331e-08 1.8313357847625538 1.3311e-08 1.7872099437597335 1.3312e-08 1.8151708425480202 1.3313e-08 1.802074681677914 1.3314e-08 1.8073465478559414 1.3315e-08 1.7535499286576097 1.3316e-08 1.8151799289622383 1.3317e-08 1.8447347165809704 1.3318e-08 1.800686124989437 1.3319e-08 1.7946259917817529 1.332e-08 1.8337792055718445 1.3320999999999999e-08 1.7321390940438277 1.3322e-08 1.8423113058198188 1.3323e-08 1.7549794602462112 1.3323999999999999e-08 1.851494276897079 1.3325e-08 1.8346727744810103 1.3326e-08 1.8292482154473266 1.3326999999999999e-08 1.7746563820139387 1.3328e-08 1.7756519986604793 1.3329e-08 1.8568788680980468 1.333e-08 1.7520992986954638 1.3331e-08 1.7002776719578048 1.3332e-08 1.7938643291716485 1.3333e-08 1.8109117520135045 1.3334e-08 1.730332102241558 1.3335e-08 1.8688857774826662 1.3336e-08 1.8193181044846336 1.3336999999999999e-08 1.8008303584704242 1.3338e-08 1.844102398112514 1.3339e-08 1.70082742506162 1.3339999999999999e-08 1.74750464826672 1.3341e-08 1.8169694066103685 1.3342e-08 1.769748822972115 1.3342999999999999e-08 1.8770965999632327 1.3344e-08 1.8049605378632412 1.3345e-08 1.9393671110478665 1.3346e-08 1.723972178553257 1.3347e-08 1.868645391431961 1.3348e-08 1.7649116695068747 1.3349e-08 1.7462727023882583 1.335e-08 1.758870197956713 1.3351e-08 1.8612589853010464 1.3352e-08 1.7890437210206758 1.3353e-08 1.8326459534256034 1.3354e-08 1.7877230996508329 1.3355e-08 1.7881780270774357 1.3355999999999999e-08 1.8087165831346406 1.3357e-08 1.759014151259522 1.3358e-08 1.8038135134417195 1.3358999999999999e-08 1.7102862305335949 1.336e-08 1.8205495497757314 1.3361e-08 1.8138393559594725 1.3361999999999999e-08 1.7670360799997433 1.3363e-08 1.751819738011939 1.3364e-08 1.778864716574957 1.3365e-08 1.8578998658522563 1.3366e-08 1.8645807466973006 1.3367e-08 1.8034993020948902 1.3368e-08 1.8147219069973788 1.3369e-08 1.780569162167239 1.337e-08 1.8529173428607868 1.3371e-08 1.8072112458250107 1.3371999999999999e-08 1.8373022541389703 1.3373e-08 1.7951110333859561 1.3374e-08 1.789874475456003 1.3374999999999999e-08 1.8605312301218584 1.3376e-08 1.8072465625413743 1.3377e-08 1.7441152484343287 1.3377999999999999e-08 1.8292761957129773 1.3379e-08 1.7668014314785525 1.338e-08 1.7486442166623597 1.3381e-08 1.8046606122296707 1.3382e-08 1.8220231935985016 1.3383e-08 1.8429447492179303 1.3384e-08 1.8802920760213206 1.3385e-08 1.7391878887429704 1.3386e-08 1.8495212683591808 1.3387e-08 1.7275278842544535 1.3388e-08 1.779906455265586 1.3389e-08 1.7563415429355966 1.339e-08 1.8318071625146348 1.3390999999999999e-08 1.8565593911451057 1.3392e-08 1.8115183803981085 1.3393e-08 1.848779625671589 1.3393999999999999e-08 1.8134228984272704 1.3395e-08 1.9034258084747673 1.3396e-08 1.8054747951220889 1.3396999999999999e-08 1.7585064698751438 1.3398e-08 1.853239937179713 1.3399e-08 1.8193539226216846 1.34e-08 1.844174487464897 1.3401e-08 1.7062549695027263 1.3402e-08 1.774153832643196 1.3403e-08 1.679310387461413 1.3404e-08 1.7544996811559808 1.3405e-08 1.791090377162509 1.3406e-08 1.9457163027420372 1.3407e-08 1.8410278121945758 1.3408e-08 1.8240181688954116 1.3409e-08 1.811034666986357 1.3409999999999999e-08 1.8464145066944717 1.3411e-08 1.8553455392699847 1.3412e-08 1.8692157857184741 1.3412999999999999e-08 1.827697559767645 1.3414e-08 1.7452767291969586 1.3415e-08 1.7715211633808112 1.3415999999999999e-08 1.7787555311503283 1.3417e-08 1.8761782334247643 1.3418e-08 1.7768297796966042 1.3419e-08 1.7750926114913108 1.342e-08 1.8156428348128342 1.3421e-08 1.7786446639629518 1.3422e-08 1.6963921599467102 1.3423e-08 1.667593932338416 1.3424e-08 1.7678009725434214 1.3425e-08 1.81334000077174 1.3425999999999999e-08 1.7271753416242226 1.3427e-08 1.7743411980977346 1.3428e-08 1.7889656701471823 1.3428999999999999e-08 1.7578443785173974 1.343e-08 1.7580328442320936 1.3431e-08 1.8051066296440816 1.3431999999999999e-08 1.7071311953711317 1.3433e-08 1.8074763993964718 1.3434e-08 1.8274612706141695 1.3435e-08 1.8105744852663943 1.3436e-08 1.8278368180433173 1.3437e-08 1.8649737612520834 1.3438e-08 1.8222807220410837 1.3439e-08 1.7894488215098756 1.344e-08 1.8601756235782725 1.3441e-08 1.7907644024652705 1.3442e-08 1.8299093093697223 1.3443e-08 1.726052887743168 1.3444e-08 1.7431055387611356 1.3444999999999999e-08 1.7574153956292426 1.3446e-08 1.8894788905735094 1.3447e-08 1.82755356391909 1.3447999999999999e-08 1.8202644155652745 1.3449e-08 1.7774596371632847 1.345e-08 1.7614249425948798 1.3450999999999999e-08 1.7485956594978933 1.3452e-08 1.8192993888314637 1.3453e-08 1.7383832636716032 1.3454e-08 1.780566804213133 1.3455e-08 1.7112593113206394 1.3456e-08 1.7550144919696131 1.3457e-08 1.8398996514653934 1.3458e-08 1.7825060138590625 1.3459e-08 1.7429317534271154 1.346e-08 1.7124729618173562 1.3460999999999999e-08 1.7683929246427137 1.3462e-08 1.8281396975379647 1.3463e-08 1.8126496179905667 1.3463999999999999e-08 1.7829241888170915 1.3465e-08 1.7753766870009609 1.3466e-08 1.8115137403744839 1.3466999999999999e-08 1.7195580788155425 1.3468e-08 1.8479134966441566 1.3469e-08 1.7110631542579435 1.347e-08 1.8253087041796914 1.3471e-08 1.7902216734221397 1.3472e-08 1.8245437333769816 1.3473e-08 1.8338308105535488 1.3474e-08 1.6580633291851983 1.3475e-08 1.784185579404993 1.3476e-08 1.7872204872226036 1.3477e-08 1.7296714299864195 1.3478e-08 1.8189483558825752 1.3479e-08 1.847393870231013 1.3479999999999999e-08 1.822508179003412 1.3481e-08 1.854737094817651 1.3482e-08 1.838937337387045 1.3482999999999999e-08 1.6509164754281538 1.3484e-08 1.841640294569725 1.3485e-08 1.6846866330829235 1.3485999999999999e-08 1.7366633288395863 1.3487e-08 1.832649618531016 1.3488e-08 1.8452849798697557 1.3489e-08 1.7300505519439948 1.349e-08 1.721070728748714 1.3491e-08 1.7939844837662065 1.3492e-08 1.8101898342901355 1.3493e-08 1.7240899452402738 1.3494e-08 1.8157376325824055 1.3495e-08 1.7864646131579336 1.3496e-08 1.8449471697305544 1.3497e-08 1.8116035053620894 1.3498e-08 1.7920252219461508 1.3498999999999999e-08 1.8775085180278015 1.35e-08 1.9213050579128728 1.3501e-08 1.7168870316990585 1.3501999999999999e-08 1.7856160454674634 1.3503e-08 1.848509465476595 1.3504e-08 1.7743571178192925 1.3504999999999999e-08 1.774343165495587 1.3506e-08 1.8629893128098427 1.3507e-08 1.8195580248855328 1.3508e-08 1.8232937525320478 1.3509e-08 1.759842987344835 1.351e-08 1.8107829462214122 1.3511e-08 1.8637101969821062 1.3512e-08 1.8823805054999556 1.3513e-08 1.7806281073953443 1.3514e-08 1.7738715165507577 1.3514999999999999e-08 1.8600268441429604 1.3516e-08 1.7962838102704934 1.3517e-08 1.8031976157751597 1.3517999999999999e-08 1.8280973843467099 1.3519e-08 1.813248990572155 1.352e-08 1.798906841051707 1.3520999999999999e-08 1.8084548597322834 1.3522e-08 1.8102450640612453 1.3523e-08 1.6743675743077675 1.3524e-08 1.8123942502133994 1.3525e-08 1.819350074358515 1.3526e-08 1.8003195252118664 1.3527e-08 1.769075968424441 1.3528e-08 1.7538508087398028 1.3529e-08 1.8588680764041077 1.353e-08 1.8248691468111222 1.3531e-08 1.7330072277608164 1.3532e-08 1.8242798183969182 1.3533e-08 1.7899837646876549 1.3533999999999999e-08 1.7683456399564914 1.3535e-08 1.819877693113365 1.3536e-08 1.7761037976407532 1.3536999999999999e-08 1.7395926958641768 1.3538e-08 1.7749414287218088 1.3539e-08 1.8181139264122015 1.3539999999999999e-08 1.8599873447826512 1.3541e-08 1.8346288744105825 1.3542e-08 1.7367076975757554 1.3543e-08 1.7585819485033332 1.3544e-08 1.8107933433383707 1.3545e-08 1.7203540811962106 1.3546e-08 1.7945648343555316 1.3547e-08 1.8020337017316663 1.3548e-08 1.837081712163377 1.3549e-08 1.7693707683975977 1.3549999999999999e-08 1.7818626380028908 1.3551e-08 1.7665661003843909 1.3552e-08 1.828586658697456 1.3552999999999999e-08 1.776234211405427 1.3554e-08 1.820327739560544 1.3555e-08 1.7986425213525759 1.3555999999999999e-08 1.7721835073544927 1.3557e-08 1.8037504826255095 1.3558e-08 1.8244092225356319 1.3559e-08 1.8145520528132542 1.356e-08 1.8417998575081436 1.3561e-08 1.789123445010105 1.3562e-08 1.8180936061197057 1.3563e-08 1.678146222176939 1.3564e-08 1.7723533913988296 1.3565e-08 1.7898709530111812 1.3566e-08 1.692211445232447 1.3567e-08 1.77944452187989 1.3568e-08 1.7600749920792993 1.3568999999999999e-08 1.7838965106998412 1.357e-08 1.774100064994803 1.3571e-08 1.9043163659189526 1.3571999999999999e-08 1.7869924647158035 1.3573e-08 1.861608774675727 1.3574e-08 1.752700622387619 1.3574999999999999e-08 1.7408940130960266 1.3576e-08 1.7750862029034764 1.3577e-08 1.7979265833631053 1.3578e-08 1.8226156453631388 1.3579e-08 1.8137447484256568 1.358e-08 1.8899458505135684 1.3581e-08 1.8292679413633557 1.3582e-08 1.8023978645374295 1.3583e-08 1.7715982014377276 1.3584e-08 1.8637404394934034 1.3585e-08 1.8175300916760149 1.3586e-08 1.8268470026591128 1.3587e-08 1.7857011381954648 1.3587999999999999e-08 1.7870012823837846 1.3589e-08 1.7449320077324069 1.359e-08 1.7656160693363314 1.3590999999999999e-08 1.8276364434922039 1.3592e-08 1.699841987874087 1.3593e-08 1.780427047554737 1.3593999999999999e-08 1.834094161222132 1.3595e-08 1.8115110761701514 1.3596e-08 1.7983083659281034 1.3597e-08 1.8199087149664428 1.3598e-08 1.8873042992336126 1.3599e-08 1.8021207292254442 1.36e-08 1.8018193822267 1.3601e-08 1.8219950513851821 1.3602e-08 1.7528188026503253 1.3603e-08 1.8227830747410134 1.3603999999999999e-08 1.7653910650866218 1.3605e-08 1.8997718606863443 1.3606e-08 1.7568730456541573 1.3606999999999999e-08 1.8282736736824474 1.3608e-08 1.8522184535700892 1.3609e-08 1.7013589032951966 1.3609999999999999e-08 1.7617291264334791 1.3611e-08 1.8570248800878417 1.3612e-08 1.865621389515996 1.3613e-08 1.733452524571243 1.3614e-08 1.772332867873254 1.3615e-08 1.8190755082063288 1.3616e-08 1.806416220811815 1.3617e-08 1.7251298126371455 1.3618e-08 1.768136657622887 1.3619e-08 1.845037661589167 1.362e-08 1.8310927683087244 1.3621e-08 1.7653898743678613 1.3622e-08 1.8192162142758521 1.3622999999999999e-08 1.7858061365358666 1.3624e-08 1.80222791851791 1.3625e-08 1.7566292464328932 1.3625999999999999e-08 1.7880897755929352 1.3627e-08 1.7396523513599726 1.3628e-08 1.7872498415742086 1.3628999999999999e-08 1.8260164687923424 1.363e-08 1.7744207689818596 1.3631e-08 1.82763574084429 1.3632e-08 1.7484852920250535 1.3633e-08 1.7365669036400846 1.3634e-08 1.8566137147243633 1.3635e-08 1.7437231093386303 1.3636e-08 1.7609829086307844 1.3637e-08 1.8340578932788034 1.3638e-08 1.8468052154682526 1.3638999999999999e-08 1.7940556780386239 1.364e-08 1.8917482604035114 1.3641e-08 1.8132532864338544 1.3641999999999999e-08 1.7520732611063319 1.3643e-08 1.721150946973796 1.3644e-08 1.851974706934599 1.3644999999999999e-08 1.7642851793137146 1.3646e-08 1.8072436140315582 1.3647e-08 1.8697748830552587 1.3648e-08 1.7296161188861963 1.3649e-08 1.777184874004505 1.365e-08 1.905547254310102 1.3651e-08 1.7540829129271815 1.3652e-08 1.7711315367727087 1.3653e-08 1.7792817969849046 1.3654e-08 1.78047241069527 1.3655e-08 1.709348615744025 1.3656e-08 1.8780124826349793 1.3657e-08 1.8519786644396805 1.3657999999999999e-08 1.7262086946373751 1.3659e-08 1.807111137101101 1.366e-08 1.8632724796409228 1.3660999999999999e-08 1.7981209106511435 1.3662e-08 1.7411008635157632 1.3663e-08 1.722823497652938 1.3663999999999999e-08 1.7913994389910841 1.3665e-08 1.76589107565545 1.3666e-08 1.708594794101813 1.3667e-08 1.7616328903257763 1.3668e-08 1.8359594391022256 1.3669e-08 1.8676335887204618 1.367e-08 1.7442337438073223 1.3671e-08 1.7654113169517716 1.3672e-08 1.854677967124353 1.3673e-08 1.756671097720145 1.3674e-08 1.7310750396102863 1.3675e-08 1.8380669596817234 1.3676e-08 1.7511723043200178 1.3676999999999999e-08 1.7349080818216986 1.3678e-08 1.76584643158733 1.3679e-08 1.7857569129196988 1.3679999999999999e-08 1.7593712764168619 1.3681e-08 1.8303698326526094 1.3682e-08 1.8022853998568449 1.3683e-08 1.7398177926838456 1.3684e-08 1.7748458899407944 1.3685e-08 1.760581001201858 1.3686e-08 1.8290756133116524 1.3687e-08 1.746416834954687 1.3688e-08 1.7422201148002532 1.3689e-08 1.7846187996520728 1.369e-08 1.8128327391215708 1.3691e-08 1.7485570056612245 1.3692e-08 1.8603161128586998 1.3692999999999999e-08 1.7615001106982735 1.3694e-08 1.8187648624973525 1.3695e-08 1.7577964663944217 1.3695999999999999e-08 1.8311669211540997 1.3697e-08 1.8401831205977912 1.3698e-08 1.9129822676126333 1.3698999999999999e-08 1.7669918370101987 1.37e-08 1.7935115119435827 1.3701e-08 1.8307236098631123 1.3702e-08 1.8361408545989 1.3703e-08 1.839491168647664 1.3704e-08 1.847975581853805 1.3705e-08 1.827556503642675 1.3706e-08 1.8252205687392815 1.3707e-08 1.7805860828128808 1.3708e-08 1.7817402425723596 1.3709e-08 1.765757956124359 1.371e-08 1.791811145849682 1.3711e-08 1.798722854122758 1.3711999999999999e-08 1.8068197038315068 1.3713e-08 1.709924016641283 1.3714e-08 1.851623639937654 1.3714999999999999e-08 1.8844178862900698 1.3716e-08 1.712556661162416 1.3717e-08 1.8488898462780916 1.3717999999999999e-08 1.7259121608771293 1.3719e-08 1.7961857670695245 1.372e-08 1.783511899423214 1.3721e-08 1.7947129564274293 1.3722e-08 1.822124970039415 1.3723e-08 1.8121011558497035 1.3724e-08 1.7559044483064858 1.3725e-08 1.8284944372422347 1.3726e-08 1.8461034111518713 1.3727e-08 1.7526577401598513 1.3727999999999999e-08 1.7889355369579893 1.3729e-08 1.7199405475363196 1.373e-08 1.799927813294711 1.3730999999999999e-08 1.9357510110424698 1.3732e-08 1.7792899516977683 1.3733e-08 1.7620256593530035 1.3733999999999999e-08 1.7554654051908731 1.3735e-08 1.8716253166419747 1.3736e-08 1.817416296377559 1.3737e-08 1.845644606119108 1.3738e-08 1.6869583036926457 1.3739e-08 1.868562856943721 1.374e-08 1.7857552300034927 1.3741e-08 1.7248364916604582 1.3742e-08 1.7571431428003383 1.3743e-08 1.747097435002765 1.3744e-08 1.8096408644792823 1.3745e-08 1.8637053683595577 1.3746e-08 1.7695193720001672 1.3746999999999999e-08 1.7811825636953436 1.3748e-08 1.844363357237002 1.3749e-08 1.7434113732552936 1.3749999999999999e-08 1.7888315831684805 1.3751e-08 1.8528171804284248 1.3752e-08 1.7862751620238124 1.3752999999999999e-08 1.8527167449979443 1.3754e-08 1.791771914784647 1.3755e-08 1.7739937054201191 1.3756e-08 1.752203057206913 1.3757e-08 1.7836840232272388 1.3758e-08 1.7969002989850007 1.3759e-08 1.8623623723368197 1.376e-08 1.7833774941224418 1.3761e-08 1.8148296558782093 1.3762e-08 1.841279126895167 1.3762999999999999e-08 1.7752181784950183 1.3764e-08 1.7996579097008374 1.3765e-08 1.8487773261519718 1.3765999999999999e-08 1.7698495609108482 1.3767e-08 1.8100873856633017 1.3768e-08 1.7699667394657168 1.3768999999999999e-08 1.7628093339704085 1.377e-08 1.8563653984824846 1.3771e-08 1.7970607448215103 1.3772e-08 1.7760570225772727 1.3773e-08 1.8402529867559727 1.3774e-08 1.8593427232387614 1.3775e-08 1.8113161717959618 1.3776e-08 1.7833075417263937 1.3777e-08 1.7733991875887118 1.3778e-08 1.8087359854552125 1.3779e-08 1.813772146727596 1.378e-08 1.8483415937688528 1.3781e-08 1.7548038366956775 1.3781999999999999e-08 1.8538120233845412 1.3783e-08 1.8093609175657823 1.3784e-08 1.7431085394002257 1.3784999999999999e-08 1.7530180752869984 1.3786e-08 1.8126649214485824 1.3787e-08 1.7121889677943831 1.3787999999999999e-08 1.880070048914616 1.3789e-08 1.8270741013588743 1.379e-08 1.7474342998417958 1.3791e-08 1.9073806871283228 1.3792e-08 1.7722866396874506 1.3793e-08 1.7251091679715354 1.3794e-08 1.7785089210339453 1.3795e-08 1.8607764113613614 1.3796e-08 1.749340782356785 1.3797e-08 1.857116336299049 1.3798e-08 1.8402557555294068 1.3799e-08 1.7617657727053315 1.38e-08 1.7185466187503966 1.3800999999999999e-08 1.7183564163570892 1.3802e-08 1.9042573016416204 1.3803e-08 1.6738052466374602 1.3803999999999999e-08 1.7663620536958569 1.3805e-08 1.7499554562050315 1.3806e-08 1.7980590871026425 1.3806999999999999e-08 1.7433374779460653 1.3808e-08 1.742799080238406 1.3809e-08 1.799610684221907 1.381e-08 1.816939359358315 1.3811e-08 1.801267128146937 1.3812e-08 1.8040521839842947 1.3813e-08 1.7987759852774907 1.3814e-08 1.7935853321010142 1.3815e-08 1.799823708578017 1.3816e-08 1.749660506460006 1.3816999999999999e-08 1.8740954694385856 1.3818e-08 1.9174078757505233 1.3819e-08 1.75141384405811 1.3819999999999999e-08 1.8781721714125057 1.3821e-08 1.8473660123088118 1.3822e-08 1.801521930288555 1.3822999999999999e-08 1.8449961168823705 1.3824e-08 1.8587660440662015 1.3825e-08 1.7891289259230487 1.3826e-08 1.7707612917398576 1.3827e-08 1.8286787991483577 1.3828e-08 1.7782212041406935 1.3829e-08 1.7869725858716352 1.383e-08 1.811840933115607 1.3831e-08 1.8239751499028543 1.3832e-08 1.826757943482412 1.3833e-08 1.7189384381040855 1.3834e-08 1.7640413057947477 1.3835e-08 1.6720926421190994 1.3835999999999999e-08 1.7241947428246127 1.3837e-08 1.8824961457414733 1.3838e-08 1.7462648100949003 1.3838999999999999e-08 1.7431862793203405 1.384e-08 1.8516892048732012 1.3841e-08 1.821165214837637 1.3841999999999999e-08 1.712200986145231 1.3843e-08 1.803199394824227 1.3844e-08 1.7558521870377357 1.3845e-08 1.7648837464006313 1.3846e-08 1.7622486828555874 1.3847e-08 1.7841445977461838 1.3848e-08 1.8361795983554552 1.3849e-08 1.8024135203988378 1.385e-08 1.8184941894184976 1.3851e-08 1.8498683863512069 1.3851999999999999e-08 1.8143497947626233 1.3853e-08 1.7237696360005572 1.3854e-08 1.8670467785846836 1.3854999999999999e-08 1.7612945647515488 1.3856e-08 1.7172571684996987 1.3857e-08 1.8040386615384265 1.3857999999999999e-08 1.781815964418342 1.3859e-08 1.7628662064479044 1.386e-08 1.7272869073869654 1.3861e-08 1.8029735521413404 1.3862e-08 1.7091679405877722 1.3863e-08 1.6653278196018344 1.3864e-08 1.7207814749840054 1.3865e-08 1.810685523053958 1.3866e-08 1.7843529881901083 1.3867e-08 1.7813472857460941 1.3868e-08 1.7276528233639112 1.3869e-08 1.8306038361581929 1.387e-08 1.7658988108792744 1.3870999999999999e-08 1.7837600485960714 1.3872e-08 1.768635746516307 1.3873e-08 1.697781229892936 1.3873999999999999e-08 1.9021946204745392 1.3875e-08 1.7469283049219697 1.3876e-08 1.7510288038162907 1.3876999999999999e-08 1.7709022986217273 1.3878e-08 1.765252167577479 1.3879e-08 1.7423004922440604 1.388e-08 1.808580388401773 1.3881e-08 1.7137811784150243 1.3882e-08 1.7005535355189931 1.3883e-08 1.8518056000242438 1.3884e-08 1.8287054815935002 1.3885e-08 1.7762911040005354 1.3886e-08 1.7936432233353952 1.3887e-08 1.8035223737272967 1.3888e-08 1.7355885245362164 1.3889e-08 1.8430534735130326 1.3889999999999999e-08 1.7668627635929768 1.3891e-08 1.822824076288682 1.3892e-08 1.8002725483569308 1.3892999999999999e-08 1.7349720159775384 1.3894e-08 1.7850450784863403 1.3895e-08 1.848459500273239 1.3895999999999999e-08 1.7776357075442628 1.3897e-08 1.716175026410856 1.3898e-08 1.7737825607464734 1.3899e-08 1.8461749205488713 1.39e-08 1.838179563866688 1.3901e-08 1.770143790799516 1.3902e-08 1.8266969435025813 1.3903e-08 1.8570756927565812 1.3904e-08 1.839642274069019 1.3905e-08 1.908308994694679 1.3905999999999999e-08 1.8429918024061778 1.3907e-08 1.8095787014526217 1.3908e-08 1.7956737646510659 1.3908999999999999e-08 1.8204276554420773 1.391e-08 1.784965172089709 1.3911e-08 1.8839040421906006 1.3911999999999999e-08 1.7635993272739334 1.3913e-08 1.7903380378040508 1.3914e-08 1.8056143654774304 1.3915e-08 1.89350634633566 1.3916e-08 1.7902875060458519 1.3917e-08 1.7727291169519759 1.3918e-08 1.6994470262754622 1.3919e-08 1.8600942070377937 1.392e-08 1.8713333729465447 1.3921e-08 1.804880128672399 1.3922e-08 1.8170144231161045 1.3923e-08 1.8812374527943072 1.3924e-08 1.7066759348504412 1.3924999999999999e-08 1.8638493989877174 1.3926e-08 1.7659688068505657 1.3927e-08 1.8349758469600512 1.3927999999999999e-08 1.7802540714106878 1.3929e-08 1.8425037079432394 1.393e-08 1.8367685994281164 1.3930999999999999e-08 1.8392713631660305 1.3932e-08 1.771475007942998 1.3933e-08 1.8745533038815132 1.3934e-08 1.8160686883845263 1.3935e-08 1.7455069280074096 1.3936e-08 1.7861769109282934 1.3937e-08 1.7846911465586972 1.3938e-08 1.7201214491027075 1.3939e-08 1.823410684588104 1.394e-08 1.7295537781263213 1.3940999999999999e-08 1.778709523717097 1.3942e-08 1.7567749397186732 1.3943e-08 1.7899050961142666 1.3943999999999999e-08 1.8001555882375857 1.3945e-08 1.7652736223799605 1.3946e-08 1.7718887493962932 1.3946999999999999e-08 1.8531956253844082 1.3948e-08 1.77318038338522 1.3949e-08 1.7529473714158923 1.395e-08 1.7838050548773623 1.3951e-08 1.8806645418859296 1.3952e-08 1.813503160272458 1.3953e-08 1.7673714670963463 1.3954e-08 1.8197413734727201 1.3955e-08 1.713208490680772 1.3956e-08 1.8935104140077696 1.3957e-08 1.8415141564606998 1.3958e-08 1.8018020217239523 1.3959e-08 1.8139407110393269 1.3959999999999999e-08 1.8476157726010278 1.3961e-08 1.8156006257218205 1.3962e-08 1.718163171213986 1.3962999999999999e-08 1.7016368257934285 1.3964e-08 1.8104837141588417 1.3965e-08 1.837992136303111 1.3965999999999999e-08 1.8042694670347643 1.3967e-08 1.8175870593741856 1.3968e-08 1.7839739148836278 1.3969e-08 1.798997212385311 1.397e-08 1.8411501133373658 1.3971e-08 1.867293589945421 1.3972e-08 1.80999209314973 1.3973e-08 1.8495530225092465 1.3974e-08 1.7803929044624542 1.3975e-08 1.8255502631947214 1.3976e-08 1.751248010489686 1.3977e-08 1.8168187339912807 1.3978e-08 1.8390806448782993 1.3978999999999999e-08 1.7364544445676842 1.398e-08 1.865964516520093 1.3981e-08 1.8407909673000422 1.3981999999999999e-08 1.7237505991053794 1.3983e-08 1.884945933502388 1.3984e-08 1.7866045358507254 1.3984999999999999e-08 1.831652458918721 1.3986e-08 1.7958294805287072 1.3987e-08 1.9557559603710588 1.3988e-08 1.7686655445110397 1.3989e-08 1.9221895211364852 1.399e-08 1.7655998862528672 1.3991e-08 1.776525563572604 1.3992e-08 1.6957668053750299 1.3993e-08 1.838354804630783 1.3994e-08 1.866788995355377 1.3994999999999999e-08 1.841312819412378 1.3996e-08 1.790229676032525 1.3997e-08 1.8586109675359106 1.3997999999999999e-08 1.771971602109018 1.3999e-08 1.8696776813959588 1.4e-08 1.752772102801245 1.4000999999999999e-08 1.7391761837190365 1.4002e-08 1.8607870756083682 1.4003e-08 1.841262064546302 1.4004e-08 1.8286537171034727 1.4005e-08 1.7650688907821634 1.4006e-08 1.7932002619307816 1.4007e-08 1.797924894710515 1.4008e-08 1.7292431448427077 1.4009e-08 1.8759796745393076 1.401e-08 1.7985567905682889 1.4011e-08 1.8145478445055787 1.4012e-08 1.7870927436871678 1.4013e-08 1.8184777061726594 1.4013999999999999e-08 1.8137356937049987 1.4015e-08 1.8166691492850433 1.4016e-08 1.8054711314459915 1.4016999999999999e-08 1.811455329641942 1.4018e-08 1.8138909149257634 1.4019e-08 1.7370522703173752 1.4019999999999999e-08 1.8094783013067888 1.4021e-08 1.834218232385039 1.4022e-08 1.8197189061371104 1.4023e-08 1.801541594824614 1.4024e-08 1.7683320054635379 1.4025e-08 1.8268389543274766 1.4026e-08 1.7743326137101803 1.4027e-08 1.73164010723317 1.4028e-08 1.8001321105509167 1.4029e-08 1.8660203245925113 1.4029999999999999e-08 1.79415237087711 1.4031e-08 1.8533338431358186 1.4032e-08 1.8326229324204828 1.4032999999999999e-08 1.7693809061872918 1.4034e-08 1.8929206393190705 1.4035e-08 1.8392929091480315 1.4035999999999999e-08 1.8495603803700353 1.4037e-08 1.7969994087837824 1.4038e-08 1.797790461095222 1.4039e-08 1.8643564324934174 1.404e-08 1.7847624345552655 1.4041e-08 1.7649466258705016 1.4042e-08 1.8174746776338313 1.4043e-08 1.868749934905106 1.4044e-08 1.84966222841855 1.4045e-08 1.9937449863376302 1.4046e-08 1.7926592068452105 1.4047e-08 1.748627740741 1.4048e-08 1.8098965325039185 1.4048999999999999e-08 1.7751394592210104 1.405e-08 1.7709090481577126 1.4051e-08 1.8175064741886933 1.4051999999999999e-08 1.76966937519677 1.4053e-08 1.7581630362167713 1.4054e-08 1.7897538637167085 1.4054999999999999e-08 1.745081245806762 1.4056e-08 1.7608175994279387 1.4057e-08 1.795856041161983 1.4058e-08 1.7758892585572195 1.4059e-08 1.7838777221272049 1.406e-08 1.8246317824342473 1.4061e-08 1.764664127686281 1.4062e-08 1.7571579226297054 1.4063e-08 1.7935263849269267 1.4064e-08 1.8012536465671003 1.4065e-08 1.782855598031865 1.4066e-08 1.7605195914199745 1.4067e-08 1.8013391327648165 1.4067999999999999e-08 1.8276884257542736 1.4069e-08 1.847119066925017 1.407e-08 1.7666209607436034 1.4070999999999999e-08 1.830842085824741 1.4072e-08 1.7837368993255385 1.4073e-08 1.8415074807439593 1.4073999999999999e-08 1.7270515138149147 1.4075e-08 1.735045536646959 1.4076e-08 1.790710156981137 1.4077e-08 1.7860665702920897 1.4078e-08 1.882381567846334 1.4079e-08 1.8623538797197572 1.408e-08 1.7748029794853968 1.4081e-08 1.8668191108770837 1.4082e-08 1.8300203221145368 1.4083e-08 1.8258419194188698 1.4083999999999999e-08 1.7541391624626574 1.4085e-08 1.833779568343517 1.4086e-08 1.7702812145804192 1.4086999999999999e-08 1.7941167589031395 1.4088e-08 1.8130482950779343 1.4089e-08 1.788632784088855 1.4089999999999999e-08 1.7294524487339906 1.4091e-08 1.830055437179038 1.4092e-08 1.8476885630876165 1.4093e-08 1.7620326272498719 1.4094e-08 1.8133206136242155 1.4095e-08 1.7855658754859585 1.4096e-08 1.8041178920265681 1.4097e-08 1.893293501491432 1.4098e-08 1.7394803246056136 1.4099e-08 1.7055738414905062 1.41e-08 1.8852523719660044 1.4101e-08 1.68940722927373 1.4102e-08 1.8016253257661468 1.4102999999999999e-08 1.8964112842100587 1.4104e-08 1.764868409913559 1.4105e-08 1.7696691705540042 1.4105999999999999e-08 1.8238199487886193 1.4107e-08 1.8685530684045462 1.4108e-08 1.8016268440748 1.4108999999999999e-08 1.8403110187892417 1.411e-08 1.7756611762641845 1.4111e-08 1.683093863014561 1.4112e-08 1.7875824477613185 1.4113e-08 1.8925475458089622 1.4114e-08 1.8150189231931555 1.4115e-08 1.7917526499313143 1.4116e-08 1.7958493465984222 1.4117e-08 1.810584838895205 1.4118e-08 1.775513824105058 1.4118999999999999e-08 1.8379622463995287 1.412e-08 1.7530993695806247 1.4121e-08 1.7572089983905685 1.4121999999999999e-08 1.7183161881544389 1.4123e-08 1.6790017615087394 1.4124e-08 1.7463732363357576 1.4124999999999999e-08 1.7746216966400132 1.4126e-08 1.8362863450288958 1.4127e-08 1.8515664915384662 1.4128e-08 1.8069738909634454 1.4129e-08 1.7546468222968004 1.413e-08 1.8241424969377227 1.4131e-08 1.7575558201156065 1.4132e-08 1.8647458082750537 1.4133e-08 1.8174050424751802 1.4134e-08 1.8477162224942871 1.4135e-08 1.8295946535267626 1.4136e-08 1.856747768193388 1.4137e-08 1.8173428400991456 1.4137999999999999e-08 1.818850749301091 1.4139e-08 1.803351613588879 1.414e-08 1.7216671271918806 1.4140999999999999e-08 1.759401773019022 1.4142e-08 1.7802325577571456 1.4143e-08 1.7706231352514026 1.4143999999999999e-08 1.7950041971301232 1.4145e-08 1.81036696639704 1.4146e-08 1.7500265683923555 1.4147e-08 1.7496058165307797 1.4148e-08 1.827170353737297 1.4149e-08 1.8034815702283926 1.415e-08 1.844965421260985 1.4151e-08 1.7557746222912274 1.4152e-08 1.8339096820336152 1.4153e-08 1.7645286274468712 1.4153999999999999e-08 1.6914517114043188 1.4155e-08 1.8953318433952926 1.4156e-08 1.7569998837890894 1.4156999999999999e-08 1.826751129493822 1.4158e-08 1.785927259808193 1.4159e-08 1.8331082408092998 1.4159999999999999e-08 1.7972342793421048 1.4161e-08 1.779765928363269 1.4162e-08 1.895998667852713 1.4162999999999999e-08 1.8479182339824956 1.4164e-08 1.834619507575913 1.4165e-08 1.805010116651963 1.4166e-08 1.7935253002467082 1.4167e-08 1.7942825332058019 1.4168e-08 1.713940106868693 1.4169e-08 1.8041357147968502 1.417e-08 1.8276798859905232 1.4171e-08 1.7408905597371118 1.4172e-08 1.7937270548654585 1.4172999999999999e-08 1.7970735515485454 1.4174e-08 1.9071298055074823 1.4175e-08 1.7075146042371552 1.4175999999999999e-08 1.8491566487023925 1.4177e-08 1.793331604959385 1.4178e-08 1.748502690810649 1.4178999999999999e-08 1.8079103528441174 1.418e-08 1.7381510615540725 1.4181e-08 1.7219340976366526 1.4182e-08 1.7182717904922449 1.4183e-08 1.8092297694764436 1.4184e-08 1.8131242657097657 1.4185e-08 1.9264667820461634 1.4186e-08 1.8766491623407582 1.4187e-08 1.83796133348373 1.4188e-08 1.8297111006775904 1.4189e-08 1.8272566663142884 1.419e-08 1.7721101611242298 1.4191e-08 1.7605828315291627 1.4191999999999999e-08 1.7609912183191092 1.4193e-08 1.8694175873973886 1.4194e-08 1.7959892489239282 1.4194999999999999e-08 1.840570728659713 1.4196e-08 1.7993797775579872 1.4197e-08 1.8462473486718816 1.4197999999999999e-08 1.7095130198736201 1.4199e-08 1.738517085586099 1.42e-08 1.7966036944090293 1.4201e-08 1.8387075435891436 1.4202e-08 1.770211527398488 1.4203e-08 1.8649816612973769 1.4204e-08 1.7683462671140324 1.4205e-08 1.79074253812205 1.4206e-08 1.8403069878791274 1.4207e-08 1.8530285516825253 1.4207999999999999e-08 1.7141095995205653 1.4209e-08 1.8888326607231138 1.421e-08 1.8109174364536544 1.4210999999999999e-08 1.7853138816244734 1.4212e-08 1.7422763289341343 1.4213e-08 1.8528670065441668 1.4213999999999999e-08 1.9378531538884052 1.4215e-08 1.6846949478302982 1.4216e-08 1.8202723860186076 1.4217e-08 1.8545408424096326 1.4218e-08 1.8271619821315657 1.4219e-08 1.813996133728298 1.422e-08 1.627531202183201 1.4221e-08 1.8391441064776424 1.4222e-08 1.787308056963287 1.4223e-08 1.836801814570399 1.4224e-08 1.906737832836498 1.4225e-08 1.7202824951225206 1.4226e-08 1.7905091152633705 1.4226999999999999e-08 1.7513169580720938 1.4228e-08 1.7945142108874508 1.4229e-08 1.8043514529010778 1.4229999999999999e-08 1.8369663637809155 1.4231e-08 1.805673219739732 1.4232e-08 1.7736433675337913 1.4232999999999999e-08 1.8240596712244548 1.4234e-08 1.8177940877178018 1.4235e-08 1.792717373661156 1.4236e-08 1.7385382032131613 1.4237e-08 1.7838742383219945 1.4238e-08 1.6809351441047122 1.4239e-08 1.8247558454875616 1.424e-08 1.7679916661574744 1.4241e-08 1.8923202036127478 1.4242e-08 1.9363399762811468 1.4242999999999999e-08 1.8863894124230223 1.4244e-08 1.821847049386265 1.4245e-08 1.7684599368087357 1.4245999999999999e-08 1.8183899734706248 1.4247e-08 1.8093990493107581 1.4248e-08 1.8221287451409498 1.4248999999999999e-08 1.772838626633831 1.425e-08 1.8519680247929509 1.4251e-08 1.8055003389179074 1.4252e-08 1.8187136263336092 1.4253e-08 1.7938139663559847 1.4254e-08 1.7878585930327855 1.4255e-08 1.856995795723927 1.4256e-08 1.8291563533383712 1.4257e-08 1.841882935420292 1.4258e-08 1.7921221989394511 1.4259e-08 1.7701650009777412 1.426e-08 1.8040674496830256 1.4261e-08 1.7724967313107294 1.4261999999999999e-08 1.7890040067318418 1.4263e-08 1.7953439922483416 1.4264e-08 1.8160895140869984 1.4264999999999999e-08 1.8230789325476722 1.4266e-08 1.8140105772911979 1.4267e-08 1.865588766606161 1.4267999999999999e-08 1.8196597492340445 1.4269e-08 1.8880315970848132 1.427e-08 1.869832547273712 1.4271e-08 1.7909027821524868 1.4272e-08 1.7545463090713584 1.4273e-08 1.7321096542015464 1.4274e-08 1.8249421745733727 1.4275e-08 1.8477222197034435 1.4276e-08 1.954194877367797 1.4277e-08 1.791495737297511 1.4278e-08 1.8209572469420514 1.4279e-08 1.8864750541134616 1.428e-08 1.9114487932907025 1.4280999999999999e-08 1.8646796761696043 1.4282e-08 1.8053480897417409 1.4283e-08 1.8990762129526424 1.4283999999999999e-08 1.7599830920141928 1.4285e-08 1.7431994673558158 1.4286e-08 1.9520417089215827 1.4286999999999999e-08 1.789561651049158 1.4288e-08 1.767306635160156 1.4289e-08 1.7659879623133976 1.429e-08 1.8768574927166555 1.4291e-08 1.7297152904571516 1.4292e-08 1.8248204758326358 1.4293e-08 1.8251202875143162 1.4294e-08 1.7807374214528584 1.4295e-08 1.7222384556961754 1.4296e-08 1.7841556199530102 1.4296999999999999e-08 1.8106035160461618 1.4298e-08 1.8347177400220471 1.4299e-08 1.7614243528461853 1.4299999999999999e-08 1.7973673816405389 1.4301e-08 1.8054276268168608 1.4302e-08 1.6743472243424407 1.4302999999999999e-08 1.7883509678932785 1.4304e-08 1.801046036421814 1.4305e-08 1.7908017227705675 1.4306e-08 1.8300521419181184 1.4307e-08 1.9022585467744832 1.4308e-08 1.7596542437785976 1.4309e-08 1.7842225909831793 1.431e-08 1.954743037916949 1.4311e-08 1.800523886520496 1.4312e-08 1.7861029698102262 1.4313e-08 1.8167797639731098 1.4314e-08 1.8584635068424384 1.4315e-08 1.6996364862100386 1.4315999999999999e-08 1.8623941112779931 1.4317e-08 1.8283316815715747 1.4318e-08 1.7405053194251972 1.4318999999999999e-08 1.906594755532674 1.432e-08 1.7265701258145354 1.4321e-08 1.7876665168255181 1.4321999999999999e-08 1.7915456107637546 1.4323e-08 1.8755651377600076 1.4324e-08 1.7247668671697791 1.4325e-08 1.8299560285083054 1.4326e-08 1.7635726867740327 1.4327e-08 1.7965237273288404 1.4328e-08 1.8196681759082793 1.4329e-08 1.8734144246501305 1.433e-08 1.816005340243134 1.4331e-08 1.8463798135464613 1.4331999999999999e-08 1.8070355396197084 1.4333e-08 1.9157796539444436 1.4334e-08 1.7949407674915854 1.4334999999999999e-08 1.755550837957202 1.4336e-08 1.8034255924793956 1.4337e-08 1.7852962721907382 1.4337999999999999e-08 1.7052855839800372 1.4339e-08 1.820851949075948 1.434e-08 1.7699978283203703 1.4341e-08 1.803672084583895 1.4342e-08 1.7502240059958465 1.4343e-08 1.8041490052549602 1.4344e-08 1.7641709793976403 1.4345e-08 1.7490824602700923 1.4346e-08 1.8023293302846979 1.4347e-08 1.8261146312180048 1.4348e-08 1.9036736572337 1.4349e-08 1.8633652754633134 1.435e-08 1.7859658945134205 1.4350999999999999e-08 1.657453313031656 1.4352e-08 1.8080904490938914 1.4353e-08 1.7684285979223668 1.4353999999999999e-08 1.840590176255823 1.4355e-08 1.967988866560261 1.4356e-08 1.82748785616437 1.4356999999999999e-08 1.8748432722487984 1.4358e-08 1.7727371553141926 1.4359e-08 1.856866994231441 1.436e-08 1.7666214825481512 1.4361e-08 1.7509132505967315 1.4362e-08 1.7830767292251297 1.4363e-08 1.8048584007102602 1.4364e-08 1.8836839581186076 1.4365e-08 1.803392816783188 1.4366e-08 1.7803506175801138 1.4367e-08 1.757595931968954 1.4368e-08 1.7049229952869913 1.4369e-08 1.8347288428954782 1.4369999999999999e-08 1.7988919012347944 1.4371e-08 1.778076269645361 1.4372e-08 1.8080095537237997 1.4372999999999999e-08 1.7801530787064457 1.4374e-08 1.8298066302517286 1.4375e-08 1.8508040987792385 1.4375999999999999e-08 1.8634797597506154 1.4377e-08 1.878037834868428 1.4378e-08 1.7773002996538059 1.4379e-08 1.8038314931890778 1.438e-08 1.787414799043039 1.4381e-08 1.7948825674249516 1.4382e-08 1.7859267654099817 1.4383e-08 1.8348342281765289 1.4384e-08 1.764309756666341 1.4385e-08 1.821683664084309 1.4385999999999999e-08 1.740592819728029 1.4387e-08 1.794950778131036 1.4388e-08 1.9179373594910851 1.4388999999999999e-08 1.8035196502431243 1.439e-08 1.692634821506273 1.4391e-08 1.8088263471712307 1.4391999999999999e-08 1.750758853201506 1.4393e-08 1.796186674971116 1.4394e-08 1.7686487283506476 1.4395e-08 1.8484818725367917 1.4396e-08 1.7619891325857473 1.4397e-08 1.8212461896961734 1.4398e-08 1.7405124660569629 1.4399e-08 1.8770986990013088 1.44e-08 1.7645002770200386 1.4401e-08 1.8122730316174769 1.4402e-08 1.7799739069728684 1.4403e-08 1.8403625570531186 1.4404e-08 1.82333095466777 1.4404999999999999e-08 1.8365519291949985 1.4406e-08 1.8698944318821211 1.4407e-08 1.8229126951837447 1.4407999999999999e-08 1.8834220568413007 1.4409e-08 1.8393013393118387 1.441e-08 1.8720791180703669 1.4410999999999999e-08 1.8644477879782477 1.4412e-08 1.7578289396708178 1.4413e-08 1.808726720974242 1.4414e-08 1.7910989299599818 1.4415e-08 1.8749031794158553 1.4416e-08 1.777017710142898 1.4417e-08 1.775362296795064 1.4418e-08 1.796442234978151 1.4419e-08 1.8027696628716978 1.442e-08 1.896109056766776 1.4420999999999999e-08 1.717631139575101 1.4422e-08 1.8369153751472962 1.4423e-08 1.7559483380168395 1.4423999999999999e-08 1.8018287692734158 1.4425e-08 1.7744020008863066 1.4426e-08 1.8287051243139727 1.4426999999999999e-08 1.7815482146934696 1.4428e-08 1.8002897218814387 1.4429e-08 1.8056638065864667 1.443e-08 1.8410714128878032 1.4431e-08 1.8814780366273338 1.4432e-08 1.7647963954651398 1.4433e-08 1.9171138936450454 1.4434e-08 1.739794891783918 1.4435e-08 1.7630558282139377 1.4436e-08 1.7733939747140297 1.4437e-08 1.7385609988916533 1.4438e-08 1.7032181290377848 1.4439e-08 1.8428968215760952 1.4439999999999999e-08 1.7810261102175522 1.4441e-08 1.8765045152219317 1.4442e-08 1.7727187928268044 1.4442999999999999e-08 1.8707672844384864 1.4444e-08 1.8316745983205431 1.4445e-08 1.7976441526618867 1.4445999999999999e-08 1.7679718317009412 1.4447e-08 1.7591668916060996 1.4448e-08 1.8174737193071706 1.4449e-08 1.8464511293044816 1.445e-08 1.880336938807253 1.4451e-08 1.6871046877877562 1.4452e-08 1.852396016464686 1.4453e-08 1.7764007997329156 1.4454e-08 1.752383194590078 1.4455e-08 1.8029982324858445 1.4455999999999999e-08 1.8198806985146372 1.4457e-08 1.873476636672702 1.4458e-08 1.803982076788068 1.4458999999999999e-08 1.7351830442960539 1.446e-08 1.8285649612040766 1.4461e-08 1.7193717723717017 1.4461999999999999e-08 1.8631117296093727 1.4463e-08 1.7320690441693856 1.4464e-08 1.7845624469236465 1.4464999999999999e-08 1.7598066765241274 1.4466e-08 1.8117474699605245 1.4467e-08 1.7927111268192846 1.4468e-08 1.8278797364122996 1.4469e-08 1.8211162259557663 1.447e-08 1.8091672616728336 1.4471e-08 1.7397059301646676 1.4472e-08 1.7810449786030507 1.4473e-08 1.8043762523675946 1.4474e-08 1.7987553658264501 1.4474999999999999e-08 1.8245136392735655 1.4476e-08 1.843766427577668 1.4477e-08 1.865318983438668 1.4477999999999999e-08 1.6806265008393548 1.4479e-08 1.8414916024180656 1.448e-08 1.7892720785216694 1.4480999999999999e-08 1.8099364166514975 1.4482e-08 1.9332839256112784 1.4483e-08 1.712785731457798 1.4484e-08 1.7443554727916208 1.4485e-08 1.7971328512720481 1.4486e-08 1.7516127597136903 1.4487e-08 1.7869649437423911 1.4488e-08 1.7932530011828953 1.4489e-08 1.757325544208894 1.449e-08 1.7244359615459426 1.4491e-08 1.865750547350362 1.4492e-08 1.8516522191201954 1.4493e-08 1.8043183908588214 1.4493999999999999e-08 1.9194002004584296 1.4495e-08 1.9159336664935045 1.4496e-08 1.7830745851664183 1.4496999999999999e-08 1.7881561995722677 1.4498e-08 1.7181918631095185 1.4499e-08 1.734658393736931 1.4499999999999999e-08 1.7312243094868323 1.4501e-08 1.7941860145719968 1.4502e-08 1.8553044084019077 1.4503e-08 1.7731457342139754 1.4504e-08 1.819604503789388 1.4505e-08 1.8540108863987064 1.4506e-08 1.8113589007691826 1.4507e-08 1.7223438396540005 1.4508e-08 1.8019526396538657 1.4509e-08 1.896961989776638 1.4509999999999999e-08 1.8494390353212984 1.4511e-08 1.7125036016810231 1.4512e-08 1.7119252478652414 1.4512999999999999e-08 1.856783648627609 1.4514e-08 1.754318032520027 1.4515e-08 1.7635197465803039 1.4515999999999999e-08 1.791096460767097 1.4517e-08 1.739646276774037 1.4518e-08 1.8406353650874638 1.4519e-08 1.7101906663435633 1.452e-08 1.8212913554048695 1.4521e-08 1.9005674743842413 1.4522e-08 1.8250574992883608 1.4523e-08 1.8196500018610742 1.4524e-08 1.7222129239349275 1.4525e-08 1.816350986522854 1.4526e-08 1.8024244768453508 1.4527e-08 1.8714884735469193 1.4528e-08 1.8060751820028524 1.4528999999999999e-08 1.77874152883948 1.453e-08 1.8506696711982638 1.4531e-08 1.765355370815114 1.4531999999999999e-08 1.7950235495550053 1.4533e-08 1.9315120516616444 1.4534e-08 1.8363792916456707 1.4534999999999999e-08 1.858264056070329 1.4536e-08 1.7982593200173744 1.4537e-08 1.8515911446902396 1.4538e-08 1.8006487255166437 1.4539e-08 1.8250939277132943 1.454e-08 1.7177065147714445 1.4541e-08 1.8375268131499858 1.4542e-08 1.8612121894218694 1.4543e-08 1.8165715203487214 1.4544e-08 1.8005583979821653 1.4544999999999999e-08 1.743063869187988 1.4546e-08 1.6854650127529809 1.4547e-08 1.746938797835445 1.4547999999999999e-08 1.7680039656620352 1.4549e-08 1.8261619802106555 1.455e-08 1.848758793855718 1.4550999999999999e-08 1.702238805486318 1.4552e-08 1.79859979607141 1.4553e-08 1.7485734457032764 1.4553999999999999e-08 1.7383188742123228 1.4555e-08 1.7431100811763744 1.4556e-08 1.8404938754827407 1.4557e-08 1.756856555691938 1.4558e-08 1.880578901530403 1.4559e-08 1.8511134897612658 1.456e-08 1.87951380558746 1.4561e-08 1.797209496611964 1.4562e-08 1.8003535471694463 1.4563e-08 1.751756332992112 1.4563999999999999e-08 1.7478363736279836 1.4565e-08 1.8273434604744836 1.4566e-08 1.7983195615945577 1.4566999999999999e-08 1.8051345503649268 1.4568e-08 1.7450276466030397 1.4569e-08 1.7743793383327564 1.4569999999999999e-08 1.7949480334259316 1.4571e-08 1.8181647029052865 1.4572e-08 1.877270844840617 1.4573e-08 1.8298779935402245 1.4574e-08 1.769151926939057 1.4575e-08 1.8027468821186736 1.4576e-08 1.920606896472146 1.4577e-08 1.7393929030485606 1.4578e-08 1.8537820078334395 1.4579e-08 1.8239364795763582 1.458e-08 1.8385164207317346 1.4581e-08 1.7640773001249936 1.4582e-08 1.7100128848446665 1.4582999999999999e-08 1.7366689035289615 1.4584e-08 1.841083999847052 1.4585e-08 1.853222406942353 1.4585999999999999e-08 1.7776590993703114 1.4587e-08 1.7549101687302555 1.4588e-08 1.7685616792009575 1.4588999999999999e-08 1.7459775109267084 1.459e-08 1.839365527531112 1.4591e-08 1.8897416602559942 1.4592e-08 1.8457449172497264 1.4593e-08 1.7622896722487036 1.4594e-08 1.8580776385683535 1.4595e-08 1.8716168471723857 1.4596e-08 1.7323234993893504 1.4597e-08 1.8529936880525983 1.4598e-08 1.8629696909745441 1.4598999999999999e-08 1.785560121854946 1.46e-08 1.7790511312331725 1.4601e-08 1.802928188031175 1.4601999999999999e-08 1.8217618018548205 1.4603e-08 1.7632978152774257 1.4604e-08 1.7603215834341623 1.4604999999999999e-08 1.7922942040128713 1.4606e-08 1.7635575501397687 1.4607e-08 1.7719975704297433 1.4608e-08 1.8074510766466636 1.4609e-08 1.802646944795142 1.461e-08 1.8641896062797498 1.4611e-08 1.7967305122196495 1.4612e-08 1.8413510215368887 1.4613e-08 1.8314015227042286 1.4614e-08 1.784156462961966 1.4615e-08 1.7408906747942452 1.4616e-08 1.7464323067654008 1.4617e-08 1.7760444235258963 1.4617999999999999e-08 1.746029480040215 1.4619e-08 1.823170947395192 1.462e-08 1.779699158159389 1.4620999999999999e-08 1.8009253312223499 1.4622e-08 1.810759629863912 1.4623e-08 1.787837326691951 1.4623999999999999e-08 1.7849305076081265 1.4625e-08 1.8140090265099764 1.4626e-08 1.799449905174895 1.4627e-08 1.7717253201678123 1.4628e-08 1.8311282318827649 1.4629e-08 1.8537597352743054 1.463e-08 1.741240293072421 1.4631e-08 1.814939117446307 1.4632e-08 1.7835676868813224 1.4633e-08 1.7747181070282512 1.4633999999999999e-08 1.8265880212045877 1.4635e-08 1.7588638833610786 1.4636e-08 1.8125878084324212 1.4636999999999999e-08 1.707268083657371 1.4638e-08 1.821588642877449 1.4639e-08 1.875040411347173 1.4639999999999999e-08 1.8305646308250647 1.4641e-08 1.784489298159973 1.4642e-08 1.834337183912201 1.4642999999999999e-08 1.8179742901979212 1.4644e-08 1.893269234572349 1.4645e-08 1.8116689041444949 1.4646e-08 1.8020753069935622 1.4647e-08 1.8063392056252952 1.4648e-08 1.84339396939576 1.4649e-08 1.7683470020912158 1.465e-08 1.8645917774319047 1.4651e-08 1.8214758617225701 1.4652e-08 1.7893961862618566 1.4652999999999999e-08 1.7605558201571763 1.4654e-08 1.7357461730545005 1.4655e-08 1.803291090757034 1.4655999999999999e-08 1.866221514366288 1.4657e-08 1.8284947512120724 1.4658e-08 1.7257575223267332 1.4658999999999999e-08 1.8409301662422313 1.466e-08 1.8513004000859032 1.4661e-08 1.7886356471752614 1.4662e-08 1.7666644201928894 1.4663e-08 1.7800375222999962 1.4664e-08 1.747230152658084 1.4665e-08 1.7407500756837502 1.4666e-08 1.7270607503271875 1.4667e-08 1.795029016538955 1.4668e-08 1.779756092688128 1.4669e-08 1.7753319130594987 1.467e-08 1.8067853037656771 1.4671e-08 1.8274047443227326 1.4671999999999999e-08 1.8104888096344505 1.4673e-08 1.7243519697682155 1.4674e-08 1.8925925203365621 1.4674999999999999e-08 1.8403008166273362 1.4676e-08 1.801387125680618 1.4677e-08 1.8535803590399873 1.4677999999999999e-08 1.7038816461122597 1.4679e-08 1.842507639804851 1.468e-08 1.833690703514674 1.4681e-08 1.7991919571335109 1.4682e-08 1.8748363126407248 1.4683e-08 1.7462631565493538 1.4684e-08 1.7831864249345437 1.4685e-08 1.7427674288909984 1.4686e-08 1.804270122158046 1.4687e-08 1.8832890128732445 1.4687999999999999e-08 1.6945654932260865 1.4689e-08 1.8150261540945376 1.469e-08 1.807586986297604 1.4690999999999999e-08 1.820066702030613 1.4692e-08 1.8213544777821393 1.4693e-08 1.8196903010264558 1.4693999999999999e-08 1.7491149526726917 1.4695e-08 1.746066942973129 1.4696e-08 1.814640990152321 1.4697e-08 1.8487300315946915 1.4698e-08 1.7702470952542748 1.4699e-08 1.787557951330021 1.47e-08 1.8475120066518376 1.4701e-08 1.840367236059019 1.4702e-08 1.7999191396864715 1.4703e-08 1.8638052527884907 1.4704e-08 1.7275155823446247 1.4705e-08 1.938177018014143 1.4706e-08 1.8370368055163024 1.4706999999999999e-08 1.8394730873541631 1.4708e-08 1.7714566748827596 1.4709e-08 1.8018254745691027 1.4709999999999999e-08 1.73794283782464 1.4711e-08 1.827980399623734 1.4712e-08 1.8259589605046629 1.4712999999999999e-08 1.769192549788837 1.4714e-08 1.7262883489241212 1.4715e-08 1.7904150581472966 1.4716e-08 1.7684413088661726 1.4717e-08 1.7397296178401558 1.4718e-08 1.7628083001075987 1.4719e-08 1.8040042315489597 1.472e-08 1.7027513879182306 1.4721e-08 1.7688691893065736 1.4722e-08 1.8411523981456979 1.4722999999999999e-08 1.9002747543286722 1.4724e-08 1.7750781128542403 1.4725e-08 1.7518241205408123 1.4725999999999999e-08 1.762726824342521 1.4727e-08 1.8506059619156838 1.4728e-08 1.8126128650381157 1.4728999999999999e-08 1.8213311458542851 1.473e-08 1.8072914212979616 1.4731e-08 1.8410648926344668 1.4731999999999999e-08 1.739378217545829 1.4733e-08 1.7543984217417108 1.4734e-08 1.844325141416407 1.4735e-08 1.8417293179472836 1.4736e-08 1.7096692445729822 1.4737e-08 1.904402476035923 1.4738e-08 1.7775108303184168 1.4739e-08 1.6766611533138613 1.474e-08 1.7489493204901598 1.4741e-08 1.8054672916410157 1.4741999999999999e-08 1.7636160569002706 1.4743e-08 1.7353997748496093 1.4744e-08 1.7740828379192295 1.4744999999999999e-08 1.8488647284982225 1.4746e-08 1.7985902368668338 1.4747e-08 1.8646016351320795 1.4747999999999999e-08 1.7687569293241456 1.4749e-08 1.8665615661214505 1.475e-08 1.8338050245692812 1.4751e-08 1.777166610982571 1.4752e-08 1.7688433634879301 1.4753e-08 1.8400531473631847 1.4754e-08 1.851969741278124 1.4755e-08 1.8170106377393875 1.4756e-08 1.7782989968214231 1.4757e-08 1.8202881351438216 1.4758e-08 1.7812130874262666 1.4759e-08 1.7607947861934066 1.476e-08 1.8432273997497675 1.4760999999999999e-08 1.7856716714158414 1.4762e-08 1.8445914636893939 1.4763e-08 1.721905223449465 1.4763999999999999e-08 1.7984383318654247 1.4765e-08 1.8264889164906384 1.4766e-08 1.7611920817602642 1.4766999999999999e-08 1.7894719375079742 1.4768e-08 1.807566806392214 1.4769e-08 1.7535234480950916 1.477e-08 1.7855355832749942 1.4771e-08 1.6774652281218767 1.4772e-08 1.842753750508823 1.4773e-08 1.8972346749242321 1.4774e-08 1.8582448972830254 1.4775e-08 1.8275297940751185 1.4776e-08 1.7212010548691874 1.4776999999999999e-08 1.8675100603559824 1.4778e-08 1.7420805159820225 1.4779e-08 1.7808898856625053 1.4779999999999999e-08 1.8024618559271801 1.4781e-08 1.7890443293874678 1.4782e-08 1.7582540513117961 1.4782999999999999e-08 1.7626284423510412 1.4784e-08 1.8179590248833997 1.4785e-08 1.8458417328322072 1.4786e-08 1.8377364472015065 1.4787e-08 1.8534069325506484 1.4788e-08 1.7429547149569438 1.4789e-08 1.8604054016327278 1.479e-08 1.7837413414279752 1.4791e-08 1.9130593579928399 1.4792e-08 1.7204592506721412 1.4793e-08 1.7753541456388071 1.4794e-08 1.7570620596845188 1.4795e-08 1.8759059521420167 1.4795999999999999e-08 1.8106954209479247 1.4797e-08 1.729711806861874 1.4798e-08 1.7305386052540397 1.4798999999999999e-08 1.7346042329169025 1.48e-08 1.8134801959275655 1.4801e-08 1.8559234215746796 1.4801999999999999e-08 1.7889299753025638 1.4803e-08 1.6859186713522039 1.4804e-08 1.9147661013016113 1.4805e-08 1.753713716460704 1.4806e-08 1.7525524495792644 1.4807e-08 1.7834504952366579 1.4808e-08 1.8067460161879372 1.4809e-08 1.777518805990434 1.481e-08 1.8738864236918202 1.4811e-08 1.836036646414951 1.4811999999999999e-08 1.84231682682474 1.4813e-08 1.826030746419148 1.4814e-08 1.814235011706567 1.4814999999999999e-08 1.8546060508024924 1.4816e-08 1.8188855027353839 1.4817e-08 1.7258861695348329 1.4817999999999999e-08 1.758144647173783 1.4819e-08 1.8505401554428555 1.482e-08 1.7825791209998134 1.4821e-08 1.796826378862526 1.4822e-08 1.747887214149314 1.4823e-08 1.8558857634246968 1.4824e-08 1.8811104065636566 1.4825e-08 1.7430511733181993 1.4826e-08 1.798678824606236 1.4827e-08 1.8346194465550814 1.4828e-08 1.8174794313065168 1.4829e-08 1.8084778881007353 1.483e-08 1.7648962131456702 1.4830999999999999e-08 1.7540220379492082 1.4832e-08 1.8389760143344218 1.4833e-08 1.8553841755610232 1.4833999999999999e-08 1.7729749946302582 1.4835e-08 1.78201176256939 1.4836e-08 1.6928140428870184 1.4836999999999999e-08 1.7194101625817477 1.4838e-08 1.820218523101112 1.4839e-08 1.8363439106587893 1.484e-08 1.8249381322085065 1.4841e-08 1.8551703923714573 1.4842e-08 1.8186035696155547 1.4843e-08 1.730799408189153 1.4844e-08 1.7407135634526838 1.4845e-08 1.7987483322237112 1.4846e-08 1.8353025721157472 1.4846999999999999e-08 1.715435475418204 1.4848e-08 1.737399072656013 1.4849e-08 1.7702097614377612 1.4849999999999999e-08 1.7332503197704043 1.4851e-08 1.8161771184830677 1.4852e-08 1.8139465778175208 1.4852999999999999e-08 1.8614841591624327 1.4854e-08 1.7909426512145559 1.4855e-08 1.7665300333121177 1.4855999999999999e-08 1.6827308470886462 1.4857e-08 1.8278098899442075 1.4858e-08 1.7359791849442079 1.4859e-08 1.8052711860098798 1.486e-08 1.8129866551742517 1.4861e-08 1.6354350327423592 1.4862e-08 1.7715793856948243 1.4863e-08 1.7916028992610482 1.4864e-08 1.7802153634577003 1.4865e-08 1.7696660376681201 1.4865999999999999e-08 1.8007011333978309 1.4867e-08 1.8354496857840057 1.4868e-08 1.8278913644694672 1.4868999999999999e-08 1.8394793328889967 1.487e-08 1.7583236688581074 1.4871e-08 1.8258741672227 1.4871999999999999e-08 1.8687942469632923 1.4873e-08 1.7841008550054342 1.4874e-08 1.7540751081705515 1.4875e-08 1.8021859347835523 1.4876e-08 1.8479721105495976 1.4877e-08 1.7623875399773592 1.4878e-08 1.8467041473260037 1.4879e-08 1.7003257927219968 1.488e-08 1.7589596104376237 1.4881e-08 1.8190354034074023 1.4882e-08 1.7877822103191254 1.4883e-08 1.792201678392747 1.4884e-08 1.9155891541270904 1.4884999999999999e-08 1.730059391172101 1.4886e-08 1.9289760033593648 1.4887e-08 1.866983694349887 1.4887999999999999e-08 1.786072355719619 1.4889e-08 1.816248362330937 1.489e-08 1.8760287133339575 1.4890999999999999e-08 1.851513971338704 1.4892e-08 1.9046783418186406 1.4893e-08 1.8191105088848727 1.4894e-08 1.7348621581932135 1.4895e-08 1.7672992709802338 1.4896e-08 1.8031053314954324 1.4897e-08 1.7830893216833268 1.4898e-08 1.8058726660004463 1.4899e-08 1.7464778575436513 1.49e-08 1.8702229965891246 1.4900999999999999e-08 1.8401987058544795 1.4902e-08 1.8280849837587363 1.4903e-08 1.8180094381639917 1.4904e-08 1.8405129487432526 1.4905e-08 1.737126027314122 1.4906e-08 1.724985052777219 1.4907e-08 1.8183915901841585 1.4908e-08 1.705437965207266 1.4909e-08 1.782084173809115 1.491e-08 1.8064959574253852 1.4911e-08 1.77143516700592 1.4911999999999998e-08 1.7994303755051542 1.4913e-08 1.7719515278694693 1.4914e-08 1.8206794176576957 1.4914999999999998e-08 1.8202064068424624 1.4916e-08 1.7854805909234663 1.4917e-08 1.7804122728937897 1.4917999999999998e-08 1.8519557153639343 1.4919e-08 1.830045724156387 1.492e-08 1.8146855223580363 1.4921e-08 1.8332060290750392 1.4922e-08 1.7948634525610423 1.4923e-08 1.7744472663755066 1.4924e-08 1.8525265694028443 1.4925e-08 1.8040355323286967 1.4926e-08 1.7860166759358642 1.4927e-08 1.8215182675435402 1.4928e-08 1.7408641687459456 1.4929e-08 1.7970178745097296 1.493e-08 1.7729234300354884 1.4931e-08 1.7875448269968037 1.4932e-08 1.8393373717425212 1.4933e-08 1.7407100433258138 1.4934e-08 1.8315360975795762 1.4935e-08 1.8032762080301286 1.4936e-08 1.8082778972519589 1.4937e-08 1.7528042764619427 1.4938e-08 1.7177652273937578 1.4939e-08 1.7681760090245853 1.494e-08 1.7909069581893295 1.4941e-08 1.8906199068122442 1.4942e-08 1.823894232273963 1.4943e-08 1.8628964658690788 1.4944e-08 1.7644307595027318 1.4945e-08 1.7823447170859812 1.4946e-08 1.8219913978509688 1.4946999999999998e-08 1.7926957884227177 1.4948e-08 1.7917087852151463 1.4949e-08 1.8384871084656595 1.4949999999999998e-08 1.803865779848556 1.4951e-08 1.8998445390080736 1.4952e-08 1.8165270792796966 1.4952999999999998e-08 1.8052073897564065 1.4954e-08 1.8086973597611289 1.4955e-08 1.8183096133670409 1.4956e-08 1.793609218672726 1.4957e-08 1.8076105947498138 1.4958e-08 1.8892976817211997 1.4959e-08 1.8676385544561558 1.496e-08 1.8438888462745275 1.4961e-08 1.768149545143836 1.4962e-08 1.8050280990987606 1.4963e-08 1.7408372279768594 1.4964e-08 1.756285477626915 1.4965e-08 1.7796050526298346 1.4966e-08 1.8341312620838517 1.4967e-08 1.7686776366384458 1.4968e-08 1.7270220597529917 1.4969e-08 1.8065716436401835 1.497e-08 1.8469559202351105 1.4971e-08 1.785114165460443 1.4972e-08 1.7465818577367793 1.4973e-08 1.737643532051827 1.4974e-08 1.7255353702951508 1.4975e-08 1.7422058716213544 1.4976e-08 1.7674356805641842 1.4977e-08 1.809806176999514 1.4978e-08 1.799654900479071 1.4979e-08 1.8202653047883859 1.498e-08 1.730987955323832 1.4981e-08 1.7893373330299123 1.4981999999999998e-08 1.7975704861226016 1.4983e-08 1.7953400430572346 1.4984e-08 1.8072695318937584 1.4984999999999998e-08 1.7490439803374065 1.4986e-08 1.73534769661282 1.4987e-08 1.7521553100511147 1.4987999999999998e-08 1.8022900834674065 1.4989e-08 1.8844901690254274 1.499e-08 1.7321529726123155 1.4991e-08 1.756111222376413 1.4992e-08 1.8207800922294564 1.4993e-08 1.7947014712783749 1.4994e-08 1.7267871352265274 1.4995e-08 1.756060485715799 1.4996e-08 1.7726124389143092 1.4997e-08 1.8142685884871945 1.4998e-08 1.7468753565837214 1.4999e-08 1.7881840237772448 1.5e-08 1.77935761227046 1.5001e-08 1.7348054980838754 1.5002e-08 1.7769647573891354 1.5003e-08 1.693362144840986 1.5004e-08 1.8050832558865233 1.5005e-08 1.9057603879370122 1.5006e-08 1.776971303467963 1.5007e-08 1.813121668924526 1.5008e-08 1.8553722340385816 1.5009e-08 1.8329991969309563 1.501e-08 1.75999660820812 1.5011e-08 1.827512056732897 1.5012e-08 1.7848503121500447 1.5013e-08 1.7248773365355619 1.5014e-08 1.7798047198089268 1.5015e-08 1.8328902278019217 1.5016e-08 1.803297561857676 1.5016999999999998e-08 1.7711982730601399 1.5018e-08 1.7765136886012842 1.5019e-08 1.764526158675366 1.5019999999999998e-08 1.8982962177801337 1.5021e-08 1.7870407373094601 1.5022e-08 1.7459620261982938 1.5022999999999998e-08 1.7290292053423189 1.5024e-08 1.914623209931156 1.5025e-08 1.7874268297089484 1.5026e-08 1.7654554292794389 1.5027e-08 1.7459830101989997 1.5028e-08 1.842271667048605 1.5029e-08 1.7753749466349082 1.503e-08 1.7273261378667462 1.5031e-08 1.8426985293747182 1.5032e-08 1.7720493205483328 1.5033e-08 1.8426109165779923 1.5034e-08 1.9088218237472134 1.5035e-08 1.8330582583467656 1.5036e-08 1.8061905446462398 1.5037e-08 1.7590486784023927 1.5038e-08 1.8558482726451793 1.5039e-08 1.6983846955534474 1.504e-08 1.7871729073687996 1.5041e-08 1.7777801999275806 1.5042e-08 1.8196490541205108 1.5043e-08 1.7731942029363172 1.5044e-08 1.8731958886769062 1.5045e-08 1.802379773409754 1.5046e-08 1.9046810396561131 1.5047e-08 1.7855810963292875 1.5048e-08 1.739284656374177 1.5049e-08 1.8414626831623446 1.505e-08 1.704081088839316 1.5051e-08 1.7657373127533433 1.5051999999999998e-08 1.7285086370931482 1.5053e-08 1.8088054653567887 1.5054e-08 1.7992444810243686 1.5054999999999998e-08 1.8073458056040654 1.5056e-08 1.8771801630131193 1.5057e-08 1.8128474297103174 1.5057999999999998e-08 1.767210053195842 1.5059e-08 1.866611845529788 1.506e-08 1.7893653674816439 1.5060999999999998e-08 1.8146587312507336 1.5062e-08 1.7842161487732742 1.5063e-08 1.8177227905154527 1.5064e-08 1.8853882435940665 1.5065e-08 1.847350107060849 1.5066e-08 1.85587892679076 1.5067e-08 1.822201306554924 1.5068e-08 1.6854005304997146 1.5069e-08 1.8151863063747478 1.507e-08 1.8006267307808024 1.5071e-08 1.8030206240751965 1.5072e-08 1.8170127623270398 1.5073e-08 1.9126376966660776 1.5074e-08 1.8010838358404762 1.5075e-08 1.7788881943907955 1.5076e-08 1.8083962530756363 1.5077e-08 1.8051130329777851 1.5078e-08 1.6675483456859193 1.5079e-08 1.7948735259749764 1.508e-08 1.8165864711885975 1.5081e-08 1.8018245244774014 1.5082e-08 1.7490790648646146 1.5083e-08 1.8157964662933779 1.5084e-08 1.7862215210727415 1.5085e-08 1.823070946241825 1.5086e-08 1.8013513768118494 1.5086999999999998e-08 1.7190647889002983 1.5088e-08 1.9060953851458344 1.5089e-08 1.8536122939827107 1.5089999999999998e-08 1.8555786951937225 1.5091e-08 1.8377289916765118 1.5092e-08 1.852370280558676 1.5092999999999998e-08 1.7843869287417355 1.5094e-08 1.801262165375925 1.5095e-08 1.84661619861613 1.5095999999999998e-08 1.7645132209108183 1.5097e-08 1.839382949943315 1.5098e-08 1.7630021772197786 1.5099e-08 1.8181098112581857 1.51e-08 1.7508373914041728 1.5101e-08 1.7723102118530583 1.5102e-08 1.9016435729710652 1.5103e-08 1.776256132519547 1.5104e-08 1.8297470262945392 1.5105e-08 1.7960626382390874 1.5106e-08 1.8446668959646 1.5107e-08 1.778500912517471 1.5108e-08 1.7961977028046687 1.5109e-08 1.7333819110759678 1.511e-08 1.8021188462871258 1.5111e-08 1.7286245532875113 1.5112e-08 1.8331477364935491 1.5113e-08 1.7828235029783954 1.5114e-08 1.8412745547880185 1.5115e-08 1.7890532654905893 1.5116e-08 1.7771483713702982 1.5117e-08 1.801605893258045 1.5118e-08 1.8205446572414157 1.5119e-08 1.7753848188048482 1.512e-08 1.7925093879115497 1.5121e-08 1.8545603669023674 1.5122e-08 1.7482385917326992 1.5123e-08 1.7762437827176807 1.5124e-08 1.7877566980836888 1.5124999999999998e-08 1.734040176958423 1.5126e-08 1.7418448822160446 1.5127e-08 1.773069775098729 1.5127999999999998e-08 1.7521141199084669 1.5129e-08 1.8824203057127944 1.513e-08 1.8207148025315631 1.5130999999999998e-08 1.7882629921434232 1.5132e-08 1.7586720023908808 1.5133e-08 1.869822086846028 1.5134e-08 1.8224586765143946 1.5135e-08 1.8811354772558515 1.5136e-08 1.8041447279717575 1.5137e-08 1.818017991656478 1.5138e-08 1.6576058463364078 1.5139e-08 1.8413500156951834 1.514e-08 1.7429266598195448 1.5141e-08 1.6927811337144412 1.5142e-08 1.80732126128939 1.5143e-08 1.7835393581841386 1.5144e-08 1.7728350751294277 1.5145e-08 1.8057841898816636 1.5146e-08 1.7922965104412214 1.5147e-08 1.8268611982089769 1.5148e-08 1.7340056584959687 1.5149e-08 1.8004068774869662 1.515e-08 1.8064154421787628 1.5151e-08 1.7512039348763022 1.5152e-08 1.754449537833256 1.5153e-08 1.8621910126538117 1.5154e-08 1.6957896018205767 1.5155e-08 1.767221326061476 1.5156e-08 1.7951261634320892 1.5157e-08 1.7612682020397463 1.5158e-08 1.7996820744302382 1.5159e-08 1.8004455885102155 1.5159999999999998e-08 1.8132903672036293 1.5161e-08 1.8230322277990951 1.5162e-08 1.7180198187866147 1.5162999999999998e-08 1.7746049398968642 1.5164e-08 1.8450928838124887 1.5165e-08 1.745675175294977 1.5165999999999998e-08 1.783461355550142 1.5167e-08 1.7919420234179688 1.5168e-08 1.731907877436472 1.5169e-08 1.663684933413663 1.517e-08 1.813447164025215 1.5171e-08 1.7730887233746944 1.5172e-08 1.7541285613283262 1.5173e-08 1.8693313199073434 1.5174e-08 1.834554945402635 1.5175e-08 1.7620978565517196 1.5176e-08 1.8926306441513914 1.5177e-08 1.826328860459195 1.5178e-08 1.7374075641310682 1.5179e-08 1.8126780581889161 1.518e-08 1.8104518513963228 1.5181e-08 1.8126337044223737 1.5182e-08 1.6914173003926294 1.5183e-08 1.819823730796632 1.5184e-08 1.8071783342602865 1.5185e-08 1.733028459946925 1.5186e-08 1.749820893308594 1.5187e-08 1.8860633480598124 1.5188e-08 1.8385749987917788 1.5189e-08 1.8453454689732192 1.519e-08 1.8328607247227173 1.5191e-08 1.867962785689145 1.5192e-08 1.7714702382039285 1.5193e-08 1.7785066471153201 1.5194e-08 1.8003014799608101 1.5194999999999998e-08 1.734232177307973 1.5196e-08 1.7792463110471153 1.5197e-08 1.839111606726204 1.5197999999999998e-08 1.8010248450006054 1.5199e-08 1.8167409834705044 1.52e-08 1.8014761078946693 1.5200999999999998e-08 1.8058743175041458 1.5202e-08 1.7577691600606584 1.5203e-08 1.7785524660937746 1.5204e-08 1.7301059552946727 1.5205e-08 1.7686972110657733 1.5206e-08 1.7686958819873777 1.5207e-08 1.831765344505581 1.5208e-08 1.7964028580220581 1.5209e-08 1.7766748894694187 1.521e-08 1.7569985670407917 1.5211e-08 1.8842638835168624 1.5212e-08 1.8369402968663413 1.5213e-08 1.7280174777913255 1.5214e-08 1.7020849151385322 1.5215e-08 1.7595115990300823 1.5216e-08 1.7954610853582484 1.5217e-08 1.765165606541052 1.5218e-08 1.774531361683907 1.5219e-08 1.793757674555635 1.522e-08 1.8747584420784567 1.5221e-08 1.6983616482769401 1.5222e-08 1.7957478478789561 1.5223e-08 1.7219226214456231 1.5224e-08 1.8694585161468766 1.5225e-08 1.7730913123650218 1.5226e-08 1.7614150421879562 1.5227e-08 1.752502435114748 1.5228e-08 1.8119920873121327 1.5229e-08 1.8249079094465963 1.5229999999999998e-08 1.7927860706875072 1.5231e-08 1.8492936532174111 1.5232e-08 1.8712231171173326 1.5232999999999998e-08 1.804977584972434 1.5234e-08 1.793852373692884 1.5235e-08 1.8652191704298848 1.5235999999999998e-08 1.8279919627222176 1.5237e-08 1.9102841130881367 1.5238e-08 1.771223726717634 1.5239e-08 1.8375279398651885 1.524e-08 1.8105166616827324 1.5241e-08 1.7682695941068598 1.5242e-08 1.7288365669048682 1.5243e-08 1.7575665086324832 1.5244e-08 1.772058742495335 1.5245e-08 1.7801766349236863 1.5246e-08 1.7434998598805023 1.5247e-08 1.728999244219739 1.5248e-08 1.7554809225782024 1.5249e-08 1.7898935343535314 1.525e-08 1.8268095110843636 1.5251e-08 1.8740528695979843 1.5252e-08 1.8276447012214767 1.5253e-08 1.8715839236898524 1.5254e-08 1.7639983424537802 1.5255e-08 1.7420383057269824 1.5256e-08 1.8864658393849765 1.5257e-08 1.836350191268665 1.5258e-08 1.8036921628710845 1.5259e-08 1.8286351741933213 1.526e-08 1.8649902104142564 1.5261e-08 1.8494002667143044 1.5262e-08 1.8082714628652878 1.5263e-08 1.8363457275815824 1.5264e-08 1.8032611644652123 1.5264999999999998e-08 1.8940768714023075 1.5266e-08 1.7522424725274943 1.5267e-08 1.9060769254359076 1.5267999999999998e-08 1.8180549634576342 1.5269e-08 1.718838409732426 1.527e-08 1.7527893650829447 1.5270999999999998e-08 1.8688670512263104 1.5272e-08 1.8401263262351948 1.5273e-08 1.671122095778764 1.5273999999999998e-08 1.6995095057389487 1.5275e-08 1.8699989534480737 1.5276e-08 1.8186544983102322 1.5277e-08 1.7637596017020003 1.5278e-08 1.791043210513987 1.5279e-08 1.8735879254313668 1.528e-08 1.8607353755613183 1.5281e-08 1.788110729108819 1.5282e-08 1.8644129901294826 1.5283e-08 1.8217231796906304 1.5284e-08 1.896775059674955 1.5285e-08 1.7514731776149026 1.5286e-08 1.876783222922469 1.5287e-08 1.7853265699244525 1.5288e-08 1.8490449435257008 1.5289e-08 1.7478028187556742 1.529e-08 1.8555424926670157 1.5291e-08 1.7716857402732011 1.5292e-08 1.7265148737205513 1.5293e-08 1.6826563405913315 1.5294e-08 1.8592447464420556 1.5295e-08 1.8880408685607197 1.5296e-08 1.7706151242467 1.5297e-08 1.7600678510507861 1.5298e-08 1.7547624185295594 1.5299e-08 1.7720658764781914 1.53e-08 1.8077218392466172 1.5301e-08 1.8013362810685454 1.5302e-08 1.7872375584599953 1.5302999999999998e-08 1.8241557323239355 1.5304e-08 1.8266539313860195 1.5305e-08 1.7960046998212127 1.5305999999999998e-08 1.860664744270198 1.5307e-08 1.8531293544193368 1.5308e-08 1.8622899420304382 1.5308999999999998e-08 1.7074280257496193 1.531e-08 1.877360781808769 1.5311e-08 1.7732329039883326 1.5312e-08 1.7998609096715623 1.5313e-08 1.7993115147652994 1.5314e-08 1.827446102401207 1.5315e-08 1.7635428828198918 1.5316e-08 1.817749125278563 1.5317e-08 1.7658446691961966 1.5318e-08 1.7753206251918394 1.5319e-08 1.797984777292415 1.532e-08 1.7562242001490838 1.5321e-08 1.8874768620804625 1.5322e-08 1.799306697735891 1.5323e-08 1.8465033055267663 1.5324e-08 1.7668103611930295 1.5325e-08 1.714742775254255 1.5326e-08 1.7343232204714287 1.5327e-08 1.8648718811319722 1.5328e-08 1.8247680549028165 1.5329e-08 1.7031685942008523 1.533e-08 1.8835704001489013 1.5331e-08 1.8016994485886615 1.5332e-08 1.7162568398120024 1.5333e-08 1.7273688921476562 1.5334e-08 1.7968786846021343 1.5335e-08 1.7351330726282714 1.5336e-08 1.828192879967647 1.5337e-08 1.7459750886482852 1.5337999999999998e-08 1.8079801736650944 1.5339e-08 1.7699594072358382 1.534e-08 1.84349774432019 1.5340999999999998e-08 1.8425629488571553 1.5342e-08 1.8161708967938652 1.5343e-08 1.7204818371037445 1.5343999999999998e-08 1.9106773804210584 1.5345e-08 1.842257257939229 1.5346e-08 1.831142029758255 1.5347e-08 1.8398859058061334 1.5348e-08 1.7707924444210115 1.5349e-08 1.8081444786788625 1.535e-08 1.8949378787431919 1.5351e-08 1.797655087495361 1.5352e-08 1.8696909300544935 1.5353e-08 1.876403985377472 1.5354e-08 1.8706555713604345 1.5355e-08 1.7877751800407857 1.5356e-08 1.901967067870979 1.5357e-08 1.6645944877259997 1.5358e-08 1.876660060090148 1.5359e-08 1.8865881294908444 1.536e-08 1.730782738492351 1.5361e-08 1.8327207136408163 1.5362e-08 1.758194415565962 1.5363e-08 1.8312802903195062 1.5364e-08 1.721181895318446 1.5365e-08 1.7985851012262115 1.5366e-08 1.7981985311102082 1.5367e-08 1.7950073993797184 1.5368e-08 1.7160115173370625 1.5369e-08 1.885522430143895 1.537e-08 1.8160223889631846 1.5371e-08 1.8555842481097515 1.5372e-08 1.8131448576460247 1.5372999999999998e-08 1.8156551970301604 1.5374e-08 1.8228212228059586 1.5375e-08 1.8238643585810923 1.5375999999999998e-08 1.7496492129666847 1.5377e-08 1.7876855544580263 1.5378e-08 1.8032668421257272 1.5378999999999998e-08 1.8322282720145786 1.538e-08 1.791561009325906 1.5381e-08 1.7575992090047992 1.5382e-08 1.8240401062047078 1.5383e-08 1.7765280772063006 1.5384e-08 1.7997946942056267 1.5385e-08 1.8216216173027595 1.5386e-08 1.8219812413361662 1.5387e-08 1.8332716713493837 1.5388e-08 1.7441205262671318 1.5389e-08 1.80060003952421 1.539e-08 1.7834968324463094 1.5391e-08 1.8104996995338556 1.5392e-08 1.74065463632546 1.5393e-08 1.8047557208171054 1.5394e-08 1.8821962719129495 1.5395e-08 1.831332256426876 1.5396e-08 1.8079095398009335 1.5397e-08 1.806734903990436 1.5398e-08 1.8045197334663712 1.5399e-08 1.804387815868858 1.54e-08 1.6965857914561475 1.5401e-08 1.7561954353061877 1.5402e-08 1.7776770546473728 1.5403e-08 1.840449549244964 1.5404e-08 1.7693333437874221 1.5405e-08 1.8358251346160286 1.5406e-08 1.8111679684751787 1.5407e-08 1.7540417015275145 1.5407999999999998e-08 1.8230614413153494 1.5409e-08 1.7133654293349814 1.541e-08 1.7661629573700046 1.5410999999999998e-08 1.8277054075135235 1.5412e-08 1.7535893514023164 1.5413e-08 1.7515023254435065 1.5413999999999998e-08 1.8495882576806975 1.5415e-08 1.8091330258741827 1.5416e-08 1.8834852672667306 1.5417e-08 1.7891101187127378 1.5418e-08 1.855868124147321 1.5419e-08 1.7836072946088681 1.542e-08 1.845857379292455 1.5421e-08 1.7512980765513393 1.5422e-08 1.7394904614394555 1.5423e-08 1.923604047930832 1.5424e-08 1.7704415247983032 1.5425e-08 1.802889150500651 1.5426e-08 1.734602135438545 1.5427e-08 1.6974786045142418 1.5428e-08 1.7722411111156775 1.5429e-08 1.774239356445914 1.543e-08 1.7967332114916525 1.5431e-08 1.7667985081688962 1.5432e-08 1.6598784098370951 1.5433e-08 1.756082258094877 1.5434e-08 1.9035953762441573 1.5435e-08 1.8723455138956155 1.5436e-08 1.83126357839619 1.5437e-08 1.8724722576826212 1.5438e-08 1.786645009541265 1.5439e-08 1.8651605605120658 1.544e-08 1.7760618543477882 1.5441e-08 1.8396106548676974 1.5442e-08 1.845291070290716 1.5442999999999998e-08 1.8045740720761614 1.5444e-08 1.8383766468295097 1.5445e-08 1.8860665944833142 1.5445999999999998e-08 1.8703460394306366 1.5447e-08 1.8429897563646334 1.5448e-08 1.8330586652071637 1.5448999999999998e-08 1.7228138025713047 1.545e-08 1.792179716105424 1.5451e-08 1.7657625722209143 1.5451999999999998e-08 1.8501083887667062 1.5453e-08 1.858820976423082 1.5454e-08 1.7856753139559924 1.5455e-08 1.7495955336615971 1.5456e-08 1.8356132923385036 1.5457e-08 1.8273317803544058 1.5458e-08 1.844266656000908 1.5459e-08 1.8297346185030094 1.546e-08 1.8226727739229196 1.5461e-08 1.771549712053124 1.5462e-08 1.742393346011617 1.5463e-08 1.7883847179100172 1.5464e-08 1.891633472088603 1.5465e-08 1.82986802085596 1.5466e-08 1.8716020145028112 1.5467e-08 1.8055898733676259 1.5468e-08 1.8120046348198688 1.5469e-08 1.836689682245425 1.547e-08 1.817090256189811 1.5471e-08 1.7806028189571057 1.5472e-08 1.7250816442132297 1.5473e-08 1.8800303854769598 1.5474e-08 1.7723715276085552 1.5475e-08 1.8298774512189544 1.5476e-08 1.8057828526761504 1.5477e-08 1.7841098247041691 1.5477999999999998e-08 1.8904996070674545 1.5479e-08 1.7145823223835974 1.548e-08 1.7656249990158617 1.5480999999999998e-08 1.7777948467672307 1.5482e-08 1.8272800054322142 1.5483e-08 1.8730430904989448 1.5483999999999998e-08 1.6699962834091897 1.5485e-08 1.8569476173639505 1.5486e-08 1.8200008242067602 1.5486999999999998e-08 1.8373302741668966 1.5488e-08 1.8603206919448225 1.5489e-08 1.802546347558253 1.549e-08 1.8430397458193633 1.5491e-08 1.7350927762495822 1.5492e-08 1.875049741406309 1.5493e-08 1.7750337216982588 1.5494e-08 1.7721672264990715 1.5495e-08 1.7870594736091534 1.5496e-08 1.8419438879147167 1.5497e-08 1.7490459593190724 1.5498e-08 1.8906923225952135 1.5499e-08 1.8007633066678381 1.55e-08 1.8194524245259647 1.5501e-08 1.7473951986325333 1.5502e-08 1.8195891291567303 1.5503e-08 1.7723955840669627 1.5504e-08 1.906888463735621 1.5505e-08 1.7494613273394373 1.5506e-08 1.7821897389477066 1.5507e-08 1.803895426186481 1.5508e-08 1.708624896832248 1.5509e-08 1.8291227979674756 1.551e-08 1.8753533454788016 1.5511e-08 1.7973031481041502 1.5512e-08 1.7779138590981396 1.5513e-08 1.845251152670699 1.5514e-08 1.7805078836317754 1.5515e-08 1.75908334909054 1.5515999999999998e-08 1.7553220633886124 1.5517e-08 1.7757684701501137 1.5518e-08 1.928041798139306 1.5518999999999998e-08 1.8806165686479657 1.552e-08 1.7697780641454024 1.5521e-08 1.8323126101485068 1.5521999999999998e-08 1.7825791641356235 1.5523e-08 1.8007810154706099 1.5524e-08 1.754404057814501 1.5525e-08 1.8106948164224494 1.5526e-08 1.8989987384701403 1.5527e-08 1.8086799452070874 1.5528e-08 1.7728530482890927 1.5529e-08 1.818430178905097 1.553e-08 1.8208517627557015 1.5531e-08 1.799030167839865 1.5532e-08 1.8503572292216242 1.5533e-08 1.7510099373155725 1.5534e-08 1.8646605981656093 1.5535e-08 1.806879113670158 1.5536e-08 1.7340266462825615 1.5537e-08 1.8760334952617117 1.5538e-08 1.788124181429043 1.5539e-08 1.9147239878882476 1.554e-08 1.7925210063433938 1.5541e-08 1.8071679905258735 1.5542e-08 1.7522903550656383 1.5543e-08 1.76198087358646 1.5544e-08 1.797837913070908 1.5545e-08 1.8629217549065766 1.5546e-08 1.7530726597704411 1.5547e-08 1.7980918413221905 1.5548e-08 1.747041555250879 1.5549e-08 1.8627120567309616 1.555e-08 1.8203597239967175 1.5550999999999998e-08 1.7909603133107022 1.5552e-08 1.7612409961808833 1.5553e-08 1.8416315519485327 1.5553999999999998e-08 1.775258345450228 1.5555e-08 1.8042229275563473 1.5556e-08 1.8550585134920126 1.5556999999999998e-08 1.8126821130239095 1.5558e-08 1.7089101162611076 1.5559e-08 1.7737916483330547 1.556e-08 1.7969812415846058 1.5561e-08 1.685232674809738 1.5562e-08 1.8034606657011387 1.5563e-08 1.7672683039824277 1.5564e-08 1.726156964307336 1.5565e-08 1.7707815437841417 1.5566e-08 1.7880897520612629 1.5567e-08 1.7766433274471638 1.5568e-08 1.8469631153426729 1.5569e-08 1.7398514206108129 1.557e-08 1.8321369620420502 1.5571e-08 1.9132655540063772 1.5572e-08 1.8578680634379863 1.5573e-08 1.7751809225474062 1.5574e-08 1.8768619542445502 1.5575e-08 1.8001842751333919 1.5576e-08 1.8219910181149968 1.5577e-08 1.8415169925759458 1.5578e-08 1.9001776330308033 1.5579e-08 1.7260704812058847 1.558e-08 1.8842803604266314 1.5581e-08 1.775511426501323 1.5582e-08 1.7982000138356293 1.5583e-08 1.830213587825133 1.5584e-08 1.8041467934152158 1.5585e-08 1.7734268760443326 1.5585999999999998e-08 1.78947199431228 1.5587e-08 1.8395594545978078 1.5588e-08 1.785757917799305 1.5588999999999998e-08 1.8340174102953994 1.559e-08 1.8257843875492783 1.5591e-08 1.747504856451258 1.5591999999999998e-08 1.7584270118795204 1.5593e-08 1.7147025873689226 1.5594e-08 1.8380947929832818 1.5595e-08 1.7510691592793861 1.5596e-08 1.8134436783793013 1.5597e-08 1.7565728763268287 1.5598e-08 1.7670103801238444 1.5599e-08 1.758681535839765 1.56e-08 1.7820883296237917 1.5601e-08 1.6987983344343807 1.5602e-08 1.8251879835957117 1.5603e-08 1.792037163574082 1.5604e-08 1.8226110330809233 1.5605e-08 1.7678457159399628 1.5606e-08 1.817297302343221 1.5607e-08 1.8246204212370292 1.5608e-08 1.732324450124791 1.5609e-08 1.7318593826823718 1.561e-08 1.7264515342367956 1.5611e-08 1.7978039754003479 1.5612e-08 1.7844557070158265 1.5613e-08 1.7630121115631168 1.5614e-08 1.7407612867221904 1.5615e-08 1.8168528718329124 1.5616e-08 1.7096347081182055 1.5617e-08 1.8050976729389543 1.5618e-08 1.7855835396803064 1.5619e-08 1.8270891541105416 1.562e-08 1.7676575360260418 1.5620999999999998e-08 1.7865048304321167 1.5622e-08 1.784282466649286 1.5623e-08 1.8146607652596112 1.5623999999999998e-08 1.7652640703340334 1.5625e-08 1.7840554626476681 1.5626e-08 1.7152940255635662 1.5626999999999998e-08 1.8365891267502565 1.5628e-08 1.8354867597753324 1.5629e-08 1.8424930595992077 1.5629999999999998e-08 1.8211366437873628 1.5631e-08 1.7457656624624407 1.5632e-08 1.8364962074563627 1.5633e-08 1.911022216312333 1.5634e-08 1.846074401046177 1.5635e-08 1.9100126301372162 1.5636e-08 1.8752350453179865 1.5637e-08 1.7313171427377232 1.5638e-08 1.7931247354121127 1.5639e-08 1.7537982376723125 1.564e-08 1.7891667193123295 1.5641e-08 1.7418223508821162 1.5642e-08 1.798054427115973 1.5643e-08 1.8497428959107842 1.5644e-08 1.79040502133126 1.5645e-08 1.7373327063140251 1.5646e-08 1.8745427576872302 1.5647e-08 1.8150995914118377 1.5648e-08 1.8631976594728337 1.5649e-08 1.8822933360231475 1.565e-08 1.8149319245971356 1.5651e-08 1.8059365561976828 1.5652e-08 1.702547157272139 1.5653e-08 1.6986011734304105 1.5654e-08 1.8021342277063193 1.5655e-08 1.858650020565607 1.5655999999999998e-08 1.857149971380366 1.5657e-08 1.884557638251764 1.5658e-08 1.7945435220760801 1.5658999999999998e-08 1.9057239218842101 1.566e-08 1.820620606562613 1.5661e-08 1.848996295003781 1.5661999999999998e-08 1.8110143113569572 1.5663e-08 1.7817825873972568 1.5664e-08 1.865127689193563 1.5664999999999998e-08 1.9193299970607887 1.5666e-08 1.852384729774007 1.5667e-08 1.789657133499666 1.5668e-08 1.740282859537146 1.5669e-08 1.7558151613130162 1.567e-08 1.7487027127026127 1.5671e-08 1.8183508719822536 1.5672e-08 1.8225429451947779 1.5673e-08 1.8899506430507815 1.5674e-08 1.7913766693261213 1.5675e-08 1.8767278632475206 1.5676e-08 1.8421522804637247 1.5677e-08 1.8872807226177397 1.5678e-08 1.8581133615330137 1.5679e-08 1.727317327992724 1.568e-08 1.746315956678006 1.5681e-08 1.7636369354799255 1.5682e-08 1.8306333284837342 1.5683e-08 1.8380216430910252 1.5684e-08 1.8105443966873362 1.5685e-08 1.8463557139436562 1.5686e-08 1.9041759759200785 1.5687e-08 1.827719082440193 1.5688e-08 1.8465219165101487 1.5689e-08 1.765361412242927 1.569e-08 1.762070905034433 1.5690999999999998e-08 1.7405332611861575 1.5692e-08 1.774087060861683 1.5693e-08 1.807061488077362 1.5693999999999998e-08 1.7717602822404763 1.5695e-08 1.7352968424775215 1.5696e-08 1.8129287236449747 1.5696999999999998e-08 1.7748594841108332 1.5698e-08 1.808270712977909 1.5699e-08 1.8527938285116399 1.5699999999999998e-08 1.8381068741252067 1.5701e-08 1.8377790198283421 1.5702e-08 1.8107506864517355 1.5703e-08 1.7459166184287338 1.5704e-08 1.830869800414137 1.5705e-08 1.7806126081680835 1.5706e-08 1.904719729919301 1.5707e-08 1.8966832325073737 1.5708e-08 1.7781971056615928 1.5709e-08 1.8565071783004314 1.571e-08 1.7443425897933902 1.5711e-08 1.885440665041649 1.5712e-08 1.7942979668818506 1.5713e-08 1.7785689231499748 1.5714e-08 1.8556620866385911 1.5715e-08 1.8065414919515366 1.5716e-08 1.8292867085862912 1.5717e-08 1.6982307174070939 1.5718e-08 1.7888078498728441 1.5719e-08 1.790400913743614 1.572e-08 1.777932701391804 1.5721e-08 1.8829276430242634 1.5722e-08 1.9256752590065993 1.5723e-08 1.8387986773493101 1.5724e-08 1.815181421998943 1.5725e-08 1.782735247090296 1.5726e-08 1.8000013903350338 1.5727e-08 1.8215625086390055 1.5728e-08 1.8433781942930991 1.5728999999999998e-08 1.8070588137464285 1.573e-08 1.8200586396030731 1.5731e-08 1.774993982462823 1.5731999999999998e-08 1.8734412816245924 1.5733e-08 1.7325861324682434 1.5734e-08 1.7973266416027356 1.5734999999999998e-08 1.879298114069162 1.5736e-08 1.7594510926481055 1.5737e-08 1.7533982413270455 1.5738e-08 1.7662522675170789 1.5739e-08 1.7546340467147612 1.574e-08 1.85157932619426 1.5741e-08 1.8388953434833617 1.5742e-08 1.8382650210502218 1.5743e-08 1.8197252469869851 1.5744e-08 1.8941393574591292 1.5745e-08 1.8085994748185161 1.5746e-08 1.9120698503413602 1.5747e-08 1.8091711937542232 1.5748e-08 1.783118416664675 1.5749e-08 1.7601291966330799 1.575e-08 1.8035559826192922 1.5751e-08 1.8404020730528983 1.5752e-08 1.759046777785836 1.5753e-08 1.850336319512575 1.5754e-08 1.7666784090381822 1.5755e-08 1.778169643201259 1.5756e-08 1.846219818753772 1.5757e-08 1.7759098945747622 1.5758e-08 1.7502163856796302 1.5759e-08 1.841867278063448 1.576e-08 1.746147717625875 1.5761e-08 1.8280039469182106 1.5762e-08 1.8144633741393452 1.5763e-08 1.7844362588276612 1.5763999999999998e-08 1.8089280848977074 1.5765e-08 1.8355700234146093 1.5766e-08 1.8013105264256228 1.5766999999999998e-08 1.848375585029254 1.5768e-08 1.817910512679739 1.5769e-08 1.7699314569701432 1.5769999999999998e-08 1.8472741766533942 1.5771e-08 1.7506754227860308 1.5772e-08 1.847365762422182 1.5773e-08 1.836406958565489 1.5774e-08 1.7730981023569627 1.5775e-08 1.8307039618993863 1.5776e-08 1.786727506584395 1.5777e-08 1.830782685295231 1.5778e-08 1.8595988206866068 1.5779e-08 1.749486396317179 1.578e-08 1.810110836941653 1.5781e-08 1.7194095887869498 1.5782e-08 1.8307715003744365 1.5783e-08 1.8573918617445724 1.5784e-08 1.766345163513563 1.5785e-08 1.7184321669700873 1.5786e-08 1.7872212042328544 1.5787e-08 1.7500347952108064 1.5788e-08 1.8427286384713737 1.5789e-08 1.7661716904353357 1.579e-08 1.882681647986969 1.5791e-08 1.8428772287262847 1.5792e-08 1.7681531180483412 1.5793e-08 1.9181663359391288 1.5794e-08 1.8125578101235178 1.5795e-08 1.7944736819181333 1.5796e-08 1.7899768519934942 1.5797e-08 1.8105704480641867 1.5798e-08 1.806234517314578 1.5798999999999998e-08 1.8165084135830976 1.58e-08 1.8589055296636803 1.5801e-08 1.7710727632123429 1.5801999999999998e-08 1.8224743770785514 1.5803e-08 1.8227509280474306 1.5804e-08 1.867409030530443 1.5804999999999998e-08 1.8921064377210397 1.5806e-08 1.7576520370488578 1.5807e-08 1.9030260981317118 1.5808e-08 1.8208125251316751 1.5809e-08 1.8124756203071606 1.581e-08 1.7536726732118333 1.5811e-08 1.8245439809066535 1.5812e-08 1.7896696944001362 1.5813e-08 1.8890221440731232 1.5814e-08 1.667756651073391 1.5815e-08 1.7909363940115066 1.5816e-08 1.7568865426754352 1.5817e-08 1.7937575785140807 1.5818e-08 1.826318155913562 1.5819e-08 1.7695152257892477 1.582e-08 1.7518415747716436 1.5821e-08 1.8205132703538967 1.5822e-08 1.7864799887807963 1.5823e-08 1.7861641019912295 1.5824e-08 1.852825389473172 1.5825e-08 1.778900816298069 1.5826e-08 1.8301569331575693 1.5827e-08 1.8600342034048774 1.5828e-08 1.7984872194302792 1.5829e-08 1.7705591025497114 1.583e-08 1.821471738161993 1.5831e-08 1.7551985658034992 1.5832e-08 1.7951283258484283 1.5833e-08 1.716211079402853 1.5833999999999998e-08 1.7909979281090171 1.5835e-08 1.7873391258462268 1.5836e-08 1.7335893537921405 1.5836999999999998e-08 1.836691363325822 1.5838e-08 1.8048688452649313 1.5839e-08 1.8043733514950606 1.5839999999999998e-08 1.842718116285085 1.5841e-08 1.8132811063004117 1.5842e-08 1.7656762791253202 1.5842999999999998e-08 1.7529701100284896 1.5844e-08 1.794645161178718 1.5845e-08 1.8361202524799423 1.5846e-08 1.7359080556131627 1.5847e-08 1.834641344449864 1.5848e-08 1.797075445988228 1.5849e-08 1.8693341320427337 1.585e-08 1.765641799761735 1.5851e-08 1.7977279747710344 1.5852e-08 1.8794278702130778 1.5853e-08 1.84631663019396 1.5854e-08 1.7684574907018833 1.5855e-08 1.8166169475733214 1.5856e-08 1.812479907244169 1.5857e-08 1.812236181623159 1.5858e-08 1.81282183287252 1.5859e-08 1.835176989999841 1.586e-08 1.6991706967371452 1.5861e-08 1.825069901195593 1.5862e-08 1.7769441560118335 1.5863e-08 1.8117519416912622 1.5864e-08 1.6650360693558468 1.5865e-08 1.8604156520530835 1.5866e-08 1.836469384326091 1.5867e-08 1.8035419695936699 1.5868e-08 1.794558664993639 1.5868999999999998e-08 1.7872728221812237 1.587e-08 1.804096406403076 1.5871e-08 1.8341642416745718 1.5871999999999998e-08 1.83402447501276 1.5873e-08 1.845160960702394 1.5874e-08 1.7817019417959257 1.5874999999999998e-08 1.818909114114768 1.5876e-08 1.7256400398121001 1.5877e-08 1.7771454179829742 1.5877999999999998e-08 1.7614887438361804 1.5879e-08 1.8164718082472207 1.588e-08 1.8316795540853552 1.5881e-08 1.8229231197376998 1.5882e-08 1.8685254532402908 1.5883e-08 1.7917811369149366 1.5884e-08 1.8001988073699309 1.5885e-08 1.9100322661940967 1.5886e-08 1.7107784494139784 1.5887e-08 1.7154734006334689 1.5888e-08 1.860266207407282 1.5889e-08 1.8379156571173585 1.589e-08 1.8629960296409152 1.5891e-08 1.8849762663883 1.5892e-08 1.8181964628984546 1.5893e-08 1.7574142347777766 1.5894e-08 1.8593160679825478 1.5895e-08 1.7586433187578259 1.5896e-08 1.7958242143962972 1.5897e-08 1.7344253936917549 1.5898e-08 1.7840100651761195 1.5899e-08 1.8398515950002006 1.59e-08 1.8248462329303332 1.5901e-08 1.7661352633175031 1.5902e-08 1.7952898644190984 1.5903e-08 1.7843534706781259 1.5904e-08 1.854491522101596 1.5905e-08 1.8038559568897143 1.5906e-08 1.8909469092243145 1.5906999999999998e-08 1.80135601331003 1.5908e-08 1.6922433698781318 1.5909e-08 1.819715548884736 1.5909999999999998e-08 1.8157388341332805 1.5911e-08 1.7785702417309828 1.5912e-08 1.8076224921994353 1.5912999999999998e-08 1.8499051093348151 1.5914e-08 1.7571072394139997 1.5915e-08 1.8086902391177946 1.5916e-08 1.7854322790596713 1.5917e-08 1.705295332695195 1.5918e-08 1.7865100322451108 1.5919e-08 1.7558446564545382 1.592e-08 1.7754434610406342 1.5921e-08 1.7916088090030977 1.5922e-08 1.7326223045030051 1.5923e-08 1.7718924038549284 1.5924e-08 1.881379709671168 1.5925e-08 1.7851830893711396 1.5926e-08 1.7495515013576837 1.5927e-08 1.8065812911732448 1.5928e-08 1.7536920475269313 1.5929e-08 1.7204834564368556 1.593e-08 1.786899979100514 1.5931e-08 1.8080293442394308 1.5932e-08 1.7482942521666198 1.5933e-08 1.7699130672973535 1.5934e-08 1.8108686855918705 1.5935e-08 1.8382776825728278 1.5936e-08 1.9189297824718163 1.5937e-08 1.7381054001746568 1.5938e-08 1.7896600479158178 1.5939e-08 1.7795415001839028 1.594e-08 1.8751415484386433 1.5941e-08 1.84224501925659 1.5941999999999998e-08 1.7788635595832347 1.5943e-08 1.8102008966952052 1.5944e-08 1.7499243691465638 1.5944999999999998e-08 1.7514199633274143 1.5946e-08 1.8312880661141693 1.5947e-08 1.804012132950653 1.5947999999999998e-08 1.8348466880913543 1.5949e-08 1.842304154982452 1.595e-08 1.7831491416309162 1.5951e-08 1.7946988947542775 1.5952e-08 1.812557998298333 1.5953e-08 1.8889637545659868 1.5954e-08 1.737124502809247 1.5955e-08 1.9013928309836772 1.5956e-08 1.7404555872126122 1.5957e-08 1.7603917045532211 1.5958e-08 1.804423359647243 1.5959e-08 1.7830428300017414 1.596e-08 1.8584336979988145 1.5961e-08 1.850412595686332 1.5962e-08 1.8366689582095415 1.5963e-08 1.6741234243827852 1.5964e-08 1.7876766295086928 1.5965e-08 1.7818633239503323 1.5966e-08 1.8420429741587094 1.5967e-08 1.8469543394812256 1.5968e-08 1.721396482832637 1.5969e-08 1.8539125620730421 1.597e-08 1.7673589930733389 1.5971e-08 1.7794950995207466 1.5972e-08 1.7189388015763474 1.5973e-08 1.8127553508816054 1.5974e-08 1.8054283418034516 1.5975e-08 1.8284156477803473 1.5976e-08 1.7733408957174521 1.5976999999999998e-08 1.8489521648806932 1.5978e-08 1.7539702244302002 1.5979e-08 1.8430063219761301 1.5979999999999998e-08 1.7582075052449293 1.5981e-08 1.7703391250919918 1.5982e-08 1.7627805200696274 1.5982999999999998e-08 1.8945299000752478 1.5984e-08 1.7037250704726934 1.5985e-08 1.852129969949306 1.5986e-08 1.723392923842705 1.5987e-08 1.8065884900817686 1.5988e-08 1.82676370677879 1.5989e-08 1.8446016380359027 1.599e-08 1.870637319847161 1.5991e-08 1.707837065009033 1.5992e-08 1.744137144651151 1.5993e-08 1.8688576054743344 1.5994e-08 1.7329842511397806 1.5995e-08 1.7943722076131334 1.5996e-08 1.7256007925358137 1.5997e-08 1.8464266298365377 1.5998e-08 1.8068395954902028 1.5999e-08 1.8271879764877708 1.6e-08 1.7518357692304523 1.6001e-08 1.843549026145485 1.6002e-08 1.8701534032681466 1.6003e-08 1.7594352650216272 1.6004e-08 1.7992365983909047 1.6005e-08 1.8212711927826708 1.6006e-08 1.8106942690568282 1.6007e-08 1.7688061473461918 1.6008e-08 1.8056905813757242 1.6009e-08 1.7921863450401705 1.601e-08 1.8094894482785011 1.6011e-08 1.7620028408764064 1.6011999999999998e-08 1.7849158275653842 1.6013e-08 1.798733255481029 1.6014e-08 1.7952200613550926 1.6014999999999998e-08 1.7742486336117176 1.6016e-08 1.8586335924154125 1.6017e-08 1.8306253122957101 1.6017999999999998e-08 1.7773467273452606 1.6019e-08 1.7762605470062804 1.602e-08 1.7980266438432984 1.6020999999999998e-08 1.801870106642909 1.6022e-08 1.6909976538181781 1.6023e-08 1.9138995097568123 1.6024e-08 1.8699988122128113 1.6025e-08 1.7842413095356604 1.6026e-08 1.7648783096218301 1.6027e-08 1.751026875100709 1.6028e-08 1.7633003362421114 1.6029e-08 1.825101600978016 1.603e-08 1.7891922574260541 1.6031e-08 1.8485413431152482 1.6032e-08 1.8437673038872209 1.6033e-08 1.808313760345726 1.6034e-08 1.72580121060693 1.6035e-08 1.7618677387449038 1.6036e-08 1.8100965097296045 1.6037e-08 1.8530855116257259 1.6038e-08 1.8732800271695764 1.6039e-08 1.8460897904839306 1.604e-08 1.8889682562522656 1.6041e-08 1.8898701318380167 1.6042e-08 1.8030778196486439 1.6043e-08 1.7835219932693522 1.6044e-08 1.834333994631354 1.6045e-08 1.8189053510197004 1.6046e-08 1.740405857043414 1.6046999999999998e-08 1.7967055873522484 1.6048e-08 1.8439457138982813 1.6049e-08 1.742729698498174 1.6049999999999998e-08 1.8185761980574193 1.6051e-08 1.7521297823979114 1.6052e-08 1.7376521385715589 1.6052999999999998e-08 1.7568685055741533 1.6054e-08 1.7493643950048126 1.6055e-08 1.8350599835612915 1.6055999999999998e-08 1.7341170923795686 1.6057e-08 1.7820361766116595 1.6058e-08 1.8357400206895658 1.6059e-08 1.8454181627022763 1.606e-08 1.8479269615937228 1.6061e-08 1.812264746064227 1.6062e-08 1.7034699669038254 1.6063e-08 1.8185918981188154 1.6064e-08 1.8252478654891864 1.6065e-08 1.6577990421722801 1.6066e-08 1.8017086445500132 1.6067e-08 1.811745140021176 1.6068e-08 1.8118359764730803 1.6069e-08 1.7554061914458114 1.607e-08 1.7979589934318747 1.6071e-08 1.836133055539105 1.6072e-08 1.8142931673789076 1.6073e-08 1.7370856570272302 1.6074e-08 1.799862510422193 1.6075e-08 1.8739546200721047 1.6076e-08 1.7813219320444618 1.6077e-08 1.844440039549318 1.6078e-08 1.805735650275532 1.6079e-08 1.7364936463180827 1.608e-08 1.827990396508382 1.6081e-08 1.8321616198090254 1.6081999999999998e-08 1.898137529817839 1.6083e-08 1.7406321609073938 1.6084e-08 1.8767151717981012 1.6084999999999998e-08 1.7935361721016945 1.6086e-08 1.8269297849218793 1.6087e-08 1.8663749518231247 1.6087999999999998e-08 1.812158247442514 1.6089e-08 1.8410183842856753 1.609e-08 1.8743801378664067 1.6090999999999998e-08 1.8838334342238927 1.6092e-08 1.8298418104964398 1.6093e-08 1.7641385573125181 1.6094e-08 1.8184425723112465 1.6095e-08 1.802337365889308 1.6096e-08 1.751895645782906 1.6097e-08 1.8785003261963056 1.6098e-08 1.8392990236210742 1.6099e-08 1.8281632546703785 1.61e-08 1.8075109925080148 1.6101e-08 1.8219973171918356 1.6102e-08 1.8048279562217526 1.6103e-08 1.8766978096592184 1.6104e-08 1.7538134471716478 1.6105e-08 1.7324460983735455 1.6106e-08 1.7950965542390385 1.6107e-08 1.8164557317006242 1.6108e-08 1.7843612592649718 1.6109e-08 1.9145401583742954 1.611e-08 1.7747655771428337 1.6111e-08 1.8092413084756058 1.6112e-08 1.8186840664269106 1.6113e-08 1.9009328509066874 1.6114e-08 1.779529163608892 1.6115e-08 1.7779179851710825 1.6116e-08 1.8117893636755344 1.6117e-08 1.7554533255064897 1.6118e-08 1.8331346794722798 1.6119e-08 1.8601447575046635 1.6119999999999998e-08 1.7963091911764788 1.6121e-08 1.7283142189930791 1.6122e-08 1.827393196165671 1.6122999999999998e-08 1.76645287384559 1.6124e-08 1.8040119124750504 1.6125e-08 1.823503104816613 1.6125999999999998e-08 1.733860901667411 1.6127e-08 1.7870784614580455 1.6128e-08 1.8593931575984566 1.6129e-08 1.747063168041985 1.613e-08 1.7725286317589921 1.6131e-08 1.8706733299247373 1.6132e-08 1.8336900170589505 1.6133e-08 1.714025270929381 1.6134e-08 1.7767180586471227 1.6135e-08 1.7797589055238783 1.6136e-08 1.7116222675847785 1.6137e-08 1.8773350032053184 1.6138e-08 1.74272757640529 1.6139e-08 1.7786170755252344 1.614e-08 1.74357932340258 1.6141e-08 1.7670265915892862 1.6142e-08 1.8657217509618058 1.6143e-08 1.7437327233674997 1.6144e-08 1.8467404508092553 1.6145e-08 1.706676139456906 1.6146e-08 1.76269360532117 1.6147e-08 1.8719763758950436 1.6148e-08 1.8487377177315345 1.6149e-08 1.7518451722598138 1.615e-08 1.712836878855496 1.6151e-08 1.7647880886173966 1.6152e-08 1.783217132988149 1.6153e-08 1.8230205164739135 1.6154e-08 1.8132527599187118 1.6154999999999998e-08 1.8370127166370167 1.6156e-08 1.8125453003983931 1.6157e-08 1.817159912040225 1.6157999999999998e-08 1.708169499369592 1.6159e-08 1.7611014312099047 1.616e-08 1.7978761251341984 1.6160999999999998e-08 1.8590135433646096 1.6162e-08 1.8103224720058846 1.6163e-08 1.8683598066578697 1.6164e-08 1.7706210679006495 1.6165e-08 1.8014386857483715 1.6166e-08 1.8436460040669835 1.6167e-08 1.9039385521112913 1.6168e-08 1.8956588388804885 1.6169e-08 1.8300874643749998 1.617e-08 1.7997843482743903 1.6171e-08 1.783680088957913 1.6172e-08 1.8663544087452855 1.6173e-08 1.7871622899598387 1.6174e-08 1.8889577335012881 1.6175e-08 1.7372523229046606 1.6176e-08 1.7918908767811834 1.6177e-08 1.7555342267793765 1.6178e-08 1.8078491662963934 1.6179e-08 1.731347683021953 1.618e-08 1.8262236767876157 1.6181e-08 1.742544869563201 1.6182e-08 1.8457796546511076 1.6183e-08 1.7987424886698244 1.6184e-08 1.7420524965566355 1.6185e-08 1.902645433456271 1.6186e-08 1.766458436606977 1.6187e-08 1.7557906821198568 1.6188e-08 1.7451295293799958 1.6189e-08 1.8820719250897058 1.6189999999999998e-08 1.7702811120287236 1.6191e-08 1.8564482460361038 1.6192e-08 1.828198295028077 1.6192999999999998e-08 1.733693227336845 1.6194e-08 1.806543380778922 1.6195e-08 1.8228927631927272 1.6195999999999998e-08 1.871782819815543 1.6197e-08 1.703251358380246 1.6198e-08 1.7664455644065544 1.6198999999999998e-08 1.8735923245840111 1.62e-08 1.828161923708811 1.6201e-08 1.6872539821897277 1.6202e-08 1.8854426876604913 1.6203e-08 1.8049971374678166 1.6204e-08 1.814938463921689 1.6205e-08 1.9030050483905017 1.6206e-08 1.742919301920446 1.6207e-08 1.811236360218649 1.6208e-08 1.8463744096208066 1.6209e-08 1.7377358858325567 1.621e-08 1.7987414766700511 1.6211e-08 1.7965672213781 1.6212e-08 1.829330727866565 1.6213e-08 1.7866566691598222 1.6214e-08 1.7783770517368047 1.6215e-08 1.8531397116160535 1.6216e-08 1.7339892267146626 1.6217e-08 1.8303676683830497 1.6218e-08 1.7417464509427905 1.6219e-08 1.8160430846272206 1.622e-08 1.7360085252209465 1.6221e-08 1.7445793504865645 1.6222e-08 1.8361808485044901 1.6223e-08 1.759694095121876 1.6224e-08 1.8536947097703644 1.6224999999999998e-08 1.8525578352137364 1.6226e-08 1.7680307476302946 1.6227e-08 1.8131808058785215 1.6227999999999998e-08 1.8812898034196583 1.6229e-08 1.8295793176582396 1.623e-08 1.771130898596784 1.6230999999999998e-08 1.7815223795214241 1.6232e-08 1.865148968283795 1.6233e-08 1.846712349008862 1.6233999999999998e-08 1.8282276503791948 1.6235e-08 1.7637294836756858 1.6236e-08 1.7370345391473556 1.6237e-08 1.756197712592794 1.6238e-08 1.8003037011056802 1.6239e-08 1.8330414364201897 1.624e-08 1.818625856764801 1.6241e-08 1.7506942922396258 1.6242e-08 1.7975728115443392 1.6243e-08 1.820991790732614 1.6244e-08 1.8302152157324034 1.6245e-08 1.7334243701821714 1.6246e-08 1.6535176930685476 1.6247e-08 1.7864425321525914 1.6248e-08 1.7571803381061468 1.6249e-08 1.711601078316183 1.625e-08 1.8357884561061784 1.6251e-08 1.7101058978531154 1.6252e-08 1.7609369183057624 1.6253e-08 1.836483211378012 1.6254e-08 1.8255729923787463 1.6255e-08 1.8435366667929496 1.6256e-08 1.8846156140933168 1.6257e-08 1.787052222886125 1.6258e-08 1.7729215971160213 1.6259e-08 1.7864269983989447 1.6259999999999998e-08 1.7993998875959782 1.6261e-08 1.8358989909588432 1.6262e-08 1.7773178424698242 1.6262999999999998e-08 1.9365189246088135 1.6264e-08 1.8053123776909192 1.6265e-08 1.8939300212664434 1.6265999999999998e-08 1.879576910214256 1.6267e-08 1.7487407235792343 1.6268e-08 1.8657783318591186 1.6268999999999998e-08 1.75082005635354 1.627e-08 1.7922612248087126 1.6271e-08 1.6697183158432563 1.6272e-08 1.7680288298955908 1.6273e-08 1.7994414245268997 1.6274e-08 1.826779110250135 1.6275e-08 1.7930710398216507 1.6276e-08 1.8382946084383485 1.6277e-08 1.8376981188389656 1.6278e-08 1.7752437265133736 1.6279e-08 1.7008017767117862 1.628e-08 1.7559368433353888 1.6281e-08 1.7589812810087289 1.6282e-08 1.8305734493608938 1.6283e-08 1.806259250404378 1.6284e-08 1.8378736310375288 1.6285e-08 1.7850757870747909 1.6286e-08 1.8328169399474774 1.6287e-08 1.7661993430002987 1.6288e-08 1.8571573565057016 1.6289e-08 1.7090453247914275 1.629e-08 1.8186087311675632 1.6291e-08 1.7730831459619076 1.6292e-08 1.783258117788072 1.6293e-08 1.7897478751824265 1.6294e-08 1.780121041614124 1.6295e-08 1.7655611932703574 1.6296e-08 1.8483743493165334 1.6297e-08 1.8910053045597846 1.6297999999999998e-08 1.846901842623501 1.6299e-08 1.767361636168156 1.63e-08 1.8609662740639072 1.6300999999999998e-08 1.7829396405299704 1.6302e-08 1.8326069670169172 1.6303e-08 1.8820967109786875 1.6303999999999998e-08 1.878291185050804 1.6305e-08 1.8852294698533494 1.6306e-08 1.8819239793633615 1.6307e-08 1.79145676120259 1.6308e-08 1.8252113487239428 1.6309e-08 1.7548784057074804 1.631e-08 1.7825254089795406 1.6311e-08 1.8531344253693451 1.6312e-08 1.8879244365901307 1.6313e-08 1.7628195859165905 1.6314e-08 1.8131130111403426 1.6315e-08 1.7729244603417582 1.6316e-08 1.8067263227504302 1.6317e-08 1.7724223115405766 1.6318e-08 1.873871381579067 1.6319e-08 1.8177632782397546 1.632e-08 1.7969870233622394 1.6321e-08 1.8793388958155781 1.6322e-08 1.8103011529303599 1.6323e-08 1.8753519512455386 1.6324e-08 1.8053664337509465 1.6325e-08 1.7940547455635505 1.6326e-08 1.7995165579132597 1.6327e-08 1.9107513157529485 1.6328e-08 1.7277685593681795 1.6329e-08 1.7873350132810146 1.633e-08 1.7763095033028782 1.6331e-08 1.7995397256302854 1.6332e-08 1.7851078606205202 1.6332999999999998e-08 1.8619144373358654 1.6334e-08 1.811377003846565 1.6335e-08 1.6936229047446465 1.6335999999999998e-08 1.7572068671576637 1.6337e-08 1.8271902096695922 1.6338e-08 1.8423094326998941 1.6338999999999998e-08 1.8269241230764288 1.634e-08 1.8314916527846792 1.6341e-08 1.800866111671457 1.6342e-08 1.836232873861142 1.6343e-08 1.8085936052665066 1.6344e-08 1.753040837778039 1.6345e-08 1.8307639242490485 1.6346e-08 1.7668356435619312 1.6347e-08 1.8306744260017014 1.6348e-08 1.85637596405476 1.6349e-08 1.8204139924258749 1.635e-08 1.8343000354111147 1.6351e-08 1.8327445492779058 1.6352e-08 1.764939702349545 1.6353e-08 1.8528996790950505 1.6354e-08 1.7807646128933783 1.6355e-08 1.7422015160097268 1.6356e-08 1.9213601242560363 1.6357e-08 1.734517314016504 1.6358e-08 1.8371708680941332 1.6359e-08 1.747813900747437 1.636e-08 1.8034126844993101 1.6361e-08 1.82510640612657 1.6362e-08 1.8003354802863603 1.6363e-08 1.8947226005954554 1.6364e-08 1.7731196935957028 1.6365e-08 1.8564533629539972 1.6366e-08 1.750520485942339 1.6367e-08 1.9267900897810117 1.6367999999999998e-08 1.776836753446104 1.6369e-08 1.8185786806548745 1.637e-08 1.8085260879854206 1.6370999999999998e-08 1.763942236091316 1.6372e-08 1.8221094918665905 1.6373e-08 1.7767477665548128 1.6373999999999998e-08 1.8457776045214616 1.6375e-08 1.7533496433080553 1.6376e-08 1.7950038549823797 1.6377e-08 1.792184500859734 1.6378e-08 1.7368676660869788 1.6379e-08 1.8711407791005614 1.638e-08 1.8722689901680123 1.6381e-08 1.7499518061555666 1.6382e-08 1.6754965052192317 1.6383e-08 1.7781521483001674 1.6384e-08 1.803963802009045 1.6385e-08 1.8257879379519124 1.6386e-08 1.8100655798025962 1.6387e-08 1.7877650192852357 1.6388e-08 1.8557218643439657 1.6389e-08 1.7103972215956382 1.639e-08 1.8666482685482748 1.6391e-08 1.7828243700924944 1.6392e-08 1.8636699029187447 1.6393e-08 1.8453193059339885 1.6394e-08 1.7704197171888403 1.6395e-08 1.7262739412563062 1.6396e-08 1.839545589764204 1.6397e-08 1.8108736563427155 1.6398e-08 1.7431565616017795 1.6399e-08 1.8273728798538673 1.64e-08 1.833748827949972 1.6401e-08 1.828480939672344 1.6402e-08 1.7845107433599137 1.6402999999999998e-08 1.8338072583717862 1.6404e-08 1.8498271872100926 1.6405e-08 1.8603940190873072 1.6405999999999998e-08 1.8415204609410423 1.6407e-08 1.7450765266344805 1.6408e-08 1.753100765320981 1.6408999999999998e-08 1.7946959765245651 1.641e-08 1.798833113973758 1.6411e-08 1.8165787797537278 1.6411999999999998e-08 1.8408252181827696 1.6413e-08 1.8036373876105167 1.6414e-08 1.8196916271523413 1.6415e-08 1.7522291697474022 1.6416e-08 1.873792946185179 1.6417e-08 1.7575804331111802 1.6418e-08 1.8709490189093185 1.6419e-08 1.8420402162593976 1.642e-08 1.8990238563013822 1.6421e-08 1.8216626750662184 1.6422e-08 1.8930890897935968 1.6423e-08 1.7791644008792904 1.6424e-08 1.7731146421926123 1.6425e-08 1.7613225626769422 1.6426e-08 1.9186574478815948 1.6427e-08 1.7715262823153968 1.6428e-08 1.7349595379516431 1.6429e-08 1.7626153252578072 1.643e-08 1.7819874303564152 1.6431e-08 1.8048571308844836 1.6432e-08 1.8578704581009984 1.6433e-08 1.7143658590302686 1.6434e-08 1.7629556945773401 1.6435e-08 1.7467523791972144 1.6436e-08 1.9318440181921048 1.6437e-08 1.7395607395190091 1.6437999999999998e-08 1.7955146735757774 1.6439e-08 1.7415051192207942 1.644e-08 1.7510441363061975 1.6440999999999998e-08 1.7702905575866548 1.6442e-08 1.7173900888664735 1.6443e-08 1.848714642411792 1.6443999999999998e-08 1.8216534579385195 1.6445e-08 1.8846495880326968 1.6446e-08 1.814527432997777 1.6446999999999998e-08 1.8045608665993864 1.6448e-08 1.703100500760355 1.6449e-08 1.8740366049261588 1.645e-08 1.7545879699394182 1.6451e-08 1.8363899074230108 1.6452e-08 1.8177231820879627 1.6453e-08 1.7437396914819747 1.6454e-08 1.7657650650492185 1.6455e-08 1.850960059171928 1.6456e-08 1.6799061963800908 1.6457e-08 1.6559821965903783 1.6458e-08 1.776556389117613 1.6459e-08 1.771865508004812 1.646e-08 1.8220100779337458 1.6461e-08 1.811488471161559 1.6462e-08 1.7738178895863603 1.6463e-08 1.7361503594213203 1.6464e-08 1.7683798989608566 1.6465e-08 1.762934412528348 1.6466e-08 1.7753689577276748 1.6467e-08 1.7431127201655185 1.6468e-08 1.7855330822783315 1.6469e-08 1.8338731188669977 1.647e-08 1.8660116338597652 1.6471e-08 1.8383747202031557 1.6472e-08 1.7991387933862777 1.6472999999999998e-08 1.7295852828712217 1.6474e-08 1.7984592254066902 1.6475e-08 1.9367023072781149 1.6475999999999998e-08 1.8150419976848453 1.6477e-08 1.8184116776834545 1.6478e-08 1.8819431776044153 1.6478999999999998e-08 1.7743568138268855 1.648e-08 1.784215530579821 1.6481e-08 1.8276349107559895 1.6481999999999998e-08 1.7071863823279498 1.6483e-08 1.7890409048664704 1.6484e-08 1.845790210688156 1.6485e-08 1.858766501063185 1.6486e-08 1.8355929739352717 1.6487e-08 1.8318029539066922 1.6488e-08 1.7540939617353841 1.6489e-08 1.8195134099551458 1.649e-08 1.681558108082986 1.6491e-08 1.7875019177115448 1.6492e-08 1.7617499054257781 1.6493e-08 1.8297462810428626 1.6494e-08 1.7980080203018736 1.6495e-08 1.8349914912645824 1.6496e-08 1.7575197462367496 1.6497e-08 1.7713641970530334 1.6498e-08 1.8291778875019613 1.6499e-08 1.9149476918190154 1.65e-08 1.7503572033165464 1.6501e-08 1.8266555916733174 1.6502e-08 1.889512646229683 1.6503e-08 1.7284862673600543 1.6504e-08 1.794745260892121 1.6505e-08 1.739461196198028 1.6506e-08 1.7298193580093622 1.6507e-08 1.719272743570918 1.6508e-08 1.7894507897590242 1.6509e-08 1.7998427227856608 1.651e-08 1.8644720331131475 1.6510999999999998e-08 1.9366454799731432 1.6512e-08 1.773846507193764 1.6513e-08 1.801975883429188 1.6513999999999998e-08 1.8404183621669692 1.6515e-08 1.734029498867513 1.6516e-08 1.8681334407091001 1.6516999999999998e-08 1.8175635966548096 1.6518e-08 1.7892042552088998 1.6519e-08 1.8466308097033466 1.652e-08 1.7819813900276484 1.6521e-08 1.77901235926244 1.6522e-08 1.7962951361033264 1.6523e-08 1.7983913823960767 1.6524e-08 1.7737129378042595 1.6525e-08 1.7725410222588143 1.6526e-08 1.8566566096264165 1.6527e-08 1.822269543782713 1.6528e-08 1.7092206510139862 1.6529e-08 1.8593371498714868 1.653e-08 1.7220159054051898 1.6531e-08 1.8063431551835394 1.6532e-08 1.7170154831648043 1.6533e-08 1.8869722190426086 1.6534e-08 1.7925000397508697 1.6535e-08 1.8249973188632596 1.6536e-08 1.7383231144293736 1.6537e-08 1.7556992695860967 1.6538e-08 1.8287784468958674 1.6539e-08 1.7975886614384953 1.654e-08 1.853634370203812 1.6541e-08 1.7533763405800793 1.6542e-08 1.813215957712728 1.6543e-08 1.7396731743471985 1.6544e-08 1.8225697788331363 1.6545e-08 1.72317501351762 1.6545999999999998e-08 1.7839531297642894 1.6547e-08 1.8376269423080127 1.6548e-08 1.7328690645294846 1.6548999999999998e-08 1.8505194586308484 1.655e-08 1.7555999264727111 1.6551e-08 1.8685323058149144 1.6551999999999998e-08 1.811834229637517 1.6553e-08 1.7925112116566162 1.6554e-08 1.8517246649961012 1.6555e-08 1.871321634016711 1.6556e-08 1.8689273339227541 1.6557e-08 1.8340525793696933 1.6558e-08 1.8340822695902712 1.6559e-08 1.8286114004289564 1.656e-08 1.8551455669329115 1.6561e-08 1.83287994330361 1.6562e-08 1.7804749779196287 1.6563e-08 1.858578979416234 1.6564e-08 1.7196510846575948 1.6565e-08 1.7826452142199192 1.6566e-08 1.8240143893709129 1.6567e-08 1.7542110267044442 1.6568e-08 1.8433380297927375 1.6569e-08 1.7964430909407345 1.657e-08 1.7612864106985795 1.6571e-08 1.7363709087038561 1.6572e-08 1.8324930318778132 1.6573e-08 1.920973906406611 1.6574e-08 1.7183531236383816 1.6575e-08 1.7750047763696282 1.6576e-08 1.7700747053402357 1.6577e-08 1.7195635376172167 1.6578e-08 1.7926741201217753 1.6579e-08 1.7947335514257794 1.658e-08 1.875171436076339 1.6580999999999998e-08 1.6992391879551305 1.6582e-08 1.7718749715103463 1.6583e-08 1.865546488285828 1.6583999999999998e-08 1.8186139506238477 1.6585e-08 1.6902404020997592 1.6586e-08 1.8047123355866457 1.6586999999999998e-08 1.8518212459942642 1.6588e-08 1.8233473667870859 1.6589e-08 1.8085163350651425 1.6589999999999998e-08 1.8017991020274526 1.6591e-08 1.790175923692966 1.6592e-08 1.7989446632854218 1.6593e-08 1.7777628835971866 1.6594e-08 1.7394621087565985 1.6595e-08 1.751113938614572 1.6596e-08 1.832798393781668 1.6597e-08 1.7861397503194598 1.6598e-08 1.7872952371462703 1.6599e-08 1.8182018526822878 1.66e-08 1.9397809918115398 1.6601e-08 1.8132606416289 1.6602e-08 1.8487001656640856 1.6603e-08 1.767305920911129 1.6604e-08 1.830630553505871 1.6605e-08 1.7808900093219893 1.6606e-08 1.7399163596814782 1.6607e-08 1.7790085365382546 1.6608e-08 1.7321843744538001 1.6609e-08 1.8622824946579803 1.661e-08 1.762228994368235 1.6611e-08 1.6793704406218308 1.6612e-08 1.8846509577638806 1.6613e-08 1.8125037910198953 1.6614e-08 1.720275749220965 1.6615e-08 1.8337117066593924 1.6615999999999998e-08 1.7389444195994521 1.6617e-08 1.7876483617226921 1.6618e-08 1.8373823248809604 1.6618999999999998e-08 1.854172572845882 1.662e-08 1.7338652989334948 1.6621e-08 1.799220634349488 1.6621999999999998e-08 1.768103878031287 1.6623e-08 1.85783635389081 1.6624e-08 1.8647683939850181 1.6624999999999998e-08 1.79204177142447 1.6626e-08 1.8533575124387727 1.6627e-08 1.8112529106507298 1.6628e-08 1.900913628957578 1.6629e-08 1.8008275115407328 1.663e-08 1.7638663492693372 1.6631e-08 1.7637820526513797 1.6632e-08 1.8201278573450208 1.6633e-08 1.7838477708923492 1.6634e-08 1.8667903536624983 1.6635e-08 1.7617127243443127 1.6636e-08 1.8299376153890698 1.6637e-08 1.8700826784190627 1.6638e-08 1.7548420538596945 1.6639e-08 1.8021332537222396 1.664e-08 1.7602023987880628 1.6641e-08 1.7891122504309982 1.6642e-08 1.7542919023285704 1.6643e-08 1.885981672619878 1.6644e-08 1.75988486438015 1.6645e-08 1.9111766810671713 1.6646e-08 1.8275007112023056 1.6647e-08 1.739237994440798 1.6648e-08 1.828369731212734 1.6649e-08 1.723591142960736 1.665e-08 1.7985898500511381 1.6650999999999998e-08 1.7305307732610977 1.6652e-08 1.8592529720498605 1.6653e-08 1.8069616475188193 1.6653999999999998e-08 1.7594693678805278 1.6655e-08 1.8163381558021463 1.6656e-08 1.752886585877717 1.6656999999999998e-08 1.8596890370421881 1.6658e-08 1.7317570670864666 1.6659e-08 1.7902867093682735 1.6659999999999998e-08 1.889350221909011 1.6661e-08 1.816353400700724 1.6662e-08 1.8506860512872303 1.6663e-08 1.8084679066416502 1.6664e-08 1.7727665439106997 1.6665e-08 1.6849565860631597 1.6666e-08 1.8518761271556925 1.6667e-08 1.6988179922050741 1.6668e-08 1.7881246938950635 1.6669e-08 1.793999275813594 1.667e-08 1.762643270473583 1.6671e-08 1.8073115528262913 1.6672e-08 1.8602644990495008 1.6673e-08 1.709861397041728 1.6674e-08 1.8058675234392112 1.6675e-08 1.8575831134481975 1.6676e-08 1.8911826034702066 1.6677e-08 1.9024224387434459 1.6678e-08 1.7791859094109532 1.6679e-08 1.8671564510112548 1.668e-08 1.7799039182028755 1.6681e-08 1.8141922698010888 1.6682e-08 1.7366368384882676 1.6683e-08 1.7852212579319604 1.6684e-08 1.75841817806096 1.6685e-08 1.8219214346654522 1.6686e-08 1.8071242627305322 1.6687e-08 1.871522752625562 1.6688e-08 1.8274466762765884 1.6688999999999998e-08 1.8745088805420331 1.669e-08 1.71131262856634 1.6691e-08 1.7819954926656418 1.6691999999999998e-08 1.7592983195420815 1.6693e-08 1.8391889880769892 1.6694e-08 1.8668312772203584 1.6694999999999998e-08 1.7597740910746336 1.6696e-08 1.8138428652401857 1.6697e-08 1.7907286998758747 1.6698e-08 1.7441503159155038 1.6699e-08 1.9129438150823082 1.67e-08 1.8113645747582414 1.6701e-08 1.8894720582412614 1.6702e-08 1.8525033755572153 1.6703e-08 1.813109783477063 1.6704e-08 1.753552740912961 1.6705e-08 1.9262079443838804 1.6706e-08 1.7423168758752345 1.6707e-08 1.9009183825947924 1.6708e-08 1.8489856720998519 1.6709e-08 1.7392643697949226 1.671e-08 1.76228588068627 1.6711e-08 1.7461092518338186 1.6712e-08 1.7791396754875115 1.6713e-08 1.8951879101660576 1.6714e-08 1.7867987905812306 1.6715e-08 1.8497228579858893 1.6716e-08 1.732864065412298 1.6717e-08 1.8148179070527812 1.6718e-08 1.76141813032227 1.6719e-08 1.768760895827384 1.672e-08 1.8809990933801732 1.6721e-08 1.78553656987805 1.6722e-08 1.758004274216781 1.6723e-08 1.8110797204949625 1.6723999999999998e-08 1.8208747363999174 1.6725e-08 1.7960701119286184 1.6726e-08 1.8631856042799468 1.6726999999999998e-08 1.8024313665036755 1.6728e-08 1.7908191672751408 1.6729e-08 1.7269663655257625 1.6729999999999998e-08 1.7372404797057996 1.6731e-08 1.791921837304388 1.6732e-08 1.770045837472244 1.6733e-08 1.7777433781597773 1.6734e-08 1.8449084607221191 1.6735e-08 1.8303210456615127 1.6736e-08 1.8470526327563128 1.6737e-08 1.819549712341562 1.6738e-08 1.8581218839616211 1.6739e-08 1.810095116386717 1.674e-08 1.7222246041275038 1.6741e-08 1.8499841249756024 1.6742e-08 1.8141315868592562 1.6743e-08 1.8350658206417685 1.6744e-08 1.8074595738192865 1.6745e-08 1.7737310934116204 1.6746e-08 1.7250112988228747 1.6747e-08 1.804334304767481 1.6748e-08 1.7678481479189472 1.6749e-08 1.8615341376959587 1.675e-08 1.8514713148024768 1.6751e-08 1.810127252184624 1.6752e-08 1.8172309281625783 1.6753e-08 1.7883982458944538 1.6754e-08 1.852886793393276 1.6755e-08 1.7572329028173568 1.6756e-08 1.8177262516375725 1.6757e-08 1.8108063497725466 1.6758e-08 1.7472931244497054 1.6758999999999998e-08 1.8456766965230214 1.676e-08 1.8583114212161065 1.6761e-08 1.769588010157777 1.6761999999999998e-08 1.780297337800512 1.6763e-08 1.7634033730201668 1.6764e-08 1.8574540910113435 1.6764999999999998e-08 1.7941176304279605 1.6766e-08 1.7771605818560117 1.6767e-08 1.751208034642832 1.6767999999999998e-08 1.8547814548142205 1.6769e-08 1.7715701531737529 1.677e-08 1.7315774558281212 1.6771e-08 1.8792587127987594 1.6772e-08 1.7937762392753762 1.6773e-08 1.8844605457504942 1.6774e-08 1.8594844103034236 1.6775e-08 1.8298927800672498 1.6776e-08 1.7786557907241096 1.6777e-08 1.79123855289472 1.6778e-08 1.7698338053008804 1.6779e-08 1.826398118222432 1.678e-08 1.859576882266555 1.6781e-08 1.880494779916838 1.6782e-08 1.6599546453361644 1.6783e-08 1.785208885760444 1.6784e-08 1.8236225053596313 1.6785e-08 1.752388732053827 1.6786e-08 1.855143293074444 1.6787e-08 1.8275664585301008 1.6788e-08 1.8073818873506207 1.6789e-08 1.7906287482071945 1.679e-08 1.7937894294844206 1.6791e-08 1.7747488988600673 1.6792e-08 1.696505052419731 1.6793e-08 1.798121857427347 1.6793999999999998e-08 1.7622002370110532 1.6795e-08 1.8127414437053955 1.6796e-08 1.8408692636810564 1.6796999999999998e-08 1.813660638739446 1.6798e-08 1.8072465835815374 1.6799e-08 1.7234204062361522 1.6799999999999998e-08 1.858090347869871 1.6801e-08 1.8036937525241983 1.6802e-08 1.8810776878075965 1.6802999999999998e-08 1.7737224906301308 1.6804e-08 1.7776725932645059 1.6805e-08 1.7703726238193234 1.6806e-08 1.77881506802829 1.6807e-08 1.807303125784137 1.6808e-08 1.7646077419207578 1.6809e-08 1.7821387625367862 1.681e-08 1.7234482130126125 1.6811e-08 1.7708317377531733 1.6812e-08 1.7631901270046288 1.6813e-08 1.8176631776989314 1.6814e-08 1.912309525083987 1.6815e-08 1.7882200205452694 1.6816e-08 1.7647628722413171 1.6817e-08 1.8613303697167614 1.6818e-08 1.7580115037735264 1.6819e-08 1.8267767239692252 1.682e-08 1.834377970464133 1.6821e-08 1.8211066326533225 1.6822e-08 1.7613893252058501 1.6823e-08 1.801459400283757 1.6824e-08 1.8567825071498594 1.6825e-08 1.8087841293156086 1.6826e-08 1.7696256250750524 1.6827e-08 1.8005003335511207 1.6828e-08 1.7761765582285836 1.6828999999999998e-08 1.7147430375938393 1.683e-08 1.844365367484641 1.6831e-08 1.8087224865352907 1.6831999999999998e-08 1.6943428282232156 1.6833e-08 1.8310961442903801 1.6834e-08 1.7562414265415478 1.6834999999999998e-08 1.7850130779869644 1.6836e-08 1.7204542268002574 1.6837e-08 1.8215648191357352 1.6837999999999998e-08 1.8517138358456287 1.6839e-08 1.7746034077922885 1.684e-08 1.8504413709660743 1.6841e-08 1.7906380967651017 1.6842e-08 1.8140645923188974 1.6843e-08 1.8269292905357484 1.6844e-08 1.8400653685558659 1.6845e-08 1.7498777952633675 1.6846e-08 1.7590781469044785 1.6847e-08 1.7315574637202078 1.6848e-08 1.7992568295773075 1.6849e-08 1.8189571436178968 1.685e-08 1.7485997265282305 1.6851e-08 1.7067270493856563 1.6852e-08 1.7489362510579947 1.6853e-08 1.7349165613097086 1.6854e-08 1.8779810816351252 1.6855e-08 1.8005136768423704 1.6856e-08 1.744944271629761 1.6857e-08 1.803626205699184 1.6858e-08 1.7947443290580427 1.6859e-08 1.7886337473568854 1.686e-08 1.8253562145398103 1.6861e-08 1.7739980909142417 1.6862e-08 1.8457434805887343 1.6863e-08 1.7963159706932599 1.6863999999999998e-08 1.8007814207046533 1.6865e-08 1.850594757914959 1.6866e-08 1.8090938516773098 1.6866999999999998e-08 1.810125526745791 1.6868e-08 1.8369969737906704 1.6869e-08 1.7409897471113065 1.6869999999999998e-08 1.7681791399768656 1.6871e-08 1.8128085392887268 1.6872e-08 1.7484470556622256 1.6872999999999998e-08 1.804989836377042 1.6874e-08 1.7176799796601614 1.6875e-08 1.7679824841921676 1.6876e-08 1.7490660484361982 1.6877e-08 1.7255541570261455 1.6878e-08 1.8208188921569977 1.6879e-08 1.7887611408188429 1.688e-08 1.7137866463065383 1.6881e-08 1.8247676101145474 1.6882e-08 1.8284821390231178 1.6883e-08 1.8058520202302593 1.6884e-08 1.8597477053674654 1.6885e-08 1.8296539165641201 1.6886e-08 1.7857013779248772 1.6887e-08 1.855242135926928 1.6888e-08 1.7551272821855906 1.6889e-08 1.898613103296125 1.689e-08 1.8417686581174646 1.6891e-08 1.78798516352025 1.6892e-08 1.8271974856394435 1.6893e-08 1.8558665485944859 1.6894e-08 1.8467037935487778 1.6895e-08 1.7009425443375794 1.6896e-08 1.8242925136307386 1.6897e-08 1.9677694637884804 1.6898e-08 1.8324263093049755 1.6899e-08 1.857261351557108 1.69e-08 1.8335519718911482 1.6901e-08 1.7279039269357201 1.6901999999999998e-08 1.768311127630627 1.6903e-08 1.7308225567176727 1.6904e-08 1.8348043829023002 1.6904999999999998e-08 1.684207131719202 1.6906e-08 1.8546556923925654 1.6907e-08 1.710295119257802 1.6907999999999998e-08 1.7356102230315795 1.6909e-08 1.819684096379164 1.691e-08 1.8274341932913465 1.6911e-08 1.8503161503411196 1.6912e-08 1.8227112996286823 1.6913e-08 1.7977291325052251 1.6914e-08 1.7608546735811244 1.6915e-08 1.7495812443175043 1.6916e-08 1.8698945392507857 1.6917e-08 1.8529268189157726 1.6918e-08 1.7500058823810711 1.6919e-08 1.8570767089264737 1.692e-08 1.8338182379722625 1.6921e-08 1.9118765811312481 1.6922e-08 1.847434661245632 1.6923e-08 1.751268746069587 1.6924e-08 1.7708949505840916 1.6925e-08 1.8250180167382992 1.6926e-08 1.7630234747821651 1.6927e-08 1.808960481920575 1.6928e-08 1.7059807102757782 1.6929e-08 1.88631063941239 1.693e-08 1.8395878124376366 1.6931e-08 1.8034542110919278 1.6932e-08 1.842337571170882 1.6933e-08 1.8298220569561672 1.6934e-08 1.7788764799697234 1.6935e-08 1.8210330730676596 1.6936e-08 1.8312435243898337 1.6936999999999998e-08 1.8450077048631377 1.6938e-08 1.7930888294651373 1.6939e-08 1.8318914843188692 1.6939999999999998e-08 1.790485617432935 1.6941e-08 1.7848466437485642 1.6942e-08 1.8727667635602585 1.6942999999999998e-08 1.7950337929888454 1.6944e-08 1.8203834014797748 1.6945e-08 1.7795917558917966 1.6946e-08 1.8499178036151291 1.6947e-08 1.8193772090307103 1.6948e-08 1.765429696448563 1.6949e-08 1.7520849184947243 1.695e-08 1.8554102753001829 1.6951e-08 1.7760944694861391 1.6952e-08 1.739966636844885 1.6953e-08 1.9057737899250067 1.6954e-08 1.8148455805510864 1.6955e-08 1.807960302460672 1.6956e-08 1.8191216343544871 1.6957e-08 1.7741951646602279 1.6958e-08 1.77632355250461 1.6959e-08 1.674427140662397 1.696e-08 1.8328576676357748 1.6961e-08 1.8164157406146613 1.6962e-08 1.8798406987256189 1.6963e-08 1.8344603352706763 1.6964e-08 1.8225468610944036 1.6965e-08 1.7470745830407763 1.6966e-08 1.7881783747387208 1.6967e-08 1.8428924737690409 1.6968e-08 1.7842152682396653 1.6969e-08 1.79027014236457 1.697e-08 1.9083315054438066 1.6971e-08 1.7529659603161207 1.6971999999999998e-08 1.798034232238146 1.6973e-08 1.6886098714794473 1.6974e-08 1.727735009264524 1.6974999999999998e-08 1.7754050736369034 1.6976e-08 1.8202602103786283 1.6977e-08 1.7814992907161065 1.6977999999999998e-08 1.7074932860787801 1.6979e-08 1.7780538338959193 1.698e-08 1.7991245611326152 1.6980999999999998e-08 1.7861801042653858 1.6982e-08 1.7682937230157159 1.6983e-08 1.765306038576383 1.6984e-08 1.7664411337294845 1.6985e-08 1.7267822045255812 1.6986e-08 1.8305607409985831 1.6987e-08 1.8269033237635786 1.6988e-08 1.7875726721376737 1.6989e-08 1.7948221432021016 1.699e-08 1.6867801610146298 1.6991e-08 1.7612008750478092 1.6992e-08 1.911533950165796 1.6993e-08 1.745117196478785 1.6994e-08 1.797480717164933 1.6995e-08 1.807503637382111 1.6996e-08 1.8115508656492785 1.6997e-08 1.7934581034688806 1.6998e-08 1.8011251900247576 1.6999e-08 1.720110338027296 1.7e-08 1.885209852029092 1.7001e-08 1.8979338649375235 1.7002e-08 1.8339081893541573 1.7003e-08 1.7401099538309204 1.7004e-08 1.8187755460342137 1.7005e-08 1.7241030011231744 1.7006e-08 1.8484534871348257 1.7006999999999998e-08 1.7943418346075162 1.7008e-08 1.7978451763920877 1.7009e-08 1.7713758753353224 1.7009999999999998e-08 1.7952230305061962 1.7011e-08 1.75666923364623 1.7012e-08 1.8320931016524673 1.7012999999999998e-08 1.8527610658118665 1.7014e-08 1.8659230811515988 1.7015e-08 1.772502395141822 1.7015999999999998e-08 1.8404523115809053 1.7017e-08 1.7319231094028025 1.7018e-08 1.8344942060384237 1.7019e-08 1.712127119881281 1.702e-08 1.7647869988379656 1.7021e-08 1.7410684356750692 1.7022e-08 1.7725927230520575 1.7023e-08 1.8285218497655722 1.7024e-08 1.760109654839131 1.7025e-08 1.7666693867392573 1.7026e-08 1.792383799539885 1.7027e-08 1.7946538722280065 1.7028e-08 1.7919409083278168 1.7029e-08 1.7636053832165801 1.703e-08 1.7340197070699361 1.7031e-08 1.7135693686700024 1.7032e-08 1.7265393494148282 1.7033e-08 1.767408665001718 1.7034e-08 1.7763674803629455 1.7035e-08 1.8132301543168585 1.7036e-08 1.8135804603987897 1.7037e-08 1.903452255136561 1.7038e-08 1.7914211690956006 1.7039e-08 1.7761634986053485 1.704e-08 1.8507439240045245 1.7041e-08 1.8699977788257343 1.7041999999999998e-08 1.7614356892185425 1.7043e-08 1.8336666520579903 1.7044e-08 1.8047177470796272 1.7044999999999998e-08 1.820902120142135 1.7046e-08 1.748898176831902 1.7047e-08 1.8380825987660023 1.7047999999999998e-08 1.7698182140170329 1.7049e-08 1.8717261713370372 1.705e-08 1.822046231941503 1.7050999999999998e-08 1.83081084735185 1.7052e-08 1.846090963103442 1.7053e-08 1.7409113572516595 1.7054e-08 1.719677499553527 1.7055e-08 1.7626250308312186 1.7056e-08 1.841423264559105 1.7057e-08 1.8475917508926527 1.7058e-08 1.7869264294016614 1.7059e-08 1.8267131186266452 1.706e-08 1.8218506898852325 1.7061e-08 1.8820591024149997 1.7062e-08 1.8280182413950459 1.7063e-08 1.7410640323690911 1.7064e-08 1.8310036893942798 1.7065e-08 1.876607936022216 1.7066e-08 1.8605947110868224 1.7067e-08 1.7751944836586615 1.7068e-08 1.733792022079672 1.7069e-08 1.821554013026114 1.707e-08 1.7538908080179363 1.7071e-08 1.7764494544783689 1.7072e-08 1.77188592566527 1.7073e-08 1.7091705629104115 1.7074e-08 1.7832541823481354 1.7075e-08 1.8228236641632687 1.7076e-08 1.7803933703382764 1.7077e-08 1.8275305706897398 1.7078e-08 1.8976130148719272 1.7079e-08 1.837782916655443 1.7079999999999998e-08 1.7474346769810363 1.7081e-08 1.8113426550581748 1.7082e-08 1.7543520635946293 1.7082999999999998e-08 1.7158390234473075 1.7084e-08 1.7956201710462527 1.7085e-08 1.8382909606888245 1.7085999999999998e-08 1.7604492842432435 1.7087e-08 1.7780343238751422 1.7088e-08 1.7780712955414537 1.7089e-08 1.8098232697167134 1.709e-08 1.775569463412821 1.7091e-08 1.8437591457760227 1.7092e-08 1.855824277440567 1.7093e-08 1.7771083645285104 1.7094e-08 1.7582261333731029 1.7095e-08 1.8129938269602595 1.7096e-08 1.766984567905938 1.7097e-08 1.8191320718933863 1.7098e-08 1.827208784342086 1.7099e-08 1.815834456311778 1.71e-08 1.7550842532469095 1.7101e-08 1.835794114011574 1.7102e-08 1.7557177079882473 1.7103e-08 1.730789056830494 1.7104e-08 1.8164373100224507 1.7105e-08 1.7910921982449235 1.7106e-08 1.8433715380431874 1.7107e-08 1.8403133732019545 1.7108e-08 1.833510463563012 1.7109e-08 1.7205724455889482 1.711e-08 1.8323854207032175 1.7111e-08 1.860587453856629 1.7112e-08 1.8528547430659335 1.7113e-08 1.8646670712944446 1.7114e-08 1.8137240378269597 1.7114999999999998e-08 1.869971340692762 1.7116e-08 1.8842733782737187 1.7117e-08 1.8489272137740993 1.7117999999999998e-08 1.7811160017520369 1.7119e-08 1.8151291922203474 1.712e-08 1.8499281807858992 1.7120999999999998e-08 1.8181508424656998 1.7122e-08 1.7685532984422365 1.7123e-08 1.7848835023172454 1.7124e-08 1.7599889730809632 1.7125e-08 1.7829703864631028 1.7126e-08 1.825210482810954 1.7127e-08 1.819003112302546 1.7128e-08 1.8858523573610615 1.7129e-08 1.8142299317107404 1.713e-08 1.7501194728597742 1.7131e-08 1.8135494763587956 1.7132e-08 1.729044153120708 1.7133e-08 1.877580049015539 1.7134e-08 1.7693053310783369 1.7135e-08 1.669968373006533 1.7136e-08 1.8419452208277856 1.7137e-08 1.8073848795095728 1.7138e-08 1.8076738050570071 1.7139e-08 1.7629911644069534 1.714e-08 1.8209189179180083 1.7141e-08 1.81450268539778 1.7142e-08 1.7442742839699783 1.7143e-08 1.7600777082144305 1.7144e-08 1.8301117161326803 1.7145e-08 1.8186101542966377 1.7146e-08 1.8930466545662585 1.7147e-08 1.805058591607381 1.7148e-08 1.8389785765116884 1.7149e-08 1.8105721143042324 1.7149999999999998e-08 1.9416061732340344 1.7151e-08 1.7871366253358978 1.7152e-08 1.7783577026064985 1.7152999999999998e-08 1.781821963041132 1.7154e-08 1.831116837815528 1.7155e-08 1.7874417028620535 1.7155999999999998e-08 1.78274817860886 1.7157e-08 1.7750616903514331 1.7158e-08 1.7550933402459135 1.7158999999999998e-08 1.8260252385208393 1.716e-08 1.8645927103308788 1.7161e-08 1.9117954536317319 1.7162e-08 1.6993452393627306 1.7163e-08 1.7714936542653246 1.7164e-08 1.9144859353176442 1.7165e-08 1.7774938582940616 1.7166e-08 1.8212726473093765 1.7167e-08 1.8773165848951254 1.7168e-08 1.7960756345005584 1.7169e-08 1.81780673054013 1.717e-08 1.7736260572768625 1.7171e-08 1.7500543173841787 1.7172e-08 1.7910936832377216 1.7173e-08 1.845891671237222 1.7174e-08 1.9597401626650681 1.7175e-08 1.8479625448948669 1.7176e-08 1.7807244448255648 1.7177e-08 1.7379121826610837 1.7178e-08 1.7290424463901184 1.7179e-08 1.8486031777186553 1.718e-08 1.8449702257072584 1.7181e-08 1.7646183605574481 1.7182e-08 1.8072763110372327 1.7183e-08 1.7041888615088074 1.7184e-08 1.7997983938109694 1.7184999999999998e-08 1.7752001433389295 1.7186e-08 1.780812969839374 1.7187e-08 1.6621201447425273 1.7187999999999998e-08 1.8063854858199178 1.7189e-08 1.762661526241135 1.719e-08 1.7716593700420682 1.7190999999999998e-08 1.8182342039420167 1.7192e-08 1.85611158925796 1.7193e-08 1.9027113246983633 1.7193999999999998e-08 1.8418891124882064 1.7195e-08 1.7241114587064315 1.7196e-08 1.8005057659663446 1.7197e-08 1.8361193388860273 1.7198e-08 1.7681154497353722 1.7199e-08 1.8634437838609288 1.72e-08 1.7513418797193634 1.7201e-08 1.8398572082175195 1.7202e-08 1.7727238928611038 1.7203e-08 1.82297252617921 1.7204e-08 1.7530442300955413 1.7205e-08 1.7755354503062237 1.7206e-08 1.7811834519043965 1.7207e-08 1.7878806246641104 1.7208e-08 1.7713772859565964 1.7209e-08 1.6963453777266408 1.721e-08 1.742611236367793 1.7211e-08 1.7489962543412456 1.7212e-08 1.7679689824603573 1.7213e-08 1.8035587352406728 1.7214e-08 1.9188421587126998 1.7215e-08 1.8330911626482866 1.7216e-08 1.8002472617577885 1.7217e-08 1.7956915714427677 1.7218e-08 1.7146185260305955 1.7219e-08 1.7988136780867212 1.7219999999999998e-08 1.834574252968787 1.7221e-08 1.8914162717022946 1.7222e-08 1.832606701293352 1.7222999999999998e-08 1.7698852771295022 1.7224e-08 1.7263023868301983 1.7225e-08 1.7109327603926832 1.7225999999999998e-08 1.7766785091995674 1.7227e-08 1.813843593695291 1.7228e-08 1.7809745429648538 1.7228999999999998e-08 1.8493043551887713 1.723e-08 1.8531584372534697 1.7231e-08 1.7984159023575075 1.7232e-08 1.7805152589927136 1.7233e-08 1.8335057205182668 1.7234e-08 1.810192981432577 1.7235e-08 1.7910458297451466 1.7236e-08 1.7457922193488278 1.7237e-08 1.7362431846207045 1.7238e-08 1.7280584310531577 1.7239e-08 1.7483498487977496 1.724e-08 1.7149122168012145 1.7241e-08 1.7348750305604925 1.7242e-08 1.8662404951266816 1.7243e-08 1.7718458404869295 1.7244e-08 1.7978864654534126 1.7245e-08 1.7724267300276024 1.7246e-08 1.8096902889005344 1.7247e-08 1.8300606446558336 1.7248e-08 1.7960627047067632 1.7249e-08 1.8141755630546728 1.725e-08 1.8007229064624066 1.7251e-08 1.8199255202981768 1.7252e-08 1.8840445456417096 1.7253e-08 1.8566238991210642 1.7254e-08 1.8218223352823826 1.7254999999999998e-08 1.8516023545167961 1.7256e-08 1.873896359043834 1.7257e-08 1.8369123774135503 1.7257999999999998e-08 1.8220076584178668 1.7259e-08 1.8278047826112729 1.726e-08 1.7799906870840343 1.7260999999999998e-08 1.8033790567701922 1.7262e-08 1.7269983106148443 1.7263e-08 1.8180216076116786 1.7263999999999998e-08 1.7842656321378874 1.7265e-08 1.7807511756025847 1.7266e-08 1.7903815740477091 1.7267e-08 1.7298924453759583 1.7268e-08 1.6457671776110636 1.7269e-08 1.8445906886716437 1.727e-08 1.8196103689528806 1.7271e-08 1.8179182589038436 1.7272e-08 1.8928882288712858 1.7273e-08 1.7647117504326353 1.7274e-08 1.7412720964190176 1.7275e-08 1.7443476292681996 1.7276e-08 1.7765186438473057 1.7277e-08 1.883541508745354 1.7278e-08 1.7783104304623043 1.7279e-08 1.830115479896351 1.728e-08 1.8727402462787799 1.7281e-08 1.9032869847704137 1.7282e-08 1.912130596035339 1.7283e-08 1.7520345138052456 1.7284e-08 1.767269977142156 1.7285e-08 1.8540128896464403 1.7286e-08 1.8207618821469813 1.7287e-08 1.8501733532498892 1.7288e-08 1.742211085980903 1.7289e-08 1.8082692322556078 1.729e-08 1.781262798250577 1.7291e-08 1.7703279747000713 1.7292e-08 1.8016598481858295 1.7292999999999998e-08 1.7707360727806938 1.7294e-08 1.737032021939783 1.7295e-08 1.8876902113594305 1.7295999999999998e-08 1.7993548517578588 1.7297e-08 1.8066742035216956 1.7298e-08 1.8081904039156662 1.7298999999999998e-08 1.837409949330668 1.73e-08 1.8154213268871138 1.7301e-08 1.763693092282452 1.7302e-08 1.7664399642605866 1.7303e-08 1.7723450756664438 1.7304e-08 1.874648112075514 1.7305e-08 1.7855068644231922 1.7306e-08 1.7079515682375062 1.7307e-08 1.861917416716754 1.7308e-08 1.7943528802431008 1.7309e-08 1.7451086960891269 1.731e-08 1.8405457396522271 1.7311e-08 1.8246676342116412 1.7312e-08 1.8089649569150654 1.7313e-08 1.798216671064133 1.7314e-08 1.791663919646533 1.7315e-08 1.8440005426303967 1.7316e-08 1.7896929503052368 1.7317e-08 1.787749625635998 1.7318e-08 1.8132005959772128 1.7319e-08 1.798897265095952 1.732e-08 1.7564802153364985 1.7321e-08 1.776920818642165 1.7322e-08 1.8563962200824053 1.7323e-08 1.8532865306436224 1.7324e-08 1.8088374876958107 1.7325e-08 1.781707563507311 1.7326e-08 1.784248604187731 1.7327e-08 1.8134430873026148 1.7327999999999998e-08 1.8635459895716244 1.7329e-08 1.7976917349032497 1.733e-08 1.8324093016842695 1.7330999999999998e-08 1.7946257620057438 1.7332e-08 1.7925930641647598 1.7333e-08 1.7683939448713342 1.7333999999999998e-08 1.746492717309714 1.7335e-08 1.6839503219711818 1.7336e-08 1.8097889794920827 1.7336999999999998e-08 1.8341688731818682 1.7338e-08 1.7496653702958913 1.7339e-08 1.8369432220206618 1.734e-08 1.765637594802424 1.7341e-08 1.8612675008278488 1.7342e-08 1.7724901874892345 1.7343e-08 1.7467653286522473 1.7344e-08 1.7761910081800976 1.7345e-08 1.812965198475214 1.7346e-08 1.8457354484797615 1.7347e-08 1.80688823711448 1.7348e-08 1.8344771942517502 1.7349e-08 1.7840894469664654 1.735e-08 1.764395713513359 1.7351e-08 1.841564774616907 1.7352e-08 1.711704985198534 1.7353e-08 1.811063376649343 1.7354e-08 1.8075987890892258 1.7355e-08 1.9147881277543866 1.7356e-08 1.8062103632543915 1.7357e-08 1.8412299322250303 1.7358e-08 1.849391863144353 1.7359e-08 1.8505536495209407 1.736e-08 1.7367817198632756 1.7361e-08 1.8197724167798346 1.7362e-08 1.7739400296342849 1.7362999999999998e-08 1.809890391177785 1.7364e-08 1.8298087235400675 1.7365e-08 1.8021194823081397 1.7365999999999998e-08 1.7786971180606603 1.7367e-08 1.7595134238483394 1.7368e-08 1.7589043988834685 1.7368999999999998e-08 1.7446020293956408 1.737e-08 1.7960414871528545 1.7371e-08 1.7477583950207933 1.7371999999999998e-08 1.7355937794304799 1.7373e-08 1.8297787313671243 1.7374e-08 1.7961200402587498 1.7375e-08 1.8044368326404663 1.7376e-08 1.7306747132112397 1.7377e-08 1.7570688615711614 1.7378e-08 1.8500909678288868 1.7379e-08 1.7268522104667356 1.738e-08 1.7942381092096047 1.7381e-08 1.8467135239814199 1.7382e-08 1.745157936094732 1.7383e-08 1.859817932997348 1.7384e-08 1.763716142515955 1.7385e-08 1.8594056182086474 1.7386e-08 1.8890445926951205 1.7387e-08 1.7076305591229053 1.7388e-08 1.8381434790000113 1.7389e-08 1.8156448319091278 1.739e-08 1.7690539992650534 1.7391e-08 1.7216605366242983 1.7392e-08 1.8585504633841403 1.7393e-08 1.7334060662958874 1.7394e-08 1.8148734420641373 1.7395e-08 1.8235712407338696 1.7396e-08 1.9265964215554672 1.7397e-08 1.8189430072294226 1.7397999999999998e-08 1.8091693211222204 1.7399e-08 1.8128551665848218 1.74e-08 1.8329252087145587 1.7400999999999998e-08 1.7870705552236723 1.7402e-08 1.8328975194890282 1.7403e-08 1.774525846951406 1.7403999999999998e-08 1.777732975290645 1.7405e-08 1.7132116657173442 1.7406e-08 1.844045477859669 1.7406999999999998e-08 1.8088952994873355 1.7408e-08 1.7317954150982298 1.7409e-08 1.8976385184314941 1.741e-08 1.8085251272204073 1.7411e-08 1.8729337060469722 1.7412e-08 1.7642646279932734 1.7413e-08 1.8358492870511676 1.7414e-08 1.7727414939028416 1.7415e-08 1.7651650714098785 1.7416e-08 1.873550467338013 1.7417e-08 1.7480931328387705 1.7418e-08 1.775584427111038 1.7419e-08 1.8331347987403994 1.742e-08 1.8490978487676706 1.7421e-08 1.7662245769498566 1.7422e-08 1.7719984019147965 1.7423e-08 1.7881116027525086 1.7424e-08 1.8108526899487998 1.7425e-08 1.8559884916563179 1.7426e-08 1.7961832389023995 1.7427e-08 1.7706782467100863 1.7428e-08 1.8282237546118636 1.7429e-08 1.7949685182308628 1.743e-08 1.8153798937062608 1.7431e-08 1.8422480383154507 1.7432e-08 1.762746151534756 1.7432999999999998e-08 1.8087336770249294 1.7434e-08 1.9416703126753427 1.7435e-08 1.8196353394716362 1.7435999999999998e-08 1.7776799939576697 1.7437e-08 1.7168149531841248 1.7438e-08 1.8300986050054575 1.7438999999999998e-08 1.8622218845228578 1.744e-08 1.7648253298846135 1.7441e-08 1.7960506474339546 1.7441999999999998e-08 1.8238007939566196 1.7443e-08 1.820737618996587 1.7444e-08 1.7319475857358977 1.7445e-08 1.8620559396653653 1.7446e-08 1.84982064672608 1.7447e-08 1.7357102054788867 1.7448e-08 1.7983740986642545 1.7449e-08 1.6766993262703334 1.745e-08 1.7834765853468608 1.7451e-08 1.8187785777773358 1.7452e-08 1.8083156006217331 1.7453e-08 1.7490463073267128 1.7454e-08 1.8540903878893509 1.7455e-08 1.81008637855656 1.7456e-08 1.7546861324362946 1.7457e-08 1.7712667003635896 1.7458e-08 1.8725684716637485 1.7459e-08 1.7071143763701448 1.746e-08 1.8289328882730203 1.7461e-08 1.754212858300922 1.7462e-08 1.8066115886286223 1.7463e-08 1.8303530228188098 1.7464e-08 1.8773433215651747 1.7465e-08 1.772291327263236 1.7466e-08 1.7287416921687595 1.7467e-08 1.7550538816868542 1.7467999999999998e-08 1.7458248416044448 1.7469e-08 1.7486003506311638 1.747e-08 1.9392452332066084 1.7470999999999998e-08 1.8130947651446137 1.7472e-08 1.7760421445796268 1.7473e-08 1.7862978912614726 1.7473999999999998e-08 1.7139542348372037 1.7475e-08 1.832028521045686 1.7476e-08 1.823117629069638 1.7476999999999998e-08 1.864171891673778 1.7478e-08 1.8046998420912763 1.7479e-08 1.8307835462304498 1.748e-08 1.8206913568305163 1.7481e-08 1.7793130082211104 1.7482e-08 1.8185948817096071 1.7483e-08 1.8638764034986763 1.7484e-08 1.8126194106459386 1.7485e-08 1.6877417527728762 1.7486e-08 1.7489865938324478 1.7487e-08 1.7368478141785257 1.7488e-08 1.7975642782384225 1.7489e-08 1.858958237282588 1.749e-08 1.8858325951374537 1.7491e-08 1.801545301676786 1.7492e-08 1.8226616393610118 1.7493e-08 1.909172435032743 1.7494e-08 1.8412965563315753 1.7495e-08 1.8034019420282394 1.7496e-08 1.768801676550414 1.7497e-08 1.8449102582995927 1.7498e-08 1.8446350860757874 1.7499e-08 1.7695709805632824 1.75e-08 1.8230095038141414 1.7501e-08 1.7701096339839402 1.7502e-08 1.8279670796332472 1.7503e-08 1.7628393550192256 1.7504e-08 1.7811784556967487 1.7505e-08 1.8689035240213314 1.7505999999999998e-08 1.829388650430994 1.7507e-08 1.8806100246856396 1.7508e-08 1.8123461402545828 1.7508999999999998e-08 1.7770805434664696 1.751e-08 1.827573191836964 1.7511e-08 1.8310335992007802 1.7511999999999998e-08 1.7390854467191639 1.7513e-08 1.8431964157120053 1.7514e-08 1.7112800306495672 1.7515e-08 1.9023800365897907 1.7516e-08 1.6732840881767523 1.7517e-08 1.8003109637484562 1.7518e-08 1.76362921800256 1.7519e-08 1.7122973916020454 1.752e-08 1.7505056952510343 1.7521e-08 1.8026934287357033 1.7522e-08 1.699629377729767 1.7523e-08 1.8081877831987396 1.7524e-08 1.7346916415204063 1.7525e-08 1.7579996758422285 1.7526e-08 1.7690983536655929 1.7527e-08 1.8458869117594594 1.7528e-08 1.8044367900840543 1.7529e-08 1.7767459295786636 1.753e-08 1.7708856644706963 1.7531e-08 1.8054418694371235 1.7532e-08 1.7082009182484412 1.7533e-08 1.8893195261293645 1.7534e-08 1.7795331208862595 1.7535e-08 1.7528949908304434 1.7536e-08 1.8236428017249255 1.7537e-08 1.8254185859595344 1.7538e-08 1.7954851194867594 1.7539e-08 1.807368747301546 1.754e-08 1.8453870888886479 1.7540999999999998e-08 1.822957696022806 1.7542e-08 1.725822478653364 1.7543e-08 1.8960736346414824 1.7543999999999998e-08 1.7646500603534059 1.7545e-08 1.7745394563720638 1.7546e-08 1.840728142854404 1.7546999999999998e-08 1.7872327367294731 1.7548e-08 1.781092616746997 1.7549e-08 1.851848575723807 1.7549999999999998e-08 1.8304972776711694 1.7551e-08 1.8145269606940968 1.7552e-08 1.7990630025008656 1.7553e-08 1.7790714462418762 1.7554e-08 1.8132753577464762 1.7555e-08 1.8109493582672544 1.7556e-08 1.753671595416849 1.7557e-08 1.7774775433966825 1.7558e-08 1.7693802086774688 1.7559e-08 1.788926199433963 1.756e-08 1.673367702477826 1.7561e-08 1.7706665674127997 1.7562e-08 1.7581819094910924 1.7563e-08 1.7869493254669089 1.7564e-08 1.7685325203890745 1.7565e-08 1.717978497195369 1.7566e-08 1.7318683991974229 1.7567e-08 1.8145888013083804 1.7568e-08 1.7655364298420941 1.7569e-08 1.8826004823753495 1.757e-08 1.7658789973584925 1.7571e-08 1.6975498639870674 1.7572e-08 1.8083827473156722 1.7573e-08 1.8490698181055856 1.7574e-08 1.7757400708756905 1.7575e-08 1.8374325209004396 1.7575999999999998e-08 1.900020103685394 1.7577e-08 1.7072900773164816 1.7578e-08 1.7897844479792255 1.7578999999999998e-08 1.754492007683691 1.758e-08 1.7656947394658604 1.7581e-08 1.7545721105433536 1.7581999999999998e-08 1.7331839998067142 1.7583e-08 1.8987505535846745 1.7584e-08 1.6936988039383984 1.7584999999999998e-08 1.809397270289243 1.7586e-08 1.823090686351697 1.7587e-08 1.8276686066154655 1.7588e-08 1.7915789585240598 1.7589e-08 1.8777771303471742 1.759e-08 1.7558587141614284 1.7591e-08 1.7097679098692273 1.7592e-08 1.7769382764273371 1.7593e-08 1.7558694772165069 1.7594e-08 1.8279159147925574 1.7595e-08 1.7422967318171485 1.7596e-08 1.8471830168011583 1.7597e-08 1.7766634308101092 1.7598e-08 1.8426172506780976 1.7599e-08 1.7926377714398913 1.76e-08 1.7563745228116612 1.7601e-08 1.8746830974139497 1.7602e-08 1.7470760186889025 1.7603e-08 1.8130678331061685 1.7604e-08 1.7827626871462012 1.7605e-08 1.6821292599885125 1.7606e-08 1.7514745880351816 1.7607e-08 1.7522081678654386 1.7608e-08 1.8143258035258618 1.7609e-08 1.8264696213473812 1.761e-08 1.7738836252476726 1.7610999999999998e-08 1.7099383377959627 1.7612e-08 1.7602960441748097 1.7613e-08 1.7111397516761653 1.7613999999999998e-08 1.8970554701312152 1.7615e-08 1.7994729871205726 1.7616e-08 1.7232925051027612 1.7616999999999998e-08 1.8472033271512822 1.7618e-08 1.8153097574816115 1.7619e-08 1.7469511624592278 1.7619999999999998e-08 1.8221537782998736 1.7621e-08 1.6841301036584477 1.7622e-08 1.849274164145935 1.7623e-08 1.7893496386585361 1.7624e-08 1.7837567810246502 1.7625e-08 1.8321682967998925 1.7626e-08 1.7868486811649396 1.7627e-08 1.862417271922537 1.7628e-08 1.724994837723865 1.7629e-08 1.7907719805377655 1.763e-08 1.7986073113337697 1.7631e-08 1.7449467700758905 1.7632e-08 1.7599259639413183 1.7633e-08 1.7388883930655779 1.7634e-08 1.7470442425739228 1.7635e-08 1.8558964229151598 1.7636e-08 1.8364675474704963 1.7637e-08 1.7940115086064543 1.7638e-08 1.7808735691056614 1.7639e-08 1.8626836250588483 1.764e-08 1.8953236506867637 1.7641e-08 1.7872472938104096 1.7642e-08 1.797106618351548 1.7643e-08 1.746277122397015 1.7644e-08 1.8915887116342127 1.7645e-08 1.7640821100052961 1.7645999999999998e-08 1.8454547241646384 1.7647e-08 1.7764827452049028 1.7648e-08 1.8619685630698435 1.7648999999999998e-08 1.7803586667740987 1.765e-08 1.7806451962044405 1.7651e-08 1.7745084800144806 1.7651999999999998e-08 1.8048727094501993 1.7653e-08 1.8250785001726095 1.7654e-08 1.813669383087185 1.7654999999999998e-08 1.8193562529435825 1.7656e-08 1.808252530636576 1.7657e-08 1.7588878205847585 1.7658e-08 1.8648468555192037 1.7659e-08 1.7327332477119342 1.766e-08 1.7688779770216456 1.7661e-08 1.7334282253121476 1.7662e-08 1.7515246925226224 1.7663e-08 1.8129137925934742 1.7664e-08 1.8144661110785187 1.7665e-08 1.7222492966323175 1.7666e-08 1.747829056091484 1.7667e-08 1.768434068210745 1.7668e-08 1.7348480882109347 1.7669e-08 1.7214905486571626 1.767e-08 1.8093757451491868 1.7671e-08 1.8762367122311496 1.7672e-08 1.8692483631658652 1.7673e-08 1.7957449197543596 1.7674e-08 1.7695660947943264 1.7675e-08 1.7631218450308341 1.7676e-08 1.731720128231714 1.7677e-08 1.7265851284953102 1.7678e-08 1.7996648334540815 1.7679e-08 1.789447345571398 1.768e-08 1.778175656059434 1.7681e-08 1.8379056861421204 1.7682e-08 1.7669546156584346 1.7683e-08 1.799505009189882 1.7683999999999998e-08 1.8128436972602977 1.7685e-08 1.8354063218540222 1.7686e-08 1.8075214507367774 1.7686999999999998e-08 1.7285722190916843 1.7688e-08 1.7639192360623832 1.7689e-08 1.7158527531374512 1.7689999999999998e-08 1.847760660032964 1.7691e-08 1.8278475283777167 1.7692e-08 1.8395580707917696 1.7693e-08 1.8449295194696664 1.7694e-08 1.789359510240214 1.7695e-08 1.8523651654557154 1.7696e-08 1.775879345379985 1.7697e-08 1.7803829265443814 1.7698e-08 1.771399664958231 1.7699e-08 1.8190541288477116 1.77e-08 1.75136712315087 1.7701e-08 1.8226444109139512 1.7702e-08 1.8541713070522174 1.7703e-08 1.8738748996052057 1.7704e-08 1.756820366731235 1.7705e-08 1.8313115716032977 1.7706e-08 1.7117172124975508 1.7707e-08 1.793536396599175 1.7708e-08 1.8091789358923047 1.7709e-08 1.7942727149692395 1.771e-08 1.828209813264012 1.7711e-08 1.8739912133327266 1.7712e-08 1.8789307532966322 1.7713e-08 1.7983792404924535 1.7714e-08 1.811002986128525 1.7715e-08 1.7670267235809571 1.7716e-08 1.7421487798492976 1.7717e-08 1.8008789981631022 1.7718e-08 1.8603600581266888 1.7718999999999998e-08 1.8288209442532233 1.772e-08 1.7593999692361204 1.7721e-08 1.7467568671820182 1.7721999999999998e-08 1.830779233729812 1.7723e-08 1.7967468762323535 1.7724e-08 1.8462048510808509 1.7724999999999998e-08 1.727315225563156 1.7726e-08 1.8584968888983182 1.7727e-08 1.7801255508816884 1.7727999999999998e-08 1.7682656934625112 1.7729e-08 1.7948135601016393 1.773e-08 1.8081703596759557 1.7731e-08 1.7675597006179138 1.7732e-08 1.790034367463857 1.7733e-08 1.794391982689264 1.7734e-08 1.8029952945124554 1.7735e-08 1.7718557376830684 1.7736e-08 1.8301964680174787 1.7737e-08 1.9316784945277745 1.7738e-08 1.8205494289560473 1.7739e-08 1.819238557568138 1.774e-08 1.8138448122345647 1.7741e-08 1.8197300783481907 1.7742e-08 1.807572224797131 1.7743e-08 1.7917262006842472 1.7744e-08 1.7941409012391176 1.7745e-08 1.7705500672193992 1.7746e-08 1.722190845531331 1.7747e-08 1.8092741979068048 1.7748e-08 1.8221187571310127 1.7749e-08 1.8282586341488873 1.775e-08 1.864040416550806 1.7751e-08 1.846630001532795 1.7752e-08 1.6698216561997652 1.7753e-08 1.8693624109086389 1.7753999999999998e-08 1.8176444451757512 1.7755e-08 1.7879840828287203 1.7756e-08 1.8049505656337883 1.7756999999999998e-08 1.7845318655705582 1.7758e-08 1.7779270287788649 1.7759e-08 1.7929385148981496 1.7759999999999998e-08 1.863479663942564 1.7761e-08 1.7987811609496331 1.7762e-08 1.7990417358557165 1.7762999999999998e-08 1.8067047182570306 1.7764e-08 1.8648389955720803 1.7765e-08 1.7956347909871626 1.7766e-08 1.8601523878022774 1.7767e-08 1.809302842976226 1.7768e-08 1.8916206684729895 1.7769e-08 1.8273863677734807 1.777e-08 1.8391361686607315 1.7771e-08 1.8035663810008946 1.7772e-08 1.7445226620046843 1.7773e-08 1.8116819974150726 1.7774e-08 1.8757577500014455 1.7775e-08 1.8251510032532374 1.7776e-08 1.8018565372683757 1.7777e-08 1.9198331362520569 1.7778e-08 1.8238111520178588 1.7779e-08 1.970265325408709 1.778e-08 1.808908649715637 1.7781e-08 1.8244682378258184 1.7782e-08 1.8403938410767111 1.7783e-08 1.8250301858962827 1.7784e-08 1.8013976563028633 1.7785e-08 1.8556357572241686 1.7786e-08 1.7540758451240137 1.7787e-08 1.8134832700857662 1.7788e-08 1.8423782557530524 1.7788999999999998e-08 1.787900652370193 1.779e-08 1.788033859714361 1.7791e-08 1.753630748779444 1.7791999999999998e-08 1.7838569182393806 1.7793e-08 1.8294631339999525 1.7794e-08 1.7115744886072732 1.7794999999999998e-08 1.7944024524841926 1.7796e-08 1.7578286805974277 1.7797e-08 1.7331606476038377 1.7797999999999998e-08 1.7915453508228643 1.7799e-08 1.7634520727998866 1.78e-08 1.732399162916275 1.7801e-08 1.801322798308403 1.7802e-08 1.7611782570407641 1.7803e-08 1.8293894834176763 1.7804e-08 1.8673676656792069 1.7805e-08 1.776400637682531 1.7806e-08 1.8195841425671808 1.7807e-08 1.7705837089332581 1.7808e-08 1.8023147384591431 1.7809e-08 1.7976104169474094 1.781e-08 1.8006538348268284 1.7811e-08 1.8257636213482609 1.7812e-08 1.7740295228502598 1.7813e-08 1.801008021948426 1.7814e-08 1.7319028833550485 1.7815e-08 1.8460585374581884 1.7816e-08 1.8215857812215792 1.7817e-08 1.8354893499707976 1.7818e-08 1.8097052791459765 1.7819e-08 1.7626975169837467 1.782e-08 1.8113410186070054 1.7821e-08 1.7904689924861081 1.7822e-08 1.7478416882102374 1.7823e-08 1.8013957083396812 1.7823999999999998e-08 1.8365496902004035 1.7825e-08 1.8252609735513774 1.7826e-08 1.7503707209801787 1.7826999999999998e-08 1.848565873710367 1.7828e-08 1.8727972446882253 1.7829e-08 1.7780090115649902 1.7829999999999998e-08 1.890640392865932 1.7831e-08 1.7759411575310124 1.7832e-08 1.7362355659251179 1.7832999999999998e-08 1.7929250111028847 1.7834e-08 1.8129144040791738 1.7835e-08 1.7923557017539964 1.7836e-08 1.8124401253531581 1.7837e-08 1.766913752441769 1.7838e-08 1.784891480482248 1.7839e-08 1.8132954319373824 1.784e-08 1.7607128638466738 1.7841e-08 1.79985809860307 1.7842e-08 1.7361052541617625 1.7843e-08 1.8538612367256944 1.7844e-08 1.738139994637967 1.7845e-08 1.8491966184978754 1.7846e-08 1.7840404056704788 1.7847e-08 1.8662015276465072 1.7848e-08 1.8288075096032326 1.7849e-08 1.9154439545560136 1.785e-08 1.8128148702073554 1.7851e-08 1.8003615428587443 1.7852e-08 1.8170649189419659 1.7853e-08 1.672440544084477 1.7854e-08 1.8128581925114489 1.7855e-08 1.682590564916068 1.7856e-08 1.7679196694849908 1.7857e-08 1.7420863235309207 1.7858e-08 1.799890704814746 1.7858999999999998e-08 1.8791035223466506 1.786e-08 1.817313265812241 1.7861e-08 1.7635369338568916 1.7861999999999998e-08 1.7992800253696433 1.7863e-08 1.7564233792095267 1.7864e-08 1.8478073468892429 1.7864999999999998e-08 1.6786798269090502 1.7866e-08 1.7583083718100512 1.7867e-08 1.7955830949693372 1.7867999999999998e-08 1.8211162396008505 1.7869e-08 1.839381196064175 1.787e-08 1.8121689883165848 1.7871e-08 1.836553138714895 1.7872e-08 1.7712150894872 1.7873e-08 1.787140643796975 1.7874e-08 1.725408537063772 1.7875e-08 1.7908208403976917 1.7876e-08 1.770626348829257 1.7877e-08 1.8489668746180061 1.7878e-08 1.740095214969004 1.7879e-08 1.7805708203399244 1.788e-08 1.7723178191106428 1.7881e-08 1.8372324547044832 1.7882e-08 1.8230606292688138 1.7883e-08 1.811195449599189 1.7884e-08 1.6958803187166653 1.7885e-08 1.8044743837052775 1.7886e-08 1.7743275920422754 1.7887e-08 1.8370752316648025 1.7888e-08 1.7406834489865701 1.7889e-08 1.7567168850216952 1.789e-08 1.7321461376766052 1.7891e-08 1.7757519526954606 1.7892e-08 1.8282675024771418 1.7893e-08 1.8511810503345996 1.7894e-08 1.760074632033302 1.7895e-08 1.7707886736418865 1.7896e-08 1.7686368900243465 1.7896999999999998e-08 1.8690089935835978 1.7898e-08 1.761702083362253 1.7899e-08 1.7835834397241752 1.7899999999999998e-08 1.8207637818859552 1.7901e-08 1.725278152079221 1.7902e-08 1.856095882331694 1.7902999999999998e-08 1.849762737779097 1.7904e-08 1.7423846309942759 1.7905e-08 1.7266015612829666 1.7905999999999998e-08 1.873078828134455 1.7907e-08 1.8946642774119624 1.7908e-08 1.8145428888609452 1.7909e-08 1.7081544931270403 1.791e-08 1.8099132100302087 1.7911e-08 1.8049758021884752 1.7912e-08 1.8190563063847949 1.7913e-08 1.74747306025124 1.7914e-08 1.7474499956673777 1.7915e-08 1.7694824901108048 1.7916e-08 1.831869778345877 1.7917e-08 1.7492506718992367 1.7918e-08 1.7644334202244614 1.7919e-08 1.7549477721312128 1.792e-08 1.776378447442743 1.7921e-08 1.7482420125502405 1.7922e-08 1.770440088102134 1.7923e-08 1.7924299072394847 1.7924e-08 1.8157906622585844 1.7925e-08 1.8049881171618898 1.7926e-08 1.8611490909496986 1.7927e-08 1.7800780151651607 1.7928e-08 1.772375091882009 1.7929e-08 1.7884096167646615 1.793e-08 1.8509417092565874 1.7931e-08 1.8034213099540604 1.7931999999999998e-08 1.7413032833856235 1.7933e-08 1.8711689863340877 1.7934e-08 1.8402465692915322 1.7934999999999998e-08 1.8016514001044068 1.7936e-08 1.8658013478880067 1.7937e-08 1.8049138559287743 1.7937999999999998e-08 1.8950211513108355 1.7939e-08 1.898383438180402 1.794e-08 1.8679275808631637 1.7940999999999998e-08 1.826878530835128 1.7942e-08 1.8635445106838353 1.7943e-08 1.6654233924865172 1.7944e-08 1.7739898654832231 1.7945e-08 1.844438442111823 1.7946e-08 1.7807128916760884 1.7947e-08 1.7308214726183877 1.7948e-08 1.775448680134076 1.7949e-08 1.7468500587139149 1.795e-08 1.8516695296546708 1.7951e-08 1.7763307206659527 1.7952e-08 1.7575832320216698 1.7953e-08 1.7976844835191792 1.7954e-08 1.8232944694938114 1.7955e-08 1.800431035944839 1.7956e-08 1.8002077145216322 1.7957e-08 1.844489950247816 1.7958e-08 1.7995583187681927 1.7959e-08 1.8006630663046774 1.796e-08 1.7820619606423234 1.7961e-08 1.8658793854141054 1.7962e-08 1.8570855461309888 1.7963e-08 1.8666163998517473 1.7964e-08 1.8081847798387718 1.7965e-08 1.7868242855010261 1.7966e-08 1.7306339681460807 1.7966999999999998e-08 1.7095446918505284 1.7968e-08 1.8342681050575815 1.7969e-08 1.829768516000102 1.7969999999999998e-08 1.8686906649931254 1.7971e-08 1.8159174486463818 1.7972e-08 1.7903107535019824 1.7972999999999998e-08 1.7797692695451852 1.7974e-08 1.7615542968324767 1.7975e-08 1.7762692837174023 1.7975999999999998e-08 1.725468144561729 1.7977e-08 1.9066947673425596 1.7978e-08 1.7933677130709924 1.7979e-08 1.7173686443884462 1.798e-08 1.8699991656277613 1.7981e-08 1.782386859173952 1.7982e-08 1.7460417458274333 1.7983e-08 1.7740625997916255 1.7984e-08 1.8250743518351982 1.7985e-08 1.7451012944364122 1.7986e-08 1.8525231882269493 1.7987e-08 1.7469258723748893 1.7988e-08 1.817249518482286 1.7989e-08 1.8896563974495864 1.799e-08 1.7953955071127312 1.7991e-08 1.7654540888856862 1.7992e-08 1.7485125831578496 1.7993e-08 1.7559485668576094 1.7994e-08 1.8470727308662362 1.7995e-08 1.9212282773025606 1.7996e-08 1.8818692751673998 1.7997e-08 1.7875321719927384 1.7998e-08 1.792780964797997 1.7999e-08 1.7892084085614381 1.8e-08 1.7527151335397007 1.8001e-08 1.8202936997870076 1.8001999999999998e-08 1.7982563559148312 1.8003e-08 1.789531822662026 1.8004e-08 1.8518855087511479 1.8004999999999998e-08 1.8780601453943364 1.8006e-08 1.7325445062355904 1.8007e-08 1.8184528304144065 1.8007999999999998e-08 1.733409304849378 1.8009e-08 1.8357497562594896 1.801e-08 1.8149438347014868 1.8010999999999998e-08 1.8386407528797633 1.8012e-08 1.8350321152301348 1.8013e-08 1.7739603904261496 1.8014e-08 1.8340709540976075 1.8015e-08 1.7912577334737827 1.8016e-08 1.7233945097800465 1.8017e-08 1.783341782977264 1.8018e-08 1.8659381434476017 1.8019e-08 1.8423689287890863 1.802e-08 1.7845087787789655 1.8021e-08 1.8583796690473489 1.8022e-08 1.807886103197107 1.8023e-08 1.8965229565340718 1.8024e-08 1.8282834062229 1.8025e-08 1.7719301695356926 1.8026e-08 1.878214975556245 1.8027e-08 1.7789400119899592 1.8028e-08 1.7682072865405012 1.8029e-08 1.853585193336149 1.803e-08 1.7972554835043415 1.8031e-08 1.766010632699554 1.8032e-08 1.7708197077077554 1.8033e-08 1.856417415788328 1.8034e-08 1.9172326378382922 1.8035e-08 1.7393854611824735 1.8036e-08 1.8267970712894017 1.8036999999999998e-08 1.7661287438262447 1.8038e-08 1.8142606299858965 1.8039e-08 1.7510851380398555 1.8039999999999998e-08 1.763311201808118 1.8041e-08 1.8071514696186752 1.8042e-08 1.7179000068815455 1.8042999999999998e-08 1.7937431266571866 1.8044e-08 1.7669501719384109 1.8045e-08 1.9121395836121855 1.8045999999999998e-08 1.776367689188677 1.8047e-08 1.7302123164037286 1.8048e-08 1.7627735798618112 1.8049e-08 1.780468421203604 1.805e-08 1.7799666996175298 1.8051e-08 1.6716729312384293 1.8052e-08 1.8429303262211076 1.8053e-08 1.827328170342169 1.8054e-08 1.842312279927619 1.8055e-08 1.8210614249260009 1.8056e-08 1.774037379441615 1.8057e-08 1.7717511145767844 1.8058e-08 1.8282456535479497 1.8059e-08 1.7801924895506798 1.806e-08 1.6981065134605127 1.8061e-08 1.8402489205253574 1.8062e-08 1.8275108597138614 1.8063e-08 1.7933827545424104 1.8064e-08 1.722575314663838 1.8065e-08 1.803589090012383 1.8066e-08 1.8217304307709672 1.8067e-08 1.8246360850315384 1.8068e-08 1.8845127885701303 1.8069e-08 1.8474576634229098 1.807e-08 1.812184412965677 1.8071e-08 1.8261228197624566 1.8072e-08 1.7559873247046365 1.8073e-08 1.9304721831548561 1.8074e-08 1.7650555417431704 1.8074999999999998e-08 1.8495208263032998 1.8076e-08 1.7519074540435449 1.8077e-08 1.8020207070588106 1.8077999999999998e-08 1.766634736123582 1.8079e-08 1.863706996925119 1.808e-08 1.881295013236169 1.8080999999999998e-08 1.8970286146158444 1.8082e-08 1.8011400822908086 1.8083e-08 1.8063897932268844 1.8084e-08 1.7936800744798542 1.8085e-08 1.848728343516871 1.8086e-08 1.7202716676085112 1.8087e-08 1.8467074629920586 1.8088e-08 1.801481489844213 1.8089e-08 1.8187012426475677 1.809e-08 1.8461343376258244 1.8091e-08 1.8904600556584277 1.8092e-08 1.8125320815011017 1.8093e-08 1.7652047736674479 1.8094e-08 1.751865311734465 1.8095e-08 1.84312521981056 1.8096e-08 1.8023284202204872 1.8097e-08 1.809691614837657 1.8098e-08 1.8225113582950994 1.8099e-08 1.805585539953271 1.81e-08 1.8708217837308432 1.8101e-08 1.6828375126968014 1.8102e-08 1.7482288849202874 1.8103e-08 1.7630583073266222 1.8104e-08 1.8240902739975862 1.8105e-08 1.8501189643791225 1.8106e-08 1.699733202750124 1.8107e-08 1.8028552809523481 1.8108e-08 1.8111046319305057 1.8109e-08 1.7778280092939969 1.8109999999999998e-08 1.857957042296011 1.8111e-08 1.8544054694446663 1.8112e-08 1.7999007186450966 1.8112999999999998e-08 1.8004376143957006 1.8114e-08 1.8395372633856208 1.8115e-08 1.779635452628527 1.8115999999999998e-08 1.7772543995322307 1.8117e-08 1.9034380323983886 1.8118e-08 1.7985414213892315 1.8118999999999998e-08 1.8499651383476825 1.812e-08 1.8261073055831585 1.8121e-08 1.8262390069150056 1.8122e-08 1.8128557009375845 1.8123e-08 1.7635364090296581 1.8124e-08 1.7655318436238925 1.8125e-08 1.8018304958937772 1.8126e-08 1.749495508985642 1.8127e-08 1.742651499010393 1.8128e-08 1.8811117294032453 1.8129e-08 1.836132927972203 1.813e-08 1.8034303240756873 1.8131e-08 1.8671908712238015 1.8132e-08 1.8219103454725603 1.8133e-08 1.7927014748302421 1.8134e-08 1.6753361286990056 1.8135e-08 1.7440848296940288 1.8136e-08 1.8445906403564465 1.8137e-08 1.7303661966328632 1.8138e-08 1.8093243553431335 1.8139e-08 1.7362449595917313 1.814e-08 1.8810440322136845 1.8141e-08 1.7624116978254418 1.8142e-08 1.6984614841899681 1.8143e-08 1.7935379884620763 1.8144e-08 1.7747135077482392 1.8144999999999998e-08 1.6963241395948687 1.8146e-08 1.7877991857346542 1.8147e-08 1.7250608081212706 1.8147999999999998e-08 1.8494285554893126 1.8149e-08 1.7172674703478696 1.815e-08 1.7632599412953502 1.8150999999999998e-08 1.8175288683300628 1.8152e-08 1.8214292620884711 1.8153e-08 1.8121723042238138 1.8153999999999998e-08 1.7215461776176002 1.8155e-08 1.8002437244544964 1.8156e-08 1.8082067155951342 1.8157e-08 1.7390639988119962 1.8158e-08 1.7857303603062042 1.8159e-08 1.776904585208722 1.816e-08 1.8345810871196144 1.8161e-08 1.7919892833516051 1.8162e-08 1.7588245607622301 1.8163e-08 1.7743393904100695 1.8164e-08 1.819868419520467 1.8165e-08 1.784862365087381 1.8166e-08 1.7622395386871108 1.8167e-08 1.8015701208730845 1.8168e-08 1.7279918290095906 1.8169e-08 1.828674696748548 1.817e-08 1.8826675178705266 1.8171e-08 1.8865192252082086 1.8172e-08 1.7713231634186035 1.8173e-08 1.8361240465011053 1.8174e-08 1.6394778180775362 1.8175e-08 1.797113660452671 1.8176e-08 1.7779675551608418 1.8177e-08 1.7967612606711292 1.8178e-08 1.7434834271265363 1.8179e-08 1.7621902967068546 1.8179999999999998e-08 1.773543277436008 1.8181e-08 1.799681491192144 1.8182e-08 1.757175728335562 1.8182999999999998e-08 1.8658283320913402 1.8184e-08 1.8013214691039974 1.8185e-08 1.7573897132907914 1.8185999999999998e-08 1.8513836678713536 1.8187e-08 1.9077877776056655 1.8188e-08 1.8179751646395703 1.8188999999999998e-08 1.6683614256505548 1.819e-08 1.793662980422248 1.8191e-08 1.7567993918285876 1.8192e-08 1.9234472547849326 1.8193e-08 1.7663230132275989 1.8194e-08 1.7981211311156373 1.8195e-08 1.7833788978297807 1.8196e-08 1.766659696452647 1.8197e-08 1.8284715307917574 1.8198e-08 1.8010500659362008 1.8199e-08 1.8394731965290563 1.82e-08 1.843359258405297 1.8201e-08 1.8050276401204939 1.8202e-08 1.7754193420300801 1.8203e-08 1.7969105147693145 1.8204e-08 1.7699324646181849 1.8205e-08 1.781596052530577 1.8206e-08 1.7931211010477799 1.8207e-08 1.6977325088616215 1.8208e-08 1.8501302032857965 1.8209e-08 1.7462575679583874 1.821e-08 1.7578364247891798 1.8211e-08 1.7611953860365035 1.8212e-08 1.8252797984020181 1.8213e-08 1.7646638866508615 1.8214e-08 1.7817569201279353 1.8214999999999998e-08 1.787714630622384 1.8216e-08 1.8120021911994408 1.8217e-08 1.836185453705681 1.8217999999999998e-08 1.8169443480544853 1.8219e-08 1.772835422649206 1.822e-08 1.8004282841466217 1.8220999999999998e-08 1.777864342462083 1.8222e-08 1.820506599893181 1.8223e-08 1.7771346595886157 1.8223999999999998e-08 1.8373822100162382 1.8225e-08 1.7432474437884642 1.8226e-08 1.820442449832109 1.8227e-08 1.81359462440694 1.8228e-08 1.8465658444093724 1.8229e-08 1.8196068081860926 1.823e-08 1.8035798977344648 1.8231e-08 1.7834795094670122 1.8232e-08 1.7748150504880262 1.8233e-08 1.8506417902130667 1.8234e-08 1.8235610884041835 1.8235e-08 1.7687935938347261 1.8236e-08 1.8390942675006203 1.8237e-08 1.7909273697256092 1.8238e-08 1.7925370142832229 1.8239e-08 1.7961650284363515 1.824e-08 1.7423404963687563 1.8241e-08 1.7802021449034071 1.8242e-08 1.7771177784791647 1.8243e-08 1.7563531568421562 1.8244e-08 1.8003274859849774 1.8245e-08 1.7850291770033493 1.8246e-08 1.8229254422448058 1.8247e-08 1.8367187533160345 1.8248e-08 1.8698354397513164 1.8249e-08 1.7708515218651861 1.8249999999999998e-08 1.7978206300405868 1.8251e-08 1.8587633052980703 1.8252e-08 1.712701298335604 1.8252999999999998e-08 1.7887036914632706 1.8254e-08 1.7376913209071203 1.8255e-08 1.762255725103902 1.8255999999999998e-08 1.8727787233173214 1.8257e-08 1.928828534622197 1.8258e-08 1.8102054759154913 1.8258999999999998e-08 1.7679056024432875 1.826e-08 1.8437373557048191 1.8261e-08 1.745094263176479 1.8262e-08 1.8038885436091439 1.8263e-08 1.815289263768204 1.8264e-08 1.741214320155116 1.8265e-08 1.7978981950286541 1.8266e-08 1.8565742501346771 1.8267e-08 1.8696995578427174 1.8268e-08 1.7443406326520479 1.8269e-08 1.7435221699917691 1.827e-08 1.8476128398069416 1.8271e-08 1.8349394831276429 1.8272e-08 1.8754871754530997 1.8273e-08 1.8265766030465997 1.8274e-08 1.8886890938749623 1.8275e-08 1.7564317578777147 1.8276e-08 1.812328882401262 1.8277e-08 1.7803099467679235 1.8278e-08 1.830976440186396 1.8279e-08 1.8482695287816813 1.828e-08 1.8985451517235363 1.8281e-08 1.8379992173786646 1.8282e-08 1.772990806333844 1.8283e-08 1.796654206980006 1.8284e-08 1.8381217784900636 1.8285e-08 1.7311995809806502 1.8286e-08 1.796261039359417 1.8287e-08 1.9032391709065775 1.8287999999999998e-08 1.8523521231422604 1.8289e-08 1.854988953664324 1.829e-08 1.7992715909771495 1.8290999999999998e-08 1.8708878399641025 1.8292e-08 1.7958935319792906 1.8293e-08 1.8272959763665158 1.8293999999999998e-08 1.801906855283672 1.8295e-08 1.8106174660629477 1.8296e-08 1.7316940608321711 1.8296999999999998e-08 1.7446403474215681 1.8298e-08 1.801036361852771 1.8299e-08 1.8298859336551008 1.83e-08 1.8368662313637594 1.8301e-08 1.7706721049210068 1.8302e-08 1.7402808428677208 1.8303e-08 1.773392480788713 1.8304e-08 1.734717424704734 1.8305e-08 1.8414849783962075 1.8306e-08 1.8926339194978685 1.8307e-08 1.7512679121479495 1.8308e-08 1.8678786462793184 1.8309e-08 1.9037159046163832 1.831e-08 1.81952886790769 1.8311e-08 1.8130526747486309 1.8312e-08 1.7844474493740161 1.8313e-08 1.757313551016395 1.8314e-08 1.7524873222057968 1.8315e-08 1.732364919881098 1.8316e-08 1.8201846145897176 1.8317e-08 1.8159757888319001 1.8318e-08 1.8272745829026784 1.8319e-08 1.777731124960352 1.832e-08 1.8273941018940434 1.8321e-08 1.737232033219264 1.8322e-08 1.8377660926005694 1.8322999999999998e-08 1.8033317884628584 1.8324e-08 1.8064567751913188 1.8325e-08 1.8077397254834935 1.8325999999999998e-08 1.7738217098275118 1.8327e-08 1.8079441780212704 1.8328e-08 1.8352073786082927 1.8328999999999998e-08 1.6731156190174405 1.833e-08 1.7357399287081485 1.8331e-08 1.8146798945500675 1.8331999999999998e-08 1.746084754120358 1.8333e-08 1.8947283181024472 1.8334e-08 1.7926240299727378 1.8335e-08 1.8627377530894775 1.8336e-08 1.85615616500197 1.8337e-08 1.70545336653282 1.8338e-08 1.7870429599827116 1.8339e-08 1.8786075365242012 1.834e-08 1.8310575363892638 1.8341e-08 1.8034183701555417 1.8342e-08 1.832405630240988 1.8343e-08 1.7733079269029857 1.8344e-08 1.8057875357516637 1.8345e-08 1.8495663522073083 1.8346e-08 1.829128368454712 1.8347e-08 1.7297482895353335 1.8348e-08 1.8065418704732434 1.8349e-08 1.8245781151550984 1.835e-08 1.7457116276426516 1.8351e-08 1.8601980102034743 1.8352e-08 1.8367741971383895 1.8353e-08 1.8038513906513935 1.8354e-08 1.8478988272220191 1.8355e-08 1.7764829650302543 1.8356e-08 1.8135997799334866 1.8357e-08 1.811867808206537 1.8357999999999998e-08 1.6720743115118617 1.8359e-08 1.9030952278994375 1.836e-08 1.801383636687564 1.8360999999999998e-08 1.8462198166631725 1.8362e-08 1.7822487049377187 1.8363e-08 1.8103181445966243 1.8363999999999998e-08 1.8067355160941112 1.8365e-08 1.7428707208009386 1.8366e-08 1.7924789918532436 1.8366999999999998e-08 1.8879594411378835 1.8368e-08 1.8076729351463912 1.8369e-08 1.7655490009266295 1.837e-08 1.7854505088443637 1.8371e-08 1.830571313075567 1.8372e-08 1.846368582122103 1.8373e-08 1.8980990276855472 1.8374e-08 1.7938626817612693 1.8375e-08 1.7583470589177992 1.8376e-08 1.846066466330441 1.8377e-08 1.752491899276124 1.8378e-08 1.7566020748593074 1.8379e-08 1.8331073547988512 1.838e-08 1.8140628469109585 1.8381e-08 1.8299623869736814 1.8382e-08 1.8352362139502056 1.8383e-08 1.8310895404754162 1.8384e-08 1.8792983673787655 1.8385e-08 1.774469522519508 1.8386e-08 1.8571025844576994 1.8387e-08 1.8677720239722548 1.8388e-08 1.75111386541839 1.8389e-08 1.7837737277627739 1.839e-08 1.7730472280282337 1.8391e-08 1.8292519219204233 1.8392e-08 1.7666316851358945 1.8392999999999998e-08 1.8375548728435658 1.8394e-08 1.8012124358514572 1.8395e-08 1.7100149005298904 1.8395999999999998e-08 1.739272658512112 1.8397e-08 1.8384934070308416 1.8398e-08 1.8509432763936617 1.8398999999999998e-08 1.7011980958834783 1.84e-08 1.800989427281793 1.8401e-08 1.725374601286744 1.8401999999999998e-08 1.7511555781132557 1.8403e-08 1.7014569366395382 1.8404e-08 1.9137772121807406 1.8405e-08 1.8184701012557998 1.8406e-08 1.757832114955222 1.8407e-08 1.8179746657031841 1.8408e-08 1.7883926800122547 1.8409e-08 1.7952034347008852 1.841e-08 1.8106607952431617 1.8411e-08 1.7827433942728328 1.8412e-08 1.7152050167717297 1.8413e-08 1.80286517471279 1.8414e-08 1.8572899204870679 1.8415e-08 1.8813435460942824 1.8416e-08 1.833081115005859 1.8417e-08 1.8082403476943247 1.8418e-08 1.7329492844470022 1.8419e-08 1.7864466847539309 1.842e-08 1.7902265897176897 1.8421e-08 1.8218595234328239 1.8422e-08 1.7408878629107598 1.8423e-08 1.7435674768712615 1.8424e-08 1.8192044591359098 1.8425e-08 1.800472357415823 1.8426e-08 1.8433887314371227 1.8427e-08 1.715381428897291 1.8427999999999998e-08 1.8109765043546384 1.8429e-08 1.8888103201763111 1.843e-08 1.9398775207548016 1.8430999999999998e-08 1.7729826503070527 1.8432e-08 1.772915350386709 1.8433e-08 1.787014190705195 1.8433999999999998e-08 1.8019535855502589 1.8435e-08 1.7736484796531842 1.8436e-08 1.708763325847166 1.8436999999999998e-08 1.721730082108065 1.8438e-08 1.8792013747925487 1.8439e-08 1.8046595867613267 1.844e-08 1.7603544981359203 1.8441e-08 1.8358659502402779 1.8442e-08 1.8275492839616745 1.8443e-08 1.8185007550076684 1.8444e-08 1.8188922569809045 1.8445e-08 1.8907793720689012 1.8446e-08 1.7859609475120513 1.8447e-08 1.801664423259092 1.8448e-08 1.7264861704153116 1.8449e-08 1.8203562605219967 1.845e-08 1.7055029343018866 1.8451e-08 1.850093557544782 1.8452e-08 1.7744850286593439 1.8453e-08 1.6988888210574282 1.8454e-08 1.8572443205183642 1.8455e-08 1.890015527712944 1.8456e-08 1.7927487478831983 1.8457e-08 1.8403454121476959 1.8458e-08 1.8480649595615164 1.8459e-08 1.7657146340921461 1.846e-08 1.8498825958685807 1.8461e-08 1.7207552996654816 1.8462e-08 1.774338143548963 1.8463e-08 1.8209757235563024 1.8464e-08 1.8756715047550485 1.8465e-08 1.800317606089267 1.8465999999999998e-08 1.8124385849977311 1.8467e-08 1.7975551744028984 1.8468e-08 1.7358870061807696 1.8468999999999998e-08 1.7574243656944522 1.847e-08 1.7484910164256895 1.8471e-08 1.9081006454587597 1.8471999999999998e-08 1.6913913192925267 1.8473e-08 1.7640061306158663 1.8474e-08 1.8000363900257894 1.8474999999999998e-08 1.8223097290569583 1.8476e-08 1.892811876430689 1.8477e-08 1.7868832884724661 1.8478e-08 1.803098625712152 1.8479e-08 1.8182724794344547 1.848e-08 1.8088313612352849 1.8481e-08 1.7732535027755745 1.8482e-08 1.8083529612447435 1.8483e-08 1.818632326685405 1.8484e-08 1.7524446150966657 1.8485e-08 1.8385956646938504 1.8486e-08 1.8183530165693405 1.8487e-08 1.75257267438489 1.8488e-08 1.8685099502945886 1.8489e-08 1.945083273265975 1.849e-08 1.7707187643274247 1.8491e-08 1.8745876818429326 1.8492e-08 1.7096285569242835 1.8493e-08 1.8580944920307008 1.8494e-08 1.7935410892223387 1.8495e-08 1.7631479997544544 1.8496e-08 1.776221529540159 1.8497e-08 1.8013295489191479 1.8498e-08 1.7558623960152855 1.8499e-08 1.8264611680479972 1.85e-08 1.781971534825474 1.8500999999999998e-08 1.8250846127460227 1.8502e-08 1.8548679911521964 1.8503e-08 1.9046355970662123 1.8503999999999998e-08 1.8691230264853629 1.8505e-08 1.8317761834871034 1.8506e-08 1.83001006890696 1.8506999999999998e-08 1.841092826571469 1.8508e-08 1.7593847066698864 1.8509e-08 1.7655464773358356 1.8509999999999998e-08 1.8425102477845359 1.8511e-08 1.8056542309916022 1.8512e-08 1.7539179183742117 1.8513e-08 1.794186721166985 1.8514e-08 1.9284025450399327 1.8515e-08 1.7779554772460873 1.8516e-08 1.8434757715401437 1.8517e-08 1.792632927234495 1.8518e-08 1.7628928189835804 1.8519e-08 1.8292833752183517 1.852e-08 1.7196664217555655 1.8521e-08 1.7435440666158677 1.8522e-08 1.8037215776426698 1.8523e-08 1.8034947403689803 1.8524e-08 1.7421886743415265 1.8525e-08 1.763177221340496 1.8526e-08 1.8133231534728211 1.8527e-08 1.872639148502378 1.8528e-08 1.8089832707310824 1.8529e-08 1.7871914232629869 1.853e-08 1.8333944340054038 1.8531e-08 1.8026937535881 1.8532e-08 1.8188667703178691 1.8533e-08 1.7356660524460756 1.8534e-08 1.7289903384617225 1.8535e-08 1.7563040130883274 1.8535999999999998e-08 1.8488578316485005 1.8537e-08 1.7386849789743228 1.8538e-08 1.7646646647531397 1.8538999999999998e-08 1.8847943039947914 1.854e-08 1.73497064355632 1.8541e-08 1.735755240431647 1.8541999999999998e-08 1.7325636862730398 1.8543e-08 1.7819421070380406 1.8544e-08 1.7787795617568471 1.8544999999999998e-08 1.7461087142149025 1.8546e-08 1.7505787112989477 1.8547e-08 1.8411214973832555 1.8548e-08 1.7602470273304085 1.8549e-08 1.8331455504760032 1.855e-08 1.7638531095472525 1.8551e-08 1.6796059345216663 1.8552e-08 1.8377083801258174 1.8553e-08 1.7957559381842743 1.8554e-08 1.8248969855620947 1.8555e-08 1.7729725221934847 1.8556e-08 1.7420289465102725 1.8557e-08 1.8520007206790046 1.8558e-08 1.8519936308379592 1.8559e-08 1.7777949263855106 1.856e-08 1.8044721868156548 1.8561e-08 1.7430784893786524 1.8562e-08 1.8409099864112357 1.8563e-08 1.8234934529301898 1.8564e-08 1.6825023110613697 1.8565e-08 1.833203867703785 1.8566e-08 1.8488325462586128 1.8567e-08 1.8230928732754403 1.8568e-08 1.7834234708275367 1.8569e-08 1.8164251055156273 1.857e-08 1.8457558472374043 1.8570999999999998e-08 1.8620390628089756 1.8572e-08 1.8136093530261543 1.8573e-08 1.8080120646902567 1.8573999999999998e-08 1.8000049134085416 1.8575e-08 1.8190764212472725 1.8576e-08 1.7160061655282637 1.8576999999999998e-08 1.7009034316833596 1.8578e-08 1.7355897805636955 1.8579e-08 1.8112036705041905 1.8579999999999998e-08 1.7522056873695033 1.8581e-08 1.853980792500818 1.8582e-08 1.7388108871245709 1.8583e-08 1.8173855869309579 1.8584e-08 1.81933073440269 1.8585e-08 1.7483599293130454 1.8586e-08 1.8013169809608778 1.8587e-08 1.8859327395500125 1.8588e-08 1.8909200766930157 1.8589e-08 1.7164367024736038 1.859e-08 1.8064593967149656 1.8591e-08 1.7780331379890144 1.8592e-08 1.7669345827339207 1.8593e-08 1.8316282230171002 1.8594e-08 1.813843597939549 1.8595e-08 1.8192306767145112 1.8596e-08 1.750281125884345 1.8597e-08 1.8541151666300606 1.8598e-08 1.9137271763742134 1.8599e-08 1.852387127420843 1.86e-08 1.7876086881765425 1.8601e-08 1.80010265326595 1.8602e-08 1.7517831253222695 1.8603e-08 1.7576374355879616 1.8604e-08 1.8446769223667614 1.8605e-08 1.7405123738654666 1.8605999999999998e-08 1.838349885818754 1.8607e-08 1.8741498032727755 1.8608e-08 1.8755345359220488 1.8608999999999998e-08 1.7559577409122653 1.861e-08 1.8284165049449206 1.8611e-08 1.782113252734603 1.8611999999999998e-08 1.7035959159224463 1.8613e-08 1.7473411735150268 1.8614e-08 1.6981599795003102 1.8614999999999998e-08 1.8914900534979366 1.8616e-08 1.8694491898852936 1.8617e-08 1.7889861301314922 1.8618e-08 1.7368166651062587 1.8619e-08 1.7428402813936705 1.862e-08 1.7596386529477346 1.8621e-08 1.9786429296960415 1.8622e-08 1.7903231918012257 1.8623e-08 1.7755012427179067 1.8624e-08 1.84097594272927 1.8625e-08 1.7440219135043895 1.8626e-08 1.747896481129368 1.8627e-08 1.7814272606143646 1.8628e-08 1.8409656141973596 1.8629e-08 1.8530173408199548 1.863e-08 1.7962362818409379 1.8631e-08 1.7926354945834333 1.8632e-08 1.7389826705914 1.8633e-08 1.8679995425828557 1.8634e-08 1.7787984497164022 1.8635e-08 1.8520921505282812 1.8636e-08 1.8079650418964723 1.8637e-08 1.7570922726164409 1.8638e-08 1.7033212061729808 1.8639e-08 1.8220003879344049 1.864e-08 1.7715406985965845 1.8640999999999998e-08 1.7698572487160373 1.8642e-08 1.8584262960290865 1.8643e-08 1.8005099429247386 1.8643999999999998e-08 1.80675203786257 1.8645e-08 1.8412043784161511 1.8646e-08 1.8078959375821109 1.8646999999999998e-08 1.7160523248076183 1.8648e-08 1.8560130010803375 1.8649e-08 1.8130607851740075 1.8649999999999998e-08 1.8704888154071506 1.8651e-08 1.8317844140220239 1.8652e-08 1.7237323837330736 1.8653e-08 1.7744816288968555 1.8654e-08 1.8696722002358628 1.8655e-08 1.8698310184323916 1.8656e-08 1.7974256477158366 1.8657e-08 1.7628433814667837 1.8658e-08 1.7650883047224608 1.8659e-08 1.8096881932250768 1.866e-08 1.7747261959009204 1.8661e-08 1.8672197974300477 1.8662e-08 1.7750386205608355 1.8663e-08 1.8247116230819376 1.8664e-08 1.757724393870667 1.8665e-08 1.8777100436793956 1.8666e-08 1.8567567935651093 1.8667e-08 1.7652918802030229 1.8668e-08 1.8053371488399224 1.8669e-08 1.7904917353523528 1.867e-08 1.7548025612924878 1.8671e-08 1.8511669529321502 1.8672e-08 1.8652182518996918 1.8673e-08 1.9058872645874079 1.8674e-08 1.816676515835275 1.8675e-08 1.799692456612045 1.8676e-08 1.8616974435220743 1.8677e-08 1.804731401802397 1.8678e-08 1.847762773081577 1.8678999999999998e-08 1.7690457175682464 1.868e-08 1.8463591414286347 1.8681e-08 1.8312778784831736 1.8681999999999998e-08 1.8802441113339456 1.8683e-08 1.7536927683644636 1.8684e-08 1.8033311998401855 1.8684999999999998e-08 1.8160759138304452 1.8686e-08 1.7842406978310497 1.8687e-08 1.8832219310811307 1.8687999999999998e-08 1.7954672981748434 1.8689e-08 1.8450104352161731 1.869e-08 1.8319570746881186 1.8691e-08 1.7520993158770435 1.8692e-08 1.8179248050698718 1.8693e-08 1.7500815775349843 1.8694e-08 1.7810730791879852 1.8695e-08 1.806343660641677 1.8696e-08 1.812170241755821 1.8697e-08 1.844126494614628 1.8698e-08 1.8174683305634665 1.8699e-08 1.7733561440110235 1.87e-08 1.851933930365401 1.8701e-08 1.7981968694077761 1.8702e-08 1.7542129631443537 1.8703e-08 1.771099860340292 1.8704e-08 1.8594781257217177 1.8705e-08 1.8143448257339871 1.8706e-08 1.9012158132741543 1.8707e-08 1.7912417247623211 1.8708e-08 1.7700517063601373 1.8709e-08 1.8264726771106932 1.871e-08 1.893742073290415 1.8711e-08 1.7570380515348976 1.8712e-08 1.7585397807662808 1.8713e-08 1.8437051347224305 1.8713999999999998e-08 1.7546126256431682 1.8715e-08 1.8208707242859896 1.8716e-08 1.849033619725337 1.8716999999999998e-08 1.7810155089421897 1.8718e-08 1.7503809196224493 1.8719e-08 1.8598602172276366 1.8719999999999998e-08 1.8712339499093118 1.8721e-08 1.8073347055264704 1.8722e-08 1.8007030255787058 1.8722999999999998e-08 1.806189734985917 1.8724e-08 1.8441519560339712 1.8725e-08 1.788228989440004 1.8726e-08 1.7508403766602665 1.8727e-08 1.8475746593619042 1.8728e-08 1.763366897257698 1.8729e-08 1.7762251906406035 1.873e-08 1.7550135056315508 1.8731e-08 1.8643184448774754 1.8732e-08 1.8311384900282792 1.8733e-08 1.714212262942278 1.8734e-08 1.8084671567745019 1.8735e-08 1.7882638446032924 1.8736e-08 1.7985252604311452 1.8737e-08 1.8159755204331944 1.8738e-08 1.742842863449525 1.8739e-08 1.8099931691144409 1.874e-08 1.8102901306235317 1.8741e-08 1.8902927892353767 1.8742e-08 1.8930864118388242 1.8743e-08 1.82059742175872 1.8744e-08 1.7384812664122136 1.8745e-08 1.7391106201263375 1.8746e-08 1.7420401542065453 1.8747e-08 1.877601668416969 1.8748e-08 1.7273282555068816 1.8748999999999998e-08 1.8291945864670653 1.875e-08 1.832204996834057 1.8751e-08 1.7503693038195034 1.8751999999999998e-08 1.8058296173673143 1.8753e-08 1.7252380728179901 1.8754e-08 1.8375825784978763 1.8754999999999998e-08 1.8198427936532873 1.8756e-08 1.8471814247140992 1.8757e-08 1.8435659538748645 1.8757999999999998e-08 1.8450002655579787 1.8759e-08 1.7913947016795493 1.876e-08 1.8072817338896434 1.8761e-08 1.786731827537392 1.8762e-08 1.8260148525509388 1.8763e-08 1.8903492588892061 1.8764e-08 1.7967142259279152 1.8765e-08 1.7442876746642748 1.8766e-08 1.8078613283132965 1.8767e-08 1.7458193956886499 1.8768e-08 1.833823603226621 1.8769e-08 1.7283991712501727 1.877e-08 1.784210581188798 1.8771e-08 1.7980280076895367 1.8772e-08 1.9045576710056773 1.8773e-08 1.8031990392006643 1.8774e-08 1.8799201718493546 1.8775e-08 1.7885699851128327 1.8776e-08 1.8065202421924467 1.8777e-08 1.7627092550712282 1.8778e-08 1.7385768050276116 1.8779e-08 1.8183305673995112 1.878e-08 1.8251802927541532 1.8781e-08 1.810000792096952 1.8782e-08 1.710252660367496 1.8783e-08 1.7205454248196468 1.8783999999999998e-08 1.808424811321972 1.8785e-08 1.756973251138607 1.8786e-08 1.7670208428146168 1.8786999999999998e-08 1.82146839903258 1.8788e-08 1.7830117618433652 1.8789e-08 1.7439720501657516 1.8789999999999998e-08 1.8504965248842966 1.8791e-08 1.687231311640969 1.8792e-08 1.783841670463182 1.8792999999999998e-08 1.7507011822815097 1.8794e-08 1.8343131571572273 1.8795e-08 1.8487786560445727 1.8796e-08 1.8722934157729696 1.8797e-08 1.767856578827478 1.8798e-08 1.8436319334175784 1.8799e-08 1.7635487582692164 1.88e-08 1.7623082565179016 1.8801e-08 1.7743730518621406 1.8802e-08 1.7742022648454125 1.8803e-08 1.7372214546513287 1.8804e-08 1.8314729261699552 1.8805e-08 1.7740491791069362 1.8806e-08 1.8333474492575477 1.8807e-08 1.790595897953501 1.8808e-08 1.82095842595315 1.8809e-08 1.9198675644717655 1.881e-08 1.8424205082769907 1.8811e-08 1.8455875594947189 1.8812e-08 1.8009694756926402 1.8813e-08 1.8049347704594765 1.8814e-08 1.8182837518547323 1.8815e-08 1.8282786772935642 1.8816e-08 1.7520701926578786 1.8817e-08 1.807037992997774 1.8818e-08 1.7961979610903775 1.8818999999999998e-08 1.773522211214042 1.882e-08 1.8675632968594658 1.8821e-08 1.8296979915503888 1.8821999999999998e-08 1.866989395361389 1.8823e-08 1.8113279651538703 1.8824e-08 1.6521248205105024 1.8824999999999998e-08 2.0146312074473336 1.8826e-08 1.767488262515789 1.8827e-08 1.752923161475004 1.8827999999999998e-08 1.948333418342547 1.8829e-08 1.8683871696681662 1.883e-08 1.8689163069479466 1.8831e-08 1.7464917414394538 1.8832e-08 1.7013048277320169 1.8833e-08 1.7927785780769456 1.8834e-08 1.73791292648382 1.8835e-08 1.7899894142220572 1.8836e-08 1.799949423549666 1.8837e-08 1.7561912478926613 1.8838e-08 1.7621073889819103 1.8839e-08 1.853614032106964 1.884e-08 1.8141548222211366 1.8841e-08 1.869207590844679 1.8842e-08 1.8500961061422996 1.8843e-08 1.741635745987673 1.8844e-08 1.8986677508578822 1.8845e-08 1.7942047757589354 1.8846e-08 1.818579594198808 1.8847e-08 1.934352061344804 1.8848e-08 1.7067090255029749 1.8849e-08 1.7847287345778995 1.885e-08 1.833866295056321 1.8851e-08 1.7573546213296922 1.8852e-08 1.788364010593924 1.8853e-08 1.797398108815984 1.8854e-08 1.8467420701115989 1.8855e-08 1.6860770461316223 1.8856e-08 1.7022052815838313 1.8856999999999998e-08 1.8121872081255153 1.8858e-08 1.7620169242520962 1.8859e-08 1.8405847848682035 1.8859999999999998e-08 1.6708124502251904 1.8861e-08 1.8235997566706228 1.8862e-08 1.6779061867906926 1.8862999999999998e-08 1.7108880757354328 1.8864e-08 1.7865175595793863 1.8865e-08 1.7206082595025625 1.8865999999999998e-08 1.8116985992500634 1.8867e-08 1.6907913813557882 1.8868e-08 1.8351716971253018 1.8869e-08 1.7137083044877444 1.887e-08 1.781887071320782 1.8871e-08 1.8086188561128453 1.8872e-08 1.815297270706461 1.8873e-08 1.7694017744836423 1.8874e-08 1.7428228433110122 1.8875e-08 1.8478283926974017 1.8876e-08 1.8003092712366948 1.8877e-08 1.7493218241267292 1.8878e-08 1.7051401842860645 1.8879e-08 1.803208699841219 1.888e-08 1.7255296418138155 1.8881e-08 1.7548054555280788 1.8882e-08 1.7958537199538442 1.8883e-08 1.8651675606823788 1.8884e-08 1.782018923995014 1.8885e-08 1.8344678409827522 1.8886e-08 1.861499425460839 1.8887e-08 1.8066042859014246 1.8888e-08 1.8122187702300887 1.8889e-08 1.7933483416429774 1.889e-08 1.7106372011189865 1.8891e-08 1.7121347320677316 1.8891999999999998e-08 1.8267325517759943 1.8893e-08 1.7227302885602493 1.8894e-08 1.7518068116563965 1.8894999999999998e-08 1.8911770892739197 1.8896e-08 1.9247554322735505 1.8897e-08 1.8440207729779525 1.8897999999999998e-08 1.7735273426240368 1.8899e-08 1.9247785786038527 1.89e-08 1.801968455419725 1.8900999999999998e-08 1.8418009352921656 1.8902e-08 1.8474440084743406 1.8903e-08 1.8132851553787366 1.8904e-08 1.7892514187523552 1.8905e-08 1.9151267719642973 1.8906e-08 1.8178867551663218 1.8907e-08 1.8224201930375237 1.8908e-08 1.7378559889046412 1.8909e-08 1.7961201766835446 1.891e-08 1.8300495468047917 1.8911e-08 1.841101504260976 1.8912e-08 1.876410501228178 1.8913e-08 1.8034267735439313 1.8914e-08 1.8199131876294552 1.8915e-08 1.7494700499395954 1.8916e-08 1.7138147016031742 1.8917e-08 1.8060479492433774 1.8918e-08 1.8541178536017766 1.8919e-08 1.8401520930803608 1.892e-08 1.8202787246068874 1.8921e-08 1.8292109724555994 1.8922e-08 1.7999320105893977 1.8923e-08 1.8009456803634183 1.8924e-08 1.7916408609248273 1.8925e-08 1.851908704812553 1.8926e-08 1.846906944866545 1.8926999999999998e-08 1.7772644638835398 1.8928e-08 1.6936913630529264 1.8929e-08 1.75362000363729 1.8929999999999998e-08 1.7015145927408921 1.8931e-08 1.7742730703184764 1.8932e-08 1.9042919477403788 1.8932999999999998e-08 1.780864618732128 1.8934e-08 1.8194575758445626 1.8935e-08 1.812162305591079 1.8935999999999998e-08 1.8968976552732484 1.8937e-08 1.7656962199702546 1.8938e-08 1.8548710159197606 1.8939e-08 1.7485472591572597 1.894e-08 1.7958096594984518 1.8941e-08 1.864069006923654 1.8942e-08 1.7642661001167845 1.8943e-08 1.7524995932032272 1.8944e-08 1.8502246518095273 1.8945e-08 1.8817769883926376 1.8946e-08 1.7337277276525938 1.8947e-08 1.7830583831909836 1.8948e-08 1.8255882389920421 1.8949e-08 1.7908382877883553 1.895e-08 1.7794600968474252 1.8951e-08 1.8254424541976 1.8952e-08 1.8349941896837205 1.8953e-08 1.781607136539574 1.8954e-08 1.7561039381371617 1.8955e-08 1.8299642647295131 1.8956e-08 1.8306337359977962 1.8957e-08 1.8682895035260438 1.8958e-08 1.6838119749247649 1.8959e-08 1.8398584197611647 1.896e-08 1.8025525448700677 1.8961e-08 1.811233190847674 1.8961999999999998e-08 1.8254613405526365 1.8963e-08 1.764932519753212 1.8964e-08 1.8538510800217374 1.8964999999999998e-08 1.7390706535110019 1.8966e-08 1.7556349753647038 1.8967e-08 1.6962415602036658 1.8967999999999998e-08 1.7962134572650243 1.8969e-08 1.8832025500820508 1.897e-08 1.8549285846150463 1.8970999999999998e-08 1.7824046163887008 1.8972e-08 1.8699449938796304 1.8973e-08 1.8217926432514484 1.8974e-08 1.861666176757351 1.8975e-08 1.759666528409029 1.8976e-08 1.7787203367965823 1.8977e-08 1.8153566739965818 1.8978e-08 1.8013020176347199 1.8979e-08 1.812213713956727 1.898e-08 1.7296265634600736 1.8981e-08 1.8620379022658835 1.8982e-08 1.713181238520938 1.8983e-08 1.802818102990793 1.8984e-08 1.8268386207611222 1.8985e-08 1.849487736008399 1.8986e-08 1.7958775812502064 1.8987e-08 1.8134608246696093 1.8988e-08 1.876356930336124 1.8989e-08 1.871204186458852 1.899e-08 1.8694208877900407 1.8991e-08 1.8037130466958282 1.8992e-08 1.8295082090656318 1.8993e-08 1.7508471121137026 1.8994e-08 1.8313939681427194 1.8995e-08 1.898742819248341 1.8996e-08 1.8050425728943003 1.8996999999999998e-08 1.7822844118141292 1.8998e-08 1.8528622988340808 1.8999e-08 1.8822982587976684 1.8999999999999998e-08 1.7377397901417715 1.9001e-08 1.7796950601430792 1.9002e-08 1.8670690964451808 1.9002999999999998e-08 1.7817436650676037 1.9004e-08 1.8663739298927549 1.9005e-08 1.7995384034826882 1.9005999999999998e-08 1.7636609113405068 1.9007e-08 1.8065982098556626 1.9008e-08 1.7828632537326847 1.9009e-08 1.7618771427570357 1.901e-08 1.8632111692767872 1.9011e-08 1.8362583048269996 1.9012e-08 1.7885310559190755 1.9013e-08 1.805031783521073 1.9014e-08 1.8881009780695286 1.9015e-08 1.8764510621053483 1.9016e-08 1.778712906000589 1.9017e-08 1.8906948999890378 1.9018e-08 1.8842124950359764 1.9019e-08 1.7827353597942215 1.902e-08 1.677569549219421 1.9021e-08 1.9048748114077823 1.9022e-08 1.8692416508721292 1.9023e-08 1.8016990854217416 1.9024e-08 1.8401783464200288 1.9025e-08 1.7711059559232663 1.9026e-08 1.8249270145199388 1.9027e-08 1.6797571515848664 1.9028e-08 1.8105980154194807 1.9029e-08 1.7425562134664039 1.903e-08 1.7611442437995375 1.9031e-08 1.718656122694504 1.9031999999999998e-08 1.7174151696204707 1.9033e-08 1.7739323425916822 1.9034e-08 1.789299612887453 1.9034999999999998e-08 1.8468410842851335 1.9036e-08 1.8237913695893286 1.9037e-08 1.781892277881045 1.9037999999999998e-08 1.8847099781781362 1.9039e-08 1.6928314063026928 1.904e-08 1.8720897065174695 1.9040999999999998e-08 1.8495616159716874 1.9042e-08 1.7516519384732832 1.9043e-08 1.7803025648222341 1.9043999999999998e-08 1.8175109604583255 1.9045e-08 1.7379385334499833 1.9046e-08 1.824315075977712 1.9047e-08 1.7155542619138269 1.9048e-08 1.711461864027312 1.9049e-08 1.821285359314249 1.905e-08 1.8519798744802825 1.9051e-08 1.7985260992231367 1.9052e-08 1.8272973424589867 1.9053e-08 1.79484996666593 1.9054e-08 1.736685458912116 1.9055e-08 1.8436935092951383 1.9056e-08 1.7895874264271177 1.9057e-08 1.7765077612270541 1.9058e-08 1.832460210985947 1.9059e-08 1.829871203687787 1.906e-08 1.89973413946992 1.9061e-08 1.833131884446442 1.9062e-08 1.916471056161326 1.9063e-08 1.8658551263751684 1.9064e-08 1.823307513086899 1.9065e-08 1.8073359227544377 1.9066e-08 1.745359515991062 1.9067e-08 1.8166318287080192 1.9068e-08 1.8245878111940124 1.9069e-08 1.7983339645439103 1.9069999999999998e-08 1.8627130470932505 1.9071e-08 1.7679051063954758 1.9072e-08 1.8135080307063423 1.9072999999999998e-08 1.7465379707098256 1.9074e-08 1.8314688024767656 1.9075e-08 1.7205828357954478 1.9075999999999998e-08 1.7808335836027955 1.9077e-08 1.8010009201787511 1.9078e-08 1.690525615454364 1.9078999999999998e-08 1.7775892043542862 1.908e-08 1.8757848487027018 1.9081e-08 1.8267460157825381 1.9082e-08 1.7409825802460712 1.9083e-08 1.7886626561299943 1.9084e-08 1.8631880584973763 1.9085e-08 1.7545040606715765 1.9086e-08 1.8488255529952051 1.9087e-08 1.8015743847385153 1.9088e-08 1.9026824559709956 1.9089e-08 1.8105594548342414 1.909e-08 1.8403703895042032 1.9091e-08 1.859692275075071 1.9092e-08 1.7382888684715379 1.9093e-08 1.7145744043528859 1.9094e-08 1.8707717516430875 1.9095e-08 1.8308654401409001 1.9096e-08 1.801089167842981 1.9097e-08 1.6963588033308599 1.9098e-08 1.8112848814991196 1.9099e-08 1.7689222793319794 1.91e-08 1.7434921050782515 1.9101e-08 1.9024211533639077 1.9102e-08 1.8216975508671216 1.9103e-08 1.7892098188986556 1.9104e-08 1.8461931249251384 1.9104999999999998e-08 1.7726211193626455 1.9106e-08 1.8397455319520695 1.9107e-08 1.7995572873536254 1.9107999999999998e-08 1.757334153592969 1.9109e-08 1.8407588222040236 1.911e-08 1.8714457279336467 1.9110999999999998e-08 1.820854525026201 1.9112e-08 1.8249555489900768 1.9113e-08 1.8017077777625559 1.9113999999999998e-08 1.7450575178349401 1.9115e-08 1.787979936672919 1.9116e-08 1.8061832253457413 1.9117e-08 1.9001426095912364 1.9118e-08 1.8220321647345 1.9119e-08 1.7659809666182433 1.912e-08 1.7214102235011748 1.9121e-08 1.801790309781888 1.9122e-08 1.829647778522835 1.9123e-08 1.79891294714464 1.9124e-08 1.7921596841235579 1.9125e-08 1.7932562193311712 1.9126e-08 1.7254792998295925 1.9127e-08 1.7903439799889282 1.9128e-08 1.8281530073502141 1.9129e-08 1.8203054177544615 1.913e-08 1.7915016403420805 1.9131e-08 1.801369414958842 1.9132e-08 1.7871437441755456 1.9133e-08 1.7715284357161338 1.9134e-08 1.9194845366810533 1.9135e-08 1.7490382008128846 1.9136e-08 1.6902488518864662 1.9137e-08 1.7961745693482285 1.9138e-08 1.8443363402407602 1.9139e-08 1.8043380355291772 1.9139999999999998e-08 1.8521964829221118 1.9141e-08 1.8837230190366496 1.9142e-08 1.7406352980927196 1.9142999999999998e-08 1.733291962386297 1.9144e-08 1.7967118033631972 1.9145e-08 1.8519781421010886 1.9145999999999998e-08 1.767455963050968 1.9147e-08 1.8589064257157493 1.9148e-08 1.7819716241795127 1.9148999999999998e-08 1.765310184479053 1.915e-08 1.7990316712124312 1.9151e-08 1.8192745696877393 1.9152e-08 1.8011864484735076 1.9153e-08 1.764253685945887 1.9154e-08 1.8256054077255124 1.9155e-08 1.720155800813041 1.9156e-08 1.805648605005258 1.9157e-08 1.6855961456657824 1.9158e-08 1.758042954073139 1.9159e-08 1.8483298685957297 1.916e-08 1.8289839194413209 1.9161e-08 1.7219175303094327 1.9162e-08 1.6791462573606035 1.9163e-08 1.766605209642621 1.9164e-08 1.7642369788937278 1.9165e-08 1.675362828041891 1.9166e-08 1.8267355312296472 1.9167e-08 1.8439107806625528 1.9168e-08 1.7545325620190488 1.9169e-08 1.769357583986704 1.917e-08 1.8237535763585104 1.9171e-08 1.7185655187237232 1.9172e-08 1.88444780411285 1.9173e-08 1.7981995049746307 1.9174e-08 1.7814027364866352 1.9174999999999998e-08 1.7634030271800512 1.9176e-08 1.8321500254573546 1.9177e-08 1.7057519007525375 1.9177999999999998e-08 1.8242864192362014 1.9179e-08 1.7079502177904153 1.918e-08 1.7460944206020834 1.9180999999999998e-08 1.7890284144307673 1.9182e-08 1.8268751451536032 1.9183e-08 1.8618047699330975 1.9183999999999998e-08 1.830830776133154 1.9185e-08 1.8381219510442353 1.9186e-08 1.7918831755945905 1.9187e-08 1.7678253166621791 1.9188e-08 1.7473680345831404 1.9189e-08 1.8490257265903967 1.919e-08 1.6825799900223903 1.9191e-08 1.8435659705686351 1.9192e-08 1.8262297867965858 1.9193e-08 1.6794838815030972 1.9194e-08 1.8919657334776432 1.9195e-08 1.8390599556315737 1.9196e-08 1.828691548966459 1.9197e-08 1.7203553142527075 1.9198e-08 1.7428147060569699 1.9199e-08 1.6993489014567102 1.92e-08 1.8322172859523407 1.9201e-08 1.8232589237066474 1.9202e-08 1.7054944174356268 1.9203e-08 1.679140814318883 1.9204e-08 1.772464345836048 1.9205e-08 1.842042755737879 1.9206e-08 1.7674997795284753 1.9207e-08 1.8511582967915157 1.9208e-08 1.7945825419216521 1.9209e-08 1.7263089987375635 1.9209999999999998e-08 1.8551867654167964 1.9211e-08 1.7877181424828559 1.9212e-08 1.7240957416560303 1.9212999999999998e-08 1.8955342208976682 1.9214e-08 1.8628572303653823 1.9215e-08 1.88649309399095 1.9215999999999998e-08 1.8916836608636143 1.9217e-08 1.8513141415228551 1.9218e-08 1.7862296461432408 1.9218999999999998e-08 1.8204314639905486 1.922e-08 1.769249146224122 1.9221e-08 1.722203790556469 1.9222e-08 1.7336030419688166 1.9223e-08 1.7727339704092209 1.9224e-08 1.8218088289646093 1.9225e-08 1.7427953102061953 1.9226e-08 1.8213944190360771 1.9227e-08 1.8350185843965097 1.9228e-08 1.7341256441554218 1.9229e-08 1.8427130205798006 1.923e-08 1.725275866952822 1.9231e-08 1.7761438604416309 1.9232e-08 1.8165304863268366 1.9233e-08 1.6928242714660966 1.9234e-08 1.8876310152833937 1.9235e-08 1.8250232747752584 1.9236e-08 1.7940466996344469 1.9237e-08 1.7843952326468715 1.9238e-08 1.8258463546588315 1.9239e-08 1.8590727607439377 1.924e-08 1.8070538824771822 1.9241e-08 1.7430616361153268 1.9242e-08 1.8115926689212112 1.9243e-08 1.743816377882334 1.9244e-08 1.838747636158069 1.9244999999999998e-08 1.8649529669414 1.9246e-08 1.8395233194762708 1.9247e-08 1.691810068141242 1.9247999999999998e-08 1.812423600005191 1.9249e-08 1.7144212703559256 1.925e-08 1.803493520554151 1.9250999999999998e-08 1.8152848618126576 1.9252e-08 1.7438173455825798 1.9253e-08 1.7521033975289333 1.9253999999999998e-08 1.81034645847627 1.9255e-08 1.7925507733228276 1.9256e-08 1.7636799715283153 1.9256999999999998e-08 1.7793190521298508 1.9258e-08 1.7449788053346968 1.9259e-08 1.7995768434459338 1.926e-08 1.8771501410837332 1.9261e-08 1.7902813949154903 1.9262e-08 1.7968531939899628 1.9263e-08 1.7163689202838377 1.9264e-08 1.793988297889141 1.9265e-08 1.752453901856853 1.9266e-08 1.822946301707312 1.9267e-08 1.7418680401675126 1.9268e-08 1.8260653658003454 1.9269e-08 1.8664639545014003 1.927e-08 1.7560111498368869 1.9271e-08 1.7131727420392622 1.9272e-08 1.840247576946731 1.9273e-08 1.7420983921015014 1.9274e-08 1.7589701373547935 1.9275e-08 1.8846869155112251 1.9276e-08 1.8019867171776849 1.9277e-08 1.8077989860531711 1.9278e-08 1.8561602671554864 1.9279e-08 1.6847610430995916 1.928e-08 1.7941542891542388 1.9281e-08 1.7058421850236767 1.9282e-08 1.8480841111533681 1.9282999999999998e-08 1.7004791052537938 1.9284e-08 1.865103234346905 1.9285e-08 1.8427152183291173 1.9285999999999998e-08 1.8474070190280094 1.9287e-08 1.847060943319174 1.9288e-08 1.8036453448123426 1.9288999999999998e-08 1.7100813429026838 1.929e-08 1.804160995293363 1.9291e-08 1.722219918234325 1.9291999999999998e-08 1.8173697771934043 1.9293e-08 1.774197455219585 1.9294e-08 1.8139986934003716 1.9295e-08 1.828612284018073 1.9296e-08 1.7841631975036572 1.9297e-08 1.8058513381491283 1.9298e-08 1.7883388921413517 1.9299e-08 1.825949718203778 1.93e-08 1.7877788524177327 1.9301e-08 1.8330000313291532 1.9302e-08 1.8311880893625734 1.9303e-08 1.7961745552822947 1.9304e-08 1.8945841846022915 1.9305e-08 1.7910682411381051 1.9306e-08 1.7741151588224815 1.9307e-08 1.7688360883912007 1.9308e-08 1.7750050208215125 1.9309e-08 1.760055561663394 1.931e-08 1.7806400032320084 1.9311e-08 1.718305438029704 1.9312e-08 1.7954911593179856 1.9313e-08 1.8368556983988342 1.9314e-08 1.747706165163248 1.9315e-08 1.7952700764139524 1.9316e-08 1.7491118610222158 1.9317e-08 1.8362622848719334 1.9317999999999998e-08 1.8264027228374544 1.9319e-08 1.7590923369200075 1.932e-08 1.741535453649739 1.9320999999999998e-08 1.8507012325845484 1.9322e-08 1.8967218247443283 1.9323e-08 1.7561075071186225 1.9323999999999998e-08 1.8533648758549324 1.9325e-08 1.8122035121106124 1.9326e-08 1.7589133026093675 1.9326999999999998e-08 1.7608757113758198 1.9328e-08 1.8602050126645393 1.9329e-08 1.786652942653349 1.933e-08 1.8532264601853634 1.9331e-08 1.782991241303845 1.9332e-08 1.8192603515942727 1.9333e-08 1.72524762412887 1.9334e-08 1.7672050919684634 1.9335e-08 1.7548276695324543 1.9336e-08 1.8355529078401631 1.9337e-08 1.7918426344917846 1.9338e-08 1.7851435201642016 1.9339e-08 1.7114424668414865 1.934e-08 1.8121157448746483 1.9341e-08 1.6883823742318826 1.9342e-08 1.780236939184737 1.9343e-08 1.7962802675125618 1.9344e-08 1.8214261193989894 1.9345e-08 1.8961728489557261 1.9346e-08 1.8136530996654912 1.9347e-08 1.8171045604023697 1.9348e-08 1.7533373481172034 1.9349e-08 1.7581956199649778 1.935e-08 1.8135312923974396 1.9351e-08 1.8357447644498774 1.9352e-08 1.8296570426646805 1.9352999999999998e-08 1.7916751871529049 1.9354e-08 1.7965963591192804 1.9355e-08 1.8280053723183822 1.9355999999999998e-08 1.7877494621843146 1.9357e-08 1.8412864760293384 1.9358e-08 1.8342805984696888 1.9358999999999998e-08 1.7707386064163997 1.936e-08 1.8663224785849828 1.9361e-08 1.7318342286866526 1.9361999999999998e-08 1.7719661873190633 1.9363e-08 1.7712891663439065 1.9364e-08 1.7629633461659728 1.9365e-08 1.8328611224870586 1.9366e-08 1.757986437533105 1.9367e-08 1.7716615061648273 1.9368e-08 1.7442645771803205 1.9369e-08 1.8018593853772353 1.937e-08 1.8175773022257575 1.9371e-08 1.7371949961550865 1.9372e-08 1.812137709213418 1.9373e-08 1.8444373865695516 1.9374e-08 1.7241375278060773 1.9375e-08 1.7999399057731613 1.9376e-08 1.82797107359004 1.9377e-08 1.8177698969371472 1.9378e-08 1.7865287645737948 1.9379e-08 1.8470873574654125 1.938e-08 1.799780961669641 1.9381e-08 1.7889218667814923 1.9382e-08 1.821278109470449 1.9383e-08 1.7704886174464367 1.9384e-08 1.7903327202997614 1.9385e-08 1.817774490981573 1.9386e-08 1.712554577449651 1.9387e-08 1.7456492915496373 1.9387999999999998e-08 1.9033567307184691 1.9389e-08 1.7721593777601796 1.939e-08 1.9063785790945627 1.9390999999999998e-08 1.8283402452514854 1.9392e-08 1.8239764884890506 1.9393e-08 1.7647473747729805 1.9393999999999998e-08 1.7388666910856174 1.9395e-08 1.8056206280549396 1.9396e-08 1.7986008251932704 1.9396999999999998e-08 1.774270167918519 1.9398e-08 1.8194466150701802 1.9399e-08 1.782746266627527 1.94e-08 1.741859694116393 1.9401e-08 1.8578636144166751 1.9402e-08 1.7535188669655932 1.9403e-08 1.7920697970584838 1.9404e-08 1.6773201671962932 1.9405e-08 1.7898122202127782 1.9406e-08 1.8609327836828689 1.9407e-08 1.8691219098239025 1.9408e-08 1.8600845675946656 1.9409e-08 1.90300893606763 1.941e-08 1.6924417076782525 1.9411e-08 1.7671147810703243 1.9412e-08 1.8044059780049213 1.9413e-08 1.8691544934628161 1.9414e-08 1.7830559495689111 1.9415e-08 1.8498650517218298 1.9416e-08 1.8346257049969312 1.9417e-08 1.7880047666548593 1.9418e-08 1.784970722853976 1.9419e-08 1.681629556881841 1.942e-08 1.7916640640841313 1.9421e-08 1.7562051591008474 1.9422e-08 1.823833933401523 1.9422999999999998e-08 1.8540954866046981 1.9424e-08 1.7321021493587008 1.9425e-08 1.7369189673757215 1.9425999999999998e-08 1.8697559057976856 1.9427e-08 1.7885896728686677 1.9428e-08 1.8152635853166779 1.9428999999999998e-08 1.77822428339124 1.943e-08 1.8160000376858623 1.9431e-08 1.858442477734769 1.9431999999999998e-08 1.780885601045557 1.9433e-08 1.903100692459446 1.9434e-08 1.817145917839146 1.9434999999999998e-08 1.787462787088533 1.9436e-08 1.7316270802168099 1.9437e-08 1.835223384709974 1.9438e-08 1.9652235646109348 1.9439e-08 1.7732496184510875 1.944e-08 1.8119826443287719 1.9441e-08 1.7453081015887921 1.9442e-08 1.8101678558904515 1.9443e-08 1.6947090388932875 1.9444e-08 1.7542251052784692 1.9445e-08 1.8281227344591653 1.9446e-08 1.7918726424347542 1.9447e-08 1.8368105823211054 1.9448e-08 1.7458410361109145 1.9449e-08 1.7095941589980144 1.945e-08 1.8765556620990014 1.9451e-08 1.8176633346189643 1.9452e-08 1.7593106026659884 1.9453e-08 1.8513445888461069 1.9454e-08 1.7822522314398106 1.9455e-08 1.6690623720998405 1.9456e-08 1.8356844620442736 1.9457e-08 1.7140553848908624 1.9458e-08 1.7969639227688168 1.9459e-08 1.8468689256777244 1.946e-08 1.7804045164917726 1.9460999999999998e-08 1.8898486552485423 1.9462e-08 1.7766649521382964 1.9463e-08 1.835034412195309 1.9463999999999998e-08 1.8010056667448928 1.9465e-08 1.8498536894974895 1.9466e-08 1.7660561028394617 1.9466999999999998e-08 1.761892868139911 1.9468e-08 1.7876483275676667 1.9469e-08 1.7836607092166628 1.9469999999999998e-08 1.6145992737432675 1.9471e-08 1.8723891324389759 1.9472e-08 1.789731277225077 1.9473e-08 1.7656799187394647 1.9474e-08 1.7580725944852837 1.9475e-08 1.8071249336712962 1.9476e-08 1.8134590157450121 1.9477e-08 1.7677221520758666 1.9478e-08 1.8059180017194856 1.9479e-08 1.858927694014484 1.948e-08 1.8231005635484432 1.9481e-08 1.8101784446090916 1.9482e-08 1.737538474804773 1.9483e-08 1.8423018618147275 1.9484e-08 1.8670979827693401 1.9485e-08 1.8099858053579274 1.9486e-08 1.8114405566091174 1.9487e-08 1.778042776823952 1.9488e-08 1.8453758510328464 1.9489e-08 1.7635915658114456 1.949e-08 1.8273844837088107 1.9491e-08 1.9006895751787583 1.9492e-08 1.848741017309328 1.9493e-08 1.77702626762556 1.9494e-08 1.8842404464799694 1.9495e-08 1.765141589953735 1.9495999999999998e-08 1.8627854862120299 1.9497e-08 1.8104967917659982 1.9498e-08 1.8169907011520998 1.9498999999999998e-08 1.834685461801174 1.95e-08 1.7778244884561667 1.9501e-08 1.8067418282854921 1.9501999999999998e-08 1.7907785653048898 1.9503e-08 1.724853869874516 1.9504e-08 1.7241215451430165 1.9504999999999998e-08 1.7397812164816036 1.9506e-08 1.7998857844910523 1.9507e-08 1.777988742128472 1.9508e-08 1.7874297121541396 1.9509e-08 1.818064107238154 1.951e-08 1.7049322637863429 1.9511e-08 1.8120622407851987 1.9512e-08 1.7726719337967183 1.9513e-08 1.7825013956052174 1.9514e-08 1.8493167449294938 1.9515e-08 1.7955090784606798 1.9516e-08 1.8972559120371622 1.9517e-08 1.8617702017766535 1.9518e-08 1.7488740519900074 1.9519e-08 1.7928921488429446 1.952e-08 1.8248387520548424 1.9521e-08 1.7796671218455091 1.9522e-08 1.8038240935408947 1.9523e-08 1.7386161608459152 1.9524e-08 1.8324365588861677 1.9525e-08 1.7418179638143758 1.9526e-08 1.7790479911039618 1.9527e-08 1.8612258721245776 1.9528e-08 1.7638260563726142 1.9529e-08 1.699028058542194 1.953e-08 1.8530618554704001 1.9530999999999998e-08 1.876533960135196 1.9532e-08 1.862671882305641 1.9533e-08 1.7772237003348699 1.9533999999999998e-08 1.8308557589114551 1.9535e-08 1.808236741777126 1.9536e-08 1.8327610552649267 1.9536999999999998e-08 1.7765307561083914 1.9538e-08 1.769792502891114 1.9539e-08 1.7452527847259678 1.9539999999999998e-08 1.8189065534681224 1.9541e-08 1.762764083602818 1.9542e-08 1.7288936754680468 1.9543e-08 1.8191257105341792 1.9544e-08 1.888477075880001 1.9545e-08 1.7928562654477023 1.9546e-08 1.850089582405084 1.9547e-08 1.7635576836457432 1.9548e-08 1.878013761397137 1.9549e-08 1.8295402014361124 1.955e-08 1.7849458562709624 1.9551e-08 1.7853205363557192 1.9552e-08 1.8837081253780659 1.9553e-08 1.862045645022357 1.9554e-08 1.7871950377909338 1.9555e-08 1.7508223425125575 1.9556e-08 1.844001497906766 1.9557e-08 1.7185263747027382 1.9558e-08 1.7420722328810485 1.9559e-08 1.8319277978781325 1.956e-08 1.8925407935581258 1.9561e-08 1.7684737076321673 1.9562e-08 1.7536955691816214 1.9563e-08 1.798857529445886 1.9564e-08 1.7706192755905434 1.9565e-08 1.85515186809247 1.9565999999999998e-08 1.7513570993565895 1.9567e-08 1.7359825566869036 1.9568e-08 1.823536892494605 1.9568999999999998e-08 1.7429107814798168 1.957e-08 1.8666756610866724 1.9571e-08 1.7984325100820935 1.9571999999999998e-08 1.7624028434935664 1.9573e-08 1.8308835856519758 1.9574e-08 1.7559855059248557 1.9574999999999998e-08 1.8164834552701155 1.9576e-08 1.7548534061442853 1.9577e-08 1.8017137920636934 1.9578e-08 1.8103560272977948 1.9579e-08 1.7918968528332133 1.958e-08 1.7925468700537746 1.9581e-08 1.7415318132547284 1.9582e-08 1.805584635384901 1.9583e-08 1.8505069819579774 1.9584e-08 1.8145350982361046 1.9585e-08 1.7966612466365581 1.9586e-08 1.7822518441272672 1.9587e-08 1.7769455285861313 1.9588e-08 1.8631296953192835 1.9589e-08 1.826856992261831 1.959e-08 1.8463463513358531 1.9591e-08 1.851770766807009 1.9592e-08 1.817316216116583 1.9593e-08 1.8836253397590579 1.9594e-08 1.7942269418980368 1.9595e-08 1.841974602393788 1.9596e-08 1.7869016621547464 1.9597e-08 1.927714916059751 1.9598e-08 1.887178517903531 1.9599e-08 1.8322112812611377 1.96e-08 1.7944419192124053 1.9600999999999998e-08 1.7593099337778857 1.9602e-08 1.8304919073959889 1.9603e-08 1.8387035016999111 1.9603999999999998e-08 1.85798780727848 1.9605e-08 1.898901194874536 1.9606e-08 1.7940361681461194 1.9606999999999998e-08 1.8359959341868837 1.9608e-08 1.8210724583988038 1.9609e-08 1.7955485733527423 1.9609999999999998e-08 1.7189324080645307 1.9611e-08 1.8024187918661259 1.9612e-08 1.814795158946554 1.9612999999999998e-08 1.8326576053917896 1.9614e-08 1.7749340821440864 1.9615e-08 1.8900826821921612 1.9616e-08 1.7748583084809377 1.9617e-08 1.8166020044393383 1.9618e-08 1.7688525943825377 1.9619e-08 1.6927565078584708 1.962e-08 1.7676085338621048 1.9621e-08 1.8075706891847938 1.9622e-08 1.7289158305694154 1.9623e-08 1.7704850035428714 1.9624e-08 1.8800152466885653 1.9625e-08 1.866321997329938 1.9626e-08 1.831781892279337 1.9627e-08 1.7922281838628562 1.9628e-08 1.8029768949599405 1.9629e-08 1.7792626529557918 1.963e-08 1.748834701543677 1.9631e-08 1.8499552374448938 1.9632e-08 1.8160134074253187 1.9633e-08 1.8357577763835056 1.9634e-08 1.7370303327866483 1.9635e-08 1.7374264518037352 1.9635999999999998e-08 1.822694010920332 1.9637e-08 1.8095932476297751 1.9638e-08 1.8830178800108903 1.9638999999999998e-08 1.8441356722936186 1.964e-08 1.8550946762916443 1.9641e-08 1.7650413578848594 1.9641999999999998e-08 1.8382401340165784 1.9643e-08 1.8401782165485798 1.9644e-08 1.795334287244319 1.9644999999999998e-08 1.7671488731242284 1.9646e-08 1.7530027301696467 1.9647e-08 1.8302332846597826 1.9647999999999998e-08 1.8444290476240677 1.9649e-08 1.7946775313554535 1.965e-08 1.7351244324116042 1.9651e-08 1.7776193908488735 1.9652e-08 1.7762087173270347 1.9653e-08 1.7553501594198382 1.9654e-08 1.7796970081833736 1.9655e-08 1.779966146797162 1.9656e-08 1.770373736083491 1.9657e-08 1.8504639708987083 1.9658e-08 1.7648229795786485 1.9659e-08 1.7486209907866188 1.966e-08 1.759724579770242 1.9661e-08 1.7648627256613745 1.9662e-08 1.7790450689027202 1.9663e-08 1.787160410109535 1.9664e-08 1.8260495080821268 1.9665e-08 1.7612099961722425 1.9666e-08 1.7252363663735681 1.9667e-08 1.8205782988928703 1.9668e-08 1.8625220683501742 1.9669e-08 1.8073538930401034 1.967e-08 1.810871330264056 1.9671e-08 1.765590743568377 1.9672e-08 1.833420440616139 1.9673e-08 1.7499447831671278 1.9673999999999998e-08 1.8781968889061085 1.9675e-08 1.8082657362698284 1.9676e-08 1.817353647248844 1.9676999999999998e-08 1.708275173460874 1.9678e-08 1.7213665308389603 1.9679e-08 1.8664950854581717 1.9679999999999998e-08 1.7211413856369715 1.9681e-08 1.742749251102404 1.9682e-08 1.8351604930902394 1.9682999999999998e-08 1.778358748773756 1.9684e-08 1.8735723325853453 1.9685e-08 1.6779912690526722 1.9686e-08 1.8038065032579669 1.9687e-08 1.9026339152610983 1.9688e-08 1.800546880225852 1.9689e-08 1.818886920293194 1.969e-08 1.8388958291125688 1.9691e-08 1.8053956953775199 1.9692e-08 1.7971093530497784 1.9693e-08 1.655880047647208 1.9694e-08 1.7531032818866503 1.9695e-08 1.7309501548038098 1.9696e-08 1.7470776215401957 1.9697e-08 1.8143355113980082 1.9698e-08 1.7735296084804262 1.9699e-08 1.8234894499356733 1.97e-08 1.7083760786131654 1.9701e-08 1.913156955852651 1.9702e-08 1.8401652695111692 1.9703e-08 1.8637146807777152 1.9704e-08 1.7134674674087378 1.9705e-08 1.7460732162432904 1.9706e-08 1.897538358217633 1.9707e-08 1.8191338832384445 1.9708e-08 1.7410151595412215 1.9708999999999998e-08 1.8482226658096252 1.971e-08 1.8468141174772472 1.9711e-08 1.7883689168299342 1.9711999999999998e-08 1.80676913909354 1.9713e-08 1.8115797188864309 1.9714e-08 1.7685333861915333 1.9714999999999998e-08 1.7419423617818424 1.9716e-08 1.8439603881840534 1.9717e-08 1.8188912575166012 1.9717999999999998e-08 1.7570986755651268 1.9719e-08 1.7655405092422338 1.972e-08 1.829949081254352 1.9721e-08 1.7680266956507324 1.9722e-08 1.8258854041162507 1.9723e-08 1.8754798561300257 1.9724e-08 1.7614916161009628 1.9725e-08 1.6803493889957877 1.9726e-08 1.8359653332549812 1.9727e-08 1.8918665180360579 1.9728e-08 1.9145399849625355 1.9729e-08 1.7249255480919814 1.973e-08 1.773427534145729 1.9731e-08 1.8183029149959948 1.9732e-08 1.8050325567230165 1.9733e-08 1.738429020661789 1.9734e-08 1.7541918510942967 1.9735e-08 1.7305689125571402 1.9736e-08 1.7198856493681658 1.9737e-08 1.8062412014608837 1.9738e-08 1.749290400943384 1.9739e-08 1.8171663849225979 1.974e-08 1.7108943771488752 1.9741e-08 1.7768384423358898 1.9742e-08 1.7977950776396383 1.9743e-08 1.8536678355599356 1.9743999999999998e-08 1.7657077096705693 1.9745e-08 1.7205893332088185 1.9746e-08 1.8033274285039858 1.9746999999999998e-08 1.8225691088357965 1.9748e-08 1.9203003120295055 1.9749e-08 1.8089765878289197 1.9749999999999998e-08 1.7571425351506769 1.9751e-08 1.7740229049826284 1.9752e-08 1.8311398217776764 1.9752999999999998e-08 1.7575177904191546 1.9754e-08 1.8049721030128079 1.9755e-08 1.8682733214538791 1.9756e-08 1.8497109030411105 1.9757e-08 1.783221569511998 1.9758e-08 1.8001217079342064 1.9759e-08 1.788656267705156 1.976e-08 1.8209756456060475 1.9761e-08 1.7026162859128768 1.9762e-08 1.8134627694169856 1.9763e-08 1.867597652036374 1.9764e-08 1.8104645208299932 1.9765e-08 1.7654876848207397 1.9766e-08 1.8187265065084357 1.9767e-08 1.825720325717463 1.9768e-08 1.7687550266729803 1.9769e-08 1.8674710602560143 1.977e-08 1.8215312631726976 1.9771e-08 1.7879687696508926 1.9772e-08 1.80707969200704 1.9773e-08 1.8465972602767369 1.9774e-08 1.7297275520572375 1.9775e-08 1.7886678349486465 1.9776e-08 1.7361993002412275 1.9777e-08 1.8762909360060307 1.9778e-08 1.8911360714898706 1.9778999999999998e-08 1.8450317946711359 1.978e-08 1.8333226507427165 1.9781e-08 1.7672304086565729 1.9781999999999998e-08 1.7739496089288749 1.9783e-08 1.6589290596329835 1.9784e-08 1.7113615555815418 1.9784999999999998e-08 1.7605762525894928 1.9786e-08 1.8226840117732 1.9787e-08 1.698623547723318 1.9787999999999998e-08 1.7612863892135406 1.9789e-08 1.7548035205071 1.979e-08 1.8010555665225028 1.9791e-08 1.939956086525996 1.9792e-08 1.8229011881761306 1.9793e-08 1.7672784656516878 1.9794e-08 1.7995755342541857 1.9795e-08 1.7876405942296199 1.9796e-08 1.7833403109810126 1.9797e-08 1.735237815267397 1.9798e-08 1.8144978632250843 1.9799e-08 1.8204264214581911 1.98e-08 1.9189775910954194 1.9801e-08 1.8582811777470363 1.9802e-08 1.8647434670906253 1.9803e-08 1.798727271310024 1.9804e-08 1.857929629773993 1.9805e-08 1.8431809622653528 1.9806e-08 1.8638914898743444 1.9807e-08 1.772774390617496 1.9808e-08 1.8068290243183636 1.9809e-08 1.7876481000357303 1.981e-08 1.76628577248287 1.9811e-08 1.7887421098330885 1.9812e-08 1.7856623221138157 1.9813e-08 1.873853168692715 1.9813999999999998e-08 1.7497525706546035 1.9815e-08 1.8292608632369123 1.9816e-08 1.7628941653549306 1.9816999999999998e-08 1.8064738014095916 1.9818e-08 1.8106614837882355 1.9819e-08 1.6988649184669837 1.9819999999999998e-08 1.8500812333807413 1.9821e-08 1.8466182045973074 1.9822e-08 1.7695662073015328 1.9822999999999998e-08 1.8319621000946884 1.9824e-08 1.7596067538253297 1.9825e-08 1.8256137620517758 1.9825999999999998e-08 1.7731609169626754 1.9827e-08 1.745938287752928 1.9828e-08 1.8656299043055597 1.9829e-08 1.8819802770891687 1.983e-08 1.8781201431017422 1.9831e-08 1.8263461116331559 1.9832e-08 1.862483366902365 1.9833e-08 1.740243198159667 1.9834e-08 1.755238803396808 1.9835e-08 1.8005303135742896 1.9836e-08 1.8799161245667118 1.9837e-08 1.805878785702826 1.9838e-08 1.8030511872598158 1.9839e-08 1.8097513390600695 1.984e-08 1.7980361600652743 1.9841e-08 1.795411088141593 1.9842e-08 1.8323267972073352 1.9843e-08 1.8137664899642076 1.9844e-08 1.7480875955787292 1.9845e-08 1.7519641190541524 1.9846e-08 1.7399054345371052 1.9847e-08 1.8125748083594844 1.9848e-08 1.8690574528139923 1.9849e-08 1.8854825830979727 1.985e-08 1.7911680996080706 1.9851e-08 1.7954338691637812 1.9851999999999998e-08 1.8077776160334857 1.9853e-08 1.7957082002469924 1.9854e-08 1.749702266241559 1.9854999999999998e-08 1.7127882978329776 1.9856e-08 1.8470007052872623 1.9857e-08 1.7654105736148382 1.9857999999999998e-08 1.7867764871596754 1.9859e-08 1.8068233263979576 1.986e-08 1.7069437876097635 1.9860999999999998e-08 1.7891006978164607 1.9862e-08 1.7509945764059012 1.9863e-08 1.889643123015622 1.9864e-08 1.7738701810516544 1.9865e-08 1.8069247280233938 1.9866e-08 1.8855739703271819 1.9867e-08 1.7781784718283462 1.9868e-08 1.7639161382250723 1.9869e-08 1.73154877511313 1.987e-08 1.8067516882943258 1.9871e-08 1.746834682185604 1.9872e-08 1.8422255417498854 1.9873e-08 1.79724958995095 1.9874e-08 1.8326428111936313 1.9875e-08 1.8005389297654255 1.9876e-08 1.8040678174751361 1.9877e-08 1.8899438459558775 1.9878e-08 1.7873047465957985 1.9879e-08 1.8566833371882547 1.988e-08 1.7523445051422917 1.9881e-08 1.8119731997126098 1.9882e-08 1.6845797915517513 1.9883e-08 1.7169128262872995 1.9884e-08 1.7501604737723897 1.9885e-08 1.8818789109479952 1.9886e-08 1.797653369985649 1.9886999999999998e-08 1.7916934598986893 1.9888e-08 1.8067964483284595 1.9889e-08 1.8521792279755391 1.9889999999999998e-08 1.8268987952427858 1.9891e-08 1.8143607471635976 1.9892e-08 1.7952436728719394 1.9892999999999998e-08 1.8799043570321958 1.9894e-08 1.7467650823398428 1.9895e-08 1.7373130871083426 1.9895999999999998e-08 1.8335631955132303 1.9897e-08 1.7302202142441525 1.9898e-08 1.7982848835909373 1.9899e-08 1.905326286450712 1.99e-08 1.8311748502704945 1.9901e-08 1.803194657892167 1.9902e-08 1.8258808509146933 1.9903e-08 1.8505366427706975 1.9904e-08 1.7510707237021275 1.9905e-08 1.7652187457502413 1.9906e-08 1.83019913675763 1.9907e-08 1.8417243452147192 1.9908e-08 1.8033898612394093 1.9909e-08 1.721628813693505 1.991e-08 1.837798358759774 1.9911e-08 1.8096002042371893 1.9912e-08 1.8272663826391675 1.9913e-08 1.8161379302062275 1.9914e-08 1.7358312642306384 1.9915e-08 1.7638267209730025 1.9916e-08 1.6802663181631232 1.9917e-08 1.8177882707986008 1.9918e-08 1.8295518837358682 1.9919e-08 1.8618554716344593 1.992e-08 1.7569443167555745 1.9921e-08 1.7691782950019928 1.9921999999999998e-08 1.8100959769474068 1.9923e-08 1.7943567686100055 1.9924e-08 1.7930651818995513 1.9924999999999998e-08 1.8055062987989017 1.9926e-08 1.7113498648392766 1.9927e-08 1.8894841364031254 1.9927999999999998e-08 1.836433012580359 1.9929e-08 1.7830569686074231 1.993e-08 1.8531138232783622 1.9930999999999998e-08 1.7582747340827451 1.9932e-08 1.7983412936719925 1.9933e-08 1.76652821247363 1.9934e-08 1.7872026881563448 1.9935e-08 1.804224312294012 1.9936e-08 1.8028294514530019 1.9937e-08 1.7855258127049083 1.9938e-08 1.730738035349901 1.9939e-08 1.8064235970637317 1.994e-08 1.8264021544620497 1.9941e-08 1.7879301279018298 1.9942e-08 1.8446601580584328 1.9943e-08 1.8119427584789716 1.9944e-08 1.8123261093447816 1.9945e-08 1.801416482337739 1.9946e-08 1.8175058275152391 1.9947e-08 1.7315668144722698 1.9948e-08 1.819627552738542 1.9949e-08 1.798037357965626 1.995e-08 1.7949274217280144 1.9951e-08 1.8053108406329987 1.9952e-08 1.765720593533762 1.9953e-08 1.7481075922718936 1.9954e-08 1.8215011988858751 1.9955e-08 1.8637509651995718 1.9956e-08 1.845344158267973 1.9956999999999998e-08 1.8359750644164219 1.9958e-08 1.8492432523959237 1.9959e-08 1.8415493131433265 1.9959999999999998e-08 1.8287569688315903 1.9961e-08 1.8159897215659808 1.9962e-08 1.7264724874156658 1.9962999999999998e-08 1.8045472219047167 1.9964e-08 1.7436372450431639 1.9965e-08 1.844264960123345 1.9965999999999998e-08 1.7807064472039948 1.9967e-08 1.7174854001399307 1.9968e-08 1.8100963048808965 1.9969e-08 1.8323095006263816 1.997e-08 1.792619715541217 1.9971e-08 1.7236199460609472 1.9972e-08 1.8459199343164532 1.9973e-08 1.822561735060301 1.9974e-08 1.7931249850097235 1.9975e-08 1.783373736688271 1.9976e-08 1.83860872929745 1.9977e-08 1.7844978274216028 1.9978e-08 1.877031111866026 1.9979e-08 1.8171627856823975 1.998e-08 1.8214539720219995 1.9981e-08 1.7704992451299384 1.9982e-08 1.8588369877568385 1.9983e-08 1.8011939161907642 1.9984e-08 1.7766894541503788 1.9985e-08 1.8361970702688415 1.9986e-08 1.8293231674474462 1.9987e-08 1.7148652915372773 1.9988e-08 1.7735055418854608 1.9989e-08 1.8165798674495102 1.999e-08 1.861868116725602 1.9991e-08 1.7824300524839125 1.9991999999999998e-08 1.8265038197100674 1.9993e-08 1.7755109113524774 1.9994e-08 1.7920384825946376 1.9994999999999998e-08 1.7635880377444304 1.9996e-08 1.7517661569868324 1.9997e-08 1.8771690639538852 1.9997999999999998e-08 1.8536947806248643 1.9999e-08 1.8617552112161313 2e-08 1.7826633874071816 2.0000999999999998e-08 1.8768143594209965 2.0002e-08 1.7907070477437221 2.0003e-08 1.8137872580065244 2.0003999999999998e-08 1.7767007602799003 2.0005e-08 1.8205877754513549 2.0006e-08 1.8404420562423207 2.0007e-08 1.744526247125775 2.0008e-08 1.7635407192200647 2.0009e-08 1.8159282757299444 2.001e-08 1.7921223005234508 2.0011e-08 1.8558967504601214 2.0012e-08 1.7946744362941578 2.0013e-08 1.856314953223571 2.0014e-08 1.9140669403543216 2.0015e-08 1.879997746654265 2.0016e-08 1.7904946196239366 2.0017e-08 1.7947346436606535 2.0018e-08 1.7504301137522553 2.0019e-08 1.7814704063645888 2.002e-08 1.84003456331119 2.0021e-08 1.8053598384488994 2.0022e-08 1.7968515378067345 2.0023e-08 1.7623047630963262 2.0024e-08 1.7679118557722049 2.0025e-08 1.85823417822606 2.0026e-08 1.8154748543223365 2.0026999999999998e-08 1.8339227160897582 2.0028e-08 1.749581291563052 2.0029e-08 1.8073928532465509 2.0029999999999998e-08 1.7251379740861028 2.0031e-08 1.7533505322422245 2.0032e-08 1.7974022241389926 2.0032999999999998e-08 1.7258093403606813 2.0034e-08 1.753058297671987 2.0035e-08 1.6955254079800337 2.0035999999999998e-08 1.8808546221879494 2.0037e-08 1.7879069501408915 2.0038e-08 1.7861350765061808 2.0038999999999998e-08 1.7910973805346329 2.004e-08 1.7959499592736092 2.0041e-08 1.8782056314374782 2.0042e-08 1.7455294175688678 2.0043e-08 1.8500949450773456 2.0044e-08 1.8206336020515355 2.0045e-08 1.8527911637640213 2.0046e-08 1.8291856945727645 2.0047e-08 1.7529805906732412 2.0048e-08 1.8546806948882846 2.0049e-08 1.7423558552941893 2.005e-08 1.8625724471856413 2.0051e-08 1.8946843120014067 2.0052e-08 1.779833916217945 2.0053e-08 1.895421173169095 2.0054e-08 1.799965417477526 2.0055e-08 1.8246581113304825 2.0056e-08 1.8485428024819912 2.0057e-08 1.880189382613251 2.0058e-08 1.7672028135128408 2.0059e-08 1.8665968042972085 2.006e-08 1.8129450945865864 2.0061e-08 1.7346985017069738 2.0062e-08 1.6158542269804714 2.0063e-08 1.7776577034201486 2.0064e-08 1.774379579333484 2.0064999999999998e-08 1.765292036774319 2.0066e-08 1.7326702218873842 2.0067e-08 1.9684330263487149 2.0067999999999998e-08 1.780221923085206 2.0069e-08 1.7431175276291455 2.007e-08 1.8813818364249377 2.0070999999999998e-08 1.7693266921998987 2.0072e-08 1.8244439104945762 2.0073e-08 1.827888201307842 2.0073999999999998e-08 1.7762395911494138 2.0075e-08 1.8081235267841569 2.0076e-08 1.7040563339123331 2.0077e-08 1.785247136462405 2.0078e-08 1.838053714559865 2.0079e-08 1.8107918400919434 2.008e-08 1.8768858852621477 2.0081e-08 1.84313853898733 2.0082e-08 1.7724657469925258 2.0083e-08 1.8141079883537345 2.0084e-08 1.857229180518563 2.0085e-08 1.8548462096820477 2.0086e-08 1.7754868699989943 2.0087e-08 1.812967626476783 2.0088e-08 1.7648282621639755 2.0089e-08 1.8219894740936755 2.009e-08 1.8210334193075322 2.0091e-08 1.7976014240451197 2.0092e-08 1.8034289703472353 2.0093e-08 1.779080953049617 2.0094e-08 1.8054895462100424 2.0095e-08 1.775634014520736 2.0096e-08 1.763555958300756 2.0097e-08 1.820269550132876 2.0098e-08 1.8418552017239695 2.0099e-08 1.7998013548134717 2.0099999999999998e-08 1.886129473097341 2.0101e-08 1.8011502851591787 2.0102e-08 1.7350542412550514 2.0102999999999998e-08 1.8578886839958288 2.0104e-08 1.9366884651446867 2.0105e-08 1.7084747793702353 2.0105999999999998e-08 1.71245344161423 2.0107e-08 1.8591739115843398 2.0108e-08 1.8945668227403525 2.0108999999999998e-08 1.6951039149188334 2.011e-08 1.8253843067126407 2.0111e-08 1.890362905387616 2.0112e-08 1.864358651674461 2.0113e-08 1.6794109984545025 2.0114e-08 1.7693716019459977 2.0115e-08 1.7436655204039702 2.0116e-08 1.5852527960313325 2.0117e-08 1.817416281669747 2.0118e-08 1.8038196342704416 2.0119e-08 1.742796755864123 2.012e-08 1.778804914629962 2.0121e-08 1.8519934490355912 2.0122e-08 1.736091157112363 2.0123e-08 1.841102906303781 2.0124e-08 1.8350643382825957 2.0125e-08 1.7407399251939235 2.0126e-08 1.815860812955918 2.0127e-08 1.880643538365961 2.0128e-08 1.7821479545279624 2.0129e-08 1.7997105467311556 2.013e-08 1.862439700398013 2.0131e-08 1.72334703885727 2.0132e-08 1.8808494779212805 2.0133e-08 1.811091069253484 2.0134e-08 1.7965081058669052 2.0134999999999998e-08 1.6464606147733511 2.0136e-08 1.7392873698139013 2.0137e-08 1.8669757857130773 2.0137999999999998e-08 1.8458233208759565 2.0139e-08 1.8280293099675826 2.014e-08 1.7732748167506824 2.0140999999999998e-08 1.9162434391810073 2.0142e-08 1.8563286933459264 2.0143e-08 1.7822967363900168 2.0143999999999998e-08 1.8703353989127982 2.0145e-08 1.8082314566077524 2.0146e-08 1.8302556111981299 2.0147e-08 1.8992775829006743 2.0148e-08 1.7736533236307934 2.0149e-08 1.8208952001762566 2.015e-08 1.8224843958656227 2.0151e-08 1.6617513063705789 2.0152e-08 1.8041514852728404 2.0153e-08 1.8314962517594953 2.0154e-08 1.744342190840657 2.0155e-08 1.6933203898029716 2.0156e-08 1.810825634733435 2.0157e-08 1.7272311148547703 2.0158e-08 1.7461910919766233 2.0159e-08 1.8156785939518545 2.016e-08 1.691634720511213 2.0161e-08 1.7535187278204487 2.0162e-08 1.7879738775302305 2.0163e-08 1.6865775596844221 2.0164e-08 1.8307510731643515 2.0165e-08 1.8214889901083247 2.0166e-08 1.7495576679775209 2.0167e-08 1.744376099593271 2.0168e-08 1.8263092987357616 2.0169e-08 1.7949797490267339 2.0169999999999998e-08 1.7600244979644797 2.0171e-08 1.8420889780940566 2.0172e-08 1.839489775573826 2.0172999999999998e-08 1.7298117479121682 2.0174e-08 1.8235511728908393 2.0175e-08 1.8838872533453777 2.0175999999999998e-08 1.8209380020699877 2.0177e-08 1.7524911840821755 2.0178e-08 1.7014062118932434 2.0178999999999998e-08 1.7344818726402966 2.018e-08 1.7463814113303158 2.0181e-08 1.822761990808526 2.0181999999999998e-08 1.7918498445876776 2.0183e-08 1.7202359325907435 2.0184e-08 1.809268971024313 2.0185e-08 1.7830657359493447 2.0186e-08 1.7781569727406366 2.0187e-08 1.8713285488623443 2.0188e-08 1.7549462703014478 2.0189e-08 1.8073359815971262 2.019e-08 1.7495463010504475 2.0191e-08 1.7442045134997044 2.0192e-08 1.7075560296613328 2.0193e-08 1.7371855858122882 2.0194e-08 1.844299010129528 2.0195e-08 1.7950581157115248 2.0196e-08 1.8007343564012586 2.0197e-08 1.7682768835030551 2.0198e-08 1.754364325538012 2.0199e-08 1.8035114070751532 2.02e-08 1.7275346382933723 2.0201e-08 1.7764907273883523 2.0202e-08 1.7311463081899119 2.0203e-08 1.7911460812139475 2.0204e-08 1.7616428010415754 2.0204999999999998e-08 1.839386834508348 2.0206e-08 1.7663922234718339 2.0207e-08 1.8708326434723337 2.0207999999999998e-08 1.8040790254263372 2.0209e-08 1.8458296995420744 2.021e-08 1.840472297002773 2.0210999999999998e-08 1.8239501859197964 2.0212e-08 1.8175025671351206 2.0213e-08 1.7978842841736042 2.0213999999999998e-08 1.8566717240757424 2.0215e-08 1.7552784273039568 2.0216e-08 1.8140896136980142 2.0216999999999998e-08 1.61636432281688 2.0218e-08 1.7148197560297571 2.0219e-08 1.7808149052347886 2.022e-08 1.779794311271508 2.0221e-08 1.8367280500054495 2.0222e-08 1.76901144379444 2.0223e-08 1.8471971465761214 2.0224e-08 1.7395632709785345 2.0225e-08 1.7326462711684019 2.0226e-08 1.8796081404598455 2.0227e-08 1.864697196178695 2.0228e-08 1.8220767378859326 2.0229e-08 1.8494317151946613 2.023e-08 1.8206355786291344 2.0231e-08 1.7984469075209883 2.0232e-08 1.8001308531629117 2.0233e-08 1.819842829049982 2.0234e-08 1.8019063669531983 2.0235e-08 1.7473438905305236 2.0236e-08 1.7854365242379469 2.0237e-08 1.7591923309151845 2.0238e-08 1.7744073246029468 2.0239e-08 1.7315159114483532 2.024e-08 1.7248754523982632 2.0241e-08 1.8483311021165003 2.0242e-08 1.8129774887217902 2.0242999999999998e-08 1.8231547982149678 2.0244e-08 1.7535568647069795 2.0245e-08 1.8266258114647027 2.0245999999999998e-08 1.7707232114770937 2.0247e-08 1.818250739194038 2.0248e-08 1.833554790688195 2.0248999999999998e-08 1.8369719558959348 2.025e-08 1.8571882160483673 2.0251e-08 1.7527461924715464 2.0251999999999998e-08 1.8697100194475758 2.0253e-08 1.870039746873775 2.0254e-08 1.737883581532081 2.0255e-08 1.819590376564304 2.0256e-08 1.8170557260422433 2.0257e-08 1.809215621911209 2.0258e-08 1.70792734443404 2.0259e-08 1.8348694670217496 2.026e-08 1.738815945745135 2.0261e-08 1.7459591419903 2.0262e-08 1.765792926860827 2.0263e-08 1.8323175157288456 2.0264e-08 1.7286304557176668 2.0265e-08 1.8515391975065292 2.0266e-08 1.7961749200305788 2.0267e-08 1.7785053411440062 2.0268e-08 1.7513545706878788 2.0269e-08 1.8429550306297369 2.027e-08 1.775705824008545 2.0271e-08 1.791591377726922 2.0272e-08 1.8813730749172697 2.0273e-08 1.8260408497781688 2.0274e-08 1.8326818566899254 2.0275e-08 1.753624273622822 2.0276e-08 1.795353097235919 2.0277e-08 1.7995802173850373 2.0277999999999998e-08 1.7364944671733968 2.0279e-08 1.7871082480200626 2.028e-08 1.7488257993784355 2.0280999999999998e-08 1.8400119701096926 2.0282e-08 1.788920413646329 2.0283e-08 1.83514828574622 2.0283999999999998e-08 1.8331160598879406 2.0285e-08 1.7846230092894584 2.0286e-08 1.865032286016085 2.0286999999999998e-08 1.7639117195564245 2.0288e-08 1.8697111916900215 2.0289e-08 1.7801173389921499 2.029e-08 1.8173501608440183 2.0291e-08 1.7792284656440522 2.0292e-08 1.8321167147366575 2.0293e-08 1.816373152796537 2.0294e-08 1.8176972935089488 2.0295e-08 1.7028307384938655 2.0296e-08 1.687380100880904 2.0297e-08 1.7909370361694634 2.0298e-08 1.7627411529189176 2.0299e-08 1.7711184808560354 2.03e-08 1.7197231775358073 2.0301e-08 1.751126949070735 2.0302e-08 1.821082001269142 2.0303e-08 1.8475433922842015 2.0304e-08 1.6979365664141417 2.0305e-08 1.74099491603127 2.0306e-08 1.8730882274199072 2.0307e-08 1.8453486597533466 2.0308e-08 1.7914799587656582 2.0309e-08 1.7363691211830719 2.031e-08 1.926929389061417 2.0311e-08 1.7644736991299197 2.0312e-08 1.7612929464139562 2.0312999999999998e-08 1.8284704177228488 2.0314e-08 1.8288872914673477 2.0315e-08 1.7837685874319358 2.0315999999999998e-08 1.7870266509741053 2.0317e-08 1.8242214071329175 2.0318e-08 1.9077016404166596 2.0318999999999998e-08 1.8062544433978214 2.032e-08 1.8507837631006505 2.0321e-08 1.811777805301 2.0321999999999998e-08 1.760073471371638 2.0323e-08 1.7632290268312738 2.0324e-08 1.8355892766448594 2.0325e-08 1.892437925361124 2.0326e-08 1.7958847426416429 2.0327e-08 1.8297480575062215 2.0328e-08 1.7065898966948472 2.0329e-08 1.809933416405001 2.033e-08 1.8129909245372435 2.0331e-08 1.7878055525738106 2.0332e-08 1.781118064426138 2.0333e-08 1.7504450190306755 2.0334e-08 1.8049819069701687 2.0335e-08 1.820103360969934 2.0336e-08 1.8347428597377673 2.0337e-08 1.7723029238195822 2.0338e-08 1.8368202207968558 2.0339e-08 1.7967799027025353 2.034e-08 1.8219324026469617 2.0341e-08 1.8180079114570564 2.0342e-08 1.8593919032415411 2.0343e-08 1.8382145472595384 2.0344e-08 1.8553725738202376 2.0345e-08 1.881923202240016 2.0346e-08 1.7977031298332 2.0347e-08 1.826971531595034 2.0347999999999998e-08 1.7806287907890028 2.0349e-08 1.8603822551333047 2.035e-08 1.671869465256742 2.0350999999999998e-08 1.899054744563094 2.0352e-08 1.741941619599606 2.0353e-08 1.774738582743001 2.0353999999999998e-08 1.769513966259091 2.0355e-08 1.7054453633353095 2.0356e-08 1.7296708733977115 2.0356999999999998e-08 1.7707527351250258 2.0358e-08 1.8104760297493854 2.0359e-08 1.7902111596177217 2.036e-08 1.7850244557481139 2.0361e-08 1.8292354641330335 2.0362e-08 1.8207434606868487 2.0363e-08 1.7449442426953472 2.0364e-08 1.7418167141321583 2.0365e-08 1.8325353110251046 2.0366e-08 1.780247869390514 2.0367e-08 1.7114213811559025 2.0368e-08 1.785318180614388 2.0369e-08 1.7617754172782494 2.037e-08 1.8130700019827817 2.0371e-08 1.8697743097149293 2.0372e-08 1.7731515977388175 2.0373e-08 1.7910602097006898 2.0374e-08 1.748954234998814 2.0375e-08 1.7733254667395975 2.0376e-08 1.8348730662606776 2.0377e-08 1.8879631138433317 2.0378e-08 1.8666504780083666 2.0379e-08 1.7578312993984082 2.038e-08 1.8225668431650126 2.0381e-08 1.7561213147585588 2.0382e-08 1.7909978496626018 2.0382999999999998e-08 1.765297474783201 2.0384e-08 1.8589141094435517 2.0385e-08 1.8547292100694965 2.0385999999999998e-08 1.8454928327591473 2.0387e-08 1.7076779571025251 2.0388e-08 1.8602684719584417 2.0388999999999998e-08 1.8294704316912367 2.039e-08 1.757692459877709 2.0391e-08 1.7877944174629932 2.0391999999999998e-08 1.8326796193078891 2.0393e-08 1.773927486880185 2.0394e-08 1.790107448969101 2.0394999999999998e-08 1.8515778964812968 2.0396e-08 1.8242387003706813 2.0397e-08 1.7907104638138092 2.0398e-08 1.7833040373968772 2.0399e-08 1.7506251617073196 2.04e-08 1.8264114082364542 2.0401e-08 1.8218121153914373 2.0402e-08 1.8438311256259483 2.0403e-08 1.7898099089870307 2.0404e-08 1.8540364606276518 2.0405e-08 1.7895411586346945 2.0406e-08 1.7379874750137811 2.0407e-08 1.8322808284165415 2.0408e-08 1.7395397637521248 2.0409e-08 1.8082136176094752 2.041e-08 1.884383390848477 2.0411e-08 1.7905079732694698 2.0412e-08 1.8208938830033174 2.0413e-08 1.7144409390194537 2.0414e-08 1.8175987467409742 2.0415e-08 1.724371612707839 2.0416e-08 1.857242250579442 2.0417e-08 1.8219277576505204 2.0417999999999998e-08 1.789097453638712 2.0419e-08 1.721649172346276 2.042e-08 1.801145973646759 2.0420999999999998e-08 1.7902758472979359 2.0422e-08 1.6847163118222648 2.0423e-08 1.7642312947336372 2.0423999999999998e-08 1.83342563774616 2.0425e-08 1.7927302394264921 2.0426e-08 1.82467090736994 2.0426999999999998e-08 1.8274367539646201 2.0428e-08 1.767675448448652 2.0429e-08 1.754150198029571 2.0429999999999998e-08 1.8557585554844904 2.0431e-08 1.8168796669175251 2.0432e-08 1.820483100534764 2.0433e-08 1.9325503408461708 2.0434e-08 1.76541839620538 2.0435e-08 1.8097976318301898 2.0436e-08 1.8423528680416006 2.0437e-08 1.7717290122863831 2.0438e-08 1.8594906565823264 2.0439e-08 1.8218654299422108 2.044e-08 1.7707745623542501 2.0441e-08 1.8095077861930864 2.0442e-08 1.7846329967055534 2.0443e-08 1.922405743545617 2.0444e-08 1.7427838473173924 2.0445e-08 1.7539340312346863 2.0446e-08 1.7683691750279986 2.0447e-08 1.7949221130388582 2.0448e-08 1.8070937563173657 2.0449e-08 1.8279008793405924 2.045e-08 1.763095586732269 2.0451e-08 1.7864130197725785 2.0452e-08 1.8138460247408583 2.0453e-08 1.897651473887752 2.0454e-08 1.8318203765141965 2.0455e-08 1.8678549633437584 2.0455999999999998e-08 1.7514262272930898 2.0457e-08 1.7115622249952789 2.0458e-08 1.778976611874795 2.0458999999999998e-08 1.7700442879062228 2.046e-08 1.7818949427739543 2.0461e-08 1.8008295633005627 2.0461999999999998e-08 1.7939962578507966 2.0463e-08 1.7569774263720452 2.0464e-08 1.8136784985314807 2.0464999999999998e-08 1.8691406308597271 2.0466e-08 1.8545282375355883 2.0467e-08 1.7106718468459157 2.0468e-08 1.9006641175216374 2.0469e-08 1.8475829685461849 2.047e-08 1.78908852536476 2.0471e-08 1.75412785759254 2.0472e-08 1.853099984847258 2.0473e-08 1.730780108604098 2.0474e-08 1.8230971020105344 2.0475e-08 1.734677811666184 2.0476e-08 1.8220004934929959 2.0477e-08 1.7541727608072288 2.0478e-08 1.871381914347507 2.0479e-08 1.750550093402367 2.048e-08 1.7669384731416866 2.0481e-08 1.8690059392111396 2.0482e-08 1.724567238035913 2.0483e-08 1.7278603727055977 2.0484e-08 1.7806220022213788 2.0485e-08 1.7846635598903648 2.0486e-08 1.7737991221241607 2.0487e-08 1.8095894592221762 2.0488e-08 1.8690375970587012 2.0489e-08 1.846381320486547 2.049e-08 1.8174995729876358 2.0490999999999998e-08 1.829331015782997 2.0492e-08 1.8154035077906792 2.0493e-08 1.7677498016144 2.0493999999999998e-08 1.8213619564782886 2.0495e-08 1.832816096384311 2.0496e-08 1.8007705491948653 2.0496999999999998e-08 1.7377252155140275 2.0498e-08 1.7411764932500113 2.0499e-08 1.855470174327274 2.0499999999999998e-08 1.843791879077906 2.0501e-08 1.7815778482958151 2.0502e-08 1.7924656464651716 2.0503e-08 1.7582896922720617 2.0504e-08 1.7637036376685649 2.0505e-08 1.809122298905516 2.0506e-08 1.8486393458833008 2.0507e-08 1.7598245489738795 2.0508e-08 1.8248551572933742 2.0509e-08 1.7854666581126155 2.051e-08 1.7955282280155773 2.0511e-08 1.767206103854268 2.0512e-08 1.738279322573589 2.0513e-08 1.8067517923701304 2.0514e-08 1.7874123923904546 2.0515e-08 1.794371632612055 2.0516e-08 1.8239792508463426 2.0517e-08 1.8288402846909975 2.0518e-08 1.818293595662638 2.0519e-08 1.8003209426752758 2.052e-08 1.7872686001457843 2.0521e-08 1.7773989687345164 2.0522e-08 1.7939558035388685 2.0523e-08 1.7944821715135582 2.0524e-08 1.7592588349598959 2.0525e-08 1.7537011050655016 2.0525999999999998e-08 1.7439115342091414 2.0527e-08 1.823232445125884 2.0528e-08 1.754835835477111 2.0528999999999998e-08 1.8248839069460552 2.053e-08 1.8449586464792804 2.0531e-08 1.7853520047291447 2.0531999999999998e-08 1.7785632394526072 2.0533e-08 1.8130487864307696 2.0534e-08 1.8007136508921546 2.0534999999999998e-08 1.8759703757412958 2.0536e-08 1.8627267825861742 2.0537e-08 1.804494409826366 2.0538e-08 1.7295820738340242 2.0539e-08 1.7254826378644437 2.054e-08 1.7790009865752219 2.0541e-08 1.7504275111611471 2.0542e-08 1.861901420050397 2.0543e-08 1.782783521052013 2.0544e-08 1.8598943755522157 2.0545e-08 1.7775707040719437 2.0546e-08 1.7430474083676062 2.0547e-08 1.7119644419528226 2.0548e-08 1.7797460847715498 2.0549e-08 1.8638475219554635 2.055e-08 1.844461369790574 2.0551e-08 1.836086940636037 2.0552e-08 1.7267168659209904 2.0553e-08 1.8003707197159955 2.0554e-08 1.8483301129275629 2.0555e-08 1.729267897669196 2.0556e-08 1.6395490859869966 2.0557e-08 1.7231385414398768 2.0558e-08 1.795081582102457 2.0559e-08 1.8592917287541353 2.056e-08 1.8312918408991792 2.0560999999999998e-08 1.828859307428939 2.0562e-08 1.8040700408370953 2.0563e-08 1.8178228828571612 2.0563999999999998e-08 1.896453078955793 2.0565e-08 1.803655398903607 2.0566e-08 1.7678466092729286 2.0566999999999998e-08 1.6783943380225366 2.0568e-08 1.7991269496087061 2.0569e-08 1.7249904551402393 2.0569999999999998e-08 1.830209293320053 2.0571e-08 1.8782703580358842 2.0572e-08 1.831292067681309 2.0572999999999998e-08 1.7488147681568664 2.0574e-08 1.8229568642391725 2.0575e-08 1.8385551817716626 2.0576e-08 1.7934394900045492 2.0577e-08 1.907249159786872 2.0578e-08 1.8290509662095393 2.0579e-08 1.6678000706624805 2.058e-08 1.7886705078566743 2.0581e-08 1.6974078049099206 2.0582e-08 1.7975610243099 2.0583e-08 1.7810894343974617 2.0584e-08 1.823136278279033 2.0585e-08 1.805798990379234 2.0586e-08 1.8144377037311101 2.0587e-08 1.7739063562717121 2.0588e-08 1.8115033470727893 2.0589e-08 1.8094673572207758 2.059e-08 1.826902191465447 2.0591e-08 1.799701094220347 2.0592e-08 1.9018798538159791 2.0593e-08 1.8142242549630843 2.0594e-08 1.8043314479580923 2.0595e-08 1.737194213268353 2.0595999999999998e-08 1.7890211786839625 2.0597e-08 1.8448798105102362 2.0598e-08 1.7610722001430925 2.0598999999999998e-08 1.8545632921643385 2.06e-08 1.8301072607397157 2.0601e-08 1.7253836281803288 2.0601999999999998e-08 1.760979483841203 2.0603e-08 1.7638353258923862 2.0604e-08 1.8385652637086438 2.0604999999999998e-08 1.8260415463884216 2.0606e-08 1.784838440056121 2.0607e-08 1.8181645588023965 2.0607999999999998e-08 1.8937066621170497 2.0609e-08 1.7022821817055918 2.061e-08 1.7780231904402855 2.0611e-08 1.8554463656431872 2.0612e-08 1.7581305644415008 2.0613e-08 1.8137814721077061 2.0614e-08 1.7843861362937652 2.0615e-08 1.7239704487571237 2.0616e-08 1.8221845251683426 2.0617e-08 1.8425363016554588 2.0618e-08 1.764500559624171 2.0619e-08 1.8842264209448154 2.062e-08 1.8245499455560001 2.0621e-08 1.8006218411854513 2.0622e-08 1.8614546419381646 2.0623e-08 1.7199285849035986 2.0624e-08 1.8322536584060756 2.0625e-08 1.7596920570565486 2.0626e-08 1.7634694810285192 2.0627e-08 1.8159559597199566 2.0628e-08 1.883276577519103 2.0629e-08 1.9020948581312611 2.063e-08 1.801346069969332 2.0631e-08 1.7736978947912074 2.0632e-08 1.815631941640606 2.0633e-08 1.743908747261982 2.0633999999999998e-08 1.7663124323699928 2.0635e-08 1.8692685129624291 2.0636e-08 1.7980256350469037 2.0636999999999998e-08 1.7957363530880173 2.0638e-08 1.8271476230599255 2.0639e-08 1.8129405578766091 2.0639999999999998e-08 1.7560961387702014 2.0641e-08 1.7686772345262058 2.0642e-08 1.8492143963549856 2.0642999999999998e-08 1.762670321531473 2.0644e-08 1.8528146530074294 2.0645e-08 1.7822799820437774 2.0646e-08 1.8756182738483946 2.0647e-08 1.692685568796303 2.0648e-08 1.721192450011397 2.0649e-08 1.7880899411359719 2.065e-08 1.7899915983833956 2.0651e-08 1.8461758480716488 2.0652e-08 1.7893467763546211 2.0653e-08 1.809285029927614 2.0654e-08 1.7774742484434882 2.0655e-08 1.7209602722417299 2.0656e-08 1.689386660350569 2.0657e-08 1.759304922435252 2.0658e-08 1.843846063739282 2.0659e-08 1.8508614175628064 2.066e-08 1.8838712172317675 2.0661e-08 1.853274194687521 2.0662e-08 1.8225265671134614 2.0663e-08 1.8585694964076251 2.0664e-08 1.8261941219910562 2.0665e-08 1.80217343984458 2.0666e-08 1.7148568903515042 2.0667e-08 1.8457251913259176 2.0668e-08 1.8179414868979704 2.0668999999999998e-08 1.7644733244099648 2.067e-08 1.7617057373868252 2.0671e-08 1.7103105078163336 2.0671999999999998e-08 1.823924509863972 2.0673e-08 1.7120715094686052 2.0674e-08 1.8164612962594056 2.0674999999999998e-08 1.7949552136527358 2.0676e-08 1.8261814205041265 2.0677e-08 1.7913223916810428 2.0677999999999998e-08 1.7044333829800085 2.0679e-08 1.7333351910288979 2.068e-08 1.8399596435822558 2.0681e-08 1.7624650451292632 2.0682e-08 1.7968474512339383 2.0683e-08 1.7674161829382213 2.0684e-08 1.8020090111475313 2.0685e-08 1.801734881639197 2.0686e-08 1.7224628837345661 2.0687e-08 1.8345122784302441 2.0688e-08 1.7974277317871503 2.0689e-08 1.8035357046851697 2.069e-08 1.8435568353870002 2.0691e-08 1.7939846477211991 2.0692e-08 1.834148550742089 2.0693e-08 1.7226228579430594 2.0694e-08 1.7583705775514011 2.0695e-08 1.7559667263673433 2.0696e-08 1.7876273483008465 2.0697e-08 1.7794744521279817 2.0698e-08 1.7969354079385094 2.0699e-08 1.8289443363059943 2.07e-08 1.8349004187705127 2.0701e-08 1.8313534863483447 2.0702e-08 1.7405915536758751 2.0703e-08 1.8263989168045986 2.0703999999999998e-08 1.7674930159417923 2.0705e-08 1.759935957710926 2.0706e-08 1.8997250801290058 2.0706999999999998e-08 1.8536522392157349 2.0708e-08 1.8148444117301885 2.0709e-08 1.8436698669338558 2.0709999999999998e-08 1.7681933142550699 2.0711e-08 1.786673775530094 2.0712e-08 1.7736966251426942 2.0712999999999998e-08 1.7907577301901516 2.0714e-08 1.7344407227066403 2.0715e-08 1.90072443699318 2.0716e-08 1.729726264855029 2.0717e-08 1.7601278456580438 2.0718e-08 1.895354998814176 2.0719e-08 1.81348588207751 2.072e-08 1.8164076384698862 2.0721e-08 1.8566159680607102 2.0722e-08 1.8870021971066255 2.0723e-08 1.6964943539127422 2.0724e-08 1.8400113040944144 2.0725e-08 1.8376656870443215 2.0726e-08 1.7986749429220914 2.0727e-08 1.8265543107051432 2.0728e-08 1.7864035536987104 2.0729e-08 1.8279721620940865 2.073e-08 1.7358513839557121 2.0731e-08 1.8081825538586378 2.0732e-08 1.761647575772251 2.0733e-08 1.7943006036099576 2.0734e-08 1.8077690635993062 2.0735e-08 1.7611815567124254 2.0736e-08 1.8362866905556245 2.0737e-08 1.7570016357218414 2.0738e-08 1.7813189742492697 2.0738999999999998e-08 1.7510865259437471 2.074e-08 1.8118945256796597 2.0741e-08 1.7391426247954531 2.0741999999999998e-08 1.7536974477023006 2.0743e-08 1.7446146888229779 2.0744e-08 1.7655765298247161 2.0744999999999998e-08 1.7582421672374484 2.0746e-08 1.8342832654082992 2.0747e-08 1.8435635970944517 2.0747999999999998e-08 1.8111916816542468 2.0749e-08 1.789623292991279 2.075e-08 1.7563901167789462 2.0750999999999998e-08 1.7870188556214452 2.0752e-08 1.7683561442710172 2.0753e-08 1.7459636767459896 2.0754e-08 1.7757216387305537 2.0755e-08 1.8547490609063984 2.0756e-08 1.7837065185740197 2.0757e-08 1.848304753773148 2.0758e-08 1.8268869897700506 2.0759e-08 1.7853919146681752 2.076e-08 1.839221124144021 2.0761e-08 1.8024449047309772 2.0762e-08 1.8114008667270738 2.0763e-08 1.8287687765142329 2.0764e-08 1.805309050624091 2.0765e-08 1.8517601529207826 2.0766e-08 1.8384893120108354 2.0767e-08 1.762631784194418 2.0768e-08 1.7441590689473991 2.0769e-08 1.7753513898055886 2.077e-08 1.7541096580979274 2.0771e-08 1.734001182918052 2.0772e-08 1.799215982898163 2.0773e-08 1.7856908174875923 2.0773999999999998e-08 1.7341237894844976 2.0775e-08 1.8378814604307236 2.0776e-08 1.8338684343624823 2.0776999999999998e-08 1.706204864743221 2.0778e-08 1.770416662032043 2.0779e-08 1.7498296559501103 2.0779999999999998e-08 1.7676505659009007 2.0781e-08 1.8358750405472182 2.0782e-08 1.8348653225600529 2.0782999999999998e-08 1.7824965473599386 2.0784e-08 1.7758678723836723 2.0785e-08 1.794900408648655 2.0785999999999998e-08 1.746220283257397 2.0787e-08 1.7982192491267601 2.0788e-08 1.9414861182941623 2.0789e-08 1.7955740277750174 2.079e-08 1.8305008193120857 2.0791e-08 1.7475446506546364 2.0792e-08 1.8485049810926444 2.0793e-08 1.8501477225129965 2.0794e-08 1.8952053488491274 2.0795e-08 1.762172673714322 2.0796e-08 1.8220543687059636 2.0797e-08 1.7767350726071776 2.0798e-08 1.7901867625639156 2.0799e-08 1.8431667864640928 2.08e-08 1.7533872547441076 2.0801e-08 1.759055229528342 2.0802e-08 1.797061926750324 2.0803e-08 1.7333500784918694 2.0804e-08 1.787030839208526 2.0805e-08 1.7476319173132733 2.0806e-08 1.7454571958671723 2.0807e-08 1.8053648509578626 2.0808e-08 1.8168002189261339 2.0808999999999998e-08 1.848904125472238 2.081e-08 1.8235568974725973 2.0811e-08 1.7202476209433901 2.0811999999999998e-08 1.8134930987928712 2.0813e-08 1.809880682918761 2.0814e-08 1.857953275359299 2.0814999999999998e-08 1.7856635708856397 2.0816e-08 1.7833278111074504 2.0817e-08 1.8162067622381903 2.0817999999999998e-08 1.8390631054495938 2.0819e-08 1.7705249328473431 2.082e-08 1.791421473148391 2.0820999999999998e-08 1.7697206354116344 2.0822e-08 1.7630055527765283 2.0823e-08 1.8375133015787244 2.0824e-08 1.8535171830430914 2.0825e-08 1.7745010432428918 2.0826e-08 1.8294470897107762 2.0827e-08 1.879556752131949 2.0828e-08 1.8989465316150984 2.0829e-08 1.783780168297071 2.083e-08 1.659044241181158 2.0831e-08 1.7209486678615835 2.0832e-08 1.7802315738270813 2.0833e-08 1.8125555588465871 2.0834e-08 1.800733572186228 2.0835e-08 1.8882398894224914 2.0836e-08 1.7798166428632105 2.0837e-08 1.7891195856362745 2.0838e-08 1.7974666984601797 2.0839e-08 1.729627181902043 2.084e-08 1.8607140861123843 2.0841e-08 1.8440478310793686 2.0842e-08 1.8112953268819887 2.0843e-08 1.792605223790549 2.0844e-08 1.8576687864746855 2.0845e-08 1.8447341686767746 2.0846e-08 1.7342550901099256 2.0846999999999998e-08 1.8659462189911897 2.0848e-08 1.7100599123322584 2.0849e-08 1.7986170862708748 2.0849999999999998e-08 1.8014239520544308 2.0851e-08 1.7918860871414353 2.0852e-08 1.7603041610828634 2.0852999999999998e-08 1.8053773210711985 2.0854e-08 1.7800031162950238 2.0855e-08 1.8583517789452262 2.0855999999999998e-08 1.7384598206511532 2.0857e-08 1.741161502025142 2.0858e-08 1.8248908283471545 2.0859e-08 1.7763974189859209 2.086e-08 1.7537950648402312 2.0861e-08 1.88304256675388 2.0862e-08 1.752567738748848 2.0863e-08 1.6610317881899608 2.0864e-08 1.8042045436571743 2.0865e-08 1.745694835847648 2.0866e-08 1.7569568980186219 2.0867e-08 1.825171199884775 2.0868e-08 1.7367803370364703 2.0869e-08 1.8192116955488487 2.087e-08 1.785934357204978 2.0871e-08 1.7489445241888182 2.0872e-08 1.7915247996936068 2.0873e-08 1.7437711759645085 2.0874e-08 1.8536031928558643 2.0875e-08 1.6785067410767989 2.0876e-08 1.7374296501322293 2.0877e-08 1.728327273358663 2.0878e-08 1.6857709909664815 2.0879e-08 1.7422206579892656 2.088e-08 1.8077199854103199 2.0881e-08 1.8830758295679955 2.0881999999999998e-08 1.7227737218083665 2.0883e-08 1.8020599321517918 2.0884e-08 1.723917300325691 2.0884999999999998e-08 1.7873308681165578 2.0886e-08 1.804809814834696 2.0887e-08 1.8099550199476377 2.0887999999999998e-08 1.7676806774083558 2.0889e-08 1.8606988436280787 2.089e-08 1.8620274739572944 2.0890999999999998e-08 1.7791788106125745 2.0892e-08 1.8323902948550659 2.0893e-08 1.8227291830244423 2.0894e-08 1.743481911232926 2.0895e-08 1.8882876382531015 2.0896e-08 1.7276282542616717 2.0897e-08 1.765493170631224 2.0898e-08 1.8241012051789265 2.0899e-08 1.8331047182222775 2.09e-08 1.7567847384749435 2.0901e-08 1.798585082364694 2.0902e-08 1.7629431471560337 2.0903e-08 1.7630985628017708 2.0904e-08 1.7871224274550173 2.0905e-08 1.8359660518041576 2.0906e-08 1.9634911994536737 2.0907e-08 1.7898474292938882 2.0908e-08 1.8157339139792614 2.0909e-08 1.7733926104085227 2.091e-08 1.8237714073663391 2.0911e-08 1.8190489007275144 2.0912e-08 1.8660368940015541 2.0913e-08 1.8203604054779257 2.0914e-08 1.6853773781888508 2.0915e-08 1.8142158442301641 2.0916e-08 1.8201477583454682 2.0916999999999998e-08 1.7614969005892778 2.0918e-08 1.7899514130820917 2.0919e-08 1.710642548331721 2.0919999999999998e-08 1.7858583633380838 2.0921e-08 1.7791189126229765 2.0922e-08 1.8080330069435548 2.0922999999999998e-08 1.906018784519405 2.0924e-08 1.8894345315835506 2.0925e-08 1.8078719440342685 2.0925999999999998e-08 1.8099228062147343 2.0927e-08 1.8426711263154691 2.0928e-08 1.838874696115883 2.0929e-08 1.8396958266100025 2.093e-08 1.872777853053006 2.0931e-08 1.8023159413202194 2.0932e-08 1.7588212518887685 2.0933e-08 1.7476398886972861 2.0934e-08 1.8934847895916922 2.0935e-08 1.7882792995176442 2.0936e-08 1.7187071024257157 2.0937e-08 1.785340443748086 2.0938e-08 1.8929107874117417 2.0939e-08 1.7853486716938771 2.094e-08 1.882370504012728 2.0941e-08 1.8216187799319878 2.0942e-08 1.7187470818807453 2.0943e-08 1.8160494284691278 2.0944e-08 1.7425868951541563 2.0945e-08 1.9069594642092678 2.0946e-08 1.762570290055352 2.0947e-08 1.7869331838791604 2.0948e-08 1.7168009662496428 2.0949e-08 1.7905463968807547 2.095e-08 1.8207286412125157 2.0951e-08 1.8646569450494854 2.0951999999999998e-08 1.791266280558133 2.0953e-08 1.7287413033447065 2.0954e-08 1.7347177174333817 2.0954999999999998e-08 1.7903817812104101 2.0956e-08 1.730549514301717 2.0957e-08 1.8313523576515434 2.0957999999999998e-08 1.7973743792651369 2.0959e-08 1.7702103358399846 2.096e-08 1.7545010357661814 2.0960999999999998e-08 1.790728581049719 2.0962e-08 1.6999083383919884 2.0963e-08 1.8317220189683856 2.0963999999999998e-08 1.8212316821597483 2.0965e-08 1.7211685792659004 2.0966e-08 1.8706805981018653 2.0967e-08 1.7265602192042802 2.0968e-08 1.8738098516654518 2.0969e-08 1.771965292738301 2.097e-08 1.7986365522245173 2.0971e-08 1.7441145007225054 2.0972e-08 1.798929464219319 2.0973e-08 1.7672147207788904 2.0974e-08 1.6909692362390298 2.0975e-08 1.8396672003848076 2.0976e-08 1.7781125064948071 2.0977e-08 1.6765791094047928 2.0978e-08 1.8703750530002665 2.0979e-08 1.7389377292490484 2.098e-08 1.8087289581645767 2.0981e-08 1.8569249113270943 2.0982e-08 1.8783057195758976 2.0983e-08 1.7781790222762497 2.0984e-08 1.7868725192722466 2.0985e-08 1.784698354591584 2.0986e-08 1.7457242910637834 2.0986999999999998e-08 1.876734555217658 2.0988e-08 1.7322366281717014 2.0989e-08 1.8920871305271774 2.0989999999999998e-08 1.79844287258051 2.0991e-08 1.801926305164071 2.0992e-08 1.8637945377625251 2.0992999999999998e-08 1.8298050050571217 2.0994e-08 1.8123282340399562 2.0995e-08 1.7632899676728389 2.0995999999999998e-08 1.7704599531642662 2.0997e-08 1.7993376247944486 2.0998e-08 1.7712717863524063 2.0998999999999998e-08 1.7313288027840263 2.1e-08 1.8143792001676622 2.1001e-08 1.773251986191656 2.1002e-08 1.7310661311627595 2.1003e-08 1.8638612847744866 2.1004e-08 1.859278659729032 2.1005e-08 1.8646628988995317 2.1006e-08 1.7968666704627199 2.1007e-08 1.8325749894993775 2.1008e-08 1.7863515072306824 2.1009e-08 1.8171757096047034 2.101e-08 1.856610123942087 2.1011e-08 1.8413286486418128 2.1012e-08 1.833468056985666 2.1013e-08 1.8287610655582247 2.1014e-08 1.7467289648849964 2.1015e-08 1.7700465843966633 2.1016e-08 1.785571766366269 2.1017e-08 1.7605952300633383 2.1018e-08 1.8107538349222272 2.1019e-08 1.8371869232248839 2.102e-08 1.8328139549490576 2.1021e-08 1.8718599825676776 2.1021999999999998e-08 1.7748364894372903 2.1023e-08 1.792716076808026 2.1024e-08 1.7639008077825349 2.1024999999999998e-08 1.749008458387092 2.1026e-08 1.8510240504219853 2.1027e-08 1.7254149879146383 2.1027999999999998e-08 1.7596054293941699 2.1029e-08 1.7586801650307842 2.103e-08 1.7641743108814347 2.1030999999999998e-08 1.6797921884189373 2.1032e-08 1.8476044840396475 2.1033e-08 1.7438158392549603 2.1033999999999998e-08 1.811570565963447 2.1035e-08 1.8040939506311324 2.1036e-08 1.7286935412758926 2.1037e-08 1.7627753458570201 2.1038e-08 1.807652163950614 2.1039e-08 1.780309050325322 2.104e-08 1.7897256895266684 2.1041e-08 1.8683268324181146 2.1042e-08 1.809941932785257 2.1043e-08 1.7764126637353816 2.1044e-08 1.8300851436896235 2.1045e-08 1.786202948844697 2.1046e-08 1.8604252691392864 2.1047e-08 1.728921542264276 2.1048e-08 1.8169401296442724 2.1049e-08 1.751761259669118 2.105e-08 1.8333273975804476 2.1051e-08 1.8360283449149373 2.1052e-08 1.819367370245944 2.1053e-08 1.835278730595608 2.1054e-08 1.8382791831583116 2.1055e-08 1.7864161733754111 2.1056e-08 1.8178764111179953 2.1057e-08 1.880594695391182 2.1058e-08 1.789719639495021 2.1059e-08 1.7776540179265623 2.1059999999999998e-08 1.8404897386394532 2.1061e-08 1.840150654919608 2.1062e-08 1.7482365596603504 2.1062999999999998e-08 1.7745364736998221 2.1064e-08 1.862119208864304 2.1065e-08 1.8011551206917622 2.1065999999999998e-08 1.932518791235475 2.1067e-08 1.8437567182841457 2.1068e-08 1.8234213521983245 2.1068999999999998e-08 1.8236856386479359 2.107e-08 1.8257908441276842 2.1071e-08 1.7910449137138233 2.1072e-08 1.7525697531253301 2.1073e-08 1.7245703341896206 2.1074e-08 1.9144042852335263 2.1075e-08 1.767359846141141 2.1076e-08 1.8360344928692482 2.1077e-08 1.7602670847021618 2.1078e-08 1.8530435682828146 2.1079e-08 1.8607119968553432 2.108e-08 1.8196265979708772 2.1081e-08 1.7969124999668737 2.1082e-08 1.708711985330951 2.1083e-08 1.7590522795890253 2.1084e-08 1.8279313232893362 2.1085e-08 1.779827411165422 2.1086e-08 1.7587678806674152 2.1087e-08 1.8126976606959924 2.1088e-08 1.7550413041376791 2.1089e-08 1.8419696725102777 2.109e-08 1.7649969029782713 2.1091e-08 1.8279177710693397 2.1092e-08 1.7708134725441729 2.1093e-08 1.7749293184773915 2.1094e-08 1.7711904726764 2.1094999999999998e-08 1.8313514260382255 2.1096e-08 1.7723938266439672 2.1097e-08 1.7638635290709455 2.1097999999999998e-08 1.764088790568843 2.1099e-08 1.784677526514024 2.11e-08 1.6969800024337738 2.1100999999999998e-08 1.7116398015198566 2.1102e-08 1.909302931050643 2.1103e-08 1.7190198108884578 2.1103999999999998e-08 1.7732973562212828 2.1105e-08 1.8113209844777292 2.1106e-08 1.7967094808610975 2.1107e-08 1.7562489870862208 2.1108e-08 1.7906963159015654 2.1109e-08 1.7353765491180864 2.111e-08 1.8684522816995897 2.1111e-08 1.7479185130751285 2.1112e-08 1.7742847441648484 2.1113e-08 1.803699133129096 2.1114e-08 1.8558054348434299 2.1115e-08 1.8287798121506995 2.1116e-08 1.8158286515027942 2.1117e-08 1.9249669058157013 2.1118e-08 1.719706738756011 2.1119e-08 1.7660116256060425 2.112e-08 1.8137146324060265 2.1121e-08 1.7680670809316823 2.1122e-08 1.875032997873541 2.1123e-08 1.8232591349765073 2.1124e-08 1.7679436715903527 2.1125e-08 1.801890504436158 2.1126e-08 1.6993554275028702 2.1127e-08 1.7625389869669177 2.1128e-08 1.8481305306379776 2.1129e-08 1.771590134788661 2.1129999999999998e-08 1.7932170247734556 2.1131e-08 1.7864339258766162 2.1132e-08 1.8321422623034336 2.1132999999999998e-08 1.7863430854492535 2.1134e-08 1.7276923987600215 2.1135e-08 1.7774592148686423 2.1135999999999998e-08 1.8010170638758727 2.1137e-08 1.8097861735164313 2.1138e-08 1.7793284043477755 2.1138999999999998e-08 1.7715479116487334 2.114e-08 1.8718486771983467 2.1141e-08 1.8023802426158626 2.1141999999999998e-08 1.8535793579029027 2.1143e-08 1.8797889393039595 2.1144e-08 1.8095619531129667 2.1145e-08 1.7383918554092261 2.1146e-08 1.7956079854681448 2.1147e-08 1.7448401392640536 2.1148e-08 1.9094641312479497 2.1149e-08 1.771462101800094 2.115e-08 1.8609816863359203 2.1151e-08 1.7469821918781305 2.1152e-08 1.764015565921526 2.1153e-08 1.8825383107865152 2.1154e-08 1.8443865397580934 2.1155e-08 1.743774404464124 2.1156e-08 1.7807490678563729 2.1157e-08 1.9294519948385211 2.1158e-08 1.8330777704583687 2.1159e-08 1.8009123960818767 2.116e-08 1.7353710163764273 2.1161e-08 1.8289534434042767 2.1162e-08 1.7428922077571072 2.1163e-08 1.7703898626296677 2.1164e-08 1.7919327156597298 2.1164999999999998e-08 1.8599126321428499 2.1166e-08 1.786783493440152 2.1167e-08 1.8224083941030014 2.1167999999999998e-08 1.7913984709770592 2.1169e-08 1.7401319289286534 2.117e-08 1.7730637101649904 2.1170999999999998e-08 1.8582309263407981 2.1172e-08 1.7815538910203434 2.1173e-08 1.8095250434810293 2.1173999999999998e-08 1.770948351026862 2.1175e-08 1.791876650164239 2.1176e-08 1.780388056476071 2.1176999999999998e-08 1.921929624177017 2.1178e-08 1.7553512634845088 2.1179e-08 1.830166035418215 2.118e-08 1.8911104919846422 2.1181e-08 1.8491908572819609 2.1182e-08 1.8358201861020786 2.1183e-08 1.7209802194745212 2.1184e-08 1.7346351278437384 2.1185e-08 1.764527540567557 2.1186e-08 1.755118800757087 2.1187e-08 1.720852576686752 2.1188e-08 1.7403386927016595 2.1189e-08 1.837747268451172 2.119e-08 1.8683632063745887 2.1191e-08 1.845014254163866 2.1192e-08 1.833271203307989 2.1193e-08 1.78705021759357 2.1194e-08 1.8163626244842757 2.1195e-08 1.7548181750422964 2.1196e-08 1.7248489711295465 2.1197e-08 1.8753396306249275 2.1198e-08 1.8607522671040762 2.1199e-08 1.7374253701827094 2.1199999999999998e-08 1.831857214492099 2.1201e-08 1.8126636541994892 2.1202e-08 1.8676557631941022 2.1202999999999998e-08 1.6861350835673519 2.1204e-08 1.9010856651731591 2.1205e-08 1.7819863918025332 2.1205999999999998e-08 1.8448134646315713 2.1207e-08 1.8573343291952402 2.1208e-08 1.9018127283721598 2.1208999999999998e-08 1.7488834668666264 2.121e-08 1.8326666869665909 2.1211e-08 1.8108718282313256 2.1211999999999998e-08 1.7985661865073754 2.1213e-08 1.8189872378333967 2.1214e-08 1.8295821659549354 2.1215e-08 1.7070336188949014 2.1216e-08 1.7387315968453885 2.1217e-08 1.7724248464134402 2.1218e-08 1.7124393449455055 2.1219e-08 1.8085656587489316 2.122e-08 1.8157374435142197 2.1221e-08 1.666628817435466 2.1222e-08 1.786203406934311 2.1223e-08 1.8666674321198855 2.1224e-08 1.8060313105563006 2.1225e-08 1.7699685119102715 2.1226e-08 1.8232226858005887 2.1227e-08 1.8194416892269567 2.1228e-08 1.855434892821183 2.1229e-08 1.8539362063180727 2.123e-08 1.7627267891203573 2.1231e-08 1.8650609283481336 2.1232e-08 1.7055880362918678 2.1233e-08 1.9097879707189995 2.1234e-08 1.8135291573195338 2.1235e-08 1.7668965280971494 2.1236e-08 1.74177881007441 2.1237e-08 1.7795781764824223 2.1237999999999998e-08 1.8171930720390896 2.1239e-08 1.853556934990972 2.124e-08 1.8192068198765976 2.1240999999999998e-08 1.7598646811859227 2.1242e-08 1.7788933169584713 2.1243e-08 1.7970233488242933 2.1243999999999998e-08 1.8189988731402593 2.1245e-08 1.8263466590453927 2.1246e-08 1.7996316250041937 2.1246999999999998e-08 1.8104301119964745 2.1248e-08 1.7336058874347235 2.1249e-08 1.760532854628928 2.125e-08 1.7471907597241885 2.1251e-08 1.8274888394709434 2.1252e-08 1.8275137867087143 2.1253e-08 1.753840847225956 2.1254e-08 1.7435089598645874 2.1255e-08 1.8397531312000197 2.1256e-08 1.864812519138929 2.1257e-08 1.8430921848469164 2.1258e-08 1.8610970938160205 2.1259e-08 1.8766406891133256 2.126e-08 1.7970067934026617 2.1261e-08 1.8083908611533006 2.1262e-08 1.7793443032778136 2.1263e-08 1.8183262763706858 2.1264e-08 1.7705086587105587 2.1265e-08 1.7125297762386054 2.1266e-08 1.7518498710231019 2.1267e-08 1.8960694788139847 2.1268e-08 1.7742660936359218 2.1269e-08 1.8394343814216514 2.127e-08 1.7471825807576349 2.1271e-08 1.7575634107084803 2.1272e-08 1.86211427045831 2.1272999999999998e-08 1.8047736227448532 2.1274e-08 1.734591654743968 2.1275e-08 1.8144853637683789 2.1275999999999998e-08 1.8929942944233928 2.1277e-08 1.8451927565379858 2.1278e-08 1.867168174873795 2.1278999999999998e-08 1.8024574511822289 2.128e-08 1.8636300082860349 2.1281e-08 1.7799613088026298 2.1281999999999998e-08 1.7560476596388825 2.1283e-08 1.7909991787495338 2.1284e-08 1.7039870185349257 2.1285e-08 1.824926026239946 2.1286e-08 1.7542824410020588 2.1287e-08 1.8094560757504154 2.1288e-08 1.761448989654885 2.1289e-08 1.919092338664289 2.129e-08 1.8335704755164524 2.1291e-08 1.750354172879255 2.1292e-08 1.8002911810266122 2.1293e-08 1.7805404095030641 2.1294e-08 1.819019613116605 2.1295e-08 1.7550360162145167 2.1296e-08 1.7744539175054004 2.1297e-08 1.7747270622086617 2.1298e-08 1.771656065624386 2.1299e-08 1.5876511302361904 2.13e-08 1.7384284801362426 2.1301e-08 1.880833349665905 2.1302e-08 1.769147199712587 2.1303e-08 1.8019364052638844 2.1304e-08 1.8495250347618817 2.1305e-08 1.8455412158858897 2.1306e-08 1.820044802318858 2.1307e-08 1.7766849623474186 2.1307999999999998e-08 1.773353643165351 2.1309e-08 1.8565488813776907 2.131e-08 1.8004341822571488 2.1310999999999998e-08 1.8281018897358174 2.1312e-08 1.7923190349446143 2.1313e-08 1.7817855572858334 2.1313999999999998e-08 1.7460216428331403 2.1315e-08 1.849323312047109 2.1316e-08 1.735562645334616 2.1316999999999998e-08 1.8036975413588192 2.1318e-08 1.733014529386913 2.1319e-08 1.7917543013360384 2.1319999999999998e-08 1.8555901717077197 2.1321e-08 1.7669696576349425 2.1322e-08 1.7297962415036934 2.1323e-08 1.7937700981454223 2.1324e-08 1.7718088301845152 2.1325e-08 1.7881409340931802 2.1326e-08 1.7648223458832468 2.1327e-08 1.774685461204924 2.1328e-08 1.744767014741278 2.1329e-08 1.7867049720916361 2.133e-08 1.7962636107537968 2.1331e-08 1.8245359758874893 2.1332e-08 1.7362011969543711 2.1333e-08 1.7821972274377185 2.1334e-08 1.7237480751808962 2.1335e-08 1.7676245401015103 2.1336e-08 1.8604403552271003 2.1337e-08 1.792978777272222 2.1338e-08 1.7386252475481625 2.1339e-08 1.8243348474803314 2.134e-08 1.8365636461849635 2.1341e-08 1.8259093049131436 2.1342e-08 1.7415844440315522 2.1342999999999998e-08 1.803624374992595 2.1344e-08 1.7498245800608117 2.1345e-08 1.771221888524836 2.1345999999999998e-08 1.6826048612060507 2.1347e-08 1.7773189984413416 2.1348e-08 1.7161706976534077 2.1348999999999998e-08 1.7952130751733217 2.135e-08 1.7928391034821454 2.1351e-08 1.709996887610689 2.1351999999999998e-08 1.7564807236717122 2.1353e-08 1.8370819954021163 2.1354e-08 1.8011091790139035 2.1354999999999998e-08 1.7786329847466729 2.1356e-08 1.8275487558969623 2.1357e-08 1.7196290908698721 2.1358e-08 1.8346138327903239 2.1359e-08 1.8324530811973778 2.136e-08 1.7396835292000628 2.1361e-08 1.7748026251922107 2.1362e-08 1.823267789091869 2.1363e-08 1.8431500906455112 2.1364e-08 1.8228640351391714 2.1365e-08 1.819246167578432 2.1366e-08 1.920221107995196 2.1367e-08 1.8656698512416376 2.1368e-08 1.792000694653849 2.1369e-08 1.814173881903472 2.137e-08 1.8027264256039917 2.1371e-08 1.8825163696924425 2.1372e-08 1.8409473158202756 2.1373e-08 1.8704646061155037 2.1374e-08 1.7417235411744971 2.1375e-08 1.8086316848271142 2.1376e-08 1.7657034003915537 2.1377e-08 1.749687317737644 2.1377999999999998e-08 1.7920361812178536 2.1379e-08 1.8783226446287933 2.138e-08 1.7362442562822962 2.1380999999999998e-08 1.7347536424645094 2.1382e-08 1.8484544272777428 2.1383e-08 1.845222584631576 2.1383999999999998e-08 1.7932861385924843 2.1385e-08 1.8188695995555029 2.1386e-08 1.8220211754166105 2.1386999999999998e-08 1.8236490136393642 2.1388e-08 1.7192585166094472 2.1389e-08 1.847191583475165 2.1389999999999998e-08 1.8721516582113944 2.1391e-08 1.7547614903182487 2.1392e-08 1.8048949289727194 2.1393e-08 1.8388866131389165 2.1394e-08 1.7212997573416797 2.1395e-08 1.764981806415665 2.1396e-08 1.8141908158790467 2.1397e-08 1.861767096717463 2.1398e-08 1.8639384361522737 2.1399e-08 1.7704308173808005 2.14e-08 1.8191552790818195 2.1401e-08 1.7024928978564282 2.1402e-08 1.7932874339630132 2.1403e-08 1.8398773133937285 2.1404e-08 1.8451148582335264 2.1405e-08 1.7566991022421012 2.1406e-08 1.834703360622553 2.1407e-08 1.8985018331459353 2.1408e-08 1.846923104495341 2.1409e-08 1.7784172520763184 2.141e-08 1.856390945617226 2.1411e-08 1.8200784815471545 2.1412e-08 1.8165001758995587 2.1412999999999998e-08 1.8374676723675154 2.1414e-08 1.7222035182683664 2.1415e-08 1.822489993686958 2.1415999999999998e-08 1.7622812287570693 2.1417e-08 1.7870619629246742 2.1418e-08 1.8421224112981371 2.1418999999999998e-08 1.8320176180462437 2.142e-08 1.7806066893072203 2.1421e-08 1.8012417950046242 2.1421999999999998e-08 1.6601641868233301 2.1423e-08 1.8314932319453507 2.1424e-08 1.72377063314657 2.1424999999999998e-08 1.744661188858926 2.1426e-08 1.7552074328088394 2.1427e-08 1.772591375212075 2.1428e-08 1.8280572481837987 2.1429e-08 1.8431246287504384 2.143e-08 1.866666197280214 2.1431e-08 1.8529986113139851 2.1432e-08 1.7815678717763812 2.1433e-08 1.8762809469247483 2.1434e-08 1.885919317725871 2.1435e-08 1.8360720351553161 2.1436e-08 1.8203837842981685 2.1437e-08 1.8032089170232155 2.1438e-08 1.8582031853424061 2.1439e-08 1.8262823918966233 2.144e-08 1.8100716488040784 2.1441e-08 1.849402432302822 2.1442e-08 1.8211458298281795 2.1443e-08 1.7789771296914099 2.1444e-08 1.8911815155846887 2.1445e-08 1.8507038750488878 2.1446e-08 1.7017308126113349 2.1447e-08 1.7762486795431547 2.1448e-08 1.844698472279334 2.1449e-08 1.7774561397568813 2.145e-08 1.7567871855682093 2.1450999999999998e-08 1.7525086766978348 2.1452e-08 1.8504500351113804 2.1453e-08 1.763456527236733 2.1453999999999998e-08 1.8544836093034758 2.1455e-08 1.8488078884144243 2.1456e-08 1.7914653479879976 2.1456999999999998e-08 1.735061017197667 2.1458e-08 1.8637833987382044 2.1459e-08 1.7583621176948343 2.1459999999999998e-08 1.830083887482401 2.1461e-08 1.8694857043597515 2.1462e-08 1.8388636713212974 2.1463e-08 1.7478947327029672 2.1464e-08 1.8103887657776834 2.1465e-08 1.7546769141876044 2.1466e-08 1.7349826043627237 2.1467e-08 1.8800005238707187 2.1468e-08 1.7740347517371287 2.1469e-08 1.8876502380013958 2.147e-08 1.79136612968805 2.1471e-08 1.8027957343470709 2.1472e-08 1.7637985322147827 2.1473e-08 1.8063084707107728 2.1474e-08 1.8042506917483574 2.1475e-08 1.7526516709564401 2.1476e-08 1.8094420140031784 2.1477e-08 1.87389656622336 2.1478e-08 1.8148032878550708 2.1479e-08 1.8141590131817094 2.148e-08 1.7857888138803337 2.1481e-08 1.7634639776399916 2.1482e-08 1.8140615136177929 2.1483e-08 1.8012827014637234 2.1484e-08 1.8193126042198209 2.1485e-08 1.7189964376449032 2.1485999999999998e-08 1.7770502821778107 2.1487e-08 1.7471668946180372 2.1488e-08 1.8125526914044856 2.1488999999999998e-08 1.741593518155728 2.149e-08 1.7573641643262077 2.1491e-08 1.7651749589869403 2.1491999999999998e-08 1.7604003645712583 2.1493e-08 1.8262411399938383 2.1494e-08 1.725539377419924 2.1494999999999998e-08 1.8809500857658907 2.1496e-08 1.829175118797979 2.1497e-08 1.799751610224892 2.1498e-08 1.688567540649342 2.1499e-08 1.887945553945412 2.15e-08 1.8394478010990567 2.1501e-08 1.9118541274912673 2.1502e-08 1.809279024848699 2.1503e-08 1.8164962121402892 2.1504e-08 1.83181644505201 2.1505e-08 1.8383875582310867 2.1506e-08 1.7845113839412343 2.1507e-08 1.8260580636647936 2.1508e-08 1.813031704351605 2.1509e-08 1.7900133427299447 2.151e-08 1.8731049066327854 2.1511e-08 1.828665751630226 2.1512e-08 1.7338986543331953 2.1513e-08 1.812005572933372 2.1514e-08 1.735575633418294 2.1515e-08 1.8018968969335911 2.1516e-08 1.7939882380391692 2.1517e-08 1.8569315734359313 2.1518e-08 1.8003311733425813 2.1519e-08 1.8278627578041977 2.152e-08 1.7634470667094522 2.1520999999999998e-08 1.7225278598896412 2.1522e-08 1.759611247505868 2.1523e-08 1.765260474132764 2.1523999999999998e-08 1.9105492027944209 2.1525e-08 1.8360640707344902 2.1526e-08 1.806678335334624 2.1526999999999998e-08 1.6810001626729059 2.1528e-08 1.7818606298669133 2.1529e-08 1.859097729863615 2.1529999999999998e-08 1.7640904244115136 2.1531e-08 1.798211230717272 2.1532e-08 1.8423128828243813 2.1532999999999998e-08 1.9280501285077734 2.1534e-08 1.8555535761020647 2.1535e-08 1.847507821421127 2.1536e-08 1.7980718669643776 2.1537e-08 1.8512594783246583 2.1538e-08 1.800336850462856 2.1539e-08 1.8058478710716888 2.154e-08 1.8473234593136552 2.1541e-08 1.8122111250830992 2.1542e-08 1.8087736204429998 2.1543e-08 1.7659458667811059 2.1544e-08 1.812899038868967 2.1545e-08 1.7832781360736714 2.1546e-08 1.8275367816555572 2.1547e-08 1.7588176329460323 2.1548e-08 1.7318055268737176 2.1549e-08 1.8156539841935544 2.155e-08 1.8053567054837634 2.1551e-08 1.8276579447167238 2.1552e-08 1.8343555026097662 2.1553e-08 1.839570628821045 2.1554e-08 1.8718202661494936 2.1555e-08 1.73321946598944 2.1555999999999998e-08 1.7950051535829543 2.1557e-08 1.7847374619105065 2.1558e-08 1.7454146362502636 2.1558999999999998e-08 1.7636779748753564 2.156e-08 1.796239712012025 2.1561e-08 1.7866646863317246 2.1561999999999998e-08 1.8088581026676664 2.1563e-08 1.7992466611313553 2.1564e-08 1.8340128814666061 2.1564999999999998e-08 1.8224672136898707 2.1566e-08 1.720746953526596 2.1567e-08 1.8001980078846949 2.1567999999999998e-08 1.8518798798669636 2.1569e-08 1.7021943697982715 2.157e-08 1.7593626731950904 2.1571e-08 1.789955313140027 2.1572e-08 1.7574863578622806 2.1573e-08 1.8400552294354493 2.1574e-08 1.8318204466173198 2.1575e-08 1.794024520959986 2.1576e-08 1.7917903120012257 2.1577e-08 1.864562225757889 2.1578e-08 1.8392813783451534 2.1579e-08 1.9352259700101864 2.158e-08 1.874187691586379 2.1581e-08 1.8286861007122766 2.1582e-08 1.7822858869512335 2.1583e-08 1.8582661286034208 2.1584e-08 1.7660405465585216 2.1585e-08 1.8157725634753858 2.1586e-08 1.743087980725894 2.1587e-08 1.7553627238557974 2.1588e-08 1.6951076575743163 2.1589e-08 1.9045131942869153 2.159e-08 1.7130698483473463 2.1590999999999998e-08 1.7971503822471353 2.1592e-08 1.7461501466761746 2.1593e-08 1.7420552413578125 2.1593999999999998e-08 1.8251265571227226 2.1595e-08 1.8354753278691325 2.1596e-08 1.843269558579029 2.1596999999999998e-08 1.8326481213853607 2.1598e-08 1.7318129315921806 2.1599e-08 1.839818794142096 2.1599999999999998e-08 1.7920100679747928 2.1601e-08 1.7678409958882306 2.1602e-08 1.8129300461790776 2.1602999999999998e-08 1.7662801125826766 2.1604e-08 1.8308090126319416 2.1605e-08 1.7630590832598907 2.1606e-08 1.839552117612468 2.1607e-08 1.8155876871813685 2.1608e-08 1.8152647735429712 2.1609e-08 1.847322995368359 2.161e-08 1.7372477706133342 2.1611e-08 1.8220757954994342 2.1612e-08 1.8461056825311466 2.1613e-08 1.8602773141388589 2.1614e-08 1.7310522326791304 2.1615e-08 1.7908301170246386 2.1616e-08 1.6890104625908051 2.1617e-08 1.8406966274148553 2.1618e-08 1.7844104879246319 2.1619e-08 1.686580986494787 2.162e-08 1.7603448179256416 2.1621e-08 1.7831386053213074 2.1622e-08 1.8179626837114429 2.1623e-08 1.7948646274682065 2.1624e-08 1.7159560925013964 2.1625e-08 1.8189311051213872 2.1626e-08 1.7840625932103833 2.1627e-08 1.7737283762018254 2.1628e-08 1.7955211908657045 2.1628999999999998e-08 1.8257960695517574 2.163e-08 1.7076528084473497 2.1631e-08 1.8328332945121455 2.1631999999999998e-08 1.9302848657825944 2.1633e-08 1.816389623379014 2.1634e-08 1.77076165678015 2.1634999999999998e-08 1.7979602601602942 2.1636e-08 1.803382014204757 2.1637e-08 1.7785464883555417 2.1637999999999998e-08 1.7453187707257856 2.1639e-08 1.7697284280673191 2.164e-08 1.8658311124357345 2.1641e-08 1.8404273329823508 2.1642e-08 1.7619516174824705 2.1643e-08 1.8420261434938254 2.1644e-08 1.6615098003502036 2.1645e-08 1.8349338883442414 2.1646e-08 1.8211516854192151 2.1647e-08 1.8015241772694683 2.1648e-08 1.8565181048495156 2.1649e-08 1.789139662533452 2.165e-08 1.804526760051077 2.1651e-08 1.8277299108100737 2.1652e-08 1.7451547642985163 2.1653e-08 1.6924951874219487 2.1654e-08 1.8214660384544201 2.1655e-08 1.8434546084064236 2.1656e-08 1.7306722856179229 2.1657e-08 1.8206764830197888 2.1658e-08 1.8175354226765088 2.1659e-08 1.8284279684159688 2.166e-08 1.7469627634003189 2.1661e-08 1.752470921931625 2.1662e-08 1.7490916884792 2.1663e-08 1.8236524869137334 2.1663999999999998e-08 1.8228416408227646 2.1665e-08 1.6940383120897065 2.1666e-08 1.7540839626674598 2.1666999999999998e-08 1.908322570846836 2.1668e-08 1.8583968401988378 2.1669e-08 1.750879936346225 2.1669999999999998e-08 1.8226003442016956 2.1671e-08 1.6816021536595325 2.1672e-08 1.813648996300568 2.1672999999999998e-08 1.6895254262597212 2.1674e-08 1.8063576825319159 2.1675e-08 1.8335886742408527 2.1676e-08 1.8233291580450082 2.1677e-08 1.8758124221768935 2.1678e-08 1.7723363452381755 2.1679e-08 1.9063980278912172 2.168e-08 1.8175744716501592 2.1681e-08 1.871613466490111 2.1682e-08 1.7721468326287544 2.1683e-08 1.9003724789341827 2.1684e-08 1.7856421221809553 2.1685e-08 1.7618449048255997 2.1686e-08 1.8039175748803629 2.1687e-08 1.743423500717754 2.1688e-08 1.7676000466018194 2.1689e-08 1.8725024404242108 2.169e-08 1.7984902564679879 2.1691e-08 1.807237790892686 2.1692e-08 1.8236654591337877 2.1693e-08 1.8381609903380118 2.1694e-08 1.8067962294567805 2.1695e-08 1.7775364854267752 2.1696e-08 1.8200575477750962 2.1697e-08 1.7576713007028195 2.1698e-08 1.809230740917393 2.1698999999999998e-08 1.8386787102764364 2.17e-08 1.7528026034744018 2.1701e-08 1.8655977214806445 2.1701999999999998e-08 1.7945860795986581 2.1703e-08 1.7237454794588478 2.1704e-08 1.700168876082538 2.1704999999999998e-08 1.8056533661613772 2.1706e-08 1.7267317028264693 2.1707e-08 1.799911319198474 2.1707999999999998e-08 1.7862643716768616 2.1709e-08 1.8256531201395794 2.171e-08 1.8389625502726703 2.1710999999999998e-08 1.853170315276092 2.1712e-08 1.8882048059221828 2.1713e-08 1.8813851709456684 2.1714e-08 1.7834168070717127 2.1715e-08 1.7809457730709264 2.1716e-08 1.872209034750566 2.1717e-08 1.8086249694207326 2.1718e-08 1.728058800100292 2.1719e-08 1.762534987391998 2.172e-08 1.7859376773375868 2.1721e-08 1.772352132630618 2.1722e-08 1.7738231191112264 2.1723e-08 1.8097232875251548 2.1724e-08 1.8432101231311442 2.1725e-08 1.8121381731357453 2.1726e-08 1.7869717465370338 2.1727e-08 1.8919683070779072 2.1728e-08 1.8815660478145142 2.1729e-08 1.7901289710968271 2.173e-08 1.7829313040509032 2.1731e-08 1.794114721108843 2.1732e-08 1.7514177641573276 2.1733e-08 1.8502856301663857 2.1733999999999998e-08 1.8103357301466514 2.1735e-08 1.79673875890402 2.1736e-08 1.7557333448293964 2.1736999999999998e-08 1.7383383227471492 2.1738e-08 1.830942346549568 2.1739e-08 1.7148435275543297 2.1739999999999998e-08 1.7576989078858054 2.1741e-08 1.7988352326469081 2.1742e-08 1.9137037573410345 2.1742999999999998e-08 1.8041885279537107 2.1744e-08 1.8224784356941062 2.1745e-08 1.8065777291057568 2.1745999999999998e-08 1.787374840505707 2.1747e-08 1.7590042138450563 2.1748e-08 1.810444174878639 2.1749e-08 1.7803043088553214 2.175e-08 1.7094196082546644 2.1751e-08 1.6839052048241985 2.1752e-08 1.9056984393816425 2.1753e-08 1.8462337425192292 2.1754e-08 1.887898953140497 2.1755e-08 1.8369798080034996 2.1756e-08 1.8281630259383392 2.1757e-08 1.870195035331341 2.1758e-08 1.7996699566646188 2.1759e-08 1.7394177561267596 2.176e-08 1.8567574185833617 2.1761e-08 1.7756389341729086 2.1762e-08 1.7804473537455225 2.1763e-08 1.8205740724447619 2.1764e-08 1.764091035289333 2.1765e-08 1.843185081849136 2.1766e-08 1.820828498099522 2.1767e-08 1.7976291266401956 2.1768e-08 1.764476088372232 2.1768999999999998e-08 1.8133977183524947 2.177e-08 1.812240266552351 2.1771e-08 1.857384905840027 2.1771999999999998e-08 1.7372221204565974 2.1773e-08 1.8486995093839371 2.1774e-08 1.8536081154701778 2.1774999999999998e-08 1.801695814374757 2.1776e-08 1.9094964863373254 2.1777e-08 1.7932910883692477 2.1777999999999998e-08 1.7872076689091985 2.1779e-08 1.8318384429448928 2.178e-08 1.900907322963611 2.1780999999999998e-08 1.8233773618305513 2.1782e-08 1.793595873505974 2.1783e-08 1.8689856770971471 2.1784e-08 1.7172949850250876 2.1785e-08 1.8440629255144785 2.1786e-08 1.7943617459944912 2.1787e-08 1.7812047491293626 2.1788e-08 1.7882735517880208 2.1789e-08 1.8936050005325882 2.179e-08 1.8029406643810828 2.1791e-08 1.7881815286387208 2.1792e-08 1.7302474288972698 2.1793e-08 1.7667629327052872 2.1794e-08 1.728597470221652 2.1795e-08 1.8909397745807888 2.1796e-08 1.8846031582513678 2.1797e-08 1.8063352308789886 2.1798e-08 1.8497271255503525 2.1799e-08 1.7185677148538019 2.18e-08 1.7471152429349972 2.1801e-08 1.8099076045181217 2.1802e-08 1.7647682441321286 2.1803e-08 1.8501333579526693 2.1803999999999998e-08 1.7525232318981727 2.1805e-08 1.828197361619387 2.1806e-08 1.7243342435783302 2.1806999999999998e-08 1.7733859383176744 2.1808e-08 1.8506226991823003 2.1809e-08 1.8548509250829677 2.1809999999999998e-08 1.8422617669198318 2.1811e-08 1.7643429580645023 2.1812e-08 1.8394546466951474 2.1812999999999998e-08 1.7705299436683024 2.1814e-08 1.8728566618948375 2.1815e-08 1.7945108946708948 2.1815999999999998e-08 1.8161291653328722 2.1817e-08 1.7925385276034937 2.1818e-08 1.7848023413219107 2.1819e-08 1.7463639242797275 2.182e-08 1.8171429195917657 2.1821e-08 1.7920400705268054 2.1822e-08 1.8114844902617397 2.1823e-08 1.8434547806375512 2.1824e-08 1.8753210239737657 2.1825e-08 1.7639803508936331 2.1826e-08 1.755438937200541 2.1827e-08 1.8994026611985764 2.1828e-08 1.780276874792444 2.1829e-08 1.788390849567367 2.183e-08 1.8009934089598951 2.1831e-08 1.8869001505951664 2.1832e-08 1.8261479562987581 2.1833e-08 1.7471996463119612 2.1834e-08 1.7824941970375785 2.1835e-08 1.7241435270359193 2.1836e-08 1.868213754085005 2.1837e-08 1.8555822790521657 2.1838e-08 1.7178262150852694 2.1839e-08 1.8167369929764094 2.184e-08 1.7958628248755373 2.1841e-08 1.8310889399615355 2.1841999999999998e-08 1.8265511518989244 2.1843e-08 1.853216213946296 2.1844e-08 1.791893548223427 2.1844999999999998e-08 1.7774029424516986 2.1846e-08 1.8496567949897196 2.1847e-08 1.7590240122248622 2.1847999999999998e-08 1.8695934680835373 2.1849e-08 1.8040691749474436 2.185e-08 1.7640365778832763 2.1850999999999998e-08 1.8549976773760741 2.1852e-08 1.7900076067360664 2.1853e-08 1.7737287003127384 2.1854e-08 1.8750928310695056 2.1855e-08 1.8545795181537224 2.1856e-08 1.7666855044095053 2.1857e-08 1.7321156858877782 2.1858e-08 1.7335847309434982 2.1859e-08 1.7900512581071881 2.186e-08 1.8071717936816603 2.1861e-08 1.8197121515183088 2.1862e-08 1.7859656278734013 2.1863e-08 1.8143071202831151 2.1864e-08 1.7789776366844454 2.1865e-08 1.785364810787803 2.1866e-08 1.7627045868114335 2.1867e-08 1.8102386942897515 2.1868e-08 1.7450405599248473 2.1869e-08 1.7185095089401226 2.187e-08 1.7905559711068602 2.1871e-08 1.720590092026095 2.1872e-08 1.7968493741576885 2.1873e-08 1.8336642702293724 2.1874e-08 1.8823781851995878 2.1875e-08 1.853492659220901 2.1876e-08 1.8242251109597682 2.1876999999999998e-08 1.8865930737960053 2.1878e-08 1.846549470164328 2.1879e-08 1.7669810843356115 2.1879999999999998e-08 1.7906582106615543 2.1881e-08 1.8620460662220784 2.1882e-08 1.7655118986858962 2.1882999999999998e-08 1.737658418435039 2.1884e-08 1.7046062947062797 2.1885e-08 1.8324003782958833 2.1885999999999998e-08 1.8592921635754003 2.1887e-08 1.8516987969708842 2.1888e-08 1.8536030065630058 2.1888999999999998e-08 1.7795570440333264 2.189e-08 1.7067749785250697 2.1891e-08 1.8614150532346831 2.1892e-08 1.7624832090204066 2.1893e-08 1.8457779966153958 2.1894e-08 1.804934348788432 2.1895e-08 1.8666937764215457 2.1896e-08 1.8880870089577608 2.1897e-08 1.818584969510083 2.1898e-08 1.7081286857592577 2.1899e-08 1.795989147624853 2.19e-08 1.8533270400874227 2.1901e-08 1.861389819331149 2.1902e-08 1.7702858411061033 2.1903e-08 1.9008129692505957 2.1904e-08 1.8076005747538233 2.1905e-08 1.9351342685563937 2.1906e-08 1.7874039802601636 2.1907e-08 1.8369802490005391 2.1908e-08 1.711608352931967 2.1909e-08 1.6692052359407235 2.191e-08 1.819298754144613 2.1911e-08 1.7608652994718579 2.1911999999999998e-08 1.7649311734096969 2.1913e-08 1.799111648787381 2.1914e-08 1.8462244788004543 2.1914999999999998e-08 1.7305040647242538 2.1916e-08 1.8391338968576108 2.1917e-08 1.7867506529801622 2.1917999999999998e-08 1.804126689756671 2.1919e-08 1.7207372254793492 2.192e-08 1.8053228750978234 2.1920999999999998e-08 1.793412941252671 2.1922e-08 1.6923697367161739 2.1923e-08 1.7757310555372847 2.1923999999999998e-08 1.7065512478453517 2.1925e-08 1.846858814016251 2.1926e-08 1.8269842140245913 2.1927e-08 1.7776123706635314 2.1928e-08 1.7918210083916812 2.1929e-08 1.715059114839024 2.193e-08 1.8085155975087404 2.1931e-08 1.7309300042910973 2.1932e-08 1.7928546333978532 2.1933e-08 1.8172320484013433 2.1934e-08 1.8009340002144618 2.1935e-08 1.8300653553716972 2.1936e-08 1.8663808224583116 2.1937e-08 1.7853916480805758 2.1938e-08 1.8521159364171351 2.1939e-08 1.7175387593436733 2.194e-08 1.8054991657881865 2.1941e-08 1.8281692355806092 2.1942e-08 1.777216712580878 2.1943e-08 1.8386930422584464 2.1944e-08 1.7856516934991704 2.1945e-08 1.821393671207376 2.1946e-08 1.8412403374381276 2.1946999999999998e-08 1.8442451480336266 2.1948e-08 1.6796073339668078 2.1949e-08 1.9045125697231726 2.1949999999999998e-08 1.798138413374322 2.1951e-08 1.8746248187280525 2.1952e-08 1.8716440557381087 2.1952999999999998e-08 1.8412283314143165 2.1954e-08 1.7663345055072222 2.1955e-08 1.807386978713887 2.1955999999999998e-08 1.8448140427925785 2.1957e-08 1.8213293885564288 2.1958e-08 1.712387016064535 2.1958999999999998e-08 1.7899963244491175 2.196e-08 1.8606451065512473 2.1961e-08 1.8541735428184785 2.1962e-08 1.8155708083932691 2.1963e-08 1.793533103340572 2.1964e-08 1.8292121922780709 2.1965e-08 1.7807117306484088 2.1966e-08 1.8439566912863445 2.1967e-08 1.783462077873719 2.1968e-08 1.857160972012077 2.1969e-08 1.8895183689989685 2.197e-08 1.8498628989382602 2.1971e-08 1.8037346869204818 2.1972e-08 1.8164746723921847 2.1973e-08 1.9175892193176065 2.1974e-08 1.8375507912404592 2.1975e-08 1.7801150101468515 2.1976e-08 1.7517805213091873 2.1977e-08 1.720727492128547 2.1978e-08 1.8140766326264963 2.1979e-08 1.832872166231121 2.198e-08 1.7806110736600735 2.1981e-08 1.7237974147161979 2.1981999999999998e-08 1.755248514364577 2.1983e-08 1.782875725464062 2.1984e-08 1.7836820638489481 2.1984999999999998e-08 1.868309244344443 2.1986e-08 1.7143002709900454 2.1987e-08 1.8185842095407043 2.1987999999999998e-08 1.682209239020802 2.1989e-08 1.7893974940316 2.199e-08 1.7971805231407405 2.1990999999999998e-08 1.7958010682856997 2.1992e-08 1.788166906352001 2.1993e-08 1.817135144435986 2.1993999999999998e-08 1.8498488889586053 2.1995e-08 1.8660553013255274 2.1996e-08 1.7977366852947738 2.1997e-08 1.783866240642467 2.1998e-08 1.7676964657643734 2.1999e-08 1.865497531018285 2.2e-08 1.8116193415479622 2.2001e-08 1.7976168652327016 2.2002e-08 1.8151136043166738 2.2003e-08 1.8152026935550423 2.2004e-08 1.7684480416529282 2.2005e-08 1.8227462730866173 2.2006e-08 1.7354425312557955 2.2007e-08 1.780181749113997 2.2008e-08 1.8416224259805765 2.2009e-08 1.792401075292323 2.201e-08 1.7440350786046168 2.2011e-08 1.7806317889751215 2.2012e-08 1.7706011293993789 2.2013e-08 1.6669132885221194 2.2014e-08 1.8305311034268863 2.2015e-08 1.7723860526210005 2.2016e-08 1.7735854729183163 2.2017e-08 1.7721111939674432 2.2018e-08 1.7592857465669662 2.2019e-08 1.772877230217025 2.2019999999999998e-08 1.908651695063457 2.2021e-08 1.7741422355882406 2.2022e-08 1.7855284739479453 2.2022999999999998e-08 1.7879731346229766 2.2024e-08 1.8765341104798838 2.2025e-08 1.8301085043271088 2.2025999999999998e-08 1.8885302212708763 2.2027e-08 1.7768430129157067 2.2028e-08 1.848054834567299 2.2028999999999998e-08 1.747682618004413 2.203e-08 1.821360147499569 2.2031e-08 1.803236075881789 2.2032e-08 1.8409687113258328 2.2033e-08 1.7796638521101742 2.2034e-08 1.7860441895570176 2.2035e-08 1.7943309477123455 2.2036e-08 1.7776926619757847 2.2037e-08 1.8285365296685936 2.2038e-08 1.8161895675305753 2.2039e-08 1.8310720459133494 2.204e-08 1.670953742148683 2.2041e-08 1.766423299319201 2.2042e-08 1.7550936002530544 2.2043e-08 1.7883352463360882 2.2044e-08 1.80364989466879 2.2045e-08 1.911217253531358 2.2046e-08 1.7758418072557853 2.2047e-08 1.7654558192742174 2.2048e-08 1.7668007030188542 2.2049e-08 1.8318792777707318 2.205e-08 1.8268593692136526 2.2051e-08 1.77386388061761 2.2052e-08 1.8807714928350643 2.2053e-08 1.8085945149264637 2.2054e-08 1.775408092496064 2.2054999999999998e-08 1.7922222546529645 2.2056e-08 1.8559937066319132 2.2057e-08 1.7724122331609047 2.2057999999999998e-08 1.8387859576870862 2.2059e-08 1.8291785612277776 2.206e-08 1.852688800131666 2.2060999999999998e-08 1.8388972852985057 2.2062e-08 1.7310563522894937 2.2063e-08 1.7794510118137719 2.2063999999999998e-08 1.8280203804015707 2.2065e-08 1.9099912347465453 2.2066e-08 1.739227055932802 2.2067e-08 1.8202603935622168 2.2068e-08 1.8457895883547404 2.2069e-08 1.8391413850056144 2.207e-08 1.807057503632135 2.2071e-08 1.7642404420960858 2.2072e-08 1.80242351824752 2.2073e-08 1.833013054178852 2.2074e-08 1.7965719230233541 2.2075e-08 1.7687796376842913 2.2076e-08 1.826344262356568 2.2077e-08 1.8087743221818875 2.2078e-08 1.7488988585848664 2.2079e-08 1.8293739726882121 2.208e-08 1.7703671187068237 2.2081e-08 1.719296572563457 2.2082e-08 1.8130081427450098 2.2083e-08 1.775811581818124 2.2084e-08 1.765935663106481 2.2085e-08 1.7813951948191962 2.2086e-08 1.7493849497938356 2.2087e-08 1.7858989511191938 2.2088e-08 1.710490865671201 2.2089e-08 1.7275038759224144 2.2089999999999998e-08 1.7968186940118096 2.2091e-08 1.8692095252842025 2.2092e-08 1.8260158264156838 2.2092999999999998e-08 1.785671985947437 2.2094e-08 1.7981827328543496 2.2095e-08 1.8030178350655701 2.2095999999999998e-08 1.8600624159774588 2.2097e-08 1.837339731276357 2.2098e-08 1.882619841514012 2.2098999999999998e-08 1.874676966543273 2.21e-08 1.8167159645693112 2.2101e-08 1.8125776576790513 2.2101999999999998e-08 1.7775415403382042 2.2103e-08 1.8753634831000432 2.2104e-08 1.9069861797795904 2.2105e-08 1.7565579819593955 2.2106e-08 1.8025821531483655 2.2107e-08 1.8231760847115064 2.2108e-08 1.8010717503251925 2.2109e-08 1.7476290105436882 2.211e-08 1.7805581942656885 2.2111e-08 1.859141770441613 2.2112e-08 1.7365807190345697 2.2113e-08 1.841227070289525 2.2114e-08 1.738431166834328 2.2115e-08 1.8409382333980655 2.2116e-08 1.8237864112943494 2.2117e-08 1.8421673092536979 2.2118e-08 1.796789125421812 2.2119e-08 1.7623352351162802 2.212e-08 1.8549368052211899 2.2121e-08 1.776361678715027 2.2122e-08 1.843526769367098 2.2123e-08 1.7767251767491195 2.2124e-08 1.8352455080689642 2.2124999999999998e-08 1.7388957342377829 2.2126e-08 1.7863105477503727 2.2127e-08 1.8255832273686323 2.2127999999999998e-08 1.8773001300174783 2.2129e-08 1.784314459008916 2.213e-08 1.8070718961275771 2.2130999999999998e-08 1.775782297860514 2.2132e-08 1.840254896085828 2.2133e-08 1.8189964557132097 2.2133999999999998e-08 1.6584397251689464 2.2135e-08 1.7806259454705666 2.2136e-08 1.772481853609839 2.2136999999999998e-08 1.8198025463269698 2.2138e-08 1.7051411319221434 2.2139e-08 1.7084990882241846 2.214e-08 1.8498249615720728 2.2141e-08 1.8407750910966139 2.2142e-08 1.788280971136178 2.2143e-08 1.8357906114145746 2.2144e-08 1.8730610294283196 2.2145e-08 1.848406188516531 2.2146e-08 1.8299663089947857 2.2147e-08 1.8624109259007784 2.2148e-08 1.7906033470924134 2.2149e-08 1.8674303794706162 2.215e-08 1.7642541729554722 2.2151e-08 1.8302061098753568 2.2152e-08 1.8521179586906678 2.2153e-08 1.8140747881857813 2.2154e-08 1.7990810420486996 2.2155e-08 1.7359137202852952 2.2156e-08 1.7311716340702068 2.2157e-08 1.8060108530014345 2.2158e-08 1.785333832835066 2.2159e-08 1.7932418097506224 2.2159999999999998e-08 1.8245741970883302 2.2161e-08 1.760115473659833 2.2162e-08 1.7888085766740947 2.2162999999999998e-08 1.686488902089245 2.2164e-08 1.8637242128140612 2.2165e-08 1.8404521771104159 2.2165999999999998e-08 1.793932557345333 2.2167e-08 1.7520284870533915 2.2168e-08 1.7781342877064468 2.2168999999999998e-08 1.8122259907586402 2.217e-08 1.738242565971541 2.2171e-08 1.7793152477805134 2.2171999999999998e-08 1.7735485845344032 2.2173e-08 1.7897510269016057 2.2174e-08 1.7990729659307825 2.2175e-08 1.8106241517679615 2.2176e-08 1.820580553442918 2.2177e-08 1.743181906277724 2.2178e-08 1.8263776929826476 2.2179e-08 1.8162894665152314 2.218e-08 1.7970498310540424 2.2181e-08 1.7948622604212123 2.2182e-08 1.8922773591007755 2.2183e-08 1.7519191466180506 2.2184e-08 1.782934464172189 2.2185e-08 1.7623300526251109 2.2186e-08 1.8432168657768402 2.2187e-08 1.7785993311999206 2.2188e-08 1.8048552472466626 2.2189e-08 1.7442047621097314 2.219e-08 1.7985507946712465 2.2191e-08 1.8240100337131118 2.2192e-08 1.8265067446529588 2.2193e-08 1.7924112674794135 2.2194e-08 1.8261308965333158 2.2194999999999998e-08 1.7410198369645686 2.2196e-08 1.7977158156037476 2.2197e-08 1.8798591499379214 2.2197999999999998e-08 1.777164812179588 2.2199e-08 1.7810073142383909 2.22e-08 1.7295302320355943 2.2200999999999998e-08 1.8155463173425763 2.2202e-08 1.8185667471396774 2.2203e-08 1.8166873194983737 2.2203999999999998e-08 1.8186397286843197 2.2205e-08 1.8425586344745657 2.2206e-08 1.8637225544822578 2.2206999999999998e-08 1.7722764313791075 2.2208e-08 1.8078423020101837 2.2209e-08 1.777597361734558 2.221e-08 1.7244283920196914 2.2211e-08 1.8158759729070026 2.2212e-08 1.7516352916271172 2.2213e-08 1.7604362046282855 2.2214e-08 1.809623320771972 2.2215e-08 1.8510945516994037 2.2216e-08 1.7307389237027464 2.2217e-08 1.7927856722616728 2.2218e-08 1.7758380981438118 2.2219e-08 1.810496236939597 2.222e-08 1.8592071161371067 2.2221e-08 1.874817113868137 2.2222e-08 1.8474757448664574 2.2223e-08 1.8676099883428232 2.2224e-08 1.7401993859871503 2.2225e-08 1.8201478179763737 2.2226e-08 1.8126198967159945 2.2227e-08 1.8723914183309764 2.2228e-08 1.8419528366381317 2.2229e-08 1.7339636193161456 2.223e-08 1.8316315155244733 2.2231e-08 1.8433660345582836 2.2232e-08 1.8473307703641881 2.2232999999999998e-08 1.735978411526386 2.2234e-08 1.8226119997031658 2.2235e-08 1.8035038796330032 2.2235999999999998e-08 1.780241871008151 2.2237e-08 1.7988640051826066 2.2238e-08 1.795467992949745 2.2238999999999998e-08 1.8979861204113226 2.224e-08 1.7490965195152313 2.2241e-08 1.7679927118510734 2.2241999999999998e-08 1.879907123295179 2.2243e-08 1.7430269677847696 2.2244e-08 1.7483152302989609 2.2245e-08 1.7815262187325327 2.2246e-08 1.8296432361401784 2.2247e-08 1.8367071006949582 2.2248e-08 1.7628340043330413 2.2249e-08 1.8581389717412031 2.225e-08 1.777920958183815 2.2251e-08 1.8105341617814366 2.2252e-08 1.7852746375962565 2.2253e-08 1.7607894892841593 2.2254e-08 1.7463394436860167 2.2255e-08 1.7898031129017218 2.2256e-08 1.7751351752937943 2.2257e-08 1.8711521094463677 2.2258e-08 1.8693950507630925 2.2259e-08 1.8806789345373651 2.226e-08 1.8315021493337176 2.2261e-08 1.8307285953098387 2.2262e-08 1.8260072704509316 2.2263e-08 1.8348341450731736 2.2264e-08 1.7743801479141175 2.2265e-08 1.8187755769667764 2.2266e-08 1.8170763794673126 2.2267e-08 1.7180616222448397 2.2267999999999998e-08 1.7914964281285397 2.2269e-08 1.8811468713664081 2.227e-08 1.7153614670075001 2.2270999999999998e-08 1.8598481225240369 2.2272e-08 1.75274842325948 2.2273e-08 1.8525550464264926 2.2273999999999998e-08 1.7736953648469826 2.2275e-08 1.8555655554221897 2.2276e-08 1.8298767612929543 2.2276999999999998e-08 1.734811654925169 2.2278e-08 1.8313678350846487 2.2279e-08 1.807145819754391 2.2279999999999998e-08 1.7545348574797672 2.2281e-08 1.8078613788815858 2.2282e-08 1.818961681570925 2.2283e-08 1.8181964087900992 2.2284e-08 1.750740520506944 2.2285e-08 1.78353999626731 2.2286e-08 1.870282825617401 2.2287e-08 1.8112015612222825 2.2288e-08 1.7884337754888227 2.2289e-08 1.8620035394018886 2.229e-08 1.7773540156884537 2.2291e-08 1.8657964593784926 2.2292e-08 1.8561619010344794 2.2293e-08 1.7727768703108535 2.2294e-08 1.8266211703855122 2.2295e-08 1.7631959641314803 2.2296e-08 1.7399407531492228 2.2297e-08 1.8033258151119926 2.2298e-08 1.743414731668397 2.2299e-08 1.749773693707871 2.23e-08 1.830974695063408 2.2301e-08 1.910959481823385 2.2302e-08 1.7299876862762884 2.2302999999999998e-08 1.8152946069183875 2.2304e-08 1.7916488725205877 2.2305e-08 1.8133955677251787 2.2305999999999998e-08 1.7575739040654834 2.2307e-08 1.7561565342110794 2.2308e-08 1.739725100404261 2.2308999999999998e-08 1.852268384142627 2.231e-08 1.6461852362668115 2.2311e-08 1.7665741941950568 2.2311999999999998e-08 1.8581292381790124 2.2313e-08 1.8174275949637675 2.2314e-08 1.809209795728424 2.2314999999999998e-08 1.8024084845215287 2.2316e-08 1.9248975838987246 2.2317e-08 1.8095474734860133 2.2318e-08 1.8162668658965042 2.2319e-08 1.7384136789410138 2.232e-08 1.7169860670511332 2.2321e-08 1.851201249704014 2.2322e-08 1.8311528863084183 2.2323e-08 1.7698841249576376 2.2324e-08 1.8977193159897876 2.2325e-08 1.7741337804967336 2.2326e-08 1.8664218813322384 2.2327e-08 1.7874424431092106 2.2328e-08 1.8213084438930867 2.2329e-08 1.8480953450895974 2.233e-08 1.8502839786537804 2.2331e-08 1.7845655224227421 2.2332e-08 1.8517076979056613 2.2333e-08 1.6724722375023258 2.2334e-08 1.8302066306234615 2.2335e-08 1.8209696842689342 2.2336e-08 1.8555513671642851 2.2337e-08 1.7691980222907682 2.2337999999999998e-08 1.7597040659858336 2.2339e-08 1.7906897836646818 2.234e-08 1.7664818142211378 2.2340999999999998e-08 1.7850548520868872 2.2342e-08 1.8122599690781755 2.2343e-08 1.6531184846211981 2.2343999999999998e-08 1.7366435632544863 2.2345e-08 1.7730110521769897 2.2346e-08 1.8021216235258912 2.2346999999999998e-08 1.8595561277300507 2.2348e-08 1.7879555473501085 2.2349e-08 1.8636725800197582 2.2349999999999998e-08 1.8197581494674253 2.2351e-08 1.8182893047272373 2.2352e-08 1.8195484655666863 2.2353e-08 1.715727884228752 2.2354e-08 1.8374809933441476 2.2355e-08 1.7300675595353672 2.2356e-08 1.8159608032170482 2.2357e-08 1.6905194170005164 2.2358e-08 1.8126832845034522 2.2359e-08 1.7738906987023255 2.236e-08 1.8528612044559016 2.2361e-08 1.7623285131309547 2.2362e-08 1.7206571961160289 2.2363e-08 1.718709451569471 2.2364e-08 1.8295253551188315 2.2365e-08 1.7863856684798547 2.2366e-08 1.8391790254045413 2.2367e-08 1.7786914099749878 2.2368e-08 1.7897261010330472 2.2369e-08 1.7976866411079515 2.237e-08 1.8349841492103494 2.2371e-08 1.8267304615729925 2.2372e-08 1.8365918270332369 2.2372999999999998e-08 1.7739496749146435 2.2374e-08 1.8906865507873953 2.2375e-08 1.8246706511447952 2.2375999999999998e-08 1.838311747826951 2.2377e-08 1.7499434456525833 2.2378e-08 1.7571043661042924 2.2378999999999998e-08 1.7696682775107373 2.238e-08 1.7549030017626963 2.2381e-08 1.70592892868476 2.2381999999999998e-08 1.8082358327315373 2.2383e-08 1.799882810288515 2.2384e-08 1.8026800865858725 2.2384999999999998e-08 1.8056885456457308 2.2386e-08 1.8142577006667437 2.2387e-08 1.8656029148872921 2.2388e-08 1.75407251044974 2.2389e-08 1.882315221341068 2.239e-08 1.8562761393067886 2.2391e-08 1.8209427255971558 2.2392e-08 1.8141074970422923 2.2393e-08 1.7944867106424474 2.2394e-08 1.7673464235753855 2.2395e-08 1.7782785997336967 2.2396e-08 1.7664832275295652 2.2397e-08 1.8642035102907033 2.2398e-08 1.84200763991511 2.2399e-08 1.805813418806861 2.24e-08 1.7993912853606193 2.2401e-08 1.7726641906712004 2.2402e-08 1.8638208353716768 2.2403e-08 1.9135591340622389 2.2404e-08 1.7556197490431154 2.2405e-08 1.7488518706111182 2.2406e-08 1.8574752397172136 2.2407e-08 1.8323834535416723 2.2408e-08 1.746497189665014 2.2409e-08 1.7836359745420896 2.241e-08 1.839121239542149 2.2410999999999998e-08 1.8103658410798946 2.2412e-08 1.844718860848166 2.2413e-08 1.8718631008716962 2.2413999999999998e-08 1.7021333700291836 2.2415e-08 1.7614913328547765 2.2416e-08 1.8323801692446344 2.2416999999999998e-08 1.8117634207250717 2.2418e-08 1.804379603649983 2.2419e-08 1.854172658045829 2.2419999999999998e-08 1.8567578938216414 2.2421e-08 1.8260796552939165 2.2422e-08 1.7650147310007938 2.2423e-08 1.8225342769033186 2.2424e-08 1.722114737847555 2.2425e-08 1.8050076571872686 2.2426e-08 1.8431414993567692 2.2427e-08 1.8110157309513673 2.2428e-08 1.863837046549208 2.2429e-08 1.8027060458688955 2.243e-08 1.8827193409365488 2.2431e-08 1.749904468430453 2.2432e-08 1.7592349519401682 2.2433e-08 1.7649202353542899 2.2434e-08 1.85908600876827 2.2435e-08 1.880674441262077 2.2436e-08 1.8632990939216314 2.2437e-08 1.823106567119099 2.2438e-08 1.7569181332637342 2.2439e-08 1.724217030983458 2.244e-08 1.7659694942863597 2.2441e-08 1.765918512202243 2.2442e-08 1.7982643691613873 2.2443e-08 1.7884234779073342 2.2444e-08 1.7729936502039536 2.2445e-08 1.7264118613818755 2.2445999999999998e-08 1.8482725587161972 2.2447e-08 1.7893770029981844 2.2448e-08 1.728445776794389 2.2448999999999998e-08 1.7524873006664692 2.245e-08 1.7250265715605706 2.2451e-08 1.7189489713001749 2.2451999999999998e-08 1.7348530781185296 2.2453e-08 1.7798507841097009 2.2454e-08 1.909488448744828 2.2454999999999998e-08 1.769390981608826 2.2456e-08 1.7447525854785506 2.2457e-08 1.8225395230481525 2.2457999999999998e-08 1.792578675530729 2.2459e-08 1.7215828309431895 2.246e-08 1.791554749878728 2.2461e-08 1.7046673797083316 2.2462e-08 1.8574088640133546 2.2463e-08 1.752725468855083 2.2464e-08 1.8512866125915266 2.2465e-08 1.8471228803553048 2.2466e-08 1.797048665397197 2.2467e-08 1.7438908584926964 2.2468e-08 1.7934910512143787 2.2469e-08 1.7701843253334018 2.247e-08 1.7950947695301036 2.2471e-08 1.8365249240371537 2.2472e-08 1.7965849035315926 2.2473e-08 1.6848001614471082 2.2474e-08 1.821313421509647 2.2475e-08 1.803077264454471 2.2476e-08 1.7946457489208274 2.2477e-08 1.8157418916731847 2.2478e-08 1.8562424002028775 2.2479e-08 1.75916126639913 2.248e-08 1.7679818456351073 2.2480999999999998e-08 1.691858442015221 2.2482e-08 1.8115298350034277 2.2483e-08 1.795291524940967 2.2483999999999998e-08 1.821140068088962 2.2485e-08 1.8540592745331848 2.2486e-08 1.7886275074211615 2.2486999999999998e-08 1.7688736061552768 2.2488e-08 1.7553211481041837 2.2489e-08 1.8822945108398712 2.2489999999999998e-08 1.7705308694845892 2.2491e-08 1.6772738907727385 2.2492e-08 1.842385138067944 2.2492999999999998e-08 1.7831692553119587 2.2494e-08 1.8057588384446528 2.2495e-08 1.7815434218047848 2.2496e-08 1.792342579617134 2.2497e-08 1.7922004569384007 2.2498e-08 1.809078699708034 2.2499e-08 1.7585570160875494 2.25e-08 1.8873208902683705 2.2501e-08 1.7973558580229838 2.2502e-08 1.8820579140522666 2.2503e-08 1.735564954338257 2.2504e-08 1.7528347062382497 2.2505e-08 1.8435867367219234 2.2506e-08 1.7894220032732648 2.2507e-08 1.8043594894451147 2.2508e-08 1.8948695463154932 2.2509e-08 1.7511660267682485 2.251e-08 1.8338032948231164 2.2511e-08 1.879736438564569 2.2512e-08 1.85506844606208 2.2513e-08 1.8047903936128122 2.2514e-08 1.7720044250767604 2.2515e-08 1.7543146015162332 2.2515999999999998e-08 1.7999876405465278 2.2517e-08 1.796133482252793 2.2518e-08 1.844649429517833 2.2518999999999998e-08 1.766269419963047 2.252e-08 1.82753671236129 2.2521e-08 1.844078468457775 2.2521999999999998e-08 1.8435236436791091 2.2523e-08 1.8394880651240642 2.2524e-08 1.8107916382783422 2.2524999999999998e-08 1.793278278866273 2.2526e-08 1.8477331525104963 2.2527e-08 1.7731008723536077 2.2527999999999998e-08 1.8785943198308606 2.2529e-08 1.8064071949452276 2.253e-08 1.8401250991653073 2.2531e-08 1.7280400750034965 2.2532e-08 1.7149781842498313 2.2533e-08 1.8144140286678885 2.2534e-08 1.8148746724202245 2.2535e-08 1.7152189353079348 2.2536e-08 1.8447224986242021 2.2537e-08 1.7599476010646322 2.2538e-08 1.7975329695830482 2.2539e-08 1.7999665924487522 2.254e-08 1.8006678346722556 2.2541e-08 1.836181838548239 2.2542e-08 1.7496768701729 2.2543e-08 1.851832944014236 2.2544e-08 1.7925898257994912 2.2545e-08 1.805846992354244 2.2546e-08 1.835023610515893 2.2547e-08 1.7898219398219488 2.2548e-08 1.7984052536936204 2.2549e-08 1.8104204857406752 2.255e-08 1.8613871079749231 2.2550999999999998e-08 1.886118969526 2.2552e-08 1.8344305244165715 2.2553e-08 1.6747850579764543 2.2553999999999998e-08 1.7771717323294156 2.2555e-08 1.836791817089285 2.2556e-08 1.7457687892097211 2.2556999999999998e-08 1.8285319093873749 2.2558e-08 1.8163155253186354 2.2559e-08 1.8162644616132937 2.2559999999999998e-08 1.8201972036395673 2.2561e-08 1.9094182750510629 2.2562e-08 1.8438831138795442 2.2562999999999998e-08 1.7548330383284498 2.2564e-08 1.754849569336399 2.2565e-08 1.8409297351875502 2.2566e-08 1.8380788646432769 2.2567e-08 1.7841849014050235 2.2568e-08 1.794549076851266 2.2569e-08 1.7254598572609592 2.257e-08 1.7343071298163988 2.2571e-08 1.8014650937386727 2.2572e-08 1.7972512689047442 2.2573e-08 1.7914683423224094 2.2574e-08 1.7537852029529517 2.2575e-08 1.7784870741916237 2.2576e-08 1.8241137219375358 2.2577e-08 1.825813832526492 2.2578e-08 1.8490453525613328 2.2579e-08 1.8171458641254254 2.258e-08 1.7869128484571453 2.2581e-08 1.7507191220041098 2.2582e-08 1.8911419752410092 2.2583e-08 1.7892448764084552 2.2584e-08 1.8022433160683489 2.2585e-08 1.8496408037267007 2.2585999999999998e-08 1.8368452622675577 2.2587e-08 1.752928164198977 2.2588e-08 1.8092117462318702 2.2588999999999998e-08 1.8629573576128033 2.259e-08 1.7850567117985559 2.2591e-08 1.7876274844408928 2.2591999999999998e-08 1.8708545253133146 2.2593e-08 1.8740100120670011 2.2594e-08 1.8687727869057917 2.2594999999999998e-08 1.8843598528979362 2.2596e-08 1.8017993740154858 2.2597e-08 1.756108324053665 2.2597999999999998e-08 1.6599238777140737 2.2599e-08 1.8569145035825967 2.26e-08 1.7560518724840501 2.2601e-08 1.7107379731583716 2.2602e-08 1.7992370184568334 2.2603e-08 1.837268054254152 2.2604e-08 1.814938508238111 2.2605e-08 1.8477737886666028 2.2606e-08 1.877242547642698 2.2607e-08 1.8475298572920116 2.2608e-08 1.7908592850695424 2.2609e-08 1.8007109262906078 2.261e-08 1.8124934500443985 2.2611e-08 1.7920313653900968 2.2612e-08 1.8469267439092218 2.2613e-08 1.7825132922623743 2.2614e-08 1.7773524259843307 2.2615e-08 1.7879312318882263 2.2616e-08 1.783673321906509 2.2617e-08 1.7855912037260333 2.2618e-08 1.8134096712634653 2.2619e-08 1.8367420369811922 2.262e-08 1.851899768069974 2.2621e-08 1.8051787592717548 2.2622e-08 1.861239843516839 2.2623e-08 1.883729585442969 2.2623999999999998e-08 1.7890935015198373 2.2625e-08 1.8356684587937253 2.2626e-08 1.8566807031511678 2.2626999999999998e-08 1.8458750411083404 2.2628e-08 1.9144919038070953 2.2629e-08 1.789390121543424 2.2629999999999998e-08 1.7563994645756618 2.2631e-08 1.7986211496843219 2.2632e-08 1.8175071601404427 2.2632999999999998e-08 1.8064054074763736 2.2634e-08 1.7283329732250252 2.2635e-08 1.8312677957665766 2.2636e-08 1.7286612836186463 2.2637e-08 1.8157990732074396 2.2638e-08 1.7257974507747307 2.2639e-08 1.8527539124248877 2.264e-08 1.8281199430497215 2.2641e-08 1.7880369940632057 2.2642e-08 1.7667979714333215 2.2643e-08 1.7462895810113144 2.2644e-08 1.794997029041728 2.2645e-08 1.8472546453894363 2.2646e-08 1.7667191365659027 2.2647e-08 1.8163233399996606 2.2648e-08 1.8876649648103074 2.2649e-08 1.7915734034572888 2.265e-08 1.7909906927696455 2.2651e-08 1.7431712790848786 2.2652e-08 1.7750738895966751 2.2653e-08 1.8582540611613128 2.2654e-08 1.7968662406287128 2.2655e-08 1.7974540152098177 2.2656e-08 1.711473133627834 2.2657e-08 1.8115717267479794 2.2658e-08 1.699587690953262 2.2658999999999998e-08 1.6399446847033832 2.266e-08 1.8077759648040077 2.2661e-08 1.858173798821083 2.2661999999999998e-08 1.8342289058174135 2.2663e-08 1.7801004837216008 2.2664e-08 1.7664614902777152 2.2664999999999998e-08 1.8155618838131538 2.2666e-08 1.781868316711287 2.2667e-08 1.7745271809371501 2.2667999999999998e-08 1.7091375147532508 2.2669e-08 1.7666010735661788 2.267e-08 1.8077723915333914 2.2670999999999998e-08 1.7392483634162241 2.2672e-08 1.8387715770031694 2.2673e-08 1.756193862614544 2.2674e-08 1.887520576817139 2.2675e-08 1.8235682192251326 2.2676e-08 1.8577266729561275 2.2677e-08 1.7664766887656247 2.2678e-08 1.7473007722335099 2.2679e-08 1.7214074935489072 2.268e-08 1.842559811773124 2.2681e-08 1.7456989964530325 2.2682e-08 1.8251226952662187 2.2683e-08 1.8340194333580087 2.2684e-08 1.8563492469196579 2.2685e-08 1.788731204883575 2.2686e-08 1.7907403260394479 2.2687e-08 1.832501961842042 2.2688e-08 1.829591202128995 2.2689e-08 1.8016494109325383 2.269e-08 1.7398702342922823 2.2691e-08 1.8049250076429588 2.2692e-08 1.797595715452463 2.2693e-08 1.7915856384242066 2.2693999999999998e-08 1.8208540798642772 2.2695e-08 1.7418225450877236 2.2696e-08 1.8338070503894697 2.2696999999999998e-08 1.7690796989303788 2.2698e-08 1.8399889647272365 2.2699e-08 1.8006084150589665 2.2699999999999998e-08 1.7615999936698232 2.2701e-08 1.7759727743301743 2.2702e-08 1.8363652847779304 2.2702999999999998e-08 1.8541048921214252 2.2704e-08 1.776571495468238 2.2705e-08 1.7316714988894717 2.2705999999999998e-08 1.6954113794775738 2.2707e-08 1.7702904414966159 2.2708e-08 1.829050058949119 2.2709e-08 1.8087118252818313 2.271e-08 1.9472506550173645 2.2711e-08 1.7648927750802756 2.2712e-08 1.7369352441999792 2.2713e-08 1.7297447749133243 2.2714e-08 1.8757938824431888 2.2715e-08 1.8217585208089364 2.2716e-08 1.6882434875400407 2.2717e-08 1.7546577513410408 2.2718e-08 1.80041013123945 2.2719e-08 1.8708014224086924 2.272e-08 1.8331926881970608 2.2721e-08 1.8287009507925542 2.2722e-08 1.8372521398818111 2.2723e-08 1.856428205042776 2.2724e-08 1.734499316911723 2.2725e-08 1.7978438228585107 2.2726e-08 1.7161851290599446 2.2727e-08 1.8846114594809942 2.2728e-08 1.8237296813973976 2.2728999999999998e-08 1.8009087786921405 2.273e-08 1.7576535789340955 2.2731e-08 1.7339759789909108 2.2731999999999998e-08 1.768505232863511 2.2733e-08 1.8619761647952062 2.2734e-08 1.8749054148730078 2.2734999999999998e-08 1.8094119395533923 2.2736e-08 1.8144365482665585 2.2737e-08 1.7877874263960736 2.2737999999999998e-08 1.8434461445337258 2.2739e-08 1.7867933640947224 2.274e-08 1.7849177384508246 2.2740999999999998e-08 1.8449711643187086 2.2742e-08 1.7794936102413181 2.2743e-08 1.773226338059042 2.2744e-08 1.8714430089187606 2.2745e-08 1.8269558516944604 2.2746e-08 1.80380089873111 2.2747e-08 1.8188029591461843 2.2748e-08 1.778821770676319 2.2749e-08 1.8154079233419373 2.275e-08 1.8026511424326432 2.2751e-08 1.7517470136941848 2.2752e-08 1.8907912943194611 2.2753e-08 1.8118693140264437 2.2754e-08 1.7540809830480377 2.2755e-08 1.7007171997374282 2.2756e-08 1.7630378449578312 2.2757e-08 1.8422409212217399 2.2758e-08 1.790240779217299 2.2759e-08 1.8426064869975072 2.276e-08 1.7969686731450654 2.2761e-08 1.8242098412859482 2.2762e-08 1.7730724771838706 2.2763e-08 1.6708123685853444 2.2763999999999998e-08 1.8404091776737188 2.2765e-08 1.8679596941493468 2.2766e-08 1.8433919913289072 2.2766999999999998e-08 1.8438994812420746 2.2768e-08 1.743162126700481 2.2769e-08 1.8116990380225575 2.2769999999999998e-08 1.8284572720776173 2.2771e-08 1.9273316634662203 2.2772e-08 1.7193513406910186 2.2772999999999998e-08 1.7847508090213382 2.2774e-08 1.8149208551533043 2.2775e-08 1.7251674977575324 2.2775999999999998e-08 1.8002412360764457 2.2777e-08 1.7711987497240975 2.2778e-08 1.7975953736046153 2.2779e-08 1.804897718910294 2.278e-08 1.8879098235088947 2.2781e-08 1.778836110943133 2.2782e-08 1.722096245863083 2.2783e-08 1.916730427212426 2.2784e-08 1.7597905140535117 2.2785e-08 1.8327279103491976 2.2786e-08 1.863380836856409 2.2787e-08 1.8418838507703648 2.2788e-08 1.7650763153748135 2.2789e-08 1.7509409328508332 2.279e-08 1.8482008875011995 2.2791e-08 1.8236712382494533 2.2792e-08 1.7983407364708488 2.2793e-08 1.9522270395288879 2.2794e-08 1.7904328607979605 2.2795e-08 1.882188767775658 2.2796e-08 1.7831106299613524 2.2797e-08 1.857632699913209 2.2798e-08 1.8084058724990215 2.2798999999999998e-08 1.8506453938192944 2.28e-08 1.8352195909255593 2.2801e-08 1.8493665935737813 2.2801999999999998e-08 1.846579344636146 2.2803e-08 1.8126596319956843 2.2804e-08 1.8294173447575435 2.2804999999999998e-08 1.8129231428727524 2.2806e-08 1.8424331962725295 2.2807e-08 1.8182813199201249 2.2807999999999998e-08 1.7944310093262574 2.2809e-08 1.780071186179552 2.281e-08 1.791858624534619 2.2810999999999998e-08 1.8216179809358855 2.2812e-08 1.8069743306413404 2.2813e-08 1.806549566299711 2.2814e-08 1.7983958372661863 2.2815e-08 1.7909587771518511 2.2816e-08 1.720877016216252 2.2817e-08 1.8115791023744596 2.2818e-08 1.679724924501289 2.2819e-08 1.80888750355931 2.282e-08 1.6939106425346082 2.2821e-08 1.8689475275255971 2.2822e-08 1.8786999371600275 2.2823e-08 1.8210141247021094 2.2824e-08 1.873014905548321 2.2825e-08 1.817387301447899 2.2826e-08 1.7732565435721068 2.2827e-08 1.8451180555335664 2.2828e-08 1.8370665120086151 2.2829e-08 1.7924382709225442 2.283e-08 1.861632324435953 2.2831e-08 1.8923335883211247 2.2832e-08 1.7453049655628652 2.2833e-08 1.7604733310958591 2.2834e-08 1.7844962703960228 2.2835e-08 1.8538713865314551 2.2836e-08 1.810068664177388 2.2836999999999998e-08 1.73917266645911 2.2838e-08 1.8310143574713804 2.2839e-08 1.7502085652058421 2.2839999999999998e-08 1.8327635844176071 2.2841e-08 1.8223391677389578 2.2842e-08 1.8165642657725398 2.2842999999999998e-08 1.8326811424675522 2.2844e-08 1.811006049424306 2.2845e-08 1.8095259886622812 2.2845999999999998e-08 1.8099452016919224 2.2847e-08 1.7620525898899917 2.2848e-08 1.840482082095854 2.2848999999999998e-08 1.8176213363006921 2.285e-08 1.7671407838267115 2.2851e-08 1.8188844660110766 2.2852e-08 1.7817853619664246 2.2853e-08 1.8552835590577383 2.2854e-08 1.6033770675794154 2.2855e-08 1.816069468708934 2.2856e-08 1.8390590976380246 2.2857e-08 1.7845657687151155 2.2858e-08 1.7646389296846652 2.2859e-08 1.8699528386238173 2.286e-08 1.883349627375958 2.2861e-08 1.8027304732318212 2.2862e-08 1.7646595802964153 2.2863e-08 1.8643302737256622 2.2864e-08 1.8748143769352212 2.2865e-08 1.808407138983465 2.2866e-08 1.839709280934388 2.2867e-08 1.7911631499770848 2.2868e-08 1.8121127581147518 2.2869e-08 1.9133837972251433 2.287e-08 1.848064233664532 2.2871e-08 1.8598589843391848 2.2871999999999998e-08 1.8483748747366164 2.2873e-08 1.8126775697070032 2.2874e-08 1.8460614433211562 2.2874999999999998e-08 1.7999858872370726 2.2876e-08 1.8410452538667537 2.2877e-08 1.8942801744300828 2.2877999999999998e-08 1.796122578361526 2.2879e-08 1.7885675815676239 2.288e-08 1.7548674210307253 2.2880999999999998e-08 1.726430253473319 2.2882e-08 1.746386308966869 2.2883e-08 1.8096945699200735 2.2883999999999998e-08 1.7839993410063875 2.2885e-08 1.6741221057787032 2.2886e-08 1.9194364473520773 2.2887e-08 1.8765115006934416 2.2888e-08 1.840627555548339 2.2889e-08 1.7250518871020406 2.289e-08 1.8122014692467796 2.2891e-08 1.803201598814765 2.2892e-08 1.8293056939834087 2.2893e-08 1.7791027147415026 2.2894e-08 1.7502096094451636 2.2895e-08 1.733634780869401 2.2896e-08 1.85528330181646 2.2897e-08 1.8142986666296257 2.2898e-08 1.8719023901495582 2.2899e-08 1.8316600810067056 2.29e-08 1.7593073848824154 2.2901e-08 1.725023813969383 2.2902e-08 1.7619282239002039 2.2903e-08 1.79475980091966 2.2904e-08 1.8277252388306793 2.2905e-08 1.78856707952014 2.2906e-08 1.8015709166541327 2.2906999999999998e-08 1.7598101675395974 2.2908e-08 1.7310087945690713 2.2909e-08 1.87715372794955 2.2909999999999998e-08 1.6801681789681595 2.2911e-08 1.7863182101577817 2.2912e-08 1.7344680663482999 2.2912999999999998e-08 1.8331880242570766 2.2914e-08 1.7667841829362712 2.2915e-08 1.8109428786772346 2.2915999999999998e-08 1.8389277231165204 2.2917e-08 1.7556200644533038 2.2918e-08 1.744804144374089 2.2918999999999998e-08 1.7208314044863469 2.292e-08 1.856608226252024 2.2921e-08 1.8408292756841282 2.2922e-08 1.8573995078050083 2.2923e-08 1.7679048934241222 2.2924e-08 1.814562028384473 2.2925e-08 1.7858003359971701 2.2926e-08 1.8077262087774848 2.2927e-08 1.8378775509377758 2.2928e-08 1.7907980183870378 2.2929e-08 1.6978983036825668 2.293e-08 1.8097967727989928 2.2931e-08 1.7625202409397827 2.2932e-08 1.8103339490840946 2.2933e-08 1.8110415886135116 2.2934e-08 1.8414219091302644 2.2935e-08 1.754739317454237 2.2936e-08 1.7740895384404962 2.2937e-08 1.753929741002505 2.2938e-08 1.8369559329841165 2.2939e-08 1.7520214548922184 2.294e-08 1.8100044222294882 2.2941e-08 1.7001737520982012 2.2941999999999998e-08 1.8132667224982655 2.2943e-08 1.8147782335418428 2.2944e-08 1.7679991375253596 2.2944999999999998e-08 1.7442102235667907 2.2946e-08 1.9428220901827484 2.2947e-08 1.8633188881078724 2.2947999999999998e-08 1.72716474361833 2.2949e-08 1.8141029558250286 2.295e-08 1.724687936277313 2.2950999999999998e-08 1.7999399953739272 2.2952e-08 1.8037062698134076 2.2953e-08 1.7918037914075937 2.2953999999999998e-08 1.8052636582741026 2.2955e-08 1.8293876710780659 2.2956e-08 1.9048472446167894 2.2957e-08 1.8789579312903575 2.2958e-08 1.755795801349577 2.2959e-08 1.8264283592930635 2.296e-08 1.7802735438031003 2.2961e-08 1.7513207990214088 2.2962e-08 1.8510694236680072 2.2963e-08 1.727675340276933 2.2964e-08 1.8383542698303974 2.2965e-08 1.7682414632377272 2.2966e-08 1.8408429307746867 2.2967e-08 1.7598876768214378 2.2968e-08 1.821762936010753 2.2969e-08 1.780123676411412 2.297e-08 1.890135261121962 2.2971e-08 1.8203534586266676 2.2972e-08 1.8253839623581325 2.2973e-08 1.7754990970054112 2.2974e-08 1.7898378519085674 2.2975e-08 1.6915384791702759 2.2976e-08 1.7076396861878966 2.2976999999999998e-08 1.82482553400164 2.2978e-08 1.7508513039259395 2.2979e-08 1.7991474594634584 2.2979999999999998e-08 1.7706936879703838 2.2981e-08 1.8419096993857833 2.2982e-08 1.7963488801143477 2.2982999999999998e-08 1.7106884210407827 2.2984e-08 1.80850671658098 2.2985e-08 1.7546494203232057 2.2985999999999998e-08 1.8014379481229448 2.2987e-08 1.8451347500856001 2.2988e-08 1.8198333887162335 2.2988999999999998e-08 1.7926655859981913 2.299e-08 1.8398997812492301 2.2991e-08 1.8460181407466445 2.2992e-08 1.8225153665054012 2.2993e-08 1.7541223687622478 2.2994e-08 1.7888506436708909 2.2995e-08 1.7771648423665753 2.2996e-08 1.7670966554125376 2.2997e-08 1.7747684701100488 2.2998e-08 1.7743126012371826 2.2999e-08 1.810958275367358 2.3e-08 1.80106238098907 2.3001e-08 1.780524197354298 2.3002e-08 1.7715589118431962 2.3003e-08 1.7822490597711476 2.3004e-08 1.759027982789887 2.3005e-08 1.7589381279065954 2.3006e-08 1.7562007850330008 2.3007e-08 1.7693602055453823 2.3008e-08 1.82493371616962 2.3009e-08 1.7750190743795387 2.301e-08 1.8035045970139179 2.3011e-08 1.7974995916488525 2.3012e-08 1.7699696910385954 2.3013e-08 1.7670676288533453 2.3014e-08 1.8111585653146132 2.3014999999999998e-08 1.798733778122968 2.3016e-08 1.8052843734821726 2.3017e-08 1.856148163337049 2.3017999999999998e-08 1.809385562714048 2.3019e-08 1.8184903089307014 2.302e-08 1.8099397644519508 2.3020999999999998e-08 1.8023003901585481 2.3022e-08 1.818194274746624 2.3023e-08 1.8825730661838682 2.3023999999999998e-08 1.809806271779197 2.3025e-08 1.7820755080419768 2.3026e-08 1.7408066355288072 2.3026999999999998e-08 1.7699141895277806 2.3028e-08 1.760172961648319 2.3029e-08 1.7303836836744122 2.303e-08 1.728208509780884 2.3031e-08 1.758228495291299 2.3032e-08 1.7907740202389775 2.3033e-08 1.7773969966174792 2.3034e-08 1.8089620719026982 2.3035e-08 1.809149872780478 2.3036e-08 1.8593029466609936 2.3037e-08 1.7753292957017708 2.3038e-08 1.7964552630200663 2.3039e-08 1.8367130764538584 2.304e-08 1.8487956301811015 2.3041e-08 1.785878211710868 2.3042e-08 1.7511006668958229 2.3043e-08 1.7792514535043158 2.3044e-08 1.8235557305934347 2.3045e-08 1.8775928623917202 2.3046e-08 1.7781993990332354 2.3047e-08 1.8251891541489145 2.3048e-08 1.7832322961826252 2.3049e-08 1.757227718632908 2.3049999999999998e-08 1.7739068445734991 2.3051e-08 1.7969446395198267 2.3052e-08 1.7941567845802124 2.3052999999999998e-08 1.7717630649987781 2.3054e-08 1.7601333145619502 2.3055e-08 1.7995761567883921 2.3055999999999998e-08 1.8154826214794593 2.3057e-08 1.8352409973880635 2.3058e-08 1.7577949338121392 2.3058999999999998e-08 1.7885557472061744 2.306e-08 1.7505146273619654 2.3061e-08 1.8710845337218145 2.3061999999999998e-08 1.8325404071142584 2.3063e-08 1.7721652431372026 2.3064e-08 1.8198115235954526 2.3065e-08 1.6913096631007505 2.3066e-08 1.8516965024502667 2.3067e-08 1.802317730815636 2.3068e-08 1.8549774427353705 2.3069e-08 1.7712562616337135 2.307e-08 1.8467563349640408 2.3071e-08 1.739183708636016 2.3072e-08 1.7739369154236455 2.3073e-08 1.7983590226447264 2.3074e-08 1.8280695508223086 2.3075e-08 1.8419903325831428 2.3076e-08 1.7634956433880893 2.3077e-08 1.7882305372677563 2.3078e-08 1.887456320738735 2.3079e-08 1.7813840911924195 2.308e-08 1.8018371568821596 2.3081e-08 1.83606937388821 2.3082e-08 1.7386060390500002 2.3083e-08 1.7317148385953631 2.3084e-08 1.7913828624458963 2.3084999999999998e-08 1.86314806448528 2.3086e-08 1.8356714401618226 2.3087e-08 1.886868559802502 2.3087999999999998e-08 1.739820075750389 2.3089e-08 1.754738078639268 2.309e-08 1.7647381031576426 2.3090999999999998e-08 1.7483520359075455 2.3092e-08 1.8107126239698441 2.3093e-08 1.8549168613262905 2.3093999999999998e-08 1.7424247106581643 2.3095e-08 1.8363150437489044 2.3096e-08 1.7441077473844047 2.3096999999999998e-08 1.799637227938459 2.3098e-08 1.7243058348352824 2.3099e-08 1.8047501281557892 2.31e-08 1.8155080139514492 2.3101e-08 1.89273209759012 2.3102e-08 1.7596509173018977 2.3103e-08 1.8718108718912843 2.3104e-08 1.7469537798843804 2.3105e-08 1.8717392551056644 2.3106e-08 1.8388694820984397 2.3107e-08 1.7293406524729307 2.3108e-08 1.781324911984002 2.3109e-08 1.8087931438114808 2.311e-08 1.7660966298320888 2.3111e-08 1.729459880637957 2.3112e-08 1.802031597266224 2.3113e-08 1.8252915767956546 2.3114e-08 1.7953642524603817 2.3115e-08 1.7100701144067618 2.3116e-08 1.7852251563899928 2.3117e-08 1.8006425169146487 2.3118e-08 1.747988845506174 2.3119e-08 1.782351716246859 2.3119999999999998e-08 1.7976590212073968 2.3121e-08 1.80846665293696 2.3122e-08 1.85021300804935 2.3122999999999998e-08 1.787534560469214 2.3124e-08 1.8073979055318428 2.3125e-08 1.7729797557074856 2.3125999999999998e-08 1.8577369177957188 2.3127e-08 1.8416812870609347 2.3128e-08 1.7504721589200045 2.3128999999999998e-08 1.8449529285021793 2.313e-08 1.816258132439062 2.3131e-08 1.7913835432442846 2.3131999999999998e-08 1.8444457727338943 2.3133e-08 1.711652723560265 2.3134e-08 1.8153874288089606 2.3135e-08 1.8473752182315695 2.3136e-08 1.8385422581436155 2.3137e-08 1.697191510693814 2.3138e-08 1.8113507131442415 2.3139e-08 1.7707506497510468 2.314e-08 1.7997793095927466 2.3141e-08 1.8391638547663043 2.3142e-08 1.7590780946777285 2.3143e-08 1.880917904275165 2.3144e-08 1.801560916230265 2.3145e-08 1.867228488337929 2.3146e-08 1.8104184408148494 2.3147e-08 1.8231266906170849 2.3148e-08 1.8022135895899662 2.3149e-08 1.7828902428931368 2.315e-08 1.8840798393598877 2.3151e-08 1.7523174709940732 2.3152e-08 1.8270986940905773 2.3153e-08 1.7159955758066952 2.3154e-08 1.7743978042365882 2.3154999999999998e-08 1.7555658164418009 2.3156e-08 1.8631743205412197 2.3157e-08 1.7322074842902866 2.3157999999999998e-08 1.8108833449405886 2.3159e-08 1.8612175397089692 2.316e-08 1.8040469953466707 2.3160999999999998e-08 1.8280794960289715 2.3162e-08 1.763974678181241 2.3163e-08 1.7486652554044018 2.3163999999999998e-08 1.7512971562056294 2.3165e-08 1.7946367041278657 2.3166e-08 1.8047464095256414 2.3166999999999998e-08 1.907671225551652 2.3168e-08 1.9035049819230079 2.3169e-08 1.8082110165572811 2.317e-08 1.7172176938056238 2.3171e-08 1.7646202802845627 2.3172e-08 1.656209703825459 2.3173e-08 1.8284080261595175 2.3174e-08 1.7629855897108984 2.3175e-08 1.8044487921860706 2.3176e-08 1.856820748212325 2.3177e-08 1.782118219158093 2.3178e-08 1.7538879120880846 2.3179e-08 1.7608608993605017 2.318e-08 1.7746259839581258 2.3181e-08 1.7098358808961125 2.3182e-08 1.7779909158035097 2.3183e-08 1.8356491935662038 2.3184e-08 1.7322230043736664 2.3185e-08 1.833895666102909 2.3186e-08 1.7626437506185337 2.3187e-08 1.7616938472234722 2.3188e-08 1.7826495451226552 2.3189e-08 1.817402862440683 2.3189999999999998e-08 1.898040746397223 2.3191e-08 1.851260619290829 2.3192e-08 1.8365913560525935 2.3192999999999998e-08 1.7120413951852624 2.3194e-08 1.8988180241022712 2.3195e-08 1.8636215381597854 2.3195999999999998e-08 1.7876281207504847 2.3197e-08 1.782684029438177 2.3198e-08 1.8240682553864958 2.3198999999999998e-08 1.8837081294606395 2.32e-08 1.7652184724166868 2.3201e-08 1.8307229930432747 2.3201999999999998e-08 1.8277583785387808 2.3203e-08 1.7472514486371407 2.3204e-08 1.7708367567561256 2.3205e-08 1.7393252461566717 2.3206e-08 1.750907714079702 2.3207e-08 1.7033251637462106 2.3208e-08 1.8202902719381298 2.3209e-08 1.7768085649362433 2.321e-08 1.7989697115119978 2.3211e-08 1.7559609108129952 2.3212e-08 1.7525560169481285 2.3213e-08 1.7780891798019423 2.3214e-08 1.8772450715923112 2.3215e-08 1.8017366215228197 2.3216e-08 1.8299536462455253 2.3217e-08 1.754749177595354 2.3218e-08 1.806811657384045 2.3219e-08 1.783035919383132 2.322e-08 1.7360218217054335 2.3221e-08 1.7249184141356162 2.3222e-08 1.8491234790627271 2.3223e-08 1.7893017874370285 2.3224e-08 1.8316023126499543 2.3225e-08 1.7565016861518146 2.3226e-08 1.7937928304938418 2.3227e-08 1.816837083670596 2.3227999999999998e-08 1.8014754884626303 2.3229e-08 1.8441493097819608 2.323e-08 1.7600586431982213 2.3230999999999998e-08 1.9064096578499925 2.3232e-08 1.7950509269727954 2.3233e-08 1.70853927384706 2.3233999999999998e-08 1.7488386671682026 2.3235e-08 1.8373523176141116 2.3236e-08 1.7867871983277948 2.3236999999999998e-08 1.8188089266895273 2.3238e-08 1.7965946994740893 2.3239e-08 1.8099665080415002 2.3239999999999998e-08 1.7355838191753383 2.3241e-08 1.8031388819781295 2.3242e-08 1.8496029794165263 2.3243e-08 1.8227725546380347 2.3244e-08 1.8325038365182924 2.3245e-08 1.8205036113808002 2.3246e-08 1.7468361880152643 2.3247e-08 1.802362270617638 2.3248e-08 1.8478475655732127 2.3249e-08 1.8818683340836904 2.325e-08 1.788135195678782 2.3251e-08 1.8012212043346298 2.3252e-08 1.91344058522318 2.3253e-08 1.7938491336938591 2.3254e-08 1.9371467328169376 2.3255e-08 1.7902580206471999 2.3256e-08 1.7407174321514796 2.3257e-08 1.7940736537733109 2.3258e-08 1.7528258887037997 2.3259e-08 1.7792647391601268 2.326e-08 1.7219278207371194 2.3261e-08 1.9078288559968568 2.3262e-08 1.7188366978661302 2.3262999999999998e-08 1.757341148705894 2.3264e-08 1.8160205179086382 2.3265e-08 1.844105856637081 2.3265999999999998e-08 1.79548661379971 2.3267e-08 1.772069370112023 2.3268e-08 1.7959161113867963 2.3268999999999998e-08 1.7882417456156543 2.327e-08 1.7953697366282988 2.3271e-08 1.7543963979308548 2.3271999999999998e-08 1.8215822636015442 2.3273e-08 1.7996319808115246 2.3274e-08 1.7288973303808413 2.3274999999999998e-08 1.7635518132649795 2.3276e-08 1.7714951635410099 2.3277e-08 1.7669226462954746 2.3278e-08 1.8816240634632604 2.3279e-08 1.8075273567281798 2.328e-08 1.8369109513018664 2.3281e-08 1.7934235401221041 2.3282e-08 1.8983818099691763 2.3283e-08 1.8573980929481673 2.3284e-08 1.805788257890386 2.3285e-08 1.8611871097339516 2.3286e-08 1.8579728783837295 2.3287e-08 1.7072444640097806 2.3288e-08 1.7995561174394497 2.3289e-08 1.847596618380974 2.329e-08 1.8373002471724968 2.3291e-08 1.7271062837832019 2.3292e-08 1.8383285866834005 2.3293e-08 1.8525323423006674 2.3294e-08 1.7695000731942088 2.3295e-08 1.8082957696602222 2.3296e-08 1.7802407091092334 2.3297e-08 1.8073721649790246 2.3297999999999998e-08 1.791718220677541 2.3299e-08 1.8729225629870945 2.33e-08 1.7869043950353405 2.3300999999999998e-08 1.8340032411283982 2.3302e-08 1.859089766921593 2.3303e-08 1.8864268929890942 2.3303999999999998e-08 1.7994192861866583 2.3305e-08 1.7722612576868466 2.3306e-08 1.8054868895553973 2.3306999999999998e-08 1.843849771005071 2.3308e-08 1.8961839649124392 2.3309e-08 1.8033305586740875 2.3309999999999998e-08 1.7693745832370855 2.3311e-08 1.7823498236266755 2.3312e-08 1.8107486325632725 2.3313e-08 1.8281203079781463 2.3314e-08 1.8304595100458616 2.3315e-08 1.8487692789567978 2.3316e-08 1.7997053923202664 2.3317e-08 1.7730821716737815 2.3318e-08 1.7342251581749786 2.3319e-08 1.8167651180704254 2.332e-08 1.8401066760879696 2.3321e-08 1.7866336898172983 2.3322e-08 1.7776066053255404 2.3323e-08 1.822317795128546 2.3324e-08 1.7603530892597126 2.3325e-08 1.782491085880079 2.3326e-08 1.7851028490959209 2.3327e-08 1.6897211100760279 2.3328e-08 1.8404784456754 2.3329e-08 1.8544800447478038 2.333e-08 1.7550549926997818 2.3331e-08 1.9121230686045243 2.3332e-08 1.8054780074590444 2.3332999999999998e-08 1.838412807636596 2.3334e-08 1.7920679682840388 2.3335e-08 1.7679849861339054 2.3335999999999998e-08 1.744550725104911 2.3337e-08 1.7254647218117403 2.3338e-08 1.7651270678214472 2.3338999999999998e-08 1.7347815211095328 2.334e-08 1.8227522729707588 2.3341e-08 1.8901921633923207 2.3341999999999998e-08 1.9120197973990392 2.3343e-08 1.8259258242049312 2.3344e-08 1.8063351573691513 2.3344999999999998e-08 1.8083969133384763 2.3346e-08 1.7736882992754408 2.3347e-08 1.7029663334241232 2.3348e-08 1.905323515051351 2.3349e-08 1.8371217117739003 2.335e-08 1.8280706321826639 2.3351e-08 1.7508201445129457 2.3352e-08 1.790237763498958 2.3353e-08 1.8036525485410404 2.3354e-08 1.8025957108869024 2.3355e-08 1.73709368027076 2.3356e-08 1.8888579917530228 2.3357e-08 1.7778077450285161 2.3358e-08 1.8230942807006114 2.3359e-08 1.8409323431194724 2.336e-08 1.8557180763230694 2.3361e-08 1.817385885706418 2.3362e-08 1.8274033410858876 2.3363e-08 1.8855600177875529 2.3364e-08 1.8400559059789392 2.3365e-08 1.8399179774596919 2.3366e-08 1.7786079323456794 2.3367e-08 1.7658426992747625 2.3367999999999998e-08 1.9302835592944905 2.3369e-08 1.8381955439671651 2.337e-08 1.8288055872509437 2.3370999999999998e-08 1.7401782233089842 2.3372e-08 1.795098236484609 2.3373e-08 1.7864600001151936 2.3373999999999998e-08 1.7660426717483106 2.3375e-08 1.788070264527237 2.3376e-08 1.7896088378538084 2.3376999999999998e-08 1.843523645199691 2.3378e-08 1.7885774768186011 2.3379e-08 1.7530310726908536 2.3379999999999998e-08 1.761086487132109 2.3381e-08 1.882210886428454 2.3382e-08 1.8591164792206987 2.3383e-08 1.84065545488807 2.3384e-08 1.796739613331793 2.3385e-08 1.828454906666943 2.3386e-08 1.8760871646742694 2.3387e-08 1.9334830107336598 2.3388e-08 1.7656072082484786 2.3389e-08 1.7657700288085252 2.339e-08 1.7247994398161541 2.3391e-08 1.8834749539569933 2.3392e-08 1.8260863973636037 2.3393e-08 1.7781739589448773 2.3394e-08 1.8288158934252379 2.3395e-08 1.8009274558290629 2.3396e-08 1.7689983330006624 2.3397e-08 1.8040475565259966 2.3398e-08 1.8418268102598783 2.3399e-08 1.8745320113545971 2.34e-08 1.7610449695314387 2.3401e-08 1.832672390512958 2.3402e-08 1.806697955346639 2.3403e-08 1.8133447001082514 2.3404e-08 1.8876754580197925 2.3405e-08 1.7847499553399686 2.3405999999999998e-08 1.7330525032993906 2.3407e-08 1.7800914744083696 2.3408e-08 1.7973197974944966 2.3408999999999998e-08 1.8679942198913044 2.341e-08 1.7636452001610214 2.3411e-08 1.7984282185574334 2.3411999999999998e-08 1.8196369759940274 2.3413e-08 1.827764857086349 2.3414e-08 1.77103888234963 2.3414999999999998e-08 1.8724607283436026 2.3416e-08 1.8300176500776102 2.3417e-08 1.8569217361681798 2.3417999999999998e-08 1.85161044712551 2.3419e-08 1.8787765990832257 2.342e-08 1.782780191394735 2.3421e-08 1.7821492761800124 2.3422e-08 1.8380550304378318 2.3423e-08 1.7584305413404204 2.3424e-08 1.8146581339294685 2.3425e-08 1.709220005567493 2.3426e-08 1.7874828986992328 2.3427e-08 1.7205877312497808 2.3428e-08 1.7967391731326048 2.3429e-08 1.8191232839254592 2.343e-08 1.9009591516080988 2.3431e-08 1.7954718822536662 2.3432e-08 1.748351068068361 2.3433e-08 1.8177918750467246 2.3434e-08 1.8586591009042506 2.3435e-08 1.8374244057775224 2.3436e-08 1.7676772294062146 2.3437e-08 1.8745015214605198 2.3438e-08 1.7646474019817626 2.3439e-08 1.8031119951089685 2.344e-08 1.8914902984185062 2.3440999999999998e-08 1.712231342484748 2.3442e-08 1.8023887908345835 2.3443e-08 1.8901262879420866 2.3443999999999998e-08 1.8946148922267374 2.3445e-08 1.816919258476582 2.3446e-08 1.786488596945011 2.3446999999999998e-08 1.7751495697206168 2.3448e-08 1.7744421949479106 2.3449e-08 1.7634552816408442 2.3449999999999998e-08 1.8180265121871877 2.3451e-08 1.9193372582505386 2.3452e-08 1.6823018315746463 2.3452999999999998e-08 1.7142649101896048 2.3454e-08 1.8382190003498426 2.3455e-08 1.7427245449497133 2.3456e-08 1.7662347694314537 2.3457e-08 1.827773522944805 2.3458e-08 1.7506374100100897 2.3459e-08 1.73703543141305 2.346e-08 1.7520223639658319 2.3461e-08 1.8476057534238446 2.3462e-08 1.8101515514202218 2.3463e-08 1.7176549899304256 2.3464e-08 1.756190786218385 2.3465e-08 1.7449391011283424 2.3466e-08 1.7894586725011747 2.3467e-08 1.7730559105980583 2.3468e-08 1.7846989597330463 2.3469e-08 1.87043793177936 2.347e-08 1.83769535441718 2.3471e-08 1.819679505807486 2.3472e-08 1.7340007018177854 2.3473e-08 1.8213956680802166 2.3474e-08 1.8610853742877436 2.3475e-08 1.863030940595843 2.3475999999999998e-08 1.8038035224017743 2.3477e-08 1.8017080419075224 2.3478e-08 1.8081233294565695 2.3478999999999998e-08 1.7288639865106588 2.348e-08 1.8366879754688863 2.3481e-08 1.7549988062387283 2.3481999999999998e-08 1.8259956273123683 2.3483e-08 1.7197876169067492 2.3484e-08 1.7334924995663679 2.3484999999999998e-08 1.779292308345282 2.3486e-08 1.8087070509991283 2.3487e-08 1.767988609760112 2.3487999999999998e-08 1.8065231243165174 2.3489e-08 1.9318331388208767 2.349e-08 1.7716183079208894 2.3491e-08 1.7692613333049205 2.3492e-08 1.8061198364154187 2.3493e-08 1.7432399285242306 2.3494e-08 1.837970596215171 2.3495e-08 1.8051113827566483 2.3496e-08 1.8875809582996588 2.3497e-08 1.7371723719773082 2.3498e-08 1.6760934227428745 2.3499e-08 1.7760792885135597 2.35e-08 1.8412684964997035 2.3501e-08 1.7612076959415799 2.3502e-08 1.7652910853745623 2.3503e-08 1.7755285557375906 2.3504e-08 1.7575875529413554 2.3505e-08 1.7512378814103908 2.3506e-08 1.8394532129070797 2.3507e-08 1.8155036327268967 2.3508e-08 1.805069621117081 2.3509e-08 1.7997083260888054 2.351e-08 1.844569817963319 2.3510999999999998e-08 1.8089290093912407 2.3512e-08 1.7722832386722027 2.3513e-08 1.858811659174212 2.3513999999999998e-08 1.778918123322471 2.3515e-08 1.8065121170823153 2.3516e-08 1.7852948434819973 2.3516999999999998e-08 1.8331263044982111 2.3518e-08 1.902209592196097 2.3519e-08 1.7787667466925317 2.3519999999999998e-08 1.7824900517262614 2.3521e-08 1.8240676359333452 2.3522e-08 1.7362916197182368 2.3522999999999998e-08 1.7486705815147854 2.3524e-08 1.7864805311777021 2.3525e-08 1.8067462690811416 2.3526e-08 1.8201130843991904 2.3527e-08 1.8507536714233144 2.3528e-08 1.863207060326738 2.3529e-08 1.7776752278211905 2.353e-08 1.8138614561378772 2.3531e-08 1.7681340465796542 2.3532e-08 1.818617054349387 2.3533e-08 1.8547743966819419 2.3534e-08 1.7852110367259542 2.3535e-08 1.7990995380352321 2.3536e-08 1.7932324161436963 2.3537e-08 1.83017747710794 2.3538e-08 1.770928117504585 2.3539e-08 1.8242093897122127 2.354e-08 1.707440662315519 2.3541e-08 1.8109550297605292 2.3542e-08 1.7243537817074825 2.3543e-08 1.92487111460159 2.3544e-08 1.720044196456602 2.3545e-08 1.8128578652882466 2.3545999999999998e-08 1.8765934627777747 2.3547e-08 1.8657679962235503 2.3548e-08 1.7756923063551775 2.3548999999999998e-08 1.8032298931389188 2.355e-08 1.7471351502947716 2.3551e-08 1.888930212347505 2.3551999999999998e-08 1.7941237044010705 2.3553e-08 1.7895052694690186 2.3554e-08 1.763433568084499 2.3554999999999998e-08 1.8260566444169726 2.3556e-08 1.8041547365118242 2.3557e-08 1.7884259649501473 2.3557999999999998e-08 1.8138401260066899 2.3559e-08 1.815865598424736 2.356e-08 1.800293173457829 2.3561e-08 1.9020800768416337 2.3562e-08 1.7730809139388428 2.3563e-08 1.7824938636749732 2.3564e-08 1.7961455383285714 2.3565e-08 1.7494495405184467 2.3566e-08 1.7952788500472239 2.3567e-08 1.8550712727581409 2.3568e-08 1.8002549688724847 2.3569e-08 1.820007081199669 2.357e-08 1.7294611196051606 2.3571e-08 1.8200204306010292 2.3572e-08 1.7529911247291476 2.3573e-08 1.7746177707344806 2.3574e-08 1.7567203925181238 2.3575e-08 1.8933187280504504 2.3576e-08 1.9016547125780914 2.3577e-08 1.8486604724125162 2.3578e-08 1.7744090458291017 2.3579e-08 1.765905345239682 2.358e-08 1.8544908001668308 2.3580999999999998e-08 1.8404567427722918 2.3582e-08 1.788454889879651 2.3583e-08 1.852983346788953 2.3583999999999998e-08 1.8016763008394234 2.3585e-08 1.8158543092704744 2.3586e-08 1.7888640925039263 2.3586999999999998e-08 1.8599151073769336 2.3588e-08 1.8005314678317779 2.3589e-08 1.8495558212484982 2.3589999999999998e-08 1.8909631000327853 2.3591e-08 1.7457495678919641 2.3592e-08 1.8324829557741806 2.3592999999999998e-08 1.8457685191208129 2.3594e-08 1.76360046157786 2.3595e-08 1.807978851033251 2.3595999999999998e-08 1.8080914522457256 2.3597e-08 1.7666360847394562 2.3598e-08 1.7977079329903778 2.3599e-08 1.7918809050337225 2.36e-08 1.7740925245122037 2.3601e-08 1.7602031708233976 2.3602e-08 1.8288036816985196 2.3603e-08 1.760960319833367 2.3604e-08 1.808418148607315 2.3605e-08 1.7611709483192606 2.3606e-08 1.7878878184555596 2.3607e-08 1.7784414052511903 2.3608e-08 1.811875844431461 2.3609e-08 1.771750521937244 2.361e-08 1.7640203146998967 2.3611e-08 1.8979474032550598 2.3612e-08 1.744930016438773 2.3613e-08 1.7390875511436306 2.3614e-08 1.8085626912473738 2.3615e-08 1.8135348164959768 2.3616e-08 1.8091018699621042 2.3617e-08 1.7811055030427991 2.3618e-08 1.8449669140561353 2.3618999999999998e-08 1.8190107875151562 2.362e-08 1.8430536159800004 2.3621e-08 1.8711512718373253 2.3621999999999998e-08 1.754262570373895 2.3623e-08 1.930415091202426 2.3624e-08 1.7796722530437672 2.3624999999999998e-08 1.8178938445451351 2.3626e-08 1.8205960493566193 2.3627e-08 1.8171505538012218 2.3627999999999998e-08 1.8649791158541222 2.3629e-08 1.7404877787628685 2.363e-08 1.7834320710197378 2.3630999999999998e-08 1.765699494629359 2.3632e-08 1.7143395906506982 2.3633e-08 1.8211539594345165 2.3634e-08 1.8407848748423485 2.3635e-08 1.8495982070415988 2.3636e-08 1.7634493748271287 2.3637e-08 1.8455936524888708 2.3638e-08 1.8755932605031207 2.3639e-08 1.865371858900117 2.364e-08 1.8097456646581422 2.3641e-08 1.8045286418472615 2.3642e-08 1.7209813362947386 2.3643e-08 1.7543256874702926 2.3644e-08 1.8009123680637122 2.3645e-08 1.7351917928114717 2.3646e-08 1.8681946316524427 2.3647e-08 1.849320276200512 2.3648e-08 1.8532771539576185 2.3649e-08 1.873042413689055 2.365e-08 1.7865077054559566 2.3651e-08 1.7669295705893133 2.3652e-08 1.8408524264463504 2.3653e-08 1.7143350158369444 2.3653999999999998e-08 1.8043699133562539 2.3655e-08 1.8479381929519585 2.3656e-08 1.8585956770661392 2.3656999999999998e-08 1.8095787032749306 2.3658e-08 1.729215468703236 2.3659e-08 1.7912920166322461 2.3659999999999998e-08 1.825251734301935 2.3661e-08 1.731825105817915 2.3662e-08 1.828553026308702 2.3662999999999998e-08 1.792126276578514 2.3664e-08 1.8207636722921625 2.3665e-08 1.7896366903442862 2.3665999999999998e-08 1.7898123038430807 2.3667e-08 1.7743146894010176 2.3668e-08 1.7893719757292659 2.3669e-08 1.8096809982918398 2.367e-08 1.7968159068727745 2.3671e-08 1.769013044953784 2.3672e-08 1.7703805260427545 2.3673e-08 1.8139012647234651 2.3674e-08 1.802009862436143 2.3675e-08 1.907059968508298 2.3676e-08 1.9008247450301998 2.3677e-08 1.7928613067004817 2.3678e-08 1.819378226526933 2.3679e-08 1.9153784806541618 2.368e-08 1.7235265274344522 2.3681e-08 1.894880738898959 2.3682e-08 1.8577369573780111 2.3683e-08 1.8094716642998856 2.3684e-08 1.785918798451212 2.3685e-08 1.8254863438679783 2.3686e-08 1.7749034322579165 2.3687e-08 1.813103095472854 2.3688e-08 1.7065629597238543 2.3688999999999998e-08 1.7440906831367178 2.369e-08 1.86345662635285 2.3691e-08 1.855155739937583 2.3691999999999998e-08 1.8183984301017269 2.3693e-08 1.7934706202920405 2.3694e-08 1.740543528680754 2.3694999999999998e-08 1.7794240636544305 2.3696e-08 1.799447090709844 2.3697e-08 1.825311253601165 2.3697999999999998e-08 1.8080621812074542 2.3699e-08 1.7928480144463164 2.37e-08 1.7893902381576532 2.3700999999999998e-08 1.8151787539309612 2.3702e-08 1.8281945633363417 2.3703e-08 1.744448128067213 2.3704e-08 1.7600818736203272 2.3705e-08 1.7886532731592484 2.3706e-08 1.8540306999782532 2.3707e-08 1.8441650430537655 2.3708e-08 1.688008084510505 2.3709e-08 1.8411710942792856 2.371e-08 1.8429274443377384 2.3711e-08 1.8479951325123456 2.3712e-08 1.7922665340903134 2.3713e-08 1.767768726282386 2.3714e-08 1.7933143459631347 2.3715e-08 1.8656714013318139 2.3716e-08 1.8506737470111618 2.3717e-08 1.8815476847872006 2.3718e-08 1.7678581446629995 2.3719e-08 1.8089697653710748 2.372e-08 1.7638851265204465 2.3721e-08 1.777897556492468 2.3722e-08 1.8701876608520718 2.3723e-08 1.7611542608783393 2.3723999999999998e-08 1.6889871565255472 2.3725e-08 1.741374088074491 2.3726e-08 1.8181453188106376 2.3726999999999998e-08 1.8471059224122741 2.3728e-08 1.7574679300436828 2.3729e-08 1.8061053970573882 2.3729999999999998e-08 1.7114974686102284 2.3731e-08 1.8641745634951243 2.3732e-08 1.833732381263074 2.3732999999999998e-08 1.8007511514818388 2.3734e-08 1.8008278893314755 2.3735e-08 1.7817736303624827 2.3735999999999998e-08 1.8333708333840721 2.3737e-08 1.7375202010934623 2.3738e-08 1.8104060990467763 2.3739e-08 1.757999420705473 2.374e-08 1.7353346891555044 2.3741e-08 1.727764603480035 2.3742e-08 1.7929526882178553 2.3743e-08 1.8193549442449692 2.3744e-08 1.7913147402334129 2.3745e-08 1.7509948395188613 2.3746e-08 1.8408327314154174 2.3747e-08 1.7507037839885293 2.3748e-08 1.7218998807635775 2.3749e-08 1.6935744488313162 2.375e-08 1.8057110755850738 2.3751e-08 1.8393476859785816 2.3752e-08 1.839565490287541 2.3753e-08 1.831014461758565 2.3754e-08 1.7715564247018731 2.3755e-08 1.7834633166944107 2.3756e-08 1.8079509518568078 2.3757e-08 1.8280597028401375 2.3758e-08 1.8069125897141458 2.3758999999999998e-08 1.8330099981642882 2.376e-08 1.7162358612614375 2.3761e-08 1.8036127052437128 2.3761999999999998e-08 1.7987344122642221 2.3763e-08 1.7651907082366853 2.3764e-08 1.7886508717783498 2.3764999999999998e-08 1.8172005360630537 2.3766e-08 1.7039505961080201 2.3767e-08 1.769230177980552 2.3767999999999998e-08 1.712924528667232 2.3769e-08 1.8268607758466184 2.377e-08 1.8025395157467845 2.3770999999999998e-08 1.8278621276901064 2.3772e-08 1.7640333173141987 2.3773e-08 1.7518367729584448 2.3774e-08 1.7999202814592266 2.3775e-08 1.8268684559010737 2.3776e-08 1.7889685241567037 2.3777e-08 1.855893075698048 2.3778e-08 1.8005417191014155 2.3779e-08 1.8656770144341277 2.378e-08 1.8042181541559117 2.3781e-08 1.8512228183985397 2.3782e-08 1.7729549852566129 2.3783e-08 1.7804351082118075 2.3784e-08 1.8217876714815553 2.3785e-08 1.80990821410088 2.3786e-08 1.8689220191126328 2.3787e-08 1.7832455653501234 2.3788e-08 1.9023518821700858 2.3789e-08 1.77452465342449 2.379e-08 1.8315374721363715 2.3791e-08 1.827714071277365 2.3792e-08 1.8657619656711801 2.3793e-08 1.787152608912322 2.3794e-08 1.7975577307523332 2.3795e-08 1.747859690659724 2.3796e-08 1.7236776562470981 2.3796999999999998e-08 1.8090727505648483 2.3798e-08 1.8092992228835818 2.3799e-08 1.7947516449434 2.3799999999999998e-08 1.7292082189674018 2.3801e-08 1.8396455039596489 2.3802e-08 1.8126390234047758 2.3802999999999998e-08 1.7782548004558898 2.3804e-08 1.8216258307659865 2.3805e-08 1.864841774594298 2.3805999999999998e-08 1.7587243799627226 2.3807e-08 1.7834088050684491 2.3808e-08 1.7653903579734083 2.3808999999999998e-08 1.7958409371455257 2.381e-08 1.812136781684794 2.3811e-08 1.795713767711847 2.3812e-08 1.7391874791568014 2.3813e-08 1.8184216184109425 2.3814e-08 1.847126586666066 2.3815e-08 1.769903012835931 2.3816e-08 1.8045712326345664 2.3817e-08 1.8410143598233528 2.3818e-08 1.8822954068100177 2.3819e-08 1.7344065742912889 2.382e-08 1.8121895142036373 2.3821e-08 1.8800432967259688 2.3822e-08 1.7597222556089054 2.3823e-08 1.8116185266260092 2.3824e-08 1.8056476355146809 2.3825e-08 1.8142208137191234 2.3826e-08 1.764153231379795 2.3827e-08 1.7833306155451274 2.3828e-08 1.8726503811818738 2.3829e-08 1.8492858264462688 2.383e-08 1.7736770633236663 2.3831e-08 1.861812425294841 2.3831999999999998e-08 1.8313221604474024 2.3833e-08 1.8613820472502312 2.3834e-08 1.8339821404478147 2.3834999999999998e-08 1.8288212598413889 2.3836e-08 1.7419865796755065 2.3837e-08 1.7949073020098265 2.3837999999999998e-08 1.7536223180719952 2.3839e-08 1.7285068390980494 2.384e-08 1.8410497725953563 2.3840999999999998e-08 1.708280028654429 2.3842e-08 1.8395218003533396 2.3843e-08 1.7300932821763455 2.3843999999999998e-08 1.7925026676226288 2.3845e-08 1.7928595141994441 2.3846e-08 1.8065256222003254 2.3847e-08 1.899738081636933 2.3848e-08 1.7944576721904109 2.3849e-08 1.8254443462569043 2.385e-08 1.7341134541550876 2.3851e-08 1.853108423462399 2.3852e-08 1.809002586819634 2.3853e-08 1.749977517562716 2.3854e-08 1.8003978501334184 2.3855e-08 1.8290204870237659 2.3856e-08 1.9226665703705423 2.3857e-08 1.8817399377478434 2.3858e-08 1.898151088287048 2.3859e-08 1.7719402314960824 2.386e-08 1.8065612808235072 2.3861e-08 1.8444473303296556 2.3862e-08 1.8734856393278339 2.3863e-08 1.8200801572346568 2.3864e-08 1.7321266812431242 2.3865e-08 1.7860270311971218 2.3866e-08 1.7977807272990927 2.3866999999999998e-08 1.7135678924991777 2.3868e-08 1.88183986892608 2.3869e-08 1.6282779396070115 2.3869999999999998e-08 1.8455753810376252 2.3871e-08 1.7634041411803385 2.3872e-08 1.80665275411493 2.3872999999999998e-08 1.854677963819654 2.3874e-08 1.7349515970480278 2.3875e-08 1.685966162141743 2.3875999999999998e-08 1.7969760709223814 2.3877e-08 1.761237616372799 2.3878e-08 1.826674643113958 2.3878999999999998e-08 1.8271832483814106 2.388e-08 1.7493949727133622 2.3881e-08 1.8794527007198083 2.3882e-08 1.7811593047645902 2.3883e-08 1.7433792643796577 2.3884e-08 1.7993720514553768 2.3885e-08 1.7481000617853895 2.3886e-08 1.826707873844323 2.3887e-08 1.775975755890324 2.3888e-08 1.777235921675799 2.3889e-08 1.8311368707001354 2.389e-08 1.8879361469449376 2.3891e-08 1.7751580282038175 2.3892e-08 1.8130929496594899 2.3893e-08 1.7606394553917575 2.3894e-08 1.8863702025234224 2.3895e-08 1.7659736156029984 2.3896e-08 1.9263532873409008 2.3897e-08 1.8014120595550238 2.3898e-08 1.809928317792476 2.3899e-08 1.820998280232164 2.39e-08 1.7617484353119988 2.3901e-08 1.8672490709804588 2.3901999999999998e-08 1.7762267167112662 2.3903e-08 1.7694571303261104 2.3904e-08 1.7321468894545706 2.3904999999999998e-08 1.8602860964005874 2.3906e-08 1.7778535721469102 2.3907e-08 1.7962612923586163 2.3907999999999998e-08 1.8071546207337306 2.3909e-08 1.8079557343392962 2.391e-08 1.8166572996412695 2.3910999999999998e-08 1.752981744047917 2.3912e-08 1.8149586095655967 2.3913e-08 1.8593362009478414 2.3913999999999998e-08 1.7755829654077802 2.3915e-08 1.8034378828556545 2.3916e-08 1.7615630327735419 2.3917e-08 1.7689115214128697 2.3918e-08 1.7550381556268986 2.3919e-08 1.8243075432510292 2.392e-08 1.8556925315545145 2.3921e-08 1.7985231338407155 2.3922e-08 1.7699764060948275 2.3923e-08 1.726755258123892 2.3924e-08 1.7975476508685537 2.3925e-08 1.7983525976975716 2.3926e-08 1.801859167292755 2.3927e-08 1.911259619695147 2.3928e-08 1.77255688329669 2.3929e-08 1.8217405061165597 2.393e-08 1.8191447394638975 2.3931e-08 1.7827972674296584 2.3932e-08 1.7544019079966056 2.3933e-08 1.7197191805718832 2.3934e-08 1.789860850406302 2.3935e-08 1.8825923247320546 2.3936e-08 1.7634582162526438 2.3936999999999998e-08 1.8240706025672266 2.3938e-08 1.88973146439646 2.3939e-08 1.8069479480963968 2.3939999999999998e-08 1.7688658908237413 2.3941e-08 1.758273954052869 2.3942e-08 1.8164874131435607 2.3942999999999998e-08 1.7997815974796314 2.3944e-08 1.7902717084217519 2.3945e-08 1.8917875185071709 2.3945999999999998e-08 1.7583992654139688 2.3947e-08 1.8332664660093252 2.3948e-08 1.8313994619604852 2.3948999999999998e-08 1.7299865028861077 2.395e-08 1.8236338194104629 2.3951e-08 1.8356177322559875 2.3952e-08 1.7626656536791676 2.3953e-08 1.8098288616980542 2.3954e-08 1.8016472970354305 2.3955e-08 1.779192058592166 2.3956e-08 1.8811365660396868 2.3957e-08 1.8364377727221317 2.3958e-08 1.7946259200749612 2.3959e-08 1.900955864335685 2.396e-08 1.8166780421255089 2.3961e-08 1.7689114636655012 2.3962e-08 1.7894109891499839 2.3963e-08 1.788222311472387 2.3964e-08 1.8707096793702322 2.3965e-08 1.857412622161036 2.3966e-08 1.8218592661737822 2.3967e-08 1.790935523686388 2.3968e-08 1.8135067745139373 2.3969e-08 1.8909128110437863 2.397e-08 1.8152116400004326 2.3971e-08 1.7967121184640045 2.3971999999999998e-08 1.9350532364965414 2.3973e-08 1.8500660248730367 2.3974e-08 1.8066940594492038 2.3974999999999998e-08 1.8001510538564078 2.3976e-08 1.735943212028603 2.3977e-08 1.8599862760848611 2.3977999999999998e-08 1.7576701986564045 2.3979e-08 1.820126735789285 2.398e-08 1.8581897174615263 2.3980999999999998e-08 1.8956078558837985 2.3982e-08 1.8337584768798825 2.3983e-08 1.7704217971727352 2.3983999999999998e-08 1.8101142750081143 2.3985e-08 1.8423541545512387 2.3986e-08 1.8165341352902893 2.3986999999999998e-08 1.7680562553317685 2.3988e-08 1.8559501655125634 2.3989e-08 1.7291968164845175 2.399e-08 1.8132850063750976 2.3991e-08 1.747718981471005 2.3992e-08 1.7407920689445866 2.3993e-08 1.7755216726323513 2.3994e-08 1.7860495151889333 2.3995e-08 1.8051678489348486 2.3996e-08 1.721153430071531 2.3997e-08 1.8066792922598294 2.3998e-08 1.7866220969025572 2.3999e-08 1.7362763930081089 2.4e-08 1.8540406753783067 2.4001e-08 1.7215997507639715 2.4002e-08 1.7834256142892737 2.4003e-08 1.7246297683054856 2.4004e-08 1.800640656632214 2.4005e-08 1.7205069867045726 2.4006e-08 1.805675758438807 2.4007e-08 1.785560430465495 2.4008e-08 1.8028180261133278 2.4009e-08 1.8540000010824267 2.4009999999999998e-08 1.809241953733969 2.4011e-08 1.7948918803713265 2.4012e-08 1.7843007547180971 2.4012999999999998e-08 1.7943192175547398 2.4014e-08 1.8401859368763553 2.4015e-08 1.7250545293958255 2.4015999999999998e-08 1.786743456302484 2.4017e-08 1.818385882557811 2.4018e-08 1.7997725680114969 2.4018999999999998e-08 1.6997265956333407 2.402e-08 1.7191890278091186 2.4021e-08 1.7782252883882945 2.4021999999999998e-08 1.7442679553585891 2.4023e-08 1.862934081089918 2.4024e-08 1.8228311819577692 2.4025e-08 1.798414615482707 2.4026e-08 1.8644651263949172 2.4027e-08 1.7642927090614617 2.4028e-08 1.8619700268774793 2.4029e-08 1.8167477928550793 2.403e-08 1.7954441347280308 2.4031e-08 1.780634738017881 2.4032e-08 1.8367397526578646 2.4033e-08 1.794947136213296 2.4034e-08 1.7590555736404232 2.4035e-08 1.8085230169658582 2.4036e-08 1.8503623362424402 2.4037e-08 1.7723269453122696 2.4038e-08 1.7544475237746662 2.4039e-08 1.806975683125212 2.404e-08 1.8288582807308982 2.4041e-08 1.825357471854952 2.4042e-08 1.8211220706261835 2.4043e-08 1.8078714705589243 2.4044e-08 1.7564424618409142 2.4044999999999998e-08 1.8114380823830611 2.4046e-08 1.8196541492823168 2.4047e-08 1.843786494220586 2.4047999999999998e-08 1.873921123265835 2.4049e-08 1.7385904552664742 2.405e-08 1.703066768530098 2.4050999999999998e-08 1.8083785326905228 2.4052e-08 1.7811440006943422 2.4053e-08 1.775481027457934 2.4053999999999998e-08 1.7616426278552364 2.4055e-08 1.7530569939175276 2.4056e-08 1.7924878474496333 2.4056999999999998e-08 1.7413926823622785 2.4058e-08 1.8082251593489815 2.4059e-08 1.735801518421424 2.406e-08 1.83801050638652 2.4061e-08 1.819156906254203 2.4062e-08 1.8594869358391444 2.4063e-08 1.8010567656780658 2.4064e-08 1.8089551948000628 2.4065e-08 1.7792671568428742 2.4066e-08 1.7559663261825071 2.4067e-08 1.8083597111148215 2.4068e-08 1.763905583340847 2.4069e-08 1.876893327706881 2.407e-08 1.8536956303578755 2.4071e-08 1.8833620263001678 2.4072e-08 1.7827420992822516 2.4073e-08 1.8233599432476717 2.4074e-08 1.8933476135496496 2.4075e-08 1.8076070436333 2.4076e-08 1.8123580453418173 2.4077e-08 1.8020365671890441 2.4078e-08 1.8100209723711451 2.4079e-08 1.8293374979096348 2.4079999999999998e-08 1.801303686230725 2.4081e-08 1.8136156534199444 2.4082e-08 1.7556067949169136 2.4082999999999998e-08 1.8541797308335464 2.4084e-08 1.8408989716640884 2.4085e-08 1.8010473513583316 2.4085999999999998e-08 1.8992043221250579 2.4087e-08 1.7075711100478763 2.4088e-08 1.8980969110215329 2.4088999999999998e-08 1.8455476599736411 2.409e-08 1.834885185403925 2.4091e-08 1.8540032377392481 2.4091999999999998e-08 1.7352525553506073 2.4093e-08 1.754356488394805 2.4094e-08 1.7871011046463081 2.4095e-08 1.8401928969381656 2.4096e-08 1.7971960851784863 2.4097e-08 1.7854060340422362 2.4098e-08 1.7332469611619576 2.4099e-08 1.8167465733790815 2.41e-08 1.784755876595216 2.4101e-08 1.7737330474317015 2.4102e-08 1.7733423243362887 2.4103e-08 1.827721086538519 2.4104e-08 1.8087956615325298 2.4105e-08 1.857359938210975 2.4106e-08 1.8292324453629236 2.4107e-08 1.7571296167194326 2.4108e-08 1.8416959132951431 2.4109e-08 1.8207676056854467 2.411e-08 1.786783956601474 2.4111e-08 1.8286344077947543 2.4112e-08 1.7229984465099868 2.4113e-08 1.8042667758351008 2.4114e-08 1.791709499012683 2.4114999999999998e-08 1.7743535729107358 2.4116e-08 1.7667149400167397 2.4117e-08 1.8033687854714657 2.4117999999999998e-08 1.7934711140403445 2.4119e-08 1.7426440854513479 2.412e-08 1.8134631522814588 2.4120999999999998e-08 1.7947233493442407 2.4122e-08 1.7283122374060653 2.4123e-08 1.7402841758153844 2.4123999999999998e-08 1.7729187985710269 2.4125e-08 1.7558332527559979 2.4126e-08 1.7413408968518873 2.4126999999999998e-08 1.7847479694951653 2.4128e-08 1.828918193783456 2.4129e-08 1.850170085116123 2.413e-08 1.8316702889482719 2.4131e-08 1.8328813485673723 2.4132e-08 1.83759522136776 2.4133e-08 1.843287970621883 2.4134e-08 1.8174270730901134 2.4135e-08 1.7420295966983306 2.4136e-08 1.7641798186737874 2.4137e-08 1.7160302409048274 2.4138e-08 1.7610193176470934 2.4139e-08 1.7601967578373223 2.414e-08 1.829396719580066 2.4141e-08 1.7466167848100318 2.4142e-08 1.7654503566831046 2.4143e-08 1.7661640575822013 2.4144e-08 1.8393295431077337 2.4145e-08 1.8269343770783053 2.4146e-08 1.7068667572001086 2.4147e-08 1.6915023777332843 2.4148e-08 1.7847388344818196 2.4149e-08 1.8297412876324988 2.4149999999999998e-08 1.8535087708257103 2.4151e-08 1.8002696126928035 2.4152e-08 1.857042863795923 2.4152999999999998e-08 1.7323241031015566 2.4154e-08 1.800535495161682 2.4155e-08 1.817612597879815 2.4155999999999998e-08 1.8703292811639414 2.4157e-08 1.7597321636365766 2.4158e-08 1.7192246617534341 2.4158999999999998e-08 1.7856457516723456 2.416e-08 1.7978575370105148 2.4161e-08 1.8324606102986838 2.4161999999999998e-08 1.8431853145178136 2.4163e-08 1.8026423782486092 2.4164e-08 1.741755838081929 2.4164999999999998e-08 1.8082421553253285 2.4166e-08 1.6812945456771058 2.4167e-08 1.82476468020034 2.4168e-08 1.7040610348650362 2.4169e-08 1.8140633417118597 2.417e-08 1.881455826819804 2.4171e-08 1.8331989445003476 2.4172e-08 1.8062957779054785 2.4173e-08 1.7496173509062733 2.4174e-08 1.7500131397945582 2.4175e-08 1.6774318668501846 2.4176e-08 1.7487404136232942 2.4177e-08 1.7122921256281534 2.4178e-08 1.8065721680244886 2.4179e-08 1.8263669597408854 2.418e-08 1.821130584959944 2.4181e-08 1.7823120443746905 2.4182e-08 1.7596184293562256 2.4183e-08 1.8029358433310336 2.4184e-08 1.8234047160150106 2.4185e-08 1.850270222980206 2.4186e-08 1.8142911992956234 2.4187e-08 1.9832721796574555 2.4187999999999998e-08 1.763955051933668 2.4189e-08 1.8026067386818894 2.419e-08 1.8326408535325873 2.4190999999999998e-08 1.83830229047134 2.4192e-08 1.8423074437822238 2.4193e-08 1.8098287015171284 2.4193999999999998e-08 1.8717185856695957 2.4195e-08 1.7601171120553454 2.4196e-08 1.7524671396793283 2.4196999999999998e-08 1.7486763225636834 2.4198e-08 1.8865713428348947 2.4199e-08 1.9085055337299406 2.4199999999999998e-08 1.7580465727051033 2.4201e-08 1.7249707119434066 2.4202e-08 1.8197980587577476 2.4203e-08 1.8232848966313342 2.4204e-08 1.8158260252418024 2.4205e-08 1.8385829163013938 2.4206e-08 1.7553406443679065 2.4207e-08 1.8856632416245436 2.4208e-08 1.830427428017039 2.4209e-08 1.8867291798195482 2.421e-08 1.8924789363950203 2.4211e-08 1.8083891172461928 2.4212e-08 1.783072568734405 2.4213e-08 1.7431144452874288 2.4214e-08 1.8189105885657402 2.4215e-08 1.7724141837994667 2.4216e-08 1.807879260543898 2.4217e-08 1.7727893403041295 2.4218e-08 1.8442316461104697 2.4219e-08 1.7793371407405558 2.422e-08 1.8462478392838801 2.4221e-08 1.7547407025405106 2.4222e-08 1.7893671471093446 2.4222999999999998e-08 1.9054681971564762 2.4224e-08 1.8052591649010747 2.4225e-08 1.8429557155130352 2.4225999999999998e-08 1.897719166178066 2.4227e-08 1.8453195625073948 2.4228e-08 1.8580535569454262 2.4228999999999998e-08 1.8030317178999142 2.423e-08 1.8183556115800712 2.4231e-08 1.7826741605471772 2.4231999999999998e-08 1.8497682955866428 2.4233e-08 1.8364510952939972 2.4234e-08 1.8452806529590804 2.4234999999999998e-08 1.8361833974290978 2.4236e-08 1.7882158145868283 2.4237e-08 1.7662841434830345 2.4238e-08 1.8479040458494755 2.4239e-08 1.8096482965040288 2.424e-08 1.797485316386473 2.4241e-08 1.7863467081328581 2.4242e-08 1.8399610569765765 2.4243e-08 1.8166877090391942 2.4244e-08 1.8666319263609321 2.4245e-08 1.7371562728844303 2.4246e-08 1.8405816080696418 2.4247e-08 1.785714742202979 2.4248e-08 1.8523565914312885 2.4249e-08 1.8652681981382007 2.425e-08 1.8296316816238274 2.4251e-08 1.779262454086384 2.4252e-08 1.805653601413527 2.4253e-08 1.7944946736175655 2.4254e-08 1.8189534211975318 2.4255e-08 1.760232742934655 2.4256e-08 1.7814980662264825 2.4257e-08 1.8216052007371402 2.4257999999999998e-08 1.7194587716898728 2.4259e-08 1.798126294954393 2.426e-08 1.8167960086465305 2.4260999999999998e-08 1.765651312037782 2.4262e-08 1.7394791522794237 2.4263e-08 1.7697595017807526 2.4263999999999998e-08 1.7819022321324463 2.4265e-08 1.8190227852377867 2.4266e-08 1.7624421704122901 2.4266999999999998e-08 1.9074402137137103 2.4268e-08 1.7988500405010666 2.4269e-08 1.95804923279834 2.4269999999999998e-08 1.8170406283996008 2.4271e-08 1.8387727427769525 2.4272e-08 1.8541904381734082 2.4273e-08 1.8086347617559182 2.4274e-08 1.7652846158987032 2.4275e-08 1.7448670892765978 2.4276e-08 1.8434455305987572 2.4277e-08 1.7982314191579427 2.4278e-08 1.8282945743101928 2.4279e-08 1.8617414167309485 2.428e-08 1.8328155770617414 2.4281e-08 1.8287314881698076 2.4282e-08 1.887967864266552 2.4283e-08 1.7164999131861942 2.4284e-08 1.7212400322549806 2.4285e-08 1.753616640334633 2.4286e-08 1.8007715507964313 2.4287e-08 1.7983203981405798 2.4288e-08 1.8017238395217277 2.4289e-08 1.7706765116798078 2.429e-08 1.724575598726508 2.4291e-08 1.8196521135300383 2.4292e-08 1.840003957260229 2.4292999999999998e-08 1.8100893302890664 2.4294e-08 1.7981513105549956 2.4295e-08 1.7800669740321515 2.4295999999999998e-08 1.7871007376546109 2.4297e-08 1.8464087770825746 2.4298e-08 1.8640414378400645 2.4298999999999998e-08 1.7671073108551196 2.43e-08 1.7835237064425082 2.4301e-08 1.7866802462329283 2.4301999999999998e-08 1.8542330726487806 2.4303e-08 1.8370726184792496 2.4304e-08 1.7948204162614203 2.4304999999999998e-08 1.8741888424993465 2.4306e-08 1.802919261638411 2.4307e-08 1.7898996540325227 2.4308e-08 1.8044739384096617 2.4309e-08 1.796473224200437 2.431e-08 1.8112575510481121 2.4311e-08 1.815353135171696 2.4312e-08 1.7548643945849605 2.4313e-08 1.8223088804480947 2.4314e-08 1.7233062557938352 2.4315e-08 1.770230185515101 2.4316e-08 1.8466873102768293 2.4317e-08 1.8193195162001345 2.4318e-08 1.8703552414412459 2.4319e-08 1.842620354126894 2.432e-08 1.8160969177960364 2.4321e-08 1.7969579181961013 2.4322e-08 1.755415901901022 2.4323e-08 1.889723228815265 2.4324e-08 1.8444166080293063 2.4325e-08 1.7573570820839528 2.4326e-08 1.8563528560374507 2.4327e-08 1.827572244211912 2.4327999999999998e-08 1.793287165978874 2.4329e-08 1.7498989902868374 2.433e-08 1.8560894683104987 2.4330999999999998e-08 1.8573358815375083 2.4332e-08 1.7934104809727016 2.4333e-08 1.8876141561168747 2.4333999999999998e-08 1.812091402356244 2.4335e-08 1.8115993538612907 2.4336e-08 1.7688628054918667 2.4336999999999998e-08 1.7737545380988962 2.4338e-08 1.8223288799281856 2.4339e-08 1.7430999483375296 2.4339999999999998e-08 1.8000074935645838 2.4341e-08 1.8295955148017797 2.4342e-08 1.7137345524171246 2.4343e-08 1.903252733031605 2.4344e-08 1.8293179063580163 2.4345e-08 1.8212026396469694 2.4346e-08 1.7663505156397876 2.4347e-08 1.8035653343261557 2.4348e-08 1.8723445019910494 2.4349e-08 1.8822915159320506 2.435e-08 1.8189704378392346 2.4351e-08 1.783007431995662 2.4352e-08 1.8604366843005322 2.4353e-08 1.7902382655218476 2.4354e-08 1.849224291363248 2.4355e-08 1.7821800313888179 2.4356e-08 1.8253530416727362 2.4357e-08 1.8537361724636057 2.4358e-08 1.9103107935338681 2.4359e-08 1.6694528841875298 2.436e-08 1.789111400046547 2.4361e-08 1.757174453380779 2.4362e-08 1.7813123424742787 2.4362999999999998e-08 1.839011953637097 2.4364e-08 1.7925213060496061 2.4365e-08 1.8191660818169684 2.4365999999999998e-08 1.8315118451145356 2.4367e-08 1.7699470717404924 2.4368e-08 1.8338179645575248 2.4368999999999998e-08 1.8236407419208074 2.437e-08 1.780999797073825 2.4371e-08 1.8101542587287152 2.4371999999999998e-08 1.7537459433783618 2.4373e-08 1.8452901813031954 2.4374e-08 1.8223920503746036 2.4374999999999998e-08 1.8905428096473025 2.4376e-08 1.7288034971030466 2.4377e-08 1.7093390857963746 2.4377999999999998e-08 1.8557519848718576 2.4379e-08 1.7274458946699909 2.438e-08 1.7956329434825304 2.4381e-08 1.8480860135855202 2.4382e-08 1.8561425542948005 2.4383e-08 1.8035180589065056 2.4384e-08 1.819209529720775 2.4385e-08 1.7023034213021586 2.4386e-08 1.8071290558583695 2.4387e-08 1.7593244728376878 2.4388e-08 1.8204071554359562 2.4389e-08 1.7596368963573537 2.439e-08 1.842862421846139 2.4391e-08 1.8251975211172975 2.4392e-08 1.7954819446657964 2.4393e-08 1.860836202329863 2.4394e-08 1.7153414813320431 2.4395e-08 1.7815911980692336 2.4396e-08 1.7671146164492835 2.4397e-08 1.779323948420946 2.4398e-08 1.7807633161382068 2.4399e-08 1.9052307224983283 2.44e-08 1.8216878570769983 2.4400999999999998e-08 1.795819449370706 2.4402e-08 1.8220939787838613 2.4403e-08 1.8085026945347051 2.4403999999999998e-08 1.7776137888505934 2.4405e-08 1.7957798125731061 2.4406e-08 1.757391570606824 2.4406999999999998e-08 1.7687235602958054 2.4408e-08 1.7793015704029072 2.4409e-08 1.80650246714681 2.4409999999999998e-08 1.8273783461841167 2.4411e-08 1.7981476287409208 2.4412e-08 1.7006978611614132 2.4412999999999998e-08 1.7992676136770875 2.4414e-08 1.7627278407532259 2.4415e-08 1.6763082714314652 2.4416e-08 1.727014340254437 2.4417e-08 1.8043654584739575 2.4418e-08 1.827254566158704 2.4419e-08 1.8037584387442835 2.442e-08 1.7662824214465125 2.4421e-08 1.7771331238367174 2.4422e-08 1.7734303481507119 2.4423e-08 1.8102186768041388 2.4424e-08 1.8321605061564938 2.4425e-08 1.7488186943096111 2.4426e-08 1.8112029566054202 2.4427e-08 1.7190410268032852 2.4428e-08 1.7900106212876201 2.4429e-08 1.8503393174511074 2.443e-08 1.8032617716420491 2.4431e-08 1.7479924209280633 2.4432e-08 1.8222014821127157 2.4433e-08 1.8045060034734657 2.4434e-08 1.7924653134965467 2.4435e-08 1.771628961182947 2.4435999999999998e-08 1.855774566478446 2.4437e-08 1.836773768277141 2.4438e-08 1.8094564140199814 2.4438999999999998e-08 1.850190876382835 2.444e-08 1.8035490024988705 2.4441e-08 1.8043313954614177 2.4441999999999998e-08 1.742138966769781 2.4443e-08 1.7683846206595941 2.4444e-08 1.7882141936250624 2.4444999999999998e-08 1.798892899370422 2.4446e-08 1.8239033107385911 2.4447e-08 1.8492391018839989 2.4447999999999998e-08 1.8367101078204142 2.4449e-08 1.7774599728352656 2.445e-08 1.8826210188266337 2.4451e-08 1.886202425442853 2.4452e-08 1.806464139267892 2.4453e-08 1.7335320751075263 2.4454e-08 1.7778126204352065 2.4455e-08 1.8048623734485403 2.4456e-08 1.8313864674219997 2.4457e-08 1.7728050085330984 2.4458e-08 1.8166340106052739 2.4459e-08 1.7567802114798352 2.446e-08 1.792329343871642 2.4461e-08 1.8227871559656197 2.4462e-08 1.7849893262736436 2.4463e-08 1.8181989290972151 2.4464e-08 1.76532440526904 2.4465e-08 1.792828501916462 2.4466e-08 1.7998146598362288 2.4467e-08 1.8587874848741768 2.4468e-08 1.790171774138132 2.4469e-08 1.8089647670130917 2.447e-08 1.8038568772730332 2.4470999999999998e-08 1.8197059290996698 2.4472e-08 1.805342739488731 2.4473e-08 1.8023150076713013 2.4473999999999998e-08 1.8286382499074507 2.4475e-08 1.720079727615936 2.4476e-08 1.7680908471856767 2.4476999999999998e-08 1.819423944175546 2.4478e-08 1.8326981334416266 2.4479e-08 1.7900919962152722 2.4479999999999998e-08 1.815937440744054 2.4481e-08 1.740323063028088 2.4482e-08 1.868212360361502 2.4482999999999998e-08 1.714502726363218 2.4484e-08 1.8133888682538932 2.4485e-08 1.8002487741026731 2.4486e-08 1.7303116720793448 2.4487e-08 1.8285769123610667 2.4488e-08 1.7874201969636456 2.4489e-08 1.7943402306973686 2.449e-08 1.7123471607642997 2.4491e-08 1.781921522726482 2.4492e-08 1.7626068339861352 2.4493e-08 1.7657383629233374 2.4494e-08 1.7481536805892581 2.4495e-08 1.8391902720073643 2.4496e-08 1.7817145264085072 2.4497e-08 1.7894536210462444 2.4498e-08 1.7983494179012496 2.4499e-08 1.8286800783674597 2.45e-08 1.787690484171848 2.4501e-08 1.8406585353826463 2.4502e-08 1.7757759232728043 2.4503e-08 1.8744272330637128 2.4504e-08 1.9264605470978502 2.4505e-08 1.75481000365596 2.4505999999999998e-08 1.7982763412275273 2.4507e-08 1.7434610985264434 2.4508e-08 1.7292133310429756 2.4508999999999998e-08 1.7759899855088552 2.451e-08 1.782426428882578 2.4511e-08 1.8107959328264889 2.4511999999999998e-08 1.8258448408660182 2.4513e-08 1.6974054337723747 2.4514e-08 1.7990383744090566 2.4514999999999998e-08 1.8808138024439103 2.4516e-08 1.7235769246695583 2.4517e-08 1.7931536429771737 2.4517999999999998e-08 1.762729489131166 2.4519e-08 1.8402264184343198 2.452e-08 1.7510784663639232 2.4521e-08 1.7549042790507758 2.4522e-08 1.7639480367323523 2.4523e-08 1.8173205459888695 2.4524e-08 1.8302075380303497 2.4525e-08 1.7584523095817035 2.4526e-08 1.8097368539305096 2.4527e-08 1.7559516066845482 2.4528e-08 1.816925538591421 2.4529e-08 1.6959585778417758 2.453e-08 1.7791332933388302 2.4531e-08 1.7458693423010723 2.4532e-08 1.818867791278144 2.4533e-08 1.7201368867487423 2.4534e-08 1.8695192590380585 2.4535e-08 1.7392052286414212 2.4536e-08 1.8061917746661127 2.4537e-08 1.7817639324316852 2.4538e-08 1.7860024002297261 2.4539e-08 1.7358417120153193 2.454e-08 1.8149691008795958 2.4540999999999998e-08 1.7895962710192381 2.4542e-08 1.774989104943739 2.4543e-08 1.7895436406162477 2.4543999999999998e-08 1.777219596410296 2.4545e-08 1.8330597513933389 2.4546e-08 1.7817479565051817 2.4546999999999998e-08 1.7368902145410061 2.4548e-08 1.807533924797061 2.4549e-08 1.7780716178068607 2.4549999999999998e-08 1.8134060606887308 2.4551e-08 1.8774083348526487 2.4552e-08 1.8103998997766206 2.4552999999999998e-08 1.9474275603548845 2.4554e-08 1.784807366464685 2.4555e-08 1.8232524155340382 2.4555999999999998e-08 1.8332865801664804 2.4557e-08 1.8592713153390497 2.4558e-08 1.75038343422722 2.4559e-08 1.6912173744399865 2.456e-08 1.8906476036110242 2.4561e-08 1.7001537529916178 2.4562e-08 1.7750916632884202 2.4563e-08 1.8504891026854549 2.4564e-08 1.8951344625232343 2.4565e-08 1.800531707462732 2.4566e-08 1.7864664129669203 2.4567e-08 1.8448466303787525 2.4568e-08 1.8638543026341459 2.4569e-08 1.7210536452464078 2.457e-08 1.7483239617619677 2.4571e-08 1.745373344329192 2.4572e-08 1.8484981261793085 2.4573e-08 1.805194046504429 2.4574e-08 1.8648065403803924 2.4575e-08 1.8061775183510838 2.4576e-08 1.7143163140619466 2.4577e-08 1.7880116015250032 2.4578e-08 1.7725361203516803 2.4578999999999998e-08 1.7861581906640158 2.458e-08 1.8664536330525203 2.4581e-08 1.8017259239003574 2.4581999999999998e-08 1.8025513637457173 2.4583e-08 1.9268680660572608 2.4584e-08 1.754130704056735 2.4584999999999998e-08 1.7582777166574264 2.4586e-08 1.7408853386547143 2.4587e-08 1.7281014690853909 2.4587999999999998e-08 1.7529997107413602 2.4589e-08 1.8683411241137111 2.459e-08 1.809121916693954 2.4590999999999998e-08 1.7960928709822774 2.4592e-08 1.86384397742383 2.4593e-08 1.686177280140292 2.4594e-08 1.8076827533738198 2.4595e-08 1.8678911822757198 2.4596e-08 1.753461630455341 2.4597e-08 1.771355360197077 2.4598e-08 1.8305556432820098 2.4599e-08 1.8909408462339719 2.46e-08 1.885415179169202 2.4601e-08 1.8495446229510655 2.4602e-08 1.8038476801623289 2.4603e-08 1.8120894483280277 2.4604e-08 1.7712170765933195 2.4605e-08 1.863388853138322 2.4606e-08 1.8051466073130036 2.4607e-08 1.8165666186584382 2.4608e-08 1.7873151216615377 2.4609e-08 1.7531082442212207 2.461e-08 1.8069785061587949 2.4611e-08 1.7908152959221535 2.4612e-08 1.706886832582983 2.4613e-08 1.8192206301869918 2.4613999999999998e-08 1.807562051719336 2.4615e-08 1.8064514262185642 2.4616e-08 1.8038510657781852 2.4616999999999998e-08 1.8151990682621695 2.4618e-08 1.8228753942153937 2.4619e-08 1.721167215294903 2.4619999999999998e-08 1.7643130464300503 2.4621e-08 1.796236424050392 2.4622e-08 1.849992545799628 2.4622999999999998e-08 1.8136525901431335 2.4624e-08 1.7729015878610797 2.4625e-08 1.8283655323791006 2.4625999999999998e-08 1.8061552428822336 2.4627e-08 1.81792617087028 2.4628e-08 1.8187037138270932 2.4629e-08 1.7737728442609746 2.463e-08 1.876187882204681 2.4631e-08 1.7440148537770517 2.4632e-08 1.751533180781659 2.4633e-08 1.744720777257996 2.4634e-08 1.8016175718031942 2.4635e-08 1.7801789079228083 2.4636e-08 1.8168897417371759 2.4637e-08 1.8027350555779378 2.4638e-08 1.8043311327038043 2.4639e-08 1.8123373969854588 2.464e-08 1.868998787747504 2.4641e-08 1.7183725545307142 2.4642e-08 1.806871339659602 2.4643e-08 1.8801122860733197 2.4644e-08 1.8023459304105933 2.4645e-08 1.7990609398943609 2.4646e-08 1.7310726311429974 2.4647e-08 1.8612802729417812 2.4648e-08 1.8822387095011222 2.4648999999999998e-08 1.7977523372393216 2.465e-08 1.8778660997596548 2.4651e-08 1.833598203445391 2.4651999999999998e-08 1.6960095166188691 2.4653e-08 1.7887776318755115 2.4654e-08 1.7960033237714486 2.4654999999999998e-08 1.8204407901012623 2.4656e-08 1.8359372128698404 2.4657e-08 1.8378265489684593 2.4657999999999998e-08 1.783369229859253 2.4659e-08 1.8554258579870029 2.466e-08 1.7926504910988186 2.4660999999999998e-08 1.818848024471777 2.4662e-08 1.7358027145322987 2.4663e-08 1.8572403979781236 2.4664e-08 1.8691938078650858 2.4665e-08 1.769409783112241 2.4666e-08 1.8224605582149622 2.4667e-08 1.8235277378736054 2.4668e-08 1.7615522643633954 2.4669e-08 1.781016384790878 2.467e-08 1.7910463396155665 2.4671e-08 1.8279771706240076 2.4672e-08 1.746051931773353 2.4673e-08 1.7969721406706372 2.4674e-08 1.8493990429838274 2.4675e-08 1.7262584808301904 2.4676e-08 1.8301387498623956 2.4677e-08 1.755024331295392 2.4678e-08 1.8328469304420352 2.4679e-08 1.7033673088279446 2.468e-08 1.798198366092017 2.4681e-08 1.851785380755305 2.4682e-08 1.7539454578099853 2.4683e-08 1.8899123648698224 2.4683999999999998e-08 1.7634689831235308 2.4685e-08 1.8855732118704962 2.4686e-08 1.8431875472202894 2.4686999999999998e-08 1.8275171045568548 2.4688e-08 1.8096499125335543 2.4689e-08 1.8974126290008946 2.4689999999999998e-08 1.9022320962766472 2.4691e-08 1.8450417068199025 2.4692e-08 1.8123945407060167 2.4692999999999998e-08 1.7930393048501652 2.4694e-08 1.7463405214206071 2.4695e-08 1.8469997402045288 2.4695999999999998e-08 1.846460745500698 2.4697e-08 1.8136267288291212 2.4698e-08 1.891903110352087 2.4699e-08 1.8889115282985138 2.47e-08 1.6506334879129871 2.4701e-08 1.8536622385884303 2.4702e-08 1.89642533967593 2.4703e-08 1.7171706349365707 2.4704e-08 1.7751561501983841 2.4705e-08 1.792303392457948 2.4706e-08 1.8989909021985734 2.4707e-08 1.758145086130407 2.4708e-08 1.7938737625725987 2.4709e-08 1.7405115746312068 2.471e-08 1.7651030789175364 2.4711e-08 1.821912821343976 2.4712e-08 1.763430101070486 2.4713e-08 1.7314913095105195 2.4714e-08 1.8139882659368258 2.4715e-08 1.8407192918744286 2.4716e-08 1.7307185953839637 2.4717e-08 1.8664273582855881 2.4718e-08 1.7844129294518027 2.4718999999999998e-08 1.7579111932167049 2.472e-08 1.8520948922560125 2.4721e-08 1.8372328682235268 2.4721999999999998e-08 1.768139540406714 2.4723e-08 1.8490833269896503 2.4724e-08 1.8145069862480359 2.4724999999999998e-08 1.7432959982542213 2.4726e-08 1.8025625395683305 2.4727e-08 1.7983564008966986 2.4727999999999998e-08 1.827606513665563 2.4729e-08 1.8339565402344729 2.473e-08 1.792472297808381 2.4730999999999998e-08 1.7552339404154076 2.4732e-08 1.7455365059721573 2.4733e-08 1.780999358036437 2.4733999999999998e-08 1.7900599590114064 2.4735e-08 1.7598755374742552 2.4736e-08 1.7359042855294118 2.4737e-08 1.775057889385408 2.4738e-08 1.8376340213074995 2.4739e-08 1.8220964693430637 2.474e-08 1.795442538000712 2.4741e-08 1.7773281436719102 2.4742e-08 1.8208270813762424 2.4743e-08 1.7400937565932622 2.4744e-08 1.6710258113669643 2.4745e-08 1.8054218595089304 2.4746e-08 1.8727388933043645 2.4747e-08 1.7200465974537233 2.4748e-08 1.761743915255535 2.4749e-08 1.7751656435441419 2.475e-08 1.8561977043504525 2.4751e-08 1.793085337710266 2.4752e-08 1.814236200005863 2.4753e-08 1.8926575645497319 2.4753999999999998e-08 1.847422717901943 2.4755e-08 1.8538581101081926 2.4756e-08 1.8062091683586898 2.4756999999999998e-08 1.879802731548185 2.4758e-08 1.7511448941588577 2.4759e-08 1.797392268894158 2.4759999999999998e-08 1.7947972060539856 2.4761e-08 1.770495630769593 2.4762e-08 1.7824698228874472 2.4762999999999998e-08 1.7862984298710003 2.4764e-08 1.8303457932459302 2.4765e-08 1.8032231209238632 2.4765999999999998e-08 1.8244885424258162 2.4767e-08 1.8308482446452714 2.4768e-08 1.803139200769328 2.4768999999999998e-08 1.7172943905346705 2.477e-08 1.86033745528702 2.4771e-08 1.9230392558170515 2.4772e-08 1.835937251906169 2.4773e-08 1.808563122468672 2.4774e-08 1.7796675539655773 2.4775e-08 1.8129582655960108 2.4776e-08 1.7788608189375028 2.4777e-08 1.7869282496926564 2.4778e-08 1.7725336192306456 2.4779e-08 1.7204212203995641 2.478e-08 1.825713926270412 2.4781e-08 1.8300756195264336 2.4782e-08 1.7803009893071746 2.4783e-08 1.848798169294596 2.4784e-08 1.8179090337246033 2.4785e-08 1.82697592384311 2.4786e-08 1.6825797496566457 2.4787e-08 1.817218164355459 2.4788e-08 1.7526110337379524 2.4789e-08 1.8152732958097804 2.479e-08 1.8402866967763845 2.4791e-08 1.8215246138015568 2.4791999999999998e-08 1.8359121972649466 2.4793e-08 1.7567027568618083 2.4794e-08 1.698282487284757 2.4794999999999998e-08 1.7916686891223215 2.4796e-08 1.8187714166722837 2.4797e-08 1.8090735699144167 2.4797999999999998e-08 1.8549759318637276 2.4799e-08 1.8641625211380741 2.48e-08 1.7890289910905328 2.4800999999999998e-08 1.7908542295059853 2.4802e-08 1.8278374653540328 2.4803e-08 1.7622120194544655 2.4803999999999998e-08 1.8313188143643326 2.4805e-08 1.7802204213384327 2.4806e-08 1.8233727060807192 2.4807e-08 1.8144615549711636 2.4808e-08 1.800139086375445 2.4809e-08 1.820620872591349 2.481e-08 1.7865146485416135 2.4811e-08 1.854120511877907 2.4812e-08 1.9249782998905567 2.4813e-08 1.7298909905146467 2.4814e-08 1.7840803230579838 2.4815e-08 1.8309868701203291 2.4816e-08 1.811990268493494 2.4817e-08 1.8487289677392675 2.4818e-08 1.8727676255389423 2.4819e-08 1.8116990002422062 2.482e-08 1.78830741049436 2.4821e-08 1.7418048144284344 2.4822e-08 1.7667672555598566 2.4823e-08 1.775151547358618 2.4824e-08 1.8038449312070106 2.4825e-08 1.727092755644634 2.4826e-08 1.7971771944191675 2.4826999999999998e-08 1.799319544618934 2.4828e-08 1.825297575554944 2.4829e-08 1.7537891017543836 2.4829999999999998e-08 1.713994204028837 2.4831e-08 1.7590706092721988 2.4832e-08 1.858481886362233 2.4832999999999998e-08 1.8601026142296564 2.4834e-08 1.7523358177729116 2.4835e-08 1.8457159841186304 2.4835999999999998e-08 1.7814111601554552 2.4837e-08 1.7809408089726895 2.4838e-08 1.753968166554295 2.4838999999999998e-08 1.7575840267181262 2.484e-08 1.7896566763029873 2.4841e-08 1.8221684418483797 2.4842e-08 1.8139861759003915 2.4843e-08 1.7407239812576072 2.4844e-08 1.674507234445444 2.4845e-08 1.8302993782133195 2.4846e-08 1.8566784146089539 2.4847e-08 1.7775412413602327 2.4848e-08 1.8454581426728873 2.4849e-08 1.9029647233496485 2.485e-08 1.83743684357466 2.4851e-08 1.7908098924660625 2.4852e-08 1.8789927712746544 2.4853e-08 1.827333172014334 2.4854e-08 1.8018965684959516 2.4855e-08 1.7631743577272483 2.4856e-08 1.805499572888711 2.4857e-08 1.7705077217992178 2.4858e-08 1.818474608167041 2.4859e-08 1.7884481771276264 2.486e-08 1.8699987246229406 2.4861e-08 1.7162378379467678 2.4861999999999998e-08 1.8161915358437566 2.4863e-08 1.76176318936366 2.4864e-08 1.763861494658665 2.4864999999999998e-08 1.7841848905708504 2.4866e-08 1.7928331442348144 2.4867e-08 1.7430704092011393 2.4867999999999998e-08 1.8646068137649747 2.4869e-08 1.761964998652813 2.487e-08 1.8770304479056317 2.4870999999999998e-08 1.807563018349868 2.4872e-08 1.8711271456541743 2.4873e-08 1.8640755710890307 2.4873999999999998e-08 1.7883441764176293 2.4875e-08 1.7983656816259694 2.4876e-08 1.7269101258647837 2.4877e-08 1.8545344963218002 2.4878e-08 1.8178067601220782 2.4879e-08 1.8184717794305099 2.488e-08 1.816341126961578 2.4881e-08 1.8589460640829005 2.4882e-08 1.8217426601820825 2.4883e-08 1.777577891691394 2.4884e-08 1.7753937752921005 2.4885e-08 1.798052474281862 2.4886e-08 1.8322538269162356 2.4887e-08 1.778681715353135 2.4888e-08 1.8448407320387294 2.4889e-08 1.7522134507636986 2.489e-08 1.874944420640578 2.4891e-08 1.8418289763654414 2.4892e-08 1.7908873078431278 2.4893e-08 1.7215021658580443 2.4894e-08 1.7745207314968972 2.4895e-08 1.8310780591753726 2.4896e-08 1.8104565242598631 2.4896999999999998e-08 1.8314625433337202 2.4898e-08 1.8071871195316835 2.4899e-08 1.807995356736391 2.4899999999999998e-08 1.7684887770973985 2.4901e-08 1.7318071266197743 2.4902e-08 1.7428363847917288 2.4902999999999998e-08 1.8047415629214565 2.4904e-08 1.7193452389853725 2.4905e-08 1.7286394358864083 2.4905999999999998e-08 1.774506288936339 2.4907e-08 1.8408968953354865 2.4908e-08 1.8106055855557277 2.4908999999999998e-08 1.8384621888563988 2.491e-08 1.8142038332677006 2.4911e-08 1.8187764094973882 2.4911999999999998e-08 1.8119162953386567 2.4913e-08 1.7581489647890334 2.4914e-08 1.8904826774136103 2.4915e-08 1.8807674239027603 2.4916e-08 1.8649937786429498 2.4917e-08 1.7622641493649551 2.4918e-08 1.712730205860759 2.4919e-08 1.819785258454433 2.492e-08 1.7818207799125092 2.4921e-08 1.7530799431476767 2.4922e-08 1.8356402584781877 2.4923e-08 1.8087064320016446 2.4924e-08 1.772239744446447 2.4925e-08 1.710550444963062 2.4926e-08 1.8216846835842053 2.4927e-08 1.7707608555895555 2.4928e-08 1.8586342078487683 2.4929e-08 1.9181920408442137 2.493e-08 1.8408957526804448 2.4931e-08 1.8599631472269889 2.4931999999999998e-08 1.7982855603134584 2.4933e-08 1.8445790354760114 2.4934e-08 1.8048157264568165 2.4934999999999998e-08 1.8664471295735874 2.4936e-08 1.7215978033367816 2.4937e-08 1.8188811970556151 2.4937999999999998e-08 1.7683965607873284 2.4939e-08 1.7203633581559183 2.494e-08 1.7887638832000083 2.4940999999999998e-08 1.7158358509694294 2.4942e-08 1.783524609975516 2.4943e-08 1.8133286661689427 2.4943999999999998e-08 1.820742993677016 2.4945e-08 1.879429755443623 2.4946e-08 1.7336121170342136 2.4946999999999998e-08 1.8606000445718438 2.4948e-08 1.8392654802825326 2.4949e-08 1.8495121596309059 2.495e-08 1.8657689789692908 2.4951e-08 1.8596342416157872 2.4952e-08 1.8238834431288804 2.4953e-08 1.807555075412302 2.4954e-08 1.906339541441223 2.4955e-08 1.7758133122050923 2.4956e-08 1.852331693477666 2.4957e-08 1.806124909810705 2.4958e-08 1.7654854805868836 2.4959e-08 1.7739304033296586 2.496e-08 1.8003425856479882 2.4961e-08 1.808113736516746 2.4962e-08 1.740768986310246 2.4963e-08 1.6969432310136519 2.4964e-08 1.8147534500271647 2.4965e-08 1.7654431847409344 2.4966e-08 1.7300495713374677 2.4966999999999998e-08 1.7957348599760568 2.4968e-08 1.8495342223322335 2.4969e-08 1.822423443997831 2.4969999999999998e-08 1.7748690106971217 2.4971e-08 1.8659482967866317 2.4972e-08 1.7422016383421928 2.4972999999999998e-08 1.8296229224372382 2.4974e-08 1.7394784913868393 2.4975e-08 1.806604774831814 2.4975999999999998e-08 1.856655045376958 2.4977e-08 1.8457313018074921 2.4978e-08 1.7858014014812824 2.4978999999999998e-08 1.8630963543304717 2.498e-08 1.8659478784604753 2.4981e-08 1.843621312880972 2.4981999999999998e-08 1.8246737299271572 2.4983e-08 1.8193467937072474 2.4984e-08 1.7816844847148439 2.4985e-08 1.7604286441575834 2.4986e-08 1.7707616177047882 2.4987e-08 1.7632121631083193 2.4988e-08 1.7169878356225632 2.4989e-08 1.790748653166728 2.499e-08 1.7110883928282472 2.4991e-08 1.7466347431605607 2.4992e-08 1.8208618463935569 2.4993e-08 1.7776418315701112 2.4994e-08 1.7137736235496004 2.4995e-08 1.8047379507464258 2.4996e-08 1.7931867840236848 2.4997e-08 1.7579409559640145 2.4998e-08 1.8744326539988432 2.4999e-08 1.7502706380583084 2.5e-08 1.8064047483475607 2.5001e-08 1.7698241056679012 2.5002e-08 1.8339849885298516 2.5003e-08 1.8160905669403689 2.5004e-08 1.83269915781899 2.5004999999999998e-08 1.7526714538561814 2.5006e-08 1.7979765939598666 2.5007e-08 1.720360346607213 2.5007999999999998e-08 1.8234668802567613 2.5009e-08 1.8662865681827099 2.501e-08 1.7639707665093713 2.5010999999999998e-08 1.792185732953423 2.5012e-08 1.839811951814444 2.5013e-08 1.791145984401318 2.5013999999999998e-08 1.7105146208611977 2.5015e-08 1.7806482413061577 2.5016e-08 1.774875883660172 2.5016999999999998e-08 1.7944802927951555 2.5018e-08 1.8305711324392937 2.5019e-08 1.7717564847948473 2.502e-08 1.7591793063862575 2.5021e-08 1.8960360951931967 2.5022e-08 1.7758178149348816 2.5023e-08 1.772093632495321 2.5024e-08 1.7361856330286758 2.5025e-08 1.8403028395255976 2.5026e-08 1.9009497280783019 2.5027e-08 1.81450890605881 2.5028e-08 1.8208858540070503 2.5029e-08 1.728393637954487 2.503e-08 1.8430204887924009 2.5031e-08 1.8360835003671048 2.5032e-08 1.6909175103080312 2.5033e-08 1.864629317864516 2.5034e-08 1.7457479403538587 2.5035e-08 1.8801724987676998 2.5036e-08 1.8472692444014718 2.5037e-08 1.9039121392798897 2.5038e-08 1.8764752974955314 2.5039e-08 1.6615057573248744 2.5039999999999998e-08 1.794727560472079 2.5041e-08 1.7747913665487305 2.5042e-08 1.799793286768484 2.5042999999999998e-08 1.745667725028269 2.5044e-08 1.787517507100595 2.5045e-08 1.7142193040294191 2.5045999999999998e-08 1.8024811349325185 2.5047e-08 1.8165230985951282 2.5048e-08 1.8372964705740047 2.5048999999999998e-08 1.8122687430380653 2.505e-08 1.870146092193319 2.5051e-08 1.8032913030275455 2.5051999999999998e-08 1.9290046799462144 2.5053e-08 1.8440216572068746 2.5054e-08 1.8308393768411584 2.5055e-08 1.7462327486895095 2.5056e-08 1.7600435823939447 2.5057e-08 1.7504867260247323 2.5058e-08 1.7703600267688362 2.5059e-08 1.803805404903207 2.506e-08 1.7861711296810177 2.5061e-08 1.6894298216748425 2.5062e-08 1.789428283903924 2.5063e-08 1.7820221244390655 2.5064e-08 1.6948100882773387 2.5065e-08 1.8132449785425813 2.5066e-08 1.6868917377093513 2.5067e-08 1.7828694297743297 2.5068e-08 1.7604340362019153 2.5069e-08 1.8572777728398688 2.507e-08 1.8611524645377173 2.5071e-08 1.8323880303168514 2.5072e-08 1.8235259695273536 2.5073e-08 1.8206827873504934 2.5074e-08 1.8488068741376444 2.5074999999999998e-08 1.7433734669011065 2.5076e-08 1.8126786214285906 2.5077e-08 1.7032677679613348 2.5077999999999998e-08 1.800952303747895 2.5079e-08 1.809663334351615 2.508e-08 1.7430185496618953 2.5080999999999998e-08 1.7797358940663024 2.5082e-08 1.776725110808263 2.5083e-08 1.8679764159732908 2.5083999999999998e-08 1.802534615017748 2.5085e-08 1.7616124422557335 2.5086e-08 1.771228781556664 2.5086999999999998e-08 1.7905894917942884 2.5088e-08 1.7472702564921512 2.5089e-08 1.7862715064339578 2.509e-08 1.7786573951862665 2.5091e-08 1.849560430393828 2.5092e-08 1.8232946803346473 2.5093e-08 1.8548108929255458 2.5094e-08 1.697398766615618 2.5095e-08 1.7613547444491369 2.5096e-08 1.7306685067883367 2.5097e-08 1.7744174057299757 2.5098e-08 1.756506738030786 2.5099e-08 1.7678087854433333 2.51e-08 1.817642886138993 2.5101e-08 1.8350525306816472 2.5102e-08 1.6756113315072807 2.5103e-08 1.8587956361525926 2.5104e-08 1.7730225559707156 2.5105e-08 1.8344447698961976 2.5106e-08 1.7879119760728064 2.5107e-08 1.8061940406478265 2.5108e-08 1.770138746268801 2.5109e-08 1.796849121880418 2.5109999999999998e-08 1.758229917088174 2.5111e-08 1.823464528315665 2.5112e-08 1.7882080319571896 2.5112999999999998e-08 1.81824653188899 2.5114e-08 1.8447746530962128 2.5115e-08 1.8432019574815794 2.5115999999999998e-08 1.818471618852607 2.5117e-08 1.786892177049766 2.5118e-08 1.7876244022674095 2.5118999999999998e-08 1.7998309777836448 2.512e-08 1.8874862880065286 2.5121e-08 1.7976488949380485 2.5121999999999998e-08 1.8397361689093183 2.5123e-08 1.8185265977747205 2.5124e-08 1.9334702326989084 2.5124999999999998e-08 1.7170759913980682 2.5126e-08 1.802384138956829 2.5127e-08 1.8234635731792492 2.5128e-08 1.7403659872845074 2.5129e-08 1.7384701080110205 2.513e-08 1.7262447270735386 2.5131e-08 1.7902550013462366 2.5132e-08 1.8186758333868769 2.5133e-08 1.8754605676002782 2.5134e-08 1.862166033636254 2.5135e-08 1.83872536207793 2.5136e-08 1.809184779369014 2.5137e-08 1.8211914273852499 2.5138e-08 1.7395232922282684 2.5139e-08 1.8789487534722766 2.514e-08 1.7991097296440794 2.5141e-08 1.8250312226311767 2.5142e-08 1.8704140081592528 2.5143e-08 1.7354595920122144 2.5144e-08 1.837913118510718 2.5144999999999998e-08 1.6948650560242409 2.5146e-08 1.7538541791179005 2.5147e-08 1.7662885507633954 2.5147999999999998e-08 1.8120119062417153 2.5149e-08 1.809562613703369 2.515e-08 1.829608344112712 2.5150999999999998e-08 1.6881346836892668 2.5152e-08 1.7585386990207683 2.5153e-08 1.8327304313831916 2.5153999999999998e-08 1.792432111395797 2.5155e-08 1.8000490788122052 2.5156e-08 1.7322266060503497 2.5156999999999998e-08 1.8119894446666844 2.5158e-08 1.796011570648911 2.5159e-08 1.8104213712170314 2.5159999999999998e-08 1.8450970440997525 2.5161e-08 1.7461859788965617 2.5162e-08 1.8130911651348152 2.5163e-08 1.759132053070273 2.5164e-08 1.810379505393691 2.5165e-08 1.7986025224829965 2.5166e-08 1.824315766970572 2.5167e-08 1.8235116185456208 2.5168e-08 1.7459256625076442 2.5169e-08 1.735309132879306 2.517e-08 1.7820545955142857 2.5171e-08 1.8317427963883708 2.5172e-08 1.7737394758487437 2.5173e-08 1.8154606412802055 2.5174e-08 1.8191327587979793 2.5175e-08 1.7978584656639698 2.5176e-08 1.8737694341635343 2.5177e-08 1.8063772280402908 2.5178e-08 1.8393215467050046 2.5179e-08 1.893193551259433 2.518e-08 1.793199346846321 2.5181e-08 1.7586878257974767 2.5182e-08 1.7419697551489115 2.5182999999999998e-08 1.873750059627778 2.5184e-08 1.753692709773918 2.5185e-08 1.8455945313224296 2.5185999999999998e-08 1.739492765351973 2.5187e-08 1.8048778261207352 2.5188e-08 1.7601589847100338 2.5188999999999998e-08 1.7869081867196248 2.519e-08 1.7719197301973317 2.5191e-08 1.8722712055680584 2.5191999999999998e-08 1.808548680342116 2.5193e-08 1.82834921538041 2.5194e-08 1.8676439280917259 2.5194999999999998e-08 1.7647393140318752 2.5196e-08 1.818070858989717 2.5197e-08 1.8242154991555464 2.5198e-08 1.7830458566952008 2.5199e-08 1.8155059292892928 2.52e-08 1.8280202111738963 2.5201e-08 1.8176643845561573 2.5202e-08 1.8225705118364979 2.5203e-08 1.8706652903232348 2.5204e-08 1.7854835588126892 2.5205e-08 1.7982276342680752 2.5206e-08 1.8142615019097739 2.5207e-08 1.7673922512813833 2.5208e-08 1.8326321953667868 2.5209e-08 1.8861572521266894 2.521e-08 1.8074339455773394 2.5211e-08 1.7869131301258911 2.5212e-08 1.7988271503861863 2.5213e-08 1.8085276231498786 2.5214e-08 1.7493620877825125 2.5215e-08 1.8399678899915608 2.5216e-08 1.7442651843342976 2.5217e-08 1.9376750592852081 2.5217999999999998e-08 1.7844060552436758 2.5219e-08 1.835831981154019 2.522e-08 1.7509364904551652 2.5220999999999998e-08 1.8412624682740395 2.5222e-08 1.8056493804458424 2.5223e-08 1.7848147185879282 2.5223999999999998e-08 1.8837878455099746 2.5225e-08 1.7915851924365034 2.5226e-08 1.8491815977406427 2.5226999999999998e-08 1.8076789676981224 2.5228e-08 1.795805137996842 2.5229e-08 1.8649753181192361 2.5229999999999998e-08 1.7767611233642597 2.5231e-08 1.7508329386316794 2.5232e-08 1.8727052364482493 2.5233e-08 1.8398436215027667 2.5234e-08 1.7783136261609305 2.5235e-08 1.8587097240874284 2.5236e-08 1.7311572735687872 2.5237e-08 1.899932757322867 2.5238e-08 1.7972564052318276 2.5239e-08 1.7431967833243998 2.524e-08 1.7958909869936486 2.5241e-08 1.7842521430009608 2.5242e-08 1.7831591356125958 2.5243e-08 1.7922994351755726 2.5244e-08 1.784939168510792 2.5245e-08 1.7738204452280193 2.5246e-08 1.7708406450093315 2.5247e-08 1.6578969112580206 2.5248e-08 1.7471902926414038 2.5249e-08 1.9092260013269045 2.525e-08 1.864756161562232 2.5251e-08 1.7755985506175664 2.5252e-08 1.790268521922093 2.5252999999999998e-08 1.6971795400465253 2.5254e-08 1.7757121311250592 2.5255e-08 1.8144475812365997 2.5255999999999998e-08 1.7970858916979873 2.5257e-08 1.788145824894498 2.5258e-08 1.786120475098682 2.5258999999999998e-08 1.8032698200798376 2.526e-08 1.7855971802319917 2.5261e-08 1.7859069737942947 2.5261999999999998e-08 1.7745726423256283 2.5263e-08 1.7115231213925899 2.5264e-08 1.7986019032248326 2.5264999999999998e-08 1.8254508242105347 2.5266e-08 1.8682689985578953 2.5267e-08 1.7478925228614102 2.5268e-08 1.7601744736107205 2.5269e-08 1.784284356091086 2.527e-08 1.7760119938863186 2.5271e-08 1.7010483457403207 2.5272e-08 1.8318449259976273 2.5273e-08 1.7505732691227935 2.5274e-08 1.885821825530754 2.5275e-08 1.7816999866317595 2.5276e-08 1.8183934056418096 2.5277e-08 1.878477029327106 2.5278e-08 1.8405623491442118 2.5279e-08 1.820884192358896 2.528e-08 1.8310611384747024 2.5281e-08 1.785477279039057 2.5282e-08 1.8265390334762734 2.5283e-08 1.8692898880969038 2.5284e-08 1.7922606985084928 2.5285e-08 1.790882387944604 2.5286e-08 1.7779549453466665 2.5287e-08 1.6902928396634314 2.5287999999999998e-08 1.793695304816566 2.5289e-08 1.7647136143583444 2.529e-08 1.77562595022411 2.5290999999999998e-08 1.7621567389451247 2.5292e-08 1.7062047399770832 2.5293e-08 1.8177068613778145 2.5293999999999998e-08 1.8547491739259074 2.5295e-08 1.8705083732678953 2.5296e-08 1.7434094404747926 2.5296999999999998e-08 1.7778900070893946 2.5298e-08 1.837513837289914 2.5299e-08 1.8893984126018122 2.5299999999999998e-08 1.8355705482868128 2.5301e-08 1.8621779361307447 2.5302e-08 1.7899871072679483 2.5302999999999998e-08 1.7435145655025428 2.5304e-08 1.8023893461666192 2.5305e-08 1.8428547811138867 2.5306e-08 1.738238202688382 2.5307e-08 1.8007792928209099 2.5308e-08 1.8159841328349708 2.5309e-08 1.8089360516972894 2.531e-08 1.7358552202352528 2.5311e-08 1.7962100726145955 2.5312e-08 1.711251748933271 2.5313e-08 1.7278480845933892 2.5314e-08 1.7343775411602258 2.5315e-08 1.8058897639462002 2.5316e-08 1.733607973708015 2.5317e-08 1.813471124414837 2.5318e-08 1.8220899000597317 2.5319e-08 1.6978792645104392 2.532e-08 1.7924499477765237 2.5321e-08 1.8314231168875608 2.5322e-08 1.7884206518019545 2.5322999999999998e-08 1.8045020036389 2.5324e-08 1.80963394373563 2.5325e-08 1.7670999375343486 2.5325999999999998e-08 1.8538763248999968 2.5327e-08 1.740531508221297 2.5328e-08 1.8223155946099383 2.5328999999999998e-08 1.9256942054999828 2.533e-08 1.6984588659873519 2.5331e-08 1.7921589388570118 2.5331999999999998e-08 1.77134455550768 2.5333e-08 1.835784801922024 2.5334e-08 1.8007510717702753 2.5334999999999998e-08 1.81041376163292 2.5336e-08 1.7827383534578363 2.5337e-08 1.819454948762022 2.5337999999999998e-08 1.7844482646259952 2.5339e-08 1.8771959204813573 2.534e-08 1.8944328452778718 2.5341e-08 1.7730054498900607 2.5342e-08 1.792089861871155 2.5343e-08 1.6961960813434032 2.5344e-08 1.8522599592538023 2.5345e-08 1.8198500986305945 2.5346e-08 1.8291211320767122 2.5347e-08 1.7534794448183968 2.5348e-08 1.7640052208769088 2.5349e-08 1.7916238721600521 2.535e-08 1.836225798641663 2.5351e-08 1.8037009095269558 2.5352e-08 1.7108460391599314 2.5353e-08 1.8285384360324168 2.5354e-08 1.785983607766538 2.5355e-08 1.814275250383553 2.5356e-08 1.845781479780566 2.5357e-08 1.8058461579209468 2.5357999999999998e-08 1.8922526178268548 2.5359e-08 1.8012877476791243 2.536e-08 1.7254372724210623 2.5360999999999998e-08 1.726052308191609 2.5362e-08 1.890826090510271 2.5363e-08 1.7641489178290874 2.5363999999999998e-08 1.8408191793759532 2.5365e-08 1.805572064691022 2.5366e-08 1.8648362279580075 2.5366999999999998e-08 1.8118684297869496 2.5368e-08 1.8188081906412168 2.5369e-08 1.7426026515674022 2.5369999999999998e-08 1.821937314357545 2.5371e-08 1.9200475898137868 2.5372e-08 1.8343891013674343 2.5372999999999998e-08 1.7862436874004102 2.5374e-08 1.8302049231781987 2.5375e-08 1.725951451362664 2.5376e-08 1.7950734508184836 2.5377e-08 1.830338857245356 2.5378e-08 1.736683238035163 2.5379e-08 1.768856067870592 2.538e-08 1.8123602419986666 2.5381e-08 1.8910876894439974 2.5382e-08 1.8274940683375402 2.5383e-08 1.7715842126984656 2.5384e-08 1.845316332463706 2.5385e-08 1.798533504656603 2.5386e-08 1.8234949136490386 2.5387e-08 1.8625614038592984 2.5388e-08 1.7946825188792 2.5389e-08 1.845734552078893 2.539e-08 1.8058129771399798 2.5391e-08 1.7153769652987982 2.5392e-08 1.8141218454623276 2.5393e-08 1.760944966528784 2.5394e-08 1.8471312955356753 2.5395e-08 1.7796947712089564 2.5395999999999998e-08 1.7273333300126759 2.5397e-08 1.88699480919939 2.5398e-08 1.7234146670855006 2.5398999999999998e-08 1.8919164293817683 2.54e-08 1.7641566733965466 2.5401e-08 1.7625423583052726 2.5401999999999998e-08 1.750951501099223 2.5403e-08 1.852209122649256 2.5404e-08 1.7825158257074227 2.5404999999999998e-08 1.8463109629060637 2.5406e-08 1.8009784489340657 2.5407e-08 1.808078975276948 2.5407999999999998e-08 1.804572005612224 2.5409e-08 1.8490716947877823 2.541e-08 1.7296779190761382 2.5411e-08 1.8211569904583376 2.5412e-08 1.7176641447025647 2.5413e-08 1.9067339403376589 2.5414e-08 1.7938378155222165 2.5415e-08 1.7778296439760959 2.5416e-08 1.7794900397149132 2.5417e-08 1.8725644180329697 2.5418e-08 1.738202819241879 2.5419e-08 1.7973733282942745 2.542e-08 1.7518002768847283 2.5421e-08 1.7722946096289622 2.5422e-08 1.8340138401397519 2.5423e-08 1.8049262706035083 2.5424e-08 1.8551590440854075 2.5425e-08 1.8784583140948456 2.5426e-08 1.7619211587385222 2.5427e-08 1.828691763712811 2.5428e-08 1.716036939118766 2.5429e-08 1.811116353477549 2.543e-08 1.829254967554019 2.5430999999999998e-08 1.79925385703827 2.5432e-08 1.8135546996488903 2.5433e-08 1.8294081309034584 2.5433999999999998e-08 1.7912539719517089 2.5435e-08 1.8069470969695829 2.5436e-08 1.8736522993348856 2.5436999999999998e-08 1.712062070814064 2.5438e-08 1.7875405746418738 2.5439e-08 1.8376215844386081 2.5439999999999998e-08 1.881525383249116 2.5441e-08 1.8600514270551134 2.5442e-08 1.8652966576953687 2.5442999999999998e-08 1.7932658141320548 2.5444e-08 1.8659547085013672 2.5445e-08 1.7689306009847998 2.5446e-08 1.7212437727298466 2.5447e-08 1.8284078525512808 2.5448e-08 1.8079535079859568 2.5449e-08 1.8519134548980587 2.545e-08 1.7876394907778421 2.5451e-08 1.7595316663390166 2.5452e-08 1.7751532875476053 2.5453e-08 1.8246817807382696 2.5454e-08 1.7978371948168368 2.5455e-08 1.7843861779148158 2.5456e-08 1.789842054638387 2.5457e-08 1.762231801436983 2.5458e-08 1.7893238544921952 2.5459e-08 1.7392986983730212 2.546e-08 1.8588230500182337 2.5461e-08 1.7052586616603311 2.5462e-08 1.7542426713103196 2.5463e-08 1.8969212218549802 2.5464e-08 1.744304156953897 2.5465e-08 1.851602345532138 2.5465999999999998e-08 1.9438908205000323 2.5467e-08 1.9407116147822199 2.5468e-08 1.9032111103676934 2.5468999999999998e-08 1.8087741130189754 2.547e-08 1.7619992655227323 2.5471e-08 1.7885859289957877 2.5471999999999998e-08 1.7491358459729203 2.5473e-08 1.7979979912316026 2.5474e-08 1.7372845787549531 2.5474999999999998e-08 1.7749258427256813 2.5476e-08 1.8436925714664045 2.5477e-08 1.8173505905660974 2.5477999999999998e-08 1.7618044712288594 2.5479e-08 1.75120943949357 2.548e-08 1.7717339218495323 2.5480999999999998e-08 1.791743055407094 2.5482e-08 1.8175638758246466 2.5483e-08 1.747773584060822 2.5484e-08 1.8526366259306692 2.5485e-08 1.8265835490296845 2.5486e-08 1.8066092152932711 2.5487e-08 1.8655763863121546 2.5488e-08 1.8614825870103078 2.5489e-08 1.8185272273299962 2.549e-08 1.8067917516090881 2.5491e-08 1.8426473701648731 2.5492e-08 1.7521661050830661 2.5493e-08 1.7522456386611427 2.5494e-08 1.823145255876579 2.5495e-08 1.8715535779526673 2.5496e-08 1.7484867393385748 2.5497e-08 1.8140626511095133 2.5498e-08 1.8633184011319868 2.5499e-08 1.721224507030268 2.55e-08 1.795692709135949 2.5500999999999998e-08 1.8556243396602239 2.5502e-08 1.7766591733426482 2.5503e-08 1.7799636436833235 2.5503999999999998e-08 1.7364366686883066 2.5505e-08 1.7364637510902656 2.5506e-08 1.7591468984317626 2.5506999999999998e-08 1.7492677690434926 2.5508e-08 1.803511514477209 2.5509e-08 1.8676240310865306 2.5509999999999998e-08 1.7792772571085793 2.5511e-08 1.78398697590358 2.5512e-08 1.7362828349118586 2.5512999999999998e-08 1.8560054219570097 2.5514e-08 1.808430880710547 2.5515e-08 1.8208463870568161 2.5515999999999998e-08 1.7754105485051033 2.5517e-08 1.89889754906614 2.5518e-08 1.833217541721304 2.5519e-08 1.8485281078371376 2.552e-08 1.817783934324261 2.5521e-08 1.7650900846463566 2.5522e-08 1.7593045065532948 2.5523e-08 1.7807979874507418 2.5524e-08 1.748780186055389 2.5525e-08 1.8377804729664136 2.5526e-08 1.840204184218022 2.5527e-08 1.8434712963699005 2.5528e-08 1.820670285179498 2.5529e-08 1.8518819697252802 2.553e-08 1.8498258109917782 2.5531e-08 1.8289813201949154 2.5532e-08 1.7838331562256884 2.5533e-08 1.7539796090222166 2.5534e-08 1.7874198771375684 2.5535e-08 1.7350391351587358 2.5535999999999998e-08 1.7306116818236914 2.5537e-08 1.8018833995303387 2.5538e-08 1.7589870508719732 2.5538999999999998e-08 1.7721395131086035 2.554e-08 1.8004863966386995 2.5541e-08 1.8222407749535365 2.5541999999999998e-08 1.7612528964612688 2.5543e-08 1.777055808414453 2.5544e-08 1.7072463373591404 2.5544999999999998e-08 1.6925518693734878 2.5546e-08 1.8117287183929434 2.5547e-08 1.7505463287919114 2.5547999999999998e-08 1.838364432713371 2.5549e-08 1.7719896695784432 2.555e-08 1.800582617295903 2.5550999999999998e-08 1.8484671013414908 2.5552e-08 1.7883041332572331 2.5553e-08 1.7727113844542965 2.5554e-08 1.7673690741428945 2.5555e-08 1.7984587653169217 2.5556e-08 1.8674463098936585 2.5557e-08 1.7943516436684899 2.5558e-08 1.8206843488363416 2.5559e-08 1.7948576507459875 2.556e-08 1.8976222067571404 2.5561e-08 1.718176661801135 2.5562e-08 1.7318930297857593 2.5563e-08 1.790530372146253 2.5564e-08 1.8113502264002936 2.5565e-08 1.716345814239918 2.5566e-08 1.808375106849861 2.5567e-08 1.790378224185152 2.5568e-08 1.7969560900110755 2.5569e-08 1.786631782864663 2.557e-08 1.8559794892083605 2.5571e-08 1.8134390817535937 2.5572e-08 1.7523354170824939 2.5573e-08 1.898640057904882 2.5573999999999998e-08 1.7790004457355 2.5575e-08 1.7971996564350006 2.5576e-08 1.895565173332064 2.5576999999999998e-08 1.745385565582265 2.5578e-08 1.8335410590398904 2.5579e-08 1.8106845680824029 2.5579999999999998e-08 1.876951885136723 2.5581e-08 1.7925547478965127 2.5582e-08 1.8888893731418506 2.5582999999999998e-08 1.7641657128150177 2.5584e-08 1.8137651912759463 2.5585e-08 1.7231962615983383 2.5585999999999998e-08 1.7736225047066743 2.5587e-08 1.8001150988292431 2.5588e-08 1.7781844188724143 2.5589e-08 1.7720411740860738 2.559e-08 1.7376071623781337 2.5591e-08 1.8051894080203728 2.5592e-08 1.7829090667776082 2.5593e-08 1.8364893238265316 2.5594e-08 1.8331815246943903 2.5595e-08 1.751763855328304 2.5596e-08 1.781249276326957 2.5597e-08 1.7715258629518802 2.5598e-08 1.772623666959136 2.5599e-08 1.8531040090671007 2.56e-08 1.7828465964400673 2.5601e-08 1.8393968740713693 2.5602e-08 1.7740496532239185 2.5603e-08 1.8712783588474893 2.5604e-08 1.8422045982437627 2.5605e-08 1.766592151664341 2.5606e-08 1.7129212863896328 2.5607e-08 1.7894679876588828 2.5608e-08 1.7715854763100505 2.5608999999999998e-08 1.7968551676334967 2.561e-08 1.7491763284409105 2.5611e-08 1.7878770704682014 2.5611999999999998e-08 1.7634842037975558 2.5613e-08 1.8859332877467638 2.5614e-08 1.8269474293669967 2.5614999999999998e-08 1.797156806019779 2.5616e-08 1.8231050916074003 2.5617e-08 1.7613799188054073 2.5617999999999998e-08 1.7614688571741355 2.5619e-08 1.8239237936268253 2.562e-08 1.8067190168540364 2.5620999999999998e-08 1.768305431964218 2.5622e-08 1.847438838981069 2.5623e-08 1.805797233093997 2.5624e-08 1.7605220227251648 2.5625e-08 1.8477017186742277 2.5626e-08 1.7358495386615655 2.5627e-08 1.7913439933358857 2.5628e-08 1.8139794294432658 2.5629e-08 1.7911675448143891 2.563e-08 1.8438238873901498 2.5631e-08 1.8170772104312212 2.5632e-08 1.7057413078059502 2.5633e-08 1.8446933659947702 2.5634e-08 1.7427790077709544 2.5635e-08 1.770000217132712 2.5636e-08 1.7730731274696705 2.5637e-08 1.8638969471184696 2.5638e-08 1.8374863101267933 2.5639e-08 1.8180760385181134 2.564e-08 1.8102176589315808 2.5641e-08 1.774801444783157 2.5642e-08 1.876969680367426 2.5643e-08 1.7631899332424656 2.5643999999999998e-08 1.743915296415583 2.5645e-08 1.769101162394504 2.5646e-08 1.804462009670232 2.5646999999999998e-08 1.7993965074257672 2.5648e-08 1.6697083897558789 2.5649e-08 1.752981647682985 2.5649999999999998e-08 1.7656099641411045 2.5651e-08 1.7734987112400413 2.5652e-08 1.734134712272186 2.5652999999999998e-08 1.8553859055877384 2.5654e-08 1.8203223196256495 2.5655e-08 1.8026610918512191 2.5655999999999998e-08 1.8031794386775823 2.5657e-08 1.7761520777653996 2.5658e-08 1.82223336441926 2.5659e-08 1.8479589518932706 2.566e-08 1.7688927585619099 2.5661e-08 1.7315789911199628 2.5662e-08 1.825538832327888 2.5663e-08 1.7352695278010566 2.5664e-08 1.8121670364269 2.5665e-08 1.8194850149464201 2.5666e-08 1.8198439201832795 2.5667e-08 1.7219776573770391 2.5668e-08 1.846676810120698 2.5669e-08 1.7443002304408008 2.567e-08 1.780114750316637 2.5671e-08 1.794049300123242 2.5672e-08 1.8611946698758919 2.5673e-08 1.8606009584368184 2.5674e-08 1.8357668024672953 2.5675e-08 1.691402353511289 2.5676e-08 1.8790095482277573 2.5677e-08 1.7526774578161557 2.5678e-08 1.8561271317098955 2.5678999999999998e-08 1.7858466334217364 2.568e-08 1.7664871253877257 2.5681e-08 1.7597515501910073 2.5681999999999998e-08 1.823907747952603 2.5683e-08 1.8453248898195422 2.5684e-08 1.8477357680322088 2.5684999999999998e-08 1.7840213716029794 2.5686e-08 1.8877942227204092 2.5687e-08 1.8658805481426832 2.5687999999999998e-08 1.8261840991917826 2.5689e-08 1.7600017745953187 2.569e-08 1.800844741766234 2.5690999999999998e-08 1.7752240021001973 2.5692e-08 1.716161742768012 2.5693e-08 1.7072249750871147 2.5693999999999998e-08 1.786301297176218 2.5695e-08 1.7667772756276054 2.5696e-08 1.8210900792387976 2.5697e-08 1.8663577496270989 2.5698e-08 1.7931928984218974 2.5699e-08 1.8397494131998249 2.57e-08 1.8186694447414562 2.5701e-08 1.7546279875616826 2.5702e-08 1.7448408284133043 2.5703e-08 1.7478106790899783 2.5704e-08 1.8093940795504688 2.5705e-08 1.711290899762869 2.5706e-08 1.7648542793903843 2.5707e-08 1.909996259342587 2.5708e-08 1.8813696471183865 2.5709e-08 1.8173298575877737 2.571e-08 1.7639480965749992 2.5711e-08 1.8003222044469898 2.5712e-08 1.807351989163722 2.5713e-08 1.7736758617382558 2.5713999999999998e-08 1.7846343291956304 2.5715e-08 1.8215306869958758 2.5716e-08 1.7813429381867134 2.5716999999999998e-08 1.8858945668021232 2.5718e-08 1.7377025738235299 2.5719e-08 1.7745391287322951 2.5719999999999998e-08 1.8574125953362841 2.5721e-08 1.8198482614583473 2.5722e-08 1.791725032920747 2.5722999999999998e-08 1.7300619222939708 2.5724e-08 1.79490900139245 2.5725e-08 1.8259571628062214 2.5725999999999998e-08 1.8040592827064958 2.5727e-08 1.7735575674607449 2.5728e-08 1.8053583753661626 2.5728999999999998e-08 1.8450738134235254 2.573e-08 1.8237299617976412 2.5731e-08 1.8392966260480397 2.5732e-08 1.878117306478258 2.5733e-08 1.8266111801756806 2.5734e-08 1.838283504037685 2.5735e-08 1.7346224878375853 2.5736e-08 1.7234122978064277 2.5737e-08 1.8109931127006371 2.5738e-08 1.7397227177099617 2.5739e-08 1.7330009478250044 2.574e-08 1.8753078800756957 2.5741e-08 1.76341219971085 2.5742e-08 1.7689167911711696 2.5743e-08 1.9408988579467104 2.5744e-08 1.7644290894572772 2.5745e-08 1.7861456028142766 2.5746e-08 1.8022840291507252 2.5747e-08 1.8512563077444602 2.5748e-08 1.8376574265530554 2.5748999999999998e-08 1.8096768136037211 2.575e-08 1.7808004572391238 2.5751e-08 1.8190367441567037 2.5751999999999998e-08 1.8503429682625783 2.5753e-08 1.761187407324676 2.5754e-08 1.8202548420087117 2.5754999999999998e-08 1.7267392419066467 2.5756e-08 1.8285016285229376 2.5757e-08 1.6912593693911844 2.5757999999999998e-08 1.853099862881027 2.5759e-08 1.7448763349153602 2.576e-08 1.7385814558933728 2.5760999999999998e-08 1.7871298695548725 2.5762e-08 1.836801957301488 2.5763e-08 1.7635248162667818 2.5763999999999998e-08 1.722528587208441 2.5765e-08 1.8537090237258949 2.5766e-08 1.7420467511153088 2.5767e-08 1.8016021368895725 2.5768e-08 1.8232137264514794 2.5769e-08 1.7887529579631771 2.577e-08 1.8490364903982677 2.5771e-08 1.895842888595596 2.5772e-08 1.8288572064091995 2.5773e-08 1.7675137140261508 2.5774e-08 1.9134527372157144 2.5775e-08 1.6872669693011222 2.5776e-08 1.7883878007251643 2.5777e-08 1.7873818388751912 2.5778e-08 1.7247177597661705 2.5779e-08 1.812123966170007 2.578e-08 1.8277825773481284 2.5781e-08 1.779560982404954 2.5782e-08 1.813025210987295 2.5783e-08 1.7662159462769684 2.5784e-08 1.813802582169285 2.5785e-08 1.932831792992064 2.5786e-08 1.804920902550864 2.5786999999999998e-08 1.8383976901067554 2.5788e-08 1.8520296111852366 2.5789e-08 1.7613761208027934 2.5789999999999998e-08 1.751972799451435 2.5791e-08 1.740393222383642 2.5792e-08 1.8118358354396291 2.5792999999999998e-08 1.7567493975237576 2.5794e-08 1.8791938996116966 2.5795e-08 1.7779836307509804 2.5795999999999998e-08 1.778817979469066 2.5797e-08 1.6637810961542885 2.5798e-08 1.872768891114249 2.5798999999999998e-08 1.8861989405958453 2.58e-08 1.7304591836383452 2.5801e-08 1.8186526058988306 2.5802e-08 1.8360944007526232 2.5803e-08 1.931598989143268 2.5804e-08 1.8280621566246362 2.5805e-08 1.832222971258196 2.5806e-08 1.7781133495511434 2.5807e-08 1.7991153415301195 2.5808e-08 1.779299883093872 2.5809e-08 1.7925461322145202 2.581e-08 1.9323268752040137 2.5811e-08 1.749552009458513 2.5812e-08 1.6645323679890458 2.5813e-08 1.8032728845605204 2.5814e-08 1.83902394642901 2.5815e-08 1.8955310910519838 2.5816e-08 1.7788228766364875 2.5817e-08 1.8247683060337045 2.5818e-08 1.7583154682228628 2.5819e-08 1.7609683143263144 2.582e-08 1.7875804752014135 2.5821e-08 1.8263217366075404 2.5821999999999998e-08 1.7890354456089357 2.5823e-08 1.7884549679828616 2.5824e-08 1.7568039913141023 2.5824999999999998e-08 1.7918102754812675 2.5826e-08 1.7691886239191636 2.5827e-08 1.824871309889172 2.5827999999999998e-08 1.7262451559136436 2.5829e-08 1.8650670786668173 2.583e-08 1.8264396625009873 2.5830999999999998e-08 1.844408036595227 2.5832e-08 1.805894577425731 2.5833e-08 1.8047629195546155 2.5833999999999998e-08 1.858087521734738 2.5835e-08 1.7568131166127579 2.5836e-08 1.7520831964042063 2.5837e-08 1.7784935902015853 2.5838e-08 1.825608683298774 2.5839e-08 1.7801102527695418 2.584e-08 1.8011757586058044 2.5841e-08 1.850555718166704 2.5842e-08 1.7786786623219795 2.5843e-08 1.9710202802427428 2.5844e-08 1.8392302359937982 2.5845e-08 1.8363355108165427 2.5846e-08 1.8128569858632277 2.5847e-08 1.78225473345166 2.5848e-08 1.7157695172163911 2.5849e-08 1.873587411403817 2.585e-08 1.8498571731312707 2.5851e-08 1.8030582418881718 2.5852e-08 1.8873676734445917 2.5853e-08 1.7817356267444049 2.5854e-08 1.8380365261880995 2.5855e-08 1.7099777424840725 2.5856e-08 1.8292179907893273 2.5856999999999998e-08 1.8515917446934589 2.5858e-08 1.7803346369467807 2.5859e-08 1.796468389710202 2.5859999999999998e-08 1.9233959576643134 2.5861e-08 1.7656882135621452 2.5862e-08 1.8266575487855798 2.5862999999999998e-08 1.7786407424477813 2.5864e-08 1.8358594095600513 2.5865e-08 1.7524132958789904 2.5865999999999998e-08 1.7787665779041528 2.5867e-08 1.8500743189049997 2.5868e-08 1.8010130135875546 2.5868999999999998e-08 1.8752228325451032 2.587e-08 1.766221254580942 2.5871e-08 1.7135873899634582 2.5871999999999998e-08 1.8323283008009008 2.5873e-08 1.821225283625587 2.5874e-08 1.728761845805441 2.5875e-08 1.768708555707133 2.5876e-08 1.793322571024982 2.5877e-08 1.8550814994350553 2.5878e-08 1.7484376683739462 2.5879e-08 1.772915762963391 2.588e-08 1.8726489592274074 2.5881e-08 1.7679723906203406 2.5882e-08 1.8222024709501194 2.5883e-08 1.8100080567969532 2.5884e-08 1.758926751118758 2.5885e-08 1.8896409592162524 2.5886e-08 1.8140561610086028 2.5887e-08 1.87752841715515 2.5888e-08 1.8688345460818114 2.5889e-08 1.7995064645781536 2.589e-08 1.8392973395653966 2.5891e-08 1.8578934102220057 2.5891999999999998e-08 1.8049834553008506 2.5893e-08 1.7297792580592097 2.5894e-08 1.8098657159486107 2.5894999999999998e-08 1.7980772522497042 2.5896e-08 1.8798173951841235 2.5897e-08 1.7154932794662112 2.5897999999999998e-08 1.8074455653803678 2.5899e-08 1.7853393898782122 2.59e-08 1.7872623175431237 2.5900999999999998e-08 1.763383793450591 2.5902e-08 1.8757321334242052 2.5903e-08 1.769505888516027 2.5903999999999998e-08 1.8010787072804024 2.5905e-08 1.7373129736176738 2.5906e-08 1.7431249037389531 2.5906999999999998e-08 1.8176011027798376 2.5908e-08 1.9064662455069183 2.5909e-08 1.8445187093114725 2.591e-08 1.8259962661330889 2.5911e-08 1.7934666094213474 2.5912e-08 1.8292093224222474 2.5913e-08 1.8519606503242951 2.5914e-08 1.9040726562310604 2.5915e-08 1.72838856913975 2.5916e-08 1.7455368420694963 2.5917e-08 1.8516139591641885 2.5918e-08 1.8602123818967198 2.5919e-08 1.7896256745258687 2.592e-08 1.7956967388138567 2.5921e-08 1.7109913881946963 2.5922e-08 1.7632586506847463 2.5923e-08 1.8303834372913905 2.5924e-08 1.8049695576805251 2.5925e-08 1.815399843682723 2.5926e-08 1.7243453136879465 2.5926999999999998e-08 1.7909823211980158 2.5928e-08 1.784763474671748 2.5929e-08 1.6757027873686496 2.5929999999999998e-08 1.6711320849384033 2.5931e-08 1.7718684389509336 2.5932e-08 1.7851991799783213 2.5932999999999998e-08 1.7694698034688874 2.5934e-08 1.863102834173363 2.5935e-08 1.8197345463139931 2.5935999999999998e-08 1.7422906209012745 2.5937e-08 1.8128090201738924 2.5938e-08 1.794958357942173 2.5938999999999998e-08 1.8215803321153514 2.594e-08 1.8291246067554938 2.5941e-08 1.752050107483383 2.5941999999999998e-08 1.6813596310641954 2.5943e-08 1.8124775771832569 2.5944e-08 1.758823430711075 2.5945e-08 1.8124694266853165 2.5946e-08 1.8934430294256523 2.5947e-08 1.7749137341535883 2.5948e-08 1.7542195443552688 2.5949e-08 1.822626567987582 2.595e-08 1.8327486299795277 2.5951e-08 1.788599414235811 2.5952e-08 1.8417443673784384 2.5953e-08 1.658273745074433 2.5954e-08 1.8092313209405637 2.5955e-08 1.8366429426883828 2.5956e-08 1.8762207474525439 2.5957e-08 1.834517156325465 2.5958e-08 1.7061778308879432 2.5959e-08 1.7825091816739491 2.596e-08 1.7530686397490975 2.5961e-08 1.8607742571979045 2.5962e-08 1.800127387563025 2.5963e-08 1.750027824208505 2.5964e-08 1.7859154462624218 2.5964999999999998e-08 1.8951747865514195 2.5966e-08 1.792057396932254 2.5967e-08 1.8249303666013839 2.5967999999999998e-08 1.7285508982037567 2.5969e-08 1.8143289990154887 2.597e-08 1.8350501731596967 2.5970999999999998e-08 1.8599448909523113 2.5972e-08 1.7720552426527598 2.5973e-08 1.7433887654828033 2.5973999999999998e-08 1.8006529176834123 2.5975e-08 1.8281915776169009 2.5976e-08 1.8482486514392384 2.5976999999999998e-08 1.7543671835004337 2.5978e-08 1.792713137403124 2.5979e-08 1.7460416680883801 2.598e-08 1.8259115691955847 2.5981e-08 1.785870790404572 2.5982e-08 1.8420612067087765 2.5983e-08 1.8263155581171386 2.5984e-08 1.8315731775589483 2.5985e-08 1.771056999051612 2.5986e-08 1.8267747870258906 2.5987e-08 1.7683244552100952 2.5988e-08 1.7462521353359566 2.5989e-08 1.7881004345838543 2.599e-08 1.877820190498948 2.5991e-08 1.8509396575027035 2.5992e-08 1.7674020244329125 2.5993e-08 1.7853896680338346 2.5994e-08 1.7358367882131582 2.5995e-08 1.770728715470881 2.5996e-08 1.864068540715145 2.5997e-08 1.7773987922678702 2.5998e-08 1.813879159780172 2.5999e-08 1.7612782273495358 2.5999999999999998e-08 1.798321061040184 2.6001e-08 1.695739690058539 2.6002e-08 1.800315843092146 2.6002999999999998e-08 1.7829120680252202 2.6004e-08 1.814671403073797 2.6005e-08 1.8481975916896625 2.6005999999999998e-08 1.8666183300149801 2.6007e-08 1.890959479859216 2.6008e-08 1.7824406878844354 2.6008999999999998e-08 1.769664291974606 2.601e-08 1.8011533833695825 2.6011e-08 1.7453038522603297 2.6011999999999998e-08 1.8290145982812789 2.6013e-08 1.7179839292925212 2.6014e-08 1.8334447776580467 2.6015e-08 1.7758799374507672 2.6016e-08 1.7967569936030088 2.6017e-08 1.7706732239070986 2.6018e-08 1.7396749425495466 2.6019e-08 1.7509228598186508 2.602e-08 1.8141880439180025 2.6021e-08 1.8290891959171192 2.6022e-08 1.827908642920324 2.6023e-08 1.7898004443618127 2.6024e-08 1.8114584803212515 2.6025e-08 1.745800410444093 2.6026e-08 1.781124437877419 2.6027e-08 1.7736992673265342 2.6028e-08 1.797018810806224 2.6029e-08 1.7326551332253521 2.603e-08 1.7895834227857093 2.6031e-08 1.8404771231967314 2.6032e-08 1.7738705795222591 2.6033e-08 1.7758494307126231 2.6034e-08 1.747318944857644 2.6034999999999998e-08 1.815213605846273 2.6036e-08 1.7807586364155468 2.6037e-08 1.750826476769511 2.6037999999999998e-08 1.805404509103038 2.6039e-08 1.860140839582103 2.604e-08 1.78343359073857 2.6040999999999998e-08 1.7978489677378233 2.6042e-08 1.8936354111665064 2.6043e-08 1.7887863072721557 2.6043999999999998e-08 1.7968864787435823 2.6045e-08 1.7565747438615167 2.6046e-08 1.7967288416979739 2.6046999999999998e-08 1.800454389779118 2.6048e-08 1.7577685499175248 2.6049e-08 1.7944050078624398 2.6049999999999998e-08 1.7079735072228184 2.6051e-08 1.7572642632949036 2.6052e-08 1.790389911063216 2.6053e-08 1.8652031502235515 2.6054e-08 1.7551450070919674 2.6055e-08 1.761356246438991 2.6056e-08 1.7541559691926103 2.6057e-08 1.814350086995711 2.6058e-08 1.8517954761500377 2.6059e-08 1.9151084461973067 2.606e-08 1.840717313392268 2.6061e-08 1.8063075180067825 2.6062e-08 1.759123068849649 2.6063e-08 1.8313437448289047 2.6064e-08 1.8076718569953911 2.6065e-08 1.8345829238333684 2.6066e-08 1.8718847585136795 2.6067e-08 1.8219264876689996 2.6068e-08 1.8440751214368838 2.6069e-08 1.8472329485672925 2.6069999999999998e-08 1.8239631483898446 2.6071e-08 1.9313453773500289 2.6072e-08 1.9047790120236539 2.6072999999999998e-08 1.7225801255185016 2.6074e-08 1.891642483222098 2.6075e-08 1.7675963615787833 2.6075999999999998e-08 1.8325670944934274 2.6077e-08 1.8515062456908307 2.6078e-08 1.7546501254011577 2.6078999999999998e-08 1.7730323313010612 2.608e-08 1.7645503790533716 2.6081e-08 1.7745901554282586 2.6081999999999998e-08 1.8636969308626845 2.6083e-08 1.8111742931920105 2.6084e-08 1.8363184712089027 2.6084999999999998e-08 1.8585549990947414 2.6086e-08 1.786601584440052 2.6087e-08 1.8092054286103925 2.6088e-08 1.8085203768859057 2.6089e-08 1.893134623847514 2.609e-08 1.7352587759946758 2.6091e-08 1.8496675644897793 2.6092e-08 1.849954609051488 2.6093e-08 1.789302324227996 2.6094e-08 1.8266119072555287 2.6095e-08 1.7621219557806842 2.6096e-08 1.6882283967311853 2.6097e-08 1.838950220485217 2.6098e-08 1.7831903071545296 2.6099e-08 1.8166427425784089 2.61e-08 1.8847525517261023 2.6101e-08 1.7617778031904663 2.6102e-08 1.8687649953336363 2.6103e-08 1.825165362939868 2.6104e-08 1.747317856209354 2.6104999999999998e-08 1.7565130706834677 2.6106e-08 1.731702232858377 2.6107e-08 1.7879795520651152 2.6107999999999998e-08 1.7488588554648195 2.6109e-08 1.6749652069911323 2.611e-08 1.8379862385636103 2.6110999999999998e-08 1.7744243900659487 2.6112e-08 1.8845677470813975 2.6113e-08 1.7809861105973972 2.6113999999999998e-08 1.7181904080580184 2.6115e-08 1.8082126765886823 2.6116e-08 1.863255967193825 2.6116999999999998e-08 1.814791930720928 2.6118e-08 1.75053647852555 2.6119e-08 1.791660191737359 2.6119999999999998e-08 1.8863221726450377 2.6121e-08 1.805473258174592 2.6122e-08 1.8294375772002924 2.6123e-08 1.815128585464487 2.6124e-08 1.8011858681897561 2.6125e-08 1.8086445641706175 2.6126e-08 1.8083984407639593 2.6127e-08 1.8182856107846632 2.6128e-08 1.7981383996809162 2.6129e-08 1.8163781669747576 2.613e-08 1.8064754128519867 2.6131e-08 1.7982719599088808 2.6132e-08 1.7474797664291073 2.6133e-08 1.8326307245794091 2.6134e-08 1.722230447408871 2.6135e-08 1.8107656253782194 2.6136e-08 1.8070471407847868 2.6137e-08 1.8639064920912711 2.6138e-08 1.8526123542595025 2.6139e-08 1.8381128286846997 2.6139999999999998e-08 1.859529290316726 2.6141e-08 1.8186325771108778 2.6142e-08 1.6975562616784503 2.6142999999999998e-08 1.7988892179013138 2.6144e-08 1.7705834400449239 2.6145e-08 1.7532978101696213 2.6145999999999998e-08 1.815946144964243 2.6147e-08 1.7817376405325072 2.6148e-08 1.7705796731575043 2.6148999999999998e-08 1.7098353586184172 2.615e-08 1.8252835876443203 2.6151e-08 1.727956953101033 2.6151999999999998e-08 1.8566524614090292 2.6153e-08 1.8008560491491281 2.6154e-08 1.8535729224674664 2.6154999999999998e-08 1.7911938920841723 2.6156e-08 1.8352436040836013 2.6157e-08 1.8218774186856372 2.6158e-08 1.7867493246437263 2.6159e-08 1.7246210123145334 2.616e-08 1.7801696365562052 2.6161e-08 1.7603755983497757 2.6162e-08 1.75315160194914 2.6163e-08 1.7889421483038561 2.6164e-08 1.749844210601688 2.6165e-08 1.7420895784466663 2.6166e-08 1.8409377922772976 2.6167e-08 1.8343429319375486 2.6168e-08 1.8031231432360728 2.6169e-08 1.7907335728113334 2.617e-08 1.8844578537438363 2.6171e-08 1.8222884502607188 2.6172e-08 1.7982477574000255 2.6173e-08 1.829615332621113 2.6174e-08 1.7551252914548223 2.6175e-08 1.8204072064638155 2.6176e-08 1.781850605690182 2.6177e-08 1.805633864512371 2.6177999999999998e-08 1.7873811736386918 2.6179e-08 1.8048521430044937 2.618e-08 1.7970710765406825 2.6180999999999998e-08 1.8406461039983517 2.6182e-08 1.9104450592515796 2.6183e-08 1.8462887225660096 2.6183999999999998e-08 1.785394349711693 2.6185e-08 1.8301114094337816 2.6186e-08 1.804991750444288 2.6186999999999998e-08 1.812008382768482 2.6188e-08 1.8137628935170513 2.6189e-08 1.7527825171145224 2.6189999999999998e-08 1.714608654667591 2.6191e-08 1.755469767963441 2.6192e-08 1.8353558340683813 2.6193e-08 1.7934229721157289 2.6194e-08 1.7588632245451952 2.6195e-08 1.898559791947066 2.6196e-08 1.7998704384485515 2.6197e-08 1.819325951601361 2.6198e-08 1.757116311407598 2.6199e-08 1.8264999100561146 2.62e-08 1.8310911540805574 2.6201e-08 1.8159727480047336 2.6202e-08 1.7991764368746639 2.6203e-08 1.852617502490235 2.6204e-08 1.787768829134984 2.6205e-08 1.8183765125927305 2.6206e-08 1.7863477269641925 2.6207e-08 1.72505708909496 2.6208e-08 1.8206915837874953 2.6209e-08 1.8217736058166407 2.621e-08 1.8235184734729164 2.6211e-08 1.8024643330798678 2.6212e-08 1.8013674574129694 2.6212999999999998e-08 1.862804138355085 2.6214e-08 1.830342278814558 2.6215e-08 1.8434873856503202 2.6215999999999998e-08 1.771838558192882 2.6217e-08 1.8480193687865245 2.6218e-08 1.7675134998674438 2.6218999999999998e-08 1.7427549465289085 2.622e-08 1.8375090039869428 2.6221e-08 1.7745657355121625 2.6221999999999998e-08 1.7295377898592432 2.6223e-08 1.75888311742689 2.6224e-08 1.8603195738419662 2.6224999999999998e-08 1.7787434850454735 2.6226e-08 1.7488302918725285 2.6227e-08 1.8238796766523349 2.6228e-08 1.7888035923649113 2.6229e-08 1.758242522606517 2.623e-08 1.9366873145801045 2.6231e-08 1.8722094946558543 2.6232e-08 1.752859710438676 2.6233e-08 1.8550519223631716 2.6234e-08 1.7975374340189831 2.6235e-08 1.6370171134500673 2.6236e-08 1.7704918544542871 2.6237e-08 1.7384111165935092 2.6238e-08 1.798478673586239 2.6239e-08 1.752496957799421 2.624e-08 1.7929012340304458 2.6241e-08 1.7822658546036052 2.6242e-08 1.833960598253423 2.6243e-08 1.828414827431751 2.6244e-08 1.7670525286204457 2.6245e-08 1.774558195822271 2.6246e-08 1.848453605389851 2.6247e-08 1.7979702602186838 2.6247999999999998e-08 1.762716500790405 2.6249e-08 1.7895250097142077 2.625e-08 1.787067816812604 2.6250999999999998e-08 1.798729364056325 2.6252e-08 1.7447439419710988 2.6253e-08 1.830318856201473 2.6253999999999998e-08 1.8481713182896533 2.6255e-08 1.8289839928140972 2.6256e-08 1.8084264141402466 2.6256999999999998e-08 1.7214641889579911 2.6258e-08 1.8685979787626688 2.6259e-08 1.8365964588944321 2.6259999999999998e-08 1.8731551557483745 2.6261e-08 1.7095036240162549 2.6262e-08 1.786521295596192 2.6262999999999998e-08 1.8108323695251953 2.6264e-08 1.880323993969318 2.6265e-08 1.7615208448708106 2.6266e-08 1.8428055690461578 2.6267e-08 1.7353419644045358 2.6268e-08 1.7509529021494519 2.6269e-08 1.818734684986468 2.627e-08 1.8466270376961675 2.6271e-08 1.8382166730920457 2.6272e-08 1.795812977894432 2.6273e-08 1.72512173252454 2.6274e-08 1.833081290087736 2.6275e-08 1.813554278512952 2.6276e-08 1.787480589532751 2.6277e-08 1.7503872555553273 2.6278e-08 1.7507686586653068 2.6279e-08 1.845867884670524 2.628e-08 1.7755401620197078 2.6281e-08 1.8290406609307792 2.6282e-08 1.7643081829400598 2.6282999999999998e-08 1.7656694515902425 2.6284e-08 1.7353655125125023 2.6285e-08 1.7797067232272046 2.6285999999999998e-08 1.8007015800217634 2.6287e-08 1.7574155218784682 2.6288e-08 1.7926812130686558 2.6288999999999998e-08 1.7075910244184833 2.629e-08 1.8623273775765563 2.6291e-08 1.6627483654465414 2.6291999999999998e-08 1.818425703236351 2.6293e-08 1.7109901923278146 2.6294e-08 1.770313161893197 2.6294999999999998e-08 1.836120449386924 2.6296e-08 1.7476024380772952 2.6297e-08 1.8270262377444682 2.6297999999999998e-08 1.8609414607697052 2.6299e-08 1.88194426593524 2.63e-08 1.7234877590410593 2.6301e-08 1.7423084509469502 2.6302e-08 1.844837971929942 2.6303e-08 1.7993766646041995 2.6304e-08 1.8110850077748983 2.6305e-08 1.8552322768160332 2.6306e-08 1.7988228954414902 2.6307e-08 1.7232076213614957 2.6308e-08 1.7350423638175978 2.6309e-08 1.797087480652753 2.631e-08 1.7823494141621654 2.6311e-08 1.8762544798495766 2.6312e-08 1.8564813773958977 2.6313e-08 1.7832096992266022 2.6314e-08 1.8409259893637424 2.6315e-08 1.8984499614368113 2.6316e-08 1.8492470767943159 2.6317e-08 1.7777505776633131 2.6317999999999998e-08 1.751973755038046 2.6319e-08 1.7976052813995602 2.632e-08 1.7158765896594552 2.6320999999999998e-08 1.7696675935303372 2.6322e-08 1.8361381264394983 2.6323e-08 1.8189353231261847 2.6323999999999998e-08 1.8321806828808647 2.6325e-08 1.7467218490920138 2.6326e-08 1.7419301532067932 2.6326999999999998e-08 1.8102027036172208 2.6328e-08 1.8345532958155102 2.6329e-08 1.7803596972823574 2.6329999999999998e-08 1.7873175929681624 2.6331e-08 1.7957647455092431 2.6332e-08 1.869882035131179 2.6332999999999998e-08 1.8420594797852778 2.6334e-08 1.7763840519844787 2.6335e-08 1.7627685241027418 2.6336e-08 1.883665744927328 2.6337e-08 1.8625869414412304 2.6338e-08 1.8306966242658842 2.6339e-08 1.7538862399277013 2.634e-08 1.8686433063972177 2.6341e-08 1.8285190272850442 2.6342e-08 1.841445553646353 2.6343e-08 1.7715225432190749 2.6344e-08 1.834880397713033 2.6345e-08 1.838051204178695 2.6346e-08 1.7247098138718364 2.6347e-08 1.82120631944346 2.6348e-08 1.78931166858863 2.6349e-08 1.8539261982761286 2.635e-08 1.7476629620965543 2.6351e-08 1.7780265427038318 2.6352e-08 1.8698125439131597 2.6353e-08 1.7094293194961367 2.6354e-08 1.7777847338577402 2.6355e-08 1.7234724856869872 2.6355999999999998e-08 1.7096484595062214 2.6357e-08 1.918988979809477 2.6358e-08 1.8387732716443026 2.6358999999999998e-08 1.8081153678499746 2.636e-08 1.8520827463713425 2.6361e-08 1.7853552377452073 2.6361999999999998e-08 1.8690992763834477 2.6363e-08 1.767898449229864 2.6364e-08 1.788767234647307 2.6364999999999998e-08 1.8057149895627114 2.6366e-08 1.7886086731422906 2.6367e-08 1.8512844350954671 2.6367999999999998e-08 1.7998627705898744 2.6369e-08 1.7419578109360685 2.637e-08 1.8506198174622153 2.6371e-08 1.8384706079884245 2.6372e-08 1.7391221588389723 2.6373e-08 1.9215730232709356 2.6374e-08 1.8378783293969614 2.6375e-08 1.8569627802083608 2.6376e-08 1.8242685835315122 2.6377e-08 1.830791234847833 2.6378e-08 1.8426719745005877 2.6379e-08 1.9096902981221286 2.638e-08 1.813886280432354 2.6381e-08 1.7925844048932358 2.6382e-08 1.7865844613955841 2.6383e-08 1.7381863587464021 2.6384e-08 1.7802449069728494 2.6385e-08 1.7714903178210308 2.6386e-08 1.9111162320968715 2.6387e-08 1.9031140434719929 2.6388e-08 1.862859333053116 2.6389e-08 1.7908392391908143 2.639e-08 1.7445863149175391 2.6390999999999998e-08 1.7488618694017795 2.6392e-08 1.763701991029895 2.6393e-08 1.7552803286635874 2.6393999999999998e-08 1.801397152171509 2.6395e-08 1.7787023232180048 2.6396e-08 1.8619964396959032 2.6396999999999998e-08 1.8058061620566668 2.6398e-08 1.833729249111811 2.6399e-08 1.7736145237344223 2.6399999999999998e-08 1.799169866305791 2.6401e-08 1.8375322043955788 2.6402e-08 1.788916918284709 2.6402999999999998e-08 1.8872027723387323 2.6404e-08 1.785165424199555 2.6405e-08 1.7473160843796407 2.6406e-08 1.7470594755358864 2.6407e-08 1.8643778347891473 2.6408e-08 1.8536667253776147 2.6409e-08 1.8118196077712856 2.641e-08 1.830953128947761 2.6411e-08 1.820673856097821 2.6412e-08 1.8205845238086749 2.6413e-08 1.7082589033621336 2.6414e-08 1.7537024210729797 2.6415e-08 1.7756844395633193 2.6416e-08 1.8449439703757662 2.6417e-08 1.7052690079700046 2.6418e-08 1.76111611149625 2.6419e-08 1.7724702873204707 2.642e-08 1.73206646056654 2.6421e-08 1.8117292738525912 2.6422e-08 1.7747433455231345 2.6423e-08 1.8298996653044286 2.6424e-08 1.8277817347613436 2.6425e-08 1.796318987400748 2.6425999999999998e-08 1.7967286610761641 2.6427e-08 1.811841875033107 2.6428e-08 1.7684544745290394 2.6428999999999998e-08 1.864864095310525 2.643e-08 1.78489531034587 2.6431e-08 1.7891312484838873 2.6431999999999998e-08 1.8264590635291316 2.6433e-08 1.7604031979125445 2.6434e-08 1.8273790187877157 2.6434999999999998e-08 1.688456631475526 2.6436e-08 1.8371692078822197 2.6437e-08 1.767804909142285 2.6437999999999998e-08 1.7580661359132435 2.6439e-08 1.7979182845397053 2.644e-08 1.7827304281968255 2.6440999999999998e-08 1.794681636674437 2.6442e-08 1.7911199497621875 2.6443e-08 1.812040389792681 2.6444e-08 1.8017982879289207 2.6445e-08 1.7742154988389511 2.6446e-08 1.7689503685451837 2.6447e-08 1.8530642125706032 2.6448e-08 1.8121646504151339 2.6449e-08 1.8408994699599104 2.645e-08 1.8854507917134125 2.6451e-08 1.7407188238721625 2.6452e-08 1.818831089595523 2.6453e-08 1.7451409053786244 2.6454e-08 1.7906848734890517 2.6455e-08 1.8005977718167836 2.6456e-08 1.792199643988445 2.6457e-08 1.796399516807804 2.6458e-08 1.8842855826014189 2.6459e-08 1.7383187976494505 2.646e-08 1.7533963719909045 2.6460999999999998e-08 1.8902238850473485 2.6462e-08 1.7614999416996628 2.6463e-08 1.7490989492434221 2.6463999999999998e-08 1.856252721964168 2.6465e-08 1.7048712694742814 2.6466e-08 1.7416660951087972 2.6466999999999998e-08 1.7051156703374755 2.6468e-08 1.8404096933636382 2.6469e-08 1.7923077641513598 2.6469999999999998e-08 1.8999436845552689 2.6471e-08 1.7432478814071974 2.6472e-08 1.772644328387081 2.6472999999999998e-08 1.8104952277729358 2.6474e-08 1.8294037859831214 2.6475e-08 1.8168382926283855 2.6475999999999998e-08 1.724849063137224 2.6477e-08 1.7513173888855158 2.6478e-08 1.7750196945459213 2.6479e-08 1.7319271669667602 2.648e-08 1.7675012081937183 2.6481e-08 1.731459680498275 2.6482e-08 1.8082614307973588 2.6483e-08 1.7757952630038274 2.6484e-08 1.7482559392942374 2.6485e-08 1.8275974709470038 2.6486e-08 1.7157112169177395 2.6487e-08 1.759204966543911 2.6488e-08 1.8012384738790175 2.6489e-08 1.7514812240655255 2.649e-08 1.7760329577177985 2.6491e-08 1.8648902285233098 2.6492e-08 1.8067595335897286 2.6493e-08 1.7704681637060538 2.6494e-08 1.6913463435942162 2.6495e-08 1.9092824287772596 2.6495999999999998e-08 1.8571716701344003 2.6497e-08 1.9454249984028558 2.6498e-08 1.7586756638931011 2.6498999999999998e-08 1.7774448786988746 2.65e-08 1.9613484129807717 2.6501e-08 1.7587315719494467 2.6501999999999998e-08 1.790944808164943 2.6503e-08 1.805963497166555 2.6504e-08 1.693321681881565 2.6504999999999998e-08 1.8732226002306127 2.6506e-08 1.809572864727025 2.6507e-08 1.7712130805949045 2.6507999999999998e-08 1.824608215491474 2.6509e-08 1.821803496563621 2.651e-08 1.8138450543443685 2.6510999999999998e-08 1.8273693994318005 2.6512e-08 1.8190980454246006 2.6513e-08 1.7259886288542614 2.6514e-08 1.744912454320151 2.6515e-08 1.829712170708536 2.6516e-08 1.7616126360651267 2.6517e-08 1.7831068318823593 2.6518e-08 1.794738368487476 2.6519e-08 1.7904378507149263 2.652e-08 1.77064287374564 2.6521e-08 1.7969713876354398 2.6522e-08 1.885748779383987 2.6523e-08 1.8103865986020682 2.6524e-08 1.7483848049757058 2.6525e-08 1.6821541437757037 2.6526e-08 1.760471013808542 2.6527e-08 1.72279575842137 2.6528e-08 1.7110909667622796 2.6529e-08 1.8227246887283595 2.653e-08 1.7404821833853208 2.6530999999999998e-08 1.8897504706840584 2.6532e-08 1.72245354481519 2.6533e-08 1.7493170358132626 2.6533999999999998e-08 1.8674156257954562 2.6535e-08 1.8055932771039946 2.6536e-08 1.8146643802719973 2.6536999999999998e-08 1.7373152157034304 2.6538e-08 1.809331863437931 2.6539e-08 1.7562588370792929 2.6539999999999998e-08 1.8428398772243306 2.6541e-08 1.8320299825588497 2.6542e-08 1.7358934578836938 2.6542999999999998e-08 1.7707458881896796 2.6544e-08 1.7379329261264658 2.6545e-08 1.8167720223938448 2.6545999999999998e-08 1.7165400135175495 2.6547e-08 1.7598420873235292 2.6548e-08 1.8368771003117883 2.6549e-08 1.8229835121416713 2.655e-08 1.7722570959967678 2.6551e-08 1.7880256313751335 2.6552e-08 1.787405313577835 2.6553e-08 1.7885399699253273 2.6554e-08 1.878399823100041 2.6555e-08 1.7297611195729243 2.6556e-08 1.7916124731509113 2.6557e-08 1.8273711748724564 2.6558e-08 1.7778401108828297 2.6559e-08 1.8076054410451137 2.656e-08 1.803083126103276 2.6561e-08 1.7761268277798852 2.6562e-08 1.8633162111491228 2.6563e-08 1.8456856949323879 2.6564e-08 1.772544429069581 2.6565e-08 1.8287497443804734 2.6566e-08 1.71415073390758 2.6567e-08 1.8639799310048812 2.6568e-08 1.8025599552484273 2.6568999999999998e-08 1.835970945339549 2.657e-08 1.7901755669465207 2.6571e-08 1.8295331399502106 2.6571999999999998e-08 1.7959569563276727 2.6573e-08 1.7691887927441552 2.6574e-08 1.83603803834015 2.6574999999999998e-08 1.7357027115298849 2.6576e-08 1.845132664829558 2.6577e-08 1.7999157450569467 2.6577999999999998e-08 1.7613816362246304 2.6579e-08 1.7396024245904484 2.658e-08 1.8297918874551031 2.6580999999999998e-08 1.8098219037634051 2.6582e-08 1.7617600845144916 2.6583e-08 1.8577102857429169 2.6584e-08 1.7307873322423855 2.6585e-08 1.8084185399533783 2.6586e-08 1.8384869176588388 2.6587e-08 1.710370618585123 2.6588e-08 1.9435831547702358 2.6589e-08 1.773874586557058 2.659e-08 1.7938979930934005 2.6591e-08 1.8464964486223694 2.6592e-08 1.840091736692765 2.6593e-08 1.8477952461565372 2.6594e-08 1.8344596051738873 2.6595e-08 1.8748521096218653 2.6596e-08 1.7941144469135726 2.6597e-08 1.8141632155047744 2.6598e-08 1.7995780452563888 2.6599e-08 1.7774072789437814 2.66e-08 1.842292636057026 2.6601e-08 1.7560566644234858 2.6602e-08 1.8096205246673087 2.6603e-08 1.7279076970116132 2.6603999999999998e-08 1.8011459510545569 2.6605e-08 1.7064504414718493 2.6606e-08 1.8449993124004815 2.6606999999999998e-08 1.7779215496520104 2.6608e-08 1.8629897841370178 2.6609e-08 1.817279904669601 2.6609999999999998e-08 1.7740149941218566 2.6611e-08 1.8632502006361447 2.6612e-08 1.7908338721289145 2.6612999999999998e-08 1.8653993835257445 2.6614e-08 1.7861208789045 2.6615e-08 1.8072042527232355 2.6615999999999998e-08 1.8506925172230078 2.6617e-08 1.7961061688473912 2.6618e-08 1.7897666655952456 2.6618999999999998e-08 1.7541360358868785 2.662e-08 1.7245044921743713 2.6621e-08 1.8506899346491 2.6622e-08 1.8577901153506802 2.6623e-08 1.8518109532084768 2.6624e-08 1.82191228833205 2.6625e-08 1.7911244437434655 2.6626e-08 1.74695870991771 2.6627e-08 1.7729316874330592 2.6628e-08 1.7948371124274083 2.6629e-08 1.8058113075092908 2.663e-08 1.8123162662209615 2.6631e-08 1.7740577221159832 2.6632e-08 1.8369257035627673 2.6633e-08 1.7765550843203153 2.6634e-08 1.8980550644451701 2.6635e-08 1.7769543402688897 2.6636e-08 1.6928422692409961 2.6637e-08 1.7026346486656976 2.6638e-08 1.771886445146277 2.6638999999999998e-08 1.739805160314878 2.664e-08 1.8608727211192735 2.6641e-08 1.7922369058082654 2.6641999999999998e-08 1.8293770414473371 2.6643e-08 1.7915618411564742 2.6644e-08 1.7325261947244792 2.6644999999999998e-08 1.859192050217906 2.6646e-08 1.7927322690534646 2.6647e-08 1.7640988660857813 2.6647999999999998e-08 1.8486222110404622 2.6649e-08 1.7547340255701482 2.665e-08 1.7646874029822754 2.6650999999999998e-08 1.837396790041057 2.6652e-08 1.8104426461309828 2.6653e-08 1.8667553321047814 2.6653999999999998e-08 1.8658464613677277 2.6655e-08 1.6860474788937725 2.6656e-08 1.8019861738759273 2.6657e-08 1.8418804426100917 2.6658e-08 1.8366562518796907 2.6659e-08 1.7665744928783058 2.666e-08 1.7191974195272577 2.6661e-08 1.8826378626689082 2.6662e-08 1.8157158451736355 2.6663e-08 1.8428533001707603 2.6664e-08 1.7606814063713512 2.6665e-08 1.7525102267496164 2.6666e-08 1.7682164245024383 2.6667e-08 1.862160872277654 2.6668e-08 1.8330880270417051 2.6669e-08 1.8573596266809653 2.667e-08 1.7798360586866189 2.6671e-08 1.869574118839391 2.6672e-08 1.8314071888293442 2.6673e-08 1.7933944291783943 2.6673999999999998e-08 1.77749662713114 2.6675e-08 1.8248128352805464 2.6676e-08 1.8180318981759604 2.6676999999999998e-08 1.8667017080414565 2.6678e-08 1.7340591469847992 2.6679e-08 1.8120247866037853 2.6679999999999998e-08 1.7722140739245005 2.6681e-08 1.7052142321832884 2.6682e-08 1.8533395589141621 2.6682999999999998e-08 1.8265959582359144 2.6684e-08 1.8386667649738804 2.6685e-08 1.7877601586281848 2.6685999999999998e-08 1.7975448680938657 2.6687e-08 1.8319355554803562 2.6688e-08 1.8971562216090643 2.6688999999999998e-08 1.8339920918019028 2.669e-08 1.733234107187552 2.6691e-08 1.7588631070311105 2.6692e-08 1.8027400018311093 2.6693e-08 1.8230467652097564 2.6694e-08 1.8358141816260292 2.6695e-08 1.8326971275347113 2.6696e-08 1.769709042898556 2.6697e-08 1.8520182717800202 2.6698e-08 1.8063750686378341 2.6699e-08 1.8128396815162975 2.67e-08 1.7753881470201374 2.6701e-08 1.755410302407905 2.6702e-08 1.7469363536212013 2.6703e-08 1.8227463124170091 2.6704e-08 1.770880690490825 2.6705e-08 1.7686466071962805 2.6706e-08 1.7323241409478696 2.6707e-08 1.7295991097814554 2.6708e-08 1.6983531126787965 2.6708999999999998e-08 1.756029400579745 2.671e-08 1.8240719939200567 2.6711e-08 1.7402179522115733 2.6711999999999998e-08 1.754718786809075 2.6713e-08 1.7840927760242693 2.6714e-08 1.8418724730466165 2.6714999999999998e-08 1.829974771163741 2.6716e-08 1.7607573118979774 2.6717e-08 1.7225870597004351 2.6717999999999998e-08 1.7438777691268377 2.6719e-08 1.8901046434841298 2.672e-08 1.8481985498516562 2.6720999999999998e-08 1.8247560535326997 2.6722e-08 1.8466651973975203 2.6723e-08 1.8190067687772231 2.6723999999999998e-08 1.82903485662979 2.6725e-08 1.8429471195386842 2.6726e-08 1.6579980820618436 2.6727e-08 1.8514820733787536 2.6728e-08 1.8296498640747316 2.6729e-08 1.910811358204193 2.673e-08 1.8000892390708596 2.6731e-08 1.708009717811223 2.6732e-08 1.7759897305206018 2.6733e-08 1.8603039883018202 2.6734e-08 1.8292958876845729 2.6735e-08 1.8610242279295062 2.6736e-08 1.7635797097597548 2.6737e-08 1.7419082970764357 2.6738e-08 1.7672406761024464 2.6739e-08 1.7916320007756261 2.674e-08 1.7913919820459083 2.6741e-08 1.709424372007994 2.6742e-08 1.8446474098823082 2.6743e-08 1.6675949523451459 2.6743999999999998e-08 1.8004654241629425 2.6745e-08 1.8508166832790975 2.6746e-08 1.7710178454842906 2.6746999999999998e-08 1.818789864030943 2.6748e-08 1.8505707203858077 2.6749e-08 1.7979409318740267 2.6749999999999998e-08 1.718009983904248 2.6751e-08 1.8642526221739328 2.6752e-08 1.7995036085927625 2.6752999999999998e-08 1.7771499529406405 2.6754e-08 1.8295265308928241 2.6755e-08 1.8056347254493446 2.6755999999999998e-08 1.7193433284187936 2.6757e-08 1.7737621765264602 2.6758e-08 1.8449989844772003 2.6758999999999998e-08 1.8107145327590008 2.676e-08 1.8151706226004363 2.6761e-08 1.8060223368182147 2.6762e-08 1.8418468335225882 2.6763e-08 1.8223470544751141 2.6764e-08 1.6949582724167662 2.6765e-08 1.7278487335438462 2.6766e-08 1.7528088865526659 2.6767e-08 1.6863942947727062 2.6768e-08 1.6905788171809202 2.6769e-08 1.8631433008898453 2.677e-08 1.7427999122279374 2.6771e-08 1.8097722904276947 2.6772e-08 1.7823389284825808 2.6773e-08 1.8229999964604726 2.6774e-08 1.7496172131154448 2.6775e-08 1.6853916593972564 2.6776e-08 1.7593205199558264 2.6777e-08 1.8305961304986305 2.6778e-08 1.7055531186932882 2.6779e-08 1.6538721044013565 2.678e-08 1.7613278286198268 2.6781e-08 1.8830276658064264 2.6781999999999998e-08 1.746332024943669 2.6783e-08 1.751594663920725 2.6784e-08 1.7957633058109168 2.6784999999999998e-08 1.83276163288517 2.6786e-08 1.7793743443782892 2.6787e-08 1.7596371841067207 2.6787999999999998e-08 1.8555066241250149 2.6789e-08 1.9265035223352371 2.679e-08 1.7820202195326114 2.6790999999999998e-08 1.8448174781043165 2.6792e-08 1.898507283841718 2.6793e-08 1.7969009784998766 2.6793999999999998e-08 1.9143436021886746 2.6795e-08 1.8028293783772942 2.6796e-08 1.7213850027784305 2.6797e-08 1.7826759382573039 2.6798e-08 1.821825022258043 2.6799e-08 1.7494502089535797 2.68e-08 1.7588946908375875 2.6801e-08 1.862663241103856 2.6802e-08 1.9195768092893863 2.6803e-08 1.7027093458028832 2.6804e-08 1.7751518091901088 2.6805e-08 1.7993201190971984 2.6806e-08 1.852743214461787 2.6807e-08 1.8057454608422103 2.6808e-08 1.7961171050843894 2.6809e-08 1.7051641434587659 2.681e-08 1.8633132640029757 2.6811e-08 1.7929079636010756 2.6812e-08 1.8747708855626513 2.6813e-08 1.746197708417224 2.6814e-08 1.8270717661169131 2.6815e-08 1.7697643783026147 2.6816e-08 1.7299207923335027 2.6816999999999998e-08 1.7042446076039914 2.6818e-08 1.8031577777993397 2.6819e-08 1.8571896272262352 2.6819999999999998e-08 1.801891624968664 2.6821e-08 1.7581505929194068 2.6822e-08 1.8004075178642216 2.6822999999999998e-08 1.802648441355216 2.6824e-08 1.8742928964538184 2.6825e-08 1.815602932974484 2.6825999999999998e-08 1.8316882005840482 2.6827e-08 1.805500293616273 2.6828e-08 1.8157829027764554 2.6828999999999998e-08 1.771387400598062 2.683e-08 1.8302888519396456 2.6831e-08 1.8132795317194004 2.6831999999999998e-08 1.7795215243026992 2.6833e-08 1.8204986225772848 2.6834e-08 1.740172717685979 2.6835e-08 1.7746106224490557 2.6836e-08 1.7035177787119493 2.6837e-08 1.790207816406995 2.6838e-08 1.719825619136566 2.6839e-08 1.799575973787586 2.684e-08 1.7764993107394003 2.6841e-08 1.8492800261434437 2.6842e-08 1.8157010741456812 2.6843e-08 1.8660281211608951 2.6844e-08 1.784812906288218 2.6845e-08 1.8898872573643832 2.6846e-08 1.7350920012107023 2.6847e-08 1.8513552108901903 2.6848e-08 1.8705174263612492 2.6849e-08 1.8097641535804043 2.685e-08 1.7882586218660015 2.6851e-08 1.919290905280417 2.6851999999999998e-08 1.7676318379862646 2.6853e-08 1.7835970358127935 2.6854e-08 1.8617003830387187 2.6854999999999998e-08 1.9008896837356324 2.6856e-08 1.8390876900579138 2.6857e-08 1.7890227176546432 2.6857999999999998e-08 1.8213391648230675 2.6859e-08 1.880450474420448 2.686e-08 1.7898375751066664 2.6860999999999998e-08 1.759648953152222 2.6862e-08 1.8311035522520624 2.6863e-08 1.778965481525614 2.6863999999999998e-08 1.7268604177521834 2.6865e-08 1.752795972975834 2.6866e-08 1.8536630577068298 2.6866999999999998e-08 1.7203813123140468 2.6868e-08 1.917604074160826 2.6869e-08 1.8427598576825979 2.687e-08 1.78422800998475 2.6871e-08 1.7474538642592754 2.6872e-08 1.8183888825190304 2.6873e-08 1.7638925877336458 2.6874e-08 1.8650122975797543 2.6875e-08 1.8389094493459157 2.6876e-08 1.8315674165436093 2.6877e-08 1.752469333247259 2.6878e-08 1.8420989691972152 2.6879e-08 1.8644907172500655 2.688e-08 1.6975093425891163 2.6881e-08 1.7878300777560117 2.6882e-08 1.8187632712674127 2.6883e-08 1.8816209522426084 2.6884e-08 1.7857635913635888 2.6885e-08 1.7650255467311629 2.6886e-08 1.8490069194259704 2.6886999999999998e-08 1.7436662369932283 2.6888e-08 1.7527947411493896 2.6889e-08 1.8670645490309428 2.6889999999999998e-08 1.8312811837883154 2.6891e-08 1.7280851088443596 2.6892e-08 1.7362406861133808 2.6892999999999998e-08 1.77859996788158 2.6894e-08 1.7941267662619127 2.6895e-08 1.8190003175658644 2.6895999999999998e-08 1.777362255702455 2.6897e-08 1.7779191583047234 2.6898e-08 1.7769705273065561 2.6898999999999998e-08 1.8166364215339315 2.69e-08 1.8530544871878025 2.6901e-08 1.8318238526954045 2.6901999999999998e-08 1.8614517064005058 2.6903e-08 1.7530307685284139 2.6904e-08 1.8158135277997085 2.6905e-08 1.8036792199707459 2.6906e-08 1.7753888340788258 2.6907e-08 1.7421155960313304 2.6908e-08 1.797068975758949 2.6909e-08 1.8003410046748198 2.691e-08 1.83913647598463 2.6911e-08 1.8335813555447855 2.6912e-08 1.8351800913645608 2.6913e-08 1.9453290366647487 2.6914e-08 1.775994436288897 2.6915e-08 1.8423866516339846 2.6916e-08 1.7645803782745801 2.6917e-08 1.8431586908334383 2.6918e-08 1.7887867436393083 2.6919e-08 1.8173509465463953 2.692e-08 1.8300809971844696 2.6921e-08 1.8755836663532834 2.6921999999999998e-08 1.7098035828597307 2.6923e-08 1.8208308050327942 2.6924e-08 1.8559370219453717 2.6924999999999998e-08 1.7950356030805703 2.6926e-08 1.8962066679579654 2.6927e-08 1.7461066852238185 2.6927999999999998e-08 1.7127483977627076 2.6929e-08 1.904147509569396 2.693e-08 1.7896730261951688 2.6930999999999998e-08 1.8411057142665017 2.6932e-08 1.8643402644953964 2.6933e-08 1.8477449296977089 2.6933999999999998e-08 1.8129507648032968 2.6935e-08 1.7504070811541472 2.6936e-08 1.8374120655040707 2.6936999999999998e-08 1.7627637647442944 2.6938e-08 1.8221941660343401 2.6939e-08 1.793308339209662 2.694e-08 1.7881134666804872 2.6941e-08 1.809779132025061 2.6942e-08 1.7998571656705955 2.6943e-08 1.6698530056916359 2.6944e-08 1.7419566791820016 2.6945e-08 1.9001901336984965 2.6946e-08 1.7296300360244852 2.6947e-08 1.861695895138569 2.6948e-08 1.7558757348965481 2.6949e-08 1.8338840894950874 2.695e-08 1.7478331772769748 2.6951e-08 1.7926257413855637 2.6952e-08 1.8503602147741296 2.6953e-08 1.7850117122903932 2.6954e-08 1.6897017526153373 2.6955e-08 1.8006116549311177 2.6956e-08 1.7545144154389016 2.6957e-08 1.7525255150566528 2.6958e-08 1.8814797512913792 2.6959e-08 1.8157091977505542 2.6959999999999998e-08 1.8181255564269208 2.6961e-08 1.8468788621661587 2.6962e-08 1.7052322750155355 2.6962999999999998e-08 1.9444181099447997 2.6964e-08 1.8876854801487224 2.6965e-08 1.8021680157032052 2.6965999999999998e-08 1.850596470958297 2.6967e-08 1.8307354701891416 2.6968e-08 1.854832189466265 2.6968999999999998e-08 1.753647870245992 2.697e-08 1.8019231106860063 2.6971e-08 1.719759288080859 2.6971999999999998e-08 1.73127002149618 2.6973e-08 1.8150587127211464 2.6974e-08 1.774748323413279 2.6975e-08 1.8151677103586787 2.6976e-08 1.7928062861383247 2.6977e-08 1.77042106511485 2.6978e-08 1.8228951000092297 2.6979e-08 1.7200953984620213 2.698e-08 1.7607162488821355 2.6981e-08 1.7763384828955064 2.6982e-08 1.7741005065532096 2.6983e-08 1.7661511582281035 2.6984e-08 1.7893720916222522 2.6985e-08 1.860027294721191 2.6986e-08 1.7939577863426925 2.6987e-08 1.809876372434203 2.6988e-08 1.8922317706106775 2.6989e-08 1.752201241784878 2.699e-08 1.7659304897417918 2.6991e-08 1.8047387983372993 2.6992e-08 1.7354214281348188 2.6993e-08 1.7548855988249623 2.6994e-08 1.797382587953675 2.6994999999999998e-08 1.7182628229694 2.6996e-08 1.784607880577343 2.6997e-08 1.83658465217214 2.6997999999999998e-08 1.6993127462468383 2.6999e-08 1.8216868231902779 2.7e-08 1.8293998188971263 2.7000999999999998e-08 1.8142598751032857 2.7002e-08 1.7964431215322652 2.7003e-08 1.8863859868715667 2.7003999999999998e-08 1.8603103294215657 2.7005e-08 1.8519087363823894 2.7006e-08 1.759465414140928 2.7006999999999998e-08 1.797713839171656 2.7008e-08 1.7577580393498036 2.7009e-08 1.7537410233234219 2.7009999999999998e-08 1.814855630872306 2.7011e-08 1.8620866301482097 2.7012e-08 1.6551190595674874 2.7013e-08 1.849906068483744 2.7014e-08 1.8822032420085968 2.7015e-08 1.7777694010131064 2.7016e-08 1.8209046135818001 2.7017e-08 1.8975159283541838 2.7018e-08 1.8097302100891215 2.7019e-08 1.7305159861687474 2.702e-08 1.8029632122880304 2.7021e-08 1.8675280800183862 2.7022e-08 1.8261382212228536 2.7023e-08 1.8013263689370818 2.7024e-08 1.7859984636925699 2.7025e-08 1.860803106219276 2.7026e-08 1.7998888826193253 2.7027e-08 1.8431245776298146 2.7028e-08 1.8868943340151532 2.7029e-08 1.849841548876931 2.7029999999999998e-08 1.7693131933099508 2.7031e-08 1.8933981988313784 2.7032e-08 1.6681856771078563 2.7032999999999998e-08 1.797093562673789 2.7034e-08 1.7961148560909557 2.7035e-08 1.7720188764070859 2.7035999999999998e-08 1.7928799866203802 2.7037e-08 1.7955769898380567 2.7038e-08 1.8672464255534886 2.7038999999999998e-08 1.7096834170742015 2.704e-08 1.8021463516099354 2.7041e-08 1.771201024825631 2.7041999999999998e-08 1.7753922574305894 2.7043e-08 1.7752642324262773 2.7044e-08 1.7506678612171367 2.7044999999999998e-08 1.7423771885367247 2.7046e-08 1.742462325704257 2.7047e-08 1.7960748262910922 2.7048e-08 1.856617209923005 2.7049e-08 1.8302121921637333 2.705e-08 1.7469306305522765 2.7051e-08 1.8397804270328186 2.7052e-08 1.8027086821255545 2.7053e-08 1.7893714750246867 2.7054e-08 1.8615505867338729 2.7055e-08 1.790376321272493 2.7056e-08 1.8045842593560084 2.7057e-08 1.7739968142099845 2.7058e-08 1.7915619575586843 2.7059e-08 1.7814517244041317 2.706e-08 1.745829452145743 2.7061e-08 1.7936225710622857 2.7062e-08 1.8395269761757262 2.7063e-08 1.7961218324304211 2.7064e-08 1.7694616114769497 2.7064999999999998e-08 1.7990653551148632 2.7066e-08 1.7678453706166095 2.7067e-08 1.7732232152970226 2.7067999999999998e-08 1.8260719075985063 2.7069e-08 1.7402684411164522 2.707e-08 1.7569964198340993 2.7070999999999998e-08 1.836175109161195 2.7072e-08 1.7842290117503146 2.7073e-08 1.820482577363001 2.7073999999999998e-08 1.7763664087607238 2.7075e-08 1.7773400408226467 2.7076e-08 1.7386810856369137 2.7076999999999998e-08 1.797746134993128 2.7078e-08 1.7910037990509429 2.7079e-08 1.7110583870772895 2.7079999999999998e-08 1.7355714363865582 2.7081e-08 1.7559139673349098 2.7082e-08 1.8173373770200465 2.7083e-08 1.7847984587340058 2.7084e-08 1.7704427316314333 2.7085e-08 1.8114261785099033 2.7086e-08 1.8245591495755753 2.7087e-08 1.891158678579956 2.7088e-08 1.7963166438809928 2.7089e-08 1.9001079687322453 2.709e-08 1.7978847232159383 2.7091e-08 1.7070563519886222 2.7092e-08 1.8032200449438682 2.7093e-08 1.7566029420814864 2.7094e-08 1.750905644609441 2.7095e-08 1.779974851904138 2.7096e-08 1.7499894789000976 2.7097e-08 1.8397778692227353 2.7098e-08 1.8508866464779252 2.7099e-08 1.861042801875971 2.7099999999999998e-08 1.8143021391458363 2.7101e-08 1.7624621954478812 2.7102e-08 1.8198887553261054 2.7102999999999998e-08 1.71628285690952 2.7104e-08 1.8499148241053163 2.7105e-08 1.7952333143655599 2.7105999999999998e-08 1.7928675878975586 2.7107e-08 1.8710574467723784 2.7108e-08 1.8764721106982096 2.7108999999999998e-08 1.8342743606153598 2.711e-08 1.72707833279454 2.7111e-08 1.7388637552686736 2.7111999999999998e-08 1.8328798346866528 2.7113e-08 1.8181405872942193 2.7114e-08 1.7960526204524752 2.7114999999999998e-08 1.8027194828232647 2.7116e-08 1.7866097282746387 2.7117e-08 1.8572828085781272 2.7118e-08 1.7554539866882146 2.7119e-08 1.7839118727616081 2.712e-08 1.8277674292082586 2.7121e-08 1.7609554674098593 2.7122e-08 1.7916970936200478 2.7123e-08 1.8360438265393273 2.7124e-08 1.7929896760943278 2.7125e-08 1.7766453301977005 2.7126e-08 1.85660577568609 2.7127e-08 1.775041116278091 2.7128e-08 1.667908800898494 2.7129e-08 1.7947718600508014 2.713e-08 1.794728021927615 2.7131e-08 1.7199336714557918 2.7132e-08 1.8326138087818886 2.7133e-08 1.8399051370731303 2.7134e-08 1.7957564359416527 2.7134999999999998e-08 1.7946942406717403 2.7136e-08 1.7534136644070408 2.7137e-08 1.7936431855960806 2.7137999999999998e-08 1.730128139419738 2.7139e-08 1.8561694759860492 2.714e-08 1.854031735103557 2.7140999999999998e-08 1.801715021348664 2.7142e-08 1.847892252431021 2.7143e-08 1.7714758587463693 2.7143999999999998e-08 1.756638783798245 2.7145e-08 1.7980337944026588 2.7146e-08 1.8323034406446053 2.7146999999999998e-08 1.8703987835746088 2.7148e-08 1.712750735575462 2.7149e-08 1.8198826833493573 2.7149999999999998e-08 1.811722783209707 2.7151e-08 1.7706222192658037 2.7152e-08 1.8104599554816878 2.7153e-08 1.8193890763711136 2.7154e-08 1.7825037726506852 2.7155e-08 1.8064369214321963 2.7156e-08 1.745838608392822 2.7157e-08 1.8614037695680712 2.7158e-08 1.6976934990062105 2.7159e-08 1.7921220367424078 2.716e-08 1.7569375283282644 2.7161e-08 1.8069002602090831 2.7162e-08 1.7671921675843718 2.7163e-08 1.8982716500289607 2.7164e-08 1.7799436499303243 2.7165e-08 1.8298763642447464 2.7166e-08 1.8357919811376602 2.7167e-08 1.8374343600994498 2.7168e-08 1.8600076204915703 2.7169e-08 1.8196563353200177 2.717e-08 1.833139980613313 2.7171e-08 1.793027659147592 2.7172e-08 1.777929129537794 2.7172999999999998e-08 1.8783836079279215 2.7174e-08 1.7126774896625312 2.7175e-08 1.8138924145362982 2.7175999999999998e-08 1.7808279042373196 2.7177e-08 1.8325391651555911 2.7178e-08 1.8003516537685065 2.7178999999999998e-08 1.7947068893153457 2.718e-08 1.7162998479180713 2.7181e-08 1.8317978169716458 2.7181999999999998e-08 1.831477247858988 2.7183e-08 1.8307188180146818 2.7184e-08 1.691500227575337 2.7184999999999998e-08 1.7876328788840548 2.7186e-08 1.7787766436348875 2.7187e-08 1.700484218024144 2.7187999999999998e-08 1.7921159597507492 2.7189e-08 1.8769893441285177 2.719e-08 1.8581117323860352 2.7191e-08 1.7788908267457617 2.7192e-08 1.7445630233238738 2.7193e-08 1.8137051385562322 2.7194e-08 1.7823902116153865 2.7195e-08 1.8451969823697625 2.7196e-08 1.8057434586330026 2.7197e-08 1.8082411907533034 2.7198e-08 1.817205362626014 2.7199e-08 1.8220027161879213 2.72e-08 1.7490659825555461 2.7201e-08 1.773310096045568 2.7202e-08 1.8546714927928456 2.7203e-08 1.7734709915783655 2.7204e-08 1.800127330566679 2.7205e-08 1.8124501109685456 2.7206e-08 1.7355505508785747 2.7207e-08 1.7950262354512905 2.7207999999999998e-08 1.807329901245473 2.7209e-08 1.7171670882689305 2.721e-08 1.8431658482511937 2.7210999999999998e-08 1.8009526753544813 2.7212e-08 1.8206568261488303 2.7213e-08 1.806282737623025 2.7213999999999998e-08 1.730600984456352 2.7215e-08 1.754881765023561 2.7216e-08 1.8018163485846364 2.7216999999999998e-08 1.7952292233528517 2.7218e-08 1.8610142514265016 2.7219e-08 1.8251845107146412 2.7219999999999998e-08 1.8369459785466238 2.7221e-08 1.778420204534483 2.7222e-08 1.798187449949716 2.7222999999999998e-08 1.8098738955140126 2.7224e-08 1.8001603258824974 2.7225e-08 1.886093594544992 2.7226e-08 1.7624198735781302 2.7227e-08 1.7544388541963443 2.7228e-08 1.771117483747754 2.7229e-08 1.8699704398321144 2.723e-08 1.7440956313982343 2.7231e-08 1.7395415751142045 2.7232e-08 1.758407141497767 2.7233e-08 1.7240696941616251 2.7234e-08 1.7992247009644116 2.7235e-08 1.8494426732713702 2.7236e-08 1.8002272928477563 2.7237e-08 1.8292511229444905 2.7238e-08 1.8766904131703788 2.7239e-08 1.8339151166649004 2.724e-08 1.8100990679959041 2.7241e-08 1.8047295776176715 2.7242e-08 1.8128916670967183 2.7242999999999998e-08 1.8037708457407569 2.7244e-08 1.8637700662903733 2.7245e-08 1.8503588445536245 2.7245999999999998e-08 1.8087434932237103 2.7247e-08 1.7463902490696113 2.7248e-08 1.8257265855243836 2.7248999999999998e-08 1.828847565206947 2.725e-08 1.769491947744255 2.7251e-08 1.763272220805525 2.7251999999999998e-08 1.8968309107222825 2.7253e-08 1.8057054798534733 2.7254e-08 1.731101730686288 2.7254999999999998e-08 1.8521435228651173 2.7256e-08 1.7968585009287552 2.7257e-08 1.7633559329936175 2.7257999999999998e-08 1.8342978138944397 2.7259e-08 1.8662711389027933 2.726e-08 1.7724559827607287 2.7261e-08 1.865749753680759 2.7262e-08 1.7823606445976539 2.7263e-08 1.8010642460650037 2.7264e-08 1.72037993858718 2.7265e-08 1.8209250884695902 2.7266e-08 1.7794893319582648 2.7267e-08 1.7579069688105124 2.7268e-08 1.778639502082417 2.7269e-08 1.7806181734954503 2.727e-08 1.7944950463347187 2.7271e-08 1.8257964778961742 2.7272e-08 1.8023542347758648 2.7273e-08 1.7917549473299927 2.7274e-08 1.7836855987403308 2.7275e-08 1.93825165276654 2.7276e-08 1.8098006295721856 2.7277e-08 1.773850568479724 2.7277999999999998e-08 1.7400226364584928 2.7279e-08 1.80663110198842 2.728e-08 1.9036088350883724 2.7280999999999998e-08 1.769257286810825 2.7282e-08 1.7131073956525231 2.7283e-08 1.8551748818094416 2.7283999999999998e-08 1.8625798572630843 2.7285e-08 1.7491769393030183 2.7286e-08 1.7395136437735041 2.7286999999999998e-08 1.7540499680652935 2.7288e-08 1.7991307098712013 2.7289e-08 1.774252267220231 2.7289999999999998e-08 1.8126678349720773 2.7291e-08 1.6923396412295373 2.7292e-08 1.8601482100788442 2.7292999999999998e-08 1.774628063957344 2.7294e-08 1.8244522201377638 2.7295e-08 1.7866749672470934 2.7296e-08 1.8234187859254738 2.7297e-08 1.846380926401121 2.7298e-08 1.8073758517739205 2.7299e-08 1.7019551908423725 2.73e-08 1.819285366666852 2.7301e-08 1.7827268248263235 2.7302e-08 1.8198764375816714 2.7303e-08 1.8697063874288213 2.7304e-08 1.8247824098771703 2.7305e-08 1.8302825212688674 2.7306e-08 1.7173615219615581 2.7307e-08 1.8275226471277544 2.7308e-08 1.8216099991376253 2.7309e-08 1.748455886453468 2.731e-08 1.9425046915418658 2.7311e-08 1.7781557692226713 2.7312e-08 1.8072250897638615 2.7312999999999998e-08 1.8128128513397266 2.7314e-08 1.8422415181221115 2.7315e-08 1.733571582107073 2.7315999999999998e-08 1.7833045342256082 2.7317e-08 1.8431192788778663 2.7318e-08 1.7664415429577542 2.7318999999999998e-08 1.8264959958489906 2.732e-08 1.7845413413729645 2.7321e-08 1.8212635703901991 2.7321999999999998e-08 1.8176180662412735 2.7323e-08 1.7921020403638783 2.7324e-08 1.794268128865046 2.7324999999999998e-08 1.8990743010258215 2.7326e-08 1.8339475325983703 2.7327e-08 1.8046862097766205 2.7327999999999998e-08 1.9357348013629085 2.7329e-08 1.8579725024326765 2.733e-08 1.7810106783858481 2.7331e-08 1.8011485188553003 2.7332e-08 1.8388165632133904 2.7333e-08 1.7606270323339122 2.7334e-08 1.792460079795883 2.7335e-08 1.8144337427195723 2.7336e-08 1.675238713164257 2.7337e-08 1.708875773134857 2.7338e-08 1.8056084841983666 2.7339e-08 1.8869017443732197 2.734e-08 1.6770745470648811 2.7341e-08 1.8005011267653037 2.7342e-08 1.714529587903246 2.7343e-08 1.8550194567346652 2.7344e-08 1.7519064223506335 2.7345e-08 1.8226875999348742 2.7346e-08 1.7457152909177724 2.7347e-08 1.774057913616508 2.7348e-08 1.799399045632618 2.7349e-08 1.868249448953915 2.735e-08 1.743357576776331 2.7350999999999998e-08 1.8791886447925032 2.7352e-08 1.8554339735214092 2.7353e-08 1.799748719486364 2.7353999999999998e-08 1.846671129674895 2.7355e-08 1.7563427944609729 2.7356e-08 1.6970426290879876 2.7356999999999998e-08 1.7726780965006517 2.7358e-08 1.7910821078345958 2.7359e-08 1.7898458434780236 2.7359999999999998e-08 1.7888884603831885 2.7361e-08 1.8059205219429966 2.7362e-08 1.7507725150692224 2.7362999999999998e-08 1.72913876732147 2.7364e-08 1.7031867379384382 2.7365e-08 1.754219327363752 2.7366e-08 1.8264357284737 2.7367e-08 1.7736166059848855 2.7368e-08 1.8254705705564869 2.7369e-08 1.7594346781597516 2.737e-08 1.7898360096629307 2.7371e-08 1.7808702971331454 2.7372e-08 1.937707606897016 2.7373e-08 1.8111417825937373 2.7374e-08 1.8321040957250676 2.7375e-08 1.8067482758226163 2.7376e-08 1.8648838344540983 2.7377e-08 1.7789600940474826 2.7378e-08 1.8153295764903834 2.7379e-08 1.8772964400552443 2.738e-08 1.8050079127844325 2.7381e-08 1.7399314059977626 2.7382e-08 1.7950400586675355 2.7383e-08 1.7260547944077052 2.7384e-08 1.7512153182795438 2.7385e-08 1.7208099907925298 2.7385999999999998e-08 1.8253621818571104 2.7387e-08 1.7883945799688294 2.7388e-08 1.8344165731737028 2.7388999999999998e-08 1.785430757360849 2.739e-08 1.7245923048679577 2.7391e-08 1.8803014587981393 2.7391999999999998e-08 1.8191123950188537 2.7393e-08 1.8426599269816133 2.7394e-08 1.7526551690968921 2.7394999999999998e-08 1.7376459204772803 2.7396e-08 1.8354518359332606 2.7397e-08 1.8861439620855116 2.7397999999999998e-08 1.8668283346201267 2.7399e-08 1.8138188475564565 2.74e-08 1.732667461635814 2.7400999999999998e-08 1.681440978247869 2.7402e-08 1.8036079835701628 2.7403e-08 1.8003902395245177 2.7404e-08 1.7924684252255998 2.7405e-08 1.7942633941579993 2.7406e-08 1.7908707844115328 2.7407e-08 1.875863525670864 2.7408e-08 1.8055426790758609 2.7409e-08 1.791501092995787 2.741e-08 1.7486789155943154 2.7411e-08 1.8170891369853956 2.7412e-08 1.7481545207543416 2.7413e-08 1.8553191635223953 2.7414e-08 1.7962952641984962 2.7415e-08 1.8570736286631548 2.7416e-08 1.7896073022205512 2.7417e-08 1.7638208242579467 2.7418e-08 1.8276184730626623 2.7419e-08 1.7862624249139065 2.742e-08 1.8659458068608077 2.7420999999999998e-08 1.8050085481783182 2.7422e-08 1.8563197343482045 2.7423e-08 1.819771633863591 2.7423999999999998e-08 1.7911520720399803 2.7425e-08 1.7623096364527524 2.7426e-08 1.8238935593117818 2.7426999999999998e-08 1.8188928263039075 2.7428e-08 1.7074080121915687 2.7429e-08 1.7712042018067065 2.7429999999999998e-08 1.8167975041201732 2.7431e-08 1.777841206656404 2.7432e-08 1.9013287078435783 2.7432999999999998e-08 1.7871363255445378 2.7434e-08 1.7808292594046136 2.7435e-08 1.7928865222180461 2.7435999999999998e-08 1.8380604004890235 2.7437e-08 1.7968190018207195 2.7438e-08 1.7864065539300469 2.7439e-08 1.8501746958479155 2.744e-08 1.768094021853891 2.7441e-08 1.8306465796435911 2.7442e-08 1.7672898629202418 2.7443e-08 1.8061875748636207 2.7444e-08 1.7922162016923773 2.7445e-08 1.707128126299052 2.7446e-08 1.8507373087936403 2.7447e-08 1.7961428471146446 2.7448e-08 1.7867346611651478 2.7449e-08 1.8626097410141633 2.745e-08 1.8511215531115388 2.7451e-08 1.8290074337403046 2.7452e-08 1.7677814284018973 2.7453e-08 1.7907730112932931 2.7454e-08 1.7590506983363359 2.7455e-08 1.7796721910201485 2.7455999999999998e-08 1.7782339767236692 2.7457e-08 1.8305257297131772 2.7458e-08 1.7977669660124957 2.7458999999999998e-08 1.7559995793191914 2.746e-08 1.8154638832360912 2.7461e-08 1.7859686752873363 2.7461999999999998e-08 1.8069886418206558 2.7463e-08 1.8758785316147595 2.7464e-08 1.7752866675842423 2.7464999999999998e-08 1.8343371108831756 2.7466e-08 1.8607240106262022 2.7467e-08 1.7546528559562131 2.7467999999999998e-08 1.7896446350946777 2.7469e-08 1.7919595828118289 2.747e-08 1.8613006622290378 2.7470999999999998e-08 1.7766298331522372 2.7472e-08 1.7514634430870537 2.7473e-08 1.7659850759861566 2.7474e-08 1.6743502368850685 2.7475e-08 1.8057937957810835 2.7476e-08 1.8029949290670593 2.7477e-08 1.7218245162628039 2.7478e-08 1.7744479501114725 2.7479e-08 1.8686784605926523 2.748e-08 1.820197151207609 2.7481e-08 1.7745041216373387 2.7482e-08 1.7982034117912382 2.7483e-08 1.8668369345913893 2.7484e-08 1.7078335308387 2.7485e-08 1.8910838875320892 2.7486e-08 1.8218852239593615 2.7487e-08 1.821013219665336 2.7488e-08 1.7885506662246735 2.7489e-08 1.8264317986185405 2.749e-08 1.7854617702297566 2.7490999999999998e-08 1.7747844261870636 2.7492e-08 1.7519695895956127 2.7493e-08 1.76842357241298 2.7493999999999998e-08 1.8231774104112561 2.7495e-08 1.7858316382568957 2.7496e-08 1.8775991157490055 2.7496999999999998e-08 1.8888490144021568 2.7498e-08 1.8135449014020493 2.7499e-08 1.8017797639992927 2.7499999999999998e-08 1.8192285067421132 2.7501e-08 1.7607369776904083 2.7502e-08 1.8130887298634921 2.7502999999999998e-08 1.829529037454714 2.7504e-08 1.760658936185404 2.7505e-08 1.7169073445461882 2.7505999999999998e-08 1.707547454622839 2.7507e-08 1.8819459663534015 2.7508e-08 1.8234760959257412 2.7509e-08 1.8504008422118505 2.751e-08 1.8505723543424186 2.7511e-08 1.732018003709929 2.7512e-08 1.7394165581528398 2.7513e-08 1.7726925826662951 2.7514e-08 1.81481170408563 2.7515e-08 1.8587049304624612 2.7516e-08 1.8973959578902433 2.7517e-08 1.7797522040801106 2.7518e-08 1.7572056205953073 2.7519e-08 1.8265913056349308 2.752e-08 1.8146013227736069 2.7521e-08 1.8312973306273077 2.7522e-08 1.8148833596303944 2.7523e-08 1.7666419374520075 2.7524e-08 1.828818188463617 2.7525e-08 1.752367540663804 2.7525999999999998e-08 1.8449433958625652 2.7527e-08 1.8373783653553002 2.7528e-08 1.7424375110500026 2.7528999999999998e-08 1.8351398929341112 2.753e-08 1.8417007055447197 2.7531e-08 1.8454804314158184 2.7531999999999998e-08 1.8157786726782752 2.7533e-08 1.8401837889506205 2.7534e-08 1.896219023145882 2.7534999999999998e-08 1.8002355583064178 2.7536e-08 1.9076932650677678 2.7537e-08 1.793678448170283 2.7537999999999998e-08 1.8498984270920893 2.7539e-08 1.7122580214768912 2.754e-08 1.822494597556648 2.7540999999999998e-08 1.728941944239563 2.7542e-08 1.7537332076054521 2.7543e-08 1.8390458670288963 2.7544e-08 1.8617467848860618 2.7545e-08 1.7425855553005458 2.7546e-08 1.7772511908028552 2.7547e-08 1.8071629395058606 2.7548e-08 1.8693096436600616 2.7549e-08 1.8062767883069166 2.755e-08 1.7801707956281416 2.7551e-08 1.8019279493688063 2.7552e-08 1.7316114700388636 2.7553e-08 1.83513955084848 2.7554e-08 1.7717545818157387 2.7555e-08 1.8027806710797365 2.7556e-08 1.761875389303532 2.7557e-08 1.7249703753733905 2.7558e-08 1.8596260162050737 2.7559e-08 1.8746532654384618 2.756e-08 1.7910587178293258 2.7561e-08 1.8202806712537143 2.7562e-08 1.7906042126419266 2.7563e-08 1.7713175748777414 2.7563999999999998e-08 1.7990290930395312 2.7565e-08 1.7821307796095631 2.7566e-08 1.8161952735484534 2.7566999999999998e-08 1.8633069746254038 2.7568e-08 1.8383275113116244 2.7569e-08 1.8155601946990314 2.7569999999999998e-08 1.8025220207714974 2.7571e-08 1.8338556817697957 2.7572e-08 1.8070788190643123 2.7572999999999998e-08 1.8401858380043474 2.7574e-08 1.7314630882787077 2.7575e-08 1.8886761015700169 2.7575999999999998e-08 1.7388871919350588 2.7577e-08 1.7751735422011623 2.7578e-08 1.7896527767693822 2.7578999999999998e-08 1.7965293020081448 2.758e-08 1.8343882138061418 2.7581e-08 1.7617544258051439 2.7582e-08 1.8601057946435389 2.7583e-08 1.7710066335988786 2.7584e-08 1.867905265802687 2.7585e-08 1.7441959592986838 2.7586e-08 1.794505428707258 2.7587e-08 1.8068338266242456 2.7588e-08 1.752776941440061 2.7589e-08 1.8281657187946865 2.759e-08 1.8422713794266659 2.7591e-08 1.802678263173726 2.7592e-08 1.8504929536601955 2.7593e-08 1.7397388080008345 2.7594e-08 1.755584517356781 2.7595e-08 1.8173769684028 2.7596e-08 1.8194096159712827 2.7597e-08 1.806600453684017 2.7598e-08 1.8507840182704125 2.7598999999999998e-08 1.858569370449764 2.76e-08 1.7384398042469003 2.7601e-08 1.9054104715412794 2.7601999999999998e-08 1.8543602248879987 2.7603e-08 1.8919011807036898 2.7604e-08 1.8583914530896113 2.7604999999999998e-08 1.7768111755110756 2.7606e-08 1.776339237499484 2.7607e-08 1.8451757830790365 2.7607999999999998e-08 1.846112372356375 2.7609e-08 1.8156191685117622 2.761e-08 1.7610009098316624 2.7610999999999998e-08 1.784586885418866 2.7612e-08 1.7688249305510197 2.7613e-08 1.8001737109688514 2.7613999999999998e-08 1.799898018553806 2.7615e-08 1.7645586250531171 2.7616e-08 1.8508370878390075 2.7617e-08 1.8044029210361567 2.7618e-08 1.7923479403084939 2.7619e-08 1.751362238686201 2.762e-08 1.866613580730088 2.7621e-08 1.7867722997262736 2.7622e-08 1.6976061013068482 2.7623e-08 1.8587565346126045 2.7624e-08 1.8067807002232064 2.7625e-08 1.738956842202619 2.7626e-08 1.7010100180143695 2.7627e-08 1.7734102093555575 2.7628e-08 1.7975462048175852 2.7629e-08 1.8089076708531235 2.763e-08 1.8475837510408772 2.7631e-08 1.7866127772460356 2.7632e-08 1.7959725879026005 2.7633e-08 1.8760549551112737 2.7633999999999998e-08 1.8272067406909265 2.7635e-08 1.8217850123060095 2.7636e-08 1.7623294725433618 2.7636999999999998e-08 1.8150913216780291 2.7638e-08 1.7740605115074144 2.7639e-08 1.8961942585028253 2.7639999999999998e-08 1.7698819472628733 2.7641e-08 1.7989712842364491 2.7642e-08 1.895232818548177 2.7642999999999998e-08 1.7159073107908556 2.7644e-08 1.7671232098681287 2.7645e-08 1.8168179678892877 2.7645999999999998e-08 1.8184369125872635 2.7647e-08 1.8218905211717793 2.7648e-08 1.7733270888058539 2.7648999999999998e-08 1.7534847120091304 2.765e-08 1.8143027327108738 2.7651e-08 1.8052979443555621 2.7652e-08 1.875223017477137 2.7653e-08 1.8883926441419912 2.7654e-08 1.7992951168592215 2.7655e-08 1.8105661546641736 2.7656e-08 1.7804278117527943 2.7657e-08 1.8206041077882187 2.7658e-08 1.756027718950849 2.7659e-08 1.7979387255613433 2.766e-08 1.7667830772469246 2.7661e-08 1.8418697368580594 2.7662e-08 1.8407473358507527 2.7663e-08 1.7919885305457444 2.7664e-08 1.8333198036973093 2.7665e-08 1.7810840416426883 2.7666e-08 1.800554197950294 2.7667e-08 1.8028143701859067 2.7668e-08 1.7107196405946543 2.7668999999999998e-08 1.904792079752378 2.767e-08 1.8481602915959627 2.7671e-08 1.782361475348982 2.7671999999999998e-08 1.749265972026789 2.7673e-08 1.8084391625907295 2.7674e-08 1.9192258743921697 2.7674999999999998e-08 1.7890255678619624 2.7676e-08 1.7828986534676594 2.7677e-08 1.7913941215501472 2.7677999999999998e-08 1.7960043899197202 2.7679e-08 1.8120201375261853 2.768e-08 1.7880020741996587 2.7680999999999998e-08 1.8335714980543718 2.7682e-08 1.813741416590983 2.7683e-08 1.7419257190644235 2.7683999999999998e-08 1.870030663052025 2.7685e-08 1.8384722855823148 2.7686e-08 1.8189475928238634 2.7687e-08 1.7775194171604352 2.7688e-08 1.772900633555512 2.7689e-08 1.8117944474792556 2.769e-08 1.7409509086174806 2.7691e-08 1.818582337946683 2.7692e-08 1.8737186847777014 2.7693e-08 1.8531281437248512 2.7694e-08 1.7197496172084792 2.7695e-08 1.7804056483788395 2.7696e-08 1.7451409962445112 2.7697e-08 1.7653722984237126 2.7698e-08 1.7223606173470107 2.7699e-08 1.8617864287332466 2.77e-08 1.7587552689039898 2.7701e-08 1.8106606181024953 2.7702e-08 1.8604042950857618 2.7703e-08 1.8162010199835448 2.7703999999999998e-08 1.8776983074140159 2.7705e-08 1.779675229913686 2.7706e-08 1.767253799128571 2.7706999999999998e-08 1.7829797213260046 2.7708e-08 1.8623973703734298 2.7709e-08 1.8198617995177087 2.7709999999999998e-08 1.8053016706902048 2.7711e-08 1.767808964691731 2.7712e-08 1.8385531702657312 2.7712999999999998e-08 1.8207763921439641 2.7714e-08 1.7775970905749834 2.7715e-08 1.8155555965486354 2.7715999999999998e-08 1.817379418443826 2.7717e-08 1.7256487259691906 2.7718e-08 1.7447769065397172 2.7718999999999998e-08 1.7971012230622958 2.772e-08 1.7859930898670964 2.7721e-08 1.8331252856021722 2.7722e-08 1.798615775943317 2.7723e-08 1.8345723562870804 2.7724e-08 1.8130606397558569 2.7725e-08 1.7443716585857554 2.7726e-08 1.8286096327984078 2.7727e-08 1.7756966715872877 2.7728e-08 1.790662836745333 2.7729e-08 1.7786741006016262 2.773e-08 1.766637090566727 2.7731e-08 1.7843811955968403 2.7732e-08 1.805844617953225 2.7733e-08 1.80299812554707 2.7734e-08 1.738154443190128 2.7735e-08 1.8479404101481944 2.7736e-08 1.7919588081529387 2.7737e-08 1.8126484771702598 2.7738e-08 1.86306981497733 2.7739e-08 1.771403986869503 2.774e-08 1.756589374929213 2.7741e-08 1.8657716364921186 2.7741999999999998e-08 1.7413103613591008 2.7743e-08 1.8013096224161194 2.7744e-08 1.8229109128471983 2.7744999999999998e-08 1.690636880087774 2.7746e-08 1.7727904715421667 2.7747e-08 1.8189732189051993 2.7747999999999998e-08 1.8379222806180582 2.7749e-08 1.7171182793722628 2.775e-08 1.8297962661689786 2.7750999999999998e-08 1.7638516654572047 2.7752e-08 1.8483038011298323 2.7753e-08 1.8146335743601771 2.7753999999999998e-08 1.8680932339873404 2.7755e-08 1.85409188569593 2.7756e-08 1.8781525804945456 2.7756999999999998e-08 1.7680199675220305 2.7758e-08 1.7874481642719426 2.7759e-08 1.7920951985415747 2.776e-08 1.8107370511585463 2.7761e-08 1.774018256497428 2.7762e-08 1.8211103714166337 2.7763e-08 1.8238984108865215 2.7764e-08 1.809547403415399 2.7765e-08 1.838444438878501 2.7766e-08 1.8214280701497556 2.7767e-08 1.7450746388888048 2.7768e-08 1.8013348831611655 2.7769e-08 1.7987700440263286 2.777e-08 1.7882574919594025 2.7771e-08 1.8022165392497038 2.7772e-08 1.8323998375776591 2.7773e-08 1.7344793096134674 2.7774e-08 1.8509432316840617 2.7775e-08 1.7570408103815254 2.7776e-08 1.8665687947457115 2.7776999999999998e-08 1.7887529928916874 2.7778e-08 1.8080868860732877 2.7779e-08 1.8505880487468953 2.7779999999999998e-08 1.8350675995687686 2.7781e-08 1.7564264447560842 2.7782e-08 1.8204755591508914 2.7782999999999998e-08 1.7578985974017423 2.7784e-08 1.8724460532879428 2.7785e-08 1.7299755762620577 2.7785999999999998e-08 1.8225519608508394 2.7787e-08 1.7599156723128133 2.7788e-08 1.846564627644621 2.7788999999999998e-08 1.8040207762494782 2.779e-08 1.8390798088614613 2.7791e-08 1.786097330481783 2.7791999999999998e-08 1.7138559177055652 2.7793e-08 1.7324472516026221 2.7794e-08 1.7625443322027379 2.7795e-08 1.8340392931738738 2.7796e-08 1.7582370835369696 2.7797e-08 1.8508008269968264 2.7798e-08 1.8403174722664613 2.7799e-08 1.769653467681586 2.78e-08 1.7542495953884154 2.7801e-08 1.835856527096288 2.7802e-08 1.7774639293126082 2.7803e-08 1.7993065405150097 2.7804e-08 1.7882940010000639 2.7805e-08 1.8300805018276771 2.7806e-08 1.732815864449226 2.7807e-08 1.7193079757968126 2.7808e-08 1.8185482389528957 2.7809e-08 1.8297221833697799 2.781e-08 1.7065083447921188 2.7811e-08 1.7536763423679926 2.7811999999999998e-08 1.8100514309930824 2.7813e-08 1.7244578895566511 2.7814e-08 1.7738040700746232 2.7814999999999998e-08 1.7566530947205625 2.7816e-08 1.8287289450359612 2.7817e-08 1.7866577342882706 2.7817999999999998e-08 1.7750416288233557 2.7819e-08 1.7758805217344347 2.782e-08 1.8089816941394288 2.7820999999999998e-08 1.8115143136901404 2.7822e-08 1.752757089687602 2.7823e-08 1.7316368003972387 2.7823999999999998e-08 1.8958153643540725 2.7825e-08 1.766920750792783 2.7826e-08 1.8127282867134962 2.7826999999999998e-08 1.7453407639579561 2.7828e-08 1.700008990171164 2.7829e-08 1.7425949535526977 2.783e-08 1.8314898854820343 2.7831e-08 1.774078873696284 2.7832e-08 1.8254177920858834 2.7833e-08 1.7327059593308574 2.7834e-08 1.777793047299945 2.7835e-08 1.8056649596936187 2.7836e-08 1.7700349655135352 2.7837e-08 1.776059800232247 2.7838e-08 1.7782101898724874 2.7839e-08 1.7691107074017325 2.784e-08 1.7904640798832254 2.7841e-08 1.873317872873802 2.7842e-08 1.7590453447252141 2.7843e-08 1.712198196661833 2.7844e-08 1.8159343722168337 2.7845e-08 1.8408142775483243 2.7846e-08 1.888916759132938 2.7846999999999998e-08 1.7156613734164023 2.7848e-08 1.8048124812989201 2.7849e-08 1.817096085141423 2.7849999999999998e-08 1.848353879625439 2.7851e-08 1.7572764873675213 2.7852e-08 1.7001298149389523 2.7852999999999998e-08 1.7733301083743638 2.7854e-08 1.793232160364249 2.7855e-08 1.817227755778715 2.7855999999999998e-08 1.8272667677948748 2.7857e-08 1.7426919853935339 2.7858e-08 1.7878973690614728 2.7858999999999998e-08 1.8008610309887536 2.786e-08 1.7743208136480326 2.7861e-08 1.8101005072285783 2.7861999999999998e-08 1.7229997300197373 2.7863e-08 1.9027176997568171 2.7864e-08 1.7725155505918746 2.7865e-08 1.8560241915077111 2.7866e-08 1.8189402063161872 2.7867e-08 1.8399460245886854 2.7868e-08 1.7503133634779378 2.7869e-08 1.7837640076664898 2.787e-08 1.8590355662371 2.7871e-08 1.8409548329888246 2.7872e-08 1.7538911671961332 2.7873e-08 1.7744064837442401 2.7874e-08 1.7828062885726677 2.7875e-08 1.8033873517570869 2.7876e-08 1.8175144402653256 2.7877e-08 1.7971085797954904 2.7878e-08 1.8368425000061117 2.7879e-08 1.7876574996011516 2.788e-08 1.7713387740145725 2.7881e-08 1.753403736452982 2.7881999999999998e-08 1.758931713293725 2.7883e-08 1.7389586967290454 2.7884e-08 1.7326321330435304 2.7884999999999998e-08 1.8274763118787016 2.7886e-08 1.8292389727050136 2.7887e-08 1.7613631334311861 2.7887999999999998e-08 1.776010947712365 2.7889e-08 1.742183120008353 2.789e-08 1.759761320748281 2.7890999999999998e-08 1.8808422401133613 2.7892e-08 1.8502335484862098 2.7893e-08 1.841567384094272 2.7893999999999998e-08 1.8470198460011034 2.7895e-08 1.809903456826924 2.7896e-08 1.8583694584899506 2.7896999999999998e-08 1.7634532082795649 2.7898e-08 1.7664016353731606 2.7899e-08 1.8311923476527627 2.79e-08 1.794643744427495 2.7901e-08 1.7546457000908247 2.7902e-08 1.75122054248594 2.7903e-08 1.7725878340227563 2.7904e-08 1.7928910801022584 2.7905e-08 1.8010849932825947 2.7906e-08 1.792987683072121 2.7907e-08 1.8317633162460218 2.7908e-08 1.719325086511547 2.7909e-08 1.9249252715321439 2.791e-08 1.879523381088986 2.7911e-08 1.7971091274103124 2.7912e-08 1.8268831138980617 2.7913e-08 1.8337414474193758 2.7914e-08 1.8404733429973452 2.7915e-08 1.7975079144022412 2.7916e-08 1.8384284492054996 2.7916999999999998e-08 1.7124293955344385 2.7918e-08 1.784476781234572 2.7919e-08 1.7972214711976884 2.7919999999999998e-08 1.7760577484805886 2.7921e-08 1.809124738023791 2.7922e-08 1.806021945736204 2.7922999999999998e-08 1.7972585089114086 2.7924e-08 1.892800083172279 2.7925e-08 1.82932764292327 2.7925999999999998e-08 1.6650066890477524 2.7927e-08 1.9078900125748048 2.7928e-08 1.8089214524590755 2.7928999999999998e-08 1.8812681151892388 2.793e-08 1.8815294351718261 2.7931e-08 1.77792415892484 2.7931999999999998e-08 1.7649910515614318 2.7933e-08 1.8147670864691618 2.7934e-08 1.7890044781066272 2.7935e-08 1.8241113335103805 2.7936e-08 1.8123792410529318 2.7937e-08 1.7466354165969102 2.7938e-08 1.8130005647212106 2.7939e-08 1.8628414768509718 2.794e-08 1.8154326525952704 2.7941e-08 1.7843313228170443 2.7942e-08 1.7686784422023223 2.7943e-08 1.8373232959712749 2.7944e-08 1.8023568970381059 2.7945e-08 1.863178443663979 2.7946e-08 1.7719120552060337 2.7947e-08 1.76321905547671 2.7948e-08 1.7420722141234184 2.7949e-08 1.9051298425054346 2.795e-08 1.7315382716562502 2.7951e-08 1.827468407766476 2.7952e-08 1.7448975604763053 2.7953e-08 1.7601893561813227 2.7954e-08 1.7259754607138478 2.7954999999999998e-08 1.9128959147734936 2.7956e-08 1.837752832346756 2.7957e-08 1.8048137003095024 2.7957999999999998e-08 1.773329756129672 2.7959e-08 1.7339579441206592 2.796e-08 1.8299039738800644 2.7960999999999998e-08 1.8525711940733356 2.7962e-08 1.7947526879318763 2.7963e-08 1.8459358098460625 2.7963999999999998e-08 1.7786829554558163 2.7965e-08 1.5660473628146385 2.7966e-08 1.7492673644090875 2.7966999999999998e-08 1.8987227372771385 2.7968e-08 1.8321030457151064 2.7969e-08 1.8818979254487491 2.7969999999999998e-08 1.8409264595816908 2.7971e-08 1.8343086781198343 2.7972e-08 1.7778205893601804 2.7973e-08 1.7860029859220512 2.7974e-08 1.7717969272973266 2.7975e-08 1.7730367191569665 2.7976e-08 1.7863660795085794 2.7977e-08 1.8719601458751325 2.7978e-08 1.8573687414722588 2.7979e-08 1.8400148437925512 2.798e-08 1.8626808170018745 2.7981e-08 1.804862191708054 2.7982e-08 1.7289247112594208 2.7983e-08 1.8447032652519229 2.7984e-08 1.7528975370770745 2.7985e-08 1.743750412128919 2.7986e-08 1.806359357346776 2.7987e-08 1.8432505796859555 2.7988e-08 1.800253371733759 2.7989e-08 1.796389023902427 2.7989999999999998e-08 1.7645472202867447 2.7991e-08 1.7681643311600628 2.7992e-08 1.8998014282274969 2.7992999999999998e-08 1.8478210369089207 2.7994e-08 1.8948186711958965 2.7995e-08 1.7416145740039224 2.7995999999999998e-08 1.7560737913328088 2.7997e-08 1.7573307542310614 2.7998e-08 1.756276508576312 2.7998999999999998e-08 1.7833748743667357 2.8e-08 1.8302968847841505 2.8001e-08 1.7555401795627226 2.8001999999999998e-08 1.7644002229449391 2.8003e-08 1.891510121072928 2.8004e-08 1.8585397244874102 2.8004999999999998e-08 1.8692720259906839 2.8006e-08 1.7772473636891974 2.8007e-08 1.8118915536383537 2.8008e-08 1.8096782355731689 2.8009e-08 1.7490731187049369 2.801e-08 1.726783347274838 2.8011e-08 1.7850822949364735 2.8012e-08 1.8589965162475715 2.8013e-08 1.750225720774674 2.8014e-08 1.7550773240612043 2.8015e-08 1.7655255590089962 2.8016e-08 1.8581406165254226 2.8017e-08 1.8483502799508156 2.8018e-08 1.7811498481978632 2.8019e-08 1.7591667903329433 2.802e-08 1.8938740427733747 2.8021e-08 1.7859411613251122 2.8022e-08 1.7237854141356075 2.8023e-08 1.7775180097262318 2.8024e-08 1.7755908252009116 2.8024999999999998e-08 1.7842621932462608 2.8026e-08 1.8787655068978513 2.8027e-08 1.7458757310084354 2.8027999999999998e-08 1.8401831696725814 2.8029e-08 1.722584189624593 2.803e-08 1.7950210172782868 2.8030999999999998e-08 1.7714601842524607 2.8032e-08 1.7583547779036215 2.8033e-08 1.8008256314745212 2.8033999999999998e-08 1.8385861489127528 2.8035e-08 1.8170029546912425 2.8036e-08 1.824831620292037 2.8036999999999998e-08 1.7457028910594723 2.8038e-08 1.865239094947697 2.8039e-08 1.8458421041669806 2.8039999999999998e-08 1.890245300216988 2.8041e-08 1.8075176100688943 2.8042e-08 1.7660250084589333 2.8043e-08 1.7902490569935194 2.8044e-08 1.8473667755054541 2.8045e-08 1.8191627805327546 2.8046e-08 1.8186498796509285 2.8047e-08 1.8435631932999261 2.8048e-08 1.7307703820555072 2.8049e-08 1.7680788218966974 2.805e-08 1.8130216860740043 2.8051e-08 1.868275197497139 2.8052e-08 1.9397137382597744 2.8053e-08 1.810512723098084 2.8054e-08 1.7957005010144647 2.8055e-08 1.7785604234151882 2.8056e-08 1.7522354131658904 2.8057e-08 1.866330517977097 2.8058e-08 1.8349071139874997 2.8059e-08 1.735629750095832 2.8059999999999998e-08 1.8360454149779128 2.8061e-08 1.8277255324478088 2.8062e-08 1.7628696933227526 2.8062999999999998e-08 1.790778634973196 2.8064e-08 1.795166966795815 2.8065e-08 1.7898797535903062 2.8065999999999998e-08 1.774902311724171 2.8067e-08 1.742038915633591 2.8068e-08 1.7552144680731798 2.8068999999999998e-08 1.82451121922366 2.807e-08 1.8298479127621985 2.8071e-08 1.8406865173825993 2.8071999999999998e-08 1.8539552316985148 2.8073e-08 1.7442653445847507 2.8074e-08 1.804222889566211 2.8074999999999998e-08 1.8397236861182784 2.8076e-08 1.8429570135801705 2.8077e-08 1.8465173506990165 2.8078e-08 1.8031621381819247 2.8079e-08 1.7704940405238534 2.808e-08 1.7919870468608234 2.8081e-08 1.8026646034494724 2.8082e-08 1.8858453325576832 2.8083e-08 1.8101618251136848 2.8084e-08 1.7681308991901832 2.8085e-08 1.8524674754289328 2.8086e-08 1.8069391069165235 2.8087e-08 1.754795303298391 2.8088e-08 1.7923527414462777 2.8089e-08 1.8014674161306174 2.809e-08 1.7557783603763246 2.8091e-08 1.8282217831789973 2.8092e-08 1.7835847941485123 2.8093e-08 1.6872206618564618 2.8094e-08 1.7494954465954777 2.8094999999999998e-08 1.8593619107547816 2.8096e-08 1.857027047348166 2.8097e-08 1.7581403979000956 2.8097999999999998e-08 1.7817683818193275 2.8099e-08 1.824849316032452 2.81e-08 1.7706502110202913 2.8100999999999998e-08 1.85728767135202 2.8102e-08 1.7258151950173337 2.8103e-08 1.781524746393896 2.8103999999999998e-08 1.8029234727931989 2.8105e-08 1.7981933500741831 2.8106e-08 1.765245109039932 2.8106999999999998e-08 1.775126114450524 2.8108e-08 1.8121586149218603 2.8109e-08 1.7809387964380905 2.8109999999999998e-08 1.8865520729081766 2.8111e-08 1.7678651854062197 2.8112e-08 1.8188777727687964 2.8113e-08 1.776348603914207 2.8114e-08 1.768148733511312 2.8115e-08 1.8314988451838392 2.8116e-08 1.8123220926069674 2.8117e-08 1.7894032116703158 2.8118e-08 1.8930821784119363 2.8119e-08 1.8149267639255013 2.812e-08 1.7852680849947937 2.8121e-08 1.87823701405832 2.8122e-08 1.7001115336191757 2.8123e-08 1.807281323358845 2.8124e-08 1.7591322126739524 2.8125e-08 1.86799279740151 2.8126e-08 1.814337123959998 2.8127e-08 1.7831393620669709 2.8128e-08 1.8825377524490614 2.8129e-08 1.807076059389214 2.813e-08 1.7971174366176026 2.8131e-08 1.863796214034452 2.8132e-08 1.881495800457913 2.8132999999999998e-08 1.8079739822756171 2.8134e-08 1.720194117836444 2.8135e-08 1.7452320779529968 2.8135999999999998e-08 1.774618424361056 2.8137e-08 1.7135660968835265 2.8138e-08 1.7976654654235353 2.8138999999999998e-08 1.7687194632081753 2.814e-08 1.8162412495006082 2.8141e-08 1.7894562243030607 2.8141999999999998e-08 1.8239558546725967 2.8143e-08 1.7792543799832015 2.8144e-08 1.8276536878414524 2.8144999999999998e-08 1.7750644297605294 2.8146e-08 1.876346446333732 2.8147e-08 1.755273320364284 2.8147999999999998e-08 1.7474239358302142 2.8149e-08 1.7618925168818513 2.815e-08 1.7421575128423274 2.8151e-08 1.7696481687584504 2.8152e-08 1.9250730094076831 2.8153e-08 1.783882140652881 2.8154e-08 1.7754381993266632 2.8155e-08 1.8473469579474018 2.8156e-08 1.915798305987917 2.8157e-08 1.740864382459709 2.8158e-08 1.8751982238023923 2.8159e-08 1.7571380120428723 2.816e-08 1.843076886010441 2.8161e-08 1.7597048864767717 2.8162e-08 1.7955473266066222 2.8163e-08 1.8605765720992546 2.8164e-08 1.7758693983370977 2.8165e-08 1.832264193809979 2.8166e-08 1.776977872952646 2.8167e-08 1.8266818297162188 2.8167999999999998e-08 1.853618974455491 2.8169e-08 1.788470917045428 2.817e-08 1.7177151428200466 2.8170999999999998e-08 1.8229456892850922 2.8172e-08 1.7751916679698911 2.8173e-08 1.7478213279695296 2.8173999999999998e-08 1.8462332076965282 2.8175e-08 1.743410604424743 2.8176e-08 1.7168461615472905 2.8176999999999998e-08 1.829088091760077 2.8178e-08 1.8128171068602745 2.8179e-08 1.9265073584159782 2.8179999999999998e-08 1.8018242479036566 2.8181e-08 1.7723051236062202 2.8182e-08 1.8309656386424487 2.8182999999999998e-08 1.8062484362229094 2.8184e-08 1.8488972511657813 2.8185e-08 1.682322111577553 2.8186e-08 1.8230207451511982 2.8187e-08 1.7953695093052102 2.8188e-08 1.8706445155951323 2.8189e-08 1.7887147763414721 2.819e-08 1.8717453218689633 2.8191e-08 1.7405651355016936 2.8192e-08 1.8043050886389893 2.8193e-08 1.7686261221466435 2.8194e-08 1.7661086483516248 2.8195e-08 1.7979093224366784 2.8196e-08 1.7736655682037132 2.8197e-08 1.7515960594208753 2.8198e-08 1.8566122108734655 2.8199e-08 1.7647419120206393 2.82e-08 1.8432897297613033 2.8201e-08 1.748066314235629 2.8202e-08 1.7185240113101412 2.8202999999999998e-08 1.783034088986348 2.8204e-08 1.8218833633275051 2.8205e-08 1.796974256133286 2.8205999999999998e-08 1.743186216909182 2.8207e-08 1.8556729955146238 2.8208e-08 1.7977264092485128 2.8208999999999998e-08 1.7820506495253592 2.821e-08 1.9443979756191547 2.8211e-08 1.7940813657546066 2.8211999999999998e-08 1.7135247269944938 2.8213e-08 1.7913729587123 2.8214e-08 1.8382792866569535 2.8214999999999998e-08 1.7900388992607215 2.8216e-08 1.787896189611855 2.8217e-08 1.826834465216346 2.8217999999999998e-08 1.7912335849196677 2.8219e-08 1.8042010783570954 2.822e-08 1.7391403228715503 2.8221e-08 1.7304374471170914 2.8222e-08 1.746305436214426 2.8223e-08 1.778172946144283 2.8224e-08 1.8306958626803398 2.8225e-08 1.9081375701847627 2.8226e-08 1.8099878216873302 2.8227e-08 1.7235426030111767 2.8228e-08 1.9025882979817572 2.8229e-08 1.7213456561196152 2.823e-08 1.8360822475795178 2.8231e-08 1.8452752459499506 2.8232e-08 1.832927871214017 2.8233e-08 1.8483929034275453 2.8234e-08 1.8513035745930164 2.8235e-08 1.8238982671310762 2.8236e-08 1.758578391705437 2.8237e-08 1.749962953054876 2.8237999999999998e-08 1.7796325211201873 2.8239e-08 1.6585410491493535 2.824e-08 1.725718889650889 2.8240999999999998e-08 1.8420564852091894 2.8242e-08 1.7968139427430776 2.8243e-08 1.8034030136601655 2.8243999999999998e-08 1.8698438918922944 2.8245e-08 1.8487505479124455 2.8246e-08 1.8550237972327985 2.8246999999999998e-08 1.8379469744590748 2.8248e-08 1.7428220993341417 2.8249e-08 1.7815325561709152 2.8249999999999998e-08 1.739658827066757 2.8251e-08 1.7406453227277965 2.8252e-08 1.7501256522544566 2.8252999999999998e-08 1.8482825830374205 2.8254e-08 1.7075758250125803 2.8255e-08 1.9121434336259293 2.8256e-08 1.7988782171965174 2.8257e-08 1.7562381077605442 2.8258e-08 1.8527325148949785 2.8259e-08 1.7971102821791793 2.826e-08 1.8043131970394408 2.8261e-08 1.7401783257820687 2.8262e-08 1.7680340708538496 2.8263e-08 1.7672026872365332 2.8264e-08 1.7950965581960285 2.8265e-08 1.797056325842541 2.8266e-08 1.87557947310998 2.8267e-08 1.7720013166596829 2.8268e-08 1.7510783077635006 2.8269e-08 1.85612636038698 2.827e-08 1.7737438516519997 2.8271e-08 1.7970008356117728 2.8272e-08 1.8211835588758387 2.8272999999999998e-08 1.8088954561199555 2.8274e-08 1.8745098992652873 2.8275e-08 1.8474425592847672 2.8275999999999998e-08 1.7403218030597813 2.8277e-08 1.8008664352318238 2.8278e-08 1.8337411050060506 2.8278999999999998e-08 1.830956834331302 2.828e-08 1.6906177539599163 2.8281e-08 1.8452392430606734 2.8281999999999998e-08 1.9222542575142538 2.8283e-08 1.8942620383850475 2.8284e-08 1.8406422919219059 2.8284999999999998e-08 1.7171686602649683 2.8286e-08 1.757866616976706 2.8287e-08 1.7620548280025485 2.8287999999999998e-08 1.9100569336947582 2.8289e-08 1.74467776615668 2.829e-08 1.8498720950102463 2.8291e-08 1.7988744919420914 2.8292e-08 1.7284272443046744 2.8293e-08 1.8187503350471699 2.8294e-08 1.826756645492215 2.8295e-08 1.9129986870545794 2.8296e-08 1.8843712188178878 2.8297e-08 1.74182467884877 2.8298e-08 1.8015936233770442 2.8299e-08 1.7980712939539012 2.83e-08 1.6771985922664663 2.8301e-08 1.8960837763540455 2.8302e-08 1.7166704801231738 2.8303e-08 1.7594160018375637 2.8304e-08 1.8569112050971766 2.8305e-08 1.8248865574405244 2.8306e-08 1.8629523744357963 2.8307e-08 1.7539813599061023 2.8307999999999998e-08 1.7566654520279639 2.8309e-08 1.8415505721766432 2.831e-08 1.8242547904646949 2.8310999999999998e-08 1.7790877818021655 2.8312e-08 1.8306211930417557 2.8313e-08 1.8423759171158414 2.8313999999999998e-08 1.77807064792949 2.8315e-08 1.8250125481120207 2.8316e-08 1.7943051129131897 2.8316999999999998e-08 1.8116671718893376 2.8318e-08 1.7617989822186033 2.8319e-08 1.7830779930634542 2.8319999999999998e-08 1.7589294023089819 2.8321e-08 1.7900811398983696 2.8322e-08 1.7779471917379825 2.8322999999999998e-08 1.8123231004617966 2.8324e-08 1.6869617807497153 2.8325e-08 1.7580752233086245 2.8325999999999998e-08 1.8528382571870463 2.8327e-08 1.8850876516953665 2.8328e-08 1.7849948234443955 2.8329e-08 1.7461368718482784 2.833e-08 1.9046663521109952 2.8331e-08 1.84119115340652 2.8332e-08 1.824648134332671 2.8333e-08 1.8521113010926473 2.8334e-08 1.746503822219444 2.8335e-08 1.7685165475866549 2.8336e-08 1.83809643976387 2.8337e-08 1.7528275976059142 2.8338e-08 1.8512874617168193 2.8339e-08 1.743012339408716 2.834e-08 1.826442547575201 2.8341e-08 1.8182116777456103 2.8342e-08 1.84971740816764 2.8343e-08 1.7839282076254304 2.8344e-08 1.7032657242798386 2.8345e-08 1.8405192135021913 2.8345999999999998e-08 1.7254944002239423 2.8347e-08 1.7467678254305357 2.8348e-08 1.8347356853729768 2.8348999999999998e-08 1.7571615067534212 2.835e-08 1.7951445886295496 2.8351e-08 1.8154410417809073 2.8351999999999998e-08 1.9055217924148982 2.8353e-08 1.896361000097711 2.8354e-08 1.7514240035588928 2.8354999999999998e-08 1.7333150840943214 2.8356e-08 1.8260051911508752 2.8357e-08 1.7979998554487473 2.8357999999999998e-08 1.7945187959733457 2.8359e-08 1.7678419290625607 2.836e-08 1.7779945502009304 2.8360999999999998e-08 1.6904048056765761 2.8362e-08 1.6951090527895514 2.8363e-08 1.8883504757749405 2.8364e-08 1.7996908334562978 2.8365e-08 1.825626486157912 2.8366e-08 1.7306508427761131 2.8367e-08 1.852323864590325 2.8368e-08 1.6746940530160213 2.8369e-08 1.8362693634015377 2.837e-08 1.8103054565307095 2.8371e-08 1.7791606755816556 2.8372e-08 1.7603574014502634 2.8373e-08 1.8261994110866606 2.8374e-08 1.7858003494753307 2.8375e-08 1.8450544445561055 2.8376e-08 1.7895568798455408 2.8377e-08 1.8437542650276597 2.8378e-08 1.8250661814810643 2.8379e-08 1.8154112252993333 2.838e-08 1.834393920278174 2.8380999999999998e-08 1.7702918142097361 2.8382e-08 1.8046757887441718 2.8383e-08 1.7817549112185667 2.8383999999999998e-08 1.8071184242838256 2.8385e-08 1.7310091729291535 2.8386e-08 1.845151444951177 2.8386999999999998e-08 1.8889640311987623 2.8388e-08 1.7259892837754456 2.8389e-08 1.7579772725665868 2.8389999999999998e-08 1.7563818897982748 2.8391e-08 1.8239437638372602 2.8392e-08 1.6989049916769134 2.8392999999999998e-08 1.7931546191114658 2.8394e-08 1.7591491994896822 2.8395e-08 1.8268385675101155 2.8395999999999998e-08 1.842439482480194 2.8397e-08 1.8248500376846972 2.8398e-08 1.810505018216681 2.8399e-08 1.7721404584020908 2.84e-08 1.913622279903939 2.8401e-08 1.8109457047401478 2.8402e-08 1.7863989056776408 2.8403e-08 1.7617891949576765 2.8404e-08 1.777033951474178 2.8405e-08 1.850858089845314 2.8406e-08 1.6898997449540296 2.8407e-08 1.7304027306010807 2.8408e-08 1.8558123333696348 2.8409e-08 1.8065585148768453 2.841e-08 1.8042506406681027 2.8411e-08 1.8683652674526139 2.8412e-08 1.7770782561204015 2.8413e-08 1.8727318895130232 2.8414e-08 1.861527729689736 2.8415e-08 1.8013454554299517 2.8415999999999998e-08 1.7371147632123844 2.8417e-08 1.8019889670806437 2.8418e-08 1.7467232565221595 2.8418999999999998e-08 1.8421695909368305 2.842e-08 1.8145861091831421 2.8421e-08 1.7921827980231 2.8421999999999998e-08 1.8660438058616489 2.8423e-08 1.8461620363758242 2.8424e-08 1.8240637714585277 2.8424999999999998e-08 1.850243010205446 2.8426e-08 1.7989055883436587 2.8427e-08 1.7566196466112636 2.8427999999999998e-08 1.8230969927744276 2.8429e-08 1.8002913455841008 2.843e-08 1.8085227775867663 2.8430999999999998e-08 1.7801598217367676 2.8432e-08 1.7217083944062308 2.8433e-08 1.8495217398380785 2.8434e-08 1.687047313648795 2.8435e-08 1.8337484558130959 2.8436e-08 1.7772684053660568 2.8437e-08 1.7679623384241279 2.8438e-08 1.8364489703034859 2.8439e-08 1.7673072154319456 2.844e-08 1.8358396356852777 2.8441e-08 1.8190684896142224 2.8442e-08 1.8461418437283892 2.8443e-08 1.7600516679380673 2.8444e-08 1.7981962366502358 2.8445e-08 1.7841985648167125 2.8446e-08 1.7802730902105048 2.8447e-08 1.8472558644377988 2.8448e-08 1.7028795261215408 2.8449e-08 1.7860211432598048 2.845e-08 1.8615001497257697 2.8450999999999998e-08 1.7520276219123534 2.8452e-08 1.805852879996953 2.8453e-08 1.7803970711323462 2.8453999999999998e-08 1.8576726059013995 2.8455e-08 1.7472949272810359 2.8456e-08 1.7915051781980127 2.8456999999999998e-08 1.7916006891048581 2.8458e-08 1.7731635443915712 2.8459e-08 1.8528159327003817 2.8459999999999998e-08 1.8102723397681826 2.8461e-08 1.8083228445356223 2.8462e-08 1.7850511980452228 2.8462999999999998e-08 1.7365837540058742 2.8464e-08 1.7949724748233777 2.8465e-08 1.7454025652465737 2.8465999999999998e-08 1.72940171388521 2.8467e-08 1.8050836066767648 2.8468e-08 1.6940610773226814 2.8469e-08 1.7333953530205295 2.847e-08 1.8027495402465745 2.8471e-08 1.7328242728142333 2.8472e-08 1.7607201220823643 2.8473e-08 1.7709491620776543 2.8474e-08 1.861121942024483 2.8475e-08 1.7911290404746039 2.8476e-08 1.8141669437931967 2.8477e-08 1.7837453785125463 2.8478e-08 1.7987004330880114 2.8479e-08 1.7886078900308282 2.848e-08 1.692724196447878 2.8481e-08 1.7767493292055634 2.8482e-08 1.7580236518837853 2.8483e-08 1.7954909091808087 2.8484e-08 1.8321064134697644 2.8485e-08 1.7836672105603975 2.8485999999999998e-08 1.7556545165214819 2.8487e-08 1.7760902080172862 2.8488e-08 1.8161601540162633 2.8488999999999998e-08 1.7751826803044246 2.849e-08 1.8332182966551425 2.8491e-08 1.7901988635733865 2.8491999999999998e-08 1.8243118066880957 2.8493e-08 1.7972821060149744 2.8494e-08 1.8289031259220576 2.8494999999999998e-08 1.7563250625199236 2.8496e-08 1.8135361410825224 2.8497e-08 1.7502338846587229 2.8497999999999998e-08 1.8289818736150767 2.8499e-08 1.8707660900530725 2.85e-08 1.7200500065441013 2.8500999999999998e-08 1.7426461136347726 2.8502e-08 1.8134380979055351 2.8503e-08 1.8092969248543276 2.8504e-08 1.7912962355654933 2.8505e-08 1.7907760177733918 2.8506e-08 1.8971030744314485 2.8507e-08 1.772609951486812 2.8508e-08 1.7807846812227281 2.8509e-08 1.7300549100140088 2.851e-08 1.7889003932679028 2.8511e-08 1.8254964801112097 2.8512e-08 1.8463457825960554 2.8513e-08 1.8818666291506672 2.8514e-08 1.7787009502245945 2.8515e-08 1.7498635675524448 2.8516e-08 1.8230452756975914 2.8517e-08 1.712108684792915 2.8518e-08 1.7948163849313699 2.8519e-08 1.7499206022732112 2.852e-08 1.8383018488624754 2.8520999999999998e-08 1.803962740972398 2.8522e-08 1.8443093136520499 2.8523e-08 1.8311601053388222 2.8523999999999998e-08 1.8075878213860412 2.8525e-08 1.7346046693914459 2.8526e-08 1.7658679886777895 2.8526999999999998e-08 1.76331685355368 2.8528e-08 1.8063960361468578 2.8529e-08 1.7845040035368944 2.8529999999999998e-08 1.8386843140040106 2.8531e-08 1.8652943287970223 2.8532e-08 1.8241634844944674 2.8532999999999998e-08 1.7948398711791231 2.8534e-08 1.7884130581712596 2.8535e-08 1.780902228898142 2.8535999999999998e-08 1.7648437745248673 2.8537e-08 1.8620135374834792 2.8538e-08 1.761915672857431 2.8538999999999998e-08 1.7351891169957743 2.854e-08 1.7425226708600026 2.8541e-08 1.8282980451289415 2.8542e-08 1.8243438853143403 2.8543e-08 1.8559580428381397 2.8544e-08 1.7469509748980965 2.8545e-08 1.8591731284087585 2.8546e-08 1.7080051276406067 2.8547e-08 1.8235730024434296 2.8548e-08 1.7241875129568054 2.8549e-08 1.7315369284957323 2.855e-08 1.718020734072231 2.8551e-08 1.8061754092125943 2.8552e-08 1.8965083337303046 2.8553e-08 1.8806083152024307 2.8554e-08 1.8026610595327635 2.8555e-08 1.8015124986588433 2.8556e-08 1.8613964181797924 2.8557e-08 1.8612537214778127 2.8558e-08 1.8447637610860934 2.8558999999999998e-08 1.743587539497304 2.856e-08 1.7249912886027539 2.8561e-08 1.875590737661878 2.8561999999999998e-08 1.8211243685763523 2.8563e-08 1.9062954371117589 2.8564e-08 1.8340138717457684 2.8564999999999998e-08 1.8448366256013855 2.8566e-08 1.7170957701990859 2.8567e-08 1.8055917743509209 2.8567999999999998e-08 1.7449882905820453 2.8569e-08 1.7818583311951885 2.857e-08 1.7817700059710115 2.8570999999999998e-08 1.8152443039768413 2.8572e-08 1.8062734376223957 2.8573e-08 1.7816004756373112 2.8573999999999998e-08 1.7778328352852193 2.8575e-08 1.8239609336428593 2.8576e-08 1.8261099679654136 2.8577e-08 1.765480104815045 2.8578e-08 1.7796029388027823 2.8579e-08 1.8234070098316373 2.858e-08 1.8747006330477833 2.8581e-08 1.868131049516601 2.8582e-08 1.8923821568732402 2.8583e-08 1.7473336727092348 2.8584e-08 1.7466526099835293 2.8585e-08 1.8257990386825398 2.8586e-08 1.8461237440083347 2.8587e-08 1.8032638512138548 2.8588e-08 1.8093441488763014 2.8589e-08 1.7624736888244943 2.859e-08 1.80215379526812 2.8591e-08 1.753030923781181 2.8592e-08 1.8094137087220734 2.8593e-08 1.8233815833706373 2.8593999999999998e-08 1.7688581388806646 2.8595e-08 1.709106897895904 2.8596e-08 1.8425481493171647 2.8596999999999998e-08 1.7277504684599578 2.8598e-08 1.7832166967590022 2.8599e-08 1.8504343016498734 2.8599999999999998e-08 1.8859130762079588 2.8601e-08 1.7129560300002167 2.8602e-08 1.7976175717655443 2.8602999999999998e-08 1.8025671916437849 2.8604e-08 1.881053388213537 2.8605e-08 1.8141768539782888 2.8605999999999998e-08 1.8252077133423412 2.8607e-08 1.7925734898807193 2.8608e-08 1.817317670699417 2.8608999999999998e-08 1.8453239877028405 2.861e-08 1.7616992609490632 2.8611e-08 1.8307668477168972 2.8612e-08 1.8605431090304148 2.8613e-08 1.8145425698678534 2.8614e-08 1.8173317338228083 2.8615e-08 1.7352264348891127 2.8616e-08 1.7959413363483288 2.8617e-08 1.8427913422982405 2.8618e-08 1.7201777659294037 2.8619e-08 1.8153592794498694 2.862e-08 1.760188247188514 2.8621e-08 1.7996443470021943 2.8622e-08 1.780340805424636 2.8623e-08 1.7616721783402358 2.8624e-08 1.7958591412483518 2.8625e-08 1.7816664806104163 2.8626e-08 1.7992104665594575 2.8627e-08 1.8730139560630155 2.8628e-08 1.7925454137135322 2.8628999999999998e-08 1.8593775833889354 2.863e-08 1.7790794618889392 2.8631e-08 1.8082793686054266 2.8631999999999998e-08 1.7144080055800917 2.8633e-08 1.8307052831753792 2.8634e-08 1.794819990188283 2.8634999999999998e-08 1.9110809848269088 2.8636e-08 1.804605482303951 2.8637e-08 1.7047704454231585 2.8637999999999998e-08 1.6720042961784076 2.8639e-08 1.8207939124970647 2.864e-08 1.7993708666132762 2.8640999999999998e-08 1.7784093604281441 2.8642e-08 1.7253124462600629 2.8643e-08 1.780075749191172 2.8643999999999998e-08 1.7621994257578706 2.8645e-08 1.694919816586116 2.8646e-08 1.7827504263699667 2.8647e-08 1.8350213241640385 2.8648e-08 1.77857466227677 2.8649e-08 1.7911483093192955 2.865e-08 1.744568672072155 2.8651e-08 1.7788269649082562 2.8652e-08 1.8641674978684097 2.8653e-08 1.8969990248433855 2.8654e-08 1.7345845158536992 2.8655e-08 1.8323769352170658 2.8656e-08 1.7179357344228974 2.8657e-08 1.7731726753998827 2.8658e-08 1.8036336737749181 2.8659e-08 1.7847109115999373 2.866e-08 1.7645604289657542 2.8661e-08 1.8183952638231238 2.8662e-08 1.853766998586076 2.8663e-08 1.7324102556816774 2.8663999999999998e-08 1.8085878907657875 2.8665e-08 1.7567723939140911 2.8666e-08 1.8399472537125694 2.8666999999999998e-08 1.8462666171339372 2.8668e-08 1.7786516219142485 2.8669e-08 1.938154195375831 2.8669999999999998e-08 1.8232739798958817 2.8671e-08 1.7977424941707305 2.8672e-08 1.7440089828112153 2.8672999999999998e-08 1.7418826153516986 2.8674e-08 1.7047194603873248 2.8675e-08 1.9070149351339611 2.8675999999999998e-08 1.6437391449734664 2.8677e-08 1.8581856068727893 2.8678e-08 1.7129202931308707 2.8678999999999998e-08 1.7716544726894499 2.868e-08 1.7034977657860666 2.8681e-08 1.8655562462532298 2.8682e-08 1.7911645540402654 2.8683e-08 1.7222509807139645 2.8684e-08 1.8397112947467493 2.8685e-08 1.7313607417865178 2.8686e-08 1.8121866672421842 2.8687e-08 1.7582569478363548 2.8688e-08 1.809911276449652 2.8689e-08 1.7662905345230417 2.869e-08 1.7221984686858458 2.8691e-08 1.799693191663274 2.8692e-08 1.7741636808410186 2.8693e-08 1.8232356362870765 2.8694e-08 1.8174674671196431 2.8695e-08 1.8472297150173935 2.8696e-08 1.7129689141999085 2.8697e-08 1.7677248705662998 2.8698e-08 1.8741400972370605 2.8698999999999998e-08 1.8368330375347943 2.87e-08 1.8928873148301442 2.8701e-08 1.8233562476110543 2.8701999999999998e-08 1.8186604136123736 2.8703e-08 1.7997591456546504 2.8704e-08 1.8564593710613355 2.8704999999999998e-08 1.8485615752277915 2.8706e-08 1.7737392206242004 2.8707e-08 1.7518178582454853 2.8707999999999998e-08 1.830156190031809 2.8709e-08 1.8356168397065862 2.871e-08 1.8386660454998818 2.8710999999999998e-08 1.7994013314237312 2.8712e-08 1.849744639282035 2.8713e-08 1.8418236592546757 2.8713999999999998e-08 1.8619467153587974 2.8715e-08 1.8166416091188533 2.8716e-08 1.8274122514128042 2.8716999999999998e-08 1.783344614450072 2.8718e-08 1.822076409821105 2.8719e-08 1.7718975930482284 2.872e-08 1.8516504611932532 2.8721e-08 1.766300317312039 2.8722e-08 1.9151729478504687 2.8723e-08 1.8552051157885638 2.8724e-08 1.842826171732335 2.8725e-08 1.9011582925869412 2.8726e-08 1.7747498027016726 2.8727e-08 1.915090550923844 2.8728e-08 1.7699621515394572 2.8729e-08 1.7834808840563328 2.873e-08 1.831022520707887 2.8731e-08 1.7353216281031771 2.8732e-08 1.7479545305095499 2.8733e-08 1.8863788682636915 2.8734e-08 1.8014224854800165 2.8735e-08 1.7624154072364184 2.8736e-08 1.7834946155868059 2.8736999999999998e-08 1.8175553885648628 2.8738e-08 1.7445140205371799 2.8739e-08 1.8657767449130076 2.8739999999999998e-08 1.8438180162012818 2.8741e-08 1.8494486969697492 2.8742e-08 1.7637187499682212 2.8742999999999998e-08 1.78032757906499 2.8744e-08 1.7927509996689484 2.8745e-08 1.8786105397931208 2.8745999999999998e-08 1.756203357825045 2.8747e-08 1.6593176270425873 2.8748e-08 1.8697024386804686 2.8748999999999998e-08 1.8575167101836112 2.875e-08 1.794936452336404 2.8751e-08 1.7967715888943272 2.8751999999999998e-08 1.7830675476747626 2.8753e-08 1.8395087766370295 2.8754e-08 1.781054396392546 2.8755e-08 1.8394244500496144 2.8756e-08 1.822730096113019 2.8757e-08 1.7572489218875493 2.8758e-08 1.7604154680782393 2.8759e-08 1.8863035819670144 2.876e-08 1.7934623629072193 2.8761e-08 1.869463931555371 2.8762e-08 1.7774519206247401 2.8763e-08 1.7826546777095809 2.8764e-08 1.7313191072645244 2.8765e-08 1.8996782943315134 2.8766e-08 1.7855778391585875 2.8767e-08 1.8343985983149291 2.8768e-08 1.76789798796239 2.8769e-08 1.7549398871554447 2.877e-08 1.8477367436694498 2.8771e-08 1.7775510370872432 2.8771999999999998e-08 1.8243917484331 2.8773e-08 1.8130972170179218 2.8774e-08 1.7895704848545542 2.8774999999999998e-08 1.8582795896233109 2.8776e-08 1.7544693005458594 2.8777e-08 1.7764616890316738 2.8777999999999998e-08 1.7740129910927038 2.8779e-08 1.6736547315507555 2.878e-08 1.775565523587564 2.8780999999999998e-08 1.8554077221244205 2.8782e-08 1.767809100762448 2.8783e-08 1.796773414725416 2.8783999999999998e-08 1.831900439896259 2.8785e-08 1.8204946484207776 2.8786e-08 1.898374683642649 2.8786999999999998e-08 1.7794347693631996 2.8788e-08 1.8303440754760958 2.8789e-08 1.7856703413269723 2.879e-08 1.6988515677297404 2.8791e-08 1.7452994324830895 2.8792e-08 1.757009212773288 2.8793e-08 1.7689100273955651 2.8794e-08 1.791270694903944 2.8795e-08 1.8140458441877458 2.8796e-08 1.8222249419342185 2.8797e-08 1.8013572962837288 2.8798e-08 1.8139051723403887 2.8799e-08 1.7041889722481982 2.88e-08 1.7853961710140913 2.8801e-08 1.7106645016850652 2.8802e-08 1.8313636385181804 2.8803e-08 1.6813136730647968 2.8804e-08 1.698720260901123 2.8805e-08 1.7862743357376283 2.8806e-08 1.8088626868296633 2.8806999999999998e-08 1.7939275918845152 2.8808e-08 1.859586382121781 2.8809e-08 1.7146381943360463 2.8809999999999998e-08 1.836848265151906 2.8811e-08 1.8854435637968212 2.8812e-08 1.793234699628246 2.8812999999999998e-08 1.825411086555609 2.8814e-08 1.7364515892314099 2.8815e-08 1.7845891927991704 2.8815999999999998e-08 1.823884250407876 2.8817e-08 1.781622089679657 2.8818e-08 1.8193410151821068 2.8818999999999998e-08 1.7599107505210134 2.882e-08 1.8073360702454466 2.8821e-08 1.7732705541478682 2.8821999999999998e-08 1.8500500641480402 2.8823e-08 1.7898819189359274 2.8824e-08 1.7700123897134519 2.8825e-08 1.7722977920127374 2.8826e-08 1.7269474546378865 2.8827e-08 1.710209567627911 2.8828e-08 1.820865110825418 2.8829e-08 1.7788439724973635 2.883e-08 1.7835756620809493 2.8831e-08 1.813363757476512 2.8832e-08 1.8331260568658019 2.8833e-08 1.8328956522161306 2.8834e-08 1.8216493194407544 2.8835e-08 1.8322892064622163 2.8836e-08 1.7671845540974696 2.8837e-08 1.906281754569649 2.8838e-08 1.8175331867863858 2.8839e-08 1.7606335585885002 2.884e-08 1.7643373287265236 2.8841e-08 1.8259461262478256 2.8841999999999998e-08 1.7831929829611672 2.8843e-08 1.8258892456655424 2.8844e-08 1.8038735284125178 2.8844999999999998e-08 1.8843324382447468 2.8846e-08 1.7740973853533841 2.8847e-08 1.8066595176329083 2.8847999999999998e-08 1.7903217194807757 2.8849e-08 1.73243205841633 2.885e-08 1.7928590788189027 2.8850999999999998e-08 1.7488717666899098 2.8852e-08 1.7939355477185215 2.8853e-08 1.732778186674039 2.8853999999999998e-08 1.8405139725295576 2.8855e-08 1.80903134156791 2.8856e-08 1.850092486888106 2.8856999999999998e-08 1.8391337779127863 2.8858e-08 1.78427515387099 2.8859e-08 1.7346570963687307 2.886e-08 1.780502897983538 2.8861e-08 1.7683370651345156 2.8862e-08 1.814216211805891 2.8863e-08 1.7942247572799948 2.8864e-08 1.7142936735093617 2.8865e-08 1.8425057764900452 2.8866e-08 1.7416391269540372 2.8867e-08 1.7774398975137364 2.8868e-08 1.8441368727224883 2.8869e-08 1.839789121344808 2.887e-08 1.7987046975252392 2.8871e-08 1.7776454485206288 2.8872e-08 1.8196825977459594 2.8873e-08 1.7757762089513365 2.8874e-08 1.8969230583393983 2.8875e-08 1.870489137206703 2.8876e-08 1.7936842979757284 2.8876999999999998e-08 1.8189924125226398 2.8878e-08 1.8028294517392582 2.8879e-08 1.7600803535464855 2.8879999999999998e-08 1.7812811141832177 2.8881e-08 1.8161034145482828 2.8882e-08 1.9302879151033039 2.8882999999999998e-08 1.777870397141388 2.8884e-08 1.766724003022995 2.8885e-08 1.8502875393642213 2.8885999999999998e-08 1.8254939212566392 2.8887e-08 1.8534207938067206 2.8888e-08 1.8284339475941542 2.8888999999999998e-08 1.8725327611524183 2.889e-08 1.8180545904487517 2.8891e-08 1.7826939510574813 2.8891999999999998e-08 1.750060739252483 2.8893e-08 1.8574360501714593 2.8894e-08 1.743831965850496 2.8894999999999998e-08 1.7810982035811633 2.8896e-08 1.8212675100291191 2.8897e-08 1.7848483570091036 2.8898e-08 1.8415559142379563 2.8899e-08 1.8828640735870874 2.89e-08 1.8624768957748856 2.8901e-08 1.8373355968772453 2.8902e-08 1.8818429121275275 2.8903e-08 1.839370157591903 2.8904e-08 1.7508252533232498 2.8905e-08 1.7782041477053923 2.8906e-08 1.7816779794331246 2.8907e-08 1.819460283193255 2.8908e-08 1.8260613838256132 2.8909e-08 1.8409769905676538 2.891e-08 1.7647204324819108 2.8911e-08 1.789502569804698 2.8911999999999998e-08 1.8335659808465505 2.8913e-08 1.790966924246476 2.8914e-08 1.8789776222097057 2.8914999999999998e-08 1.7502871440400412 2.8916e-08 1.8056372794092221 2.8917e-08 1.888773312383052 2.8917999999999998e-08 1.7724582031481806 2.8919e-08 1.678418284443431 2.892e-08 1.856707213260861 2.8920999999999998e-08 1.826430743057432 2.8922e-08 1.8375462181599043 2.8923e-08 1.7503864216889904 2.8923999999999998e-08 1.7855323671577084 2.8925e-08 1.854122923064139 2.8926e-08 1.8180692680879043 2.8926999999999998e-08 1.8020720963435926 2.8928e-08 1.7890318051892495 2.8929e-08 1.837353645253144 2.8929999999999998e-08 1.8264643271017742 2.8931e-08 1.7566669601108524 2.8932e-08 1.7577953368250534 2.8933e-08 1.7947624696828026 2.8934e-08 1.8433046948913658 2.8935e-08 1.8166331559583353 2.8936e-08 1.8321432979852657 2.8937e-08 1.8494130418036485 2.8938e-08 1.7968644021446754 2.8939e-08 1.8327532830685909 2.894e-08 1.7273172208907772 2.8941e-08 1.8457672785696446 2.8942e-08 1.811161536479085 2.8943e-08 1.8130535875906864 2.8944e-08 1.8079941374528437 2.8945e-08 1.7612330361121862 2.8946e-08 1.7975277869488435 2.8947e-08 1.8274763401718745 2.8948e-08 1.8709467080368367 2.8949e-08 1.915686749923681 2.8949999999999998e-08 1.7962844668384983 2.8951e-08 1.799497251071712 2.8952e-08 1.8016162004127705 2.8952999999999998e-08 1.7539695309288388 2.8954e-08 1.859487153675619 2.8955e-08 1.739529794212233 2.8955999999999998e-08 1.7067314508695046 2.8957e-08 1.7476816129945416 2.8958e-08 1.8082329581626395 2.8958999999999998e-08 1.8020383443930634 2.896e-08 1.8655702189590313 2.8961e-08 1.7264959694989463 2.8961999999999998e-08 1.821334934493089 2.8963e-08 1.8388316476643924 2.8964e-08 1.8165589148631083 2.8964999999999998e-08 1.8864131598243992 2.8966e-08 1.7499935367899078 2.8967e-08 1.896891453779034 2.8968e-08 1.807089473001679 2.8969e-08 1.8556641087456525 2.897e-08 1.8105066901084526 2.8971e-08 1.868956120589765 2.8972e-08 1.7054113002539002 2.8973e-08 1.7956227842319543 2.8974e-08 1.7635715093171718 2.8975e-08 1.7843252181841631 2.8976e-08 1.8691130315878934 2.8977e-08 1.891692917703585 2.8978e-08 1.9179008919443847 2.8979e-08 1.8246017650032775 2.898e-08 1.7781902172786348 2.8981e-08 1.7369786596353611 2.8982e-08 1.8030608071978522 2.8983e-08 1.8775525606139678 2.8984e-08 1.791907941278384 2.8984999999999998e-08 1.8358077919336662 2.8986e-08 1.8372125159858832 2.8987e-08 1.883745399314271 2.8987999999999998e-08 1.7436068940268017 2.8989e-08 1.788812349667216 2.899e-08 1.8653288224232356 2.8990999999999998e-08 1.8011097917093026 2.8992e-08 1.8435523374257643 2.8993e-08 1.7501502913961278 2.8993999999999998e-08 1.7684796649302115 2.8995e-08 1.8425423884686887 2.8996e-08 1.7053802044996602 2.8996999999999998e-08 1.8139033403219 2.8998e-08 1.8623691355044407 2.8999e-08 1.7433067494070182 2.8999999999999998e-08 1.8074158088725272 2.9001e-08 1.8088389483748935 2.9002e-08 1.88696657572819 2.9003e-08 1.8705042567102295 2.9004e-08 1.8574842487052898 2.9005e-08 1.907466082456648 2.9006e-08 1.7961738526630364 2.9007e-08 1.7436156181031206 2.9008e-08 1.8672704886901923 2.9009e-08 1.7970036679316224 2.901e-08 1.8013084390755472 2.9011e-08 1.7970183498348218 2.9012e-08 1.7957712049796353 2.9013e-08 1.7774043749275499 2.9014e-08 1.796156227328703 2.9015e-08 1.8665617949420954 2.9016e-08 1.772421862110872 2.9017e-08 1.8106930465909097 2.9018e-08 1.7914281834594414 2.9019e-08 1.7760027511612866 2.9019999999999998e-08 1.7557794653026648 2.9021e-08 1.7929803079512399 2.9022e-08 1.717717797199326 2.9022999999999998e-08 1.7963830804614793 2.9024e-08 1.8333124371011909 2.9025e-08 1.8175355317631174 2.9025999999999998e-08 1.7956400983900285 2.9027e-08 1.7275528992029465 2.9028e-08 1.7729870582048115 2.9028999999999998e-08 1.7636294324709838 2.903e-08 1.7087674114519842 2.9031e-08 1.8297452711544242 2.9031999999999998e-08 1.83515467678378 2.9033e-08 1.8558647853911718 2.9034e-08 1.8567163140580454 2.9034999999999998e-08 1.7892474512712646 2.9036e-08 1.7957944051810646 2.9037e-08 1.8729525039263126 2.9038e-08 1.7751679458348704 2.9039e-08 1.879987733122258 2.904e-08 1.8381433692865656 2.9041e-08 1.8473164200111842 2.9042e-08 1.8928419689661407 2.9043e-08 1.7751302205003254 2.9044e-08 1.8163670223979076 2.9045e-08 1.8086078301143202 2.9046e-08 1.7390139383570618 2.9047e-08 1.8546431334423603 2.9048e-08 1.7808261093889675 2.9049e-08 1.834313115727035 2.905e-08 1.7539735468248263 2.9051e-08 1.8656188208173383 2.9052e-08 1.7344532721741568 2.9053e-08 1.798771365538526 2.9054e-08 1.722668101693482 2.9054999999999998e-08 1.8381780031228554 2.9056e-08 1.7429460580575307 2.9057e-08 1.890327886137929 2.9057999999999998e-08 1.7946528431020947 2.9059e-08 1.7066824566756016 2.906e-08 1.7990215223559307 2.9060999999999998e-08 1.8086701232812916 2.9062e-08 1.7188403210391947 2.9063e-08 1.7179348509344332 2.9063999999999998e-08 1.8466145519517274 2.9065e-08 1.7651640366680579 2.9066e-08 1.7693706824528441 2.9066999999999998e-08 1.7020849200190722 2.9068e-08 1.8630381442112238 2.9069e-08 1.7377479746353317 2.9069999999999998e-08 1.7649615479590428 2.9071e-08 1.8461937456486084 2.9072e-08 1.7805985061987788 2.9073e-08 1.840121927344686 2.9074e-08 1.7362450378236616 2.9075e-08 1.85761719204881 2.9076e-08 1.8050046592285751 2.9077e-08 1.7894441070337321 2.9078e-08 1.7550026452137961 2.9079e-08 1.7382545514061878 2.908e-08 1.796026263290256 2.9081e-08 1.834138907435891 2.9082e-08 1.7415316777689063 2.9083e-08 1.8871001385647288 2.9084e-08 1.7503670553143171 2.9085e-08 1.7413418158664555 2.9086e-08 1.8191876399460416 2.9087e-08 1.8079304940876855 2.9088e-08 1.7542015624687626 2.9089e-08 1.8556462917768966 2.9089999999999998e-08 1.783116511028164 2.9091e-08 1.7816687284794466 2.9092e-08 1.8199966842806268 2.9092999999999998e-08 1.8576132949183812 2.9094e-08 1.7947555579433123 2.9095e-08 1.824713436137788 2.9095999999999998e-08 1.7078369305234533 2.9097e-08 1.7480424079858825 2.9098e-08 1.8485441107004226 2.9098999999999998e-08 1.7461494058937639 2.91e-08 1.829974465761175 2.9101e-08 1.8347628091631552 2.9101999999999998e-08 1.8484957226099694 2.9103e-08 1.8289797171165434 2.9104e-08 1.8096123484106892 2.9104999999999998e-08 1.781303612857525 2.9106e-08 1.8056481585092297 2.9107e-08 1.8702994855037196 2.9107999999999998e-08 1.8132074013480466 2.9109e-08 1.7689233147197216 2.911e-08 1.7718966580531217 2.9111e-08 1.8484143521413727 2.9112e-08 1.7132350185669303 2.9113e-08 1.8283460616903562 2.9114e-08 1.801047218826696 2.9115e-08 1.8475097719520657 2.9116e-08 1.8538494304108175 2.9117e-08 1.9241224255993272 2.9118e-08 1.7760821002143883 2.9119e-08 1.807262476154442 2.912e-08 1.8817988175121112 2.9121e-08 1.8432578292748922 2.9122e-08 1.8100120601155494 2.9123e-08 1.7563873324201642 2.9124e-08 1.8229149384183616 2.9125e-08 1.7942347792599194 2.9126e-08 1.8389325683053963 2.9127e-08 1.7896200930937332 2.9127999999999998e-08 1.7731317075705815 2.9129e-08 1.8704701513085935 2.913e-08 1.6995999241822057 2.9130999999999998e-08 1.776556027084033 2.9132e-08 1.7168947707307685 2.9133e-08 1.8510867412060945 2.9133999999999998e-08 1.667938600532978 2.9135e-08 1.7932359147937014 2.9136e-08 1.767262924058762 2.9136999999999998e-08 1.7832645169299075 2.9138e-08 1.7999079420856268 2.9139e-08 1.8863282770671959 2.9139999999999998e-08 1.8550510132314726 2.9141e-08 1.824027445225264 2.9142e-08 1.7546103072797152 2.9142999999999998e-08 1.814802290550933 2.9144e-08 1.8247435913665289 2.9145e-08 1.7969968202239692 2.9146e-08 1.8299285610328613 2.9147e-08 1.8241642015669024 2.9148e-08 1.84342769384166 2.9149e-08 1.8586526919815833 2.915e-08 1.8009056435123942 2.9151e-08 1.747666989526384 2.9152e-08 1.7799331720995828 2.9153e-08 1.733358969245345 2.9154e-08 1.743659993841712 2.9155e-08 1.769387045510887 2.9156e-08 1.7883930388095814 2.9157e-08 1.8438045484598755 2.9158e-08 1.8335726637678758 2.9159e-08 1.837169779409189 2.916e-08 1.8324017697909918 2.9161e-08 1.8086034307579892 2.9162e-08 1.797578170437514 2.9162999999999998e-08 1.8364696907218148 2.9164e-08 1.7849607023006635 2.9165e-08 1.774937338934589 2.9165999999999998e-08 1.8865964062412222 2.9167e-08 1.7622977936621276 2.9168e-08 1.8370991197469126 2.9168999999999998e-08 1.8377073143828297 2.917e-08 1.828178979288704 2.9171e-08 1.9128168117861222 2.9171999999999998e-08 1.8061649761023348 2.9173e-08 1.8096531561610858 2.9174e-08 1.855752771467023 2.9174999999999998e-08 1.8081849192313502 2.9176e-08 1.8147659501042304 2.9177e-08 1.8021098863623388 2.9177999999999998e-08 1.8043702613920471 2.9179e-08 1.8319858712807666 2.918e-08 1.9066358255594762 2.9181e-08 1.7814593123935551 2.9182e-08 1.8442695221660317 2.9183e-08 1.8020531115610976 2.9184e-08 1.8320014045749864 2.9185e-08 1.7835540713381224 2.9186e-08 1.820961395650497 2.9187e-08 1.8290808911165959 2.9188e-08 1.8624125592869096 2.9189e-08 1.8375022359729525 2.919e-08 1.8394888229531177 2.9191e-08 1.8812589852961745 2.9192e-08 1.7376892957119567 2.9193e-08 1.8267148730796494 2.9194e-08 1.8329068683057257 2.9195e-08 1.7162200850385958 2.9196e-08 1.800301391581242 2.9197e-08 1.7522632862709495 2.9197999999999998e-08 1.793027652506084 2.9199e-08 1.7829293274092137 2.92e-08 1.8217894651312334 2.9200999999999998e-08 1.7980854586604158 2.9202e-08 1.7814861386230023 2.9203e-08 1.8150430371126096 2.9203999999999998e-08 1.7849260014025095 2.9205e-08 1.8539993731549211 2.9206e-08 1.806740535666919 2.9206999999999998e-08 1.830663422152013 2.9208e-08 1.783236216403189 2.9209e-08 1.8027608060845892 2.9209999999999998e-08 1.8382762962289798 2.9211e-08 1.764208022032697 2.9212e-08 1.7387888896149584 2.9212999999999998e-08 1.7670286194762563 2.9214e-08 1.8746434569143617 2.9215e-08 1.831965063315539 2.9216e-08 1.7938413211107767 2.9217e-08 1.7838724551450627 2.9218e-08 1.8162778221188598 2.9219e-08 1.7258774036244813 2.922e-08 1.7839553955525138 2.9221e-08 1.81217970788412 2.9222e-08 1.8262857376533883 2.9223e-08 1.8602751364537453 2.9224e-08 1.7141414083984658 2.9225e-08 1.79075187304 2.9226e-08 1.7627587178541309 2.9227e-08 1.7445812235800906 2.9228e-08 1.8447996844168415 2.9229e-08 1.7632941173631806 2.923e-08 1.7176105734243912 2.9231e-08 1.7752064856628849 2.9232e-08 1.8161790327051097 2.9232999999999998e-08 1.7884275938425536 2.9234e-08 1.7411120180125246 2.9235e-08 1.744728984571432 2.9235999999999998e-08 1.8817384997697473 2.9237e-08 1.7901368734845047 2.9238e-08 1.8899347045744324 2.9238999999999998e-08 1.7731989200448932 2.924e-08 1.7642582500468103 2.9241e-08 1.7503272427730043 2.9241999999999998e-08 1.8310550106929269 2.9243e-08 1.8162710659152446 2.9244e-08 1.7880385085845896 2.9244999999999998e-08 1.8741591610683348 2.9246e-08 1.8501577730087801 2.9247e-08 1.8252422305383564 2.9247999999999998e-08 1.830660602002993 2.9249e-08 1.857558765522386 2.925e-08 1.8013474730250512 2.9251e-08 1.8505832651632779 2.9252e-08 1.8738173876941067 2.9253e-08 1.763784620692138 2.9254e-08 1.825702816150961 2.9255e-08 1.7836821435761516 2.9256e-08 1.8618212513189996 2.9257e-08 1.8828833123366073 2.9258e-08 1.8172317243681633 2.9259e-08 1.8073901670189962 2.926e-08 1.768638183645222 2.9261e-08 1.726486462247631 2.9262e-08 1.7844107975012111 2.9263e-08 1.9052547270470201 2.9264e-08 1.8117897121588555 2.9265e-08 1.8336775519852475 2.9266e-08 1.8473106580974188 2.9267e-08 1.8405702321245123 2.9267999999999998e-08 1.7962392420834836 2.9269e-08 1.7465140796641756 2.927e-08 1.849557979544189 2.9270999999999998e-08 1.7808418787002223 2.9272e-08 1.8474954014535072 2.9273e-08 1.754394040887867 2.9273999999999998e-08 1.7012906751945203 2.9275e-08 1.8222016812020283 2.9276e-08 1.8119649597441196 2.9276999999999998e-08 1.8129701211474445 2.9278e-08 1.7442361637073953 2.9279e-08 1.751266750559959 2.9279999999999998e-08 1.8086672762237739 2.9281e-08 1.8349505162064415 2.9282e-08 1.842369752788252 2.9282999999999998e-08 1.8256655664691472 2.9284e-08 1.7709698544738055 2.9285e-08 1.882638999410819 2.9285999999999998e-08 1.8271771275793776 2.9287e-08 1.7983832594334337 2.9288e-08 1.7868979965696101 2.9289e-08 1.7605901525273246 2.929e-08 1.788727118914128 2.9291e-08 1.792179473234385 2.9292e-08 1.853086525265168 2.9293e-08 1.7822143548782432 2.9294e-08 1.8296683756315146 2.9295e-08 1.8137617630794314 2.9296e-08 1.9079160094366627 2.9297e-08 1.7400257855189905 2.9298e-08 1.8597897056742154 2.9299e-08 1.7927984611243748 2.93e-08 1.785060221150784 2.9301e-08 1.8420116126988444 2.9302e-08 1.7211489033444611 2.9302999999999998e-08 1.8076539309206112 2.9304e-08 1.8080824847207306 2.9305e-08 1.8093999396669578 2.9305999999999998e-08 1.7320677348305897 2.9307e-08 1.7767234756237211 2.9308e-08 1.7705187903893609 2.9308999999999998e-08 1.8066912385942033 2.931e-08 1.7170495011305382 2.9311e-08 1.7901433900697319 2.9311999999999998e-08 1.8118616662411045 2.9313e-08 1.8191590606787276 2.9314e-08 1.7336489279120715 2.9314999999999998e-08 1.7708465928447308 2.9316e-08 1.817260308902085 2.9317e-08 1.7799266175120219 2.9317999999999998e-08 1.6821121217638249 2.9319e-08 1.833878281453363 2.932e-08 1.8605313138443265 2.9320999999999998e-08 1.7753287956407477 2.9322e-08 1.80277048378021 2.9323e-08 1.7949592609884946 2.9324e-08 1.7778840862222087 2.9325e-08 1.8502137738786348 2.9326e-08 1.775390083967441 2.9327e-08 1.8956819497878175 2.9328e-08 1.8281250251792858 2.9329e-08 1.7429892511482592 2.933e-08 1.7125796859672509 2.9331e-08 1.7574285905864453 2.9332e-08 1.8069757718681 2.9333e-08 1.7603938521352644 2.9334e-08 1.8561254683363693 2.9335e-08 1.8071670031076088 2.9336e-08 1.7930295033678196 2.9337e-08 1.818743862854402 2.9338e-08 1.8413833584278154 2.9339e-08 1.7445315609791194 2.934e-08 1.8155373232246643 2.9340999999999998e-08 1.802724919381727 2.9342e-08 1.7564993402501543 2.9343e-08 1.7210031359797453 2.9343999999999998e-08 1.7592863750386727 2.9345e-08 1.8008449960410993 2.9346e-08 1.7970550678689625 2.9346999999999998e-08 1.839960474182517 2.9348e-08 1.861144611278678 2.9349e-08 1.8362655954292755 2.9349999999999998e-08 1.8397220837060848 2.9351e-08 1.796822866601699 2.9352e-08 1.7314231881580067 2.9352999999999998e-08 1.7885970068468569 2.9354e-08 1.7942050053324337 2.9355e-08 1.755735250698327 2.9355999999999998e-08 1.7638835574884422 2.9357e-08 1.848131994003832 2.9358e-08 1.8117525313658294 2.9359e-08 1.7787120725197958 2.936e-08 1.7583787596102782 2.9361e-08 1.8435748321277554 2.9362e-08 1.8268466086041444 2.9363e-08 1.7331350570280502 2.9364e-08 1.7755038690413976 2.9365e-08 1.76394596560787 2.9366e-08 1.89111629611341 2.9367e-08 1.909918646841442 2.9368e-08 1.825059986686674 2.9369e-08 1.8293766806148228 2.937e-08 1.844039913696295 2.9371e-08 1.7767453108048015 2.9372e-08 1.7825106436601759 2.9373e-08 1.8591046604143524 2.9374e-08 1.7420823007157873 2.9375e-08 1.7044606615159994 2.9375999999999998e-08 1.8615108071444375 2.9377e-08 1.7980725838681981 2.9378e-08 1.69593332859962 2.9378999999999998e-08 1.8239463391226616 2.938e-08 1.8376585116707804 2.9381e-08 1.8503240522052002 2.9381999999999998e-08 1.7894421466608834 2.9383e-08 1.7945126442849895 2.9384e-08 1.816487583329205 2.9384999999999998e-08 1.8247540649561347 2.9386e-08 1.7688412076832443 2.9387e-08 1.7549579677400726 2.9387999999999998e-08 1.8894720410314743 2.9389e-08 1.7874091126690734 2.939e-08 1.859113233187834 2.9390999999999998e-08 1.812941813181029 2.9392e-08 1.8229707534362274 2.9393e-08 1.8827277742189685 2.9394e-08 1.738821503896971 2.9395e-08 1.7084107636803685 2.9396e-08 1.7753669094722047 2.9397e-08 1.8419521566677344 2.9398e-08 1.9631689936684924 2.9399e-08 1.770324034299122 2.94e-08 1.8798183988340027 2.9401e-08 1.8311823425689864 2.9402e-08 1.8475292725841228 2.9403e-08 1.742586982953852 2.9404e-08 1.7715148383076238 2.9405e-08 1.798527767487559 2.9406e-08 1.7318029135480328 2.9407e-08 1.8090379061395279 2.9408e-08 1.7581066312587659 2.9409e-08 1.8029656841529216 2.941e-08 1.815074563581303 2.9410999999999998e-08 1.819435142414041 2.9412e-08 1.7648553639606037 2.9413e-08 1.799744156190583 2.9413999999999998e-08 1.8340726948239052 2.9415e-08 1.8342883316634986 2.9416e-08 1.8706393477256007 2.9416999999999998e-08 1.8279530712439025 2.9418e-08 1.7929215910879743 2.9419e-08 1.6607153599763211 2.9419999999999998e-08 1.790217979705674 2.9421e-08 1.8113838233883819 2.9422e-08 1.792353846164673 2.9422999999999998e-08 1.7027239969243788 2.9424e-08 1.7832726432023123 2.9425e-08 1.7834197104410467 2.9425999999999998e-08 1.8701793226689425 2.9427e-08 1.7350674370217147 2.9428e-08 1.826660098091229 2.9429e-08 1.7443596585056103 2.943e-08 1.8002806609317865 2.9431e-08 1.7709616521196636 2.9432e-08 1.8162774054325026 2.9433e-08 1.7785116141343087 2.9434e-08 1.765416491604274 2.9435e-08 1.7126822017556655 2.9436e-08 1.7523022883461075 2.9437e-08 1.8443115148562834 2.9438e-08 1.8838000673023545 2.9439e-08 1.7560516194091873 2.944e-08 1.7209370694123725 2.9441e-08 1.6907253875495991 2.9442e-08 1.772851816124216 2.9443e-08 1.7743459235147463 2.9444e-08 1.7679349278473901 2.9445e-08 1.8614071201354887 2.9445999999999998e-08 1.7847907611200546 2.9447e-08 1.7533467012617883 2.9448e-08 1.7927511961810096 2.9448999999999998e-08 1.726393813755756 2.945e-08 1.8616667102204392 2.9451e-08 1.7407335037748655 2.9451999999999998e-08 1.8173393418386936 2.9453e-08 1.7236565067528606 2.9454e-08 1.7928475639292603 2.9454999999999998e-08 1.8515653586593523 2.9456e-08 1.823972127093285 2.9457e-08 1.8366833984210722 2.9457999999999998e-08 1.7014286014943398 2.9459e-08 1.8490517751336202 2.946e-08 1.9038276118450481 2.9460999999999998e-08 1.6913892998266695 2.9462e-08 1.812768241224515 2.9463e-08 1.7779854206756536 2.9463999999999998e-08 1.752052401769503 2.9465e-08 1.8507132203958756 2.9466e-08 1.8678797817544828 2.9467e-08 1.8562517908497818 2.9468e-08 1.7310418531169638 2.9469e-08 1.7724004035618592 2.947e-08 1.808152828707673 2.9471e-08 1.7414926423425325 2.9472e-08 1.7993332313986314 2.9473e-08 1.8177474692439974 2.9474e-08 1.8781476829115682 2.9475e-08 1.844845635110669 2.9476e-08 1.8582361598339363 2.9477e-08 1.7992558103709329 2.9478e-08 1.752591622194948 2.9479e-08 1.8059857385541573 2.948e-08 1.8070643886723543 2.9480999999999998e-08 1.826993470350075 2.9482e-08 1.874591442653007 2.9483e-08 1.7296637899979497 2.9483999999999998e-08 1.7357096564803252 2.9485e-08 1.832187959304565 2.9486e-08 1.8949518384595203 2.9486999999999998e-08 1.775781415259531 2.9488e-08 1.7041487745761443 2.9489e-08 1.7495363634228003 2.9489999999999998e-08 1.8539338641165788 2.9491e-08 1.8468193947671216 2.9492e-08 1.805512259623778 2.9492999999999998e-08 1.7487805512665033 2.9494e-08 1.785891437603029 2.9495e-08 1.7778812293105923 2.9495999999999998e-08 1.831584494947086 2.9497e-08 1.7887935167727937 2.9498e-08 1.8883389249252471 2.9498999999999998e-08 1.714247391283041 2.95e-08 1.7827863617375301 2.9501e-08 1.8143211770445875 2.9502e-08 1.8023250169345546 2.9503e-08 1.7149981115005173 2.9504e-08 1.790851694829152 2.9505e-08 1.8376932165065807 2.9506e-08 1.8344717100819676 2.9507e-08 1.7744151549515488 2.9508e-08 1.8118715428001069 2.9509e-08 1.6905273168360573 2.951e-08 1.8224167371787527 2.9511e-08 1.804382974699646 2.9512e-08 1.7603771711581186 2.9513e-08 1.7284790439235507 2.9514e-08 1.7923735631637323 2.9515e-08 1.7345981406868294 2.9516e-08 1.8115038776983723 2.9517e-08 1.817585514862386 2.9518e-08 1.740834368531458 2.9518999999999998e-08 1.809889964485307 2.952e-08 1.7305006547431256 2.9521e-08 1.765963914822838 2.9521999999999998e-08 1.7809092410843057 2.9523e-08 1.7857984711295127 2.9524e-08 1.866264144358723 2.9524999999999998e-08 1.8697978771858486 2.9526e-08 1.9267366346332835 2.9527e-08 1.8358636880319958 2.9527999999999998e-08 1.7988318329599695 2.9529e-08 1.8019913944024577 2.953e-08 1.840718769115959 2.9530999999999998e-08 1.7867016946751766 2.9532e-08 1.7941596881327218 2.9533e-08 1.7999974561276393 2.9533999999999998e-08 1.8456477635847561 2.9535e-08 1.8238660431017841 2.9536e-08 1.7338377649067134 2.9537e-08 1.754916312016763 2.9538e-08 1.81061667548762 2.9539e-08 1.8542095127121374 2.954e-08 1.7701328765788797 2.9541e-08 1.8199500149543832 2.9542e-08 1.7819949263752957 2.9543e-08 1.78704089329621 2.9544e-08 1.8301070459497424 2.9545e-08 1.6634426590690012 2.9546e-08 1.8211093330851398 2.9547e-08 1.7827189609700893 2.9548e-08 1.8514897982987244 2.9549e-08 1.8081851567407559 2.955e-08 1.8193472106358015 2.9551e-08 1.9048486514796665 2.9552e-08 1.7442632051227038 2.9553e-08 1.7426733553652385 2.9553999999999998e-08 1.8021921682849764 2.9555e-08 1.8071909097475227 2.9556e-08 1.837810184535753 2.9556999999999998e-08 1.7900678294272556 2.9558e-08 1.7768396076108472 2.9559e-08 1.7251424391394987 2.9559999999999998e-08 1.7540163418196228 2.9561e-08 1.8945524899170731 2.9562e-08 1.8444578773326408 2.9562999999999998e-08 1.8411655520541506 2.9564e-08 1.7282079793940603 2.9565e-08 1.773002646730135 2.9565999999999998e-08 1.7046608595028423 2.9567e-08 1.7669473809515726 2.9568e-08 1.787677814634982 2.9568999999999998e-08 1.8307526282325979 2.957e-08 1.7912125718467085 2.9571e-08 1.7062138430844063 2.9572e-08 1.8117033037497616 2.9573e-08 1.7677328102295682 2.9574e-08 1.8443180988801218 2.9575e-08 1.6705107139811992 2.9576e-08 1.799162403004946 2.9577e-08 1.8597976353604286 2.9578e-08 1.7808473681497954 2.9579e-08 1.7640346284309072 2.958e-08 1.8218555004426753 2.9581e-08 1.696922532073219 2.9582e-08 1.7738915796892025 2.9583e-08 1.886849291526599 2.9584e-08 1.8283339109158978 2.9585e-08 1.7657119459538053 2.9586e-08 1.8233353015080331 2.9587e-08 1.8946854883077002 2.9588e-08 1.7732673980108649 2.9588999999999998e-08 1.7624004999377856 2.959e-08 1.8534585946022482 2.9591e-08 1.7688244377020914 2.9591999999999998e-08 1.8160243160313787 2.9593e-08 1.6970183429197805 2.9594e-08 1.8694630508356147 2.9594999999999998e-08 1.797493612535435 2.9596e-08 1.831454213678316 2.9597e-08 1.7684733949549394 2.9597999999999998e-08 1.7987654109396134 2.9599e-08 1.7538334384061147 2.96e-08 1.8435836335191367 2.9600999999999998e-08 1.7923843620983042 2.9602e-08 1.8150098224612365 2.9603e-08 1.8592212669605588 2.9603999999999998e-08 1.8358410384900277 2.9605e-08 1.8377597546416742 2.9606e-08 1.8689409949017557 2.9607e-08 1.7987510437090066 2.9608e-08 1.8434038244791238 2.9609e-08 1.8388021000354104 2.961e-08 1.8746802460424563 2.9611e-08 1.762808318259574 2.9612e-08 1.8674523242000884 2.9613e-08 1.8639530094904202 2.9614e-08 1.8350419635386683 2.9615e-08 1.7917576905590942 2.9616e-08 1.740184157131463 2.9617e-08 1.780691370390067 2.9618e-08 1.7825380388534537 2.9619e-08 1.8290958487789117 2.962e-08 1.7500594492400947 2.9621e-08 1.7258978010972719 2.9622e-08 1.7507611433374868 2.9623e-08 1.7573638379841467 2.9623999999999998e-08 1.8418671994264908 2.9625e-08 1.8154530444771766 2.9626e-08 1.784213296886224 2.9626999999999998e-08 1.7792273745319849 2.9628e-08 1.796821514290184 2.9629e-08 1.8819705573903511 2.9629999999999998e-08 1.8131519143589265 2.9631e-08 1.7198838941420822 2.9632e-08 1.811086295051792 2.9632999999999998e-08 1.7813956372576005 2.9634e-08 1.7997537744719805 2.9635e-08 1.847131654920086 2.9635999999999998e-08 1.7976345986312272 2.9637e-08 1.7391916062443735 2.9638e-08 1.8186116009426998 2.9638999999999998e-08 1.7716750815709765 2.964e-08 1.8136072159851255 2.9641e-08 1.8395667901864077 2.9642e-08 1.7644112835317267 2.9643e-08 1.7776424180643577 2.9644e-08 1.7643753467230268 2.9645e-08 1.8303160530136637 2.9646e-08 1.786036776767341 2.9647e-08 1.8669548635035533 2.9648e-08 1.9374796503978957 2.9649e-08 1.7776714523491532 2.965e-08 1.7747941059666978 2.9651e-08 1.7572127090305956 2.9652e-08 1.7946380721596036 2.9653e-08 1.8270873671645584 2.9654e-08 1.8551275975737407 2.9655e-08 1.791677170067362 2.9656e-08 1.8113840590771004 2.9657e-08 1.7864650942230833 2.9658e-08 1.7560818942081406 2.9658999999999998e-08 1.7640808814928204 2.966e-08 1.7753459924352606 2.9661e-08 1.7718928094948994 2.9661999999999998e-08 1.7209361848240472 2.9663e-08 1.640754451743686 2.9664e-08 1.7853733038611426 2.9664999999999998e-08 1.7234201788191232 2.9666e-08 1.8377681250692943 2.9667e-08 1.8717230795598456 2.9667999999999998e-08 1.8102887727579535 2.9669e-08 1.7066705167223124 2.967e-08 1.829823170092875 2.9670999999999998e-08 1.818385615544698 2.9672e-08 1.8670442306151822 2.9673e-08 1.8658056652494606 2.9673999999999998e-08 1.8566690501907792 2.9675e-08 1.806097976969375 2.9676e-08 1.7793712675775832 2.9676999999999998e-08 1.7032354598658936 2.9678e-08 1.7634809711046298 2.9679e-08 1.8089670953908144 2.968e-08 1.7947018695977714 2.9681e-08 1.789422717733379 2.9682e-08 1.790808083230043 2.9683e-08 1.8339676060844505 2.9684e-08 1.7888292890860717 2.9685e-08 1.86632727577575 2.9686e-08 1.821383537654179 2.9687e-08 1.773177240958194 2.9688e-08 1.753817955723792 2.9689e-08 1.7625926369495166 2.969e-08 1.8022606178709306 2.9691e-08 1.7790897656624376 2.9692e-08 1.850586452892745 2.9693e-08 1.837558579787801 2.9693999999999998e-08 1.8421047226020923 2.9695e-08 1.7655950032914782 2.9696e-08 1.864139541476929 2.9696999999999998e-08 1.7747552079241324 2.9698e-08 1.7875768034106778 2.9699e-08 1.8470766570784836 2.9699999999999998e-08 1.70806913258096 2.9701e-08 1.7591165313888715 2.9702e-08 1.8402712068530072 2.9702999999999998e-08 1.7289604924908266 2.9704e-08 1.6877178005915452 2.9705e-08 1.8150154690892026 2.9705999999999998e-08 1.8461290805146928 2.9707e-08 1.8994546361488258 2.9708e-08 1.811054922273044 2.9708999999999998e-08 1.6987818104202157 2.971e-08 1.684015876492094 2.9711e-08 1.8230216459955646 2.9711999999999998e-08 1.8454901834260877 2.9713e-08 1.8527438176051023 2.9714e-08 1.8139720268805137 2.9715e-08 1.8233023409319007 2.9716e-08 1.8257500742904467 2.9717e-08 1.7079333296208896 2.9718e-08 1.8267783927001577 2.9719e-08 1.7372017314372123 2.972e-08 1.7558435437445472 2.9721e-08 1.7879588067526497 2.9722e-08 1.789671194937474 2.9723e-08 1.7606353228770424 2.9724e-08 1.784455416845104 2.9725e-08 1.8252220624190285 2.9726e-08 1.8145743715270437 2.9727e-08 1.838504930541949 2.9728e-08 1.8242446816740165 2.9729e-08 1.7522039421172437 2.973e-08 1.7975015431458419 2.9731e-08 1.798891755720687 2.9731999999999998e-08 1.882800096277502 2.9733e-08 1.736576277985423 2.9734e-08 1.7701776186476335 2.9734999999999998e-08 1.917720695812187 2.9736e-08 1.77969559959821 2.9737e-08 1.822726100400316 2.9737999999999998e-08 1.731599271265168 2.9739e-08 1.7064657983722276 2.974e-08 1.869472151423817 2.9740999999999998e-08 1.853176818246089 2.9742e-08 1.7915114913283603 2.9743e-08 1.7044506700020574 2.9743999999999998e-08 1.8232616719732686 2.9745e-08 1.8466925128162166 2.9746e-08 1.7601898765794937 2.9746999999999998e-08 1.8173465734503558 2.9748e-08 1.806204736648216 2.9749e-08 1.7880204653087866 2.975e-08 1.8495106703781239 2.9751e-08 1.7888781527902644 2.9752e-08 1.791726663353143 2.9753e-08 1.817746023921029 2.9754e-08 1.8303683453114479 2.9755e-08 1.817936994503774 2.9756e-08 1.7735461872754177 2.9757e-08 1.814608477883438 2.9758e-08 1.7358357078690267 2.9759e-08 1.7727445172945138 2.976e-08 1.8800733501314768 2.9761e-08 1.9449264239923527 2.9762e-08 1.7911670084725977 2.9763e-08 1.7618161027207278 2.9764e-08 1.7389896305787595 2.9765e-08 1.8627617904423093 2.9766e-08 1.7992787986434473 2.9766999999999998e-08 1.7773878679097255 2.9768e-08 1.835629087500101 2.9769e-08 1.7257900940469204 2.9769999999999998e-08 1.743374553088413 2.9771e-08 1.8328965605877718 2.9772e-08 1.6893885169652731 2.9772999999999998e-08 1.768793749590732 2.9774e-08 1.7843301531390614 2.9775e-08 1.7748133274797901 2.9775999999999998e-08 1.7745213088423317 2.9777e-08 1.7993389082732674 2.9778e-08 1.7971670377627436 2.9778999999999998e-08 1.830171888647183 2.978e-08 1.7114387218685745 2.9781e-08 1.7963508415521248 2.9781999999999998e-08 1.8264567534702754 2.9783e-08 1.8324712252685773 2.9784e-08 1.7023705030283633 2.9785e-08 1.7593649097047428 2.9786e-08 1.8067863429368998 2.9787e-08 1.8569790297873425 2.9788e-08 1.8187822208862683 2.9789e-08 1.797905387329762 2.979e-08 1.8005930676843906 2.9791e-08 1.7731550768524689 2.9792e-08 1.7534569962981255 2.9793e-08 1.7423605975751486 2.9794e-08 1.845326361560544 2.9795e-08 1.8091106831707577 2.9796e-08 1.811995904144605 2.9797e-08 1.7575505609301723 2.9798e-08 1.8349165445848326 2.9799e-08 1.8362876782292095 2.98e-08 1.9134177324035533 2.9801e-08 1.7674067130932545 2.9801999999999998e-08 1.7889358364646062 2.9803e-08 1.7990126829957693 2.9804e-08 1.880512535653395 2.9805e-08 1.813460526631688 2.9806e-08 1.823321278754615 2.9807e-08 1.753850892667964 2.9808e-08 1.827459878524299 2.9809e-08 1.8051539893099082 2.981e-08 1.7766745748546224 2.9811e-08 1.828581994922976 2.9812e-08 1.7948884138695607 2.9813e-08 1.8439663923531402 2.9814e-08 1.8003952985469243 2.9815e-08 1.7464828611560246 2.9816e-08 1.8772414857574846 2.9817e-08 1.7488033427580456 2.9818e-08 1.7976479760614827 2.9819e-08 1.7896151328999723 2.982e-08 1.800821302412415 2.9821e-08 1.7606066090736952 2.9822e-08 1.7267884367766724 2.9823e-08 1.8757950270200245 2.9823999999999996e-08 1.8840374481558249 2.9825e-08 1.8655720873574277 2.9826e-08 1.7614510742097889 2.9827e-08 1.7640144687213672 2.9828e-08 1.7645660808402406 2.9829e-08 1.8154340373211184 2.9829999999999996e-08 1.7535004488834234 2.9831e-08 1.7032773239247077 2.9832e-08 1.8413505694249024 2.9833e-08 1.7633386745141384 2.9834e-08 1.7981747509676989 2.9835e-08 1.8202486009111827 2.9835999999999997e-08 1.7797728151884569 2.9837e-08 1.7220473041280004 2.9838e-08 1.8254929018059725 2.9839e-08 1.8169526885258909 2.984e-08 1.8194043630647176 2.9841e-08 1.6803468508741932 2.9842e-08 1.764942275860347 2.9843e-08 1.7543971849128182 2.9844e-08 1.8061595484349968 2.9845e-08 1.785669484917831 2.9846e-08 1.7373844383589103 2.9847e-08 1.8256191897121474 2.9848e-08 1.8046801069955705 2.9849e-08 1.7678245085865325 2.985e-08 1.760551851246479 2.9851e-08 1.7157436891931166 2.9852e-08 1.7075415018133402 2.9853e-08 1.7545796437656174 2.9854e-08 1.7837116142474034 2.9855e-08 1.8519861771757558 2.9856e-08 1.7576092081623182 2.9857e-08 1.860128904298766 2.9858e-08 1.8389039315249482 2.9858999999999996e-08 1.8170313065705996 2.986e-08 1.7524277741643604 2.9861e-08 1.77104733213901 2.9862e-08 1.8672456081304436 2.9863e-08 1.7683486879721455 2.9864e-08 1.7306808458333338 2.9864999999999996e-08 1.8929884873211966 2.9866e-08 1.7616031566870316 2.9867e-08 1.7462587525172868 2.9868e-08 1.7972376834676085 2.9869e-08 1.8380434155009688 2.987e-08 1.8140226024854622 2.9870999999999997e-08 1.8162459341935158 2.9872e-08 1.80621347764155 2.9873e-08 1.7885805519080327 2.9874e-08 1.7894298327475846 2.9875e-08 1.7539468828160194 2.9876e-08 1.8269421611489098 2.9877e-08 1.8580640142289255 2.9878e-08 1.7797693396372445 2.9879e-08 1.8089644326541403 2.988e-08 1.894709523557029 2.9881e-08 1.657008736050212 2.9882e-08 1.79052663695294 2.9883e-08 1.7573865237999575 2.9884e-08 1.8945064995268432 2.9885e-08 1.8333257134754513 2.9886e-08 1.8423087296043092 2.9887e-08 1.7173522524704736 2.9888e-08 1.7812003708581003 2.9889e-08 1.7857864217201558 2.989e-08 1.778777617277111 2.9891e-08 1.772757170945903 2.9892e-08 1.7961362174514024 2.9893e-08 1.76252372490829 2.9893999999999996e-08 1.7368248534972508 2.9895e-08 1.735198410558104 2.9896e-08 1.8332648205994726 2.9897e-08 1.83233585595843 2.9898e-08 1.810680821643706 2.9899e-08 1.811665805756362 2.9899999999999996e-08 1.7600767354293887 2.9901e-08 1.82830350915094 2.9902e-08 1.8088449497461514 2.9903e-08 1.7870141475917185 2.9904e-08 1.8484568162509736 2.9905e-08 1.7579614983121017 2.9905999999999997e-08 1.8275359997958216 2.9907e-08 1.7358414880465338 2.9908e-08 1.7509488612821154 2.9909e-08 1.8309154017312483 2.991e-08 1.818246086247737 2.9911e-08 1.8071840599577589 2.9912e-08 1.771261827626345 2.9913e-08 1.7932122787895333 2.9914e-08 1.8213435057582272 2.9915e-08 1.79410146888971 2.9916e-08 1.8825296159506637 2.9917e-08 1.7681506487247596 2.9918e-08 1.7595389167389346 2.9919e-08 1.7518184199471105 2.992e-08 1.8544144045576143 2.9921e-08 1.8431647984036772 2.9922e-08 1.9291363516776487 2.9923e-08 1.8215086153909272 2.9924e-08 1.974597236984574 2.9925e-08 1.8000731640685217 2.9926e-08 1.7539384537668121 2.9927e-08 1.8621987684664436 2.9928e-08 1.7464685109355869 2.9928999999999996e-08 1.884990859650752 2.993e-08 1.7518933289657639 2.9931e-08 1.7710131410979648 2.9932e-08 1.777775566079411 2.9933e-08 1.8136101023610989 2.9934e-08 1.8484216518560428 2.9934999999999996e-08 1.8420122479197385 2.9936e-08 1.7869003433417756 2.9937e-08 1.796235530567994 2.9938e-08 1.7542574214896127 2.9939e-08 1.7966028636056326 2.994e-08 1.7554146051309663 2.9940999999999997e-08 1.7500923420415955 2.9942e-08 1.6661205723509218 2.9943e-08 1.8683835396422137 2.9944e-08 1.7717523143623006 2.9945e-08 1.7805576829061343 2.9946e-08 1.7724582678352503 2.9947e-08 1.7653190311363556 2.9948e-08 1.7266281934507988 2.9949e-08 1.8789213286365702 2.995e-08 1.7247365307048175 2.9951e-08 1.9512552457889123 2.9952e-08 1.8543138396548908 2.9953e-08 1.8104275298151857 2.9954e-08 1.8882491448948786 2.9955e-08 1.8941457490794076 2.9956e-08 1.7844557738807054 2.9957e-08 1.7908536719265598 2.9958e-08 1.7760356243974962 2.9959e-08 1.7508601330986535 2.996e-08 1.8060755286281702 2.9961e-08 1.7772928510346742 2.9962e-08 1.8710372168185727 2.9963e-08 1.81263690941238 2.9963999999999996e-08 1.7993542437002361 2.9965e-08 1.8010920089876796 2.9966e-08 1.7831675084748948 2.9967e-08 1.8332026588817252 2.9968e-08 1.7813321343403683 2.9969e-08 1.7225049917442687 2.9969999999999996e-08 1.8404851121366161 2.9971e-08 1.7330863772289533 2.9972e-08 1.8531184517051613 2.9973e-08 1.7315175775381486 2.9974e-08 1.743307116659538 2.9975e-08 1.8091479551338876 2.9975999999999997e-08 1.7806213927076648 2.9977e-08 1.8610489803881922 2.9978e-08 1.765554940926753 2.9979e-08 1.8658251308663967 2.998e-08 1.7677840998423788 2.9981e-08 1.829492961668335 2.9982e-08 1.7998968959567307 2.9983e-08 1.801950549066446 2.9984e-08 1.9212774406166049 2.9985e-08 1.8031298811272194 2.9986e-08 1.7918266587575413 2.9987e-08 1.82995802192256 2.9988e-08 1.7364008770858665 2.9989e-08 1.6868758501815864 2.999e-08 1.7486109619473986 2.9991e-08 1.8169124215399115 2.9992e-08 1.6975427370857523 2.9993e-08 1.8230385943435512 2.9994e-08 1.939445629954557 2.9995e-08 1.7882712572382438 2.9996e-08 1.8350015031270523 2.9997e-08 1.7970685304447735 2.9998e-08 1.8376500052008125 2.9998999999999996e-08 1.7742823294772054 )
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/ss.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/ss/specialized_cells.spice




.option method=gear
.option wnflag=1
.option savecurrents


.save
+@m.xm1.msky130_fd_pr__nfet_01v8[gm]
+@m.xm2.msky130_fd_pr__pfet_01v8[gm]
+@m.xm3.msky130_fd_pr__nfet_01v8[gm]
+@m.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.xm5.msky130_fd_pr__nfet_01v8[gm]
+@m.xm6.msky130_fd_pr__pfet_01v8[gm]

.temp 75
.ic v(osc)=0

.control
  save all
  tran 1ps 30ns
  remzerovec
  linearize v(osc) v(vdd)
  write test_inverter_speed.raw
  wrdata /foss/designs/my_design/projects/pll/bandgapref/xschem_ngspice/oscillator.txt v(osc)
  set appendwrite
.endc




**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
