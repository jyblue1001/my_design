magic
tech sky130A
timestamp 1737651475
<< nwell >>
rect -468 88 1054 464
<< nmos >>
rect 0 -5 22 38
rect -130 -145 -115 -45
rect -65 -145 -50 -45
rect 419 -5 441 38
rect 77 -145 92 -102
rect 354 -145 369 -45
rect 838 -5 860 38
rect 496 -145 511 -102
rect 773 -145 788 -45
rect 915 -145 931 -102
<< pmos >>
rect -400 229 -250 429
rect -200 229 -50 429
rect 77 229 92 315
rect 219 229 369 429
rect 496 229 511 315
rect 638 229 788 429
rect 915 229 930 315
rect 0 106 22 192
rect 419 106 441 192
rect 838 106 860 192
<< ndiff >>
rect -50 30 0 38
rect -50 5 -35 30
rect -15 5 0 30
rect -50 -5 0 5
rect 22 30 72 38
rect 22 5 37 30
rect 57 5 72 30
rect 22 -5 72 5
rect -180 -55 -130 -45
rect -180 -135 -165 -55
rect -145 -135 -130 -55
rect -180 -145 -130 -135
rect -115 -55 -65 -45
rect -115 -135 -100 -55
rect -80 -135 -65 -55
rect -115 -145 -65 -135
rect -50 -55 0 -45
rect -50 -135 -35 -55
rect -15 -135 0 -55
rect 369 30 419 38
rect 369 5 384 30
rect 404 5 419 30
rect 369 -5 419 5
rect 441 30 491 38
rect 441 5 456 30
rect 476 5 491 30
rect 441 -5 491 5
rect 304 -55 354 -45
rect -50 -145 0 -135
rect 27 -112 77 -102
rect 27 -135 42 -112
rect 62 -135 77 -112
rect 27 -145 77 -135
rect 92 -112 142 -102
rect 92 -135 107 -112
rect 127 -135 142 -112
rect 92 -145 142 -135
rect 304 -135 319 -55
rect 339 -135 354 -55
rect 304 -145 354 -135
rect 369 -55 419 -45
rect 369 -135 384 -55
rect 404 -135 419 -55
rect 788 30 838 38
rect 788 5 803 30
rect 823 5 838 30
rect 788 -5 838 5
rect 860 30 910 38
rect 860 5 875 30
rect 895 5 910 30
rect 860 -5 910 5
rect 723 -55 773 -45
rect 369 -145 419 -135
rect 446 -112 496 -102
rect 446 -135 461 -112
rect 481 -135 496 -112
rect 446 -145 496 -135
rect 511 -112 561 -102
rect 511 -135 526 -112
rect 546 -135 561 -112
rect 511 -145 561 -135
rect 723 -135 738 -55
rect 758 -135 773 -55
rect 723 -145 773 -135
rect 788 -55 839 -45
rect 788 -135 803 -55
rect 823 -135 839 -55
rect 788 -145 839 -135
rect 866 -112 915 -102
rect 866 -135 881 -112
rect 901 -135 915 -112
rect 866 -145 915 -135
rect 931 -112 980 -102
rect 931 -135 945 -112
rect 966 -135 980 -112
rect 931 -145 980 -135
<< pdiff >>
rect -450 419 -400 429
rect -450 239 -435 419
rect -415 239 -400 419
rect -450 229 -400 239
rect -250 419 -200 429
rect -250 239 -235 419
rect -215 239 -200 419
rect -250 229 -200 239
rect -50 419 0 429
rect -50 239 -35 419
rect -15 239 0 419
rect 169 419 219 429
rect -50 229 0 239
rect 27 305 77 315
rect 27 239 42 305
rect 62 239 77 305
rect 27 229 77 239
rect 92 305 142 315
rect 92 239 107 305
rect 127 239 142 305
rect 92 229 142 239
rect 169 239 184 419
rect 204 239 219 419
rect 169 229 219 239
rect 369 419 419 429
rect 369 239 384 419
rect 404 239 419 419
rect 588 419 638 429
rect 369 229 419 239
rect 446 305 496 315
rect 446 239 461 305
rect 481 239 496 305
rect 446 229 496 239
rect 511 305 561 315
rect 511 239 526 305
rect 546 239 561 305
rect 511 229 561 239
rect 588 239 603 419
rect 623 239 638 419
rect 588 229 638 239
rect 788 419 838 429
rect 788 239 803 419
rect 823 239 838 419
rect 788 229 838 239
rect 865 305 915 315
rect 865 239 880 305
rect 900 239 915 305
rect 865 229 915 239
rect 930 305 980 315
rect 930 239 945 305
rect 965 239 980 305
rect 930 229 980 239
rect -50 184 0 192
rect -50 116 -35 184
rect -15 116 0 184
rect -50 106 0 116
rect 22 184 72 192
rect 22 116 37 184
rect 57 116 72 184
rect 22 106 72 116
rect 369 184 419 192
rect 369 116 384 184
rect 404 116 419 184
rect 369 106 419 116
rect 441 184 491 192
rect 441 116 456 184
rect 476 116 491 184
rect 441 106 491 116
rect 788 184 838 192
rect 788 116 803 184
rect 823 116 838 184
rect 788 106 838 116
rect 860 184 910 192
rect 860 116 875 184
rect 895 116 910 184
rect 860 106 910 116
<< ndiffc >>
rect -35 5 -15 30
rect 37 5 57 30
rect -165 -135 -145 -55
rect -100 -135 -80 -55
rect -35 -135 -15 -55
rect 384 5 404 30
rect 456 5 476 30
rect 42 -135 62 -112
rect 107 -135 127 -112
rect 319 -135 339 -55
rect 384 -135 404 -55
rect 803 5 823 30
rect 875 5 895 30
rect 461 -135 481 -112
rect 526 -135 546 -112
rect 738 -135 758 -55
rect 803 -135 823 -55
rect 881 -135 901 -112
rect 945 -135 966 -112
<< pdiffc >>
rect -435 239 -415 419
rect -235 239 -215 419
rect -35 239 -15 419
rect 42 239 62 305
rect 107 239 127 305
rect 184 239 204 419
rect 384 239 404 419
rect 461 239 481 305
rect 526 239 546 305
rect 603 239 623 419
rect 803 239 823 419
rect 880 239 900 305
rect 945 239 965 305
rect -35 116 -15 184
rect 37 116 57 184
rect 384 116 404 184
rect 456 116 476 184
rect 803 116 823 184
rect 875 116 895 184
<< psubdiff >>
rect 254 -55 304 -45
rect 142 -112 192 -102
rect 142 -135 157 -112
rect 177 -135 192 -112
rect 142 -145 192 -135
rect 254 -135 269 -55
rect 289 -135 304 -55
rect 254 -145 304 -135
rect 561 -112 611 -102
rect 561 -135 576 -112
rect 596 -135 611 -112
rect 561 -145 611 -135
rect 980 -112 1030 -102
rect 980 -135 995 -112
rect 1015 -135 1030 -112
rect 980 -145 1030 -135
<< nsubdiff >>
rect 980 305 1030 315
rect 980 239 995 305
rect 1015 239 1030 305
rect 980 229 1030 239
<< psubdiffcont >>
rect 157 -135 177 -112
rect 269 -135 289 -55
rect 576 -135 596 -112
rect 995 -135 1015 -112
<< nsubdiffcont >>
rect 995 239 1015 305
<< poly >>
rect -400 444 788 464
rect -400 429 -250 444
rect -200 429 -50 444
rect 219 429 369 444
rect 638 429 788 444
rect 77 315 92 330
rect 496 315 511 330
rect 915 315 930 330
rect -400 214 -250 229
rect -200 214 -50 229
rect 77 214 92 229
rect 219 214 369 229
rect 496 214 511 229
rect 638 214 788 229
rect 915 214 930 229
rect -400 204 -360 214
rect -400 184 -389 204
rect -369 184 -360 204
rect 0 192 22 207
rect 77 199 177 214
rect -400 174 -360 184
rect 92 168 132 178
rect 92 148 102 168
rect 122 148 132 168
rect 92 138 132 148
rect 0 87 22 106
rect -40 82 22 87
rect -280 62 -30 82
rect -10 62 22 82
rect -280 -152 -260 62
rect -40 57 22 62
rect 0 38 22 57
rect 0 -20 22 -5
rect -130 -45 -115 -30
rect -65 -45 -50 -30
rect 92 -72 107 138
rect 162 -47 177 199
rect 419 192 441 207
rect 496 199 596 214
rect 511 168 551 178
rect 511 148 521 168
rect 541 148 551 168
rect 511 138 551 148
rect 419 87 441 106
rect 379 82 441 87
rect 379 62 389 82
rect 409 62 441 82
rect 379 57 441 62
rect 419 38 441 57
rect 419 -20 441 -5
rect 354 -45 369 -30
rect 77 -87 107 -72
rect 137 -57 177 -47
rect 137 -77 147 -57
rect 167 -77 177 -57
rect 137 -87 177 -77
rect 77 -102 92 -87
rect 511 -72 526 138
rect 581 -47 596 199
rect 838 192 860 207
rect 915 199 1015 214
rect 930 168 970 178
rect 930 148 940 168
rect 960 148 970 168
rect 930 138 970 148
rect 838 87 860 106
rect 798 82 860 87
rect 798 62 808 82
rect 828 62 860 82
rect 798 57 860 62
rect 838 38 860 57
rect 838 -20 860 -5
rect 773 -45 788 -30
rect 496 -87 526 -72
rect 556 -57 596 -47
rect 556 -77 566 -57
rect 586 -77 596 -57
rect 556 -87 596 -77
rect 496 -102 511 -87
rect 930 -72 945 138
rect 1000 -47 1015 199
rect 915 -87 945 -72
rect 975 -57 1015 -47
rect 975 -77 985 -57
rect 1005 -77 1015 -57
rect 975 -87 1015 -77
rect 915 -102 931 -87
rect -290 -162 -250 -152
rect -290 -182 -280 -162
rect -260 -182 -250 -162
rect -290 -192 -250 -182
rect -130 -213 -115 -145
rect -65 -213 -50 -145
rect 77 -160 92 -145
rect 354 -213 369 -145
rect 496 -160 511 -145
rect 773 -213 788 -145
rect 915 -160 931 -145
rect -339 -228 788 -213
<< polycont >>
rect -389 184 -369 204
rect 102 148 122 168
rect -30 62 -10 82
rect 521 148 541 168
rect 389 62 409 82
rect 147 -77 167 -57
rect 940 148 960 168
rect 808 62 828 82
rect 566 -77 586 -57
rect 985 -77 1005 -57
rect -280 -182 -260 -162
<< locali >>
rect -445 419 -405 429
rect -445 239 -435 419
rect -415 239 -405 419
rect -445 214 -405 239
rect -245 419 -205 429
rect -245 239 -235 419
rect -215 239 -205 419
rect -245 229 -205 239
rect -45 419 -5 429
rect -45 239 -35 419
rect -15 239 -5 419
rect 174 419 214 429
rect -45 229 -5 239
rect 32 305 72 315
rect 32 239 42 305
rect 62 239 72 305
rect 32 229 72 239
rect -445 204 -360 214
rect -445 184 -389 204
rect -369 184 -360 204
rect -445 174 -360 184
rect -45 209 72 229
rect 97 305 137 315
rect 97 239 107 305
rect 127 239 137 305
rect 97 229 137 239
rect 174 239 184 419
rect 204 239 214 419
rect 174 229 214 239
rect 374 419 414 429
rect 374 239 384 419
rect 404 239 414 419
rect 593 419 633 429
rect 374 229 414 239
rect 451 305 491 315
rect 451 239 461 305
rect 481 239 491 305
rect 451 229 491 239
rect -45 184 -5 209
rect -445 -5 -405 174
rect -45 116 -35 184
rect -15 116 -5 184
rect -45 106 -5 116
rect 27 184 67 192
rect 27 116 37 184
rect 57 116 67 184
rect 97 178 117 229
rect 374 209 491 229
rect 516 305 556 315
rect 516 239 526 305
rect 546 239 556 305
rect 516 229 556 239
rect 593 239 603 419
rect 623 239 633 419
rect 593 229 633 239
rect 793 419 833 429
rect 793 239 803 419
rect 823 239 833 419
rect 793 229 833 239
rect 870 305 910 315
rect 870 239 880 305
rect 900 239 910 305
rect 870 229 910 239
rect 374 184 414 209
rect 92 168 132 178
rect 92 148 102 168
rect 122 148 132 168
rect 92 138 132 148
rect -40 82 0 87
rect -40 62 -30 82
rect -10 62 0 82
rect -40 57 0 62
rect 27 82 67 116
rect 374 116 384 184
rect 404 116 414 184
rect 374 106 414 116
rect 446 184 486 192
rect 446 116 456 184
rect 476 116 486 184
rect 516 178 536 229
rect 793 209 910 229
rect 935 305 1025 315
rect 935 239 945 305
rect 965 239 995 305
rect 1015 239 1025 305
rect 935 229 1025 239
rect 793 184 833 209
rect 511 168 551 178
rect 511 148 521 168
rect 541 148 551 168
rect 511 138 551 148
rect 379 82 419 87
rect 27 62 389 82
rect 409 62 419 82
rect -45 30 -5 38
rect -45 5 -35 30
rect -15 5 -5 30
rect -445 -45 -135 -5
rect -45 -22 -5 5
rect 27 30 67 62
rect 379 57 419 62
rect 446 82 486 116
rect 793 116 803 184
rect 823 116 833 184
rect 793 106 833 116
rect 865 184 905 192
rect 865 116 875 184
rect 895 116 905 184
rect 935 178 955 229
rect 930 168 970 178
rect 930 148 940 168
rect 960 148 970 168
rect 930 138 970 148
rect 798 82 838 87
rect 446 62 808 82
rect 828 62 838 82
rect 27 5 37 30
rect 57 5 67 30
rect 27 -5 67 5
rect 374 30 414 38
rect 374 5 384 30
rect 404 5 414 30
rect 374 -5 414 5
rect 446 30 486 62
rect 798 57 838 62
rect 865 82 905 116
rect 865 62 1082 82
rect 446 5 456 30
rect 476 5 486 30
rect 446 -5 486 5
rect 793 30 833 38
rect 793 5 803 30
rect 823 5 833 30
rect 374 -22 415 -5
rect 793 -22 833 5
rect 865 30 905 62
rect 865 5 875 30
rect 895 5 905 30
rect 865 -5 905 5
rect -45 -42 72 -22
rect -175 -55 -135 -45
rect -175 -135 -165 -55
rect -145 -135 -135 -55
rect -175 -145 -135 -135
rect -110 -55 -70 -45
rect -110 -135 -100 -55
rect -80 -135 -70 -55
rect -110 -145 -70 -135
rect -45 -55 -5 -42
rect -45 -135 -35 -55
rect -15 -135 -5 -55
rect -45 -145 -5 -135
rect 32 -112 72 -42
rect 374 -42 491 -22
rect 137 -57 177 -47
rect 137 -77 147 -57
rect 167 -77 177 -57
rect 137 -102 177 -77
rect 259 -55 349 -45
rect 32 -135 42 -112
rect 62 -135 72 -112
rect 32 -145 72 -135
rect 97 -112 187 -102
rect 97 -135 107 -112
rect 127 -135 157 -112
rect 177 -135 187 -112
rect 97 -145 187 -135
rect 259 -135 269 -55
rect 289 -135 319 -55
rect 339 -135 349 -55
rect 259 -145 349 -135
rect 374 -55 414 -42
rect 374 -135 384 -55
rect 404 -135 414 -55
rect 374 -145 414 -135
rect 451 -112 491 -42
rect 793 -42 911 -22
rect 556 -57 596 -47
rect 556 -77 566 -57
rect 586 -77 596 -57
rect 556 -102 596 -77
rect 728 -55 768 -45
rect 451 -135 461 -112
rect 481 -135 491 -112
rect 451 -145 491 -135
rect 516 -112 606 -102
rect 516 -135 526 -112
rect 546 -135 576 -112
rect 596 -135 606 -112
rect 516 -145 606 -135
rect 728 -135 738 -55
rect 758 -135 768 -55
rect 728 -145 768 -135
rect 793 -55 833 -42
rect 793 -135 803 -55
rect 823 -135 833 -55
rect 793 -145 833 -135
rect 871 -112 911 -42
rect 975 -57 1015 -47
rect 975 -77 985 -57
rect 1005 -77 1015 -57
rect 975 -102 1015 -77
rect 871 -135 881 -112
rect 901 -135 911 -112
rect 871 -145 911 -135
rect 935 -112 1025 -102
rect 935 -135 945 -112
rect 966 -135 995 -112
rect 1015 -135 1025 -112
rect 935 -145 1025 -135
rect -290 -162 -250 -152
rect 1042 -162 1062 62
rect -290 -182 -280 -162
rect -260 -182 1062 -162
rect -290 -192 -250 -182
<< viali >>
rect -235 239 -215 419
rect 107 239 127 305
rect 184 239 204 419
rect 526 239 546 305
rect 603 239 623 419
rect 945 239 965 305
rect 995 239 1015 305
rect -100 -135 -80 -55
rect 107 -135 127 -112
rect 157 -135 177 -112
rect 269 -135 289 -55
rect 319 -135 339 -55
rect 526 -135 546 -112
rect 576 -135 596 -112
rect 738 -135 758 -55
rect 945 -135 966 -112
rect 995 -135 1015 -112
<< metal1 >>
rect -450 419 1054 429
rect -450 239 -235 419
rect -215 305 184 419
rect -215 239 107 305
rect 127 239 184 305
rect 204 305 603 419
rect 204 239 526 305
rect 546 239 603 305
rect 623 305 1054 419
rect 623 239 945 305
rect 965 239 995 305
rect 1015 239 1054 305
rect -450 229 1054 239
rect -180 -55 1062 -45
rect -180 -135 -100 -55
rect -80 -112 269 -55
rect -80 -135 107 -112
rect 127 -135 157 -112
rect 177 -135 269 -112
rect 289 -135 319 -55
rect 339 -112 738 -55
rect 339 -135 526 -112
rect 546 -135 576 -112
rect 596 -135 738 -112
rect 758 -112 1062 -55
rect 758 -135 945 -112
rect 966 -135 995 -112
rect 1015 -135 1062 -112
rect -180 -145 1062 -135
<< labels >>
flabel metal1 -450 329 -450 329 7 FreeSans 64 0 0 0 VDDA
port 1 w
flabel poly -339 -221 -339 -221 7 FreeSans 80 0 0 0 V_CONT
port 3 w
flabel locali 1082 71 1082 71 3 FreeSans 80 0 0 0 V_OSC
port 2 e
<< end >>
