** sch_path: /foss/designs/my_design/projects/mim_capacitor/xschem_ngspice/mimcap_1pF_xschem.sch
**.subckt mimcap_1pF_xschem
XC1 top bot sky130_fd_pr__cap_mim_m3_1 W=25 L=20 MF=1 m=1
**.ends
.end
