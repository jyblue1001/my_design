** sch_path: /foss/designs/projects/opamp/xschem_ngspice/vds_vgs_sweep_pfet.sch
**.subckt vds_vgs_sweep_pfet
VGS GND VGS 1.05
VDS GND VDS 1.8
XM1 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.6 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.3 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.15 W=104 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 VDS VGS GND GND sky130_fd_pr__pfet_01v8 L=0.2 W=35 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.option method=gear
.option wnflag=1
.option savecurrents
*.temp = 120

.save
+@m.xm1.msky130_fd_pr__pfet_01v8[gm]
+@m.xm2.msky130_fd_pr__pfet_01v8[gm]
+@m.xm3.msky130_fd_pr__pfet_01v8[gm]
+@m.xm4.msky130_fd_pr__pfet_01v8[gm]
+@m.xm5.msky130_fd_pr__pfet_01v8[gm]
+@m.xm6.msky130_fd_pr__pfet_01v8[gm]
+@m.xm7.msky130_fd_pr__pfet_01v8[gm]
+@m.xm8.msky130_fd_pr__pfet_01v8[gm]
+@m.xm9.msky130_fd_pr__pfet_01v8[gm]
+@m.xm10.msky130_fd_pr__pfet_01v8[gm]
+@m.xm1.msky130_fd_pr__pfet_01v8[gds]
+@m.xm2.msky130_fd_pr__pfet_01v8[gds]
+@m.xm2.msky130_fd_pr__pfet_01v8[vth]
+@m.xm3.msky130_fd_pr__pfet_01v8[gds]
+@m.xm4.msky130_fd_pr__pfet_01v8[gds]
+@m.xm5.msky130_fd_pr__pfet_01v8[gds]
+@m.xm6.msky130_fd_pr__pfet_01v8[gds]
+@m.xm7.msky130_fd_pr__pfet_01v8[gds]


.control
  save all
  * dc VGS 0 1.8 0.1 VDS 0 1.8 0.1
  * dc VDS 0 1.0 0.001 VGS 0.0 1.13 1.13
  dc VDS 0 0.6 0.001 VGS 0.8 1.1 0.01
  remzerovec
  write vds_vgs_sweep_pfet.raw
  set appendwrite
  let rout1 = deriv(vds)/deriv(@m.xm1.msky130_fd_pr__pfet_01v8[id])
  let rout2 = deriv(vds)/deriv(@m.xm2.msky130_fd_pr__pfet_01v8[id])
  let rout3 = deriv(vds)/deriv(@m.xm3.msky130_fd_pr__pfet_01v8[id])
  let rout4 = deriv(vds)/deriv(@m.xm4.msky130_fd_pr__pfet_01v8[id])
  let rout5 = deriv(vds)/deriv(@m.xm5.msky130_fd_pr__pfet_01v8[id])
  show
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
