* PEX produced on Sun Jun 22 03:49:02 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from ref_volt_cur_gen_dummy.ext - technology: sky130A

.subckt ref_volt_cur_gen_dummy VB1_CUR_BIAS GNDA ERR_AMP_REF VDDA VB2_CUR_BIAS VB3_CUR_BIAS
+ ERR_AMP_CUR_BIAS V_CMFB_S2 TAIL_CUR_MIR_BIAS V_CMFB_S1 V_CMFB_S4 V_CMFB_S3
X0 VDDA.t213 VDDA.t211 V_CMFB_S1.t5 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X1 VDDA.t117 V_TOP.t14 Vin+.t5 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X2 GNDA.t110 VDDA.t214 V_p_1.t10 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X3 VDDA.t28 PFET_GATE_10uA.t10 TAIL_CUR_MIR_BIAS.t7 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X4 VDDA.t210 VDDA.t208 V_TOP.t13 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X5 1st_Vout_1.t11 cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t90 GNDA.t88 VB3_CUR_BIAS.t4 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X7 1st_Vout_2.t11 cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VDDA.t32 V_TOP.t15 START_UP.t3 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X9 V_mir2.t16 V_mir2.t15 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X10 GNDA.t68 GNDA.t93 Vbe2.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X11 GNDA.t31 a_4400_6480.t0 GNDA.t30 sky130_fd_pr__res_xhigh_po_0p35 l=6
X12 VDDA.t128 V_mir2.t13 V_mir2.t14 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X13 VB2_CUR_BIAS.t7 NFET_GATE_10uA.t5 GNDA.t29 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X14 GNDA.t72 GNDA.t92 Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X15 a_2792_6360.t1 a_4400_6480.t1 GNDA.t5 sky130_fd_pr__res_xhigh_po_0p35 l=6
X16 1st_Vout_1.t12 cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 GNDA.t50 START_UP_NFET1.t1 START_UP_NFET1.t0 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X18 V_TOP.t1 START_UP.t6 Vin-.t7 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X19 TAIL_CUR_MIR_BIAS.t6 PFET_GATE_10uA.t11 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X20 VB1_CUR_BIAS.t1 PFET_GATE_10uA.t12 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X21 1st_Vout_2.t12 cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 GNDA.t70 GNDA.t91 Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X23 VB2_CUR_BIAS.t6 NFET_GATE_10uA.t6 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X24 VDDA.t49 V_mir2.t17 1st_Vout_2.t6 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X25 1st_Vout_2.t8 V_CUR_REF_REG.t3 V_p_2.t9 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X26 1st_Vout_1.t13 cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 VB2_CUR_BIAS.t5 NFET_GATE_10uA.t7 GNDA.t25 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X28 Vin-.t4 V_TOP.t16 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X29 1st_Vout_2.t13 cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 TAIL_CUR_MIR_BIAS.t5 PFET_GATE_10uA.t13 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X31 VDDA.t207 VDDA.t205 PFET_GATE_10uA.t9 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X32 V_TOP.t5 1st_Vout_1.t14 VDDA.t115 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X33 1st_Vout_1.t15 cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 V_TOP.t12 VDDA.t202 VDDA.t204 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X35 ERR_AMP_REF.t4 V_TOP.t17 VDDA.t152 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X36 V_TOP.t18 VDDA.t158 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 1st_Vout_2.t14 cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 1st_Vout_1.t16 cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 NFET_GATE_10uA.t0 GNDA.t94 GNDA.t96 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X40 V_mir2.t0 ERR_AMP_REF.t7 V_p_2.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X41 V_TOP.t19 VDDA.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 GNDA.t87 GNDA.t85 VB2_CUR_BIAS.t1 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X43 VDDA.t109 V_mir2.t11 V_mir2.t12 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X44 PFET_GATE_10uA.t6 1st_Vout_2.t15 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X45 1st_Vout_2.t16 cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 V_TOP.t20 VDDA.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 GNDA.t42 NFET_GATE_10uA.t8 VB2_CUR_BIAS.t4 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X48 VB3_CUR_BIAS.t1 NFET_GATE_10uA.t9 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X49 VDDA.t113 V_mir1.t17 1st_Vout_1.t4 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 V_p_1.t8 Vin+.t6 1st_Vout_1.t10 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X51 V_p_2.t3 ERR_AMP_REF.t8 V_mir2.t3 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X52 VDDA.t65 PFET_GATE_10uA.t14 TAIL_CUR_MIR_BIAS.t4 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X53 VDDA.t136 V_TOP.t21 Vin-.t3 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X54 V_TOP.t22 VDDA.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VDDA.t84 1st_Vout_1.t17 V_TOP.t2 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X56 1st_Vout_2.t17 cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 VB2_CUR_BIAS.t0 GNDA.t82 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X58 VDDA.t15 V_TOP.t23 START_UP.t2 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X59 V_p_1.t2 Vin-.t8 V_mir1.t16 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X60 V_TOP.t9 VDDA.t215 GNDA.t109 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X61 V_p_2.t8 V_CUR_REF_REG.t4 1st_Vout_2.t3 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X62 VDDA.t201 VDDA.t199 ERR_AMP_REF.t6 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X63 V_TOP.t24 VDDA.t146 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 GNDA.t68 GNDA.t73 Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X65 1st_Vout_2.t18 cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 GNDA.t72 GNDA.t71 Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X67 VDDA.t145 1st_Vout_1.t18 V_TOP.t7 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X68 V_CMFB_S1.t1 PFET_GATE_10uA.t15 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X69 1st_Vout_1.t19 cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 V_p_1.t6 Vin+.t7 1st_Vout_1.t9 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X71 GNDA.t106 NFET_GATE_10uA.t10 VB3_CUR_BIAS.t5 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X72 VDDA.t157 1st_Vout_1.t20 V_TOP.t8 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X73 V_TOP.t25 VDDA.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 V_CMFB_S4.t3 NFET_GATE_10uA.t11 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X75 V_p_2.t4 ERR_AMP_REF.t9 V_mir2.t4 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X76 V_TOP.t11 VDDA.t196 VDDA.t198 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X77 V_CUR_REF_REG.t1 PFET_GATE_10uA.t16 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X78 V_mir2.t10 V_mir2.t9 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 GNDA.t108 VDDA.t216 PFET_GATE_10uA.t7 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X80 1st_Vout_1.t21 cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 PFET_GATE_10uA.t4 1st_Vout_2.t19 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X82 1st_Vout_2.t20 cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 GNDA.t54 NFET_GATE_10uA.t12 VB2_CUR_BIAS.t3 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X84 VDDA.t91 PFET_GATE_10uA.t17 V_CMFB_S3.t3 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X85 NFET_GATE_10uA.t4 VDDA.t169 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X86 Vin-.t2 V_TOP.t26 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X87 V_mir1.t15 Vin-.t9 V_p_1.t4 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X88 1st_Vout_2.t5 V_CUR_REF_REG.t5 V_p_2.t7 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X89 1st_Vout_1.t22 cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 1st_Vout_2.t21 cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 1st_Vout_2.t22 cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 V_mir1.t11 V_mir1.t10 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X93 ERR_AMP_REF.t3 V_TOP.t27 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X94 1st_Vout_1.t8 Vin+.t8 V_p_1.t5 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X95 VDDA.t161 PFET_GATE_10uA.t18 V_CMFB_S1.t3 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X96 1st_Vout_1.t23 cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 GNDA.t18 a_1830_6460.t0 GNDA.t17 sky130_fd_pr__res_xhigh_po_0p35 l=6
X98 VDDA.t195 VDDA.t193 VB1_CUR_BIAS.t3 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X99 GNDA.t81 GNDA.t79 V_CMFB_S4.t0 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X100 V_mir1.t9 V_mir1.t8 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X101 1st_Vout_1.t7 Vin+.t9 V_p_1.t9 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X102 1st_Vout_2.t23 cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 V_CMFB_S3.t2 PFET_GATE_10uA.t19 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X104 V_TOP.t28 VDDA.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 V_CMFB_S4.t2 NFET_GATE_10uA.t13 GNDA.t58 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X106 V_mir1.t7 V_mir1.t6 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X107 V_mir1.t14 Vin-.t10 V_p_1.t3 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X108 1st_Vout_2.t7 V_CUR_REF_REG.t6 V_p_2.t6 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X109 VDDA.t101 PFET_GATE_10uA.t20 NFET_GATE_10uA.t1 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X110 GNDA.t100 NFET_GATE_10uA.t14 VB2_CUR_BIAS.t2 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X111 VDDA.t17 V_mir2.t7 V_mir2.t8 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X112 1st_Vout_2.t24 cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 V_TOP.t29 VDDA.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 V_CUR_REF_REG.t0 a_1830_6460.t1 GNDA.t32 sky130_fd_pr__res_xhigh_po_0p35 l=6
X115 V_TOP.t30 VDDA.t159 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VDDA.t174 VDDA.t172 V_TOP.t10 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X117 VDDA.t86 V_TOP.t31 ERR_AMP_REF.t2 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X118 VDDA.t61 PFET_GATE_10uA.t21 TAIL_CUR_MIR_BIAS.t3 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X119 V_p_1.t0 Vin-.t11 V_mir1.t13 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X120 1st_Vout_2.t25 cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 1st_Vout_2.t26 cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 GNDA.t11 NFET_GATE_10uA.t2 NFET_GATE_10uA.t3 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X123 1st_Vout_1.t3 V_mir1.t18 VDDA.t111 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X124 cap_res1.t0 V_TOP.t6 GNDA.t59 sky130_fd_pr__res_high_po_0p35 l=2.05
X125 VDDA.t89 V_mir1.t4 V_mir1.t5 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X126 1st_Vout_1.t24 cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 V_CMFB_S2.t0 GNDA.t76 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X128 1st_Vout_2.t2 V_mir2.t18 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X129 V_TOP.t32 VDDA.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VDDA.t107 PFET_GATE_10uA.t22 V_CMFB_S3.t1 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X131 ERR_AMP_REF.t5 VDDA.t190 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X132 VDDA.t96 V_mir1.t2 V_mir1.t3 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X133 V_p_1.t7 Vin+.t10 1st_Vout_1.t6 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X134 1st_Vout_1.t25 cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 V_p_2.t10 VDDA.t217 GNDA.t107 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X136 Vin-.t6 START_UP.t7 V_TOP.t3 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X137 V_TOP.t33 VDDA.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 V_CMFB_S2.t3 NFET_GATE_10uA.t15 GNDA.t102 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X139 GNDA.t70 GNDA.t75 Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X140 PFET_GATE_10uA.t8 VDDA.t187 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X141 V_p_2.t5 V_CUR_REF_REG.t7 1st_Vout_2.t9 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X142 1st_Vout_1.t26 cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 TAIL_CUR_MIR_BIAS.t2 PFET_GATE_10uA.t23 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X144 VDDA.t13 V_mir1.t0 V_mir1.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X145 V_TOP.t34 VDDA.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 1st_Vout_2.t27 cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 V_TOP.t35 VDDA.t153 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 ERR_AMP_CUR_BIAS.t1 NFET_GATE_10uA.t16 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X149 PFET_GATE_10uA.t0 1st_Vout_2.t28 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X150 VDDA.t139 1st_Vout_2.t29 PFET_GATE_10uA.t3 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X151 START_UP.t1 V_TOP.t36 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X152 VDDA.t11 V_mir1.t19 1st_Vout_1.t2 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X153 1st_Vout_1.t27 cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 1st_Vout_1.t28 cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VB3_CUR_BIAS.t3 NFET_GATE_10uA.t17 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X156 VDDA.t74 V_TOP.t37 ERR_AMP_REF.t1 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X157 V_CMFB_S3.t0 PFET_GATE_10uA.t24 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X158 VDDA.t130 V_mir1.t20 1st_Vout_1.t5 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X159 1st_Vout_1.t0 V_mir1.t21 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X160 GNDA.t48 NFET_GATE_10uA.t18 V_CMFB_S2.t2 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X161 VDDA.t82 V_TOP.t38 Vin-.t1 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X162 VDDA.t3 V_mir2.t19 1st_Vout_2.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X163 1st_Vout_1.t29 cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 1st_Vout_2.t30 cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 V_mir1.t12 Vin-.t12 V_p_1.t1 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X166 GNDA.t46 NFET_GATE_10uA.t19 ERR_AMP_CUR_BIAS.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X167 cap_res2.t0 PFET_GATE_10uA.t2 GNDA.t59 sky130_fd_pr__res_high_po_0p35 l=2.05
X168 Vbe2.t0 Vin+.t0 GNDA.t37 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X169 1st_Vout_1.t1 V_mir1.t22 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 V_TOP.t39 VDDA.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VDDA.t122 1st_Vout_2.t31 PFET_GATE_10uA.t1 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X172 1st_Vout_2.t32 cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 1st_Vout_2.t33 cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 V_mir2.t2 ERR_AMP_REF.t10 V_p_2.t2 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X175 VDDA.t186 VDDA.t184 V_CUR_REF_REG.t2 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X176 GNDA.t44 NFET_GATE_10uA.t20 VB3_CUR_BIAS.t2 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X177 START_UP.t0 V_TOP.t40 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X178 GNDA.t68 GNDA.t67 Vin-.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X179 VDDA.t183 VDDA.t181 V_CMFB_S3.t5 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.5
X180 GNDA.t72 GNDA.t74 Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X181 VDDA.t163 1st_Vout_2.t34 PFET_GATE_10uA.t5 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X182 V_CMFB_S1.t4 VDDA.t178 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X183 V_TOP.t4 1st_Vout_1.t30 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X184 1st_Vout_2.t35 cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 GNDA.t61 NFET_GATE_10uA.t21 V_CMFB_S4.t1 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X186 GNDA.t70 GNDA.t69 Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X187 Vin+.t4 V_TOP.t41 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X188 1st_Vout_1.t31 cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 TAIL_CUR_MIR_BIAS.t1 PFET_GATE_10uA.t25 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X190 V_CMFB_S3.t4 VDDA.t175 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X191 VB1_CUR_BIAS.t2 VDDA.t166 VDDA.t168 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.5
X192 ERR_AMP_REF.t0 a_1890_6990.t1 GNDA.t16 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X193 V_TOP.t42 VDDA.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 V_CMFB_S1.t2 PFET_GATE_10uA.t26 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X195 V_TOP.t0 1st_Vout_1.t32 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X196 VDDA.t34 V_mir2.t20 1st_Vout_2.t4 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X197 1st_Vout_1.t33 cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 1st_Vout_1.t34 cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 START_UP_NFET1.t0 START_UP.t4 START_UP.t5 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X200 a_2792_6240.t0 a_4400_6600.t0 GNDA.t8 sky130_fd_pr__res_xhigh_po_0p35 l=6
X201 Vin+.t3 V_TOP.t43 VDDA.t120 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X202 V_mir2.t6 V_mir2.t5 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X203 a_2792_6240.t1 Vin+.t1 GNDA.t5 sky130_fd_pr__res_xhigh_po_0p35 l=6
X204 V_TOP.t44 VDDA.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 V_TOP.t45 VDDA.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 VB3_CUR_BIAS.t0 NFET_GATE_10uA.t22 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X207 V_TOP.t46 VDDA.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 1st_Vout_1.t35 cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 1st_Vout_1.t36 cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 GNDA.t36 NFET_GATE_10uA.t23 V_CMFB_S2.t1 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X211 1st_Vout_2.t10 V_mir2.t21 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X212 V_TOP.t47 VDDA.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 VDDA.t67 PFET_GATE_10uA.t27 V_CMFB_S1.t0 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X214 V_p_2.t1 ERR_AMP_REF.t11 V_mir2.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X215 VDDA.t42 V_TOP.t48 Vin+.t2 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X216 1st_Vout_2.t36 cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 V_TOP.t49 VDDA.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 GNDA.t20 a_4400_6600.t1 GNDA.t19 sky130_fd_pr__res_xhigh_po_0p35 l=6
X219 VDDA.t71 PFET_GATE_10uA.t28 TAIL_CUR_MIR_BIAS.t0 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X220 VDDA.t76 PFET_GATE_10uA.t29 VB1_CUR_BIAS.t0 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.5
X221 GNDA.t7 a_1890_6990.t0 GNDA.t6 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X222 a_2792_6360.t0 Vin-.t0 GNDA.t5 sky130_fd_pr__res_xhigh_po_0p35 l=6
X223 1st_Vout_2.t1 V_mir2.t22 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 VDDA.n121 VDDA.n117 6600
R1 VDDA.n121 VDDA.n118 6600
R2 VDDA.n123 VDDA.n117 6570
R3 VDDA.n123 VDDA.n118 6570
R4 VDDA.n66 VDDA.n13 4710
R5 VDDA.n66 VDDA.n14 4710
R6 VDDA.n64 VDDA.n13 4710
R7 VDDA.n64 VDDA.n14 4710
R8 VDDA.n42 VDDA.n35 4710
R9 VDDA.n44 VDDA.n35 4710
R10 VDDA.n42 VDDA.n41 4710
R11 VDDA.n44 VDDA.n41 4710
R12 VDDA.n188 VDDA.n182 4350
R13 VDDA.n188 VDDA.n183 4350
R14 VDDA.n186 VDDA.n182 4350
R15 VDDA.n186 VDDA.n183 4350
R16 VDDA.n202 VDDA.n196 2730
R17 VDDA.n202 VDDA.n197 2730
R18 VDDA.n200 VDDA.n196 2730
R19 VDDA.n200 VDDA.n197 2730
R20 VDDA.n174 VDDA.n168 2730
R21 VDDA.n174 VDDA.n169 2730
R22 VDDA.n172 VDDA.n168 2730
R23 VDDA.n172 VDDA.n169 2730
R24 VDDA.n136 VDDA.n131 2190
R25 VDDA.n138 VDDA.n131 2190
R26 VDDA.n136 VDDA.n134 2190
R27 VDDA.n138 VDDA.n134 2190
R28 VDDA.n108 VDDA.n103 1770
R29 VDDA.n110 VDDA.n103 1770
R30 VDDA.n108 VDDA.n106 1770
R31 VDDA.n110 VDDA.n106 1770
R32 VDDA.n120 VDDA.n119 704
R33 VDDA.n120 VDDA.n86 704
R34 VDDA.n125 VDDA.n124 518.4
R35 VDDA.n124 VDDA.n116 518.4
R36 VDDA.n46 VDDA.n45 496
R37 VDDA.n46 VDDA.n34 496
R38 VDDA.n185 VDDA.n184 464
R39 VDDA.n185 VDDA.n152 464
R40 VDDA.n101 VDDA.t172 413.084
R41 VDDA.n104 VDDA.t202 413.084
R42 VDDA.t182 VDDA.n196 394.774
R43 VDDA.t176 VDDA.n197 394.774
R44 VDDA.t194 VDDA.n136 394.774
R45 VDDA.n138 VDDA.t167 394.774
R46 VDDA.t185 VDDA.n182 390.262
R47 VDDA.t170 VDDA.n183 390.262
R48 VDDA.t212 VDDA.n168 390.262
R49 VDDA.t179 VDDA.n169 390.262
R50 VDDA.n129 VDDA.t195 389.185
R51 VDDA.n132 VDDA.t168 389.185
R52 VDDA.n205 VDDA.t183 387.051
R53 VDDA.n194 VDDA.t177 387.051
R54 VDDA.n191 VDDA.t186 387.051
R55 VDDA.n180 VDDA.t171 387.051
R56 VDDA.n177 VDDA.t213 387.051
R57 VDDA.n166 VDDA.t180 387.051
R58 VDDA.n101 VDDA.t174 384.918
R59 VDDA.n104 VDDA.t204 384.918
R60 VDDA.n15 VDDA.t207 384.918
R61 VDDA.n17 VDDA.t189 384.918
R62 VDDA.n38 VDDA.t210 384.918
R63 VDDA.n36 VDDA.t198 384.918
R64 VDDA.n63 VDDA.n16 384
R65 VDDA.n63 VDDA.n62 384
R66 VDDA.n40 VDDA.n39 384
R67 VDDA.n40 VDDA.n37 384
R68 VDDA.n115 VDDA.t190 360.868
R69 VDDA.n126 VDDA.t199 360.868
R70 VDDA.n15 VDDA.t205 358.858
R71 VDDA.n17 VDDA.t187 358.858
R72 VDDA.n38 VDDA.t208 358.858
R73 VDDA.n36 VDDA.t196 358.858
R74 VDDA.t206 VDDA.n13 351.591
R75 VDDA.t188 VDDA.n14 351.591
R76 VDDA.t209 VDDA.n42 351.591
R77 VDDA.n44 VDDA.t197 351.591
R78 VDDA.n190 VDDA.n189 345.601
R79 VDDA.n189 VDDA.n181 345.601
R80 VDDA.t173 VDDA.n108 344.394
R81 VDDA.n110 VDDA.t203 344.394
R82 VDDA.n29 VDDA.n27 342.301
R83 VDDA.n57 VDDA.n56 341.676
R84 VDDA.n55 VDDA.n54 341.676
R85 VDDA.n53 VDDA.n52 341.676
R86 VDDA.n51 VDDA.n50 341.676
R87 VDDA.n33 VDDA.n32 341.676
R88 VDDA.n31 VDDA.n30 341.676
R89 VDDA.n29 VDDA.n28 341.676
R90 VDDA.n146 VDDA.n145 339.272
R91 VDDA.n149 VDDA.n148 339.272
R92 VDDA.n151 VDDA.n150 339.272
R93 VDDA.n154 VDDA.n153 339.272
R94 VDDA.n156 VDDA.n155 339.272
R95 VDDA.n158 VDDA.n157 339.272
R96 VDDA.n160 VDDA.n159 339.272
R97 VDDA.n162 VDDA.n161 339.272
R98 VDDA.n165 VDDA.n164 339.272
R99 VDDA.n25 VDDA.n24 337.176
R100 VDDA.n22 VDDA.n20 337.176
R101 VDDA.n11 VDDA.n10 337.176
R102 VDDA.n68 VDDA.n9 337.176
R103 VDDA.n71 VDDA.n70 337.176
R104 VDDA.n75 VDDA.n74 337.176
R105 VDDA.n78 VDDA.n77 337.176
R106 VDDA.n81 VDDA.n5 337.176
R107 VDDA.n59 VDDA.n19 337.176
R108 VDDA.n48 VDDA.n47 337.176
R109 VDDA.n142 VDDA.n128 335.022
R110 VDDA.n199 VDDA.n198 291.2
R111 VDDA.n199 VDDA.n147 291.2
R112 VDDA.n171 VDDA.n170 291.2
R113 VDDA.n171 VDDA.n163 291.2
R114 VDDA.t200 VDDA.n117 278.95
R115 VDDA.t191 VDDA.n118 278.95
R116 VDDA.n129 VDDA.t193 274.509
R117 VDDA.n132 VDDA.t166 274.509
R118 VDDA.n126 VDDA.t201 270.705
R119 VDDA.n115 VDDA.t192 270.705
R120 VDDA.n194 VDDA.t175 264.467
R121 VDDA.n205 VDDA.t181 264.467
R122 VDDA.n180 VDDA.t169 264.467
R123 VDDA.n191 VDDA.t184 264.467
R124 VDDA.n166 VDDA.t178 264.467
R125 VDDA.n177 VDDA.t211 264.467
R126 VDDA.t35 VDDA.t182 259.091
R127 VDDA.t106 VDDA.t35 259.091
R128 VDDA.t0 VDDA.t90 259.091
R129 VDDA.t90 VDDA.t176 259.091
R130 VDDA.t102 VDDA.t194 259.091
R131 VDDA.t167 VDDA.t75 259.091
R132 VDDA.t154 VDDA.t185 255.225
R133 VDDA.t64 VDDA.t154 255.225
R134 VDDA.t62 VDDA.t64 255.225
R135 VDDA.t27 VDDA.t62 255.225
R136 VDDA.t77 VDDA.t27 255.225
R137 VDDA.t60 VDDA.t22 255.225
R138 VDDA.t22 VDDA.t70 255.225
R139 VDDA.t70 VDDA.t20 255.225
R140 VDDA.t20 VDDA.t100 255.225
R141 VDDA.t100 VDDA.t170 255.225
R142 VDDA.t149 VDDA.t212 255.225
R143 VDDA.t160 VDDA.t149 255.225
R144 VDDA.t142 VDDA.t66 255.225
R145 VDDA.t66 VDDA.t179 255.225
R146 VDDA.n139 VDDA.n133 233.601
R147 VDDA.n135 VDDA.n133 233.601
R148 VDDA.n111 VDDA.n105 188.8
R149 VDDA.n107 VDDA.n105 188.8
R150 VDDA.n61 VDDA.n60 188.8
R151 VDDA.n80 VDDA.n6 188.8
R152 VDDA.n119 VDDA.n116 182.4
R153 VDDA.n125 VDDA.n86 182.4
R154 VDDA.n204 VDDA.n203 172.8
R155 VDDA.n203 VDDA.n195 172.8
R156 VDDA.n176 VDDA.n175 172.8
R157 VDDA.n175 VDDA.n167 172.8
R158 VDDA.t164 VDDA.t206 172.727
R159 VDDA.t127 VDDA.t164 172.727
R160 VDDA.t123 VDDA.t127 172.727
R161 VDDA.t2 VDDA.t123 172.727
R162 VDDA.t18 VDDA.t2 172.727
R163 VDDA.t138 VDDA.t18 172.727
R164 VDDA.t140 VDDA.t138 172.727
R165 VDDA.t108 VDDA.t140 172.727
R166 VDDA.t92 VDDA.t108 172.727
R167 VDDA.t33 VDDA.t6 172.727
R168 VDDA.t6 VDDA.t162 172.727
R169 VDDA.t162 VDDA.t50 172.727
R170 VDDA.t50 VDDA.t16 172.727
R171 VDDA.t16 VDDA.t125 172.727
R172 VDDA.t125 VDDA.t48 172.727
R173 VDDA.t48 VDDA.t147 172.727
R174 VDDA.t147 VDDA.t121 172.727
R175 VDDA.t121 VDDA.t188 172.727
R176 VDDA.t29 VDDA.t209 172.727
R177 VDDA.t129 VDDA.t29 172.727
R178 VDDA.t110 VDDA.t129 172.727
R179 VDDA.t12 VDDA.t110 172.727
R180 VDDA.t58 VDDA.t12 172.727
R181 VDDA.t156 VDDA.t58 172.727
R182 VDDA.t104 VDDA.t156 172.727
R183 VDDA.t10 VDDA.t104 172.727
R184 VDDA.t8 VDDA.t10 172.727
R185 VDDA.t56 VDDA.t95 172.727
R186 VDDA.t144 VDDA.t56 172.727
R187 VDDA.t114 VDDA.t144 172.727
R188 VDDA.t112 VDDA.t114 172.727
R189 VDDA.t4 VDDA.t112 172.727
R190 VDDA.t88 VDDA.t4 172.727
R191 VDDA.t133 VDDA.t88 172.727
R192 VDDA.t83 VDDA.t133 172.727
R193 VDDA.t197 VDDA.t83 172.727
R194 VDDA.n85 VDDA.n84 168.435
R195 VDDA.n88 VDDA.n87 168.435
R196 VDDA.n90 VDDA.n89 168.435
R197 VDDA.n92 VDDA.n91 168.435
R198 VDDA.n94 VDDA.n93 168.435
R199 VDDA.n96 VDDA.n95 168.435
R200 VDDA.n98 VDDA.n97 168.435
R201 VDDA.n100 VDDA.n99 168.435
R202 VDDA.t151 VDDA.t200 159.814
R203 VDDA.t31 VDDA.t151 159.814
R204 VDDA.t68 VDDA.t31 159.814
R205 VDDA.t135 VDDA.t68 159.814
R206 VDDA.t24 VDDA.t135 159.814
R207 VDDA.t116 VDDA.t24 159.814
R208 VDDA.t119 VDDA.t116 159.814
R209 VDDA.t85 VDDA.t119 159.814
R210 VDDA.t44 VDDA.t41 159.814
R211 VDDA.t41 VDDA.t54 159.814
R212 VDDA.t54 VDDA.t81 159.814
R213 VDDA.t81 VDDA.t52 159.814
R214 VDDA.t52 VDDA.t14 159.814
R215 VDDA.t14 VDDA.t38 159.814
R216 VDDA.t38 VDDA.t73 159.814
R217 VDDA.t73 VDDA.t191 159.814
R218 VDDA.t43 VDDA.t173 158.333
R219 VDDA.t203 VDDA.t94 158.333
R220 VDDA.n201 VDDA.t106 129.546
R221 VDDA.n201 VDDA.t0 129.546
R222 VDDA.n137 VDDA.t102 129.546
R223 VDDA.t75 VDDA.n137 129.546
R224 VDDA.n187 VDDA.t77 127.612
R225 VDDA.n187 VDDA.t60 127.612
R226 VDDA.n173 VDDA.t160 127.612
R227 VDDA.n173 VDDA.t142 127.612
R228 VDDA.n198 VDDA.n195 118.4
R229 VDDA.n204 VDDA.n147 118.4
R230 VDDA.n184 VDDA.n181 118.4
R231 VDDA.n190 VDDA.n152 118.4
R232 VDDA.n170 VDDA.n167 118.4
R233 VDDA.n176 VDDA.n163 118.4
R234 VDDA.n140 VDDA.n139 118.4
R235 VDDA.n135 VDDA.n130 118.4
R236 VDDA.n112 VDDA.n111 118.4
R237 VDDA.n107 VDDA.n102 118.4
R238 VDDA.n62 VDDA.n61 118.4
R239 VDDA.n16 VDDA.n6 118.4
R240 VDDA.n45 VDDA.n37 118.4
R241 VDDA.n39 VDDA.n34 118.4
R242 VDDA.n141 VDDA.n140 107.52
R243 VDDA.n141 VDDA.n130 107.52
R244 VDDA.n198 VDDA.n197 92.5005
R245 VDDA.n200 VDDA.n199 92.5005
R246 VDDA.n201 VDDA.n200 92.5005
R247 VDDA.n196 VDDA.n147 92.5005
R248 VDDA.n203 VDDA.n202 92.5005
R249 VDDA.n202 VDDA.n201 92.5005
R250 VDDA.n184 VDDA.n183 92.5005
R251 VDDA.n186 VDDA.n185 92.5005
R252 VDDA.n187 VDDA.n186 92.5005
R253 VDDA.n182 VDDA.n152 92.5005
R254 VDDA.n189 VDDA.n188 92.5005
R255 VDDA.n188 VDDA.n187 92.5005
R256 VDDA.n170 VDDA.n169 92.5005
R257 VDDA.n172 VDDA.n171 92.5005
R258 VDDA.n173 VDDA.n172 92.5005
R259 VDDA.n168 VDDA.n163 92.5005
R260 VDDA.n175 VDDA.n174 92.5005
R261 VDDA.n174 VDDA.n173 92.5005
R262 VDDA.n139 VDDA.n138 92.5005
R263 VDDA.n136 VDDA.n135 92.5005
R264 VDDA.n119 VDDA.n118 92.5005
R265 VDDA.n121 VDDA.n120 92.5005
R266 VDDA.n122 VDDA.n121 92.5005
R267 VDDA.n117 VDDA.n86 92.5005
R268 VDDA.n124 VDDA.n123 92.5005
R269 VDDA.n123 VDDA.n122 92.5005
R270 VDDA.n111 VDDA.n110 92.5005
R271 VDDA.n106 VDDA.n105 92.5005
R272 VDDA.n109 VDDA.n106 92.5005
R273 VDDA.n108 VDDA.n107 92.5005
R274 VDDA.n113 VDDA.n103 92.5005
R275 VDDA.n109 VDDA.n103 92.5005
R276 VDDA.n61 VDDA.n14 92.5005
R277 VDDA.n64 VDDA.n63 92.5005
R278 VDDA.n65 VDDA.n64 92.5005
R279 VDDA.n13 VDDA.n6 92.5005
R280 VDDA.n67 VDDA.n66 92.5005
R281 VDDA.n66 VDDA.n65 92.5005
R282 VDDA.n45 VDDA.n44 92.5005
R283 VDDA.n41 VDDA.n40 92.5005
R284 VDDA.n43 VDDA.n41 92.5005
R285 VDDA.n42 VDDA.n34 92.5005
R286 VDDA.n46 VDDA.n35 92.5005
R287 VDDA.n43 VDDA.n35 92.5005
R288 VDDA.n65 VDDA.t92 86.3641
R289 VDDA.n65 VDDA.t33 86.3641
R290 VDDA.n43 VDDA.t8 86.3641
R291 VDDA.t95 VDDA.n43 86.3641
R292 VDDA.n122 VDDA.t85 79.907
R293 VDDA.n122 VDDA.t44 79.907
R294 VDDA.n109 VDDA.t43 79.1672
R295 VDDA.t94 VDDA.n109 79.1672
R296 VDDA.n113 VDDA.n112 64.0005
R297 VDDA.n113 VDDA.n102 64.0005
R298 VDDA.n80 VDDA.n79 64.0005
R299 VDDA.n79 VDDA.n76 64.0005
R300 VDDA.n76 VDDA.n7 64.0005
R301 VDDA.n67 VDDA.n7 64.0005
R302 VDDA.n67 VDDA.n12 64.0005
R303 VDDA.n21 VDDA.n12 64.0005
R304 VDDA.n21 VDDA.n18 64.0005
R305 VDDA.n60 VDDA.n18 64.0005
R306 VDDA.n0 VDDA.t215 59.5681
R307 VDDA.n1 VDDA.t216 59.5681
R308 VDDA.n0 VDDA.t214 51.8887
R309 VDDA.n2 VDDA.t217 48.9557
R310 VDDA.n134 VDDA.n133 46.2505
R311 VDDA.n137 VDDA.n134 46.2505
R312 VDDA.n141 VDDA.n131 46.2505
R313 VDDA.n137 VDDA.n131 46.2505
R314 VDDA.n145 VDDA.t36 39.4005
R315 VDDA.n145 VDDA.t107 39.4005
R316 VDDA.n148 VDDA.t1 39.4005
R317 VDDA.n148 VDDA.t91 39.4005
R318 VDDA.n150 VDDA.t155 39.4005
R319 VDDA.n150 VDDA.t65 39.4005
R320 VDDA.n153 VDDA.t63 39.4005
R321 VDDA.n153 VDDA.t28 39.4005
R322 VDDA.n155 VDDA.t78 39.4005
R323 VDDA.n155 VDDA.t61 39.4005
R324 VDDA.n157 VDDA.t23 39.4005
R325 VDDA.n157 VDDA.t71 39.4005
R326 VDDA.n159 VDDA.t21 39.4005
R327 VDDA.n159 VDDA.t101 39.4005
R328 VDDA.n161 VDDA.t150 39.4005
R329 VDDA.n161 VDDA.t161 39.4005
R330 VDDA.n164 VDDA.t143 39.4005
R331 VDDA.n164 VDDA.t67 39.4005
R332 VDDA.n128 VDDA.t103 39.4005
R333 VDDA.n128 VDDA.t76 39.4005
R334 VDDA.n24 VDDA.t126 39.4005
R335 VDDA.n24 VDDA.t49 39.4005
R336 VDDA.n20 VDDA.t51 39.4005
R337 VDDA.n20 VDDA.t17 39.4005
R338 VDDA.n10 VDDA.t7 39.4005
R339 VDDA.n10 VDDA.t163 39.4005
R340 VDDA.n9 VDDA.t93 39.4005
R341 VDDA.n9 VDDA.t34 39.4005
R342 VDDA.n70 VDDA.t141 39.4005
R343 VDDA.n70 VDDA.t109 39.4005
R344 VDDA.n74 VDDA.t19 39.4005
R345 VDDA.n74 VDDA.t139 39.4005
R346 VDDA.n77 VDDA.t124 39.4005
R347 VDDA.n77 VDDA.t3 39.4005
R348 VDDA.n5 VDDA.t165 39.4005
R349 VDDA.n5 VDDA.t128 39.4005
R350 VDDA.n19 VDDA.t148 39.4005
R351 VDDA.n19 VDDA.t122 39.4005
R352 VDDA.n56 VDDA.t30 39.4005
R353 VDDA.n56 VDDA.t130 39.4005
R354 VDDA.n54 VDDA.t111 39.4005
R355 VDDA.n54 VDDA.t13 39.4005
R356 VDDA.n52 VDDA.t59 39.4005
R357 VDDA.n52 VDDA.t157 39.4005
R358 VDDA.n50 VDDA.t105 39.4005
R359 VDDA.n50 VDDA.t11 39.4005
R360 VDDA.n47 VDDA.t9 39.4005
R361 VDDA.n47 VDDA.t96 39.4005
R362 VDDA.n32 VDDA.t57 39.4005
R363 VDDA.n32 VDDA.t145 39.4005
R364 VDDA.n30 VDDA.t115 39.4005
R365 VDDA.n30 VDDA.t113 39.4005
R366 VDDA.n28 VDDA.t5 39.4005
R367 VDDA.n28 VDDA.t89 39.4005
R368 VDDA.n27 VDDA.t134 39.4005
R369 VDDA.n27 VDDA.t84 39.4005
R370 VDDA VDDA.n3 32.4135
R371 VDDA.n130 VDDA.n129 21.3338
R372 VDDA.n140 VDDA.n132 21.3338
R373 VDDA.n102 VDDA.n101 21.3338
R374 VDDA.n112 VDDA.n104 21.3338
R375 VDDA.n16 VDDA.n15 21.3338
R376 VDDA.n62 VDDA.n17 21.3338
R377 VDDA.n39 VDDA.n38 21.3338
R378 VDDA.n37 VDDA.n36 21.3338
R379 VDDA.n205 VDDA.n204 19.2005
R380 VDDA.n195 VDDA.n194 19.2005
R381 VDDA.n191 VDDA.n190 19.2005
R382 VDDA.n181 VDDA.n180 19.2005
R383 VDDA.n177 VDDA.n176 19.2005
R384 VDDA.n167 VDDA.n166 19.2005
R385 VDDA.n126 VDDA.n125 19.2005
R386 VDDA.n116 VDDA.n115 19.2005
R387 VDDA.n114 VDDA.n113 16.363
R388 VDDA.n212 VDDA.t40 15.0181
R389 VDDA.n166 VDDA.n165 14.8005
R390 VDDA.n194 VDDA.n193 13.8005
R391 VDDA.n180 VDDA.n179 13.8005
R392 VDDA.n178 VDDA.n177 13.8005
R393 VDDA.n192 VDDA.n191 13.8005
R394 VDDA.n206 VDDA.n205 13.8005
R395 VDDA.n115 VDDA.n114 13.8005
R396 VDDA.n127 VDDA.n126 13.8005
R397 VDDA.n84 VDDA.t152 13.1338
R398 VDDA.n84 VDDA.t32 13.1338
R399 VDDA.n87 VDDA.t69 13.1338
R400 VDDA.n87 VDDA.t136 13.1338
R401 VDDA.n89 VDDA.t25 13.1338
R402 VDDA.n89 VDDA.t117 13.1338
R403 VDDA.n91 VDDA.t120 13.1338
R404 VDDA.n91 VDDA.t86 13.1338
R405 VDDA.n93 VDDA.t45 13.1338
R406 VDDA.n93 VDDA.t42 13.1338
R407 VDDA.n95 VDDA.t55 13.1338
R408 VDDA.n95 VDDA.t82 13.1338
R409 VDDA.n97 VDDA.t53 13.1338
R410 VDDA.n97 VDDA.t15 13.1338
R411 VDDA.n99 VDDA.t39 13.1338
R412 VDDA.n99 VDDA.t74 13.1338
R413 VDDA.n142 VDDA.n141 9.3005
R414 VDDA.n81 VDDA.n80 9.3005
R415 VDDA.n79 VDDA.n78 9.3005
R416 VDDA.n76 VDDA.n75 9.3005
R417 VDDA.n71 VDDA.n7 9.3005
R418 VDDA.n68 VDDA.n67 9.3005
R419 VDDA.n12 VDDA.n11 9.3005
R420 VDDA.n22 VDDA.n21 9.3005
R421 VDDA.n25 VDDA.n18 9.3005
R422 VDDA.n60 VDDA.n59 9.3005
R423 VDDA.n48 VDDA.n46 9.3005
R424 VDDA.n3 VDDA.n2 8.03219
R425 VDDA.n83 VDDA.n82 6.098
R426 VDDA.n144 VDDA.n143 5.69621
R427 VDDA.n207 VDDA.n206 5.1605
R428 VDDA.n143 VDDA.n142 4.50831
R429 VDDA.n49 VDDA.n48 4.5005
R430 VDDA.n59 VDDA.n58 4.5005
R431 VDDA.n26 VDDA.n25 4.5005
R432 VDDA.n23 VDDA.n22 4.5005
R433 VDDA.n11 VDDA.n8 4.5005
R434 VDDA.n69 VDDA.n68 4.5005
R435 VDDA.n72 VDDA.n71 4.5005
R436 VDDA.n75 VDDA.n73 4.5005
R437 VDDA.n78 VDDA.n4 4.5005
R438 VDDA.n82 VDDA.n81 4.5005
R439 VDDA.n1 VDDA.n0 4.12334
R440 VDDA.n58 VDDA.n57 3.3755
R441 VDDA.n2 VDDA.n1 2.93377
R442 VDDA.n143 VDDA.n127 2.91121
R443 VDDA.n179 VDDA.n178 1.813
R444 VDDA.n193 VDDA.n192 1.813
R445 VDDA VDDA.n212 1.0815
R446 VDDA.n165 VDDA.n162 1.0005
R447 VDDA.n178 VDDA.n162 1.0005
R448 VDDA.n179 VDDA.n160 1.0005
R449 VDDA.n160 VDDA.n158 1.0005
R450 VDDA.n158 VDDA.n156 1.0005
R451 VDDA.n156 VDDA.n154 1.0005
R452 VDDA.n154 VDDA.n151 1.0005
R453 VDDA.n192 VDDA.n151 1.0005
R454 VDDA.n193 VDDA.n149 1.0005
R455 VDDA.n149 VDDA.n146 1.0005
R456 VDDA.n206 VDDA.n146 1.0005
R457 VDDA.n114 VDDA.n100 1.0005
R458 VDDA.n100 VDDA.n98 1.0005
R459 VDDA.n98 VDDA.n96 1.0005
R460 VDDA.n96 VDDA.n94 1.0005
R461 VDDA.n94 VDDA.n92 1.0005
R462 VDDA.n92 VDDA.n90 1.0005
R463 VDDA.n90 VDDA.n88 1.0005
R464 VDDA.n88 VDDA.n85 1.0005
R465 VDDA.n127 VDDA.n85 1.0005
R466 VDDA.n83 VDDA.n3 0.840625
R467 VDDA.n144 VDDA.n83 0.74075
R468 VDDA.n31 VDDA.n29 0.6255
R469 VDDA.n33 VDDA.n31 0.6255
R470 VDDA.n49 VDDA.n33 0.6255
R471 VDDA.n51 VDDA.n49 0.6255
R472 VDDA.n53 VDDA.n51 0.6255
R473 VDDA.n55 VDDA.n53 0.6255
R474 VDDA.n57 VDDA.n55 0.6255
R475 VDDA.n58 VDDA.n26 0.6255
R476 VDDA.n26 VDDA.n23 0.6255
R477 VDDA.n23 VDDA.n8 0.6255
R478 VDDA.n69 VDDA.n8 0.6255
R479 VDDA.n72 VDDA.n69 0.6255
R480 VDDA.n73 VDDA.n72 0.6255
R481 VDDA.n73 VDDA.n4 0.6255
R482 VDDA.n82 VDDA.n4 0.6255
R483 VDDA.n207 VDDA.n144 0.546875
R484 VDDA.n212 VDDA.n207 0.370625
R485 VDDA.t132 VDDA.t37 0.1603
R486 VDDA.t72 VDDA.t87 0.1603
R487 VDDA.t47 VDDA.t26 0.1603
R488 VDDA.t118 VDDA.t98 0.1603
R489 VDDA.t158 VDDA.t99 0.1603
R490 VDDA.t137 VDDA.t80 0.1603
R491 VDDA.t46 VDDA.t153 0.1603
R492 VDDA.t159 VDDA.t79 0.1603
R493 VDDA.n209 VDDA.t146 0.159278
R494 VDDA.n210 VDDA.t97 0.159278
R495 VDDA.n211 VDDA.t131 0.159278
R496 VDDA.n211 VDDA.t132 0.1368
R497 VDDA.n211 VDDA.t72 0.1368
R498 VDDA.n210 VDDA.t47 0.1368
R499 VDDA.n210 VDDA.t118 0.1368
R500 VDDA.n209 VDDA.t158 0.1368
R501 VDDA.n209 VDDA.t137 0.1368
R502 VDDA.n208 VDDA.t46 0.1368
R503 VDDA.n208 VDDA.t159 0.1368
R504 VDDA.t146 VDDA.n208 0.00152174
R505 VDDA.t97 VDDA.n209 0.00152174
R506 VDDA.t131 VDDA.n210 0.00152174
R507 VDDA.t40 VDDA.n211 0.00152174
R508 V_CMFB_S1.n2 V_CMFB_S1.n0 340.272
R509 V_CMFB_S1.n2 V_CMFB_S1.n1 339.272
R510 V_CMFB_S1.n4 V_CMFB_S1.n3 287.264
R511 V_CMFB_S1 V_CMFB_S1.n4 70.9787
R512 V_CMFB_S1.n4 V_CMFB_S1.n2 53.01
R513 V_CMFB_S1.n3 V_CMFB_S1.t5 39.4005
R514 V_CMFB_S1.n3 V_CMFB_S1.t2 39.4005
R515 V_CMFB_S1.n1 V_CMFB_S1.t3 39.4005
R516 V_CMFB_S1.n1 V_CMFB_S1.t1 39.4005
R517 V_CMFB_S1.n0 V_CMFB_S1.t0 39.4005
R518 V_CMFB_S1.n0 V_CMFB_S1.t4 39.4005
R519 V_TOP.n0 V_TOP.t37 369.534
R520 V_TOP.n10 V_TOP.n8 339.959
R521 V_TOP.n7 V_TOP.n6 339.272
R522 V_TOP.n15 V_TOP.n14 339.272
R523 V_TOP.n17 V_TOP.n16 339.272
R524 V_TOP.n10 V_TOP.n9 339.272
R525 V_TOP.n12 V_TOP.n11 334.772
R526 V_TOP.n1 V_TOP.n0 224.934
R527 V_TOP.n2 V_TOP.n1 224.934
R528 V_TOP.n3 V_TOP.n2 224.934
R529 V_TOP.n4 V_TOP.n3 224.934
R530 V_TOP.n5 V_TOP.n4 224.934
R531 V_TOP.n27 V_TOP.n26 224.934
R532 V_TOP.n26 V_TOP.n25 224.934
R533 V_TOP.n25 V_TOP.n24 224.934
R534 V_TOP.n24 V_TOP.n23 224.934
R535 V_TOP.n23 V_TOP.n22 224.934
R536 V_TOP.n22 V_TOP.n21 224.934
R537 V_TOP.n21 V_TOP.n20 224.934
R538 V_TOP V_TOP.t17 214.222
R539 V_TOP V_TOP.n40 203.69
R540 V_TOP.n7 V_TOP.t6 176.114
R541 V_TOP.n19 V_TOP.n18 163.175
R542 V_TOP.n0 V_TOP.t40 144.601
R543 V_TOP.n1 V_TOP.t23 144.601
R544 V_TOP.n2 V_TOP.t26 144.601
R545 V_TOP.n3 V_TOP.t38 144.601
R546 V_TOP.n4 V_TOP.t41 144.601
R547 V_TOP.n5 V_TOP.t48 144.601
R548 V_TOP.n27 V_TOP.t15 144.601
R549 V_TOP.n26 V_TOP.t36 144.601
R550 V_TOP.n25 V_TOP.t21 144.601
R551 V_TOP.n24 V_TOP.t16 144.601
R552 V_TOP.n23 V_TOP.t14 144.601
R553 V_TOP.n22 V_TOP.t43 144.601
R554 V_TOP.n21 V_TOP.t31 144.601
R555 V_TOP.n20 V_TOP.t27 144.601
R556 V_TOP.n18 V_TOP.t9 95.447
R557 V_TOP.n19 V_TOP.n5 69.6227
R558 V_TOP V_TOP.n27 69.6227
R559 V_TOP.n20 V_TOP.n19 69.6227
R560 V_TOP.n6 V_TOP.t2 39.4005
R561 V_TOP.n6 V_TOP.t11 39.4005
R562 V_TOP.n11 V_TOP.t7 39.4005
R563 V_TOP.n11 V_TOP.t5 39.4005
R564 V_TOP.n9 V_TOP.t10 39.4005
R565 V_TOP.n9 V_TOP.t1 39.4005
R566 V_TOP.n8 V_TOP.t3 39.4005
R567 V_TOP.n8 V_TOP.t12 39.4005
R568 V_TOP.n14 V_TOP.t8 39.4005
R569 V_TOP.n14 V_TOP.t4 39.4005
R570 V_TOP.n16 V_TOP.t13 39.4005
R571 V_TOP.n16 V_TOP.t0 39.4005
R572 V_TOP.n12 V_TOP.n10 8.313
R573 V_TOP.n18 V_TOP.n17 5.188
R574 V_TOP.n28 V_TOP.t49 4.8295
R575 V_TOP.n29 V_TOP.t35 4.8295
R576 V_TOP.n31 V_TOP.t20 4.8295
R577 V_TOP.n32 V_TOP.t44 4.8295
R578 V_TOP.n34 V_TOP.t46 4.8295
R579 V_TOP.n35 V_TOP.t33 4.8295
R580 V_TOP.n37 V_TOP.t25 4.8295
R581 V_TOP.n28 V_TOP.t30 4.5005
R582 V_TOP.n30 V_TOP.t24 4.5005
R583 V_TOP.n29 V_TOP.t45 4.5005
R584 V_TOP.n31 V_TOP.t39 4.5005
R585 V_TOP.n33 V_TOP.t29 4.5005
R586 V_TOP.n32 V_TOP.t18 4.5005
R587 V_TOP.n34 V_TOP.t28 4.5005
R588 V_TOP.n36 V_TOP.t22 4.5005
R589 V_TOP.n35 V_TOP.t42 4.5005
R590 V_TOP.n40 V_TOP.t34 4.5005
R591 V_TOP.n39 V_TOP.t19 4.5005
R592 V_TOP.n38 V_TOP.t47 4.5005
R593 V_TOP.n37 V_TOP.t32 4.5005
R594 V_TOP.n13 V_TOP.n12 4.5005
R595 V_TOP.n17 V_TOP.n15 2.1255
R596 V_TOP.n15 V_TOP.n13 2.1255
R597 V_TOP.n13 V_TOP.n7 2.1255
R598 V_TOP.n30 V_TOP.n28 0.3295
R599 V_TOP.n30 V_TOP.n29 0.3295
R600 V_TOP.n33 V_TOP.n31 0.3295
R601 V_TOP.n33 V_TOP.n32 0.3295
R602 V_TOP.n36 V_TOP.n34 0.3295
R603 V_TOP.n36 V_TOP.n35 0.3295
R604 V_TOP.n40 V_TOP.n39 0.3295
R605 V_TOP.n39 V_TOP.n38 0.3295
R606 V_TOP.n38 V_TOP.n37 0.3295
R607 V_TOP.n33 V_TOP.n30 0.2825
R608 V_TOP.n36 V_TOP.n33 0.2825
R609 V_TOP.n38 V_TOP.n36 0.2825
R610 Vin+.n3 Vin+.n2 526.183
R611 Vin+.n1 Vin+.n0 514.134
R612 Vin+.n0 Vin+.t7 303.259
R613 Vin+.n7 Vin+.n3 215.732
R614 Vin+.n0 Vin+.t8 174.726
R615 Vin+.n1 Vin+.t10 174.726
R616 Vin+.n2 Vin+.t9 174.726
R617 Vin+.n6 Vin+.n4 170.56
R618 Vin+.n6 Vin+.n5 168.435
R619 Vin+.t0 Vin+.n8 158.796
R620 Vin+.n8 Vin+.t1 147.981
R621 Vin+.n2 Vin+.n1 128.534
R622 Vin+.n3 Vin+.t6 96.4005
R623 Vin+.n7 Vin+.n6 13.5005
R624 Vin+.n5 Vin+.t2 13.1338
R625 Vin+.n5 Vin+.t4 13.1338
R626 Vin+.n4 Vin+.t5 13.1338
R627 Vin+.n4 Vin+.t3 13.1338
R628 Vin+.n8 Vin+.n7 1.438
R629 V_p_1.n0 V_p_1.n1 229.562
R630 V_p_1.n0 V_p_1.n4 228.939
R631 V_p_1.n0 V_p_1.n3 228.939
R632 V_p_1.n0 V_p_1.n2 228.939
R633 V_p_1.n5 V_p_1.n0 228.938
R634 V_p_1.n0 V_p_1.t10 100.103
R635 V_p_1.n4 V_p_1.t4 48.0005
R636 V_p_1.n4 V_p_1.t8 48.0005
R637 V_p_1.n3 V_p_1.t1 48.0005
R638 V_p_1.n3 V_p_1.t7 48.0005
R639 V_p_1.n2 V_p_1.t5 48.0005
R640 V_p_1.n2 V_p_1.t2 48.0005
R641 V_p_1.n1 V_p_1.t3 48.0005
R642 V_p_1.n1 V_p_1.t6 48.0005
R643 V_p_1.n5 V_p_1.t9 48.0005
R644 V_p_1.t0 V_p_1.n5 48.0005
R645 GNDA.n1974 GNDA.n1973 46964.7
R646 GNDA.n1976 GNDA.n1975 29808.3
R647 GNDA.n1976 GNDA.n88 26648.4
R648 GNDA.n2000 GNDA.n82 12361.8
R649 GNDA.n1996 GNDA.n82 12312.5
R650 GNDA.n2000 GNDA.n83 11918.5
R651 GNDA.n1996 GNDA.n83 11869.2
R652 GNDA.n1975 GNDA.n1974 11754
R653 GNDA.n1974 GNDA.n90 11338.5
R654 GNDA.n1973 GNDA.n1972 11169.2
R655 GNDA.n91 GNDA.n88 11169.2
R656 GNDA.n1980 GNDA.n1976 10371.4
R657 GNDA.n1971 GNDA.n91 9642.55
R658 GNDA.n1970 GNDA.n88 8207.69
R659 GNDA.n1484 GNDA.n1474 8175.5
R660 GNDA.n1506 GNDA.n1474 8126.25
R661 GNDA.n1973 GNDA.n91 7898.5
R662 GNDA.n1978 GNDA.n70 7880
R663 GNDA.n2003 GNDA.n70 7880
R664 GNDA.n1989 GNDA.n87 7880
R665 GNDA.n1989 GNDA.n1982 7880
R666 GNDA.n1978 GNDA.n71 7830.75
R667 GNDA.n2003 GNDA.n71 7830.75
R668 GNDA.n87 GNDA.n86 7830.75
R669 GNDA.n1982 GNDA.n86 7830.75
R670 GNDA.n1484 GNDA.n1475 7732.25
R671 GNDA.n1506 GNDA.n1475 7683
R672 GNDA.n1488 GNDA.n1480 6845.75
R673 GNDA.n1488 GNDA.n1481 6845.75
R674 GNDA.n1493 GNDA.n1480 6796.5
R675 GNDA.n1493 GNDA.n1481 6796.5
R676 GNDA.n1502 GNDA.n1497 6698
R677 GNDA.n1500 GNDA.n1497 6698
R678 GNDA.n1502 GNDA.n1501 6648.75
R679 GNDA.n1501 GNDA.n1500 6648.75
R680 GNDA.n1972 GNDA.n1971 6291.31
R681 GNDA.n1959 GNDA.n67 6254.75
R682 GNDA.n2018 GNDA.n67 6254.75
R683 GNDA.n1959 GNDA.n68 6254.75
R684 GNDA.n2018 GNDA.n68 6254.75
R685 GNDA.n63 GNDA.n58 5368.25
R686 GNDA.n2025 GNDA.n58 5368.25
R687 GNDA.n63 GNDA.n59 5368.25
R688 GNDA.n2025 GNDA.n59 5368.25
R689 GNDA.n1968 GNDA.n93 5368.25
R690 GNDA.n1962 GNDA.n93 5368.25
R691 GNDA.n1968 GNDA.n94 5368.25
R692 GNDA.n1962 GNDA.n94 5368.25
R693 GNDA.n1971 GNDA.n1970 5223.84
R694 GNDA.n2014 GNDA.n72 4974.25
R695 GNDA.n2014 GNDA.n73 4974.25
R696 GNDA.n1738 GNDA.n242 4678.75
R697 GNDA.n1734 GNDA.n242 4629.5
R698 GNDA.n1738 GNDA.n243 4629.5
R699 GNDA.n1563 GNDA.n1307 4580.25
R700 GNDA.n1563 GNDA.n1308 4580.25
R701 GNDA.n1734 GNDA.n243 4580.25
R702 GNDA.n1566 GNDA.n1565 4580.25
R703 GNDA.n1565 GNDA.n1314 4580.25
R704 GNDA.n72 GNDA.n69 4531
R705 GNDA.n73 GNDA.n69 4531
R706 GNDA.n1570 GNDA.n1307 4481.75
R707 GNDA.n1570 GNDA.n1308 4481.75
R708 GNDA.n1566 GNDA.n1203 4481.75
R709 GNDA.n1314 GNDA.n1203 4481.75
R710 GNDA.n1970 GNDA.n1969 4375.88
R711 GNDA.n1972 GNDA.n90 3484.9
R712 GNDA.n1487 GNDA.n90 3260.59
R713 GNDA.n1975 GNDA.n89 2543.73
R714 GNDA.n1033 GNDA.n876 2429.06
R715 GNDA.n1993 GNDA.n85 2371.15
R716 GNDA.n1957 GNDA.n85 2371.15
R717 GNDA.n1740 GNDA.n89 2026.18
R718 GNDA.n2078 GNDA.n2077 1748.05
R719 GNDA.n1305 GNDA.n1204 1323.19
R720 GNDA.n1991 GNDA.n85 1301.55
R721 GNDA.n1739 GNDA.n241 1285.24
R722 GNDA.n589 GNDA.t70 1012.05
R723 GNDA.n886 GNDA.t70 1012.05
R724 GNDA.n2166 GNDA.t70 990.407
R725 GNDA.n607 GNDA.t70 990.407
R726 GNDA.n1835 GNDA.n199 949.682
R727 GNDA.n1931 GNDA.n1930 949.682
R728 GNDA.n1999 GNDA.n75 803.201
R729 GNDA.n1997 GNDA.n75 800
R730 GNDA.n1999 GNDA.n1998 774.4
R731 GNDA.n1998 GNDA.n1997 771.201
R732 GNDA.n1948 GNDA.n1947 669.307
R733 GNDA.n1835 GNDA.n1834 662.155
R734 GNDA.n1930 GNDA.n1929 662.155
R735 GNDA.n1835 GNDA.n200 623.755
R736 GNDA.n1930 GNDA.n134 623.755
R737 GNDA.n1836 GNDA.n197 588.271
R738 GNDA.n56 GNDA.n54 588.271
R739 GNDA.n2169 GNDA.n2168 585
R740 GNDA.n2170 GNDA.n29 585
R741 GNDA.n2172 GNDA.n2171 585
R742 GNDA.n2174 GNDA.n27 585
R743 GNDA.n2176 GNDA.n2175 585
R744 GNDA.n2177 GNDA.n26 585
R745 GNDA.n2179 GNDA.n2178 585
R746 GNDA.n2181 GNDA.n24 585
R747 GNDA.n2183 GNDA.n2182 585
R748 GNDA.n2184 GNDA.n23 585
R749 GNDA.n2186 GNDA.n2185 585
R750 GNDA.n2188 GNDA.n13 585
R751 GNDA.n1063 GNDA.n860 585
R752 GNDA.n1064 GNDA.n858 585
R753 GNDA.n1065 GNDA.n857 585
R754 GNDA.n855 GNDA.n852 585
R755 GNDA.n1070 GNDA.n851 585
R756 GNDA.n1071 GNDA.n849 585
R757 GNDA.n1072 GNDA.n848 585
R758 GNDA.n846 GNDA.n843 585
R759 GNDA.n1077 GNDA.n842 585
R760 GNDA.n1078 GNDA.n840 585
R761 GNDA.n1079 GNDA.n839 585
R762 GNDA.n920 GNDA.n837 585
R763 GNDA.n835 GNDA.n21 585
R764 GNDA.n2190 GNDA.n21 585
R765 GNDA.n1063 GNDA.n1062 585
R766 GNDA.n1064 GNDA.n854 585
R767 GNDA.n1066 GNDA.n1065 585
R768 GNDA.n1068 GNDA.n852 585
R769 GNDA.n1070 GNDA.n1069 585
R770 GNDA.n1071 GNDA.n845 585
R771 GNDA.n1073 GNDA.n1072 585
R772 GNDA.n1075 GNDA.n843 585
R773 GNDA.n1077 GNDA.n1076 585
R774 GNDA.n1078 GNDA.n838 585
R775 GNDA.n1080 GNDA.n1079 585
R776 GNDA.n1082 GNDA.n837 585
R777 GNDA.n830 GNDA.n829 585
R778 GNDA.n827 GNDA.n663 585
R779 GNDA.n826 GNDA.n664 585
R780 GNDA.n824 GNDA.n823 585
R781 GNDA.n666 GNDA.n665 585
R782 GNDA.n815 GNDA.n814 585
R783 GNDA.n812 GNDA.n668 585
R784 GNDA.n810 GNDA.n809 585
R785 GNDA.n670 GNDA.n669 585
R786 GNDA.n803 GNDA.n802 585
R787 GNDA.n800 GNDA.n672 585
R788 GNDA.n798 GNDA.n797 585
R789 GNDA.n2192 GNDA.n2191 585
R790 GNDA.n2191 GNDA.n2190 585
R791 GNDA.n444 GNDA.n20 585
R792 GNDA.n2190 GNDA.n20 585
R793 GNDA.n831 GNDA.n830 585
R794 GNDA.n819 GNDA.n663 585
R795 GNDA.n820 GNDA.n664 585
R796 GNDA.n823 GNDA.n822 585
R797 GNDA.n818 GNDA.n666 585
R798 GNDA.n816 GNDA.n815 585
R799 GNDA.n668 GNDA.n667 585
R800 GNDA.n809 GNDA.n808 585
R801 GNDA.n806 GNDA.n670 585
R802 GNDA.n804 GNDA.n803 585
R803 GNDA.n672 GNDA.n671 585
R804 GNDA.n797 GNDA.n796 585
R805 GNDA.n484 GNDA.n483 585
R806 GNDA.n480 GNDA.n479 585
R807 GNDA.n556 GNDA.n555 585
R808 GNDA.n558 GNDA.n478 585
R809 GNDA.n561 GNDA.n560 585
R810 GNDA.n475 GNDA.n474 585
R811 GNDA.n570 GNDA.n569 585
R812 GNDA.n574 GNDA.n573 585
R813 GNDA.n572 GNDA.n470 585
R814 GNDA.n581 GNDA.n580 585
R815 GNDA.n583 GNDA.n582 585
R816 GNDA.n586 GNDA.n585 585
R817 GNDA.n613 GNDA.n612 585
R818 GNDA.n615 GNDA.n452 585
R819 GNDA.n617 GNDA.n616 585
R820 GNDA.n618 GNDA.n451 585
R821 GNDA.n620 GNDA.n619 585
R822 GNDA.n622 GNDA.n449 585
R823 GNDA.n624 GNDA.n623 585
R824 GNDA.n625 GNDA.n448 585
R825 GNDA.n627 GNDA.n626 585
R826 GNDA.n629 GNDA.n447 585
R827 GNDA.n630 GNDA.n445 585
R828 GNDA.n633 GNDA.n632 585
R829 GNDA.n924 GNDA.n923 585
R830 GNDA.n918 GNDA.n917 585
R831 GNDA.n983 GNDA.n982 585
R832 GNDA.n985 GNDA.n916 585
R833 GNDA.n988 GNDA.n987 585
R834 GNDA.n914 GNDA.n913 585
R835 GNDA.n995 GNDA.n994 585
R836 GNDA.n997 GNDA.n911 585
R837 GNDA.n1000 GNDA.n999 585
R838 GNDA.n890 GNDA.n889 585
R839 GNDA.n1008 GNDA.n1007 585
R840 GNDA.n1011 GNDA.n1010 585
R841 GNDA.n2167 GNDA.n30 585
R842 GNDA.n2167 GNDA.n2166 585
R843 GNDA.n2161 GNDA.n32 585
R844 GNDA.n2165 GNDA.n32 585
R845 GNDA.n2163 GNDA.n2162 585
R846 GNDA.n2164 GNDA.n2163 585
R847 GNDA.n2160 GNDA.n34 585
R848 GNDA.n34 GNDA.n33 585
R849 GNDA.n2159 GNDA.n2158 585
R850 GNDA.n2158 GNDA.n2157 585
R851 GNDA.n36 GNDA.n35 585
R852 GNDA.n2156 GNDA.n36 585
R853 GNDA.n2067 GNDA.n2065 585
R854 GNDA.n2065 GNDA.n37 585
R855 GNDA.n2069 GNDA.n2068 585
R856 GNDA.n2070 GNDA.n2069 585
R857 GNDA.n2066 GNDA.n2063 585
R858 GNDA.n2071 GNDA.n2063 585
R859 GNDA.n2073 GNDA.n2064 585
R860 GNDA.n2073 GNDA.n2072 585
R861 GNDA.n611 GNDA.n454 585
R862 GNDA.n607 GNDA.n454 585
R863 GNDA.n610 GNDA.n609 585
R864 GNDA.n609 GNDA.n608 585
R865 GNDA.n456 GNDA.n455 585
R866 GNDA.n606 GNDA.n456 585
R867 GNDA.n604 GNDA.n603 585
R868 GNDA.n605 GNDA.n604 585
R869 GNDA.n602 GNDA.n458 585
R870 GNDA.n458 GNDA.n457 585
R871 GNDA.n601 GNDA.n600 585
R872 GNDA.n600 GNDA.n599 585
R873 GNDA.n460 GNDA.n459 585
R874 GNDA.n598 GNDA.n460 585
R875 GNDA.n596 GNDA.n595 585
R876 GNDA.n597 GNDA.n596 585
R877 GNDA.n594 GNDA.n463 585
R878 GNDA.n463 GNDA.n462 585
R879 GNDA.n593 GNDA.n592 585
R880 GNDA.n592 GNDA.n591 585
R881 GNDA.n590 GNDA.n465 585
R882 GNDA.n589 GNDA.n588 585
R883 GNDA.n1035 GNDA.n1034 585
R884 GNDA.n1034 GNDA.n1033 585
R885 GNDA.n879 GNDA.n878 585
R886 GNDA.n1032 GNDA.n879 585
R887 GNDA.n1030 GNDA.n1029 585
R888 GNDA.n1031 GNDA.n1030 585
R889 GNDA.n1028 GNDA.n881 585
R890 GNDA.n881 GNDA.n880 585
R891 GNDA.n1027 GNDA.n1026 585
R892 GNDA.n1026 GNDA.n1025 585
R893 GNDA.n1024 GNDA.n882 585
R894 GNDA.n1024 GNDA.n871 585
R895 GNDA.n1023 GNDA.n1022 585
R896 GNDA.n1023 GNDA.n870 585
R897 GNDA.n1021 GNDA.n883 585
R898 GNDA.n1017 GNDA.n883 585
R899 GNDA.n1020 GNDA.n1019 585
R900 GNDA.n1019 GNDA.n1018 585
R901 GNDA.n885 GNDA.n884 585
R902 GNDA.n1016 GNDA.n885 585
R903 GNDA.n1015 GNDA.n1014 585
R904 GNDA.n887 GNDA.n886 585
R905 GNDA.n1060 GNDA.n1059 585
R906 GNDA.n1059 GNDA.n134 585
R907 GNDA.n1036 GNDA.n877 585
R908 GNDA.n877 GNDA.n876 585
R909 GNDA.n1038 GNDA.n1037 585
R910 GNDA.n1039 GNDA.n1038 585
R911 GNDA.n875 GNDA.n874 585
R912 GNDA.n1040 GNDA.n875 585
R913 GNDA.n1043 GNDA.n1042 585
R914 GNDA.n1042 GNDA.n1041 585
R915 GNDA.n1044 GNDA.n873 585
R916 GNDA.n873 GNDA.n872 585
R917 GNDA.n1046 GNDA.n1045 585
R918 GNDA.n1047 GNDA.n1046 585
R919 GNDA.n868 GNDA.n867 585
R920 GNDA.n1048 GNDA.n868 585
R921 GNDA.n1051 GNDA.n1050 585
R922 GNDA.n1050 GNDA.n1049 585
R923 GNDA.n1052 GNDA.n865 585
R924 GNDA.n865 GNDA.n864 585
R925 GNDA.n1054 GNDA.n1053 585
R926 GNDA.n1055 GNDA.n1054 585
R927 GNDA.n866 GNDA.n862 585
R928 GNDA.n1056 GNDA.n862 585
R929 GNDA.n1058 GNDA.n863 585
R930 GNDA.n1058 GNDA.n1057 585
R931 GNDA.n124 GNDA.n123 585
R932 GNDA.n1945 GNDA.n1944 585
R933 GNDA.n1946 GNDA.n1945 585
R934 GNDA.n1280 GNDA.n1215 585
R935 GNDA.n1280 GNDA.n199 585
R936 GNDA.n1283 GNDA.n1282 585
R937 GNDA.n1282 GNDA.n1281 585
R938 GNDA.n1284 GNDA.n1213 585
R939 GNDA.n1213 GNDA.n1212 585
R940 GNDA.n1286 GNDA.n1285 585
R941 GNDA.n1287 GNDA.n1286 585
R942 GNDA.n1214 GNDA.n1211 585
R943 GNDA.n1288 GNDA.n1211 585
R944 GNDA.n1290 GNDA.n1210 585
R945 GNDA.n1290 GNDA.n1289 585
R946 GNDA.n1293 GNDA.n1292 585
R947 GNDA.n1292 GNDA.n1291 585
R948 GNDA.n1294 GNDA.n1209 585
R949 GNDA.n1209 GNDA.n1208 585
R950 GNDA.n1296 GNDA.n1295 585
R951 GNDA.n1297 GNDA.n1296 585
R952 GNDA.n1207 GNDA.n1206 585
R953 GNDA.n1298 GNDA.n1207 585
R954 GNDA.n1301 GNDA.n1300 585
R955 GNDA.n1300 GNDA.n1299 585
R956 GNDA.n1302 GNDA.n1205 585
R957 GNDA.n1205 GNDA.n1204 585
R958 GNDA.n133 GNDA.n132 585
R959 GNDA.n1931 GNDA.n133 585
R960 GNDA.n1934 GNDA.n1933 585
R961 GNDA.n1933 GNDA.n1932 585
R962 GNDA.n1935 GNDA.n131 585
R963 GNDA.n131 GNDA.n130 585
R964 GNDA.n1937 GNDA.n1936 585
R965 GNDA.n1938 GNDA.n1937 585
R966 GNDA.n129 GNDA.n127 585
R967 GNDA.n1939 GNDA.n129 585
R968 GNDA.n1942 GNDA.n1941 585
R969 GNDA.n1941 GNDA.n1940 585
R970 GNDA.n128 GNDA.n126 585
R971 GNDA.n128 GNDA.n125 585
R972 GNDA.n1268 GNDA.n1267 585
R973 GNDA.n1267 GNDA.n1266 585
R974 GNDA.n1269 GNDA.n1264 585
R975 GNDA.n1264 GNDA.n1263 585
R976 GNDA.n1271 GNDA.n1270 585
R977 GNDA.n1272 GNDA.n1271 585
R978 GNDA.n1265 GNDA.n1261 585
R979 GNDA.n1273 GNDA.n1261 585
R980 GNDA.n1275 GNDA.n1262 585
R981 GNDA.n1275 GNDA.n1274 585
R982 GNDA.n1277 GNDA.n1276 585
R983 GNDA.n1276 GNDA.n200 585
R984 GNDA.n1597 GNDA.n1596 585
R985 GNDA.n1185 GNDA.n1184 585
R986 GNDA.n1656 GNDA.n1655 585
R987 GNDA.n1658 GNDA.n1183 585
R988 GNDA.n1661 GNDA.n1660 585
R989 GNDA.n1181 GNDA.n1180 585
R990 GNDA.n1668 GNDA.n1667 585
R991 GNDA.n1670 GNDA.n1178 585
R992 GNDA.n1673 GNDA.n1672 585
R993 GNDA.n1157 GNDA.n1156 585
R994 GNDA.n1681 GNDA.n1680 585
R995 GNDA.n1684 GNDA.n1683 585
R996 GNDA.n1435 GNDA.n1434 585
R997 GNDA.n1437 GNDA.n1356 585
R998 GNDA.n1439 GNDA.n1438 585
R999 GNDA.n1440 GNDA.n1355 585
R1000 GNDA.n1442 GNDA.n1441 585
R1001 GNDA.n1444 GNDA.n1353 585
R1002 GNDA.n1446 GNDA.n1445 585
R1003 GNDA.n1447 GNDA.n1352 585
R1004 GNDA.n1449 GNDA.n1448 585
R1005 GNDA.n1451 GNDA.n1350 585
R1006 GNDA.n1453 GNDA.n1452 585
R1007 GNDA.n1454 GNDA.n1349 585
R1008 GNDA.n1728 GNDA.n1727 585
R1009 GNDA.n1725 GNDA.n1724 585
R1010 GNDA.n253 GNDA.n252 585
R1011 GNDA.n336 GNDA.n335 585
R1012 GNDA.n338 GNDA.n337 585
R1013 GNDA.n343 GNDA.n342 585
R1014 GNDA.n346 GNDA.n345 585
R1015 GNDA.n328 GNDA.n327 585
R1016 GNDA.n353 GNDA.n352 585
R1017 GNDA.n355 GNDA.n275 585
R1018 GNDA.n1717 GNDA.n1716 585
R1019 GNDA.n1714 GNDA.n1713 585
R1020 GNDA.n1549 GNDA.n382 585
R1021 GNDA.n1551 GNDA.n1550 585
R1022 GNDA.n1548 GNDA.n1529 585
R1023 GNDA.n1547 GNDA.n1546 585
R1024 GNDA.n1545 GNDA.n1544 585
R1025 GNDA.n1543 GNDA.n1542 585
R1026 GNDA.n1541 GNDA.n1540 585
R1027 GNDA.n1539 GNDA.n1538 585
R1028 GNDA.n1537 GNDA.n1536 585
R1029 GNDA.n1535 GNDA.n1534 585
R1030 GNDA.n1533 GNDA.n1532 585
R1031 GNDA.n1531 GNDA.n1530 585
R1032 GNDA.n2074 GNDA.n2060 585
R1033 GNDA.n2077 GNDA.n2076 585
R1034 GNDA.n2197 GNDA.n8 585
R1035 GNDA.n2198 GNDA.n7 585
R1036 GNDA.n2199 GNDA.n6 585
R1037 GNDA.n16 GNDA.n2 585
R1038 GNDA.n2204 GNDA.n1 585
R1039 GNDA.n149 GNDA.n0 585
R1040 GNDA.n153 GNDA.n152 585
R1041 GNDA.n150 GNDA.n145 585
R1042 GNDA.n158 GNDA.n144 585
R1043 GNDA.n159 GNDA.n142 585
R1044 GNDA.n160 GNDA.n141 585
R1045 GNDA.n139 GNDA.n137 585
R1046 GNDA.n2189 GNDA.n9 585
R1047 GNDA.n2190 GNDA.n2189 585
R1048 GNDA.n2197 GNDA.n2196 585
R1049 GNDA.n2198 GNDA.n5 585
R1050 GNDA.n2200 GNDA.n2199 585
R1051 GNDA.n2202 GNDA.n2 585
R1052 GNDA.n2204 GNDA.n2203 585
R1053 GNDA.n147 GNDA.n0 585
R1054 GNDA.n154 GNDA.n153 585
R1055 GNDA.n156 GNDA.n145 585
R1056 GNDA.n158 GNDA.n157 585
R1057 GNDA.n159 GNDA.n138 585
R1058 GNDA.n161 GNDA.n160 585
R1059 GNDA.n163 GNDA.n137 585
R1060 GNDA.n2195 GNDA.n2194 585
R1061 GNDA.n1414 GNDA.n12 585
R1062 GNDA.n1416 GNDA.n1415 585
R1063 GNDA.n1417 GNDA.n1412 585
R1064 GNDA.n1419 GNDA.n1418 585
R1065 GNDA.n1421 GNDA.n1410 585
R1066 GNDA.n1423 GNDA.n1422 585
R1067 GNDA.n1424 GNDA.n1409 585
R1068 GNDA.n1426 GNDA.n1425 585
R1069 GNDA.n1428 GNDA.n1408 585
R1070 GNDA.n1429 GNDA.n1406 585
R1071 GNDA.n1432 GNDA.n1431 585
R1072 GNDA.n689 GNDA.n357 585
R1073 GNDA.n692 GNDA.n691 585
R1074 GNDA.n761 GNDA.n760 585
R1075 GNDA.n763 GNDA.n687 585
R1076 GNDA.n766 GNDA.n765 585
R1077 GNDA.n684 GNDA.n683 585
R1078 GNDA.n776 GNDA.n775 585
R1079 GNDA.n778 GNDA.n682 585
R1080 GNDA.n781 GNDA.n780 585
R1081 GNDA.n679 GNDA.n675 585
R1082 GNDA.n792 GNDA.n791 585
R1083 GNDA.n794 GNDA.n673 585
R1084 GNDA.n833 GNDA.n832 585
R1085 GNDA.n635 GNDA.n634 585
R1086 GNDA.n658 GNDA.n657 585
R1087 GNDA.n656 GNDA.n640 585
R1088 GNDA.n655 GNDA.n654 585
R1089 GNDA.n653 GNDA.n652 585
R1090 GNDA.n651 GNDA.n650 585
R1091 GNDA.n649 GNDA.n648 585
R1092 GNDA.n647 GNDA.n646 585
R1093 GNDA.n645 GNDA.n644 585
R1094 GNDA.n643 GNDA.n642 585
R1095 GNDA.n641 GNDA.n387 585
R1096 GNDA.n1151 GNDA.n1150 585
R1097 GNDA.n398 GNDA.n392 585
R1098 GNDA.n1146 GNDA.n1145 585
R1099 GNDA.n400 GNDA.n397 585
R1100 GNDA.n428 GNDA.n427 585
R1101 GNDA.n432 GNDA.n431 585
R1102 GNDA.n430 GNDA.n421 585
R1103 GNDA.n439 GNDA.n438 585
R1104 GNDA.n441 GNDA.n440 585
R1105 GNDA.n1086 GNDA.n443 585
R1106 GNDA.n1088 GNDA.n1087 585
R1107 GNDA.n1084 GNDA.n1083 585
R1108 GNDA.n1404 GNDA.n1403 585
R1109 GNDA.n1401 GNDA.n1359 585
R1110 GNDA.n1400 GNDA.n1399 585
R1111 GNDA.n1390 GNDA.n1361 585
R1112 GNDA.n1392 GNDA.n1391 585
R1113 GNDA.n1388 GNDA.n1387 585
R1114 GNDA.n1364 GNDA.n1363 585
R1115 GNDA.n1382 GNDA.n1381 585
R1116 GNDA.n1379 GNDA.n1366 585
R1117 GNDA.n1377 GNDA.n1376 585
R1118 GNDA.n1371 GNDA.n1367 585
R1119 GNDA.n1370 GNDA.n1369 585
R1120 GNDA.n1405 GNDA.n388 585
R1121 GNDA.n1688 GNDA.n388 585
R1122 GNDA.n1691 GNDA.n385 585
R1123 GNDA.n383 GNDA.n380 585
R1124 GNDA.n1696 GNDA.n379 585
R1125 GNDA.n1697 GNDA.n377 585
R1126 GNDA.n1698 GNDA.n376 585
R1127 GNDA.n374 GNDA.n371 585
R1128 GNDA.n1703 GNDA.n370 585
R1129 GNDA.n1704 GNDA.n368 585
R1130 GNDA.n1705 GNDA.n367 585
R1131 GNDA.n365 GNDA.n362 585
R1132 GNDA.n1710 GNDA.n361 585
R1133 GNDA.n1711 GNDA.n359 585
R1134 GNDA.n389 GNDA.n358 585
R1135 GNDA.n1688 GNDA.n389 585
R1136 GNDA.n1690 GNDA.n1689 585
R1137 GNDA.n1689 GNDA.n1688 585
R1138 GNDA.n1278 GNDA.n1259 585
R1139 GNDA.n1257 GNDA.n1217 585
R1140 GNDA.n1256 GNDA.n1255 585
R1141 GNDA.n1247 GNDA.n1219 585
R1142 GNDA.n1249 GNDA.n1248 585
R1143 GNDA.n1245 GNDA.n1244 585
R1144 GNDA.n1222 GNDA.n1221 585
R1145 GNDA.n1239 GNDA.n1238 585
R1146 GNDA.n1236 GNDA.n1224 585
R1147 GNDA.n1234 GNDA.n1233 585
R1148 GNDA.n1228 GNDA.n1227 585
R1149 GNDA.n1225 GNDA.n1152 585
R1150 GNDA.n1687 GNDA.n1686 585
R1151 GNDA.n1688 GNDA.n1687 585
R1152 GNDA.n1404 GNDA.n1358 585
R1153 GNDA.n1397 GNDA.n1359 585
R1154 GNDA.n1399 GNDA.n1398 585
R1155 GNDA.n1394 GNDA.n1361 585
R1156 GNDA.n1393 GNDA.n1392 585
R1157 GNDA.n1387 GNDA.n1386 585
R1158 GNDA.n1385 GNDA.n1364 585
R1159 GNDA.n1383 GNDA.n1382 585
R1160 GNDA.n1366 GNDA.n1365 585
R1161 GNDA.n1376 GNDA.n1375 585
R1162 GNDA.n1373 GNDA.n1371 585
R1163 GNDA.n1370 GNDA.n205 585
R1164 GNDA.n1692 GNDA.n1691 585
R1165 GNDA.n1694 GNDA.n380 585
R1166 GNDA.n1696 GNDA.n1695 585
R1167 GNDA.n1697 GNDA.n373 585
R1168 GNDA.n1699 GNDA.n1698 585
R1169 GNDA.n1701 GNDA.n371 585
R1170 GNDA.n1703 GNDA.n1702 585
R1171 GNDA.n1704 GNDA.n364 585
R1172 GNDA.n1706 GNDA.n1705 585
R1173 GNDA.n1708 GNDA.n362 585
R1174 GNDA.n1710 GNDA.n1709 585
R1175 GNDA.n1711 GNDA.n356 585
R1176 GNDA.n1279 GNDA.n1278 585
R1177 GNDA.n1253 GNDA.n1217 585
R1178 GNDA.n1255 GNDA.n1254 585
R1179 GNDA.n1251 GNDA.n1219 585
R1180 GNDA.n1250 GNDA.n1249 585
R1181 GNDA.n1244 GNDA.n1243 585
R1182 GNDA.n1242 GNDA.n1222 585
R1183 GNDA.n1240 GNDA.n1239 585
R1184 GNDA.n1224 GNDA.n1223 585
R1185 GNDA.n1233 GNDA.n1232 585
R1186 GNDA.n1230 GNDA.n1228 585
R1187 GNDA.n1154 GNDA.n1152 585
R1188 GNDA.n57 GNDA.n56 585
R1189 GNDA.n2030 GNDA.n2029 585
R1190 GNDA.n2029 GNDA.n2028 585
R1191 GNDA.n52 GNDA.n51 585
R1192 GNDA.n51 GNDA.n50 585
R1193 GNDA.n2139 GNDA.n2138 585
R1194 GNDA.n2140 GNDA.n2139 585
R1195 GNDA.n49 GNDA.n48 585
R1196 GNDA.n2141 GNDA.n49 585
R1197 GNDA.n2144 GNDA.n2143 585
R1198 GNDA.n2143 GNDA.n2142 585
R1199 GNDA.n45 GNDA.n40 585
R1200 GNDA.n40 GNDA.n38 585
R1201 GNDA.n2154 GNDA.n2153 585
R1202 GNDA.n2155 GNDA.n2154 585
R1203 GNDA.n43 GNDA.n41 585
R1204 GNDA.n41 GNDA.n39 585
R1205 GNDA.n2057 GNDA.n2056 585
R1206 GNDA.n2058 GNDA.n2057 585
R1207 GNDA.n2052 GNDA.n2050 585
R1208 GNDA.n2059 GNDA.n2052 585
R1209 GNDA.n2081 GNDA.n2080 585
R1210 GNDA.n2080 GNDA.n2079 585
R1211 GNDA.n2061 GNDA.n2053 585
R1212 GNDA.n2078 GNDA.n2053 585
R1213 GNDA.n1837 GNDA.n1836 585
R1214 GNDA.n1840 GNDA.n1839 585
R1215 GNDA.n1839 GNDA.n1838 585
R1216 GNDA.n196 GNDA.n195 585
R1217 GNDA.n195 GNDA.n194 585
R1218 GNDA.n1899 GNDA.n1898 585
R1219 GNDA.n1900 GNDA.n1899 585
R1220 GNDA.n1894 GNDA.n193 585
R1221 GNDA.n1901 GNDA.n193 585
R1222 GNDA.n1905 GNDA.n1904 585
R1223 GNDA.n1904 GNDA.n1903 585
R1224 GNDA.n191 GNDA.n190 585
R1225 GNDA.n1902 GNDA.n190 585
R1226 GNDA.n1912 GNDA.n1911 585
R1227 GNDA.n1913 GNDA.n1912 585
R1228 GNDA.n188 GNDA.n186 585
R1229 GNDA.n1914 GNDA.n188 585
R1230 GNDA.n1918 GNDA.n1917 585
R1231 GNDA.n1917 GNDA.n1916 585
R1232 GNDA.n189 GNDA.n165 585
R1233 GNDA.n1915 GNDA.n189 585
R1234 GNDA.n1925 GNDA.n136 585
R1235 GNDA.n136 GNDA.n135 585
R1236 GNDA.n1928 GNDA.n1927 585
R1237 GNDA.n1929 GNDA.n1928 585
R1238 GNDA.n1810 GNDA.n1809 585
R1239 GNDA.n1809 GNDA.n1808 585
R1240 GNDA.n233 GNDA.n232 585
R1241 GNDA.n1807 GNDA.n232 585
R1242 GNDA.n1817 GNDA.n1816 585
R1243 GNDA.n1818 GNDA.n1817 585
R1244 GNDA.n230 GNDA.n228 585
R1245 GNDA.n1819 GNDA.n230 585
R1246 GNDA.n1823 GNDA.n1822 585
R1247 GNDA.n1822 GNDA.n1821 585
R1248 GNDA.n231 GNDA.n207 585
R1249 GNDA.n1820 GNDA.n231 585
R1250 GNDA.n1830 GNDA.n204 585
R1251 GNDA.n204 GNDA.n203 585
R1252 GNDA.n1833 GNDA.n1832 585
R1253 GNDA.n1834 GNDA.n1833 585
R1254 GNDA.n1744 GNDA.n1743 585
R1255 GNDA.n1743 GNDA.n1742 585
R1256 GNDA.n237 GNDA.n236 585
R1257 GNDA.n1741 GNDA.n236 585
R1258 GNDA.n1803 GNDA.n1802 585
R1259 GNDA.n1804 GNDA.n1803 585
R1260 GNDA.n1798 GNDA.n235 585
R1261 GNDA.n1805 GNDA.n235 585
R1262 GNDA.n1457 GNDA.n1348 585
R1263 GNDA.n1458 GNDA.n1457 585
R1264 GNDA.n1461 GNDA.n1460 585
R1265 GNDA.n1460 GNDA.n1459 585
R1266 GNDA.n1462 GNDA.n1346 585
R1267 GNDA.n1346 GNDA.n1345 585
R1268 GNDA.n1464 GNDA.n1463 585
R1269 GNDA.n1465 GNDA.n1464 585
R1270 GNDA.n1347 GNDA.n1344 585
R1271 GNDA.n1466 GNDA.n1344 585
R1272 GNDA.n1469 GNDA.n1468 585
R1273 GNDA.n1468 GNDA.n1467 585
R1274 GNDA.n1470 GNDA.n1333 585
R1275 GNDA.n1333 GNDA.n1331 585
R1276 GNDA.n1472 GNDA.n1471 585
R1277 GNDA.n1473 GNDA.n1472 585
R1278 GNDA.n1343 GNDA.n1332 585
R1279 GNDA.n1332 GNDA.n1330 585
R1280 GNDA.n1342 GNDA.n1341 585
R1281 GNDA.n1341 GNDA.n1340 585
R1282 GNDA.n1339 GNDA.n1335 585
R1283 GNDA.n1338 GNDA.n1337 585
R1284 GNDA.n240 GNDA.n238 585
R1285 GNDA.n241 GNDA.n240 585
R1286 GNDA.n1456 GNDA.n1455 585
R1287 GNDA.n1456 GNDA.n245 585
R1288 GNDA.n1558 GNDA.n1557 585
R1289 GNDA.n1557 GNDA.n1556 585
R1290 GNDA.n1559 GNDA.n1318 585
R1291 GNDA.n1318 GNDA.n1316 585
R1292 GNDA.n1561 GNDA.n1560 585
R1293 GNDA.n1562 GNDA.n1561 585
R1294 GNDA.n1521 GNDA.n1317 585
R1295 GNDA.n1317 GNDA.n1315 585
R1296 GNDA.n1520 GNDA.n1519 585
R1297 GNDA.n1519 GNDA.n1518 585
R1298 GNDA.n1513 GNDA.n1319 585
R1299 GNDA.n1517 GNDA.n1319 585
R1300 GNDA.n1515 GNDA.n1514 585
R1301 GNDA.n1516 GNDA.n1515 585
R1302 GNDA.n1512 GNDA.n1321 585
R1303 GNDA.n1321 GNDA.n1320 585
R1304 GNDA.n1511 GNDA.n1510 585
R1305 GNDA.n1510 GNDA.n1509 585
R1306 GNDA.n1323 GNDA.n1322 585
R1307 GNDA.n1328 GNDA.n1323 585
R1308 GNDA.n1327 GNDA.n1326 585
R1309 GNDA.n1324 GNDA.n248 585
R1310 GNDA.n1730 GNDA.n1729 585
R1311 GNDA.n1731 GNDA.n1730 585
R1312 GNDA.n1523 GNDA.n1522 585
R1313 GNDA.n1555 GNDA.n1523 585
R1314 GNDA.n1202 GNDA.n1201 585
R1315 GNDA.n1306 GNDA.n1202 585
R1316 GNDA.n1574 GNDA.n1573 585
R1317 GNDA.n1573 GNDA.n1572 585
R1318 GNDA.n1575 GNDA.n1199 585
R1319 GNDA.n1199 GNDA.n1198 585
R1320 GNDA.n1577 GNDA.n1576 585
R1321 GNDA.n1578 GNDA.n1577 585
R1322 GNDA.n1200 GNDA.n1197 585
R1323 GNDA.n1579 GNDA.n1197 585
R1324 GNDA.n1582 GNDA.n1581 585
R1325 GNDA.n1581 GNDA.n1580 585
R1326 GNDA.n1583 GNDA.n1195 585
R1327 GNDA.n1195 GNDA.n1194 585
R1328 GNDA.n1585 GNDA.n1584 585
R1329 GNDA.n1586 GNDA.n1585 585
R1330 GNDA.n1196 GNDA.n1190 585
R1331 GNDA.n1587 GNDA.n1190 585
R1332 GNDA.n1589 GNDA.n1192 585
R1333 GNDA.n1589 GNDA.n1588 585
R1334 GNDA.n1591 GNDA.n1590 585
R1335 GNDA.n1593 GNDA.n1592 585
R1336 GNDA.n1187 GNDA.n1186 585
R1337 GNDA.n1189 GNDA.n1187 585
R1338 GNDA.n1304 GNDA.n1303 585
R1339 GNDA.n1305 GNDA.n1304 585
R1340 GNDA.n1483 GNDA.n1476 531.201
R1341 GNDA.n1505 GNDA.n1476 528
R1342 GNDA.n2005 GNDA.n78 512
R1343 GNDA.n2005 GNDA.n2004 512
R1344 GNDA.n1988 GNDA.n1983 512
R1345 GNDA.n1988 GNDA.n1985 512
R1346 GNDA.n79 GNDA.n78 508.8
R1347 GNDA.n2004 GNDA.n79 508.8
R1348 GNDA.n1984 GNDA.n1983 508.8
R1349 GNDA.n1985 GNDA.n1984 508.8
R1350 GNDA.n1299 GNDA.n1204 505.748
R1351 GNDA.n1299 GNDA.n1298 505.748
R1352 GNDA.n1298 GNDA.n1297 505.748
R1353 GNDA.n1297 GNDA.n1208 505.748
R1354 GNDA.n1291 GNDA.n1208 505.748
R1355 GNDA.n1289 GNDA.n1288 505.748
R1356 GNDA.n1288 GNDA.n1287 505.748
R1357 GNDA.n1287 GNDA.n1212 505.748
R1358 GNDA.n1281 GNDA.n1212 505.748
R1359 GNDA.n1281 GNDA.n199 505.748
R1360 GNDA.n1274 GNDA.n200 505.748
R1361 GNDA.n1274 GNDA.n1273 505.748
R1362 GNDA.n1273 GNDA.n1272 505.748
R1363 GNDA.n1272 GNDA.n1263 505.748
R1364 GNDA.n1266 GNDA.n1263 505.748
R1365 GNDA.n1266 GNDA.n125 505.748
R1366 GNDA.n1940 GNDA.n1939 505.748
R1367 GNDA.n1939 GNDA.n1938 505.748
R1368 GNDA.n1938 GNDA.n130 505.748
R1369 GNDA.n1932 GNDA.n130 505.748
R1370 GNDA.n1932 GNDA.n1931 505.748
R1371 GNDA.n1057 GNDA.n134 505.748
R1372 GNDA.n1057 GNDA.n1056 505.748
R1373 GNDA.n1056 GNDA.n1055 505.748
R1374 GNDA.n1055 GNDA.n864 505.748
R1375 GNDA.n1049 GNDA.n864 505.748
R1376 GNDA.n1049 GNDA.n1048 505.748
R1377 GNDA.n1047 GNDA.n872 505.748
R1378 GNDA.n1041 GNDA.n872 505.748
R1379 GNDA.n1041 GNDA.n1040 505.748
R1380 GNDA.n1040 GNDA.n1039 505.748
R1381 GNDA.n1039 GNDA.n876 505.748
R1382 GNDA.n1483 GNDA.n1477 499.2
R1383 GNDA.n1806 GNDA.t72 496.098
R1384 GNDA.n2077 GNDA.n2060 487.086
R1385 GNDA.n2072 GNDA.n2060 487.086
R1386 GNDA.n2072 GNDA.n2071 487.086
R1387 GNDA.n2071 GNDA.n2070 487.086
R1388 GNDA.n2070 GNDA.n37 487.086
R1389 GNDA.n2157 GNDA.n2156 487.086
R1390 GNDA.n2157 GNDA.n33 487.086
R1391 GNDA.n2164 GNDA.n33 487.086
R1392 GNDA.n2165 GNDA.n2164 487.086
R1393 GNDA.n2166 GNDA.n2165 487.086
R1394 GNDA.n590 GNDA.n589 487.086
R1395 GNDA.n591 GNDA.n590 487.086
R1396 GNDA.n591 GNDA.n462 487.086
R1397 GNDA.n597 GNDA.n462 487.086
R1398 GNDA.n598 GNDA.n597 487.086
R1399 GNDA.n599 GNDA.n457 487.086
R1400 GNDA.n605 GNDA.n457 487.086
R1401 GNDA.n606 GNDA.n605 487.086
R1402 GNDA.n608 GNDA.n606 487.086
R1403 GNDA.n608 GNDA.n607 487.086
R1404 GNDA.n1015 GNDA.n886 487.086
R1405 GNDA.n1016 GNDA.n1015 487.086
R1406 GNDA.n1018 GNDA.n1016 487.086
R1407 GNDA.n1018 GNDA.n1017 487.086
R1408 GNDA.n1017 GNDA.n870 487.086
R1409 GNDA.n1025 GNDA.n871 487.086
R1410 GNDA.n1025 GNDA.n880 487.086
R1411 GNDA.n1031 GNDA.n880 487.086
R1412 GNDA.n1032 GNDA.n1031 487.086
R1413 GNDA.n1033 GNDA.n1032 487.086
R1414 GNDA.n1505 GNDA.n1504 486.401
R1415 GNDA.n1740 GNDA.n1739 467.039
R1416 GNDA.n1489 GNDA.n1482 444.8
R1417 GNDA.n1490 GNDA.n1489 444.8
R1418 GNDA.n1993 GNDA.n1992 444.695
R1419 GNDA.n1492 GNDA.n1482 441.601
R1420 GNDA.n1491 GNDA.n1490 438.401
R1421 GNDA.n1499 GNDA.n1498 435.2
R1422 GNDA.n1837 GNDA.n1835 434.906
R1423 GNDA.n1930 GNDA.n57 434.906
R1424 GNDA.n1499 GNDA.n1479 425.601
R1425 GNDA.n1503 GNDA.n1478 422.401
R1426 GNDA.n1503 GNDA.n1479 419.2
R1427 GNDA.n1956 GNDA.n64 406.401
R1428 GNDA.n2019 GNDA.n64 406.401
R1429 GNDA.n1992 GNDA.n1991 377.149
R1430 GNDA.n1554 GNDA.n1553 370.214
R1431 GNDA.n1732 GNDA.n246 370.214
R1432 GNDA.n1554 GNDA.n1155 365.957
R1433 GNDA.n1732 GNDA.n247 365.957
R1434 GNDA.n1338 GNDA.n241 354.67
R1435 GNDA.n1731 GNDA.n248 354.67
R1436 GNDA.n1592 GNDA.n1189 354.67
R1437 GNDA.n1808 GNDA.n1807 352.627
R1438 GNDA.n1819 GNDA.n1818 352.627
R1439 GNDA.n1821 GNDA.n1819 352.627
R1440 GNDA.n1821 GNDA.n1820 352.627
R1441 GNDA.n1820 GNDA.n203 352.627
R1442 GNDA.n1834 GNDA.n203 352.627
R1443 GNDA.n1838 GNDA.n1837 352.627
R1444 GNDA.n1838 GNDA.n194 352.627
R1445 GNDA.n1900 GNDA.n194 352.627
R1446 GNDA.n1901 GNDA.n1900 352.627
R1447 GNDA.n1903 GNDA.n1901 352.627
R1448 GNDA.n1903 GNDA.n1902 352.627
R1449 GNDA.n1914 GNDA.n1913 352.627
R1450 GNDA.n1916 GNDA.n1914 352.627
R1451 GNDA.n1916 GNDA.n1915 352.627
R1452 GNDA.n1915 GNDA.n135 352.627
R1453 GNDA.n1929 GNDA.n135 352.627
R1454 GNDA.n2028 GNDA.n57 352.627
R1455 GNDA.n2140 GNDA.n50 352.627
R1456 GNDA.n2141 GNDA.n2140 352.627
R1457 GNDA.n2142 GNDA.n2141 352.627
R1458 GNDA.n2142 GNDA.n38 352.627
R1459 GNDA.n2155 GNDA.n39 352.627
R1460 GNDA.n2058 GNDA.n39 352.627
R1461 GNDA.n2059 GNDA.n2058 352.627
R1462 GNDA.n2079 GNDA.n2059 352.627
R1463 GNDA.n2079 GNDA.n2078 352.627
R1464 GNDA.n2020 GNDA.n60 348.8
R1465 GNDA.n2024 GNDA.n60 348.8
R1466 GNDA.n1967 GNDA.n95 348.8
R1467 GNDA.n1963 GNDA.n95 348.8
R1468 GNDA.n1742 GNDA.n1741 343.452
R1469 GNDA.n1805 GNDA.n1804 343.452
R1470 GNDA.n1289 GNDA.t72 342.784
R1471 GNDA.n1940 GNDA.t68 342.784
R1472 GNDA.t70 GNDA.n1047 342.784
R1473 GNDA.n1458 GNDA.n245 337.111
R1474 GNDA.n1556 GNDA.n1555 337.111
R1475 GNDA.n1306 GNDA.n1305 337.111
R1476 GNDA.t70 GNDA.n461 172.876
R1477 GNDA.t70 GNDA.n869 172.876
R1478 GNDA.n1155 GNDA.t72 327.661
R1479 GNDA.n247 GNDA.t72 327.661
R1480 GNDA.t70 GNDA.n22 172.615
R1481 GNDA.t70 GNDA.n446 172.615
R1482 GNDA.n1553 GNDA.t72 323.404
R1483 GNDA.n246 GNDA.t72 323.404
R1484 GNDA.n2013 GNDA.n2012 323.2
R1485 GNDA.n2013 GNDA.n2010 316.8
R1486 GNDA.n1339 GNDA.n1338 316.043
R1487 GNDA.n1340 GNDA.n1339 316.043
R1488 GNDA.n1340 GNDA.n1330 316.043
R1489 GNDA.n1473 GNDA.n1331 316.043
R1490 GNDA.n1467 GNDA.n1466 316.043
R1491 GNDA.n1466 GNDA.n1465 316.043
R1492 GNDA.n1465 GNDA.n1345 316.043
R1493 GNDA.n1459 GNDA.n1345 316.043
R1494 GNDA.n1459 GNDA.n1458 316.043
R1495 GNDA.n1327 GNDA.n248 316.043
R1496 GNDA.n1328 GNDA.n1327 316.043
R1497 GNDA.n1509 GNDA.n1328 316.043
R1498 GNDA.n1516 GNDA.n1320 316.043
R1499 GNDA.n1518 GNDA.n1517 316.043
R1500 GNDA.n1518 GNDA.n1315 316.043
R1501 GNDA.n1562 GNDA.n1316 316.043
R1502 GNDA.n1556 GNDA.n1316 316.043
R1503 GNDA.n1592 GNDA.n1591 316.043
R1504 GNDA.n1588 GNDA.n1587 316.043
R1505 GNDA.n1587 GNDA.n1586 316.043
R1506 GNDA.n1586 GNDA.n1194 316.043
R1507 GNDA.n1580 GNDA.n1579 316.043
R1508 GNDA.n1579 GNDA.n1578 316.043
R1509 GNDA.n1578 GNDA.n1198 316.043
R1510 GNDA.n1572 GNDA.n1198 316.043
R1511 GNDA.n1555 GNDA.n1554 305.507
R1512 GNDA.n1737 GNDA.n244 304
R1513 GNDA.n1732 GNDA.n1731 301.995
R1514 GNDA.n1554 GNDA.n1189 301.995
R1515 GNDA.n1806 GNDA.n1805 301.474
R1516 GNDA.n1735 GNDA.n244 300.8
R1517 GNDA.n1737 GNDA.n1736 300.8
R1518 GNDA.n1736 GNDA.n1735 297.601
R1519 GNDA.n1310 GNDA.n1309 297.601
R1520 GNDA.n1568 GNDA.n1310 297.601
R1521 GNDA.n1567 GNDA.n1311 297.601
R1522 GNDA.n1313 GNDA.n1311 297.601
R1523 GNDA.n2012 GNDA.n2011 294.401
R1524 GNDA.n1953 GNDA.t88 292.584
R1525 GNDA.n65 GNDA.t94 292.584
R1526 GNDA.n61 GNDA.t76 292.584
R1527 GNDA.n62 GNDA.t85 292.584
R1528 GNDA.n1951 GNDA.t79 292.584
R1529 GNDA.n1952 GNDA.t82 292.584
R1530 GNDA.n1963 GNDA.n1962 292.5
R1531 GNDA.n1962 GNDA.n1961 292.5
R1532 GNDA.n1965 GNDA.n94 292.5
R1533 GNDA.n94 GNDA.n84 292.5
R1534 GNDA.n1968 GNDA.n1967 292.5
R1535 GNDA.n1969 GNDA.n1968 292.5
R1536 GNDA.n95 GNDA.n93 292.5
R1537 GNDA.n93 GNDA.n84 292.5
R1538 GNDA.n2019 GNDA.n2018 292.5
R1539 GNDA.n2018 GNDA.n2017 292.5
R1540 GNDA.n1954 GNDA.n68 292.5
R1541 GNDA.n1980 GNDA.n68 292.5
R1542 GNDA.n1959 GNDA.n1956 292.5
R1543 GNDA.n1960 GNDA.n1959 292.5
R1544 GNDA.n67 GNDA.n64 292.5
R1545 GNDA.n1980 GNDA.n67 292.5
R1546 GNDA.n2025 GNDA.n2024 292.5
R1547 GNDA.n2026 GNDA.n2025 292.5
R1548 GNDA.n2022 GNDA.n59 292.5
R1549 GNDA.n80 GNDA.n59 292.5
R1550 GNDA.n2020 GNDA.n63 292.5
R1551 GNDA.n2016 GNDA.n63 292.5
R1552 GNDA.n60 GNDA.n58 292.5
R1553 GNDA.n80 GNDA.n58 292.5
R1554 GNDA.n2000 GNDA.n1999 292.5
R1555 GNDA.n2001 GNDA.n2000 292.5
R1556 GNDA.n1998 GNDA.n83 292.5
R1557 GNDA.n1980 GNDA.n83 292.5
R1558 GNDA.n1997 GNDA.n1996 292.5
R1559 GNDA.n1996 GNDA.n1995 292.5
R1560 GNDA.n82 GNDA.n75 292.5
R1561 GNDA.n1980 GNDA.n82 292.5
R1562 GNDA.n1985 GNDA.n1982 292.5
R1563 GNDA.n1982 GNDA.n1981 292.5
R1564 GNDA.n1989 GNDA.n1988 292.5
R1565 GNDA.n1990 GNDA.n1989 292.5
R1566 GNDA.n1983 GNDA.n87 292.5
R1567 GNDA.n92 GNDA.n87 292.5
R1568 GNDA.n1984 GNDA.n86 292.5
R1569 GNDA.n1990 GNDA.n86 292.5
R1570 GNDA.n2004 GNDA.n2003 292.5
R1571 GNDA.n2003 GNDA.n2002 292.5
R1572 GNDA.n2005 GNDA.n70 292.5
R1573 GNDA.n2015 GNDA.n70 292.5
R1574 GNDA.n1978 GNDA.n78 292.5
R1575 GNDA.n1979 GNDA.n1978 292.5
R1576 GNDA.n79 GNDA.n71 292.5
R1577 GNDA.n2015 GNDA.n71 292.5
R1578 GNDA.n1957 GNDA.n74 292.5
R1579 GNDA.n1958 GNDA.n1957 292.5
R1580 GNDA.n1994 GNDA.n1993 292.5
R1581 GNDA.n1991 GNDA.n1990 292.5
R1582 GNDA.n2012 GNDA.n73 292.5
R1583 GNDA.n81 GNDA.n73 292.5
R1584 GNDA.n2011 GNDA.n69 292.5
R1585 GNDA.n2015 GNDA.n69 292.5
R1586 GNDA.n2010 GNDA.n72 292.5
R1587 GNDA.n1977 GNDA.n72 292.5
R1588 GNDA.n2014 GNDA.n2013 292.5
R1589 GNDA.n2015 GNDA.n2014 292.5
R1590 GNDA.n1312 GNDA.n1203 292.5
R1591 GNDA.n1571 GNDA.n1203 292.5
R1592 GNDA.n1314 GNDA.n1313 292.5
R1593 GNDA.n1314 GNDA.n1193 292.5
R1594 GNDA.n1565 GNDA.n1311 292.5
R1595 GNDA.n1565 GNDA.n1564 292.5
R1596 GNDA.n1567 GNDA.n1566 292.5
R1597 GNDA.n1566 GNDA.n1193 292.5
R1598 GNDA.n1735 GNDA.n1734 292.5
R1599 GNDA.n1734 GNDA.n1733 292.5
R1600 GNDA.n1736 GNDA.n243 292.5
R1601 GNDA.n1507 GNDA.n243 292.5
R1602 GNDA.n1738 GNDA.n1737 292.5
R1603 GNDA.n1739 GNDA.n1738 292.5
R1604 GNDA.n244 GNDA.n242 292.5
R1605 GNDA.n1507 GNDA.n242 292.5
R1606 GNDA.n1570 GNDA.n1569 292.5
R1607 GNDA.n1571 GNDA.n1570 292.5
R1608 GNDA.n1568 GNDA.n1308 292.5
R1609 GNDA.n1308 GNDA.n1193 292.5
R1610 GNDA.n1563 GNDA.n1310 292.5
R1611 GNDA.n1564 GNDA.n1563 292.5
R1612 GNDA.n1309 GNDA.n1307 292.5
R1613 GNDA.n1307 GNDA.n1193 292.5
R1614 GNDA.n1506 GNDA.n1505 292.5
R1615 GNDA.n1507 GNDA.n1506 292.5
R1616 GNDA.n1477 GNDA.n1475 292.5
R1617 GNDA.n1495 GNDA.n1475 292.5
R1618 GNDA.n1476 GNDA.n1474 292.5
R1619 GNDA.n1495 GNDA.n1474 292.5
R1620 GNDA.n1484 GNDA.n1483 292.5
R1621 GNDA.n1485 GNDA.n1484 292.5
R1622 GNDA.n1490 GNDA.n1481 292.5
R1623 GNDA.n1486 GNDA.n1481 292.5
R1624 GNDA.n1493 GNDA.n1492 292.5
R1625 GNDA.n1494 GNDA.n1493 292.5
R1626 GNDA.n1482 GNDA.n1480 292.5
R1627 GNDA.n1486 GNDA.n1480 292.5
R1628 GNDA.n1489 GNDA.n1488 292.5
R1629 GNDA.n1488 GNDA.n1487 292.5
R1630 GNDA.n1500 GNDA.n1499 292.5
R1631 GNDA.n1500 GNDA.n1329 292.5
R1632 GNDA.n1498 GNDA.n1497 292.5
R1633 GNDA.n1497 GNDA.n1496 292.5
R1634 GNDA.n1503 GNDA.n1502 292.5
R1635 GNDA.n1502 GNDA.n1329 292.5
R1636 GNDA.n1501 GNDA.n1479 292.5
R1637 GNDA.n1501 GNDA.n1193 292.5
R1638 GNDA.n1509 GNDA.n1508 291.462
R1639 GNDA.n1569 GNDA.n1309 291.2
R1640 GNDA.n1569 GNDA.n1568 291.2
R1641 GNDA.n1567 GNDA.n1312 291.2
R1642 GNDA.n1313 GNDA.n1312 291.2
R1643 GNDA.n2011 GNDA.n2010 288
R1644 GNDA.n1955 GNDA.n1954 288
R1645 GNDA.n1954 GNDA.n66 288
R1646 GNDA.n1564 GNDA.n1562 270.392
R1647 GNDA.n1969 GNDA.t80 262.5
R1648 GNDA.n2026 GNDA.t77 262.5
R1649 GNDA.n2101 GNDA.n2042 258.334
R1650 GNDA.n1856 GNDA.n176 258.334
R1651 GNDA.n1614 GNDA.n1168 258.334
R1652 GNDA.n518 GNDA.n496 258.334
R1653 GNDA.n723 GNDA.n705 258.334
R1654 GNDA.n941 GNDA.n901 258.334
R1655 GNDA.n1108 GNDA.n413 258.334
R1656 GNDA.n1760 GNDA.n218 258.334
R1657 GNDA.n309 GNDA.n264 258.334
R1658 GNDA.n1928 GNDA.n163 257.466
R1659 GNDA.n2076 GNDA.n2053 257.466
R1660 GNDA.n796 GNDA.n794 257.466
R1661 GNDA.n588 GNDA.n586 257.466
R1662 GNDA.n1083 GNDA.n1082 257.466
R1663 GNDA.n1010 GNDA.n887 257.466
R1664 GNDA.n1683 GNDA.n1154 257.466
R1665 GNDA.n1833 GNDA.n205 257.466
R1666 GNDA.n1714 GNDA.n356 257.466
R1667 GNDA.n2075 GNDA.n2062 254.442
R1668 GNDA.n2156 GNDA.t70 254.368
R1669 GNDA.n599 GNDA.t70 254.368
R1670 GNDA.t70 GNDA.n871 254.368
R1671 GNDA.n31 GNDA.n22 254.34
R1672 GNDA.n2173 GNDA.n22 254.34
R1673 GNDA.n28 GNDA.n22 254.34
R1674 GNDA.n2180 GNDA.n22 254.34
R1675 GNDA.n25 GNDA.n22 254.34
R1676 GNDA.n2187 GNDA.n22 254.34
R1677 GNDA.n859 GNDA.n19 254.34
R1678 GNDA.n856 GNDA.n19 254.34
R1679 GNDA.n850 GNDA.n19 254.34
R1680 GNDA.n847 GNDA.n19 254.34
R1681 GNDA.n841 GNDA.n19 254.34
R1682 GNDA.n919 GNDA.n19 254.34
R1683 GNDA.n1061 GNDA.n4 254.34
R1684 GNDA.n1067 GNDA.n4 254.34
R1685 GNDA.n853 GNDA.n4 254.34
R1686 GNDA.n1074 GNDA.n4 254.34
R1687 GNDA.n844 GNDA.n4 254.34
R1688 GNDA.n1081 GNDA.n4 254.34
R1689 GNDA.n828 GNDA.n19 254.34
R1690 GNDA.n825 GNDA.n19 254.34
R1691 GNDA.n813 GNDA.n19 254.34
R1692 GNDA.n811 GNDA.n19 254.34
R1693 GNDA.n801 GNDA.n19 254.34
R1694 GNDA.n799 GNDA.n19 254.34
R1695 GNDA.n662 GNDA.n4 254.34
R1696 GNDA.n821 GNDA.n4 254.34
R1697 GNDA.n817 GNDA.n4 254.34
R1698 GNDA.n807 GNDA.n4 254.34
R1699 GNDA.n805 GNDA.n4 254.34
R1700 GNDA.n795 GNDA.n4 254.34
R1701 GNDA.n482 GNDA.n461 254.34
R1702 GNDA.n557 GNDA.n461 254.34
R1703 GNDA.n559 GNDA.n461 254.34
R1704 GNDA.n571 GNDA.n461 254.34
R1705 GNDA.n469 GNDA.n461 254.34
R1706 GNDA.n466 GNDA.n461 254.34
R1707 GNDA.n614 GNDA.n446 254.34
R1708 GNDA.n453 GNDA.n446 254.34
R1709 GNDA.n621 GNDA.n446 254.34
R1710 GNDA.n450 GNDA.n446 254.34
R1711 GNDA.n628 GNDA.n446 254.34
R1712 GNDA.n631 GNDA.n446 254.34
R1713 GNDA.n922 GNDA.n869 254.34
R1714 GNDA.n984 GNDA.n869 254.34
R1715 GNDA.n986 GNDA.n869 254.34
R1716 GNDA.n996 GNDA.n869 254.34
R1717 GNDA.n998 GNDA.n869 254.34
R1718 GNDA.n1009 GNDA.n869 254.34
R1719 GNDA.n587 GNDA.n464 254.34
R1720 GNDA.n1013 GNDA.n1012 254.34
R1721 GNDA.n1595 GNDA.n1155 254.34
R1722 GNDA.n1657 GNDA.n1155 254.34
R1723 GNDA.n1659 GNDA.n1155 254.34
R1724 GNDA.n1669 GNDA.n1155 254.34
R1725 GNDA.n1671 GNDA.n1155 254.34
R1726 GNDA.n1682 GNDA.n1155 254.34
R1727 GNDA.n1436 GNDA.n246 254.34
R1728 GNDA.n1357 GNDA.n246 254.34
R1729 GNDA.n1443 GNDA.n246 254.34
R1730 GNDA.n1354 GNDA.n246 254.34
R1731 GNDA.n1450 GNDA.n246 254.34
R1732 GNDA.n1351 GNDA.n246 254.34
R1733 GNDA.n1726 GNDA.n247 254.34
R1734 GNDA.n333 GNDA.n247 254.34
R1735 GNDA.n330 GNDA.n247 254.34
R1736 GNDA.n344 GNDA.n247 254.34
R1737 GNDA.n354 GNDA.n247 254.34
R1738 GNDA.n1715 GNDA.n247 254.34
R1739 GNDA.n1553 GNDA.n1552 254.34
R1740 GNDA.n1553 GNDA.n1528 254.34
R1741 GNDA.n1553 GNDA.n1527 254.34
R1742 GNDA.n1553 GNDA.n1526 254.34
R1743 GNDA.n1553 GNDA.n1525 254.34
R1744 GNDA.n1553 GNDA.n1524 254.34
R1745 GNDA.n19 GNDA.n18 254.34
R1746 GNDA.n19 GNDA.n17 254.34
R1747 GNDA.n148 GNDA.n19 254.34
R1748 GNDA.n151 GNDA.n19 254.34
R1749 GNDA.n143 GNDA.n19 254.34
R1750 GNDA.n140 GNDA.n19 254.34
R1751 GNDA.n10 GNDA.n4 254.34
R1752 GNDA.n2201 GNDA.n4 254.34
R1753 GNDA.n4 GNDA.n3 254.34
R1754 GNDA.n155 GNDA.n4 254.34
R1755 GNDA.n146 GNDA.n4 254.34
R1756 GNDA.n162 GNDA.n4 254.34
R1757 GNDA.n1407 GNDA.n11 254.34
R1758 GNDA.n1413 GNDA.n1407 254.34
R1759 GNDA.n1420 GNDA.n1407 254.34
R1760 GNDA.n1411 GNDA.n1407 254.34
R1761 GNDA.n1427 GNDA.n1407 254.34
R1762 GNDA.n1430 GNDA.n1407 254.34
R1763 GNDA.n690 GNDA.n674 254.34
R1764 GNDA.n762 GNDA.n674 254.34
R1765 GNDA.n764 GNDA.n674 254.34
R1766 GNDA.n777 GNDA.n674 254.34
R1767 GNDA.n779 GNDA.n674 254.34
R1768 GNDA.n793 GNDA.n674 254.34
R1769 GNDA.n661 GNDA.n660 254.34
R1770 GNDA.n660 GNDA.n659 254.34
R1771 GNDA.n660 GNDA.n639 254.34
R1772 GNDA.n660 GNDA.n638 254.34
R1773 GNDA.n660 GNDA.n637 254.34
R1774 GNDA.n660 GNDA.n636 254.34
R1775 GNDA.n1149 GNDA.n1148 254.34
R1776 GNDA.n1148 GNDA.n1147 254.34
R1777 GNDA.n1148 GNDA.n396 254.34
R1778 GNDA.n1148 GNDA.n395 254.34
R1779 GNDA.n1148 GNDA.n394 254.34
R1780 GNDA.n1148 GNDA.n393 254.34
R1781 GNDA.n1402 GNDA.n202 254.34
R1782 GNDA.n1360 GNDA.n202 254.34
R1783 GNDA.n1389 GNDA.n202 254.34
R1784 GNDA.n1380 GNDA.n202 254.34
R1785 GNDA.n1378 GNDA.n202 254.34
R1786 GNDA.n1368 GNDA.n202 254.34
R1787 GNDA.n384 GNDA.n202 254.34
R1788 GNDA.n378 GNDA.n202 254.34
R1789 GNDA.n375 GNDA.n202 254.34
R1790 GNDA.n369 GNDA.n202 254.34
R1791 GNDA.n366 GNDA.n202 254.34
R1792 GNDA.n360 GNDA.n202 254.34
R1793 GNDA.n1258 GNDA.n202 254.34
R1794 GNDA.n1218 GNDA.n202 254.34
R1795 GNDA.n1246 GNDA.n202 254.34
R1796 GNDA.n1237 GNDA.n202 254.34
R1797 GNDA.n1235 GNDA.n202 254.34
R1798 GNDA.n1226 GNDA.n202 254.34
R1799 GNDA.n1396 GNDA.n201 254.34
R1800 GNDA.n1395 GNDA.n201 254.34
R1801 GNDA.n1362 GNDA.n201 254.34
R1802 GNDA.n1384 GNDA.n201 254.34
R1803 GNDA.n1374 GNDA.n201 254.34
R1804 GNDA.n1372 GNDA.n201 254.34
R1805 GNDA.n1693 GNDA.n201 254.34
R1806 GNDA.n381 GNDA.n201 254.34
R1807 GNDA.n1700 GNDA.n201 254.34
R1808 GNDA.n372 GNDA.n201 254.34
R1809 GNDA.n1707 GNDA.n201 254.34
R1810 GNDA.n363 GNDA.n201 254.34
R1811 GNDA.n1216 GNDA.n201 254.34
R1812 GNDA.n1252 GNDA.n201 254.34
R1813 GNDA.n1220 GNDA.n201 254.34
R1814 GNDA.n1241 GNDA.n201 254.34
R1815 GNDA.n1231 GNDA.n201 254.34
R1816 GNDA.n1229 GNDA.n201 254.34
R1817 GNDA.n1336 GNDA.n1334 254.34
R1818 GNDA.n1325 GNDA.n250 254.34
R1819 GNDA.n1191 GNDA.n1188 254.34
R1820 GNDA.n1741 GNDA.n89 251.865
R1821 GNDA.n2196 GNDA.n2195 251.614
R1822 GNDA.n2168 GNDA.n2167 251.614
R1823 GNDA.n832 GNDA.n831 251.614
R1824 GNDA.n613 GNDA.n454 251.614
R1825 GNDA.n1062 GNDA.n133 251.614
R1826 GNDA.n1034 GNDA.n877 251.614
R1827 GNDA.n1280 GNDA.n1279 251.614
R1828 GNDA.n1435 GNDA.n1358 251.614
R1829 GNDA.n1692 GNDA.n382 251.614
R1830 GNDA.n1947 GNDA.n1946 250.349
R1831 GNDA.n1818 GNDA.t72 239.004
R1832 GNDA.n1913 GNDA.t68 239.004
R1833 GNDA.t70 GNDA.n2155 239.004
R1834 GNDA.t70 GNDA.n37 232.719
R1835 GNDA.t70 GNDA.n598 232.719
R1836 GNDA.t70 GNDA.n870 232.719
R1837 GNDA.t41 GNDA.t24 225
R1838 GNDA.t43 GNDA.t55 225
R1839 GNDA.t55 GNDA.t105 225
R1840 GNDA.t33 GNDA.t45 225
R1841 GNDA.t45 GNDA.t12 225
R1842 GNDA.t28 GNDA.t99 225
R1843 GNDA.n2023 GNDA.n2022 224
R1844 GNDA.n2022 GNDA.n2021 224
R1845 GNDA.n1966 GNDA.n1965 224
R1846 GNDA.n1965 GNDA.n1964 224
R1847 GNDA.n1995 GNDA.t103 212.5
R1848 GNDA.n1733 GNDA.n245 200.161
R1849 GNDA.n1591 GNDA.t17 200.161
R1850 GNDA.n1571 GNDA.n1306 200.161
R1851 GNDA.t35 GNDA.n2001 200
R1852 GNDA.n1945 GNDA.n124 197
R1853 GNDA.n1369 GNDA.n198 195.049
R1854 GNDA.n139 GNDA.n55 195.049
R1855 GNDA.n688 GNDA.n359 195.049
R1856 GNDA.n798 GNDA.n15 195.049
R1857 GNDA.n1225 GNDA.n390 195.049
R1858 GNDA.n921 GNDA.n920 195.049
R1859 GNDA.n1594 GNDA.n1593 195.049
R1860 GNDA.n1337 GNDA.n239 195.049
R1861 GNDA.n1324 GNDA.n249 195.049
R1862 GNDA.n2028 GNDA.n2027 191.987
R1863 GNDA.n1403 GNDA.n388 187.249
R1864 GNDA.n2189 GNDA.n8 187.249
R1865 GNDA.n1689 GNDA.n385 187.249
R1866 GNDA.n829 GNDA.n20 187.249
R1867 GNDA.n1276 GNDA.n1259 187.249
R1868 GNDA.n1059 GNDA.n860 187.249
R1869 GNDA.n1304 GNDA.n1202 187.249
R1870 GNDA.n1457 GNDA.n1456 187.249
R1871 GNDA.n1557 GNDA.n1523 187.249
R1872 GNDA.n2099 GNDA.n2042 185
R1873 GNDA.n2042 GNDA.t91 185
R1874 GNDA.n2098 GNDA.n2097 185
R1875 GNDA.n2095 GNDA.n2043 185
R1876 GNDA.n2094 GNDA.n2044 185
R1877 GNDA.n2092 GNDA.n2091 185
R1878 GNDA.n2090 GNDA.n2045 185
R1879 GNDA.n2089 GNDA.n2088 185
R1880 GNDA.n2086 GNDA.n2046 185
R1881 GNDA.n2086 GNDA.t91 185
R1882 GNDA.n2085 GNDA.n2047 185
R1883 GNDA.n2101 GNDA.n2100 185
R1884 GNDA.n2103 GNDA.n2040 185
R1885 GNDA.n2105 GNDA.n2104 185
R1886 GNDA.n2106 GNDA.n2039 185
R1887 GNDA.n2108 GNDA.n2107 185
R1888 GNDA.n2110 GNDA.n2037 185
R1889 GNDA.n2112 GNDA.n2111 185
R1890 GNDA.n2113 GNDA.n2036 185
R1891 GNDA.n2115 GNDA.n2114 185
R1892 GNDA.n2117 GNDA.n2035 185
R1893 GNDA.n2119 GNDA.n2118 185
R1894 GNDA.n2121 GNDA.n2120 185
R1895 GNDA.n2124 GNDA.n2123 185
R1896 GNDA.n2125 GNDA.n2033 185
R1897 GNDA.n2127 GNDA.n2126 185
R1898 GNDA.n2129 GNDA.n2032 185
R1899 GNDA.n2131 GNDA.n2130 185
R1900 GNDA.n2133 GNDA.n2132 185
R1901 GNDA.n1855 GNDA.n176 185
R1902 GNDA.t73 GNDA.n176 185
R1903 GNDA.n1854 GNDA.n1853 185
R1904 GNDA.n1852 GNDA.n1851 185
R1905 GNDA.n1850 GNDA.n1849 185
R1906 GNDA.n1848 GNDA.n1847 185
R1907 GNDA.n1846 GNDA.n1845 185
R1908 GNDA.n1844 GNDA.n1843 185
R1909 GNDA.n1842 GNDA.n181 185
R1910 GNDA.t73 GNDA.n181 185
R1911 GNDA.n167 GNDA.n164 185
R1912 GNDA.n1857 GNDA.n1856 185
R1913 GNDA.n1859 GNDA.n1858 185
R1914 GNDA.n1861 GNDA.n1860 185
R1915 GNDA.n1863 GNDA.n1862 185
R1916 GNDA.n1865 GNDA.n1864 185
R1917 GNDA.n1867 GNDA.n1866 185
R1918 GNDA.n1869 GNDA.n1868 185
R1919 GNDA.n1871 GNDA.n1870 185
R1920 GNDA.n1873 GNDA.n1872 185
R1921 GNDA.n1875 GNDA.n1874 185
R1922 GNDA.n1877 GNDA.n1876 185
R1923 GNDA.n1879 GNDA.n1878 185
R1924 GNDA.n1881 GNDA.n1880 185
R1925 GNDA.n1883 GNDA.n1882 185
R1926 GNDA.n1885 GNDA.n1884 185
R1927 GNDA.n1887 GNDA.n1886 185
R1928 GNDA.n1889 GNDA.n1888 185
R1929 GNDA.n1891 GNDA.n1890 185
R1930 GNDA.n1613 GNDA.n1168 185
R1931 GNDA.t92 GNDA.n1168 185
R1932 GNDA.n1612 GNDA.n1611 185
R1933 GNDA.n1610 GNDA.n1609 185
R1934 GNDA.n1608 GNDA.n1607 185
R1935 GNDA.n1606 GNDA.n1605 185
R1936 GNDA.n1604 GNDA.n1603 185
R1937 GNDA.n1602 GNDA.n1601 185
R1938 GNDA.n1600 GNDA.n1173 185
R1939 GNDA.t92 GNDA.n1173 185
R1940 GNDA.n1599 GNDA.n1159 185
R1941 GNDA.n1615 GNDA.n1614 185
R1942 GNDA.n1617 GNDA.n1616 185
R1943 GNDA.n1619 GNDA.n1618 185
R1944 GNDA.n1621 GNDA.n1620 185
R1945 GNDA.n1623 GNDA.n1622 185
R1946 GNDA.n1625 GNDA.n1624 185
R1947 GNDA.n1627 GNDA.n1626 185
R1948 GNDA.n1629 GNDA.n1628 185
R1949 GNDA.n1631 GNDA.n1630 185
R1950 GNDA.n1633 GNDA.n1632 185
R1951 GNDA.n1635 GNDA.n1634 185
R1952 GNDA.n1637 GNDA.n1636 185
R1953 GNDA.n1639 GNDA.n1638 185
R1954 GNDA.n1641 GNDA.n1640 185
R1955 GNDA.n1643 GNDA.n1642 185
R1956 GNDA.n1645 GNDA.n1644 185
R1957 GNDA.n1647 GNDA.n1646 185
R1958 GNDA.n1649 GNDA.n1648 185
R1959 GNDA.n516 GNDA.n496 185
R1960 GNDA.n496 GNDA.t75 185
R1961 GNDA.n515 GNDA.n514 185
R1962 GNDA.n512 GNDA.n497 185
R1963 GNDA.n511 GNDA.n498 185
R1964 GNDA.n509 GNDA.n508 185
R1965 GNDA.n507 GNDA.n499 185
R1966 GNDA.n506 GNDA.n505 185
R1967 GNDA.n503 GNDA.n500 185
R1968 GNDA.n503 GNDA.t75 185
R1969 GNDA.n502 GNDA.n467 185
R1970 GNDA.n518 GNDA.n517 185
R1971 GNDA.n520 GNDA.n494 185
R1972 GNDA.n522 GNDA.n521 185
R1973 GNDA.n523 GNDA.n493 185
R1974 GNDA.n525 GNDA.n524 185
R1975 GNDA.n527 GNDA.n491 185
R1976 GNDA.n529 GNDA.n528 185
R1977 GNDA.n530 GNDA.n490 185
R1978 GNDA.n532 GNDA.n531 185
R1979 GNDA.n534 GNDA.n489 185
R1980 GNDA.n536 GNDA.n535 185
R1981 GNDA.n538 GNDA.n537 185
R1982 GNDA.n541 GNDA.n540 185
R1983 GNDA.n542 GNDA.n487 185
R1984 GNDA.n544 GNDA.n543 185
R1985 GNDA.n546 GNDA.n486 185
R1986 GNDA.n548 GNDA.n547 185
R1987 GNDA.n550 GNDA.n549 185
R1988 GNDA.n721 GNDA.n705 185
R1989 GNDA.n705 GNDA.t67 185
R1990 GNDA.n720 GNDA.n719 185
R1991 GNDA.n717 GNDA.n706 185
R1992 GNDA.n716 GNDA.n707 185
R1993 GNDA.n714 GNDA.n713 185
R1994 GNDA.n712 GNDA.n708 185
R1995 GNDA.n711 GNDA.n710 185
R1996 GNDA.n678 GNDA.n677 185
R1997 GNDA.t67 GNDA.n678 185
R1998 GNDA.n789 GNDA.n788 185
R1999 GNDA.n723 GNDA.n722 185
R2000 GNDA.n725 GNDA.n703 185
R2001 GNDA.n727 GNDA.n726 185
R2002 GNDA.n728 GNDA.n702 185
R2003 GNDA.n730 GNDA.n729 185
R2004 GNDA.n732 GNDA.n700 185
R2005 GNDA.n734 GNDA.n733 185
R2006 GNDA.n735 GNDA.n699 185
R2007 GNDA.n737 GNDA.n736 185
R2008 GNDA.n739 GNDA.n698 185
R2009 GNDA.n741 GNDA.n740 185
R2010 GNDA.n743 GNDA.n742 185
R2011 GNDA.n746 GNDA.n745 185
R2012 GNDA.n747 GNDA.n696 185
R2013 GNDA.n749 GNDA.n748 185
R2014 GNDA.n751 GNDA.n695 185
R2015 GNDA.n753 GNDA.n752 185
R2016 GNDA.n755 GNDA.n754 185
R2017 GNDA.n758 GNDA.n757 185
R2018 GNDA.n759 GNDA.n686 185
R2019 GNDA.n768 GNDA.n767 185
R2020 GNDA.n770 GNDA.n685 185
R2021 GNDA.n773 GNDA.n772 185
R2022 GNDA.n774 GNDA.n681 185
R2023 GNDA.n783 GNDA.n782 185
R2024 GNDA.n785 GNDA.n680 185
R2025 GNDA.n786 GNDA.n676 185
R2026 GNDA.n940 GNDA.n901 185
R2027 GNDA.t69 GNDA.n901 185
R2028 GNDA.n939 GNDA.n938 185
R2029 GNDA.n937 GNDA.n936 185
R2030 GNDA.n935 GNDA.n934 185
R2031 GNDA.n933 GNDA.n932 185
R2032 GNDA.n931 GNDA.n930 185
R2033 GNDA.n929 GNDA.n928 185
R2034 GNDA.n927 GNDA.n906 185
R2035 GNDA.t69 GNDA.n906 185
R2036 GNDA.n926 GNDA.n892 185
R2037 GNDA.n942 GNDA.n941 185
R2038 GNDA.n944 GNDA.n943 185
R2039 GNDA.n946 GNDA.n945 185
R2040 GNDA.n948 GNDA.n947 185
R2041 GNDA.n950 GNDA.n949 185
R2042 GNDA.n952 GNDA.n951 185
R2043 GNDA.n954 GNDA.n953 185
R2044 GNDA.n956 GNDA.n955 185
R2045 GNDA.n958 GNDA.n957 185
R2046 GNDA.n960 GNDA.n959 185
R2047 GNDA.n962 GNDA.n961 185
R2048 GNDA.n964 GNDA.n963 185
R2049 GNDA.n966 GNDA.n965 185
R2050 GNDA.n968 GNDA.n967 185
R2051 GNDA.n970 GNDA.n969 185
R2052 GNDA.n972 GNDA.n971 185
R2053 GNDA.n974 GNDA.n973 185
R2054 GNDA.n976 GNDA.n975 185
R2055 GNDA.n1106 GNDA.n413 185
R2056 GNDA.n413 GNDA.t93 185
R2057 GNDA.n1105 GNDA.n1104 185
R2058 GNDA.n1102 GNDA.n414 185
R2059 GNDA.n1101 GNDA.n415 185
R2060 GNDA.n1099 GNDA.n1098 185
R2061 GNDA.n1097 GNDA.n416 185
R2062 GNDA.n1096 GNDA.n1095 185
R2063 GNDA.n1093 GNDA.n417 185
R2064 GNDA.n1093 GNDA.t93 185
R2065 GNDA.n1092 GNDA.n418 185
R2066 GNDA.n1108 GNDA.n1107 185
R2067 GNDA.n1110 GNDA.n411 185
R2068 GNDA.n1112 GNDA.n1111 185
R2069 GNDA.n1113 GNDA.n410 185
R2070 GNDA.n1115 GNDA.n1114 185
R2071 GNDA.n1117 GNDA.n408 185
R2072 GNDA.n1119 GNDA.n1118 185
R2073 GNDA.n1120 GNDA.n407 185
R2074 GNDA.n1122 GNDA.n1121 185
R2075 GNDA.n1124 GNDA.n406 185
R2076 GNDA.n1126 GNDA.n1125 185
R2077 GNDA.n1128 GNDA.n1127 185
R2078 GNDA.n1131 GNDA.n1130 185
R2079 GNDA.n1132 GNDA.n404 185
R2080 GNDA.n1134 GNDA.n1133 185
R2081 GNDA.n1136 GNDA.n403 185
R2082 GNDA.n1138 GNDA.n1137 185
R2083 GNDA.n1140 GNDA.n1139 185
R2084 GNDA.n1141 GNDA.n399 185
R2085 GNDA.n1144 GNDA.n1143 185
R2086 GNDA.n426 GNDA.n401 185
R2087 GNDA.n429 GNDA.n425 185
R2088 GNDA.n434 GNDA.n433 185
R2089 GNDA.n437 GNDA.n436 185
R2090 GNDA.n423 GNDA.n420 185
R2091 GNDA.n442 GNDA.n419 185
R2092 GNDA.n1090 GNDA.n1089 185
R2093 GNDA.n978 GNDA.n977 185
R2094 GNDA.n981 GNDA.n980 185
R2095 GNDA.n979 GNDA.n915 185
R2096 GNDA.n990 GNDA.n989 185
R2097 GNDA.n992 GNDA.n991 185
R2098 GNDA.n993 GNDA.n910 185
R2099 GNDA.n1002 GNDA.n1001 185
R2100 GNDA.n912 GNDA.n891 185
R2101 GNDA.n1006 GNDA.n1005 185
R2102 GNDA.n553 GNDA.n552 185
R2103 GNDA.n554 GNDA.n477 185
R2104 GNDA.n563 GNDA.n562 185
R2105 GNDA.n565 GNDA.n476 185
R2106 GNDA.n568 GNDA.n567 185
R2107 GNDA.n473 GNDA.n472 185
R2108 GNDA.n576 GNDA.n575 185
R2109 GNDA.n579 GNDA.n578 185
R2110 GNDA.n471 GNDA.n468 185
R2111 GNDA.n1651 GNDA.n1650 185
R2112 GNDA.n1654 GNDA.n1653 185
R2113 GNDA.n1652 GNDA.n1182 185
R2114 GNDA.n1663 GNDA.n1662 185
R2115 GNDA.n1665 GNDA.n1664 185
R2116 GNDA.n1666 GNDA.n1177 185
R2117 GNDA.n1675 GNDA.n1674 185
R2118 GNDA.n1179 GNDA.n1158 185
R2119 GNDA.n1679 GNDA.n1678 185
R2120 GNDA.n1759 GNDA.n218 185
R2121 GNDA.t71 GNDA.n218 185
R2122 GNDA.n1758 GNDA.n1757 185
R2123 GNDA.n1756 GNDA.n1755 185
R2124 GNDA.n1754 GNDA.n1753 185
R2125 GNDA.n1752 GNDA.n1751 185
R2126 GNDA.n1750 GNDA.n1749 185
R2127 GNDA.n1748 GNDA.n1747 185
R2128 GNDA.n1746 GNDA.n223 185
R2129 GNDA.t71 GNDA.n223 185
R2130 GNDA.n209 GNDA.n206 185
R2131 GNDA.n1761 GNDA.n1760 185
R2132 GNDA.n1763 GNDA.n1762 185
R2133 GNDA.n1765 GNDA.n1764 185
R2134 GNDA.n1767 GNDA.n1766 185
R2135 GNDA.n1769 GNDA.n1768 185
R2136 GNDA.n1771 GNDA.n1770 185
R2137 GNDA.n1773 GNDA.n1772 185
R2138 GNDA.n1775 GNDA.n1774 185
R2139 GNDA.n1777 GNDA.n1776 185
R2140 GNDA.n1779 GNDA.n1778 185
R2141 GNDA.n1781 GNDA.n1780 185
R2142 GNDA.n1783 GNDA.n1782 185
R2143 GNDA.n1785 GNDA.n1784 185
R2144 GNDA.n1787 GNDA.n1786 185
R2145 GNDA.n1789 GNDA.n1788 185
R2146 GNDA.n1791 GNDA.n1790 185
R2147 GNDA.n1793 GNDA.n1792 185
R2148 GNDA.n1795 GNDA.n1794 185
R2149 GNDA.n1797 GNDA.n1796 185
R2150 GNDA.n1801 GNDA.n1800 185
R2151 GNDA.n1799 GNDA.n234 185
R2152 GNDA.n1812 GNDA.n1811 185
R2153 GNDA.n1814 GNDA.n1813 185
R2154 GNDA.n1815 GNDA.n227 185
R2155 GNDA.n1825 GNDA.n1824 185
R2156 GNDA.n229 GNDA.n208 185
R2157 GNDA.n1829 GNDA.n1828 185
R2158 GNDA.n311 GNDA.n264 185
R2159 GNDA.t74 GNDA.n264 185
R2160 GNDA.n313 GNDA.n312 185
R2161 GNDA.n315 GNDA.n314 185
R2162 GNDA.n317 GNDA.n316 185
R2163 GNDA.n319 GNDA.n318 185
R2164 GNDA.n321 GNDA.n320 185
R2165 GNDA.n323 GNDA.n322 185
R2166 GNDA.n324 GNDA.n269 185
R2167 GNDA.t74 GNDA.n269 185
R2168 GNDA.n325 GNDA.n273 185
R2169 GNDA.n310 GNDA.n309 185
R2170 GNDA.n308 GNDA.n307 185
R2171 GNDA.n306 GNDA.n305 185
R2172 GNDA.n304 GNDA.n303 185
R2173 GNDA.n302 GNDA.n301 185
R2174 GNDA.n300 GNDA.n299 185
R2175 GNDA.n298 GNDA.n297 185
R2176 GNDA.n296 GNDA.n295 185
R2177 GNDA.n294 GNDA.n293 185
R2178 GNDA.n292 GNDA.n291 185
R2179 GNDA.n290 GNDA.n289 185
R2180 GNDA.n288 GNDA.n287 185
R2181 GNDA.n286 GNDA.n285 185
R2182 GNDA.n284 GNDA.n283 185
R2183 GNDA.n282 GNDA.n281 185
R2184 GNDA.n280 GNDA.n279 185
R2185 GNDA.n278 GNDA.n277 185
R2186 GNDA.n276 GNDA.n254 185
R2187 GNDA.n1723 GNDA.n1722 185
R2188 GNDA.n334 GNDA.n255 185
R2189 GNDA.n332 GNDA.n331 185
R2190 GNDA.n341 GNDA.n340 185
R2191 GNDA.n339 GNDA.n329 185
R2192 GNDA.n348 GNDA.n347 185
R2193 GNDA.n350 GNDA.n349 185
R2194 GNDA.n351 GNDA.n274 185
R2195 GNDA.n1719 GNDA.n1718 185
R2196 GNDA.n1893 GNDA.n1892 185
R2197 GNDA.n1897 GNDA.n1896 185
R2198 GNDA.n1895 GNDA.n192 185
R2199 GNDA.n1907 GNDA.n1906 185
R2200 GNDA.n1909 GNDA.n1908 185
R2201 GNDA.n1910 GNDA.n185 185
R2202 GNDA.n1920 GNDA.n1919 185
R2203 GNDA.n187 GNDA.n166 185
R2204 GNDA.n1924 GNDA.n1923 185
R2205 GNDA.n2136 GNDA.n2135 185
R2206 GNDA.n2137 GNDA.n47 185
R2207 GNDA.n2146 GNDA.n2145 185
R2208 GNDA.n2148 GNDA.n46 185
R2209 GNDA.n2149 GNDA.n42 185
R2210 GNDA.n2152 GNDA.n2151 185
R2211 GNDA.n2054 GNDA.n44 185
R2212 GNDA.n2055 GNDA.n2049 185
R2213 GNDA.n2083 GNDA.n2082 185
R2214 GNDA.n1839 GNDA.n195 175.546
R2215 GNDA.n1899 GNDA.n195 175.546
R2216 GNDA.n1899 GNDA.n193 175.546
R2217 GNDA.n1904 GNDA.n193 175.546
R2218 GNDA.n1904 GNDA.n190 175.546
R2219 GNDA.n1912 GNDA.n190 175.546
R2220 GNDA.n1912 GNDA.n188 175.546
R2221 GNDA.n1917 GNDA.n188 175.546
R2222 GNDA.n1917 GNDA.n189 175.546
R2223 GNDA.n189 GNDA.n136 175.546
R2224 GNDA.n1928 GNDA.n136 175.546
R2225 GNDA.n1377 GNDA.n1367 175.546
R2226 GNDA.n1381 GNDA.n1379 175.546
R2227 GNDA.n1388 GNDA.n1363 175.546
R2228 GNDA.n1391 GNDA.n1390 175.546
R2229 GNDA.n1401 GNDA.n1400 175.546
R2230 GNDA.n1429 GNDA.n1428 175.546
R2231 GNDA.n1426 GNDA.n1409 175.546
R2232 GNDA.n1422 GNDA.n1421 175.546
R2233 GNDA.n1419 GNDA.n1412 175.546
R2234 GNDA.n1415 GNDA.n1414 175.546
R2235 GNDA.n161 GNDA.n138 175.546
R2236 GNDA.n157 GNDA.n156 175.546
R2237 GNDA.n154 GNDA.n147 175.546
R2238 GNDA.n2203 GNDA.n2202 175.546
R2239 GNDA.n2200 GNDA.n5 175.546
R2240 GNDA.n142 GNDA.n141 175.546
R2241 GNDA.n150 GNDA.n144 175.546
R2242 GNDA.n152 GNDA.n149 175.546
R2243 GNDA.n16 GNDA.n1 175.546
R2244 GNDA.n7 GNDA.n6 175.546
R2245 GNDA.n2029 GNDA.n51 175.546
R2246 GNDA.n2139 GNDA.n51 175.546
R2247 GNDA.n2139 GNDA.n49 175.546
R2248 GNDA.n2143 GNDA.n49 175.546
R2249 GNDA.n2143 GNDA.n40 175.546
R2250 GNDA.n2154 GNDA.n40 175.546
R2251 GNDA.n2154 GNDA.n41 175.546
R2252 GNDA.n2057 GNDA.n41 175.546
R2253 GNDA.n2057 GNDA.n2052 175.546
R2254 GNDA.n2080 GNDA.n2052 175.546
R2255 GNDA.n2080 GNDA.n2053 175.546
R2256 GNDA.n2074 GNDA.n2073 175.546
R2257 GNDA.n2073 GNDA.n2063 175.546
R2258 GNDA.n2069 GNDA.n2063 175.546
R2259 GNDA.n2069 GNDA.n2065 175.546
R2260 GNDA.n2065 GNDA.n36 175.546
R2261 GNDA.n2158 GNDA.n36 175.546
R2262 GNDA.n2158 GNDA.n34 175.546
R2263 GNDA.n2163 GNDA.n34 175.546
R2264 GNDA.n2163 GNDA.n32 175.546
R2265 GNDA.n2167 GNDA.n32 175.546
R2266 GNDA.n2186 GNDA.n23 175.546
R2267 GNDA.n2182 GNDA.n2181 175.546
R2268 GNDA.n2179 GNDA.n26 175.546
R2269 GNDA.n2175 GNDA.n2174 175.546
R2270 GNDA.n2172 GNDA.n29 175.546
R2271 GNDA.n761 GNDA.n691 175.546
R2272 GNDA.n765 GNDA.n763 175.546
R2273 GNDA.n776 GNDA.n683 175.546
R2274 GNDA.n780 GNDA.n778 175.546
R2275 GNDA.n792 GNDA.n675 175.546
R2276 GNDA.n365 GNDA.n361 175.546
R2277 GNDA.n368 GNDA.n367 175.546
R2278 GNDA.n374 GNDA.n370 175.546
R2279 GNDA.n377 GNDA.n376 175.546
R2280 GNDA.n383 GNDA.n379 175.546
R2281 GNDA.n644 GNDA.n643 175.546
R2282 GNDA.n648 GNDA.n647 175.546
R2283 GNDA.n652 GNDA.n651 175.546
R2284 GNDA.n654 GNDA.n640 175.546
R2285 GNDA.n658 GNDA.n635 175.546
R2286 GNDA.n804 GNDA.n671 175.546
R2287 GNDA.n808 GNDA.n806 175.546
R2288 GNDA.n816 GNDA.n667 175.546
R2289 GNDA.n822 GNDA.n818 175.546
R2290 GNDA.n820 GNDA.n819 175.546
R2291 GNDA.n630 GNDA.n629 175.546
R2292 GNDA.n627 GNDA.n448 175.546
R2293 GNDA.n623 GNDA.n622 175.546
R2294 GNDA.n620 GNDA.n451 175.546
R2295 GNDA.n616 GNDA.n615 175.546
R2296 GNDA.n592 GNDA.n465 175.546
R2297 GNDA.n592 GNDA.n463 175.546
R2298 GNDA.n596 GNDA.n463 175.546
R2299 GNDA.n596 GNDA.n460 175.546
R2300 GNDA.n600 GNDA.n460 175.546
R2301 GNDA.n600 GNDA.n458 175.546
R2302 GNDA.n604 GNDA.n458 175.546
R2303 GNDA.n604 GNDA.n456 175.546
R2304 GNDA.n609 GNDA.n456 175.546
R2305 GNDA.n609 GNDA.n454 175.546
R2306 GNDA.n556 GNDA.n479 175.546
R2307 GNDA.n560 GNDA.n558 175.546
R2308 GNDA.n570 GNDA.n474 175.546
R2309 GNDA.n573 GNDA.n572 175.546
R2310 GNDA.n582 GNDA.n581 175.546
R2311 GNDA.n802 GNDA.n800 175.546
R2312 GNDA.n810 GNDA.n669 175.546
R2313 GNDA.n814 GNDA.n812 175.546
R2314 GNDA.n824 GNDA.n665 175.546
R2315 GNDA.n827 GNDA.n826 175.546
R2316 GNDA.n1146 GNDA.n392 175.546
R2317 GNDA.n427 GNDA.n397 175.546
R2318 GNDA.n431 GNDA.n430 175.546
R2319 GNDA.n440 GNDA.n439 175.546
R2320 GNDA.n1087 GNDA.n1086 175.546
R2321 GNDA.n1234 GNDA.n1227 175.546
R2322 GNDA.n1238 GNDA.n1236 175.546
R2323 GNDA.n1245 GNDA.n1221 175.546
R2324 GNDA.n1248 GNDA.n1247 175.546
R2325 GNDA.n1257 GNDA.n1256 175.546
R2326 GNDA.n1275 GNDA.n1261 175.546
R2327 GNDA.n1271 GNDA.n1261 175.546
R2328 GNDA.n1271 GNDA.n1264 175.546
R2329 GNDA.n1267 GNDA.n1264 175.546
R2330 GNDA.n1267 GNDA.n128 175.546
R2331 GNDA.n1941 GNDA.n128 175.546
R2332 GNDA.n1941 GNDA.n129 175.546
R2333 GNDA.n1937 GNDA.n129 175.546
R2334 GNDA.n1937 GNDA.n131 175.546
R2335 GNDA.n1933 GNDA.n131 175.546
R2336 GNDA.n1933 GNDA.n133 175.546
R2337 GNDA.n1080 GNDA.n838 175.546
R2338 GNDA.n1076 GNDA.n1075 175.546
R2339 GNDA.n1073 GNDA.n845 175.546
R2340 GNDA.n1069 GNDA.n1068 175.546
R2341 GNDA.n1066 GNDA.n854 175.546
R2342 GNDA.n1058 GNDA.n862 175.546
R2343 GNDA.n1054 GNDA.n862 175.546
R2344 GNDA.n1054 GNDA.n865 175.546
R2345 GNDA.n1050 GNDA.n865 175.546
R2346 GNDA.n1050 GNDA.n868 175.546
R2347 GNDA.n1046 GNDA.n868 175.546
R2348 GNDA.n1046 GNDA.n873 175.546
R2349 GNDA.n1042 GNDA.n873 175.546
R2350 GNDA.n1042 GNDA.n875 175.546
R2351 GNDA.n1038 GNDA.n875 175.546
R2352 GNDA.n1038 GNDA.n877 175.546
R2353 GNDA.n1014 GNDA.n885 175.546
R2354 GNDA.n1019 GNDA.n885 175.546
R2355 GNDA.n1019 GNDA.n883 175.546
R2356 GNDA.n1023 GNDA.n883 175.546
R2357 GNDA.n1024 GNDA.n1023 175.546
R2358 GNDA.n1026 GNDA.n1024 175.546
R2359 GNDA.n1026 GNDA.n881 175.546
R2360 GNDA.n1030 GNDA.n881 175.546
R2361 GNDA.n1030 GNDA.n879 175.546
R2362 GNDA.n1034 GNDA.n879 175.546
R2363 GNDA.n983 GNDA.n917 175.546
R2364 GNDA.n987 GNDA.n985 175.546
R2365 GNDA.n995 GNDA.n913 175.546
R2366 GNDA.n999 GNDA.n997 175.546
R2367 GNDA.n1008 GNDA.n889 175.546
R2368 GNDA.n840 GNDA.n839 175.546
R2369 GNDA.n846 GNDA.n842 175.546
R2370 GNDA.n849 GNDA.n848 175.546
R2371 GNDA.n855 GNDA.n851 175.546
R2372 GNDA.n858 GNDA.n857 175.546
R2373 GNDA.n1590 GNDA.n1589 175.546
R2374 GNDA.n1589 GNDA.n1190 175.546
R2375 GNDA.n1585 GNDA.n1190 175.546
R2376 GNDA.n1585 GNDA.n1195 175.546
R2377 GNDA.n1581 GNDA.n1195 175.546
R2378 GNDA.n1581 GNDA.n1197 175.546
R2379 GNDA.n1577 GNDA.n1197 175.546
R2380 GNDA.n1577 GNDA.n1199 175.546
R2381 GNDA.n1573 GNDA.n1199 175.546
R2382 GNDA.n1573 GNDA.n1202 175.546
R2383 GNDA.n1656 GNDA.n1184 175.546
R2384 GNDA.n1660 GNDA.n1658 175.546
R2385 GNDA.n1668 GNDA.n1180 175.546
R2386 GNDA.n1672 GNDA.n1670 175.546
R2387 GNDA.n1681 GNDA.n1156 175.546
R2388 GNDA.n1232 GNDA.n1230 175.546
R2389 GNDA.n1240 GNDA.n1223 175.546
R2390 GNDA.n1243 GNDA.n1242 175.546
R2391 GNDA.n1251 GNDA.n1250 175.546
R2392 GNDA.n1254 GNDA.n1253 175.546
R2393 GNDA.n1300 GNDA.n1205 175.546
R2394 GNDA.n1300 GNDA.n1207 175.546
R2395 GNDA.n1296 GNDA.n1207 175.546
R2396 GNDA.n1296 GNDA.n1209 175.546
R2397 GNDA.n1292 GNDA.n1209 175.546
R2398 GNDA.n1292 GNDA.n1290 175.546
R2399 GNDA.n1290 GNDA.n1211 175.546
R2400 GNDA.n1286 GNDA.n1211 175.546
R2401 GNDA.n1286 GNDA.n1213 175.546
R2402 GNDA.n1282 GNDA.n1213 175.546
R2403 GNDA.n1282 GNDA.n1280 175.546
R2404 GNDA.n1341 GNDA.n1335 175.546
R2405 GNDA.n1341 GNDA.n1332 175.546
R2406 GNDA.n1472 GNDA.n1332 175.546
R2407 GNDA.n1472 GNDA.n1333 175.546
R2408 GNDA.n1468 GNDA.n1333 175.546
R2409 GNDA.n1468 GNDA.n1344 175.546
R2410 GNDA.n1464 GNDA.n1344 175.546
R2411 GNDA.n1464 GNDA.n1346 175.546
R2412 GNDA.n1460 GNDA.n1346 175.546
R2413 GNDA.n1460 GNDA.n1457 175.546
R2414 GNDA.n1743 GNDA.n236 175.546
R2415 GNDA.n1803 GNDA.n236 175.546
R2416 GNDA.n1803 GNDA.n235 175.546
R2417 GNDA.n1809 GNDA.n235 175.546
R2418 GNDA.n1809 GNDA.n232 175.546
R2419 GNDA.n1817 GNDA.n232 175.546
R2420 GNDA.n1817 GNDA.n230 175.546
R2421 GNDA.n1822 GNDA.n230 175.546
R2422 GNDA.n1822 GNDA.n231 175.546
R2423 GNDA.n231 GNDA.n204 175.546
R2424 GNDA.n1833 GNDA.n204 175.546
R2425 GNDA.n1375 GNDA.n1373 175.546
R2426 GNDA.n1383 GNDA.n1365 175.546
R2427 GNDA.n1386 GNDA.n1385 175.546
R2428 GNDA.n1394 GNDA.n1393 175.546
R2429 GNDA.n1398 GNDA.n1397 175.546
R2430 GNDA.n1452 GNDA.n1451 175.546
R2431 GNDA.n1449 GNDA.n1352 175.546
R2432 GNDA.n1445 GNDA.n1444 175.546
R2433 GNDA.n1442 GNDA.n1355 175.546
R2434 GNDA.n1438 GNDA.n1437 175.546
R2435 GNDA.n1326 GNDA.n1323 175.546
R2436 GNDA.n1510 GNDA.n1323 175.546
R2437 GNDA.n1510 GNDA.n1321 175.546
R2438 GNDA.n1515 GNDA.n1321 175.546
R2439 GNDA.n1515 GNDA.n1319 175.546
R2440 GNDA.n1519 GNDA.n1319 175.546
R2441 GNDA.n1519 GNDA.n1317 175.546
R2442 GNDA.n1561 GNDA.n1317 175.546
R2443 GNDA.n1561 GNDA.n1318 175.546
R2444 GNDA.n1557 GNDA.n1318 175.546
R2445 GNDA.n1534 GNDA.n1533 175.546
R2446 GNDA.n1538 GNDA.n1537 175.546
R2447 GNDA.n1542 GNDA.n1541 175.546
R2448 GNDA.n1546 GNDA.n1545 175.546
R2449 GNDA.n1551 GNDA.n1529 175.546
R2450 GNDA.n1709 GNDA.n1708 175.546
R2451 GNDA.n1706 GNDA.n364 175.546
R2452 GNDA.n1702 GNDA.n1701 175.546
R2453 GNDA.n1699 GNDA.n373 175.546
R2454 GNDA.n1695 GNDA.n1694 175.546
R2455 GNDA.n1725 GNDA.n252 175.546
R2456 GNDA.n337 GNDA.n336 175.546
R2457 GNDA.n345 GNDA.n343 175.546
R2458 GNDA.n353 GNDA.n327 175.546
R2459 GNDA.n1716 GNDA.n355 175.546
R2460 GNDA.t80 GNDA.n92 175
R2461 GNDA.n2002 GNDA.t77 175
R2462 GNDA.n674 GNDA.t68 172.876
R2463 GNDA.n1148 GNDA.t68 172.876
R2464 GNDA.n1407 GNDA.t68 172.615
R2465 GNDA.n660 GNDA.t68 172.615
R2466 GNDA.n1467 GNDA.t72 165.044
R2467 GNDA.n1517 GNDA.t72 165.044
R2468 GNDA.n1580 GNDA.t72 165.044
R2469 GNDA.n2135 GNDA.n2133 163.333
R2470 GNDA.n1892 GNDA.n1891 163.333
R2471 GNDA.n1650 GNDA.n1649 163.333
R2472 GNDA.n552 GNDA.n550 163.333
R2473 GNDA.n757 GNDA.n755 163.333
R2474 GNDA.n977 GNDA.n976 163.333
R2475 GNDA.n1141 GNDA.n1140 163.333
R2476 GNDA.n1796 GNDA.n1795 163.333
R2477 GNDA.n1722 GNDA.n254 163.333
R2478 GNDA.n1291 GNDA.t72 162.964
R2479 GNDA.n1048 GNDA.t70 162.964
R2480 GNDA.n1953 GNDA.t90 160.725
R2481 GNDA.n65 GNDA.t96 160.725
R2482 GNDA.n61 GNDA.t78 160.725
R2483 GNDA.n62 GNDA.t87 160.725
R2484 GNDA.n1951 GNDA.t81 160.725
R2485 GNDA.n1952 GNDA.t84 160.725
R2486 GNDA.n2027 GNDA.n50 160.642
R2487 GNDA.n120 GNDA.t7 157.555
R2488 GNDA.n121 GNDA.t18 157.555
R2489 GNDA.n116 GNDA.t50 153.294
R2490 GNDA.t72 GNDA.n1331 150.999
R2491 GNDA.t72 GNDA.n1516 150.999
R2492 GNDA.t72 GNDA.n1194 150.999
R2493 GNDA.n2146 GNDA.n47 150
R2494 GNDA.n2149 GNDA.n2148 150
R2495 GNDA.n2151 GNDA.n44 150
R2496 GNDA.n2083 GNDA.n2049 150
R2497 GNDA.n2130 GNDA.n2129 150
R2498 GNDA.n2127 GNDA.n2033 150
R2499 GNDA.n2123 GNDA.n2121 150
R2500 GNDA.n2118 GNDA.n2117 150
R2501 GNDA.n2115 GNDA.n2036 150
R2502 GNDA.n2111 GNDA.n2110 150
R2503 GNDA.n2108 GNDA.n2039 150
R2504 GNDA.n2104 GNDA.n2103 150
R2505 GNDA.n2086 GNDA.n2085 150
R2506 GNDA.n2088 GNDA.n2086 150
R2507 GNDA.n2092 GNDA.n2045 150
R2508 GNDA.n2095 GNDA.n2094 150
R2509 GNDA.n2097 GNDA.n2042 150
R2510 GNDA.n1896 GNDA.n1895 150
R2511 GNDA.n1908 GNDA.n1907 150
R2512 GNDA.n1920 GNDA.n185 150
R2513 GNDA.n1923 GNDA.n166 150
R2514 GNDA.n1888 GNDA.n1887 150
R2515 GNDA.n1884 GNDA.n1883 150
R2516 GNDA.n1880 GNDA.n1879 150
R2517 GNDA.n1876 GNDA.n1875 150
R2518 GNDA.n1872 GNDA.n1871 150
R2519 GNDA.n1868 GNDA.n1867 150
R2520 GNDA.n1864 GNDA.n1863 150
R2521 GNDA.n1860 GNDA.n1859 150
R2522 GNDA.n181 GNDA.n167 150
R2523 GNDA.n1843 GNDA.n181 150
R2524 GNDA.n1847 GNDA.n1846 150
R2525 GNDA.n1851 GNDA.n1850 150
R2526 GNDA.n1853 GNDA.n176 150
R2527 GNDA.n1653 GNDA.n1652 150
R2528 GNDA.n1664 GNDA.n1663 150
R2529 GNDA.n1675 GNDA.n1177 150
R2530 GNDA.n1678 GNDA.n1158 150
R2531 GNDA.n1646 GNDA.n1645 150
R2532 GNDA.n1642 GNDA.n1641 150
R2533 GNDA.n1638 GNDA.n1637 150
R2534 GNDA.n1634 GNDA.n1633 150
R2535 GNDA.n1630 GNDA.n1629 150
R2536 GNDA.n1626 GNDA.n1625 150
R2537 GNDA.n1622 GNDA.n1621 150
R2538 GNDA.n1618 GNDA.n1617 150
R2539 GNDA.n1173 GNDA.n1159 150
R2540 GNDA.n1601 GNDA.n1173 150
R2541 GNDA.n1605 GNDA.n1604 150
R2542 GNDA.n1609 GNDA.n1608 150
R2543 GNDA.n1611 GNDA.n1168 150
R2544 GNDA.n563 GNDA.n477 150
R2545 GNDA.n567 GNDA.n565 150
R2546 GNDA.n576 GNDA.n472 150
R2547 GNDA.n578 GNDA.n471 150
R2548 GNDA.n547 GNDA.n546 150
R2549 GNDA.n544 GNDA.n487 150
R2550 GNDA.n540 GNDA.n538 150
R2551 GNDA.n535 GNDA.n534 150
R2552 GNDA.n532 GNDA.n490 150
R2553 GNDA.n528 GNDA.n527 150
R2554 GNDA.n525 GNDA.n493 150
R2555 GNDA.n521 GNDA.n520 150
R2556 GNDA.n503 GNDA.n502 150
R2557 GNDA.n505 GNDA.n503 150
R2558 GNDA.n509 GNDA.n499 150
R2559 GNDA.n512 GNDA.n511 150
R2560 GNDA.n514 GNDA.n496 150
R2561 GNDA.n768 GNDA.n686 150
R2562 GNDA.n772 GNDA.n770 150
R2563 GNDA.n783 GNDA.n681 150
R2564 GNDA.n786 GNDA.n785 150
R2565 GNDA.n752 GNDA.n751 150
R2566 GNDA.n749 GNDA.n696 150
R2567 GNDA.n745 GNDA.n743 150
R2568 GNDA.n740 GNDA.n739 150
R2569 GNDA.n737 GNDA.n699 150
R2570 GNDA.n733 GNDA.n732 150
R2571 GNDA.n730 GNDA.n702 150
R2572 GNDA.n726 GNDA.n725 150
R2573 GNDA.n788 GNDA.n678 150
R2574 GNDA.n710 GNDA.n678 150
R2575 GNDA.n714 GNDA.n708 150
R2576 GNDA.n717 GNDA.n716 150
R2577 GNDA.n719 GNDA.n705 150
R2578 GNDA.n980 GNDA.n979 150
R2579 GNDA.n991 GNDA.n990 150
R2580 GNDA.n1002 GNDA.n910 150
R2581 GNDA.n1005 GNDA.n891 150
R2582 GNDA.n973 GNDA.n972 150
R2583 GNDA.n969 GNDA.n968 150
R2584 GNDA.n965 GNDA.n964 150
R2585 GNDA.n961 GNDA.n960 150
R2586 GNDA.n957 GNDA.n956 150
R2587 GNDA.n953 GNDA.n952 150
R2588 GNDA.n949 GNDA.n948 150
R2589 GNDA.n945 GNDA.n944 150
R2590 GNDA.n906 GNDA.n892 150
R2591 GNDA.n928 GNDA.n906 150
R2592 GNDA.n932 GNDA.n931 150
R2593 GNDA.n936 GNDA.n935 150
R2594 GNDA.n938 GNDA.n901 150
R2595 GNDA.n1143 GNDA.n401 150
R2596 GNDA.n434 GNDA.n425 150
R2597 GNDA.n436 GNDA.n423 150
R2598 GNDA.n1090 GNDA.n419 150
R2599 GNDA.n1137 GNDA.n1136 150
R2600 GNDA.n1134 GNDA.n404 150
R2601 GNDA.n1130 GNDA.n1128 150
R2602 GNDA.n1125 GNDA.n1124 150
R2603 GNDA.n1122 GNDA.n407 150
R2604 GNDA.n1118 GNDA.n1117 150
R2605 GNDA.n1115 GNDA.n410 150
R2606 GNDA.n1111 GNDA.n1110 150
R2607 GNDA.n1093 GNDA.n1092 150
R2608 GNDA.n1095 GNDA.n1093 150
R2609 GNDA.n1099 GNDA.n416 150
R2610 GNDA.n1102 GNDA.n1101 150
R2611 GNDA.n1104 GNDA.n413 150
R2612 GNDA.n1800 GNDA.n1799 150
R2613 GNDA.n1813 GNDA.n1812 150
R2614 GNDA.n1825 GNDA.n227 150
R2615 GNDA.n1828 GNDA.n208 150
R2616 GNDA.n1792 GNDA.n1791 150
R2617 GNDA.n1788 GNDA.n1787 150
R2618 GNDA.n1784 GNDA.n1783 150
R2619 GNDA.n1780 GNDA.n1779 150
R2620 GNDA.n1776 GNDA.n1775 150
R2621 GNDA.n1772 GNDA.n1771 150
R2622 GNDA.n1768 GNDA.n1767 150
R2623 GNDA.n1764 GNDA.n1763 150
R2624 GNDA.n223 GNDA.n209 150
R2625 GNDA.n1747 GNDA.n223 150
R2626 GNDA.n1751 GNDA.n1750 150
R2627 GNDA.n1755 GNDA.n1754 150
R2628 GNDA.n1757 GNDA.n218 150
R2629 GNDA.n331 GNDA.n255 150
R2630 GNDA.n340 GNDA.n339 150
R2631 GNDA.n349 GNDA.n348 150
R2632 GNDA.n1719 GNDA.n274 150
R2633 GNDA.n279 GNDA.n278 150
R2634 GNDA.n283 GNDA.n282 150
R2635 GNDA.n287 GNDA.n286 150
R2636 GNDA.n291 GNDA.n290 150
R2637 GNDA.n295 GNDA.n294 150
R2638 GNDA.n299 GNDA.n298 150
R2639 GNDA.n303 GNDA.n302 150
R2640 GNDA.n307 GNDA.n306 150
R2641 GNDA.n273 GNDA.n269 150
R2642 GNDA.n322 GNDA.n269 150
R2643 GNDA.n320 GNDA.n319 150
R2644 GNDA.n316 GNDA.n315 150
R2645 GNDA.n312 GNDA.n264 150
R2646 GNDA.t2 GNDA.t23 150
R2647 GNDA.t98 GNDA.t27 150
R2648 GNDA.t65 GNDA.t64 150
R2649 GNDA.t52 GNDA.t26 150
R2650 GNDA.n1992 GNDA.n74 149.181
R2651 GNDA.n118 GNDA.t20 148.906
R2652 GNDA.n118 GNDA.t31 148.653
R2653 GNDA.n1742 GNDA.n1740 145.013
R2654 GNDA.t5 GNDA.t37 140.464
R2655 GNDA.n98 GNDA.n96 140.077
R2656 GNDA.n114 GNDA.n113 139.077
R2657 GNDA.n112 GNDA.n111 139.077
R2658 GNDA.n110 GNDA.n109 139.077
R2659 GNDA.n108 GNDA.n107 139.077
R2660 GNDA.n106 GNDA.n105 139.077
R2661 GNDA.n104 GNDA.n103 139.077
R2662 GNDA.n102 GNDA.n101 139.077
R2663 GNDA.n100 GNDA.n99 139.077
R2664 GNDA.n98 GNDA.n97 139.077
R2665 GNDA.n1431 GNDA.n388 126.782
R2666 GNDA.n2189 GNDA.n2188 126.782
R2667 GNDA.n1689 GNDA.n387 126.782
R2668 GNDA.n632 GNDA.n20 126.782
R2669 GNDA.n1276 GNDA.n1275 126.782
R2670 GNDA.n1059 GNDA.n1058 126.782
R2671 GNDA.n1304 GNDA.n1205 126.782
R2672 GNDA.n1456 GNDA.n1349 126.782
R2673 GNDA.n1530 GNDA.n1523 126.782
R2674 GNDA.t57 GNDA.t40 125.001
R2675 GNDA.t83 GNDA.t15 125.001
R2676 GNDA.t63 GNDA.t86 125.001
R2677 GNDA.t66 GNDA.t47 125.001
R2678 GNDA.n1839 GNDA.n198 124.832
R2679 GNDA.n2029 GNDA.n55 124.832
R2680 GNDA.n689 GNDA.n688 124.832
R2681 GNDA.n483 GNDA.n15 124.832
R2682 GNDA.n1150 GNDA.n390 124.832
R2683 GNDA.n923 GNDA.n921 124.832
R2684 GNDA.n1596 GNDA.n1594 124.832
R2685 GNDA.n1743 GNDA.n239 124.832
R2686 GNDA.n1727 GNDA.n249 124.832
R2687 GNDA.n1487 GNDA.t16 121.787
R2688 GNDA.n2024 GNDA.n2023 118.4
R2689 GNDA.n2021 GNDA.n2020 118.4
R2690 GNDA.n2019 GNDA.n66 118.4
R2691 GNDA.n1956 GNDA.n1955 118.4
R2692 GNDA.n1967 GNDA.n1966 118.4
R2693 GNDA.n1964 GNDA.n1963 118.4
R2694 GNDA.t6 GNDA.t30 117.858
R2695 GNDA.n1572 GNDA.n1571 115.882
R2696 GNDA.n1807 GNDA.t72 113.624
R2697 GNDA.n1902 GNDA.t68 113.624
R2698 GNDA.t70 GNDA.n38 113.624
R2699 GNDA.t60 GNDA.n84 112.501
R2700 GNDA.t89 GNDA.t14 112.501
R2701 GNDA.t14 GNDA.t0 112.501
R2702 GNDA.t0 GNDA.n1958 112.501
R2703 GNDA.n1958 GNDA.t43 112.501
R2704 GNDA.t12 GNDA.n1977 112.501
R2705 GNDA.n1977 GNDA.t10 112.501
R2706 GNDA.t10 GNDA.t51 112.501
R2707 GNDA.t51 GNDA.t95 112.501
R2708 GNDA.n80 GNDA.t101 112.501
R2709 GNDA.n2027 GNDA.n2026 112.501
R2710 GNDA.n1946 GNDA.t68 112.388
R2711 GNDA.n1733 GNDA.n1732 105.347
R2712 GNDA.n1930 GNDA.n19 103.144
R2713 GNDA.n1835 GNDA.n202 103.144
R2714 GNDA.t24 GNDA.n1994 100.001
R2715 GNDA.t40 GNDA.t60 100.001
R2716 GNDA.t15 GNDA.t53 100.001
R2717 GNDA.t21 GNDA.t63 100.001
R2718 GNDA.t101 GNDA.t66 100.001
R2719 GNDA.t99 GNDA.n81 100.001
R2720 GNDA.n1930 GNDA.n4 99.6276
R2721 GNDA.n1835 GNDA.n201 99.6276
R2722 GNDA.t5 GNDA.n1330 94.813
R2723 GNDA.t19 GNDA.t8 94.2862
R2724 GNDA.n1804 GNDA.n89 91.5877
R2725 GNDA.t68 GNDA.n4 91.423
R2726 GNDA.t72 GNDA.n201 91.423
R2727 GNDA.n1961 GNDA.t3 87.5005
R2728 GNDA.n2016 GNDA.t38 87.5005
R2729 GNDA.n2006 GNDA.n77 85.2842
R2730 GNDA.n1987 GNDA.n1986 85.2842
R2731 GNDA.n1947 GNDA.n124 84.306
R2732 GNDA.n1496 GNDA.n1494 78.5719
R2733 GNDA.n1368 GNDA.n1367 76.3222
R2734 GNDA.n1379 GNDA.n1378 76.3222
R2735 GNDA.n1380 GNDA.n1363 76.3222
R2736 GNDA.n1391 GNDA.n1389 76.3222
R2737 GNDA.n1400 GNDA.n1360 76.3222
R2738 GNDA.n1403 GNDA.n1402 76.3222
R2739 GNDA.n1430 GNDA.n1429 76.3222
R2740 GNDA.n1427 GNDA.n1426 76.3222
R2741 GNDA.n1422 GNDA.n1411 76.3222
R2742 GNDA.n1420 GNDA.n1419 76.3222
R2743 GNDA.n1415 GNDA.n1413 76.3222
R2744 GNDA.n2195 GNDA.n11 76.3222
R2745 GNDA.n162 GNDA.n161 76.3222
R2746 GNDA.n157 GNDA.n146 76.3222
R2747 GNDA.n155 GNDA.n154 76.3222
R2748 GNDA.n2203 GNDA.n3 76.3222
R2749 GNDA.n2201 GNDA.n2200 76.3222
R2750 GNDA.n2196 GNDA.n10 76.3222
R2751 GNDA.n140 GNDA.n139 76.3222
R2752 GNDA.n143 GNDA.n142 76.3222
R2753 GNDA.n151 GNDA.n150 76.3222
R2754 GNDA.n149 GNDA.n148 76.3222
R2755 GNDA.n17 GNDA.n16 76.3222
R2756 GNDA.n18 GNDA.n8 76.3222
R2757 GNDA.n2075 GNDA.n2074 76.3222
R2758 GNDA.n2187 GNDA.n2186 76.3222
R2759 GNDA.n2182 GNDA.n25 76.3222
R2760 GNDA.n2180 GNDA.n2179 76.3222
R2761 GNDA.n2175 GNDA.n28 76.3222
R2762 GNDA.n2173 GNDA.n2172 76.3222
R2763 GNDA.n2168 GNDA.n31 76.3222
R2764 GNDA.n31 GNDA.n29 76.3222
R2765 GNDA.n2174 GNDA.n2173 76.3222
R2766 GNDA.n28 GNDA.n26 76.3222
R2767 GNDA.n2181 GNDA.n2180 76.3222
R2768 GNDA.n25 GNDA.n23 76.3222
R2769 GNDA.n2188 GNDA.n2187 76.3222
R2770 GNDA.n690 GNDA.n689 76.3222
R2771 GNDA.n762 GNDA.n761 76.3222
R2772 GNDA.n765 GNDA.n764 76.3222
R2773 GNDA.n777 GNDA.n776 76.3222
R2774 GNDA.n780 GNDA.n779 76.3222
R2775 GNDA.n793 GNDA.n792 76.3222
R2776 GNDA.n361 GNDA.n360 76.3222
R2777 GNDA.n367 GNDA.n366 76.3222
R2778 GNDA.n370 GNDA.n369 76.3222
R2779 GNDA.n376 GNDA.n375 76.3222
R2780 GNDA.n379 GNDA.n378 76.3222
R2781 GNDA.n385 GNDA.n384 76.3222
R2782 GNDA.n643 GNDA.n636 76.3222
R2783 GNDA.n647 GNDA.n637 76.3222
R2784 GNDA.n651 GNDA.n638 76.3222
R2785 GNDA.n654 GNDA.n639 76.3222
R2786 GNDA.n659 GNDA.n658 76.3222
R2787 GNDA.n832 GNDA.n661 76.3222
R2788 GNDA.n795 GNDA.n671 76.3222
R2789 GNDA.n806 GNDA.n805 76.3222
R2790 GNDA.n807 GNDA.n667 76.3222
R2791 GNDA.n818 GNDA.n817 76.3222
R2792 GNDA.n821 GNDA.n820 76.3222
R2793 GNDA.n831 GNDA.n662 76.3222
R2794 GNDA.n631 GNDA.n630 76.3222
R2795 GNDA.n628 GNDA.n627 76.3222
R2796 GNDA.n623 GNDA.n450 76.3222
R2797 GNDA.n621 GNDA.n620 76.3222
R2798 GNDA.n616 GNDA.n453 76.3222
R2799 GNDA.n614 GNDA.n613 76.3222
R2800 GNDA.n588 GNDA.n587 76.3222
R2801 GNDA.n482 GNDA.n479 76.3222
R2802 GNDA.n558 GNDA.n557 76.3222
R2803 GNDA.n559 GNDA.n474 76.3222
R2804 GNDA.n573 GNDA.n571 76.3222
R2805 GNDA.n581 GNDA.n469 76.3222
R2806 GNDA.n586 GNDA.n466 76.3222
R2807 GNDA.n799 GNDA.n798 76.3222
R2808 GNDA.n802 GNDA.n801 76.3222
R2809 GNDA.n811 GNDA.n810 76.3222
R2810 GNDA.n814 GNDA.n813 76.3222
R2811 GNDA.n825 GNDA.n824 76.3222
R2812 GNDA.n829 GNDA.n828 76.3222
R2813 GNDA.n1150 GNDA.n1149 76.3222
R2814 GNDA.n1147 GNDA.n1146 76.3222
R2815 GNDA.n427 GNDA.n396 76.3222
R2816 GNDA.n430 GNDA.n395 76.3222
R2817 GNDA.n440 GNDA.n394 76.3222
R2818 GNDA.n1087 GNDA.n393 76.3222
R2819 GNDA.n1227 GNDA.n1226 76.3222
R2820 GNDA.n1236 GNDA.n1235 76.3222
R2821 GNDA.n1237 GNDA.n1221 76.3222
R2822 GNDA.n1248 GNDA.n1246 76.3222
R2823 GNDA.n1256 GNDA.n1218 76.3222
R2824 GNDA.n1259 GNDA.n1258 76.3222
R2825 GNDA.n1081 GNDA.n1080 76.3222
R2826 GNDA.n1076 GNDA.n844 76.3222
R2827 GNDA.n1074 GNDA.n1073 76.3222
R2828 GNDA.n1069 GNDA.n853 76.3222
R2829 GNDA.n1067 GNDA.n1066 76.3222
R2830 GNDA.n1062 GNDA.n1061 76.3222
R2831 GNDA.n1014 GNDA.n1013 76.3222
R2832 GNDA.n923 GNDA.n922 76.3222
R2833 GNDA.n984 GNDA.n983 76.3222
R2834 GNDA.n987 GNDA.n986 76.3222
R2835 GNDA.n996 GNDA.n995 76.3222
R2836 GNDA.n999 GNDA.n998 76.3222
R2837 GNDA.n1009 GNDA.n1008 76.3222
R2838 GNDA.n920 GNDA.n919 76.3222
R2839 GNDA.n841 GNDA.n840 76.3222
R2840 GNDA.n847 GNDA.n846 76.3222
R2841 GNDA.n850 GNDA.n849 76.3222
R2842 GNDA.n856 GNDA.n855 76.3222
R2843 GNDA.n859 GNDA.n858 76.3222
R2844 GNDA.n860 GNDA.n859 76.3222
R2845 GNDA.n857 GNDA.n856 76.3222
R2846 GNDA.n851 GNDA.n850 76.3222
R2847 GNDA.n848 GNDA.n847 76.3222
R2848 GNDA.n842 GNDA.n841 76.3222
R2849 GNDA.n919 GNDA.n839 76.3222
R2850 GNDA.n1061 GNDA.n854 76.3222
R2851 GNDA.n1068 GNDA.n1067 76.3222
R2852 GNDA.n853 GNDA.n845 76.3222
R2853 GNDA.n1075 GNDA.n1074 76.3222
R2854 GNDA.n844 GNDA.n838 76.3222
R2855 GNDA.n1082 GNDA.n1081 76.3222
R2856 GNDA.n828 GNDA.n827 76.3222
R2857 GNDA.n826 GNDA.n825 76.3222
R2858 GNDA.n813 GNDA.n665 76.3222
R2859 GNDA.n812 GNDA.n811 76.3222
R2860 GNDA.n801 GNDA.n669 76.3222
R2861 GNDA.n800 GNDA.n799 76.3222
R2862 GNDA.n819 GNDA.n662 76.3222
R2863 GNDA.n822 GNDA.n821 76.3222
R2864 GNDA.n817 GNDA.n816 76.3222
R2865 GNDA.n808 GNDA.n807 76.3222
R2866 GNDA.n805 GNDA.n804 76.3222
R2867 GNDA.n796 GNDA.n795 76.3222
R2868 GNDA.n483 GNDA.n482 76.3222
R2869 GNDA.n557 GNDA.n556 76.3222
R2870 GNDA.n560 GNDA.n559 76.3222
R2871 GNDA.n571 GNDA.n570 76.3222
R2872 GNDA.n572 GNDA.n469 76.3222
R2873 GNDA.n582 GNDA.n466 76.3222
R2874 GNDA.n615 GNDA.n614 76.3222
R2875 GNDA.n453 GNDA.n451 76.3222
R2876 GNDA.n622 GNDA.n621 76.3222
R2877 GNDA.n450 GNDA.n448 76.3222
R2878 GNDA.n629 GNDA.n628 76.3222
R2879 GNDA.n632 GNDA.n631 76.3222
R2880 GNDA.n922 GNDA.n917 76.3222
R2881 GNDA.n985 GNDA.n984 76.3222
R2882 GNDA.n986 GNDA.n913 76.3222
R2883 GNDA.n997 GNDA.n996 76.3222
R2884 GNDA.n998 GNDA.n889 76.3222
R2885 GNDA.n1010 GNDA.n1009 76.3222
R2886 GNDA.n587 GNDA.n465 76.3222
R2887 GNDA.n1013 GNDA.n887 76.3222
R2888 GNDA.n1590 GNDA.n1188 76.3222
R2889 GNDA.n1596 GNDA.n1595 76.3222
R2890 GNDA.n1657 GNDA.n1656 76.3222
R2891 GNDA.n1660 GNDA.n1659 76.3222
R2892 GNDA.n1669 GNDA.n1668 76.3222
R2893 GNDA.n1672 GNDA.n1671 76.3222
R2894 GNDA.n1682 GNDA.n1681 76.3222
R2895 GNDA.n1230 GNDA.n1229 76.3222
R2896 GNDA.n1231 GNDA.n1223 76.3222
R2897 GNDA.n1242 GNDA.n1241 76.3222
R2898 GNDA.n1250 GNDA.n1220 76.3222
R2899 GNDA.n1254 GNDA.n1252 76.3222
R2900 GNDA.n1279 GNDA.n1216 76.3222
R2901 GNDA.n1595 GNDA.n1184 76.3222
R2902 GNDA.n1658 GNDA.n1657 76.3222
R2903 GNDA.n1659 GNDA.n1180 76.3222
R2904 GNDA.n1670 GNDA.n1669 76.3222
R2905 GNDA.n1671 GNDA.n1156 76.3222
R2906 GNDA.n1683 GNDA.n1682 76.3222
R2907 GNDA.n1336 GNDA.n1335 76.3222
R2908 GNDA.n1373 GNDA.n1372 76.3222
R2909 GNDA.n1374 GNDA.n1365 76.3222
R2910 GNDA.n1385 GNDA.n1384 76.3222
R2911 GNDA.n1393 GNDA.n1362 76.3222
R2912 GNDA.n1398 GNDA.n1395 76.3222
R2913 GNDA.n1396 GNDA.n1358 76.3222
R2914 GNDA.n1452 GNDA.n1351 76.3222
R2915 GNDA.n1450 GNDA.n1449 76.3222
R2916 GNDA.n1445 GNDA.n1354 76.3222
R2917 GNDA.n1443 GNDA.n1442 76.3222
R2918 GNDA.n1438 GNDA.n1357 76.3222
R2919 GNDA.n1436 GNDA.n1435 76.3222
R2920 GNDA.n1437 GNDA.n1436 76.3222
R2921 GNDA.n1357 GNDA.n1355 76.3222
R2922 GNDA.n1444 GNDA.n1443 76.3222
R2923 GNDA.n1354 GNDA.n1352 76.3222
R2924 GNDA.n1451 GNDA.n1450 76.3222
R2925 GNDA.n1351 GNDA.n1349 76.3222
R2926 GNDA.n1326 GNDA.n1325 76.3222
R2927 GNDA.n1530 GNDA.n1524 76.3222
R2928 GNDA.n1534 GNDA.n1525 76.3222
R2929 GNDA.n1538 GNDA.n1526 76.3222
R2930 GNDA.n1542 GNDA.n1527 76.3222
R2931 GNDA.n1546 GNDA.n1528 76.3222
R2932 GNDA.n1552 GNDA.n1551 76.3222
R2933 GNDA.n1709 GNDA.n363 76.3222
R2934 GNDA.n1707 GNDA.n1706 76.3222
R2935 GNDA.n1702 GNDA.n372 76.3222
R2936 GNDA.n1700 GNDA.n1699 76.3222
R2937 GNDA.n1695 GNDA.n381 76.3222
R2938 GNDA.n1693 GNDA.n1692 76.3222
R2939 GNDA.n1726 GNDA.n1725 76.3222
R2940 GNDA.n336 GNDA.n333 76.3222
R2941 GNDA.n343 GNDA.n330 76.3222
R2942 GNDA.n344 GNDA.n327 76.3222
R2943 GNDA.n355 GNDA.n354 76.3222
R2944 GNDA.n1715 GNDA.n1714 76.3222
R2945 GNDA.n1727 GNDA.n1726 76.3222
R2946 GNDA.n333 GNDA.n252 76.3222
R2947 GNDA.n337 GNDA.n330 76.3222
R2948 GNDA.n345 GNDA.n344 76.3222
R2949 GNDA.n354 GNDA.n353 76.3222
R2950 GNDA.n1716 GNDA.n1715 76.3222
R2951 GNDA.n1552 GNDA.n382 76.3222
R2952 GNDA.n1529 GNDA.n1528 76.3222
R2953 GNDA.n1545 GNDA.n1527 76.3222
R2954 GNDA.n1541 GNDA.n1526 76.3222
R2955 GNDA.n1537 GNDA.n1525 76.3222
R2956 GNDA.n1533 GNDA.n1524 76.3222
R2957 GNDA.n2076 GNDA.n2075 76.3222
R2958 GNDA.n18 GNDA.n7 76.3222
R2959 GNDA.n17 GNDA.n6 76.3222
R2960 GNDA.n148 GNDA.n1 76.3222
R2961 GNDA.n152 GNDA.n151 76.3222
R2962 GNDA.n144 GNDA.n143 76.3222
R2963 GNDA.n141 GNDA.n140 76.3222
R2964 GNDA.n10 GNDA.n5 76.3222
R2965 GNDA.n2202 GNDA.n2201 76.3222
R2966 GNDA.n147 GNDA.n3 76.3222
R2967 GNDA.n156 GNDA.n155 76.3222
R2968 GNDA.n146 GNDA.n138 76.3222
R2969 GNDA.n163 GNDA.n162 76.3222
R2970 GNDA.n1414 GNDA.n11 76.3222
R2971 GNDA.n1413 GNDA.n1412 76.3222
R2972 GNDA.n1421 GNDA.n1420 76.3222
R2973 GNDA.n1411 GNDA.n1409 76.3222
R2974 GNDA.n1428 GNDA.n1427 76.3222
R2975 GNDA.n1431 GNDA.n1430 76.3222
R2976 GNDA.n691 GNDA.n690 76.3222
R2977 GNDA.n763 GNDA.n762 76.3222
R2978 GNDA.n764 GNDA.n683 76.3222
R2979 GNDA.n778 GNDA.n777 76.3222
R2980 GNDA.n779 GNDA.n675 76.3222
R2981 GNDA.n794 GNDA.n793 76.3222
R2982 GNDA.n661 GNDA.n635 76.3222
R2983 GNDA.n659 GNDA.n640 76.3222
R2984 GNDA.n652 GNDA.n639 76.3222
R2985 GNDA.n648 GNDA.n638 76.3222
R2986 GNDA.n644 GNDA.n637 76.3222
R2987 GNDA.n636 GNDA.n387 76.3222
R2988 GNDA.n1149 GNDA.n392 76.3222
R2989 GNDA.n1147 GNDA.n397 76.3222
R2990 GNDA.n431 GNDA.n396 76.3222
R2991 GNDA.n439 GNDA.n395 76.3222
R2992 GNDA.n1086 GNDA.n394 76.3222
R2993 GNDA.n1083 GNDA.n393 76.3222
R2994 GNDA.n1402 GNDA.n1401 76.3222
R2995 GNDA.n1390 GNDA.n1360 76.3222
R2996 GNDA.n1389 GNDA.n1388 76.3222
R2997 GNDA.n1381 GNDA.n1380 76.3222
R2998 GNDA.n1378 GNDA.n1377 76.3222
R2999 GNDA.n1369 GNDA.n1368 76.3222
R3000 GNDA.n384 GNDA.n383 76.3222
R3001 GNDA.n378 GNDA.n377 76.3222
R3002 GNDA.n375 GNDA.n374 76.3222
R3003 GNDA.n369 GNDA.n368 76.3222
R3004 GNDA.n366 GNDA.n365 76.3222
R3005 GNDA.n360 GNDA.n359 76.3222
R3006 GNDA.n1258 GNDA.n1257 76.3222
R3007 GNDA.n1247 GNDA.n1218 76.3222
R3008 GNDA.n1246 GNDA.n1245 76.3222
R3009 GNDA.n1238 GNDA.n1237 76.3222
R3010 GNDA.n1235 GNDA.n1234 76.3222
R3011 GNDA.n1226 GNDA.n1225 76.3222
R3012 GNDA.n1397 GNDA.n1396 76.3222
R3013 GNDA.n1395 GNDA.n1394 76.3222
R3014 GNDA.n1386 GNDA.n1362 76.3222
R3015 GNDA.n1384 GNDA.n1383 76.3222
R3016 GNDA.n1375 GNDA.n1374 76.3222
R3017 GNDA.n1372 GNDA.n205 76.3222
R3018 GNDA.n1694 GNDA.n1693 76.3222
R3019 GNDA.n381 GNDA.n373 76.3222
R3020 GNDA.n1701 GNDA.n1700 76.3222
R3021 GNDA.n372 GNDA.n364 76.3222
R3022 GNDA.n1708 GNDA.n1707 76.3222
R3023 GNDA.n363 GNDA.n356 76.3222
R3024 GNDA.n1253 GNDA.n1216 76.3222
R3025 GNDA.n1252 GNDA.n1251 76.3222
R3026 GNDA.n1243 GNDA.n1220 76.3222
R3027 GNDA.n1241 GNDA.n1240 76.3222
R3028 GNDA.n1232 GNDA.n1231 76.3222
R3029 GNDA.n1229 GNDA.n1154 76.3222
R3030 GNDA.n1337 GNDA.n1336 76.3222
R3031 GNDA.n1325 GNDA.n1324 76.3222
R3032 GNDA.n1593 GNDA.n1188 76.3222
R3033 GNDA.n1990 GNDA.t97 75.0005
R3034 GNDA.n1990 GNDA.t3 75.0005
R3035 GNDA.n1960 GNDA.t98 75.0005
R3036 GNDA.n1981 GNDA.n1980 75.0005
R3037 GNDA.n1980 GNDA.n1979 75.0005
R3038 GNDA.n2017 GNDA.t64 75.0005
R3039 GNDA.t38 GNDA.n2015 75.0005
R3040 GNDA.n2015 GNDA.t62 75.0005
R3041 GNDA.n2084 GNDA.n2083 74.5978
R3042 GNDA.n2085 GNDA.n2084 74.5978
R3043 GNDA.n1923 GNDA.n1922 74.5978
R3044 GNDA.n1922 GNDA.n167 74.5978
R3045 GNDA.n1678 GNDA.n1677 74.5978
R3046 GNDA.n1677 GNDA.n1159 74.5978
R3047 GNDA.n501 GNDA.n471 74.5978
R3048 GNDA.n502 GNDA.n501 74.5978
R3049 GNDA.n787 GNDA.n786 74.5978
R3050 GNDA.n788 GNDA.n787 74.5978
R3051 GNDA.n1005 GNDA.n1004 74.5978
R3052 GNDA.n1004 GNDA.n892 74.5978
R3053 GNDA.n1091 GNDA.n1090 74.5978
R3054 GNDA.n1092 GNDA.n1091 74.5978
R3055 GNDA.n1828 GNDA.n1827 74.5978
R3056 GNDA.n1827 GNDA.n209 74.5978
R3057 GNDA.n1720 GNDA.n1719 74.5978
R3058 GNDA.n1720 GNDA.n273 74.5978
R3059 GNDA.n2117 GNDA.n2116 69.3109
R3060 GNDA.n2116 GNDA.n2115 69.3109
R3061 GNDA.n1875 GNDA.n175 69.3109
R3062 GNDA.n1872 GNDA.n175 69.3109
R3063 GNDA.n1633 GNDA.n1167 69.3109
R3064 GNDA.n1630 GNDA.n1167 69.3109
R3065 GNDA.n534 GNDA.n533 69.3109
R3066 GNDA.n533 GNDA.n532 69.3109
R3067 GNDA.n739 GNDA.n738 69.3109
R3068 GNDA.n738 GNDA.n737 69.3109
R3069 GNDA.n960 GNDA.n900 69.3109
R3070 GNDA.n957 GNDA.n900 69.3109
R3071 GNDA.n1124 GNDA.n1123 69.3109
R3072 GNDA.n1123 GNDA.n1122 69.3109
R3073 GNDA.n1779 GNDA.n217 69.3109
R3074 GNDA.n1776 GNDA.n217 69.3109
R3075 GNDA.n291 GNDA.n263 69.3109
R3076 GNDA.n294 GNDA.n263 69.3109
R3077 GNDA.n2096 GNDA.t91 65.8183
R3078 GNDA.n2093 GNDA.t91 65.8183
R3079 GNDA.n2087 GNDA.t91 65.8183
R3080 GNDA.n2102 GNDA.t91 65.8183
R3081 GNDA.n2041 GNDA.t91 65.8183
R3082 GNDA.n2109 GNDA.t91 65.8183
R3083 GNDA.n2038 GNDA.t91 65.8183
R3084 GNDA.n2034 GNDA.t91 65.8183
R3085 GNDA.n2122 GNDA.t91 65.8183
R3086 GNDA.n2128 GNDA.t91 65.8183
R3087 GNDA.n53 GNDA.t91 65.8183
R3088 GNDA.t73 GNDA.n174 65.8183
R3089 GNDA.t73 GNDA.n172 65.8183
R3090 GNDA.t73 GNDA.n170 65.8183
R3091 GNDA.t73 GNDA.n177 65.8183
R3092 GNDA.t73 GNDA.n178 65.8183
R3093 GNDA.t73 GNDA.n179 65.8183
R3094 GNDA.t73 GNDA.n180 65.8183
R3095 GNDA.t73 GNDA.n173 65.8183
R3096 GNDA.t73 GNDA.n171 65.8183
R3097 GNDA.t73 GNDA.n169 65.8183
R3098 GNDA.t73 GNDA.n168 65.8183
R3099 GNDA.t92 GNDA.n1166 65.8183
R3100 GNDA.t92 GNDA.n1164 65.8183
R3101 GNDA.t92 GNDA.n1162 65.8183
R3102 GNDA.t92 GNDA.n1169 65.8183
R3103 GNDA.t92 GNDA.n1170 65.8183
R3104 GNDA.t92 GNDA.n1171 65.8183
R3105 GNDA.t92 GNDA.n1172 65.8183
R3106 GNDA.t92 GNDA.n1165 65.8183
R3107 GNDA.t92 GNDA.n1163 65.8183
R3108 GNDA.t92 GNDA.n1161 65.8183
R3109 GNDA.t92 GNDA.n1160 65.8183
R3110 GNDA.n513 GNDA.t75 65.8183
R3111 GNDA.n510 GNDA.t75 65.8183
R3112 GNDA.n504 GNDA.t75 65.8183
R3113 GNDA.n519 GNDA.t75 65.8183
R3114 GNDA.n495 GNDA.t75 65.8183
R3115 GNDA.n526 GNDA.t75 65.8183
R3116 GNDA.n492 GNDA.t75 65.8183
R3117 GNDA.n488 GNDA.t75 65.8183
R3118 GNDA.n539 GNDA.t75 65.8183
R3119 GNDA.n545 GNDA.t75 65.8183
R3120 GNDA.n481 GNDA.t75 65.8183
R3121 GNDA.n718 GNDA.t67 65.8183
R3122 GNDA.n715 GNDA.t67 65.8183
R3123 GNDA.n709 GNDA.t67 65.8183
R3124 GNDA.n724 GNDA.t67 65.8183
R3125 GNDA.n704 GNDA.t67 65.8183
R3126 GNDA.n731 GNDA.t67 65.8183
R3127 GNDA.n701 GNDA.t67 65.8183
R3128 GNDA.n697 GNDA.t67 65.8183
R3129 GNDA.n744 GNDA.t67 65.8183
R3130 GNDA.n750 GNDA.t67 65.8183
R3131 GNDA.n693 GNDA.t67 65.8183
R3132 GNDA.n756 GNDA.t67 65.8183
R3133 GNDA.n769 GNDA.t67 65.8183
R3134 GNDA.n771 GNDA.t67 65.8183
R3135 GNDA.n784 GNDA.t67 65.8183
R3136 GNDA.t69 GNDA.n899 65.8183
R3137 GNDA.t69 GNDA.n897 65.8183
R3138 GNDA.t69 GNDA.n895 65.8183
R3139 GNDA.t69 GNDA.n902 65.8183
R3140 GNDA.t69 GNDA.n903 65.8183
R3141 GNDA.t69 GNDA.n904 65.8183
R3142 GNDA.t69 GNDA.n905 65.8183
R3143 GNDA.t69 GNDA.n898 65.8183
R3144 GNDA.t69 GNDA.n896 65.8183
R3145 GNDA.t69 GNDA.n894 65.8183
R3146 GNDA.t69 GNDA.n893 65.8183
R3147 GNDA.n1103 GNDA.t93 65.8183
R3148 GNDA.n1100 GNDA.t93 65.8183
R3149 GNDA.n1094 GNDA.t93 65.8183
R3150 GNDA.n1109 GNDA.t93 65.8183
R3151 GNDA.n412 GNDA.t93 65.8183
R3152 GNDA.n1116 GNDA.t93 65.8183
R3153 GNDA.n409 GNDA.t93 65.8183
R3154 GNDA.n405 GNDA.t93 65.8183
R3155 GNDA.n1129 GNDA.t93 65.8183
R3156 GNDA.n1135 GNDA.t93 65.8183
R3157 GNDA.n402 GNDA.t93 65.8183
R3158 GNDA.n1142 GNDA.t93 65.8183
R3159 GNDA.n424 GNDA.t93 65.8183
R3160 GNDA.n435 GNDA.t93 65.8183
R3161 GNDA.n422 GNDA.t93 65.8183
R3162 GNDA.t69 GNDA.n907 65.8183
R3163 GNDA.t69 GNDA.n908 65.8183
R3164 GNDA.t69 GNDA.n909 65.8183
R3165 GNDA.t69 GNDA.n1003 65.8183
R3166 GNDA.n551 GNDA.t75 65.8183
R3167 GNDA.n564 GNDA.t75 65.8183
R3168 GNDA.n566 GNDA.t75 65.8183
R3169 GNDA.n577 GNDA.t75 65.8183
R3170 GNDA.t92 GNDA.n1174 65.8183
R3171 GNDA.t92 GNDA.n1175 65.8183
R3172 GNDA.t92 GNDA.n1176 65.8183
R3173 GNDA.t92 GNDA.n1676 65.8183
R3174 GNDA.t71 GNDA.n216 65.8183
R3175 GNDA.t71 GNDA.n214 65.8183
R3176 GNDA.t71 GNDA.n212 65.8183
R3177 GNDA.t71 GNDA.n219 65.8183
R3178 GNDA.t71 GNDA.n220 65.8183
R3179 GNDA.t71 GNDA.n221 65.8183
R3180 GNDA.t71 GNDA.n222 65.8183
R3181 GNDA.t71 GNDA.n215 65.8183
R3182 GNDA.t71 GNDA.n213 65.8183
R3183 GNDA.t71 GNDA.n211 65.8183
R3184 GNDA.t71 GNDA.n210 65.8183
R3185 GNDA.t71 GNDA.n224 65.8183
R3186 GNDA.t71 GNDA.n225 65.8183
R3187 GNDA.t71 GNDA.n226 65.8183
R3188 GNDA.t71 GNDA.n1826 65.8183
R3189 GNDA.t74 GNDA.n262 65.8183
R3190 GNDA.t74 GNDA.n260 65.8183
R3191 GNDA.t74 GNDA.n258 65.8183
R3192 GNDA.t74 GNDA.n265 65.8183
R3193 GNDA.t74 GNDA.n266 65.8183
R3194 GNDA.t74 GNDA.n267 65.8183
R3195 GNDA.t74 GNDA.n268 65.8183
R3196 GNDA.t74 GNDA.n261 65.8183
R3197 GNDA.t74 GNDA.n259 65.8183
R3198 GNDA.t74 GNDA.n257 65.8183
R3199 GNDA.t74 GNDA.n256 65.8183
R3200 GNDA.n1721 GNDA.t74 65.8183
R3201 GNDA.t74 GNDA.n270 65.8183
R3202 GNDA.t74 GNDA.n271 65.8183
R3203 GNDA.t74 GNDA.n272 65.8183
R3204 GNDA.t73 GNDA.n182 65.8183
R3205 GNDA.t73 GNDA.n183 65.8183
R3206 GNDA.t73 GNDA.n184 65.8183
R3207 GNDA.t73 GNDA.n1921 65.8183
R3208 GNDA.n2134 GNDA.t91 65.8183
R3209 GNDA.n2147 GNDA.t91 65.8183
R3210 GNDA.n2150 GNDA.t91 65.8183
R3211 GNDA.n2048 GNDA.t91 65.8183
R3212 GNDA.n1961 GNDA.t4 62.5005
R3213 GNDA.t39 GNDA.n2016 62.5005
R3214 GNDA.n2190 GNDA.t70 60.9488
R3215 GNDA.n1688 GNDA.t68 60.9488
R3216 GNDA.n1507 GNDA.n1473 59.6972
R3217 GNDA.n1588 GNDA.n1193 59.6972
R3218 GNDA.n2116 GNDA.t91 57.8461
R3219 GNDA.t73 GNDA.n175 57.8461
R3220 GNDA.t92 GNDA.n1167 57.8461
R3221 GNDA.n533 GNDA.t75 57.8461
R3222 GNDA.n738 GNDA.t67 57.8461
R3223 GNDA.t69 GNDA.n900 57.8461
R3224 GNDA.n1123 GNDA.t93 57.8461
R3225 GNDA.t71 GNDA.n217 57.8461
R3226 GNDA.t74 GNDA.n263 57.8461
R3227 GNDA.n787 GNDA.t67 55.2026
R3228 GNDA.n1091 GNDA.t93 55.2026
R3229 GNDA.n1004 GNDA.t69 55.2026
R3230 GNDA.n501 GNDA.t75 55.2026
R3231 GNDA.n1677 GNDA.t92 55.2026
R3232 GNDA.n1827 GNDA.t71 55.2026
R3233 GNDA.t74 GNDA.n1720 55.2026
R3234 GNDA.n1922 GNDA.t73 55.2026
R3235 GNDA.n2084 GNDA.t91 55.2026
R3236 GNDA.n2135 GNDA.n2134 53.3664
R3237 GNDA.n2147 GNDA.n2146 53.3664
R3238 GNDA.n2150 GNDA.n2149 53.3664
R3239 GNDA.n2048 GNDA.n44 53.3664
R3240 GNDA.n2133 GNDA.n53 53.3664
R3241 GNDA.n2129 GNDA.n2128 53.3664
R3242 GNDA.n2122 GNDA.n2033 53.3664
R3243 GNDA.n2121 GNDA.n2034 53.3664
R3244 GNDA.n2111 GNDA.n2038 53.3664
R3245 GNDA.n2109 GNDA.n2108 53.3664
R3246 GNDA.n2104 GNDA.n2041 53.3664
R3247 GNDA.n2102 GNDA.n2101 53.3664
R3248 GNDA.n2088 GNDA.n2087 53.3664
R3249 GNDA.n2093 GNDA.n2092 53.3664
R3250 GNDA.n2096 GNDA.n2095 53.3664
R3251 GNDA.n2097 GNDA.n2096 53.3664
R3252 GNDA.n2094 GNDA.n2093 53.3664
R3253 GNDA.n2087 GNDA.n2045 53.3664
R3254 GNDA.n2103 GNDA.n2102 53.3664
R3255 GNDA.n2041 GNDA.n2039 53.3664
R3256 GNDA.n2110 GNDA.n2109 53.3664
R3257 GNDA.n2038 GNDA.n2036 53.3664
R3258 GNDA.n2118 GNDA.n2034 53.3664
R3259 GNDA.n2123 GNDA.n2122 53.3664
R3260 GNDA.n2128 GNDA.n2127 53.3664
R3261 GNDA.n2130 GNDA.n53 53.3664
R3262 GNDA.n1892 GNDA.n182 53.3664
R3263 GNDA.n1895 GNDA.n183 53.3664
R3264 GNDA.n1908 GNDA.n184 53.3664
R3265 GNDA.n1921 GNDA.n1920 53.3664
R3266 GNDA.n1891 GNDA.n168 53.3664
R3267 GNDA.n1887 GNDA.n169 53.3664
R3268 GNDA.n1883 GNDA.n171 53.3664
R3269 GNDA.n1879 GNDA.n173 53.3664
R3270 GNDA.n1868 GNDA.n180 53.3664
R3271 GNDA.n1864 GNDA.n179 53.3664
R3272 GNDA.n1860 GNDA.n178 53.3664
R3273 GNDA.n1856 GNDA.n177 53.3664
R3274 GNDA.n1843 GNDA.n170 53.3664
R3275 GNDA.n1847 GNDA.n172 53.3664
R3276 GNDA.n1851 GNDA.n174 53.3664
R3277 GNDA.n1853 GNDA.n174 53.3664
R3278 GNDA.n1850 GNDA.n172 53.3664
R3279 GNDA.n1846 GNDA.n170 53.3664
R3280 GNDA.n1859 GNDA.n177 53.3664
R3281 GNDA.n1863 GNDA.n178 53.3664
R3282 GNDA.n1867 GNDA.n179 53.3664
R3283 GNDA.n1871 GNDA.n180 53.3664
R3284 GNDA.n1876 GNDA.n173 53.3664
R3285 GNDA.n1880 GNDA.n171 53.3664
R3286 GNDA.n1884 GNDA.n169 53.3664
R3287 GNDA.n1888 GNDA.n168 53.3664
R3288 GNDA.n1650 GNDA.n1174 53.3664
R3289 GNDA.n1652 GNDA.n1175 53.3664
R3290 GNDA.n1664 GNDA.n1176 53.3664
R3291 GNDA.n1676 GNDA.n1675 53.3664
R3292 GNDA.n1649 GNDA.n1160 53.3664
R3293 GNDA.n1645 GNDA.n1161 53.3664
R3294 GNDA.n1641 GNDA.n1163 53.3664
R3295 GNDA.n1637 GNDA.n1165 53.3664
R3296 GNDA.n1626 GNDA.n1172 53.3664
R3297 GNDA.n1622 GNDA.n1171 53.3664
R3298 GNDA.n1618 GNDA.n1170 53.3664
R3299 GNDA.n1614 GNDA.n1169 53.3664
R3300 GNDA.n1601 GNDA.n1162 53.3664
R3301 GNDA.n1605 GNDA.n1164 53.3664
R3302 GNDA.n1609 GNDA.n1166 53.3664
R3303 GNDA.n1611 GNDA.n1166 53.3664
R3304 GNDA.n1608 GNDA.n1164 53.3664
R3305 GNDA.n1604 GNDA.n1162 53.3664
R3306 GNDA.n1617 GNDA.n1169 53.3664
R3307 GNDA.n1621 GNDA.n1170 53.3664
R3308 GNDA.n1625 GNDA.n1171 53.3664
R3309 GNDA.n1629 GNDA.n1172 53.3664
R3310 GNDA.n1634 GNDA.n1165 53.3664
R3311 GNDA.n1638 GNDA.n1163 53.3664
R3312 GNDA.n1642 GNDA.n1161 53.3664
R3313 GNDA.n1646 GNDA.n1160 53.3664
R3314 GNDA.n552 GNDA.n551 53.3664
R3315 GNDA.n564 GNDA.n563 53.3664
R3316 GNDA.n567 GNDA.n566 53.3664
R3317 GNDA.n577 GNDA.n576 53.3664
R3318 GNDA.n550 GNDA.n481 53.3664
R3319 GNDA.n546 GNDA.n545 53.3664
R3320 GNDA.n539 GNDA.n487 53.3664
R3321 GNDA.n538 GNDA.n488 53.3664
R3322 GNDA.n528 GNDA.n492 53.3664
R3323 GNDA.n526 GNDA.n525 53.3664
R3324 GNDA.n521 GNDA.n495 53.3664
R3325 GNDA.n519 GNDA.n518 53.3664
R3326 GNDA.n505 GNDA.n504 53.3664
R3327 GNDA.n510 GNDA.n509 53.3664
R3328 GNDA.n513 GNDA.n512 53.3664
R3329 GNDA.n514 GNDA.n513 53.3664
R3330 GNDA.n511 GNDA.n510 53.3664
R3331 GNDA.n504 GNDA.n499 53.3664
R3332 GNDA.n520 GNDA.n519 53.3664
R3333 GNDA.n495 GNDA.n493 53.3664
R3334 GNDA.n527 GNDA.n526 53.3664
R3335 GNDA.n492 GNDA.n490 53.3664
R3336 GNDA.n535 GNDA.n488 53.3664
R3337 GNDA.n540 GNDA.n539 53.3664
R3338 GNDA.n545 GNDA.n544 53.3664
R3339 GNDA.n547 GNDA.n481 53.3664
R3340 GNDA.n757 GNDA.n756 53.3664
R3341 GNDA.n769 GNDA.n768 53.3664
R3342 GNDA.n772 GNDA.n771 53.3664
R3343 GNDA.n784 GNDA.n783 53.3664
R3344 GNDA.n755 GNDA.n693 53.3664
R3345 GNDA.n751 GNDA.n750 53.3664
R3346 GNDA.n744 GNDA.n696 53.3664
R3347 GNDA.n743 GNDA.n697 53.3664
R3348 GNDA.n733 GNDA.n701 53.3664
R3349 GNDA.n731 GNDA.n730 53.3664
R3350 GNDA.n726 GNDA.n704 53.3664
R3351 GNDA.n724 GNDA.n723 53.3664
R3352 GNDA.n710 GNDA.n709 53.3664
R3353 GNDA.n715 GNDA.n714 53.3664
R3354 GNDA.n718 GNDA.n717 53.3664
R3355 GNDA.n719 GNDA.n718 53.3664
R3356 GNDA.n716 GNDA.n715 53.3664
R3357 GNDA.n709 GNDA.n708 53.3664
R3358 GNDA.n725 GNDA.n724 53.3664
R3359 GNDA.n704 GNDA.n702 53.3664
R3360 GNDA.n732 GNDA.n731 53.3664
R3361 GNDA.n701 GNDA.n699 53.3664
R3362 GNDA.n740 GNDA.n697 53.3664
R3363 GNDA.n745 GNDA.n744 53.3664
R3364 GNDA.n750 GNDA.n749 53.3664
R3365 GNDA.n752 GNDA.n693 53.3664
R3366 GNDA.n756 GNDA.n686 53.3664
R3367 GNDA.n770 GNDA.n769 53.3664
R3368 GNDA.n771 GNDA.n681 53.3664
R3369 GNDA.n785 GNDA.n784 53.3664
R3370 GNDA.n977 GNDA.n907 53.3664
R3371 GNDA.n979 GNDA.n908 53.3664
R3372 GNDA.n991 GNDA.n909 53.3664
R3373 GNDA.n1003 GNDA.n1002 53.3664
R3374 GNDA.n976 GNDA.n893 53.3664
R3375 GNDA.n972 GNDA.n894 53.3664
R3376 GNDA.n968 GNDA.n896 53.3664
R3377 GNDA.n964 GNDA.n898 53.3664
R3378 GNDA.n953 GNDA.n905 53.3664
R3379 GNDA.n949 GNDA.n904 53.3664
R3380 GNDA.n945 GNDA.n903 53.3664
R3381 GNDA.n941 GNDA.n902 53.3664
R3382 GNDA.n928 GNDA.n895 53.3664
R3383 GNDA.n932 GNDA.n897 53.3664
R3384 GNDA.n936 GNDA.n899 53.3664
R3385 GNDA.n938 GNDA.n899 53.3664
R3386 GNDA.n935 GNDA.n897 53.3664
R3387 GNDA.n931 GNDA.n895 53.3664
R3388 GNDA.n944 GNDA.n902 53.3664
R3389 GNDA.n948 GNDA.n903 53.3664
R3390 GNDA.n952 GNDA.n904 53.3664
R3391 GNDA.n956 GNDA.n905 53.3664
R3392 GNDA.n961 GNDA.n898 53.3664
R3393 GNDA.n965 GNDA.n896 53.3664
R3394 GNDA.n969 GNDA.n894 53.3664
R3395 GNDA.n973 GNDA.n893 53.3664
R3396 GNDA.n1142 GNDA.n1141 53.3664
R3397 GNDA.n424 GNDA.n401 53.3664
R3398 GNDA.n435 GNDA.n434 53.3664
R3399 GNDA.n423 GNDA.n422 53.3664
R3400 GNDA.n1140 GNDA.n402 53.3664
R3401 GNDA.n1136 GNDA.n1135 53.3664
R3402 GNDA.n1129 GNDA.n404 53.3664
R3403 GNDA.n1128 GNDA.n405 53.3664
R3404 GNDA.n1118 GNDA.n409 53.3664
R3405 GNDA.n1116 GNDA.n1115 53.3664
R3406 GNDA.n1111 GNDA.n412 53.3664
R3407 GNDA.n1109 GNDA.n1108 53.3664
R3408 GNDA.n1095 GNDA.n1094 53.3664
R3409 GNDA.n1100 GNDA.n1099 53.3664
R3410 GNDA.n1103 GNDA.n1102 53.3664
R3411 GNDA.n1104 GNDA.n1103 53.3664
R3412 GNDA.n1101 GNDA.n1100 53.3664
R3413 GNDA.n1094 GNDA.n416 53.3664
R3414 GNDA.n1110 GNDA.n1109 53.3664
R3415 GNDA.n412 GNDA.n410 53.3664
R3416 GNDA.n1117 GNDA.n1116 53.3664
R3417 GNDA.n409 GNDA.n407 53.3664
R3418 GNDA.n1125 GNDA.n405 53.3664
R3419 GNDA.n1130 GNDA.n1129 53.3664
R3420 GNDA.n1135 GNDA.n1134 53.3664
R3421 GNDA.n1137 GNDA.n402 53.3664
R3422 GNDA.n1143 GNDA.n1142 53.3664
R3423 GNDA.n425 GNDA.n424 53.3664
R3424 GNDA.n436 GNDA.n435 53.3664
R3425 GNDA.n422 GNDA.n419 53.3664
R3426 GNDA.n980 GNDA.n907 53.3664
R3427 GNDA.n990 GNDA.n908 53.3664
R3428 GNDA.n910 GNDA.n909 53.3664
R3429 GNDA.n1003 GNDA.n891 53.3664
R3430 GNDA.n551 GNDA.n477 53.3664
R3431 GNDA.n565 GNDA.n564 53.3664
R3432 GNDA.n566 GNDA.n472 53.3664
R3433 GNDA.n578 GNDA.n577 53.3664
R3434 GNDA.n1653 GNDA.n1174 53.3664
R3435 GNDA.n1663 GNDA.n1175 53.3664
R3436 GNDA.n1177 GNDA.n1176 53.3664
R3437 GNDA.n1676 GNDA.n1158 53.3664
R3438 GNDA.n1796 GNDA.n224 53.3664
R3439 GNDA.n1799 GNDA.n225 53.3664
R3440 GNDA.n1813 GNDA.n226 53.3664
R3441 GNDA.n1826 GNDA.n1825 53.3664
R3442 GNDA.n1795 GNDA.n210 53.3664
R3443 GNDA.n1791 GNDA.n211 53.3664
R3444 GNDA.n1787 GNDA.n213 53.3664
R3445 GNDA.n1783 GNDA.n215 53.3664
R3446 GNDA.n1772 GNDA.n222 53.3664
R3447 GNDA.n1768 GNDA.n221 53.3664
R3448 GNDA.n1764 GNDA.n220 53.3664
R3449 GNDA.n1760 GNDA.n219 53.3664
R3450 GNDA.n1747 GNDA.n212 53.3664
R3451 GNDA.n1751 GNDA.n214 53.3664
R3452 GNDA.n1755 GNDA.n216 53.3664
R3453 GNDA.n1757 GNDA.n216 53.3664
R3454 GNDA.n1754 GNDA.n214 53.3664
R3455 GNDA.n1750 GNDA.n212 53.3664
R3456 GNDA.n1763 GNDA.n219 53.3664
R3457 GNDA.n1767 GNDA.n220 53.3664
R3458 GNDA.n1771 GNDA.n221 53.3664
R3459 GNDA.n1775 GNDA.n222 53.3664
R3460 GNDA.n1780 GNDA.n215 53.3664
R3461 GNDA.n1784 GNDA.n213 53.3664
R3462 GNDA.n1788 GNDA.n211 53.3664
R3463 GNDA.n1792 GNDA.n210 53.3664
R3464 GNDA.n1800 GNDA.n224 53.3664
R3465 GNDA.n1812 GNDA.n225 53.3664
R3466 GNDA.n227 GNDA.n226 53.3664
R3467 GNDA.n1826 GNDA.n208 53.3664
R3468 GNDA.n1722 GNDA.n1721 53.3664
R3469 GNDA.n331 GNDA.n270 53.3664
R3470 GNDA.n339 GNDA.n271 53.3664
R3471 GNDA.n349 GNDA.n272 53.3664
R3472 GNDA.n256 GNDA.n254 53.3664
R3473 GNDA.n279 GNDA.n257 53.3664
R3474 GNDA.n283 GNDA.n259 53.3664
R3475 GNDA.n287 GNDA.n261 53.3664
R3476 GNDA.n298 GNDA.n268 53.3664
R3477 GNDA.n302 GNDA.n267 53.3664
R3478 GNDA.n306 GNDA.n266 53.3664
R3479 GNDA.n309 GNDA.n265 53.3664
R3480 GNDA.n322 GNDA.n258 53.3664
R3481 GNDA.n319 GNDA.n260 53.3664
R3482 GNDA.n315 GNDA.n262 53.3664
R3483 GNDA.n312 GNDA.n262 53.3664
R3484 GNDA.n316 GNDA.n260 53.3664
R3485 GNDA.n320 GNDA.n258 53.3664
R3486 GNDA.n307 GNDA.n265 53.3664
R3487 GNDA.n303 GNDA.n266 53.3664
R3488 GNDA.n299 GNDA.n267 53.3664
R3489 GNDA.n295 GNDA.n268 53.3664
R3490 GNDA.n290 GNDA.n261 53.3664
R3491 GNDA.n286 GNDA.n259 53.3664
R3492 GNDA.n282 GNDA.n257 53.3664
R3493 GNDA.n278 GNDA.n256 53.3664
R3494 GNDA.n1721 GNDA.n255 53.3664
R3495 GNDA.n340 GNDA.n270 53.3664
R3496 GNDA.n348 GNDA.n271 53.3664
R3497 GNDA.n274 GNDA.n272 53.3664
R3498 GNDA.n1896 GNDA.n182 53.3664
R3499 GNDA.n1907 GNDA.n183 53.3664
R3500 GNDA.n185 GNDA.n184 53.3664
R3501 GNDA.n1921 GNDA.n166 53.3664
R3502 GNDA.n2134 GNDA.n47 53.3664
R3503 GNDA.n2148 GNDA.n2147 53.3664
R3504 GNDA.n2151 GNDA.n2150 53.3664
R3505 GNDA.n2049 GNDA.n2048 53.3664
R3506 GNDA.t16 GNDA.n1486 51.0719
R3507 GNDA.n1946 GNDA.n125 50.5752
R3508 GNDA.n92 GNDA.t103 50.0005
R3509 GNDA.t53 GNDA.t2 50.0005
R3510 GNDA.t4 GNDA.t49 50.0005
R3511 GNDA.t9 GNDA.t39 50.0005
R3512 GNDA.t26 GNDA.t21 50.0005
R3513 GNDA.n2002 GNDA.t35 50.0005
R3514 GNDA.n1564 GNDA.n1315 45.6509
R3515 GNDA.n1808 GNDA.n1806 43.0993
R3516 GNDA.n1486 GNDA.n1485 39.2862
R3517 GNDA.t27 GNDA.t89 37.5005
R3518 GNDA.n1981 GNDA.t105 37.5005
R3519 GNDA.n1979 GNDA.t33 37.5005
R3520 GNDA.t95 GNDA.t65 37.5005
R3521 GNDA.t32 GNDA.n1495 35.3576
R3522 GNDA.n1193 GNDA.t59 31.6047
R3523 GNDA.n1504 GNDA.n1503 28.1318
R3524 GNDA.n2020 GNDA.n2019 27.8193
R3525 GNDA.n1963 GNDA.n1956 27.8193
R3526 GNDA.n2100 GNDA.n2099 27.5561
R3527 GNDA.n1857 GNDA.n1855 27.5561
R3528 GNDA.n1615 GNDA.n1613 27.5561
R3529 GNDA.n517 GNDA.n516 27.5561
R3530 GNDA.n722 GNDA.n721 27.5561
R3531 GNDA.n942 GNDA.n940 27.5561
R3532 GNDA.n1107 GNDA.n1106 27.5561
R3533 GNDA.n1761 GNDA.n1759 27.5561
R3534 GNDA.n311 GNDA.n310 27.5561
R3535 GNDA.n2190 GNDA.n19 26.9584
R3536 GNDA.n1688 GNDA.n202 26.9584
R3537 GNDA.t23 GNDA.t57 25.0005
R3538 GNDA.t97 GNDA.t83 25.0005
R3539 GNDA.t49 GNDA.n1960 25.0005
R3540 GNDA.n2017 GNDA.t9 25.0005
R3541 GNDA.t86 GNDA.t62 25.0005
R3542 GNDA.t47 GNDA.t52 25.0005
R3543 GNDA.n2001 GNDA.t28 25.0005
R3544 GNDA.n1508 GNDA.n1320 24.5815
R3545 GNDA.t59 GNDA.t17 24.5815
R3546 GNDA.n113 GNDA.t104 24.0005
R3547 GNDA.n113 GNDA.t42 24.0005
R3548 GNDA.n111 GNDA.t25 24.0005
R3549 GNDA.n111 GNDA.t61 24.0005
R3550 GNDA.n109 GNDA.t58 24.0005
R3551 GNDA.n109 GNDA.t54 24.0005
R3552 GNDA.n107 GNDA.t1 24.0005
R3553 GNDA.n107 GNDA.t44 24.0005
R3554 GNDA.n105 GNDA.t56 24.0005
R3555 GNDA.n105 GNDA.t106 24.0005
R3556 GNDA.n103 GNDA.t34 24.0005
R3557 GNDA.n103 GNDA.t46 24.0005
R3558 GNDA.n101 GNDA.t13 24.0005
R3559 GNDA.n101 GNDA.t11 24.0005
R3560 GNDA.n99 GNDA.t22 24.0005
R3561 GNDA.n99 GNDA.t48 24.0005
R3562 GNDA.n97 GNDA.t102 24.0005
R3563 GNDA.n97 GNDA.t100 24.0005
R3564 GNDA.n96 GNDA.t29 24.0005
R3565 GNDA.n96 GNDA.t36 24.0005
R3566 GNDA.n2114 GNDA.n2035 23.6449
R3567 GNDA.n1874 GNDA.n1873 23.6449
R3568 GNDA.n1632 GNDA.n1631 23.6449
R3569 GNDA.n531 GNDA.n489 23.6449
R3570 GNDA.n736 GNDA.n698 23.6449
R3571 GNDA.n959 GNDA.n958 23.6449
R3572 GNDA.n1121 GNDA.n406 23.6449
R3573 GNDA.n1778 GNDA.n1777 23.6449
R3574 GNDA.n293 GNDA.n292 23.6449
R3575 GNDA.n1508 GNDA.n1329 23.5719
R3576 GNDA.n1479 GNDA.n122 21.4917
R3577 GNDA.n1955 GNDA.n1953 21.3338
R3578 GNDA.n66 GNDA.n65 21.3338
R3579 GNDA.n2023 GNDA.n61 21.3338
R3580 GNDA.n2021 GNDA.n62 21.3338
R3581 GNDA.n1966 GNDA.n1951 21.3338
R3582 GNDA.n1964 GNDA.n1952 21.3338
R3583 GNDA.t37 GNDA.n1507 21.0699
R3584 GNDA.n119 GNDA.n118 19.4279
R3585 GNDA.n1491 GNDA.n1478 19.2005
R3586 GNDA.n1479 GNDA.n1309 19.2005
R3587 GNDA.n1505 GNDA.n244 19.2005
R3588 GNDA.n1568 GNDA.n1567 19.2005
R3589 GNDA.n2006 GNDA.n2005 19.2005
R3590 GNDA.n1988 GNDA.n1987 19.2005
R3591 GNDA.n1967 GNDA.n1950 18.3355
R3592 GNDA.n2007 GNDA.n2006 17.613
R3593 GNDA.n1949 GNDA.n1948 17.4917
R3594 GNDA.n1036 GNDA.n1035 17.0672
R3595 GNDA.n2169 GNDA.n30 17.0672
R3596 GNDA.n612 GNDA.n611 17.0672
R3597 GNDA.n1944 GNDA.n1943 16.9605
R3598 GNDA.n2047 GNDA.n2046 16.0005
R3599 GNDA.n2089 GNDA.n2046 16.0005
R3600 GNDA.n2090 GNDA.n2089 16.0005
R3601 GNDA.n2091 GNDA.n2090 16.0005
R3602 GNDA.n2091 GNDA.n2044 16.0005
R3603 GNDA.n2044 GNDA.n2043 16.0005
R3604 GNDA.n2098 GNDA.n2043 16.0005
R3605 GNDA.n2099 GNDA.n2098 16.0005
R3606 GNDA.n2114 GNDA.n2113 16.0005
R3607 GNDA.n2113 GNDA.n2112 16.0005
R3608 GNDA.n2112 GNDA.n2037 16.0005
R3609 GNDA.n2107 GNDA.n2037 16.0005
R3610 GNDA.n2107 GNDA.n2106 16.0005
R3611 GNDA.n2106 GNDA.n2105 16.0005
R3612 GNDA.n2105 GNDA.n2040 16.0005
R3613 GNDA.n2100 GNDA.n2040 16.0005
R3614 GNDA.n2132 GNDA.n2131 16.0005
R3615 GNDA.n2131 GNDA.n2032 16.0005
R3616 GNDA.n2126 GNDA.n2032 16.0005
R3617 GNDA.n2126 GNDA.n2125 16.0005
R3618 GNDA.n2125 GNDA.n2124 16.0005
R3619 GNDA.n2120 GNDA.n2119 16.0005
R3620 GNDA.n2119 GNDA.n2035 16.0005
R3621 GNDA.n1842 GNDA.n164 16.0005
R3622 GNDA.n1844 GNDA.n1842 16.0005
R3623 GNDA.n1845 GNDA.n1844 16.0005
R3624 GNDA.n1848 GNDA.n1845 16.0005
R3625 GNDA.n1849 GNDA.n1848 16.0005
R3626 GNDA.n1852 GNDA.n1849 16.0005
R3627 GNDA.n1854 GNDA.n1852 16.0005
R3628 GNDA.n1855 GNDA.n1854 16.0005
R3629 GNDA.n1873 GNDA.n1870 16.0005
R3630 GNDA.n1870 GNDA.n1869 16.0005
R3631 GNDA.n1869 GNDA.n1866 16.0005
R3632 GNDA.n1866 GNDA.n1865 16.0005
R3633 GNDA.n1865 GNDA.n1862 16.0005
R3634 GNDA.n1862 GNDA.n1861 16.0005
R3635 GNDA.n1861 GNDA.n1858 16.0005
R3636 GNDA.n1858 GNDA.n1857 16.0005
R3637 GNDA.n1890 GNDA.n1889 16.0005
R3638 GNDA.n1889 GNDA.n1886 16.0005
R3639 GNDA.n1886 GNDA.n1885 16.0005
R3640 GNDA.n1885 GNDA.n1882 16.0005
R3641 GNDA.n1882 GNDA.n1881 16.0005
R3642 GNDA.n1878 GNDA.n1877 16.0005
R3643 GNDA.n1877 GNDA.n1874 16.0005
R3644 GNDA.n1600 GNDA.n1599 16.0005
R3645 GNDA.n1602 GNDA.n1600 16.0005
R3646 GNDA.n1603 GNDA.n1602 16.0005
R3647 GNDA.n1606 GNDA.n1603 16.0005
R3648 GNDA.n1607 GNDA.n1606 16.0005
R3649 GNDA.n1610 GNDA.n1607 16.0005
R3650 GNDA.n1612 GNDA.n1610 16.0005
R3651 GNDA.n1613 GNDA.n1612 16.0005
R3652 GNDA.n1631 GNDA.n1628 16.0005
R3653 GNDA.n1628 GNDA.n1627 16.0005
R3654 GNDA.n1627 GNDA.n1624 16.0005
R3655 GNDA.n1624 GNDA.n1623 16.0005
R3656 GNDA.n1623 GNDA.n1620 16.0005
R3657 GNDA.n1620 GNDA.n1619 16.0005
R3658 GNDA.n1619 GNDA.n1616 16.0005
R3659 GNDA.n1616 GNDA.n1615 16.0005
R3660 GNDA.n1648 GNDA.n1647 16.0005
R3661 GNDA.n1647 GNDA.n1644 16.0005
R3662 GNDA.n1644 GNDA.n1643 16.0005
R3663 GNDA.n1643 GNDA.n1640 16.0005
R3664 GNDA.n1640 GNDA.n1639 16.0005
R3665 GNDA.n1636 GNDA.n1635 16.0005
R3666 GNDA.n1635 GNDA.n1632 16.0005
R3667 GNDA.n1944 GNDA.n123 16.0005
R3668 GNDA.n1948 GNDA.n123 16.0005
R3669 GNDA.n500 GNDA.n467 16.0005
R3670 GNDA.n506 GNDA.n500 16.0005
R3671 GNDA.n507 GNDA.n506 16.0005
R3672 GNDA.n508 GNDA.n507 16.0005
R3673 GNDA.n508 GNDA.n498 16.0005
R3674 GNDA.n498 GNDA.n497 16.0005
R3675 GNDA.n515 GNDA.n497 16.0005
R3676 GNDA.n516 GNDA.n515 16.0005
R3677 GNDA.n531 GNDA.n530 16.0005
R3678 GNDA.n530 GNDA.n529 16.0005
R3679 GNDA.n529 GNDA.n491 16.0005
R3680 GNDA.n524 GNDA.n491 16.0005
R3681 GNDA.n524 GNDA.n523 16.0005
R3682 GNDA.n523 GNDA.n522 16.0005
R3683 GNDA.n522 GNDA.n494 16.0005
R3684 GNDA.n517 GNDA.n494 16.0005
R3685 GNDA.n549 GNDA.n548 16.0005
R3686 GNDA.n548 GNDA.n486 16.0005
R3687 GNDA.n543 GNDA.n486 16.0005
R3688 GNDA.n543 GNDA.n542 16.0005
R3689 GNDA.n542 GNDA.n541 16.0005
R3690 GNDA.n537 GNDA.n536 16.0005
R3691 GNDA.n536 GNDA.n489 16.0005
R3692 GNDA.n789 GNDA.n677 16.0005
R3693 GNDA.n711 GNDA.n677 16.0005
R3694 GNDA.n712 GNDA.n711 16.0005
R3695 GNDA.n713 GNDA.n712 16.0005
R3696 GNDA.n713 GNDA.n707 16.0005
R3697 GNDA.n707 GNDA.n706 16.0005
R3698 GNDA.n720 GNDA.n706 16.0005
R3699 GNDA.n721 GNDA.n720 16.0005
R3700 GNDA.n736 GNDA.n735 16.0005
R3701 GNDA.n735 GNDA.n734 16.0005
R3702 GNDA.n734 GNDA.n700 16.0005
R3703 GNDA.n729 GNDA.n700 16.0005
R3704 GNDA.n729 GNDA.n728 16.0005
R3705 GNDA.n728 GNDA.n727 16.0005
R3706 GNDA.n727 GNDA.n703 16.0005
R3707 GNDA.n722 GNDA.n703 16.0005
R3708 GNDA.n754 GNDA.n753 16.0005
R3709 GNDA.n753 GNDA.n695 16.0005
R3710 GNDA.n748 GNDA.n695 16.0005
R3711 GNDA.n748 GNDA.n747 16.0005
R3712 GNDA.n747 GNDA.n746 16.0005
R3713 GNDA.n742 GNDA.n741 16.0005
R3714 GNDA.n741 GNDA.n698 16.0005
R3715 GNDA.n927 GNDA.n926 16.0005
R3716 GNDA.n929 GNDA.n927 16.0005
R3717 GNDA.n930 GNDA.n929 16.0005
R3718 GNDA.n933 GNDA.n930 16.0005
R3719 GNDA.n934 GNDA.n933 16.0005
R3720 GNDA.n937 GNDA.n934 16.0005
R3721 GNDA.n939 GNDA.n937 16.0005
R3722 GNDA.n940 GNDA.n939 16.0005
R3723 GNDA.n958 GNDA.n955 16.0005
R3724 GNDA.n955 GNDA.n954 16.0005
R3725 GNDA.n954 GNDA.n951 16.0005
R3726 GNDA.n951 GNDA.n950 16.0005
R3727 GNDA.n950 GNDA.n947 16.0005
R3728 GNDA.n947 GNDA.n946 16.0005
R3729 GNDA.n946 GNDA.n943 16.0005
R3730 GNDA.n943 GNDA.n942 16.0005
R3731 GNDA.n975 GNDA.n974 16.0005
R3732 GNDA.n974 GNDA.n971 16.0005
R3733 GNDA.n971 GNDA.n970 16.0005
R3734 GNDA.n970 GNDA.n967 16.0005
R3735 GNDA.n967 GNDA.n966 16.0005
R3736 GNDA.n963 GNDA.n962 16.0005
R3737 GNDA.n962 GNDA.n959 16.0005
R3738 GNDA.n418 GNDA.n417 16.0005
R3739 GNDA.n1096 GNDA.n417 16.0005
R3740 GNDA.n1097 GNDA.n1096 16.0005
R3741 GNDA.n1098 GNDA.n1097 16.0005
R3742 GNDA.n1098 GNDA.n415 16.0005
R3743 GNDA.n415 GNDA.n414 16.0005
R3744 GNDA.n1105 GNDA.n414 16.0005
R3745 GNDA.n1106 GNDA.n1105 16.0005
R3746 GNDA.n1121 GNDA.n1120 16.0005
R3747 GNDA.n1120 GNDA.n1119 16.0005
R3748 GNDA.n1119 GNDA.n408 16.0005
R3749 GNDA.n1114 GNDA.n408 16.0005
R3750 GNDA.n1114 GNDA.n1113 16.0005
R3751 GNDA.n1113 GNDA.n1112 16.0005
R3752 GNDA.n1112 GNDA.n411 16.0005
R3753 GNDA.n1107 GNDA.n411 16.0005
R3754 GNDA.n1139 GNDA.n1138 16.0005
R3755 GNDA.n1138 GNDA.n403 16.0005
R3756 GNDA.n1133 GNDA.n403 16.0005
R3757 GNDA.n1133 GNDA.n1132 16.0005
R3758 GNDA.n1132 GNDA.n1131 16.0005
R3759 GNDA.n1127 GNDA.n1126 16.0005
R3760 GNDA.n1126 GNDA.n406 16.0005
R3761 GNDA.n1746 GNDA.n206 16.0005
R3762 GNDA.n1748 GNDA.n1746 16.0005
R3763 GNDA.n1749 GNDA.n1748 16.0005
R3764 GNDA.n1752 GNDA.n1749 16.0005
R3765 GNDA.n1753 GNDA.n1752 16.0005
R3766 GNDA.n1756 GNDA.n1753 16.0005
R3767 GNDA.n1758 GNDA.n1756 16.0005
R3768 GNDA.n1759 GNDA.n1758 16.0005
R3769 GNDA.n1777 GNDA.n1774 16.0005
R3770 GNDA.n1774 GNDA.n1773 16.0005
R3771 GNDA.n1773 GNDA.n1770 16.0005
R3772 GNDA.n1770 GNDA.n1769 16.0005
R3773 GNDA.n1769 GNDA.n1766 16.0005
R3774 GNDA.n1766 GNDA.n1765 16.0005
R3775 GNDA.n1765 GNDA.n1762 16.0005
R3776 GNDA.n1762 GNDA.n1761 16.0005
R3777 GNDA.n1794 GNDA.n1793 16.0005
R3778 GNDA.n1793 GNDA.n1790 16.0005
R3779 GNDA.n1790 GNDA.n1789 16.0005
R3780 GNDA.n1789 GNDA.n1786 16.0005
R3781 GNDA.n1786 GNDA.n1785 16.0005
R3782 GNDA.n1782 GNDA.n1781 16.0005
R3783 GNDA.n1781 GNDA.n1778 16.0005
R3784 GNDA.n325 GNDA.n324 16.0005
R3785 GNDA.n324 GNDA.n323 16.0005
R3786 GNDA.n323 GNDA.n321 16.0005
R3787 GNDA.n321 GNDA.n318 16.0005
R3788 GNDA.n318 GNDA.n317 16.0005
R3789 GNDA.n317 GNDA.n314 16.0005
R3790 GNDA.n314 GNDA.n313 16.0005
R3791 GNDA.n313 GNDA.n311 16.0005
R3792 GNDA.n296 GNDA.n293 16.0005
R3793 GNDA.n297 GNDA.n296 16.0005
R3794 GNDA.n300 GNDA.n297 16.0005
R3795 GNDA.n301 GNDA.n300 16.0005
R3796 GNDA.n304 GNDA.n301 16.0005
R3797 GNDA.n305 GNDA.n304 16.0005
R3798 GNDA.n308 GNDA.n305 16.0005
R3799 GNDA.n310 GNDA.n308 16.0005
R3800 GNDA.n277 GNDA.n276 16.0005
R3801 GNDA.n280 GNDA.n277 16.0005
R3802 GNDA.n281 GNDA.n280 16.0005
R3803 GNDA.n284 GNDA.n281 16.0005
R3804 GNDA.n285 GNDA.n284 16.0005
R3805 GNDA.n289 GNDA.n288 16.0005
R3806 GNDA.n292 GNDA.n289 16.0005
R3807 GNDA.t8 GNDA.t32 15.7148
R3808 GNDA.n1495 GNDA.n1329 15.7148
R3809 GNDA.t5 GNDA.t17 15.7148
R3810 GNDA.n1686 GNDA.n386 15.5383
R3811 GNDA.n835 GNDA.n834 15.5383
R3812 GNDA.n2193 GNDA.n2192 15.5383
R3813 GNDA.n1433 GNDA.n358 15.5383
R3814 GNDA.n2010 GNDA.n2009 15.363
R3815 GNDA.n2009 GNDA.n74 15.363
R3816 GNDA.n119 GNDA 14.6989
R3817 GNDA.n1987 GNDA.n76 13.8005
R3818 GNDA.n1950 GNDA.n1949 13.7706
R3819 GNDA.n2120 GNDA 12.9783
R3820 GNDA.n1878 GNDA 12.9783
R3821 GNDA.n1636 GNDA 12.9783
R3822 GNDA.n537 GNDA 12.9783
R3823 GNDA.n742 GNDA 12.9783
R3824 GNDA.n963 GNDA 12.9783
R3825 GNDA.n1127 GNDA 12.9783
R3826 GNDA.n1782 GNDA 12.9783
R3827 GNDA.n288 GNDA 12.9783
R3828 GNDA.n1995 GNDA.t41 12.5005
R3829 GNDA.n1994 GNDA.n84 12.5005
R3830 GNDA.n81 GNDA.n80 12.5005
R3831 GNDA.n1303 GNDA.n1201 12.4126
R3832 GNDA.n1455 GNDA.n1348 12.4126
R3833 GNDA.n1558 GNDA.n1522 12.4126
R3834 GNDA.n1496 GNDA.t19 11.7862
R3835 GNDA.n866 GNDA.n863 11.6369
R3836 GNDA.n1053 GNDA.n866 11.6369
R3837 GNDA.n1053 GNDA.n1052 11.6369
R3838 GNDA.n1052 GNDA.n1051 11.6369
R3839 GNDA.n1051 GNDA.n867 11.6369
R3840 GNDA.n1045 GNDA.n867 11.6369
R3841 GNDA.n1045 GNDA.n1044 11.6369
R3842 GNDA.n1044 GNDA.n1043 11.6369
R3843 GNDA.n1043 GNDA.n874 11.6369
R3844 GNDA.n1037 GNDA.n874 11.6369
R3845 GNDA.n1037 GNDA.n1036 11.6369
R3846 GNDA.n1020 GNDA.n884 11.6369
R3847 GNDA.n1021 GNDA.n1020 11.6369
R3848 GNDA.n1022 GNDA.n1021 11.6369
R3849 GNDA.n1022 GNDA.n882 11.6369
R3850 GNDA.n1027 GNDA.n882 11.6369
R3851 GNDA.n1028 GNDA.n1027 11.6369
R3852 GNDA.n1029 GNDA.n1028 11.6369
R3853 GNDA.n1029 GNDA.n878 11.6369
R3854 GNDA.n1035 GNDA.n878 11.6369
R3855 GNDA.n2066 GNDA.n2064 11.6369
R3856 GNDA.n2068 GNDA.n2066 11.6369
R3857 GNDA.n2068 GNDA.n2067 11.6369
R3858 GNDA.n2067 GNDA.n35 11.6369
R3859 GNDA.n2159 GNDA.n35 11.6369
R3860 GNDA.n2160 GNDA.n2159 11.6369
R3861 GNDA.n2162 GNDA.n2160 11.6369
R3862 GNDA.n2162 GNDA.n2161 11.6369
R3863 GNDA.n2161 GNDA.n30 11.6369
R3864 GNDA.n2185 GNDA.n13 11.6369
R3865 GNDA.n2185 GNDA.n2184 11.6369
R3866 GNDA.n2184 GNDA.n2183 11.6369
R3867 GNDA.n2183 GNDA.n24 11.6369
R3868 GNDA.n2178 GNDA.n24 11.6369
R3869 GNDA.n2178 GNDA.n2177 11.6369
R3870 GNDA.n2177 GNDA.n2176 11.6369
R3871 GNDA.n2176 GNDA.n27 11.6369
R3872 GNDA.n2171 GNDA.n27 11.6369
R3873 GNDA.n2171 GNDA.n2170 11.6369
R3874 GNDA.n2170 GNDA.n2169 11.6369
R3875 GNDA.n594 GNDA.n593 11.6369
R3876 GNDA.n595 GNDA.n594 11.6369
R3877 GNDA.n595 GNDA.n459 11.6369
R3878 GNDA.n601 GNDA.n459 11.6369
R3879 GNDA.n602 GNDA.n601 11.6369
R3880 GNDA.n603 GNDA.n602 11.6369
R3881 GNDA.n603 GNDA.n455 11.6369
R3882 GNDA.n610 GNDA.n455 11.6369
R3883 GNDA.n611 GNDA.n610 11.6369
R3884 GNDA.n633 GNDA.n445 11.6369
R3885 GNDA.n447 GNDA.n445 11.6369
R3886 GNDA.n626 GNDA.n447 11.6369
R3887 GNDA.n626 GNDA.n625 11.6369
R3888 GNDA.n625 GNDA.n624 11.6369
R3889 GNDA.n624 GNDA.n449 11.6369
R3890 GNDA.n619 GNDA.n449 11.6369
R3891 GNDA.n619 GNDA.n618 11.6369
R3892 GNDA.n618 GNDA.n617 11.6369
R3893 GNDA.n617 GNDA.n452 11.6369
R3894 GNDA.n612 GNDA.n452 11.6369
R3895 GNDA.n1196 GNDA.n1192 11.6369
R3896 GNDA.n1584 GNDA.n1196 11.6369
R3897 GNDA.n1584 GNDA.n1583 11.6369
R3898 GNDA.n1583 GNDA.n1582 11.6369
R3899 GNDA.n1576 GNDA.n1200 11.6369
R3900 GNDA.n1576 GNDA.n1575 11.6369
R3901 GNDA.n1575 GNDA.n1574 11.6369
R3902 GNDA.n1574 GNDA.n1201 11.6369
R3903 GNDA.n1302 GNDA.n1301 11.6369
R3904 GNDA.n1301 GNDA.n1206 11.6369
R3905 GNDA.n1295 GNDA.n1206 11.6369
R3906 GNDA.n1295 GNDA.n1294 11.6369
R3907 GNDA.n1294 GNDA.n1293 11.6369
R3908 GNDA.n1293 GNDA.n1210 11.6369
R3909 GNDA.n1214 GNDA.n1210 11.6369
R3910 GNDA.n1285 GNDA.n1214 11.6369
R3911 GNDA.n1285 GNDA.n1284 11.6369
R3912 GNDA.n1284 GNDA.n1283 11.6369
R3913 GNDA.n1283 GNDA.n1215 11.6369
R3914 GNDA.n1265 GNDA.n1262 11.6369
R3915 GNDA.n1270 GNDA.n1265 11.6369
R3916 GNDA.n1270 GNDA.n1269 11.6369
R3917 GNDA.n1269 GNDA.n1268 11.6369
R3918 GNDA.n1268 GNDA.n126 11.6369
R3919 GNDA.n1942 GNDA.n127 11.6369
R3920 GNDA.n1936 GNDA.n127 11.6369
R3921 GNDA.n1936 GNDA.n1935 11.6369
R3922 GNDA.n1935 GNDA.n1934 11.6369
R3923 GNDA.n1934 GNDA.n132 11.6369
R3924 GNDA.n1343 GNDA.n1342 11.6369
R3925 GNDA.n1471 GNDA.n1343 11.6369
R3926 GNDA.n1471 GNDA.n1470 11.6369
R3927 GNDA.n1470 GNDA.n1469 11.6369
R3928 GNDA.n1463 GNDA.n1347 11.6369
R3929 GNDA.n1463 GNDA.n1462 11.6369
R3930 GNDA.n1462 GNDA.n1461 11.6369
R3931 GNDA.n1461 GNDA.n1348 11.6369
R3932 GNDA.n1454 GNDA.n1453 11.6369
R3933 GNDA.n1453 GNDA.n1350 11.6369
R3934 GNDA.n1448 GNDA.n1350 11.6369
R3935 GNDA.n1448 GNDA.n1447 11.6369
R3936 GNDA.n1447 GNDA.n1446 11.6369
R3937 GNDA.n1446 GNDA.n1353 11.6369
R3938 GNDA.n1441 GNDA.n1353 11.6369
R3939 GNDA.n1441 GNDA.n1440 11.6369
R3940 GNDA.n1440 GNDA.n1439 11.6369
R3941 GNDA.n1439 GNDA.n1356 11.6369
R3942 GNDA.n1434 GNDA.n1356 11.6369
R3943 GNDA.n1511 GNDA.n1322 11.6369
R3944 GNDA.n1512 GNDA.n1511 11.6369
R3945 GNDA.n1514 GNDA.n1512 11.6369
R3946 GNDA.n1514 GNDA.n1513 11.6369
R3947 GNDA.n1521 GNDA.n1520 11.6369
R3948 GNDA.n1560 GNDA.n1521 11.6369
R3949 GNDA.n1560 GNDA.n1559 11.6369
R3950 GNDA.n1559 GNDA.n1558 11.6369
R3951 GNDA.n1532 GNDA.n1531 11.6369
R3952 GNDA.n1535 GNDA.n1532 11.6369
R3953 GNDA.n1536 GNDA.n1535 11.6369
R3954 GNDA.n1539 GNDA.n1536 11.6369
R3955 GNDA.n1540 GNDA.n1539 11.6369
R3956 GNDA.n1543 GNDA.n1540 11.6369
R3957 GNDA.n1544 GNDA.n1543 11.6369
R3958 GNDA.n1547 GNDA.n1544 11.6369
R3959 GNDA.n1548 GNDA.n1547 11.6369
R3960 GNDA.n1550 GNDA.n1548 11.6369
R3961 GNDA.n1550 GNDA.n1549 11.6369
R3962 GNDA.n642 GNDA.n641 11.6369
R3963 GNDA.n645 GNDA.n642 11.6369
R3964 GNDA.n646 GNDA.n645 11.6369
R3965 GNDA.n649 GNDA.n646 11.6369
R3966 GNDA.n650 GNDA.n649 11.6369
R3967 GNDA.n653 GNDA.n650 11.6369
R3968 GNDA.n655 GNDA.n653 11.6369
R3969 GNDA.n656 GNDA.n655 11.6369
R3970 GNDA.n657 GNDA.n656 11.6369
R3971 GNDA.n657 GNDA.n634 11.6369
R3972 GNDA.n833 GNDA.n634 11.6369
R3973 GNDA.n1432 GNDA.n1406 11.6369
R3974 GNDA.n1408 GNDA.n1406 11.6369
R3975 GNDA.n1425 GNDA.n1408 11.6369
R3976 GNDA.n1425 GNDA.n1424 11.6369
R3977 GNDA.n1424 GNDA.n1423 11.6369
R3978 GNDA.n1423 GNDA.n1410 11.6369
R3979 GNDA.n1418 GNDA.n1410 11.6369
R3980 GNDA.n1418 GNDA.n1417 11.6369
R3981 GNDA.n1417 GNDA.n1416 11.6369
R3982 GNDA.n1416 GNDA.n12 11.6369
R3983 GNDA.n2194 GNDA.n12 11.6369
R3984 GNDA.n1192 GNDA.n1191 11.3514
R3985 GNDA.n1342 GNDA.n1334 11.3514
R3986 GNDA.n1322 GNDA.n250 11.3514
R3987 GNDA.n1012 GNDA.n884 11.249
R3988 GNDA.n2064 GNDA.n2062 11.249
R3989 GNDA.n593 GNDA.n464 11.249
R3990 GNDA.n1943 GNDA.n1942 10.4732
R3991 GNDA.n1200 GNDA 10.3439
R3992 GNDA.n1347 GNDA 10.3439
R3993 GNDA.n1520 GNDA 10.3439
R3994 GNDA.n2008 GNDA.n75 9.78488
R3995 GNDA.n77 GNDA.t109 9.6005
R3996 GNDA.n77 GNDA.t110 9.6005
R3997 GNDA.n1986 GNDA.t107 9.6005
R3998 GNDA.n1986 GNDA.t108 9.6005
R3999 GNDA.n117 GNDA.n76 9.37925
R4000 GNDA.n1303 GNDA.n1302 8.79242
R4001 GNDA.n1455 GNDA.n1454 8.79242
R4002 GNDA.n1531 GNDA.n1522 8.79242
R4003 GNDA.n863 GNDA.n861 8.53383
R4004 GNDA.n2193 GNDA.n13 8.53383
R4005 GNDA.n834 GNDA.n633 8.53383
R4006 GNDA.n1262 GNDA.n1260 8.53383
R4007 GNDA.n641 GNDA.n386 8.53383
R4008 GNDA.n1433 GNDA.n1432 8.53383
R4009 GNDA.n2051 GNDA.n2047 8.35606
R4010 GNDA.n1926 GNDA.n164 8.35606
R4011 GNDA.n1599 GNDA.n1153 8.35606
R4012 GNDA.n584 GNDA.n467 8.35606
R4013 GNDA.n790 GNDA.n789 8.35606
R4014 GNDA.n926 GNDA.n888 8.35606
R4015 GNDA.n1085 GNDA.n418 8.35606
R4016 GNDA.n1831 GNDA.n206 8.35606
R4017 GNDA.n326 GNDA.n325 8.35606
R4018 GNDA.n2009 GNDA.n2008 7.71925
R4019 GNDA.n1498 GNDA.n1478 6.4005
R4020 GNDA.n115 GNDA.n114 6.0355
R4021 GNDA.n1597 GNDA.n1186 4.6085
R4022 GNDA.n1744 GNDA.n238 4.6085
R4023 GNDA.n1729 GNDA.n1728 4.6085
R4024 GNDA.n1063 GNDA.n1060 4.55161
R4025 GNDA.n830 GNDA.n444 4.55161
R4026 GNDA.n1278 GNDA.n1277 4.55161
R4027 GNDA.n1691 GNDA.n1690 4.55161
R4028 GNDA.n1405 GNDA.n1404 4.55161
R4029 GNDA.n2197 GNDA.n9 4.55161
R4030 GNDA.n2008 GNDA.n2007 4.5005
R4031 GNDA.n1260 GNDA.n1215 4.39646
R4032 GNDA.n861 GNDA.n132 4.39646
R4033 GNDA.n1434 GNDA.n1433 4.39646
R4034 GNDA.n1549 GNDA.n386 4.39646
R4035 GNDA.n834 GNDA.n833 4.39646
R4036 GNDA.n2194 GNDA.n2193 4.39646
R4037 GNDA.n1012 GNDA.n1011 4.3013
R4038 GNDA.n585 GNDA.n464 4.3013
R4039 GNDA.n1079 GNDA.n837 4.26717
R4040 GNDA.n1079 GNDA.n1078 4.26717
R4041 GNDA.n1078 GNDA.n1077 4.26717
R4042 GNDA.n1077 GNDA.n843 4.26717
R4043 GNDA.n1072 GNDA.n843 4.26717
R4044 GNDA.n1072 GNDA.n1071 4.26717
R4045 GNDA.n1070 GNDA.n852 4.26717
R4046 GNDA.n1065 GNDA.n852 4.26717
R4047 GNDA.n1065 GNDA.n1064 4.26717
R4048 GNDA.n1064 GNDA.n1063 4.26717
R4049 GNDA.n797 GNDA.n672 4.26717
R4050 GNDA.n803 GNDA.n672 4.26717
R4051 GNDA.n803 GNDA.n670 4.26717
R4052 GNDA.n809 GNDA.n670 4.26717
R4053 GNDA.n809 GNDA.n668 4.26717
R4054 GNDA.n815 GNDA.n668 4.26717
R4055 GNDA.n823 GNDA.n666 4.26717
R4056 GNDA.n823 GNDA.n664 4.26717
R4057 GNDA.n664 GNDA.n663 4.26717
R4058 GNDA.n830 GNDA.n663 4.26717
R4059 GNDA.n1228 GNDA.n1152 4.26717
R4060 GNDA.n1233 GNDA.n1228 4.26717
R4061 GNDA.n1233 GNDA.n1224 4.26717
R4062 GNDA.n1239 GNDA.n1224 4.26717
R4063 GNDA.n1239 GNDA.n1222 4.26717
R4064 GNDA.n1244 GNDA.n1222 4.26717
R4065 GNDA.n1249 GNDA.n1219 4.26717
R4066 GNDA.n1255 GNDA.n1219 4.26717
R4067 GNDA.n1255 GNDA.n1217 4.26717
R4068 GNDA.n1278 GNDA.n1217 4.26717
R4069 GNDA.n1711 GNDA.n1710 4.26717
R4070 GNDA.n1710 GNDA.n362 4.26717
R4071 GNDA.n1705 GNDA.n362 4.26717
R4072 GNDA.n1705 GNDA.n1704 4.26717
R4073 GNDA.n1704 GNDA.n1703 4.26717
R4074 GNDA.n1703 GNDA.n371 4.26717
R4075 GNDA.n1698 GNDA.n1697 4.26717
R4076 GNDA.n1697 GNDA.n1696 4.26717
R4077 GNDA.n1696 GNDA.n380 4.26717
R4078 GNDA.n1691 GNDA.n380 4.26717
R4079 GNDA.n1371 GNDA.n1370 4.26717
R4080 GNDA.n1376 GNDA.n1371 4.26717
R4081 GNDA.n1376 GNDA.n1366 4.26717
R4082 GNDA.n1382 GNDA.n1366 4.26717
R4083 GNDA.n1382 GNDA.n1364 4.26717
R4084 GNDA.n1387 GNDA.n1364 4.26717
R4085 GNDA.n1392 GNDA.n1361 4.26717
R4086 GNDA.n1399 GNDA.n1361 4.26717
R4087 GNDA.n1399 GNDA.n1359 4.26717
R4088 GNDA.n1404 GNDA.n1359 4.26717
R4089 GNDA.n160 GNDA.n137 4.26717
R4090 GNDA.n160 GNDA.n159 4.26717
R4091 GNDA.n159 GNDA.n158 4.26717
R4092 GNDA.n158 GNDA.n145 4.26717
R4093 GNDA.n153 GNDA.n145 4.26717
R4094 GNDA.n153 GNDA.n0 4.26717
R4095 GNDA.n2204 GNDA.n2 4.26717
R4096 GNDA.n2199 GNDA.n2 4.26717
R4097 GNDA.n2199 GNDA.n2198 4.26717
R4098 GNDA.n2198 GNDA.n2197 4.26717
R4099 GNDA.n2062 GNDA.n2061 4.1989
R4100 GNDA.n1485 GNDA.t6 3.92907
R4101 GNDA.n1494 GNDA.t30 3.92907
R4102 GNDA.n1508 GNDA.t5 3.92907
R4103 GNDA.n2007 GNDA.n76 3.813
R4104 GNDA GNDA.n1070 3.79309
R4105 GNDA GNDA.n666 3.79309
R4106 GNDA.n1249 GNDA 3.79309
R4107 GNDA.n1698 GNDA 3.79309
R4108 GNDA.n1392 GNDA 3.79309
R4109 GNDA GNDA.n2204 3.79309
R4110 GNDA GNDA.n117 3.68412
R4111 GNDA.n760 GNDA.n758 3.5845
R4112 GNDA.n759 GNDA.n687 3.5845
R4113 GNDA.n767 GNDA.n766 3.5845
R4114 GNDA.n685 GNDA.n684 3.5845
R4115 GNDA.n775 GNDA.n773 3.5845
R4116 GNDA.n774 GNDA.n682 3.5845
R4117 GNDA.n782 GNDA.n781 3.5845
R4118 GNDA.n680 GNDA.n679 3.5845
R4119 GNDA.n791 GNDA.n676 3.5845
R4120 GNDA.n1145 GNDA.n399 3.5845
R4121 GNDA.n1144 GNDA.n400 3.5845
R4122 GNDA.n428 GNDA.n426 3.5845
R4123 GNDA.n432 GNDA.n429 3.5845
R4124 GNDA.n433 GNDA.n421 3.5845
R4125 GNDA.n438 GNDA.n437 3.5845
R4126 GNDA.n441 GNDA.n420 3.5845
R4127 GNDA.n443 GNDA.n442 3.5845
R4128 GNDA.n1089 GNDA.n1088 3.5845
R4129 GNDA.n982 GNDA.n978 3.5845
R4130 GNDA.n981 GNDA.n916 3.5845
R4131 GNDA.n988 GNDA.n915 3.5845
R4132 GNDA.n989 GNDA.n914 3.5845
R4133 GNDA.n994 GNDA.n992 3.5845
R4134 GNDA.n993 GNDA.n911 3.5845
R4135 GNDA.n1001 GNDA.n1000 3.5845
R4136 GNDA.n912 GNDA.n890 3.5845
R4137 GNDA.n1007 GNDA.n1006 3.5845
R4138 GNDA.n555 GNDA.n553 3.5845
R4139 GNDA.n554 GNDA.n478 3.5845
R4140 GNDA.n562 GNDA.n561 3.5845
R4141 GNDA.n476 GNDA.n475 3.5845
R4142 GNDA.n569 GNDA.n568 3.5845
R4143 GNDA.n574 GNDA.n473 3.5845
R4144 GNDA.n575 GNDA.n470 3.5845
R4145 GNDA.n580 GNDA.n579 3.5845
R4146 GNDA.n583 GNDA.n468 3.5845
R4147 GNDA.n1655 GNDA.n1651 3.5845
R4148 GNDA.n1654 GNDA.n1183 3.5845
R4149 GNDA.n1661 GNDA.n1182 3.5845
R4150 GNDA.n1662 GNDA.n1181 3.5845
R4151 GNDA.n1667 GNDA.n1665 3.5845
R4152 GNDA.n1666 GNDA.n1178 3.5845
R4153 GNDA.n1674 GNDA.n1673 3.5845
R4154 GNDA.n1179 GNDA.n1157 3.5845
R4155 GNDA.n1680 GNDA.n1679 3.5845
R4156 GNDA.n1802 GNDA.n1797 3.5845
R4157 GNDA.n1801 GNDA.n1798 3.5845
R4158 GNDA.n1810 GNDA.n234 3.5845
R4159 GNDA.n1811 GNDA.n233 3.5845
R4160 GNDA.n1816 GNDA.n1814 3.5845
R4161 GNDA.n1815 GNDA.n228 3.5845
R4162 GNDA.n1824 GNDA.n1823 3.5845
R4163 GNDA.n229 GNDA.n207 3.5845
R4164 GNDA.n1830 GNDA.n1829 3.5845
R4165 GNDA.n1723 GNDA.n253 3.5845
R4166 GNDA.n335 GNDA.n334 3.5845
R4167 GNDA.n338 GNDA.n332 3.5845
R4168 GNDA.n342 GNDA.n341 3.5845
R4169 GNDA.n346 GNDA.n329 3.5845
R4170 GNDA.n347 GNDA.n328 3.5845
R4171 GNDA.n352 GNDA.n350 3.5845
R4172 GNDA.n351 GNDA.n275 3.5845
R4173 GNDA.n1718 GNDA.n1717 3.5845
R4174 GNDA.n1898 GNDA.n1893 3.5845
R4175 GNDA.n1897 GNDA.n1894 3.5845
R4176 GNDA.n1905 GNDA.n192 3.5845
R4177 GNDA.n1906 GNDA.n191 3.5845
R4178 GNDA.n1911 GNDA.n1909 3.5845
R4179 GNDA.n1910 GNDA.n186 3.5845
R4180 GNDA.n1919 GNDA.n1918 3.5845
R4181 GNDA.n187 GNDA.n165 3.5845
R4182 GNDA.n1925 GNDA.n1924 3.5845
R4183 GNDA.n2138 GNDA.n2136 3.5845
R4184 GNDA.n2137 GNDA.n48 3.5845
R4185 GNDA.n2145 GNDA.n2144 3.5845
R4186 GNDA.n46 GNDA.n45 3.5845
R4187 GNDA.n2153 GNDA.n42 3.5845
R4188 GNDA.n2152 GNDA.n43 3.5845
R4189 GNDA.n2056 GNDA.n2054 3.5845
R4190 GNDA.n2055 GNDA.n2050 3.5845
R4191 GNDA.n2082 GNDA.n2081 3.5845
R4192 GNDA.n1712 GNDA.n357 3.3797
R4193 GNDA.n790 GNDA.n673 3.3797
R4194 GNDA.n1685 GNDA.n1151 3.3797
R4195 GNDA.n1085 GNDA.n1084 3.3797
R4196 GNDA.n924 GNDA.n836 3.3797
R4197 GNDA.n1011 GNDA.n888 3.3797
R4198 GNDA.n484 GNDA.n14 3.3797
R4199 GNDA.n585 GNDA.n584 3.3797
R4200 GNDA.n1684 GNDA.n1153 3.3797
R4201 GNDA.n1832 GNDA.n1831 3.3797
R4202 GNDA.n1713 GNDA.n326 3.3797
R4203 GNDA.n1840 GNDA.n197 3.3797
R4204 GNDA.n1927 GNDA.n1926 3.3797
R4205 GNDA.n2030 GNDA.n54 3.3797
R4206 GNDA.n2061 GNDA.n2051 3.3797
R4207 GNDA.n836 GNDA.n835 3.27161
R4208 GNDA.n2192 GNDA.n14 3.27161
R4209 GNDA.n1686 GNDA.n1685 3.27161
R4210 GNDA.n1712 GNDA.n358 3.27161
R4211 GNDA.n102 GNDA.n100 3.21925
R4212 GNDA.n110 GNDA.n108 3.21925
R4213 GNDA.n1492 GNDA.n1491 3.2005
R4214 GNDA.n1504 GNDA.n1477 3.2005
R4215 GNDA.n2124 GNDA 3.02272
R4216 GNDA.n1881 GNDA 3.02272
R4217 GNDA.n1639 GNDA 3.02272
R4218 GNDA.n541 GNDA 3.02272
R4219 GNDA.n746 GNDA 3.02272
R4220 GNDA.n966 GNDA 3.02272
R4221 GNDA.n1131 GNDA 3.02272
R4222 GNDA.n1785 GNDA 3.02272
R4223 GNDA.n285 GNDA 3.02272
R4224 GNDA.n694 GNDA.n692 2.8677
R4225 GNDA.n398 GNDA.n391 2.8677
R4226 GNDA.n925 GNDA.n918 2.8677
R4227 GNDA.n485 GNDA.n480 2.8677
R4228 GNDA.n1598 GNDA.n1185 2.8677
R4229 GNDA.n1745 GNDA.n237 2.8677
R4230 GNDA.n1724 GNDA.n251 2.8677
R4231 GNDA.n1841 GNDA.n196 2.8677
R4232 GNDA.n2031 GNDA.n52 2.8677
R4233 GNDA.n2132 GNDA.n2031 2.31161
R4234 GNDA.n1890 GNDA.n1841 2.31161
R4235 GNDA.n1648 GNDA.n1598 2.31161
R4236 GNDA.n549 GNDA.n485 2.31161
R4237 GNDA.n754 GNDA.n694 2.31161
R4238 GNDA.n975 GNDA.n925 2.31161
R4239 GNDA.n1139 GNDA.n391 2.31161
R4240 GNDA.n1794 GNDA.n1745 2.31161
R4241 GNDA.n276 GNDA.n251 2.31161
R4242 GNDA.n1836 GNDA.n198 1.951
R4243 GNDA.n56 GNDA.n55 1.951
R4244 GNDA.n688 GNDA.n389 1.951
R4245 GNDA.n2191 GNDA.n15 1.951
R4246 GNDA.n1687 GNDA.n390 1.951
R4247 GNDA.n921 GNDA.n21 1.951
R4248 GNDA.n1594 GNDA.n1187 1.951
R4249 GNDA.n240 GNDA.n239 1.951
R4250 GNDA.n1730 GNDA.n249 1.951
R4251 GNDA.n694 GNDA.n357 1.7413
R4252 GNDA.n673 GNDA.n14 1.7413
R4253 GNDA.n1151 GNDA.n391 1.7413
R4254 GNDA.n1084 GNDA.n836 1.7413
R4255 GNDA.n925 GNDA.n924 1.7413
R4256 GNDA.n485 GNDA.n484 1.7413
R4257 GNDA.n1598 GNDA.n1597 1.7413
R4258 GNDA.n1685 GNDA.n1684 1.7413
R4259 GNDA.n1745 GNDA.n1744 1.7413
R4260 GNDA.n1832 GNDA.n197 1.7413
R4261 GNDA.n1728 GNDA.n251 1.7413
R4262 GNDA.n1713 GNDA.n1712 1.7413
R4263 GNDA.n1841 GNDA.n1840 1.7413
R4264 GNDA.n1927 GNDA.n54 1.7413
R4265 GNDA.n2031 GNDA.n2030 1.7413
R4266 GNDA.n1949 GNDA.n122 1.73362
R4267 GNDA.n837 GNDA.n836 1.51754
R4268 GNDA.n797 GNDA.n14 1.51754
R4269 GNDA.n1685 GNDA.n1152 1.51754
R4270 GNDA.n1712 GNDA.n1711 1.51754
R4271 GNDA.n1370 GNDA.n197 1.51754
R4272 GNDA.n137 GNDA.n54 1.51754
R4273 GNDA.n1582 GNDA 1.29343
R4274 GNDA.n1469 GNDA 1.29343
R4275 GNDA.n1513 GNDA 1.29343
R4276 GNDA.n791 GNDA.n790 1.2293
R4277 GNDA.n1088 GNDA.n1085 1.2293
R4278 GNDA.n1007 GNDA.n888 1.2293
R4279 GNDA.n584 GNDA.n583 1.2293
R4280 GNDA.n1680 GNDA.n1153 1.2293
R4281 GNDA.n1831 GNDA.n1830 1.2293
R4282 GNDA.n1717 GNDA.n326 1.2293
R4283 GNDA.n1926 GNDA.n1925 1.2293
R4284 GNDA.n2081 GNDA.n2051 1.2293
R4285 GNDA.n1191 GNDA.n1186 1.1781
R4286 GNDA.n1334 GNDA.n238 1.1781
R4287 GNDA.n1729 GNDA.n250 1.1781
R4288 GNDA.n1943 GNDA.n126 1.16414
R4289 GNDA.n758 GNDA.n692 1.0245
R4290 GNDA.n760 GNDA.n759 1.0245
R4291 GNDA.n767 GNDA.n687 1.0245
R4292 GNDA.n766 GNDA.n685 1.0245
R4293 GNDA.n773 GNDA.n684 1.0245
R4294 GNDA.n775 GNDA.n774 1.0245
R4295 GNDA.n782 GNDA.n682 1.0245
R4296 GNDA.n781 GNDA.n680 1.0245
R4297 GNDA.n679 GNDA.n676 1.0245
R4298 GNDA.n399 GNDA.n398 1.0245
R4299 GNDA.n1145 GNDA.n1144 1.0245
R4300 GNDA.n426 GNDA.n400 1.0245
R4301 GNDA.n429 GNDA.n428 1.0245
R4302 GNDA.n433 GNDA.n432 1.0245
R4303 GNDA.n437 GNDA.n421 1.0245
R4304 GNDA.n438 GNDA.n420 1.0245
R4305 GNDA.n442 GNDA.n441 1.0245
R4306 GNDA.n1089 GNDA.n443 1.0245
R4307 GNDA.n978 GNDA.n918 1.0245
R4308 GNDA.n982 GNDA.n981 1.0245
R4309 GNDA.n916 GNDA.n915 1.0245
R4310 GNDA.n989 GNDA.n988 1.0245
R4311 GNDA.n992 GNDA.n914 1.0245
R4312 GNDA.n994 GNDA.n993 1.0245
R4313 GNDA.n1001 GNDA.n911 1.0245
R4314 GNDA.n1000 GNDA.n912 1.0245
R4315 GNDA.n1006 GNDA.n890 1.0245
R4316 GNDA.n553 GNDA.n480 1.0245
R4317 GNDA.n555 GNDA.n554 1.0245
R4318 GNDA.n562 GNDA.n478 1.0245
R4319 GNDA.n561 GNDA.n476 1.0245
R4320 GNDA.n568 GNDA.n475 1.0245
R4321 GNDA.n569 GNDA.n473 1.0245
R4322 GNDA.n575 GNDA.n574 1.0245
R4323 GNDA.n579 GNDA.n470 1.0245
R4324 GNDA.n580 GNDA.n468 1.0245
R4325 GNDA.n1651 GNDA.n1185 1.0245
R4326 GNDA.n1655 GNDA.n1654 1.0245
R4327 GNDA.n1183 GNDA.n1182 1.0245
R4328 GNDA.n1662 GNDA.n1661 1.0245
R4329 GNDA.n1665 GNDA.n1181 1.0245
R4330 GNDA.n1667 GNDA.n1666 1.0245
R4331 GNDA.n1674 GNDA.n1178 1.0245
R4332 GNDA.n1673 GNDA.n1179 1.0245
R4333 GNDA.n1679 GNDA.n1157 1.0245
R4334 GNDA.n1797 GNDA.n237 1.0245
R4335 GNDA.n1802 GNDA.n1801 1.0245
R4336 GNDA.n1798 GNDA.n234 1.0245
R4337 GNDA.n1811 GNDA.n1810 1.0245
R4338 GNDA.n1814 GNDA.n233 1.0245
R4339 GNDA.n1816 GNDA.n1815 1.0245
R4340 GNDA.n1824 GNDA.n228 1.0245
R4341 GNDA.n1823 GNDA.n229 1.0245
R4342 GNDA.n1829 GNDA.n207 1.0245
R4343 GNDA.n1724 GNDA.n1723 1.0245
R4344 GNDA.n334 GNDA.n253 1.0245
R4345 GNDA.n335 GNDA.n332 1.0245
R4346 GNDA.n341 GNDA.n338 1.0245
R4347 GNDA.n342 GNDA.n329 1.0245
R4348 GNDA.n347 GNDA.n346 1.0245
R4349 GNDA.n350 GNDA.n328 1.0245
R4350 GNDA.n352 GNDA.n351 1.0245
R4351 GNDA.n1718 GNDA.n275 1.0245
R4352 GNDA.n1893 GNDA.n196 1.0245
R4353 GNDA.n1898 GNDA.n1897 1.0245
R4354 GNDA.n1894 GNDA.n192 1.0245
R4355 GNDA.n1906 GNDA.n1905 1.0245
R4356 GNDA.n1909 GNDA.n191 1.0245
R4357 GNDA.n1911 GNDA.n1910 1.0245
R4358 GNDA.n1919 GNDA.n186 1.0245
R4359 GNDA.n1918 GNDA.n187 1.0245
R4360 GNDA.n1924 GNDA.n165 1.0245
R4361 GNDA.n2136 GNDA.n52 1.0245
R4362 GNDA.n2138 GNDA.n2137 1.0245
R4363 GNDA.n2145 GNDA.n48 1.0245
R4364 GNDA.n2144 GNDA.n46 1.0245
R4365 GNDA.n45 GNDA.n42 1.0245
R4366 GNDA.n2153 GNDA.n2152 1.0245
R4367 GNDA.n2054 GNDA.n43 1.0245
R4368 GNDA.n2056 GNDA.n2055 1.0245
R4369 GNDA.n2082 GNDA.n2050 1.0245
R4370 GNDA.n100 GNDA.n98 1.0005
R4371 GNDA.n104 GNDA.n102 1.0005
R4372 GNDA.n106 GNDA.n104 1.0005
R4373 GNDA.n108 GNDA.n106 1.0005
R4374 GNDA.n112 GNDA.n110 1.0005
R4375 GNDA.n114 GNDA.n112 1.0005
R4376 GNDA.n1071 GNDA 0.474574
R4377 GNDA.n815 GNDA 0.474574
R4378 GNDA.n1244 GNDA 0.474574
R4379 GNDA GNDA.n371 0.474574
R4380 GNDA.n1387 GNDA 0.474574
R4381 GNDA GNDA.n0 0.474574
R4382 GNDA.n120 GNDA.n119 0.41175
R4383 GNDA.n121 GNDA.n120 0.311875
R4384 GNDA.n117 GNDA.n116 0.276625
R4385 GNDA.n116 GNDA.n115 0.22375
R4386 GNDA.n1950 GNDA.n115 0.100375
R4387 GNDA.n1060 GNDA.n861 0.0953148
R4388 GNDA.n834 GNDA.n444 0.0953148
R4389 GNDA.n1277 GNDA.n1260 0.0953148
R4390 GNDA.n1690 GNDA.n386 0.0953148
R4391 GNDA.n1433 GNDA.n1405 0.0953148
R4392 GNDA.n2193 GNDA.n9 0.0953148
R4393 GNDA.n122 GNDA.n121 0.076875
R4394 PFET_GATE_10uA.n23 PFET_GATE_10uA.n21 341.397
R4395 PFET_GATE_10uA.n25 PFET_GATE_10uA.n24 339.272
R4396 PFET_GATE_10uA.n23 PFET_GATE_10uA.n22 339.272
R4397 PFET_GATE_10uA.n28 PFET_GATE_10uA.n27 334.772
R4398 PFET_GATE_10uA.n11 PFET_GATE_10uA.t20 273.134
R4399 PFET_GATE_10uA.n8 PFET_GATE_10uA.t16 273.134
R4400 PFET_GATE_10uA.n5 PFET_GATE_10uA.t27 273.134
R4401 PFET_GATE_10uA.n4 PFET_GATE_10uA.t26 273.134
R4402 PFET_GATE_10uA.n2 PFET_GATE_10uA.t17 273.134
R4403 PFET_GATE_10uA.n1 PFET_GATE_10uA.t24 273.134
R4404 PFET_GATE_10uA.n12 PFET_GATE_10uA.n11 224.934
R4405 PFET_GATE_10uA.n13 PFET_GATE_10uA.n12 224.934
R4406 PFET_GATE_10uA.n9 PFET_GATE_10uA.n8 224.934
R4407 PFET_GATE_10uA.n10 PFET_GATE_10uA.n9 224.934
R4408 PFET_GATE_10uA.n16 PFET_GATE_10uA.n15 224.934
R4409 PFET_GATE_10uA.t2 PFET_GATE_10uA.n29 194.895
R4410 PFET_GATE_10uA.n7 PFET_GATE_10uA.n6 172.363
R4411 PFET_GATE_10uA.n20 PFET_GATE_10uA.n0 169.832
R4412 PFET_GATE_10uA.n19 PFET_GATE_10uA.n3 168.863
R4413 PFET_GATE_10uA.n18 PFET_GATE_10uA.n17 166.05
R4414 PFET_GATE_10uA.n14 PFET_GATE_10uA.n7 166.05
R4415 PFET_GATE_10uA.n0 PFET_GATE_10uA.t29 117.823
R4416 PFET_GATE_10uA.n0 PFET_GATE_10uA.t12 117.823
R4417 PFET_GATE_10uA.n26 PFET_GATE_10uA.t7 100.635
R4418 PFET_GATE_10uA.n14 PFET_GATE_10uA.n13 69.6227
R4419 PFET_GATE_10uA.n17 PFET_GATE_10uA.n10 69.6227
R4420 PFET_GATE_10uA.n17 PFET_GATE_10uA.n16 69.6227
R4421 PFET_GATE_10uA.n15 PFET_GATE_10uA.n14 69.6227
R4422 PFET_GATE_10uA.n6 PFET_GATE_10uA.n5 69.6227
R4423 PFET_GATE_10uA.n6 PFET_GATE_10uA.n4 69.6227
R4424 PFET_GATE_10uA.n3 PFET_GATE_10uA.n2 69.6227
R4425 PFET_GATE_10uA.n3 PFET_GATE_10uA.n1 69.6227
R4426 PFET_GATE_10uA.n11 PFET_GATE_10uA.t25 48.2005
R4427 PFET_GATE_10uA.n12 PFET_GATE_10uA.t28 48.2005
R4428 PFET_GATE_10uA.n13 PFET_GATE_10uA.t11 48.2005
R4429 PFET_GATE_10uA.n8 PFET_GATE_10uA.t14 48.2005
R4430 PFET_GATE_10uA.n9 PFET_GATE_10uA.t13 48.2005
R4431 PFET_GATE_10uA.n10 PFET_GATE_10uA.t10 48.2005
R4432 PFET_GATE_10uA.n16 PFET_GATE_10uA.t23 48.2005
R4433 PFET_GATE_10uA.n15 PFET_GATE_10uA.t21 48.2005
R4434 PFET_GATE_10uA.n5 PFET_GATE_10uA.t15 48.2005
R4435 PFET_GATE_10uA.n4 PFET_GATE_10uA.t18 48.2005
R4436 PFET_GATE_10uA.n2 PFET_GATE_10uA.t19 48.2005
R4437 PFET_GATE_10uA.n1 PFET_GATE_10uA.t22 48.2005
R4438 PFET_GATE_10uA.n27 PFET_GATE_10uA.t1 39.4005
R4439 PFET_GATE_10uA.n27 PFET_GATE_10uA.t8 39.4005
R4440 PFET_GATE_10uA.n24 PFET_GATE_10uA.t5 39.4005
R4441 PFET_GATE_10uA.n24 PFET_GATE_10uA.t0 39.4005
R4442 PFET_GATE_10uA.n22 PFET_GATE_10uA.t3 39.4005
R4443 PFET_GATE_10uA.n22 PFET_GATE_10uA.t4 39.4005
R4444 PFET_GATE_10uA.n21 PFET_GATE_10uA.t9 39.4005
R4445 PFET_GATE_10uA.n21 PFET_GATE_10uA.t6 39.4005
R4446 PFET_GATE_10uA.n20 PFET_GATE_10uA.n19 26.0005
R4447 PFET_GATE_10uA.n29 PFET_GATE_10uA.n28 5.15675
R4448 PFET_GATE_10uA.n28 PFET_GATE_10uA.n26 4.5005
R4449 PFET_GATE_10uA.n29 PFET_GATE_10uA.n20 4.188
R4450 PFET_GATE_10uA.n19 PFET_GATE_10uA.n18 3.3755
R4451 PFET_GATE_10uA.n25 PFET_GATE_10uA.n23 2.1255
R4452 PFET_GATE_10uA.n26 PFET_GATE_10uA.n25 2.1255
R4453 PFET_GATE_10uA.n18 PFET_GATE_10uA.n7 1.0005
R4454 TAIL_CUR_MIR_BIAS.n2 TAIL_CUR_MIR_BIAS.n0 340.272
R4455 TAIL_CUR_MIR_BIAS.n4 TAIL_CUR_MIR_BIAS.n3 339.272
R4456 TAIL_CUR_MIR_BIAS.n2 TAIL_CUR_MIR_BIAS.n1 339.272
R4457 TAIL_CUR_MIR_BIAS.n6 TAIL_CUR_MIR_BIAS.n5 334.772
R4458 TAIL_CUR_MIR_BIAS.n5 TAIL_CUR_MIR_BIAS.t4 39.4005
R4459 TAIL_CUR_MIR_BIAS.n5 TAIL_CUR_MIR_BIAS.t5 39.4005
R4460 TAIL_CUR_MIR_BIAS.n3 TAIL_CUR_MIR_BIAS.t7 39.4005
R4461 TAIL_CUR_MIR_BIAS.n3 TAIL_CUR_MIR_BIAS.t2 39.4005
R4462 TAIL_CUR_MIR_BIAS.n1 TAIL_CUR_MIR_BIAS.t3 39.4005
R4463 TAIL_CUR_MIR_BIAS.n1 TAIL_CUR_MIR_BIAS.t6 39.4005
R4464 TAIL_CUR_MIR_BIAS.n0 TAIL_CUR_MIR_BIAS.t0 39.4005
R4465 TAIL_CUR_MIR_BIAS.n0 TAIL_CUR_MIR_BIAS.t1 39.4005
R4466 TAIL_CUR_MIR_BIAS TAIL_CUR_MIR_BIAS.n6 16.7193
R4467 TAIL_CUR_MIR_BIAS.n6 TAIL_CUR_MIR_BIAS.n4 5.5005
R4468 TAIL_CUR_MIR_BIAS.n4 TAIL_CUR_MIR_BIAS.n2 1.0005
R4469 1st_Vout_1.n9 1st_Vout_1.t32 355.293
R4470 1st_Vout_1.n11 1st_Vout_1.t17 346.8
R4471 1st_Vout_1.n2 1st_Vout_1.n12 339.522
R4472 1st_Vout_1.n9 1st_Vout_1.n8 339.522
R4473 1st_Vout_1.n14 1st_Vout_1.n7 335.022
R4474 1st_Vout_1.t10 1st_Vout_1.n17 275.909
R4475 1st_Vout_1.n17 1st_Vout_1.n6 227.909
R4476 1st_Vout_1.n16 1st_Vout_1.n15 222.034
R4477 1st_Vout_1.n13 1st_Vout_1.t14 184.097
R4478 1st_Vout_1.n13 1st_Vout_1.t18 184.097
R4479 1st_Vout_1.n10 1st_Vout_1.t30 184.097
R4480 1st_Vout_1.n10 1st_Vout_1.t20 184.097
R4481 1st_Vout_1.n2 1st_Vout_1.n13 166.05
R4482 1st_Vout_1.n3 1st_Vout_1.n10 166.05
R4483 1st_Vout_1.n15 1st_Vout_1.t6 48.0005
R4484 1st_Vout_1.n15 1st_Vout_1.t7 48.0005
R4485 1st_Vout_1.n6 1st_Vout_1.t9 48.0005
R4486 1st_Vout_1.n6 1st_Vout_1.t8 48.0005
R4487 1st_Vout_1.n12 1st_Vout_1.t4 39.4005
R4488 1st_Vout_1.n12 1st_Vout_1.t0 39.4005
R4489 1st_Vout_1.n8 1st_Vout_1.t5 39.4005
R4490 1st_Vout_1.n8 1st_Vout_1.t3 39.4005
R4491 1st_Vout_1.n7 1st_Vout_1.t2 39.4005
R4492 1st_Vout_1.n7 1st_Vout_1.t1 39.4005
R4493 1st_Vout_1.n11 1st_Vout_1.n5 33.1711
R4494 1st_Vout_1.n0 1st_Vout_1.t36 4.8295
R4495 1st_Vout_1.n4 1st_Vout_1.t34 4.8295
R4496 1st_Vout_1.n0 1st_Vout_1.t16 4.8295
R4497 1st_Vout_1.n0 1st_Vout_1.t15 4.8295
R4498 1st_Vout_1.n1 1st_Vout_1.t33 4.8295
R4499 1st_Vout_1.n1 1st_Vout_1.t31 4.8295
R4500 1st_Vout_1.n1 1st_Vout_1.t24 4.8295
R4501 1st_Vout_1.n0 1st_Vout_1.t28 4.5005
R4502 1st_Vout_1.n0 1st_Vout_1.t23 4.5005
R4503 1st_Vout_1.n4 1st_Vout_1.t12 4.5005
R4504 1st_Vout_1.n0 1st_Vout_1.t35 4.5005
R4505 1st_Vout_1.n0 1st_Vout_1.t27 4.5005
R4506 1st_Vout_1.n0 1st_Vout_1.t19 4.5005
R4507 1st_Vout_1.n1 1st_Vout_1.t26 4.5005
R4508 1st_Vout_1.n1 1st_Vout_1.t22 4.5005
R4509 1st_Vout_1.n1 1st_Vout_1.t11 4.5005
R4510 1st_Vout_1.n5 1st_Vout_1.t25 4.5005
R4511 1st_Vout_1.n5 1st_Vout_1.t21 4.5005
R4512 1st_Vout_1.n1 1st_Vout_1.t13 4.5005
R4513 1st_Vout_1.n1 1st_Vout_1.t29 4.5005
R4514 1st_Vout_1.n14 1st_Vout_1.n3 4.5005
R4515 1st_Vout_1.n17 1st_Vout_1.n16 4.5005
R4516 1st_Vout_1.n3 1st_Vout_1.n2 2.0005
R4517 1st_Vout_1.n2 1st_Vout_1.n11 1.813
R4518 1st_Vout_1.n1 1st_Vout_1.n0 1.5515
R4519 1st_Vout_1.n3 1st_Vout_1.n9 1.3755
R4520 1st_Vout_1.n0 1st_Vout_1.n4 1.2695
R4521 1st_Vout_1.n5 1st_Vout_1.n1 0.9875
R4522 1st_Vout_1.n16 1st_Vout_1.n14 0.78175
R4523 cap_res1.t0 cap_res1.t18 178.633
R4524 cap_res1.t6 cap_res1.t11 0.1603
R4525 cap_res1.t14 cap_res1.t10 0.1603
R4526 cap_res1.t20 cap_res1.t5 0.1603
R4527 cap_res1.t9 cap_res1.t4 0.1603
R4528 cap_res1.t15 cap_res1.t17 0.1603
R4529 cap_res1.t2 cap_res1.t16 0.1603
R4530 cap_res1.t19 cap_res1.t3 0.1603
R4531 cap_res1.t7 cap_res1.t1 0.1603
R4532 cap_res1.n1 cap_res1.t12 0.159278
R4533 cap_res1.n2 cap_res1.t8 0.159278
R4534 cap_res1.n3 cap_res1.t13 0.159278
R4535 cap_res1.n3 cap_res1.t6 0.1368
R4536 cap_res1.n3 cap_res1.t14 0.1368
R4537 cap_res1.n2 cap_res1.t20 0.1368
R4538 cap_res1.n2 cap_res1.t9 0.1368
R4539 cap_res1.n1 cap_res1.t15 0.1368
R4540 cap_res1.n1 cap_res1.t2 0.1368
R4541 cap_res1.n0 cap_res1.t19 0.1368
R4542 cap_res1.n0 cap_res1.t7 0.1368
R4543 cap_res1.t12 cap_res1.n0 0.00152174
R4544 cap_res1.t8 cap_res1.n1 0.00152174
R4545 cap_res1.t13 cap_res1.n2 0.00152174
R4546 cap_res1.t18 cap_res1.n3 0.00152174
R4547 VB3_CUR_BIAS.n2 VB3_CUR_BIAS.n1 140.077
R4548 VB3_CUR_BIAS.n2 VB3_CUR_BIAS.n0 140.077
R4549 VB3_CUR_BIAS.n4 VB3_CUR_BIAS.n3 134.577
R4550 VB3_CUR_BIAS.n3 VB3_CUR_BIAS.t2 24.0005
R4551 VB3_CUR_BIAS.n3 VB3_CUR_BIAS.t3 24.0005
R4552 VB3_CUR_BIAS.n1 VB3_CUR_BIAS.t5 24.0005
R4553 VB3_CUR_BIAS.n1 VB3_CUR_BIAS.t1 24.0005
R4554 VB3_CUR_BIAS.n0 VB3_CUR_BIAS.t4 24.0005
R4555 VB3_CUR_BIAS.n0 VB3_CUR_BIAS.t0 24.0005
R4556 VB3_CUR_BIAS.n4 VB3_CUR_BIAS.n2 4.5005
R4557 VB3_CUR_BIAS VB3_CUR_BIAS.n4 2.5005
R4558 1st_Vout_2 1st_Vout_2.t31 354.854
R4559 1st_Vout_2.n0 1st_Vout_2.t15 346.8
R4560 1st_Vout_2 1st_Vout_2.n11 339.522
R4561 1st_Vout_2.n0 1st_Vout_2.n4 339.522
R4562 1st_Vout_2.n3 1st_Vout_2.n6 335.022
R4563 1st_Vout_2.n8 1st_Vout_2.t7 275.909
R4564 1st_Vout_2.n8 1st_Vout_2.n7 227.909
R4565 1st_Vout_2.n3 1st_Vout_2.n9 222.034
R4566 1st_Vout_2.n5 1st_Vout_2.t19 184.097
R4567 1st_Vout_2.n5 1st_Vout_2.t29 184.097
R4568 1st_Vout_2.n10 1st_Vout_2.t28 184.097
R4569 1st_Vout_2.n10 1st_Vout_2.t34 184.097
R4570 1st_Vout_2.n0 1st_Vout_2.n5 166.05
R4571 1st_Vout_2 1st_Vout_2.n10 166.05
R4572 1st_Vout_2.n0 1st_Vout_2.n2 57.7228
R4573 1st_Vout_2.n9 1st_Vout_2.t3 48.0005
R4574 1st_Vout_2.n9 1st_Vout_2.t8 48.0005
R4575 1st_Vout_2.n7 1st_Vout_2.t9 48.0005
R4576 1st_Vout_2.n7 1st_Vout_2.t5 48.0005
R4577 1st_Vout_2.n6 1st_Vout_2.t4 39.4005
R4578 1st_Vout_2.n6 1st_Vout_2.t1 39.4005
R4579 1st_Vout_2.n11 1st_Vout_2.t6 39.4005
R4580 1st_Vout_2.n11 1st_Vout_2.t10 39.4005
R4581 1st_Vout_2.n4 1st_Vout_2.t0 39.4005
R4582 1st_Vout_2.n4 1st_Vout_2.t2 39.4005
R4583 1st_Vout_2 1st_Vout_2.n0 5.6255
R4584 1st_Vout_2 1st_Vout_2.n3 5.28175
R4585 1st_Vout_2.n1 1st_Vout_2.t22 4.8295
R4586 1st_Vout_2.n1 1st_Vout_2.t18 4.8295
R4587 1st_Vout_2.n1 1st_Vout_2.t27 4.8295
R4588 1st_Vout_2.n1 1st_Vout_2.t25 4.8295
R4589 1st_Vout_2.n2 1st_Vout_2.t20 4.8295
R4590 1st_Vout_2.n2 1st_Vout_2.t17 4.8295
R4591 1st_Vout_2.n2 1st_Vout_2.t36 4.8295
R4592 1st_Vout_2.n3 1st_Vout_2.n8 4.5005
R4593 1st_Vout_2.n1 1st_Vout_2.t14 4.5005
R4594 1st_Vout_2.n1 1st_Vout_2.t33 4.5005
R4595 1st_Vout_2.n1 1st_Vout_2.t26 4.5005
R4596 1st_Vout_2.n1 1st_Vout_2.t21 4.5005
R4597 1st_Vout_2.n1 1st_Vout_2.t11 4.5005
R4598 1st_Vout_2.n1 1st_Vout_2.t32 4.5005
R4599 1st_Vout_2.n2 1st_Vout_2.t13 4.5005
R4600 1st_Vout_2.n2 1st_Vout_2.t30 4.5005
R4601 1st_Vout_2.n2 1st_Vout_2.t24 4.5005
R4602 1st_Vout_2.n2 1st_Vout_2.t12 4.5005
R4603 1st_Vout_2.n2 1st_Vout_2.t35 4.5005
R4604 1st_Vout_2.n2 1st_Vout_2.t23 4.5005
R4605 1st_Vout_2.n2 1st_Vout_2.t16 4.5005
R4606 1st_Vout_2.n2 1st_Vout_2.n1 3.8075
R4607 cap_res2.t0 cap_res2.t10 188.573
R4608 cap_res2.t16 cap_res2.t1 0.1603
R4609 cap_res2.t2 cap_res2.t19 0.1603
R4610 cap_res2.t9 cap_res2.t15 0.1603
R4611 cap_res2.t18 cap_res2.t13 0.1603
R4612 cap_res2.t4 cap_res2.t8 0.1603
R4613 cap_res2.t12 cap_res2.t6 0.1603
R4614 cap_res2.t7 cap_res2.t14 0.1603
R4615 cap_res2.t17 cap_res2.t11 0.1603
R4616 cap_res2.n1 cap_res2.t3 0.159278
R4617 cap_res2.n2 cap_res2.t20 0.159278
R4618 cap_res2.n3 cap_res2.t5 0.159278
R4619 cap_res2.n3 cap_res2.t16 0.1368
R4620 cap_res2.n3 cap_res2.t2 0.1368
R4621 cap_res2.n2 cap_res2.t9 0.1368
R4622 cap_res2.n2 cap_res2.t18 0.1368
R4623 cap_res2.n1 cap_res2.t4 0.1368
R4624 cap_res2.n1 cap_res2.t12 0.1368
R4625 cap_res2.n0 cap_res2.t7 0.1368
R4626 cap_res2.n0 cap_res2.t17 0.1368
R4627 cap_res2.t3 cap_res2.n0 0.00152174
R4628 cap_res2.t20 cap_res2.n1 0.00152174
R4629 cap_res2.t5 cap_res2.n2 0.00152174
R4630 cap_res2.t10 cap_res2.n3 0.00152174
R4631 START_UP.n1 START_UP.t7 238.322
R4632 START_UP.n1 START_UP.t6 238.322
R4633 START_UP.n5 START_UP.n4 175.558
R4634 START_UP.n4 START_UP.n3 168.935
R4635 START_UP.n2 START_UP.n1 166.925
R4636 START_UP.n0 START_UP.t5 130.001
R4637 START_UP.n0 START_UP.t4 81.7084
R4638 START_UP.n2 START_UP.n0 53.0427
R4639 START_UP.n3 START_UP.t2 13.1338
R4640 START_UP.n3 START_UP.t0 13.1338
R4641 START_UP.t3 START_UP.n5 13.1338
R4642 START_UP.n5 START_UP.t1 13.1338
R4643 START_UP.n4 START_UP.n2 4.21925
R4644 V_mir2.n4 V_mir2.n0 325.473
R4645 V_mir2.n9 V_mir2.n5 325.471
R4646 V_mir2.n20 V_mir2.n19 325.471
R4647 V_mir2.n16 V_mir2.t18 310.488
R4648 V_mir2.n6 V_mir2.t22 310.488
R4649 V_mir2.n1 V_mir2.t21 310.488
R4650 V_mir2.n12 V_mir2.t3 278.312
R4651 V_mir2.n12 V_mir2.n11 228.939
R4652 V_mir2.n13 V_mir2.n10 224.439
R4653 V_mir2.n18 V_mir2.t13 184.097
R4654 V_mir2.n8 V_mir2.t11 184.097
R4655 V_mir2.n3 V_mir2.t7 184.097
R4656 V_mir2.n17 V_mir2.n16 167.094
R4657 V_mir2.n7 V_mir2.n6 167.094
R4658 V_mir2.n2 V_mir2.n1 167.094
R4659 V_mir2.n9 V_mir2.n8 152
R4660 V_mir2.n4 V_mir2.n3 152
R4661 V_mir2.n19 V_mir2.n18 152
R4662 V_mir2.n16 V_mir2.t19 120.501
R4663 V_mir2.n17 V_mir2.t5 120.501
R4664 V_mir2.n6 V_mir2.t20 120.501
R4665 V_mir2.n7 V_mir2.t15 120.501
R4666 V_mir2.n1 V_mir2.t17 120.501
R4667 V_mir2.n2 V_mir2.t9 120.501
R4668 V_mir2.n11 V_mir2.t1 48.0005
R4669 V_mir2.n11 V_mir2.t2 48.0005
R4670 V_mir2.n10 V_mir2.t4 48.0005
R4671 V_mir2.n10 V_mir2.t0 48.0005
R4672 V_mir2.n18 V_mir2.n17 40.7027
R4673 V_mir2.n8 V_mir2.n7 40.7027
R4674 V_mir2.n3 V_mir2.n2 40.7027
R4675 V_mir2.n5 V_mir2.t12 39.4005
R4676 V_mir2.n5 V_mir2.t16 39.4005
R4677 V_mir2.n0 V_mir2.t8 39.4005
R4678 V_mir2.n0 V_mir2.t10 39.4005
R4679 V_mir2.t14 V_mir2.n20 39.4005
R4680 V_mir2.n20 V_mir2.t6 39.4005
R4681 V_mir2.n15 V_mir2.n4 15.8005
R4682 V_mir2.n19 V_mir2.n15 15.8005
R4683 V_mir2.n14 V_mir2.n9 9.3005
R4684 V_mir2.n13 V_mir2.n12 5.8755
R4685 V_mir2.n15 V_mir2.n14 4.5005
R4686 V_mir2.n14 V_mir2.n13 0.78175
R4687 Vbe2.n102 Vbe2.t0 162.458
R4688 Vbe2.n117 Vbe2.n116 83.5719
R4689 Vbe2.n115 Vbe2.n9 83.5719
R4690 Vbe2.n114 Vbe2.n113 83.5719
R4691 Vbe2.n105 Vbe2.n12 83.5719
R4692 Vbe2.n97 Vbe2.n13 83.5719
R4693 Vbe2.n99 Vbe2.n98 83.5719
R4694 Vbe2.n91 Vbe2.n17 83.5719
R4695 Vbe2.n81 Vbe2.n80 83.5719
R4696 Vbe2.n79 Vbe2.n78 83.5719
R4697 Vbe2.n77 Vbe2.n76 83.5719
R4698 Vbe2.n38 Vbe2.n37 83.5719
R4699 Vbe2.n36 Vbe2.n34 83.5719
R4700 Vbe2.n44 Vbe2.n33 83.5719
R4701 Vbe2.n52 Vbe2.n51 83.5719
R4702 Vbe2.n31 Vbe2.n29 83.5719
R4703 Vbe2.n57 Vbe2.n28 83.5719
R4704 Vbe2.n65 Vbe2.n64 83.5719
R4705 Vbe2.n130 Vbe2.n0 83.5719
R4706 Vbe2.n132 Vbe2.n131 83.5719
R4707 Vbe2.n134 Vbe2.n133 83.5719
R4708 Vbe2.n116 Vbe2.n8 73.682
R4709 Vbe2.n37 Vbe2.n35 73.682
R4710 Vbe2.n114 Vbe2.n10 73.3165
R4711 Vbe2.n98 Vbe2.n96 73.3165
R4712 Vbe2.n77 Vbe2.n24 73.3165
R4713 Vbe2.n46 Vbe2.n33 73.3165
R4714 Vbe2.n59 Vbe2.n28 73.3165
R4715 Vbe2.n135 Vbe2.n134 73.3165
R4716 Vbe2.n107 Vbe2.n12 73.19
R4717 Vbe2.n93 Vbe2.n17 73.19
R4718 Vbe2.n82 Vbe2.n81 73.19
R4719 Vbe2.n51 Vbe2.n50 73.19
R4720 Vbe2.n64 Vbe2.n63 73.19
R4721 Vbe2.n130 Vbe2.n4 73.19
R4722 Vbe2.n18 Vbe2.t4 36.6632
R4723 Vbe2.t6 Vbe2.n25 36.6632
R4724 Vbe2.n115 Vbe2.n114 26.074
R4725 Vbe2.n98 Vbe2.n97 26.074
R4726 Vbe2.n79 Vbe2.n77 26.074
R4727 Vbe2.n36 Vbe2.n33 26.074
R4728 Vbe2.n31 Vbe2.n28 26.074
R4729 Vbe2.n134 Vbe2.n132 26.074
R4730 Vbe2.n116 Vbe2.t7 25.7843
R4731 Vbe2.t2 Vbe2.n12 25.7843
R4732 Vbe2.t4 Vbe2.n17 25.7843
R4733 Vbe2.n81 Vbe2.t5 25.7843
R4734 Vbe2.n37 Vbe2.t1 25.7843
R4735 Vbe2.n51 Vbe2.t3 25.7843
R4736 Vbe2.n64 Vbe2.t6 25.7843
R4737 Vbe2.t8 Vbe2.n130 25.7843
R4738 Vbe2.n138 Vbe2.n3 9.3005
R4739 Vbe2.n124 Vbe2.n3 9.3005
R4740 Vbe2.n129 Vbe2.n3 9.3005
R4741 Vbe2.n136 Vbe2.n3 9.3005
R4742 Vbe2.n138 Vbe2.n5 9.3005
R4743 Vbe2.n124 Vbe2.n5 9.3005
R4744 Vbe2.n129 Vbe2.n5 9.3005
R4745 Vbe2.n136 Vbe2.n5 9.3005
R4746 Vbe2.n138 Vbe2.n2 9.3005
R4747 Vbe2.n124 Vbe2.n2 9.3005
R4748 Vbe2.n129 Vbe2.n2 9.3005
R4749 Vbe2.n136 Vbe2.n2 9.3005
R4750 Vbe2.n138 Vbe2.n6 9.3005
R4751 Vbe2.n124 Vbe2.n6 9.3005
R4752 Vbe2.n129 Vbe2.n6 9.3005
R4753 Vbe2.n136 Vbe2.n6 9.3005
R4754 Vbe2.n138 Vbe2.n1 9.3005
R4755 Vbe2.n124 Vbe2.n1 9.3005
R4756 Vbe2.n129 Vbe2.n1 9.3005
R4757 Vbe2.n123 Vbe2.n1 9.3005
R4758 Vbe2.n136 Vbe2.n1 9.3005
R4759 Vbe2.n138 Vbe2.n137 9.3005
R4760 Vbe2.n137 Vbe2.n124 9.3005
R4761 Vbe2.n137 Vbe2.n129 9.3005
R4762 Vbe2.n137 Vbe2.n123 9.3005
R4763 Vbe2.n137 Vbe2.n136 9.3005
R4764 Vbe2.n71 Vbe2.n22 9.3005
R4765 Vbe2.n71 Vbe2.n20 9.3005
R4766 Vbe2.n71 Vbe2.n23 9.3005
R4767 Vbe2.n86 Vbe2.n71 9.3005
R4768 Vbe2.n73 Vbe2.n22 9.3005
R4769 Vbe2.n73 Vbe2.n20 9.3005
R4770 Vbe2.n73 Vbe2.n23 9.3005
R4771 Vbe2.n86 Vbe2.n73 9.3005
R4772 Vbe2.n70 Vbe2.n22 9.3005
R4773 Vbe2.n70 Vbe2.n20 9.3005
R4774 Vbe2.n70 Vbe2.n23 9.3005
R4775 Vbe2.n86 Vbe2.n70 9.3005
R4776 Vbe2.n85 Vbe2.n22 9.3005
R4777 Vbe2.n85 Vbe2.n20 9.3005
R4778 Vbe2.n85 Vbe2.n23 9.3005
R4779 Vbe2.n86 Vbe2.n85 9.3005
R4780 Vbe2.n69 Vbe2.n22 9.3005
R4781 Vbe2.n69 Vbe2.n20 9.3005
R4782 Vbe2.n69 Vbe2.n23 9.3005
R4783 Vbe2.n69 Vbe2.n19 9.3005
R4784 Vbe2.n86 Vbe2.n69 9.3005
R4785 Vbe2.n87 Vbe2.n22 9.3005
R4786 Vbe2.n87 Vbe2.n20 9.3005
R4787 Vbe2.n87 Vbe2.n23 9.3005
R4788 Vbe2.n87 Vbe2.n19 9.3005
R4789 Vbe2.n87 Vbe2.n86 9.3005
R4790 Vbe2.n123 Vbe2.n121 4.64654
R4791 Vbe2.n127 Vbe2.n126 4.64654
R4792 Vbe2.n123 Vbe2.n122 4.64654
R4793 Vbe2.n127 Vbe2.n125 4.64654
R4794 Vbe2.n128 Vbe2.n127 4.64654
R4795 Vbe2.n72 Vbe2.n19 4.64654
R4796 Vbe2.n83 Vbe2.n75 4.64654
R4797 Vbe2.n74 Vbe2.n19 4.64654
R4798 Vbe2.n84 Vbe2.n83 4.64654
R4799 Vbe2.n83 Vbe2.n21 4.64654
R4800 Vbe2.n108 Vbe2.n107 2.36206
R4801 Vbe2.n94 Vbe2.n93 2.36206
R4802 Vbe2.n50 Vbe2.n48 2.36206
R4803 Vbe2.n63 Vbe2.n61 2.36206
R4804 Vbe2.n109 Vbe2.n10 2.19742
R4805 Vbe2.n96 Vbe2.n95 2.19742
R4806 Vbe2.n47 Vbe2.n46 2.19742
R4807 Vbe2.n60 Vbe2.n59 2.19742
R4808 Vbe2.n90 Vbe2.n18 1.80777
R4809 Vbe2.n66 Vbe2.n25 1.80777
R4810 Vbe2.n62 Vbe2.n26 1.5505
R4811 Vbe2.n67 Vbe2.n66 1.5505
R4812 Vbe2.n49 Vbe2.n30 1.5505
R4813 Vbe2.n54 Vbe2.n53 1.5505
R4814 Vbe2.n56 Vbe2.n55 1.5505
R4815 Vbe2.n58 Vbe2.n27 1.5505
R4816 Vbe2.n40 Vbe2.n39 1.5505
R4817 Vbe2.n43 Vbe2.n42 1.5505
R4818 Vbe2.n45 Vbe2.n32 1.5505
R4819 Vbe2.n92 Vbe2.n16 1.5505
R4820 Vbe2.n90 Vbe2.n89 1.5505
R4821 Vbe2.n106 Vbe2.n11 1.5505
R4822 Vbe2.n104 Vbe2.n103 1.5505
R4823 Vbe2.n101 Vbe2.n100 1.5505
R4824 Vbe2.n15 Vbe2.n14 1.5505
R4825 Vbe2.n119 Vbe2.n118 1.5505
R4826 Vbe2.n112 Vbe2.n7 1.5505
R4827 Vbe2.n111 Vbe2.n110 1.5505
R4828 Vbe2.n111 Vbe2.n10 1.19225
R4829 Vbe2.n96 Vbe2.n15 1.19225
R4830 Vbe2.n24 Vbe2.n19 1.19225
R4831 Vbe2.n46 Vbe2.n45 1.19225
R4832 Vbe2.n59 Vbe2.n58 1.19225
R4833 Vbe2.n135 Vbe2.n123 1.19225
R4834 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14.Emitter Vbe2.n8 1.07742
R4835 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12.Emitter Vbe2.n35 1.07742
R4836 Vbe2.n118 Vbe2.n9 1.07024
R4837 Vbe2.n104 Vbe2.n13 1.07024
R4838 Vbe2.n78 Vbe2.n20 1.07024
R4839 Vbe2.n39 Vbe2.n34 1.07024
R4840 Vbe2.n53 Vbe2.n29 1.07024
R4841 Vbe2.n131 Vbe2.n124 1.07024
R4842 Vbe2.n68 Vbe2.n25 1.04793
R4843 Vbe2.n88 Vbe2.n18 1.04793
R4844 Vbe2.n107 Vbe2.n106 1.0237
R4845 Vbe2.n93 Vbe2.n92 1.0237
R4846 Vbe2.n82 Vbe2.n22 1.0237
R4847 Vbe2.n50 Vbe2.n49 1.0237
R4848 Vbe2.n63 Vbe2.n62 1.0237
R4849 Vbe2.n138 Vbe2.n4 1.0237
R4850 Vbe2.n113 Vbe2.n111 0.959578
R4851 Vbe2.n99 Vbe2.n15 0.959578
R4852 Vbe2.n76 Vbe2.n19 0.959578
R4853 Vbe2.n45 Vbe2.n44 0.959578
R4854 Vbe2.n58 Vbe2.n57 0.959578
R4855 Vbe2.n133 Vbe2.n123 0.959578
R4856 Vbe2.n113 Vbe2.n112 0.885803
R4857 Vbe2.n100 Vbe2.n99 0.885803
R4858 Vbe2.n76 Vbe2.n23 0.885803
R4859 Vbe2.n44 Vbe2.n43 0.885803
R4860 Vbe2.n57 Vbe2.n56 0.885803
R4861 Vbe2.n133 Vbe2.n129 0.885803
R4862 Vbe2.n83 Vbe2.n82 0.812055
R4863 Vbe2.n127 Vbe2.n4 0.812055
R4864 Vbe2.n112 Vbe2.n9 0.77514
R4865 Vbe2.n100 Vbe2.n13 0.77514
R4866 Vbe2.n78 Vbe2.n23 0.77514
R4867 Vbe2.n43 Vbe2.n34 0.77514
R4868 Vbe2.n56 Vbe2.n29 0.77514
R4869 Vbe2.n131 Vbe2.n129 0.77514
R4870 Vbe2.n40 Vbe2.n35 0.763532
R4871 Vbe2.n119 Vbe2.n8 0.763532
R4872 Vbe2.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16.Emitter 0.756696
R4873 Vbe2.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11.Emitter 0.756696
R4874 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9.Emitter Vbe2.n22 0.756696
R4875 Vbe2.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15.Emitter 0.756696
R4876 Vbe2.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10.Emitter 0.756696
R4877 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13.Emitter Vbe2.n138 0.756696
R4878 Vbe2.n86 Vbe2.n24 0.647417
R4879 Vbe2.n136 Vbe2.n135 0.647417
R4880 Vbe2.n118 Vbe2.n117 0.590702
R4881 Vbe2.n105 Vbe2.n104 0.590702
R4882 Vbe2.n91 Vbe2.n90 0.590702
R4883 Vbe2.n80 Vbe2.n20 0.590702
R4884 Vbe2.n39 Vbe2.n38 0.590702
R4885 Vbe2.n53 Vbe2.n52 0.590702
R4886 Vbe2.n66 Vbe2.n65 0.590702
R4887 Vbe2.n124 Vbe2.n0 0.590702
R4888 Vbe2.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14.Emitter 0.498483
R4889 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16.Emitter Vbe2.n105 0.498483
R4890 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11.Emitter Vbe2.n91 0.498483
R4891 Vbe2.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9.Emitter 0.498483
R4892 Vbe2.n38 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12.Emitter 0.498483
R4893 Vbe2.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15.Emitter 0.498483
R4894 Vbe2.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10.Emitter 0.498483
R4895 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13.Emitter Vbe2.n0 0.498483
R4896 Vbe2.t7 Vbe2.n115 0.290206
R4897 Vbe2.n97 Vbe2.t2 0.290206
R4898 Vbe2.t5 Vbe2.n79 0.290206
R4899 Vbe2.t1 Vbe2.n36 0.290206
R4900 Vbe2.t3 Vbe2.n31 0.290206
R4901 Vbe2.n132 Vbe2.t8 0.290206
R4902 Vbe2.n61 Vbe2.n60 0.154071
R4903 Vbe2.n48 Vbe2.n47 0.154071
R4904 Vbe2.n95 Vbe2.n94 0.154071
R4905 Vbe2.n109 Vbe2.n108 0.154071
R4906 Vbe2.n137 Vbe2.n120 0.137464
R4907 Vbe2.n88 Vbe2.n87 0.137464
R4908 Vbe2.n41 Vbe2.n1 0.134964
R4909 Vbe2.n69 Vbe2.n68 0.134964
R4910 Vbe2.n67 Vbe2.n26 0.0183571
R4911 Vbe2.n61 Vbe2.n26 0.0183571
R4912 Vbe2.n60 Vbe2.n27 0.0183571
R4913 Vbe2.n55 Vbe2.n27 0.0183571
R4914 Vbe2.n55 Vbe2.n54 0.0183571
R4915 Vbe2.n54 Vbe2.n30 0.0183571
R4916 Vbe2.n48 Vbe2.n30 0.0183571
R4917 Vbe2.n47 Vbe2.n32 0.0183571
R4918 Vbe2.n42 Vbe2.n32 0.0183571
R4919 Vbe2.n89 Vbe2.n16 0.0183571
R4920 Vbe2.n94 Vbe2.n16 0.0183571
R4921 Vbe2.n95 Vbe2.n14 0.0183571
R4922 Vbe2.n101 Vbe2.n14 0.0183571
R4923 Vbe2.n103 Vbe2.n11 0.0183571
R4924 Vbe2.n108 Vbe2.n11 0.0183571
R4925 Vbe2.n110 Vbe2.n109 0.0183571
R4926 Vbe2.n110 Vbe2.n7 0.0183571
R4927 Vbe2.n68 Vbe2.n67 0.0106786
R4928 Vbe2.n41 Vbe2.n40 0.0106786
R4929 Vbe2.n89 Vbe2.n88 0.0106786
R4930 Vbe2.n120 Vbe2.n119 0.0106786
R4931 Vbe2.n102 Vbe2.n101 0.00996429
R4932 Vbe2.n137 Vbe2.n128 0.00992001
R4933 Vbe2.n121 Vbe2.n5 0.00992001
R4934 Vbe2.n126 Vbe2.n2 0.00992001
R4935 Vbe2.n122 Vbe2.n6 0.00992001
R4936 Vbe2.n125 Vbe2.n1 0.00992001
R4937 Vbe2.n128 Vbe2.n3 0.00992001
R4938 Vbe2.n121 Vbe2.n3 0.00992001
R4939 Vbe2.n126 Vbe2.n5 0.00992001
R4940 Vbe2.n122 Vbe2.n2 0.00992001
R4941 Vbe2.n125 Vbe2.n6 0.00992001
R4942 Vbe2.n87 Vbe2.n21 0.00992001
R4943 Vbe2.n73 Vbe2.n72 0.00992001
R4944 Vbe2.n75 Vbe2.n70 0.00992001
R4945 Vbe2.n85 Vbe2.n74 0.00992001
R4946 Vbe2.n84 Vbe2.n69 0.00992001
R4947 Vbe2.n71 Vbe2.n21 0.00992001
R4948 Vbe2.n72 Vbe2.n71 0.00992001
R4949 Vbe2.n75 Vbe2.n73 0.00992001
R4950 Vbe2.n74 Vbe2.n70 0.00992001
R4951 Vbe2.n85 Vbe2.n84 0.00992001
R4952 Vbe2.n103 Vbe2.n102 0.00889286
R4953 Vbe2.n42 Vbe2.n41 0.00817857
R4954 Vbe2.n120 Vbe2.n7 0.00817857
R4955 a_4400_6480.t0 a_4400_6480.t1 376.99
R4956 NFET_GATE_10uA.n19 NFET_GATE_10uA.n0 392.666
R4957 NFET_GATE_10uA.n10 NFET_GATE_10uA.t23 273.134
R4958 NFET_GATE_10uA.n9 NFET_GATE_10uA.t6 273.134
R4959 NFET_GATE_10uA.n7 NFET_GATE_10uA.t12 273.134
R4960 NFET_GATE_10uA.n4 NFET_GATE_10uA.t11 273.134
R4961 NFET_GATE_10uA.n1 NFET_GATE_10uA.t22 273.134
R4962 NFET_GATE_10uA.t2 NFET_GATE_10uA.n18 273.134
R4963 NFET_GATE_10uA.n11 NFET_GATE_10uA.n10 224.934
R4964 NFET_GATE_10uA.n12 NFET_GATE_10uA.n11 224.934
R4965 NFET_GATE_10uA.n5 NFET_GATE_10uA.n4 224.934
R4966 NFET_GATE_10uA.n6 NFET_GATE_10uA.n5 224.934
R4967 NFET_GATE_10uA.n2 NFET_GATE_10uA.n1 224.934
R4968 NFET_GATE_10uA.n3 NFET_GATE_10uA.n2 224.934
R4969 NFET_GATE_10uA.n17 NFET_GATE_10uA.n16 224.934
R4970 NFET_GATE_10uA.n18 NFET_GATE_10uA.n17 224.934
R4971 NFET_GATE_10uA.n19 NFET_GATE_10uA.t2 200.201
R4972 NFET_GATE_10uA.n14 NFET_GATE_10uA.n13 171.582
R4973 NFET_GATE_10uA.n14 NFET_GATE_10uA.n8 171.582
R4974 NFET_GATE_10uA.n15 NFET_GATE_10uA.n14 166.113
R4975 NFET_GATE_10uA.n20 NFET_GATE_10uA.n19 150.876
R4976 NFET_GATE_10uA.n13 NFET_GATE_10uA.n12 69.6227
R4977 NFET_GATE_10uA.n13 NFET_GATE_10uA.n9 69.6227
R4978 NFET_GATE_10uA.n8 NFET_GATE_10uA.n7 69.6227
R4979 NFET_GATE_10uA.n8 NFET_GATE_10uA.n6 69.6227
R4980 NFET_GATE_10uA.n15 NFET_GATE_10uA.n3 69.6227
R4981 NFET_GATE_10uA.n16 NFET_GATE_10uA.n15 69.6227
R4982 NFET_GATE_10uA.n10 NFET_GATE_10uA.t5 48.2005
R4983 NFET_GATE_10uA.n11 NFET_GATE_10uA.t14 48.2005
R4984 NFET_GATE_10uA.n12 NFET_GATE_10uA.t15 48.2005
R4985 NFET_GATE_10uA.n9 NFET_GATE_10uA.t18 48.2005
R4986 NFET_GATE_10uA.n7 NFET_GATE_10uA.t13 48.2005
R4987 NFET_GATE_10uA.n4 NFET_GATE_10uA.t8 48.2005
R4988 NFET_GATE_10uA.n5 NFET_GATE_10uA.t7 48.2005
R4989 NFET_GATE_10uA.n6 NFET_GATE_10uA.t21 48.2005
R4990 NFET_GATE_10uA.n1 NFET_GATE_10uA.t20 48.2005
R4991 NFET_GATE_10uA.n2 NFET_GATE_10uA.t17 48.2005
R4992 NFET_GATE_10uA.n3 NFET_GATE_10uA.t10 48.2005
R4993 NFET_GATE_10uA.n16 NFET_GATE_10uA.t9 48.2005
R4994 NFET_GATE_10uA.n17 NFET_GATE_10uA.t19 48.2005
R4995 NFET_GATE_10uA.n18 NFET_GATE_10uA.t16 48.2005
R4996 NFET_GATE_10uA.n0 NFET_GATE_10uA.t1 39.4005
R4997 NFET_GATE_10uA.n0 NFET_GATE_10uA.t4 39.4005
R4998 NFET_GATE_10uA.n20 NFET_GATE_10uA.t3 24.0005
R4999 NFET_GATE_10uA.t0 NFET_GATE_10uA.n20 24.0005
R5000 VB2_CUR_BIAS.n5 VB2_CUR_BIAS.n3 141.422
R5001 VB2_CUR_BIAS.n2 VB2_CUR_BIAS.n0 141.421
R5002 VB2_CUR_BIAS.n5 VB2_CUR_BIAS.n4 139.296
R5003 VB2_CUR_BIAS.n2 VB2_CUR_BIAS.n1 139.296
R5004 VB2_CUR_BIAS.n4 VB2_CUR_BIAS.t1 24.0005
R5005 VB2_CUR_BIAS.n4 VB2_CUR_BIAS.t6 24.0005
R5006 VB2_CUR_BIAS.n3 VB2_CUR_BIAS.t2 24.0005
R5007 VB2_CUR_BIAS.n3 VB2_CUR_BIAS.t7 24.0005
R5008 VB2_CUR_BIAS.n1 VB2_CUR_BIAS.t3 24.0005
R5009 VB2_CUR_BIAS.n1 VB2_CUR_BIAS.t0 24.0005
R5010 VB2_CUR_BIAS.n0 VB2_CUR_BIAS.t4 24.0005
R5011 VB2_CUR_BIAS.n0 VB2_CUR_BIAS.t5 24.0005
R5012 VB2_CUR_BIAS VB2_CUR_BIAS.n6 6.8755
R5013 VB2_CUR_BIAS.n6 VB2_CUR_BIAS.n5 4.34425
R5014 VB2_CUR_BIAS.n6 VB2_CUR_BIAS.n2 4.34425
R5015 a_2792_6360.t0 a_2792_6360.t1 258.591
R5016 START_UP_NFET1.t0 START_UP_NFET1.t1 178.194
R5017 Vin-.n11 Vin-.t10 688.859
R5018 Vin-.n13 Vin-.n12 514.134
R5019 Vin-.n9 Vin-.n8 345.116
R5020 Vin-.n15 Vin-.n14 214.713
R5021 Vin-.n11 Vin-.t8 174.726
R5022 Vin-.n12 Vin-.t12 174.726
R5023 Vin-.n13 Vin-.t11 174.726
R5024 Vin-.n14 Vin-.t9 174.726
R5025 Vin-.n7 Vin-.n5 173.029
R5026 Vin-.n7 Vin-.n6 168.654
R5027 Vin-.n9 Vin-.t0 162.921
R5028 Vin-.n12 Vin-.n11 128.534
R5029 Vin-.n14 Vin-.n13 128.534
R5030 Vin-.n1 Vin-.n0 83.5719
R5031 Vin-.n22 Vin-.n21 83.5719
R5032 Vin-.n20 Vin-.n19 83.5719
R5033 Vin-.n25 Vin-.n1 73.682
R5034 Vin-.n20 Vin-.n4 73.3165
R5035 Vin-.n8 Vin-.t7 39.4005
R5036 Vin-.n8 Vin-.t6 39.4005
R5037 Vin-.n21 Vin-.n20 26.074
R5038 Vin-.t5 Vin-.n1 25.7843
R5039 Vin-.n16 Vin-.n15 17.526
R5040 Vin-.n6 Vin-.t1 13.1338
R5041 Vin-.n6 Vin-.t2 13.1338
R5042 Vin-.n5 Vin-.t3 13.1338
R5043 Vin-.n5 Vin-.t4 13.1338
R5044 Vin-.n15 Vin-.n10 12.5317
R5045 Vin-.n10 Vin-.n9 6.40675
R5046 Vin-.n10 Vin-.n7 3.8755
R5047 Vin-.n16 Vin-.n4 2.19742
R5048 Vin-.n24 Vin-.n23 1.5505
R5049 Vin-.n3 Vin-.n2 1.5505
R5050 Vin-.n18 Vin-.n17 1.5505
R5051 Vin-.n18 Vin-.n4 1.19225
R5052 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter Vin-.n25 1.07742
R5053 Vin-.n23 Vin-.n22 1.07024
R5054 Vin-.n19 Vin-.n18 0.959578
R5055 Vin-.n19 Vin-.n3 0.885803
R5056 Vin-.n22 Vin-.n3 0.77514
R5057 Vin-.n25 Vin-.n24 0.763532
R5058 Vin-.n23 Vin-.n0 0.590702
R5059 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter Vin-.n0 0.498483
R5060 Vin-.n21 Vin-.t5 0.290206
R5061 Vin-.n17 Vin-.n16 0.0183571
R5062 Vin-.n17 Vin-.n2 0.0183571
R5063 Vin-.n24 Vin-.n2 0.0183571
R5064 VB1_CUR_BIAS.n2 VB1_CUR_BIAS.n0 340.397
R5065 VB1_CUR_BIAS.n2 VB1_CUR_BIAS.n1 339.272
R5066 VB1_CUR_BIAS.n1 VB1_CUR_BIAS.t3 39.4005
R5067 VB1_CUR_BIAS.n1 VB1_CUR_BIAS.t1 39.4005
R5068 VB1_CUR_BIAS.n0 VB1_CUR_BIAS.t0 39.4005
R5069 VB1_CUR_BIAS.n0 VB1_CUR_BIAS.t2 39.4005
R5070 VB1_CUR_BIAS VB1_CUR_BIAS.n2 3.813
R5071 V_CUR_REF_REG.n3 V_CUR_REF_REG.n2 526.183
R5072 V_CUR_REF_REG.n1 V_CUR_REF_REG.n0 514.134
R5073 V_CUR_REF_REG.n0 V_CUR_REF_REG.t5 303.259
R5074 V_CUR_REF_REG.n5 V_CUR_REF_REG.n4 287.264
R5075 V_CUR_REF_REG.n5 V_CUR_REF_REG.n3 282.522
R5076 V_CUR_REF_REG.t0 V_CUR_REF_REG.n5 244.567
R5077 V_CUR_REF_REG.n0 V_CUR_REF_REG.t7 174.726
R5078 V_CUR_REF_REG.n1 V_CUR_REF_REG.t3 174.726
R5079 V_CUR_REF_REG.n2 V_CUR_REF_REG.t4 174.726
R5080 V_CUR_REF_REG.n2 V_CUR_REF_REG.n1 128.534
R5081 V_CUR_REF_REG.n3 V_CUR_REF_REG.t6 96.4005
R5082 V_CUR_REF_REG.n4 V_CUR_REF_REG.t2 39.4005
R5083 V_CUR_REF_REG.n4 V_CUR_REF_REG.t1 39.4005
R5084 V_p_2.n1 V_p_2.n4 229.562
R5085 V_p_2.n1 V_p_2.n5 228.939
R5086 V_p_2.n0 V_p_2.n3 228.939
R5087 V_p_2.n0 V_p_2.n2 228.939
R5088 V_p_2.n6 V_p_2.n0 228.938
R5089 V_p_2.n0 V_p_2.t10 98.2282
R5090 V_p_2.n5 V_p_2.t2 48.0005
R5091 V_p_2.n5 V_p_2.t5 48.0005
R5092 V_p_2.n4 V_p_2.t7 48.0005
R5093 V_p_2.n4 V_p_2.t3 48.0005
R5094 V_p_2.n3 V_p_2.t0 48.0005
R5095 V_p_2.n3 V_p_2.t8 48.0005
R5096 V_p_2.n2 V_p_2.t6 48.0005
R5097 V_p_2.n2 V_p_2.t4 48.0005
R5098 V_p_2.t9 V_p_2.n6 48.0005
R5099 V_p_2.n6 V_p_2.t1 48.0005
R5100 V_p_2.n0 V_p_2.n1 1.8755
R5101 ERR_AMP_REF.n0 ERR_AMP_REF.t8 688.859
R5102 ERR_AMP_REF.n2 ERR_AMP_REF.n1 514.134
R5103 ERR_AMP_REF.n10 ERR_AMP_REF.n3 208.838
R5104 ERR_AMP_REF.n5 ERR_AMP_REF.t0 197.964
R5105 ERR_AMP_REF.n0 ERR_AMP_REF.t10 174.726
R5106 ERR_AMP_REF.n1 ERR_AMP_REF.t11 174.726
R5107 ERR_AMP_REF.n2 ERR_AMP_REF.t7 174.726
R5108 ERR_AMP_REF.n3 ERR_AMP_REF.t9 174.726
R5109 ERR_AMP_REF.n9 ERR_AMP_REF.n8 169.215
R5110 ERR_AMP_REF.n7 ERR_AMP_REF.n6 169.215
R5111 ERR_AMP_REF.n5 ERR_AMP_REF.n4 169.215
R5112 ERR_AMP_REF.n1 ERR_AMP_REF.n0 128.534
R5113 ERR_AMP_REF.n3 ERR_AMP_REF.n2 128.534
R5114 ERR_AMP_REF.n10 ERR_AMP_REF.n9 16.8443
R5115 ERR_AMP_REF.n8 ERR_AMP_REF.t6 13.1338
R5116 ERR_AMP_REF.n8 ERR_AMP_REF.t4 13.1338
R5117 ERR_AMP_REF.n6 ERR_AMP_REF.t2 13.1338
R5118 ERR_AMP_REF.n6 ERR_AMP_REF.t3 13.1338
R5119 ERR_AMP_REF.n4 ERR_AMP_REF.t1 13.1338
R5120 ERR_AMP_REF.n4 ERR_AMP_REF.t5 13.1338
R5121 ERR_AMP_REF.n7 ERR_AMP_REF.n5 4.3755
R5122 ERR_AMP_REF.n9 ERR_AMP_REF.n7 4.3755
R5123 ERR_AMP_REF ERR_AMP_REF.n10 3.1255
R5124 V_mir1.n20 V_mir1.n19 325.473
R5125 V_mir1.n9 V_mir1.n5 325.471
R5126 V_mir1.n4 V_mir1.n0 325.471
R5127 V_mir1.n16 V_mir1.t17 310.488
R5128 V_mir1.n6 V_mir1.t19 310.488
R5129 V_mir1.n1 V_mir1.t20 310.488
R5130 V_mir1.n12 V_mir1.t14 278.312
R5131 V_mir1.n12 V_mir1.n11 228.939
R5132 V_mir1.n13 V_mir1.n10 224.439
R5133 V_mir1.n18 V_mir1.t10 184.097
R5134 V_mir1.n8 V_mir1.t8 184.097
R5135 V_mir1.n3 V_mir1.t6 184.097
R5136 V_mir1.n17 V_mir1.n16 167.094
R5137 V_mir1.n7 V_mir1.n6 167.094
R5138 V_mir1.n2 V_mir1.n1 167.094
R5139 V_mir1.n9 V_mir1.n8 152
R5140 V_mir1.n4 V_mir1.n3 152
R5141 V_mir1.n19 V_mir1.n18 152
R5142 V_mir1.n16 V_mir1.t21 120.501
R5143 V_mir1.n17 V_mir1.t4 120.501
R5144 V_mir1.n6 V_mir1.t22 120.501
R5145 V_mir1.n7 V_mir1.t2 120.501
R5146 V_mir1.n1 V_mir1.t18 120.501
R5147 V_mir1.n2 V_mir1.t0 120.501
R5148 V_mir1.n11 V_mir1.t16 48.0005
R5149 V_mir1.n11 V_mir1.t12 48.0005
R5150 V_mir1.n10 V_mir1.t13 48.0005
R5151 V_mir1.n10 V_mir1.t15 48.0005
R5152 V_mir1.n18 V_mir1.n17 40.7027
R5153 V_mir1.n8 V_mir1.n7 40.7027
R5154 V_mir1.n3 V_mir1.n2 40.7027
R5155 V_mir1.n5 V_mir1.t3 39.4005
R5156 V_mir1.n5 V_mir1.t9 39.4005
R5157 V_mir1.n0 V_mir1.t1 39.4005
R5158 V_mir1.n0 V_mir1.t7 39.4005
R5159 V_mir1.n20 V_mir1.t5 39.4005
R5160 V_mir1.t11 V_mir1.n20 39.4005
R5161 V_mir1.n15 V_mir1.n4 15.8005
R5162 V_mir1.n19 V_mir1.n15 15.8005
R5163 V_mir1.n14 V_mir1.n9 9.3005
R5164 V_mir1.n13 V_mir1.n12 5.8755
R5165 V_mir1.n15 V_mir1.n14 4.5005
R5166 V_mir1.n14 V_mir1.n13 0.78175
R5167 V_CMFB_S4.n2 V_CMFB_S4.n0 145.702
R5168 V_CMFB_S4.n2 V_CMFB_S4.n1 134.577
R5169 V_CMFB_S4.n1 V_CMFB_S4.t0 24.0005
R5170 V_CMFB_S4.n1 V_CMFB_S4.t3 24.0005
R5171 V_CMFB_S4.n0 V_CMFB_S4.t1 24.0005
R5172 V_CMFB_S4.n0 V_CMFB_S4.t2 24.0005
R5173 V_CMFB_S4 V_CMFB_S4.n2 2.71925
R5174 V_CMFB_S3.n2 V_CMFB_S3.n0 340.272
R5175 V_CMFB_S3.n4 V_CMFB_S3.n3 339.272
R5176 V_CMFB_S3.n2 V_CMFB_S3.n1 339.272
R5177 V_CMFB_S3.n3 V_CMFB_S3.t5 39.4005
R5178 V_CMFB_S3.n3 V_CMFB_S3.t0 39.4005
R5179 V_CMFB_S3.n1 V_CMFB_S3.t1 39.4005
R5180 V_CMFB_S3.n1 V_CMFB_S3.t2 39.4005
R5181 V_CMFB_S3.n0 V_CMFB_S3.t3 39.4005
R5182 V_CMFB_S3.n0 V_CMFB_S3.t4 39.4005
R5183 V_CMFB_S3 V_CMFB_S3.n4 4.438
R5184 V_CMFB_S3.n4 V_CMFB_S3.n2 1.0005
R5185 a_1830_6460.t0 a_1830_6460.t1 258.591
R5186 V_CMFB_S2.n2 V_CMFB_S2.n0 145.702
R5187 V_CMFB_S2.n2 V_CMFB_S2.n1 134.577
R5188 V_CMFB_S2.n1 V_CMFB_S2.t1 24.0005
R5189 V_CMFB_S2.n1 V_CMFB_S2.t0 24.0005
R5190 V_CMFB_S2.n0 V_CMFB_S2.t2 24.0005
R5191 V_CMFB_S2.n0 V_CMFB_S2.t3 24.0005
R5192 V_CMFB_S2 V_CMFB_S2.n2 2.71925
R5193 ERR_AMP_CUR_BIAS ERR_AMP_CUR_BIAS.n0 137.077
R5194 ERR_AMP_CUR_BIAS.n0 ERR_AMP_CUR_BIAS.t0 24.0005
R5195 ERR_AMP_CUR_BIAS.n0 ERR_AMP_CUR_BIAS.t1 24.0005
R5196 a_1890_6990.t0 a_1890_6990.t1 258.591
R5197 a_2792_6240.t0 a_2792_6240.t1 376.99
R5198 a_4400_6600.t0 a_4400_6600.t1 258.591
C0 VDDA VB2_CUR_BIAS 0.039226f
C1 ERR_AMP_REF 1st_Vout_2 1.2502f
C2 1st_Vout_2 m2_8800_4340# 0.075543f
C3 V_TOP m2_7440_4340# 0.012f
C4 V_CMFB_S1 1st_Vout_2 0.152732f
C5 VDDA ERR_AMP_REF 1.92277f
C6 ERR_AMP_REF VB1_CUR_BIAS 0.030389f
C7 V_CMFB_S1 V_CMFB_S3 0.054662f
C8 VDDA m2_8800_4340# 0.010446f
C9 1st_Vout_2 V_CMFB_S3 0.046453f
C10 TAIL_CUR_MIR_BIAS 1st_Vout_2 0.030187f
C11 VDDA V_CMFB_S1 1.56408f
C12 TAIL_CUR_MIR_BIAS V_CMFB_S3 0.09066f
C13 VDDA 1st_Vout_2 2.88327f
C14 1st_Vout_2 VB1_CUR_BIAS 0.11484f
C15 VDDA VB3_CUR_BIAS 0.014806f
C16 VDDA V_CMFB_S3 1.00211f
C17 VDDA TAIL_CUR_MIR_BIAS 2.67038f
C18 TAIL_CUR_MIR_BIAS VB1_CUR_BIAS 0.047171f
C19 ERR_AMP_CUR_BIAS VB2_CUR_BIAS 0.151486f
C20 VDDA VB1_CUR_BIAS 0.713685f
C21 V_CMFB_S4 VB2_CUR_BIAS 0.31039f
C22 VDDA li_8890_7630# 0.02401f
C23 V_TOP li_10290_7530# 0.019775f
C24 V_CMFB_S2 VB2_CUR_BIAS 0.31039f
C25 ERR_AMP_REF V_TOP 1.14179f
C26 VDDA m2_7440_4340# 0.010446f
C27 ERR_AMP_CUR_BIAS VB3_CUR_BIAS 0.023067f
C28 V_CMFB_S1 V_TOP 0.168893f
C29 V_TOP 1st_Vout_2 1.35794f
C30 V_TOP V_CMFB_S3 0.023065f
C31 VDDA ERR_AMP_CUR_BIAS 0.013734f
C32 TAIL_CUR_MIR_BIAS V_TOP 0.033074f
C33 VDDA V_CMFB_S4 0.021014f
C34 VDDA V_TOP 15.985599f
C35 VB3_CUR_BIAS VB2_CUR_BIAS 0.531334f
C36 VDDA V_CMFB_S2 0.017706f
C37 1st_Vout_2 li_6790_7420# 0.020658f
C38 ERR_AMP_REF V_CMFB_S1 0.019012f
C39 V_CMFB_S4 GNDA 1.08175f
C40 VB3_CUR_BIAS GNDA 1.07445f
C41 ERR_AMP_CUR_BIAS GNDA 0.46336f
C42 VB2_CUR_BIAS GNDA 2.64778f
C43 V_CMFB_S2 GNDA 0.970371f
C44 VB1_CUR_BIAS GNDA 0.335187f
C45 V_CMFB_S3 GNDA 0.320585f
C46 TAIL_CUR_MIR_BIAS GNDA 1.084837f
C47 V_CMFB_S1 GNDA 1.834906f
C48 ERR_AMP_REF GNDA 4.434041f
C49 VDDA GNDA 90.56943f
C50 li_6790_7420# GNDA 0.048841f $ **FLOATING
C51 li_5390_7420# GNDA 0.043891f $ **FLOATING
C52 li_10290_7530# GNDA 0.047034f $ **FLOATING
C53 li_3290_7530# GNDA 0.049721f $ **FLOATING
C54 li_1890_7530# GNDA 0.050514f $ **FLOATING
C55 li_8890_7630# GNDA 0.047886f $ **FLOATING
C56 1st_Vout_2 GNDA 5.057145f
C57 V_TOP GNDA 6.756155f
C58 V_mir1.t5 GNDA 0.03537f
C59 V_mir1.t1 GNDA 0.03537f
C60 V_mir1.t7 GNDA 0.03537f
C61 V_mir1.n0 GNDA 0.08097f
C62 V_mir1.t0 GNDA 0.042444f
C63 V_mir1.t18 GNDA 0.042444f
C64 V_mir1.t20 GNDA 0.06851f
C65 V_mir1.n1 GNDA 0.076506f
C66 V_mir1.n2 GNDA 0.052264f
C67 V_mir1.t6 GNDA 0.053881f
C68 V_mir1.n3 GNDA 0.081315f
C69 V_mir1.n4 GNDA 0.201563f
C70 V_mir1.t3 GNDA 0.03537f
C71 V_mir1.t9 GNDA 0.03537f
C72 V_mir1.n5 GNDA 0.08097f
C73 V_mir1.t2 GNDA 0.042444f
C74 V_mir1.t22 GNDA 0.042444f
C75 V_mir1.t19 GNDA 0.06851f
C76 V_mir1.n6 GNDA 0.076506f
C77 V_mir1.n7 GNDA 0.052264f
C78 V_mir1.t8 GNDA 0.053881f
C79 V_mir1.n8 GNDA 0.081315f
C80 V_mir1.n9 GNDA 0.156007f
C81 V_mir1.t13 GNDA 0.017685f
C82 V_mir1.t15 GNDA 0.017685f
C83 V_mir1.n10 GNDA 0.046242f
C84 V_mir1.t14 GNDA 0.075466f
C85 V_mir1.t16 GNDA 0.017685f
C86 V_mir1.t12 GNDA 0.017685f
C87 V_mir1.n11 GNDA 0.050199f
C88 V_mir1.n12 GNDA 0.827814f
C89 V_mir1.n13 GNDA 0.268286f
C90 V_mir1.n14 GNDA 0.09373f
C91 V_mir1.n15 GNDA 0.699157f
C92 V_mir1.t4 GNDA 0.042444f
C93 V_mir1.t21 GNDA 0.042444f
C94 V_mir1.t17 GNDA 0.06851f
C95 V_mir1.n16 GNDA 0.076506f
C96 V_mir1.n17 GNDA 0.052264f
C97 V_mir1.t10 GNDA 0.053881f
C98 V_mir1.n18 GNDA 0.081315f
C99 V_mir1.n19 GNDA 0.203577f
C100 V_mir1.n20 GNDA 0.08097f
C101 V_mir1.t11 GNDA 0.03537f
C102 ERR_AMP_REF.t8 GNDA 0.055552f
C103 ERR_AMP_REF.t10 GNDA 0.020773f
C104 ERR_AMP_REF.n0 GNDA 0.065156f
C105 ERR_AMP_REF.t11 GNDA 0.020773f
C106 ERR_AMP_REF.n1 GNDA 0.053336f
C107 ERR_AMP_REF.t7 GNDA 0.020773f
C108 ERR_AMP_REF.n2 GNDA 0.053336f
C109 ERR_AMP_REF.t9 GNDA 0.020773f
C110 ERR_AMP_REF.n3 GNDA 0.081827f
C111 ERR_AMP_REF.t0 GNDA 0.530484f
C112 ERR_AMP_REF.t1 GNDA 0.067372f
C113 ERR_AMP_REF.t5 GNDA 0.067372f
C114 ERR_AMP_REF.n4 GNDA 0.225764f
C115 ERR_AMP_REF.n5 GNDA 2.54385f
C116 ERR_AMP_REF.t2 GNDA 0.067372f
C117 ERR_AMP_REF.t3 GNDA 0.067372f
C118 ERR_AMP_REF.n6 GNDA 0.225764f
C119 ERR_AMP_REF.n7 GNDA 0.609647f
C120 ERR_AMP_REF.t6 GNDA 0.067372f
C121 ERR_AMP_REF.t4 GNDA 0.067372f
C122 ERR_AMP_REF.n8 GNDA 0.225764f
C123 ERR_AMP_REF.n9 GNDA 0.871595f
C124 ERR_AMP_REF.n10 GNDA 0.758181f
C125 V_CUR_REF_REG.t5 GNDA 0.014159f
C126 V_CUR_REF_REG.n0 GNDA 0.030368f
C127 V_CUR_REF_REG.n1 GNDA 0.023632f
C128 V_CUR_REF_REG.n2 GNDA 0.023951f
C129 V_CUR_REF_REG.n3 GNDA 0.219126f
C130 V_CUR_REF_REG.n4 GNDA 0.0199f
C131 V_CUR_REF_REG.n5 GNDA 1.48046f
C132 V_CUR_REF_REG.t0 GNDA 0.434924f
C133 Vin-.n0 GNDA 0.048818f
C134 Vin-.n1 GNDA 0.333648f
C135 Vin-.n2 GNDA 0.166915f
C136 Vin-.n3 GNDA 0.074468f
C137 Vin-.n4 GNDA 0.338979f
C138 Vin-.t3 GNDA 0.028614f
C139 Vin-.t4 GNDA 0.028614f
C140 Vin-.n5 GNDA 0.099613f
C141 Vin-.t1 GNDA 0.028614f
C142 Vin-.t2 GNDA 0.028614f
C143 Vin-.n6 GNDA 0.095121f
C144 Vin-.n7 GNDA 0.408067f
C145 Vin-.t0 GNDA 0.098662f
C146 Vin-.n8 GNDA 0.025702f
C147 Vin-.n9 GNDA 0.469862f
C148 Vin-.n10 GNDA 0.222852f
C149 Vin-.t10 GNDA 0.023594f
C150 Vin-.n11 GNDA 0.027673f
C151 Vin-.n12 GNDA 0.022653f
C152 Vin-.n13 GNDA 0.022653f
C153 Vin-.n14 GNDA 0.040466f
C154 Vin-.n15 GNDA 0.524007f
C155 Vin-.n16 GNDA 0.461299f
C156 Vin-.n17 GNDA 0.166915f
C157 Vin-.n18 GNDA 0.10855f
C158 Vin-.n19 GNDA 0.082742f
C159 Vin-.n20 GNDA 0.331333f
C160 Vin-.t5 GNDA 0.072966f
C161 Vin-.n21 GNDA 0.073776f
C162 Vin-.n22 GNDA 0.082742f
C163 Vin-.n23 GNDA 0.074468f
C164 Vin-.n24 GNDA 0.656866f
C165 Vin-.n25 GNDA 0.389111f
C166 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.086659f
C167 V_mir2.t6 GNDA 0.03537f
C168 V_mir2.t8 GNDA 0.03537f
C169 V_mir2.t10 GNDA 0.03537f
C170 V_mir2.n0 GNDA 0.08097f
C171 V_mir2.t7 GNDA 0.053881f
C172 V_mir2.t9 GNDA 0.042444f
C173 V_mir2.t17 GNDA 0.042444f
C174 V_mir2.t21 GNDA 0.06851f
C175 V_mir2.n1 GNDA 0.076506f
C176 V_mir2.n2 GNDA 0.052264f
C177 V_mir2.n3 GNDA 0.081315f
C178 V_mir2.n4 GNDA 0.201563f
C179 V_mir2.t12 GNDA 0.03537f
C180 V_mir2.t16 GNDA 0.03537f
C181 V_mir2.n5 GNDA 0.08097f
C182 V_mir2.t11 GNDA 0.053881f
C183 V_mir2.t15 GNDA 0.042444f
C184 V_mir2.t20 GNDA 0.042444f
C185 V_mir2.t22 GNDA 0.06851f
C186 V_mir2.n6 GNDA 0.076506f
C187 V_mir2.n7 GNDA 0.052264f
C188 V_mir2.n8 GNDA 0.081315f
C189 V_mir2.n9 GNDA 0.156007f
C190 V_mir2.t4 GNDA 0.017685f
C191 V_mir2.t0 GNDA 0.017685f
C192 V_mir2.n10 GNDA 0.046242f
C193 V_mir2.t3 GNDA 0.075466f
C194 V_mir2.t1 GNDA 0.017685f
C195 V_mir2.t2 GNDA 0.017685f
C196 V_mir2.n11 GNDA 0.050199f
C197 V_mir2.n12 GNDA 0.827814f
C198 V_mir2.n13 GNDA 0.268286f
C199 V_mir2.n14 GNDA 0.09373f
C200 V_mir2.n15 GNDA 0.699157f
C201 V_mir2.t13 GNDA 0.053881f
C202 V_mir2.t5 GNDA 0.042444f
C203 V_mir2.t19 GNDA 0.042444f
C204 V_mir2.t18 GNDA 0.06851f
C205 V_mir2.n16 GNDA 0.076506f
C206 V_mir2.n17 GNDA 0.052264f
C207 V_mir2.n18 GNDA 0.081315f
C208 V_mir2.n19 GNDA 0.203577f
C209 V_mir2.n20 GNDA 0.08097f
C210 V_mir2.t14 GNDA 0.03537f
C211 START_UP.t1 GNDA 0.041701f
C212 START_UP.t4 GNDA 1.6623f
C213 START_UP.t5 GNDA 0.043697f
C214 START_UP.n0 GNDA 1.28651f
C215 START_UP.t6 GNDA 0.01567f
C216 START_UP.t7 GNDA 0.01567f
C217 START_UP.n1 GNDA 0.044238f
C218 START_UP.n2 GNDA 0.853868f
C219 START_UP.t2 GNDA 0.041701f
C220 START_UP.t0 GNDA 0.041701f
C221 START_UP.n3 GNDA 0.139173f
C222 START_UP.n4 GNDA 0.720786f
C223 START_UP.n5 GNDA 0.151283f
C224 START_UP.t3 GNDA 0.041701f
C225 cap_res2.t19 GNDA 0.406156f
C226 cap_res2.t2 GNDA 0.407628f
C227 cap_res2.t1 GNDA 0.406156f
C228 cap_res2.t16 GNDA 0.407628f
C229 cap_res2.t13 GNDA 0.406156f
C230 cap_res2.t18 GNDA 0.407628f
C231 cap_res2.t15 GNDA 0.406156f
C232 cap_res2.t9 GNDA 0.407628f
C233 cap_res2.t6 GNDA 0.406156f
C234 cap_res2.t12 GNDA 0.407628f
C235 cap_res2.t8 GNDA 0.406156f
C236 cap_res2.t4 GNDA 0.407628f
C237 cap_res2.t11 GNDA 0.406156f
C238 cap_res2.t17 GNDA 0.407628f
C239 cap_res2.t14 GNDA 0.406156f
C240 cap_res2.t7 GNDA 0.407628f
C241 cap_res2.n0 GNDA 0.272247f
C242 cap_res2.t3 GNDA 0.216805f
C243 cap_res2.n1 GNDA 0.295394f
C244 cap_res2.t20 GNDA 0.216805f
C245 cap_res2.n2 GNDA 0.295394f
C246 cap_res2.t5 GNDA 0.216805f
C247 cap_res2.n3 GNDA 0.295394f
C248 cap_res2.t10 GNDA 0.846971f
C249 cap_res2.t0 GNDA 0.133907f
C250 1st_Vout_2.n0 GNDA 0.708804f
C251 1st_Vout_2.n1 GNDA 1.48853f
C252 1st_Vout_2.n2 GNDA 2.06173f
C253 1st_Vout_2.n3 GNDA 0.130779f
C254 1st_Vout_2.t12 GNDA 0.36135f
C255 1st_Vout_2.t22 GNDA 0.367505f
C256 1st_Vout_2.t14 GNDA 0.36135f
C257 1st_Vout_2.t33 GNDA 0.36135f
C258 1st_Vout_2.t18 GNDA 0.367505f
C259 1st_Vout_2.t26 GNDA 0.36135f
C260 1st_Vout_2.t27 GNDA 0.367505f
C261 1st_Vout_2.t21 GNDA 0.36135f
C262 1st_Vout_2.t11 GNDA 0.36135f
C263 1st_Vout_2.t25 GNDA 0.367505f
C264 1st_Vout_2.t32 GNDA 0.36135f
C265 1st_Vout_2.t20 GNDA 0.367505f
C266 1st_Vout_2.t13 GNDA 0.36135f
C267 1st_Vout_2.t30 GNDA 0.36135f
C268 1st_Vout_2.t17 GNDA 0.367505f
C269 1st_Vout_2.t24 GNDA 0.36135f
C270 1st_Vout_2.t36 GNDA 0.367505f
C271 1st_Vout_2.t16 GNDA 0.36135f
C272 1st_Vout_2.t23 GNDA 0.36135f
C273 1st_Vout_2.t35 GNDA 0.36135f
C274 1st_Vout_2.t15 GNDA 0.023606f
C275 1st_Vout_2.n4 GNDA 0.022772f
C276 1st_Vout_2.t29 GNDA 0.013762f
C277 1st_Vout_2.t19 GNDA 0.013762f
C278 1st_Vout_2.n5 GNDA 0.030615f
C279 1st_Vout_2.n6 GNDA 0.021829f
C280 1st_Vout_2.t7 GNDA 0.019027f
C281 1st_Vout_2.n7 GNDA 0.013049f
C282 1st_Vout_2.n8 GNDA 0.197381f
C283 1st_Vout_2.n9 GNDA 0.011807f
C284 1st_Vout_2.t34 GNDA 0.013762f
C285 1st_Vout_2.t28 GNDA 0.013762f
C286 1st_Vout_2.n10 GNDA 0.030615f
C287 1st_Vout_2.n11 GNDA 0.022772f
C288 1st_Vout_2.t31 GNDA 0.0216f
C289 cap_res1.t10 GNDA 0.417173f
C290 cap_res1.t14 GNDA 0.418684f
C291 cap_res1.t11 GNDA 0.417173f
C292 cap_res1.t6 GNDA 0.418684f
C293 cap_res1.t4 GNDA 0.417173f
C294 cap_res1.t9 GNDA 0.418684f
C295 cap_res1.t5 GNDA 0.417173f
C296 cap_res1.t20 GNDA 0.418684f
C297 cap_res1.t16 GNDA 0.417173f
C298 cap_res1.t2 GNDA 0.418684f
C299 cap_res1.t17 GNDA 0.417173f
C300 cap_res1.t15 GNDA 0.418684f
C301 cap_res1.t1 GNDA 0.417173f
C302 cap_res1.t7 GNDA 0.418684f
C303 cap_res1.t3 GNDA 0.417173f
C304 cap_res1.t19 GNDA 0.418684f
C305 cap_res1.n0 GNDA 0.279631f
C306 cap_res1.t12 GNDA 0.222685f
C307 cap_res1.n1 GNDA 0.303406f
C308 cap_res1.t8 GNDA 0.222685f
C309 cap_res1.n2 GNDA 0.303406f
C310 cap_res1.t13 GNDA 0.222685f
C311 cap_res1.n3 GNDA 0.303406f
C312 cap_res1.t18 GNDA 0.649059f
C313 cap_res1.t0 GNDA 0.10618f
C314 1st_Vout_1.n0 GNDA 1.19655f
C315 1st_Vout_1.n1 GNDA 1.19655f
C316 1st_Vout_1.n2 GNDA 0.184254f
C317 1st_Vout_1.n3 GNDA 0.119384f
C318 1st_Vout_1.n4 GNDA 0.23261f
C319 1st_Vout_1.n5 GNDA 0.588341f
C320 1st_Vout_1.n6 GNDA 0.012529f
C321 1st_Vout_1.n7 GNDA 0.020958f
C322 1st_Vout_1.t32 GNDA 0.020816f
C323 1st_Vout_1.n8 GNDA 0.021864f
C324 1st_Vout_1.n9 GNDA 0.166349f
C325 1st_Vout_1.t20 GNDA 0.013213f
C326 1st_Vout_1.t30 GNDA 0.013213f
C327 1st_Vout_1.n10 GNDA 0.029393f
C328 1st_Vout_1.t25 GNDA 0.346936f
C329 1st_Vout_1.t36 GNDA 0.352846f
C330 1st_Vout_1.t28 GNDA 0.346936f
C331 1st_Vout_1.t23 GNDA 0.346936f
C332 1st_Vout_1.t34 GNDA 0.352846f
C333 1st_Vout_1.t12 GNDA 0.346936f
C334 1st_Vout_1.t16 GNDA 0.352846f
C335 1st_Vout_1.t35 GNDA 0.346936f
C336 1st_Vout_1.t27 GNDA 0.346936f
C337 1st_Vout_1.t15 GNDA 0.352846f
C338 1st_Vout_1.t19 GNDA 0.346936f
C339 1st_Vout_1.t33 GNDA 0.352846f
C340 1st_Vout_1.t26 GNDA 0.346936f
C341 1st_Vout_1.t22 GNDA 0.346936f
C342 1st_Vout_1.t31 GNDA 0.352846f
C343 1st_Vout_1.t11 GNDA 0.346936f
C344 1st_Vout_1.t24 GNDA 0.352846f
C345 1st_Vout_1.t29 GNDA 0.346936f
C346 1st_Vout_1.t13 GNDA 0.346936f
C347 1st_Vout_1.t21 GNDA 0.346936f
C348 1st_Vout_1.t17 GNDA 0.022665f
C349 1st_Vout_1.n11 GNDA 0.389472f
C350 1st_Vout_1.n12 GNDA 0.021864f
C351 1st_Vout_1.t18 GNDA 0.013213f
C352 1st_Vout_1.t14 GNDA 0.013213f
C353 1st_Vout_1.n13 GNDA 0.029393f
C354 1st_Vout_1.n14 GNDA 0.077485f
C355 1st_Vout_1.n15 GNDA 0.011336f
C356 1st_Vout_1.n16 GNDA 0.048077f
C357 1st_Vout_1.n17 GNDA 0.189508f
C358 1st_Vout_1.t10 GNDA 0.018268f
C359 TAIL_CUR_MIR_BIAS.t0 GNDA 0.027636f
C360 TAIL_CUR_MIR_BIAS.t1 GNDA 0.027636f
C361 TAIL_CUR_MIR_BIAS.n0 GNDA 0.069525f
C362 TAIL_CUR_MIR_BIAS.t3 GNDA 0.027636f
C363 TAIL_CUR_MIR_BIAS.t6 GNDA 0.027636f
C364 TAIL_CUR_MIR_BIAS.n1 GNDA 0.068809f
C365 TAIL_CUR_MIR_BIAS.n2 GNDA 0.524921f
C366 TAIL_CUR_MIR_BIAS.t7 GNDA 0.027636f
C367 TAIL_CUR_MIR_BIAS.t2 GNDA 0.027636f
C368 TAIL_CUR_MIR_BIAS.n3 GNDA 0.068809f
C369 TAIL_CUR_MIR_BIAS.n4 GNDA 0.349996f
C370 TAIL_CUR_MIR_BIAS.t4 GNDA 0.027636f
C371 TAIL_CUR_MIR_BIAS.t5 GNDA 0.027636f
C372 TAIL_CUR_MIR_BIAS.n5 GNDA 0.066651f
C373 TAIL_CUR_MIR_BIAS.n6 GNDA 0.659828f
C374 PFET_GATE_10uA.t12 GNDA 0.183848f
C375 PFET_GATE_10uA.t29 GNDA 0.183848f
C376 PFET_GATE_10uA.n0 GNDA 0.18877f
C377 PFET_GATE_10uA.t22 GNDA 0.124467f
C378 PFET_GATE_10uA.t24 GNDA 0.220136f
C379 PFET_GATE_10uA.n1 GNDA 0.133438f
C380 PFET_GATE_10uA.t19 GNDA 0.124467f
C381 PFET_GATE_10uA.t17 GNDA 0.220136f
C382 PFET_GATE_10uA.n2 GNDA 0.133438f
C383 PFET_GATE_10uA.n3 GNDA 0.098427f
C384 PFET_GATE_10uA.t18 GNDA 0.124467f
C385 PFET_GATE_10uA.t26 GNDA 0.220136f
C386 PFET_GATE_10uA.n4 GNDA 0.133438f
C387 PFET_GATE_10uA.t15 GNDA 0.124467f
C388 PFET_GATE_10uA.t27 GNDA 0.220136f
C389 PFET_GATE_10uA.n5 GNDA 0.133438f
C390 PFET_GATE_10uA.n6 GNDA 0.115937f
C391 PFET_GATE_10uA.n7 GNDA 1.39925f
C392 PFET_GATE_10uA.t10 GNDA 0.124467f
C393 PFET_GATE_10uA.t13 GNDA 0.124467f
C394 PFET_GATE_10uA.t14 GNDA 0.124467f
C395 PFET_GATE_10uA.t16 GNDA 0.220136f
C396 PFET_GATE_10uA.n8 GNDA 0.149116f
C397 PFET_GATE_10uA.n9 GNDA 0.128616f
C398 PFET_GATE_10uA.n10 GNDA 0.112938f
C399 PFET_GATE_10uA.t23 GNDA 0.124467f
C400 PFET_GATE_10uA.t21 GNDA 0.124467f
C401 PFET_GATE_10uA.t11 GNDA 0.124467f
C402 PFET_GATE_10uA.t28 GNDA 0.124467f
C403 PFET_GATE_10uA.t25 GNDA 0.124467f
C404 PFET_GATE_10uA.t20 GNDA 0.220136f
C405 PFET_GATE_10uA.n11 GNDA 0.149116f
C406 PFET_GATE_10uA.n12 GNDA 0.128616f
C407 PFET_GATE_10uA.n13 GNDA 0.112938f
C408 PFET_GATE_10uA.n14 GNDA 0.09092f
C409 PFET_GATE_10uA.n15 GNDA 0.112938f
C410 PFET_GATE_10uA.n16 GNDA 0.112938f
C411 PFET_GATE_10uA.n17 GNDA 0.09092f
C412 PFET_GATE_10uA.n18 GNDA 0.546176f
C413 PFET_GATE_10uA.n19 GNDA 1.54777f
C414 PFET_GATE_10uA.n20 GNDA 1.84483f
C415 PFET_GATE_10uA.t9 GNDA 0.041489f
C416 PFET_GATE_10uA.t6 GNDA 0.041489f
C417 PFET_GATE_10uA.n21 GNDA 0.106043f
C418 PFET_GATE_10uA.t3 GNDA 0.041489f
C419 PFET_GATE_10uA.t4 GNDA 0.041489f
C420 PFET_GATE_10uA.n22 GNDA 0.103303f
C421 PFET_GATE_10uA.n23 GNDA 1.01043f
C422 PFET_GATE_10uA.t5 GNDA 0.041489f
C423 PFET_GATE_10uA.t0 GNDA 0.041489f
C424 PFET_GATE_10uA.n24 GNDA 0.103303f
C425 PFET_GATE_10uA.n25 GNDA 0.572968f
C426 PFET_GATE_10uA.t7 GNDA 0.606053f
C427 PFET_GATE_10uA.n26 GNDA 1.16968f
C428 PFET_GATE_10uA.t1 GNDA 0.041489f
C429 PFET_GATE_10uA.t8 GNDA 0.041489f
C430 PFET_GATE_10uA.n27 GNDA 0.100062f
C431 PFET_GATE_10uA.n28 GNDA 0.368273f
C432 PFET_GATE_10uA.n29 GNDA 3.97508f
C433 PFET_GATE_10uA.t2 GNDA 0.806816f
C434 Vin+.t1 GNDA 0.125873f
C435 Vin+.t7 GNDA 0.020459f
C436 Vin+.t8 GNDA 0.013299f
C437 Vin+.n0 GNDA 0.04388f
C438 Vin+.t10 GNDA 0.013299f
C439 Vin+.n1 GNDA 0.034146f
C440 Vin+.t9 GNDA 0.013299f
C441 Vin+.n2 GNDA 0.034607f
C442 Vin+.n3 GNDA 0.074523f
C443 Vin+.t5 GNDA 0.043132f
C444 Vin+.t3 GNDA 0.043132f
C445 Vin+.n4 GNDA 0.144858f
C446 Vin+.t2 GNDA 0.043132f
C447 Vin+.t4 GNDA 0.043132f
C448 Vin+.n5 GNDA 0.142496f
C449 Vin+.n6 GNDA 0.656763f
C450 Vin+.n7 GNDA 0.71769f
C451 Vin+.n8 GNDA 0.446219f
C452 Vin+.t0 GNDA 0.137433f
C453 V_TOP.t17 GNDA 0.132312f
C454 V_TOP.t15 GNDA 0.114819f
C455 V_TOP.t36 GNDA 0.114819f
C456 V_TOP.t21 GNDA 0.114819f
C457 V_TOP.t16 GNDA 0.114819f
C458 V_TOP.t14 GNDA 0.114819f
C459 V_TOP.t43 GNDA 0.114819f
C460 V_TOP.t31 GNDA 0.114819f
C461 V_TOP.t27 GNDA 0.114819f
C462 V_TOP.t48 GNDA 0.114819f
C463 V_TOP.t41 GNDA 0.114819f
C464 V_TOP.t38 GNDA 0.114819f
C465 V_TOP.t26 GNDA 0.114819f
C466 V_TOP.t23 GNDA 0.114819f
C467 V_TOP.t40 GNDA 0.114819f
C468 V_TOP.t37 GNDA 0.150097f
C469 V_TOP.n0 GNDA 0.083915f
C470 V_TOP.n1 GNDA 0.061237f
C471 V_TOP.n2 GNDA 0.061237f
C472 V_TOP.n3 GNDA 0.061237f
C473 V_TOP.n4 GNDA 0.061237f
C474 V_TOP.n5 GNDA 0.057104f
C475 V_TOP.t9 GNDA 0.147656f
C476 V_TOP.t6 GNDA 0.155466f
C477 V_TOP.t2 GNDA 0.010935f
C478 V_TOP.t11 GNDA 0.010935f
C479 V_TOP.n6 GNDA 0.027227f
C480 V_TOP.n7 GNDA 0.725415f
C481 V_TOP.t3 GNDA 0.010935f
C482 V_TOP.t12 GNDA 0.010935f
C483 V_TOP.n8 GNDA 0.027411f
C484 V_TOP.t10 GNDA 0.010935f
C485 V_TOP.t1 GNDA 0.010935f
C486 V_TOP.n9 GNDA 0.027227f
C487 V_TOP.n10 GNDA 0.252327f
C488 V_TOP.t7 GNDA 0.010935f
C489 V_TOP.t5 GNDA 0.010935f
C490 V_TOP.n11 GNDA 0.026373f
C491 V_TOP.n12 GNDA 0.153275f
C492 V_TOP.n13 GNDA 0.087481f
C493 V_TOP.t8 GNDA 0.010935f
C494 V_TOP.t4 GNDA 0.010935f
C495 V_TOP.n14 GNDA 0.027227f
C496 V_TOP.n15 GNDA 0.151015f
C497 V_TOP.t13 GNDA 0.010935f
C498 V_TOP.t0 GNDA 0.010935f
C499 V_TOP.n16 GNDA 0.027227f
C500 V_TOP.n17 GNDA 0.149579f
C501 V_TOP.n18 GNDA 0.3288f
C502 V_TOP.n19 GNDA 0.023138f
C503 V_TOP.n20 GNDA 0.057104f
C504 V_TOP.n21 GNDA 0.061237f
C505 V_TOP.n22 GNDA 0.061237f
C506 V_TOP.n23 GNDA 0.061237f
C507 V_TOP.n24 GNDA 0.061237f
C508 V_TOP.n25 GNDA 0.061237f
C509 V_TOP.n26 GNDA 0.061237f
C510 V_TOP.n27 GNDA 0.057104f
C511 V_TOP.t34 GNDA 0.437405f
C512 V_TOP.t49 GNDA 0.444855f
C513 V_TOP.t30 GNDA 0.437405f
C514 V_TOP.n28 GNDA 0.293266f
C515 V_TOP.t24 GNDA 0.437405f
C516 V_TOP.t35 GNDA 0.444855f
C517 V_TOP.t45 GNDA 0.437405f
C518 V_TOP.n29 GNDA 0.293266f
C519 V_TOP.n30 GNDA 0.273378f
C520 V_TOP.t20 GNDA 0.444855f
C521 V_TOP.t39 GNDA 0.437405f
C522 V_TOP.n31 GNDA 0.293266f
C523 V_TOP.t29 GNDA 0.437405f
C524 V_TOP.t44 GNDA 0.444855f
C525 V_TOP.t18 GNDA 0.437405f
C526 V_TOP.n32 GNDA 0.293266f
C527 V_TOP.n33 GNDA 0.355392f
C528 V_TOP.t46 GNDA 0.444855f
C529 V_TOP.t28 GNDA 0.437405f
C530 V_TOP.n34 GNDA 0.293266f
C531 V_TOP.t22 GNDA 0.437405f
C532 V_TOP.t33 GNDA 0.444855f
C533 V_TOP.t42 GNDA 0.437405f
C534 V_TOP.n35 GNDA 0.293266f
C535 V_TOP.n36 GNDA 0.355392f
C536 V_TOP.t25 GNDA 0.444855f
C537 V_TOP.t32 GNDA 0.437405f
C538 V_TOP.n37 GNDA 0.293266f
C539 V_TOP.t47 GNDA 0.437405f
C540 V_TOP.n38 GNDA 0.273378f
C541 V_TOP.t19 GNDA 0.437405f
C542 V_TOP.n39 GNDA 0.191365f
C543 V_TOP.n40 GNDA 0.836546f
C544 V_CMFB_S1.t0 GNDA 0.020333f
C545 V_CMFB_S1.t4 GNDA 0.020333f
C546 V_CMFB_S1.n0 GNDA 0.051153f
C547 V_CMFB_S1.t3 GNDA 0.020333f
C548 V_CMFB_S1.t1 GNDA 0.020333f
C549 V_CMFB_S1.n1 GNDA 0.050626f
C550 V_CMFB_S1.n2 GNDA 0.507984f
C551 V_CMFB_S1.t5 GNDA 0.020333f
C552 V_CMFB_S1.t2 GNDA 0.020333f
C553 V_CMFB_S1.n3 GNDA 0.040665f
C554 V_CMFB_S1.n4 GNDA 0.276616f
C555 VDDA.t217 GNDA 0.57636f
C556 VDDA.t214 GNDA 0.589048f
C557 VDDA.t215 GNDA 0.614289f
C558 VDDA.n0 GNDA 0.41176f
C559 VDDA.t216 GNDA 0.614289f
C560 VDDA.n1 GNDA 0.199909f
C561 VDDA.n2 GNDA 0.256296f
C562 VDDA.n3 GNDA 2.36961f
C563 VDDA.n4 GNDA 0.016683f
C564 VDDA.n5 GNDA 0.012627f
C565 VDDA.n6 GNDA 0.026016f
C566 VDDA.n7 GNDA 0.016683f
C567 VDDA.n8 GNDA 0.016683f
C568 VDDA.n9 GNDA 0.012627f
C569 VDDA.n10 GNDA 0.012627f
C570 VDDA.n11 GNDA 0.0369f
C571 VDDA.n12 GNDA 0.016683f
C572 VDDA.n13 GNDA 0.178687f
C573 VDDA.n14 GNDA 0.178687f
C574 VDDA.t206 GNDA 0.162978f
C575 VDDA.t164 GNDA 0.103225f
C576 VDDA.t127 GNDA 0.103225f
C577 VDDA.t123 GNDA 0.103225f
C578 VDDA.t2 GNDA 0.103225f
C579 VDDA.t18 GNDA 0.103225f
C580 VDDA.t138 GNDA 0.103225f
C581 VDDA.t140 GNDA 0.103225f
C582 VDDA.t108 GNDA 0.103225f
C583 VDDA.t92 GNDA 0.077419f
C584 VDDA.t207 GNDA 0.019584f
C585 VDDA.t205 GNDA 0.012905f
C586 VDDA.n15 GNDA 0.030723f
C587 VDDA.n16 GNDA 0.043715f
C588 VDDA.t189 GNDA 0.019584f
C589 VDDA.t187 GNDA 0.012905f
C590 VDDA.n17 GNDA 0.030723f
C591 VDDA.n18 GNDA 0.016683f
C592 VDDA.n19 GNDA 0.012627f
C593 VDDA.n20 GNDA 0.012627f
C594 VDDA.n21 GNDA 0.016683f
C595 VDDA.n22 GNDA 0.0369f
C596 VDDA.n23 GNDA 0.016683f
C597 VDDA.n24 GNDA 0.012627f
C598 VDDA.n25 GNDA 0.0369f
C599 VDDA.n26 GNDA 0.016683f
C600 VDDA.n27 GNDA 0.013202f
C601 VDDA.n28 GNDA 0.013113f
C602 VDDA.n29 GNDA 0.101934f
C603 VDDA.n30 GNDA 0.013113f
C604 VDDA.n31 GNDA 0.053097f
C605 VDDA.n32 GNDA 0.013113f
C606 VDDA.n33 GNDA 0.053097f
C607 VDDA.n34 GNDA 0.051281f
C608 VDDA.n35 GNDA 0.082182f
C609 VDDA.t198 GNDA 0.019584f
C610 VDDA.t196 GNDA 0.012905f
C611 VDDA.n36 GNDA 0.030723f
C612 VDDA.n37 GNDA 0.043715f
C613 VDDA.t210 GNDA 0.019584f
C614 VDDA.t208 GNDA 0.012905f
C615 VDDA.n38 GNDA 0.030723f
C616 VDDA.n39 GNDA 0.043715f
C617 VDDA.n40 GNDA 0.062561f
C618 VDDA.n41 GNDA 0.082182f
C619 VDDA.n42 GNDA 0.178687f
C620 VDDA.t209 GNDA 0.162978f
C621 VDDA.t29 GNDA 0.103225f
C622 VDDA.t129 GNDA 0.103225f
C623 VDDA.t110 GNDA 0.103225f
C624 VDDA.t12 GNDA 0.103225f
C625 VDDA.t58 GNDA 0.103225f
C626 VDDA.t156 GNDA 0.103225f
C627 VDDA.t104 GNDA 0.103225f
C628 VDDA.t10 GNDA 0.103225f
C629 VDDA.t8 GNDA 0.077419f
C630 VDDA.n43 GNDA 0.051612f
C631 VDDA.t95 GNDA 0.077419f
C632 VDDA.t56 GNDA 0.103225f
C633 VDDA.t144 GNDA 0.103225f
C634 VDDA.t114 GNDA 0.103225f
C635 VDDA.t112 GNDA 0.103225f
C636 VDDA.t4 GNDA 0.103225f
C637 VDDA.t88 GNDA 0.103225f
C638 VDDA.t133 GNDA 0.103225f
C639 VDDA.t83 GNDA 0.103225f
C640 VDDA.t197 GNDA 0.162978f
C641 VDDA.n44 GNDA 0.178687f
C642 VDDA.n45 GNDA 0.051281f
C643 VDDA.n46 GNDA 0.087359f
C644 VDDA.n47 GNDA 0.012627f
C645 VDDA.n48 GNDA 0.0369f
C646 VDDA.n49 GNDA 0.016683f
C647 VDDA.n50 GNDA 0.013113f
C648 VDDA.n51 GNDA 0.053097f
C649 VDDA.n52 GNDA 0.013113f
C650 VDDA.n53 GNDA 0.053097f
C651 VDDA.n54 GNDA 0.013113f
C652 VDDA.n55 GNDA 0.053097f
C653 VDDA.n56 GNDA 0.013113f
C654 VDDA.n57 GNDA 0.076036f
C655 VDDA.n58 GNDA 0.039622f
C656 VDDA.n59 GNDA 0.0369f
C657 VDDA.n60 GNDA 0.027238f
C658 VDDA.n61 GNDA 0.026016f
C659 VDDA.n62 GNDA 0.043715f
C660 VDDA.n63 GNDA 0.062561f
C661 VDDA.n64 GNDA 0.082182f
C662 VDDA.t188 GNDA 0.162978f
C663 VDDA.t121 GNDA 0.103225f
C664 VDDA.t147 GNDA 0.103225f
C665 VDDA.t48 GNDA 0.103225f
C666 VDDA.t125 GNDA 0.103225f
C667 VDDA.t16 GNDA 0.103225f
C668 VDDA.t50 GNDA 0.103225f
C669 VDDA.t162 GNDA 0.103225f
C670 VDDA.t6 GNDA 0.103225f
C671 VDDA.t33 GNDA 0.077419f
C672 VDDA.n65 GNDA 0.051612f
C673 VDDA.n66 GNDA 0.082182f
C674 VDDA.n67 GNDA 0.016683f
C675 VDDA.n68 GNDA 0.0369f
C676 VDDA.n69 GNDA 0.016683f
C677 VDDA.n70 GNDA 0.012627f
C678 VDDA.n71 GNDA 0.0369f
C679 VDDA.n72 GNDA 0.016683f
C680 VDDA.n73 GNDA 0.016683f
C681 VDDA.n74 GNDA 0.012627f
C682 VDDA.n75 GNDA 0.0369f
C683 VDDA.n76 GNDA 0.016683f
C684 VDDA.n77 GNDA 0.012627f
C685 VDDA.n78 GNDA 0.0369f
C686 VDDA.n79 GNDA 0.016683f
C687 VDDA.n80 GNDA 0.027238f
C688 VDDA.n81 GNDA 0.0369f
C689 VDDA.n82 GNDA 0.050506f
C690 VDDA.n83 GNDA 0.153337f
C691 VDDA.t152 GNDA 0.01564f
C692 VDDA.t32 GNDA 0.01564f
C693 VDDA.n84 GNDA 0.05167f
C694 VDDA.n85 GNDA 0.066673f
C695 VDDA.n86 GNDA 0.073249f
C696 VDDA.t190 GNDA 0.074578f
C697 VDDA.t192 GNDA 0.047931f
C698 VDDA.t69 GNDA 0.01564f
C699 VDDA.t136 GNDA 0.01564f
C700 VDDA.n87 GNDA 0.05167f
C701 VDDA.n88 GNDA 0.066673f
C702 VDDA.t25 GNDA 0.01564f
C703 VDDA.t117 GNDA 0.01564f
C704 VDDA.n89 GNDA 0.05167f
C705 VDDA.n90 GNDA 0.066673f
C706 VDDA.t120 GNDA 0.01564f
C707 VDDA.t86 GNDA 0.01564f
C708 VDDA.n91 GNDA 0.05167f
C709 VDDA.n92 GNDA 0.066673f
C710 VDDA.t45 GNDA 0.01564f
C711 VDDA.t42 GNDA 0.01564f
C712 VDDA.n93 GNDA 0.05167f
C713 VDDA.n94 GNDA 0.066673f
C714 VDDA.t55 GNDA 0.01564f
C715 VDDA.t82 GNDA 0.01564f
C716 VDDA.n95 GNDA 0.05167f
C717 VDDA.n96 GNDA 0.066673f
C718 VDDA.t53 GNDA 0.01564f
C719 VDDA.t15 GNDA 0.01564f
C720 VDDA.n97 GNDA 0.05167f
C721 VDDA.n98 GNDA 0.066673f
C722 VDDA.t39 GNDA 0.01564f
C723 VDDA.t74 GNDA 0.01564f
C724 VDDA.n99 GNDA 0.05167f
C725 VDDA.n100 GNDA 0.066673f
C726 VDDA.t174 GNDA 0.019584f
C727 VDDA.n101 GNDA 0.030877f
C728 VDDA.n102 GNDA 0.017804f
C729 VDDA.n103 GNDA 0.031643f
C730 VDDA.t204 GNDA 0.019584f
C731 VDDA.n104 GNDA 0.030877f
C732 VDDA.n105 GNDA 0.031643f
C733 VDDA.n106 GNDA 0.031643f
C734 VDDA.n107 GNDA 0.025963f
C735 VDDA.n108 GNDA 0.131054f
C736 VDDA.t173 GNDA 0.158968f
C737 VDDA.t43 GNDA 0.070967f
C738 VDDA.n109 GNDA 0.047311f
C739 VDDA.t94 GNDA 0.070967f
C740 VDDA.t203 GNDA 0.156658f
C741 VDDA.n110 GNDA 0.124763f
C742 VDDA.n111 GNDA 0.025963f
C743 VDDA.n112 GNDA 0.017804f
C744 VDDA.n113 GNDA 0.025013f
C745 VDDA.n114 GNDA 0.073615f
C746 VDDA.n115 GNDA 0.089006f
C747 VDDA.n116 GNDA 0.059995f
C748 VDDA.n117 GNDA 0.269888f
C749 VDDA.n118 GNDA 0.269888f
C750 VDDA.t200 GNDA 0.348246f
C751 VDDA.t151 GNDA 0.251024f
C752 VDDA.t31 GNDA 0.251024f
C753 VDDA.t68 GNDA 0.251024f
C754 VDDA.t135 GNDA 0.251024f
C755 VDDA.t24 GNDA 0.251024f
C756 VDDA.t116 GNDA 0.251024f
C757 VDDA.t119 GNDA 0.251024f
C758 VDDA.t85 GNDA 0.188268f
C759 VDDA.n119 GNDA 0.073249f
C760 VDDA.n120 GNDA 0.11513f
C761 VDDA.n121 GNDA 0.11513f
C762 VDDA.t191 GNDA 0.348246f
C763 VDDA.t73 GNDA 0.251024f
C764 VDDA.t38 GNDA 0.251024f
C765 VDDA.t14 GNDA 0.251024f
C766 VDDA.t52 GNDA 0.251024f
C767 VDDA.t81 GNDA 0.251024f
C768 VDDA.t54 GNDA 0.251024f
C769 VDDA.t41 GNDA 0.251024f
C770 VDDA.t44 GNDA 0.188268f
C771 VDDA.n122 GNDA 0.125512f
C772 VDDA.n123 GNDA 0.114601f
C773 VDDA.n124 GNDA 0.084457f
C774 VDDA.n125 GNDA 0.059995f
C775 VDDA.t201 GNDA 0.047931f
C776 VDDA.t199 GNDA 0.074578f
C777 VDDA.n126 GNDA 0.089006f
C778 VDDA.n127 GNDA 0.044506f
C779 VDDA.n128 GNDA 0.012591f
C780 VDDA.t195 GNDA 0.01973f
C781 VDDA.t193 GNDA 0.030994f
C782 VDDA.n129 GNDA 0.029171f
C783 VDDA.n130 GNDA 0.021297f
C784 VDDA.n131 GNDA 0.038772f
C785 VDDA.t168 GNDA 0.01973f
C786 VDDA.t166 GNDA 0.030994f
C787 VDDA.n132 GNDA 0.029171f
C788 VDDA.n133 GNDA 0.038772f
C789 VDDA.n134 GNDA 0.038772f
C790 VDDA.n135 GNDA 0.029697f
C791 VDDA.n136 GNDA 0.154692f
C792 VDDA.t194 GNDA 0.203013f
C793 VDDA.t102 GNDA 0.116128f
C794 VDDA.n137 GNDA 0.077419f
C795 VDDA.t75 GNDA 0.116128f
C796 VDDA.t167 GNDA 0.200997f
C797 VDDA.n138 GNDA 0.148106f
C798 VDDA.n139 GNDA 0.029697f
C799 VDDA.n140 GNDA 0.021297f
C800 VDDA.n141 GNDA 0.026067f
C801 VDDA.n142 GNDA 0.03484f
C802 VDDA.n143 GNDA 0.072535f
C803 VDDA.n144 GNDA 0.124757f
C804 VDDA.n145 GNDA 0.012981f
C805 VDDA.n146 GNDA 0.053229f
C806 VDDA.n147 GNDA 0.03446f
C807 VDDA.t175 GNDA 0.032051f
C808 VDDA.t177 GNDA 0.019635f
C809 VDDA.n148 GNDA 0.012981f
C810 VDDA.n149 GNDA 0.053229f
C811 VDDA.n150 GNDA 0.012981f
C812 VDDA.n151 GNDA 0.053229f
C813 VDDA.n152 GNDA 0.048643f
C814 VDDA.t169 GNDA 0.032051f
C815 VDDA.t171 GNDA 0.019635f
C816 VDDA.n153 GNDA 0.012981f
C817 VDDA.n154 GNDA 0.053229f
C818 VDDA.n155 GNDA 0.012981f
C819 VDDA.n156 GNDA 0.053229f
C820 VDDA.n157 GNDA 0.012981f
C821 VDDA.n158 GNDA 0.053229f
C822 VDDA.n159 GNDA 0.012981f
C823 VDDA.n160 GNDA 0.053229f
C824 VDDA.n161 GNDA 0.012981f
C825 VDDA.n162 GNDA 0.053229f
C826 VDDA.n163 GNDA 0.03446f
C827 VDDA.t178 GNDA 0.032051f
C828 VDDA.t180 GNDA 0.019635f
C829 VDDA.n164 GNDA 0.012981f
C830 VDDA.n165 GNDA 0.073054f
C831 VDDA.n166 GNDA 0.036146f
C832 VDDA.n167 GNDA 0.026511f
C833 VDDA.n168 GNDA 0.158888f
C834 VDDA.n169 GNDA 0.158888f
C835 VDDA.t212 GNDA 0.204433f
C836 VDDA.t149 GNDA 0.157183f
C837 VDDA.t160 GNDA 0.117887f
C838 VDDA.n170 GNDA 0.03446f
C839 VDDA.n171 GNDA 0.048015f
C840 VDDA.n172 GNDA 0.048015f
C841 VDDA.t179 GNDA 0.204433f
C842 VDDA.t66 GNDA 0.157183f
C843 VDDA.t142 GNDA 0.117887f
C844 VDDA.n173 GNDA 0.078592f
C845 VDDA.n174 GNDA 0.048015f
C846 VDDA.n175 GNDA 0.028152f
C847 VDDA.n176 GNDA 0.026511f
C848 VDDA.t213 GNDA 0.019635f
C849 VDDA.t211 GNDA 0.032051f
C850 VDDA.n177 GNDA 0.034709f
C851 VDDA.n178 GNDA 0.035338f
C852 VDDA.n179 GNDA 0.035338f
C853 VDDA.n180 GNDA 0.034709f
C854 VDDA.n181 GNDA 0.040587f
C855 VDDA.n182 GNDA 0.187253f
C856 VDDA.n183 GNDA 0.187253f
C857 VDDA.t185 GNDA 0.204433f
C858 VDDA.t154 GNDA 0.157183f
C859 VDDA.t64 GNDA 0.157183f
C860 VDDA.t62 GNDA 0.157183f
C861 VDDA.t27 GNDA 0.157183f
C862 VDDA.t77 GNDA 0.117887f
C863 VDDA.n184 GNDA 0.048643f
C864 VDDA.n185 GNDA 0.075953f
C865 VDDA.n186 GNDA 0.075953f
C866 VDDA.t170 GNDA 0.204433f
C867 VDDA.t100 GNDA 0.157183f
C868 VDDA.t20 GNDA 0.157183f
C869 VDDA.t70 GNDA 0.157183f
C870 VDDA.t22 GNDA 0.157183f
C871 VDDA.t60 GNDA 0.117887f
C872 VDDA.n187 GNDA 0.078592f
C873 VDDA.n188 GNDA 0.075953f
C874 VDDA.n189 GNDA 0.056304f
C875 VDDA.n190 GNDA 0.040587f
C876 VDDA.t186 GNDA 0.019635f
C877 VDDA.t184 GNDA 0.032051f
C878 VDDA.n191 GNDA 0.034709f
C879 VDDA.n192 GNDA 0.035338f
C880 VDDA.n193 GNDA 0.035338f
C881 VDDA.n194 GNDA 0.034709f
C882 VDDA.n195 GNDA 0.026511f
C883 VDDA.n196 GNDA 0.157631f
C884 VDDA.n197 GNDA 0.157631f
C885 VDDA.t182 GNDA 0.200997f
C886 VDDA.t35 GNDA 0.154837f
C887 VDDA.t106 GNDA 0.116128f
C888 VDDA.n198 GNDA 0.03446f
C889 VDDA.n199 GNDA 0.048015f
C890 VDDA.n200 GNDA 0.048015f
C891 VDDA.t176 GNDA 0.200997f
C892 VDDA.t90 GNDA 0.154837f
C893 VDDA.t0 GNDA 0.116128f
C894 VDDA.n201 GNDA 0.077419f
C895 VDDA.n202 GNDA 0.048015f
C896 VDDA.n203 GNDA 0.028152f
C897 VDDA.n204 GNDA 0.026511f
C898 VDDA.t183 GNDA 0.019635f
C899 VDDA.t181 GNDA 0.032051f
C900 VDDA.n205 GNDA 0.034709f
C901 VDDA.n206 GNDA 0.049286f
C902 VDDA.n207 GNDA 0.088755f
C903 VDDA.t87 GNDA 0.291427f
C904 VDDA.t72 GNDA 0.292484f
C905 VDDA.t37 GNDA 0.291427f
C906 VDDA.t132 GNDA 0.292484f
C907 VDDA.t98 GNDA 0.291427f
C908 VDDA.t118 GNDA 0.292484f
C909 VDDA.t26 GNDA 0.291427f
C910 VDDA.t47 GNDA 0.292484f
C911 VDDA.t80 GNDA 0.291427f
C912 VDDA.t137 GNDA 0.292484f
C913 VDDA.t99 GNDA 0.291427f
C914 VDDA.t158 GNDA 0.292484f
C915 VDDA.t79 GNDA 0.291427f
C916 VDDA.t159 GNDA 0.292484f
C917 VDDA.t153 GNDA 0.291427f
C918 VDDA.t46 GNDA 0.292484f
C919 VDDA.n208 GNDA 0.195344f
C920 VDDA.t146 GNDA 0.155563f
C921 VDDA.n209 GNDA 0.211953f
C922 VDDA.t97 GNDA 0.155563f
C923 VDDA.n210 GNDA 0.211953f
C924 VDDA.t131 GNDA 0.155563f
C925 VDDA.n211 GNDA 0.211953f
C926 VDDA.t40 GNDA 0.232131f
C927 VDDA.n212 GNDA 0.202273f
.ends

