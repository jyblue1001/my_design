* PEX produced on Sat Jan 25 03:13:23 PM CET 2025 using ./iic-pex.sh with m=2 and s=1
* NGSPICE file created from pfd_3.ext - technology: sky130A

.subckt pfd_3
X0 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_4.Y a_3115_297# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_4.B a_1593_47# sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4 sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_3115_297# sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X13 a_135_297# sky130_fd_sc_hd__nor2_1_4.A sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X14 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_1099_n953# sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X17 a_135_n953# sky130_fd_sc_hd__nor2_1_0.A sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X18 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_4.A sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X23 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X26 sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_5.B a_625_297# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X27 a_3115_n953# sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X28 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_1.Y a_1099_297# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X29 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_1593_47# sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X32 a_625_n953# sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X33 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_1.Y a_1099_n953# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X34 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.Y a_3115_n953# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X35 a_625_297# sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X36 sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X37 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.A sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.B a_135_n953# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X39 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X41 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_4.B a_135_297# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X42 a_1099_297# sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X43 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X44 sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_2.B a_625_n953# sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X45 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__nor2_1_7.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
C0 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.25991f
C1 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_1.A 0.060251f
C2 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__nor2_1_0.Y 0.015649f
C3 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_4.B 0.428538f
C4 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_5.Y 0.193757f
C5 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_2.B 0.301379f
C6 sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.687357f
C7 sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_0.VGND 0.204585f
C8 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_4.A 0.06019f
C9 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_4.A 0.064249f
C10 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_2.Y 0.193177f
C11 sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__inv_1_1.Y 0.051591f
C12 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_4.A 0.058413f
C13 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_0.VPB 0.127396f
C14 sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.665829f
C15 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_0.VPWR 1.45635f
C16 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.175327f
C17 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.VGND 0.886022f
C18 sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_0.Y 0.085339f
C19 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_4.B 0.280668f
C20 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_0.B 0.238995f
C21 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.A 0.064207f
C22 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_5.Y 0.021511f
C23 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.VGND 0.538795f
C24 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_0.VGND 0.48823f
C25 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__nor2_1_5.Y 0.110928f
C26 sky130_fd_sc_hd__nor2_1_4.Y a_135_297# 0.011374f
C27 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.A 0.058413f
C28 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__nor2_1_2.Y 0.014764f
C29 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_2.Y 0.130437f
C30 a_3115_n953# sky130_fd_sc_hd__nor2_1_0.B 0.01129f
C31 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_1.A 0.196269f
C32 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.Y 1.31604f
C33 a_135_n953# sky130_fd_sc_hd__nor2_1_0.Y 0.011374f
C34 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_4.A 0.048086f
C35 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nand2_1_1.Y 0.061816f
C36 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.VPWR 0.259501f
C37 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__nor2_1_2.Y 0.130172f
C38 sky130_fd_sc_hd__nor2_1_4.A sky130_fd_sc_hd__nor2_1_0.VGND 0.049683f
C39 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_5.B 0.085332f
C40 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_4.A 0.054114f
C41 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_0.Y 0.349326f
C42 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_4.A 0.197834f
C43 sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__inv_1_1.Y 0.092839f
C44 sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__inv_1_1.Y 0.053871f
C45 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.B 0.05302f
C46 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_4.B 0.213728f
C47 a_625_n953# sky130_fd_sc_hd__nor2_1_2.Y 0.0113f
C48 a_1099_n953# sky130_fd_sc_hd__nor2_1_2.B 0.011338f
C49 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_0.VGND 0.181232f
C50 sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_5.Y 0.299059f
C51 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__inv_1_4.A 0.024648f
C52 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__inv_1_4.A 0.028663f
C53 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_0.A 0.045926f
C54 sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_2.Y 0.100358f
C55 sky130_fd_sc_hd__nor2_1_0.A sky130_fd_sc_hd__nor2_1_0.VGND 0.049683f
C56 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_1.Y 0.268597f
C57 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__inv_1_1.A 0.127725f
C58 sky130_fd_sc_hd__nor2_1_5.B a_1099_297# 0.01129f
C59 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_5.B 0.159438f
C60 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__inv_1_1.Y 0.017081f
C61 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__inv_1_1.Y 0.252155f
C62 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_0.Y 0.467302f
C63 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__nor2_1_0.VGND 0.174115f
C64 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.260124f
C65 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.VPB 0.081018f
C66 sky130_fd_sc_hd__nor2_1_4.B a_3115_297# 0.01129f
C67 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__nor2_1_2.Y 0.014874f
C68 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_5.Y 0.130618f
C69 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.227252f
C70 sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_4.B 0.011732f
C71 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__inv_1_4.A 0.125052f
C72 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__inv_1_0.A 0.196292f
C73 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_0.A 0.047251f
C74 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__nor2_1_0.VGND 0.31793f
C75 sky130_fd_sc_hd__nor2_1_5.Y a_625_297# 0.0113f
C76 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__nor2_1_0.Y 0.015525f
C77 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_4.Y 0.015545f
C78 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_0.VPWR 1.33441f
C79 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__inv_1_1.Y 0.17549f
C80 sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_0.VGND 0.423942f
C81 sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_2.Y 0.016719f
C82 sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_2.Y 0.298166f
C83 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_4.B 0.358704f
C84 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_5.B 0.302178f
C85 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_5.Y 0.02609f
C86 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_5.Y 0.187607f
C87 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_2.B 0.159412f
C88 sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_0.VGND 0.204379f
C89 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_5.Y 0.032475f
C90 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_5.Y 0.804239f
C91 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__inv_1_0.A 0.128036f
C92 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_2.B 0.010272f
C93 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__nor2_1_0.VGND 0.1765f
C94 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__inv_1_1.Y 0.061228f
C95 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_2.Y 0.187294f
C96 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_4.A 0.047251f
C97 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__inv_1_1.Y 0.015497f
C98 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_0.VPWR 0.196439f
C99 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_2.Y 0.741418f
C100 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_0.VPB 0.50148f
C101 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_0.B 0.182946f
C102 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_4.B 0.187715f
C103 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__nor2_1_7.VNB 0.212781f
C104 sky130_fd_sc_hd__inv_1_1.A sky130_fd_sc_hd__nor2_1_7.VNB 0.211599f
C105 sky130_fd_sc_hd__nor2_1_2.B sky130_fd_sc_hd__nor2_1_7.VNB 0.180291f
C106 sky130_fd_sc_hd__nor2_1_2.Y sky130_fd_sc_hd__nor2_1_7.VNB 1.31564f
C107 sky130_fd_sc_hd__nor2_1_0.Y sky130_fd_sc_hd__nor2_1_7.VNB 1.22213f
C108 sky130_fd_sc_hd__nor2_1_0.A sky130_fd_sc_hd__nor2_1_7.VNB 0.142405f
C109 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__nor2_1_7.VNB 0.366837f
C110 sky130_fd_sc_hd__nor2_1_0.VGND sky130_fd_sc_hd__nor2_1_7.VNB 2.10724f
C111 sky130_fd_sc_hd__nor2_1_0.VPWR sky130_fd_sc_hd__nor2_1_7.VNB 2.06194f
C112 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__nor2_1_7.VNB 0.209443f
C113 sky130_fd_sc_hd__nand2_1_1.Y sky130_fd_sc_hd__nor2_1_7.VNB 0.190018f
C114 sky130_fd_sc_hd__nor2_1_0.B sky130_fd_sc_hd__nor2_1_7.VNB 2.15242f
C115 sky130_fd_sc_hd__inv_1_1.Y sky130_fd_sc_hd__nor2_1_7.VNB 0.458688f
C116 sky130_fd_sc_hd__nor2_1_5.Y sky130_fd_sc_hd__nor2_1_7.VNB 1.25998f
C117 sky130_fd_sc_hd__nor2_1_5.B sky130_fd_sc_hd__nor2_1_7.VNB 0.177353f
C118 sky130_fd_sc_hd__nor2_1_4.B sky130_fd_sc_hd__nor2_1_7.VNB 2.27583f
C119 sky130_fd_sc_hd__nor2_1_4.A sky130_fd_sc_hd__nor2_1_7.VNB 0.140245f
C120 sky130_fd_sc_hd__nor2_1_4.Y sky130_fd_sc_hd__nor2_1_7.VNB 1.18392f
C121 sky130_fd_sc_hd__nor2_1_0.VPB sky130_fd_sc_hd__nor2_1_7.VNB 8.02312f
.ends

