* PEX produced on Fri Jul  4 11:27:02 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t308 bgr_0.V_TOP.t14 bgr_0.Vin-.t4 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 a_9610_5930.t8 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 bgr_0.V_TOP.t15 VDDA.t306 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t174 GNDA.t176 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X5 two_stage_opamp_dummy_magic_0.VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t96 GNDA.t173 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 two_stage_opamp_dummy_magic_0.X.t13 GNDA.t185 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X8 two_stage_opamp_dummy_magic_0.VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 two_stage_opamp_dummy_magic_0.VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 bgr_0.NFET_GATE_10uA.t2 bgr_0.NFET_GATE_10uA.t1 GNDA.t278 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X11 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 bgr_0.V_TOP.t16 VDDA.t305 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 VDDA.t115 bgr_0.V_mir2.t14 bgr_0.V_mir2.t15 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X14 two_stage_opamp_dummy_magic_0.V_err_gate.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 two_stage_opamp_dummy_magic_0.VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 two_stage_opamp_dummy_magic_0.VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 a_8420_8490.t10 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD3.t7 w_8160_8260.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X18 VDDA.t154 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.VOUT+.t13 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X19 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X20 two_stage_opamp_dummy_magic_0.VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 two_stage_opamp_dummy_magic_0.VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t168 two_stage_opamp_dummy_magic_0.Y.t14 two_stage_opamp_dummy_magic_0.VOUT+.t12 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X23 VDDA.t230 bgr_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 VDDA.t229 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X24 two_stage_opamp_dummy_magic_0.VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 a_14520_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X26 bgr_0.V_TOP.t17 VDDA.t304 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 two_stage_opamp_dummy_magic_0.VOUT-.t8 GNDA.t170 GNDA.t172 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X28 VDDA.t166 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X29 VDDA.t3 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X30 two_stage_opamp_dummy_magic_0.VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X32 two_stage_opamp_dummy_magic_0.VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_0.VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 two_stage_opamp_dummy_magic_0.VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 two_stage_opamp_dummy_magic_0.VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 two_stage_opamp_dummy_magic_0.VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 two_stage_opamp_dummy_magic_0.VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 two_stage_opamp_dummy_magic_0.V_p_mir.t3 bgr_0.TAIL_CUR_MIR_BIAS.t12 GNDA.t46 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X40 VDDA.t13 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.VOUT-.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X41 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_0.Y.t15 VDDA.t226 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X42 two_stage_opamp_dummy_magic_0.VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 bgr_0.V_mir2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 bgr_0.V_p_2.t4 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X44 bgr_0.Vin-.t7 bgr_0.V_TOP.t18 VDDA.t303 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X45 VDDA.t423 VDDA.t421 two_stage_opamp_dummy_magic_0.V_err_gate.t12 VDDA.t422 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X46 GNDA.t284 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t283 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X47 GNDA.t50 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 two_stage_opamp_dummy_magic_0.V_err_p.t17 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t160 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X49 two_stage_opamp_dummy_magic_0.VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 two_stage_opamp_dummy_magic_0.VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 a_8420_8490.t9 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD3.t13 w_8160_8260.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X52 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X53 two_stage_opamp_dummy_magic_0.Y.t4 a_10530_5140# two_stage_opamp_dummy_magic_0.VD1.t17 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X54 two_stage_opamp_dummy_magic_0.VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 two_stage_opamp_dummy_magic_0.VOUT-.t16 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA.t280 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X56 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 two_stage_opamp_dummy_magic_0.Y.t16 GNDA.t190 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X57 bgr_0.1st_Vout_1.t10 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t337 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X58 two_stage_opamp_dummy_magic_0.VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 GNDA.t72 bgr_0.TAIL_CUR_MIR_BIAS.t13 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X61 VDDA.t420 VDDA.t418 bgr_0.V_TOP.t5 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X62 GNDA.t314 bgr_0.TAIL_CUR_MIR_BIAS.t14 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA.t313 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X63 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 two_stage_opamp_dummy_magic_0.X.t15 VDDA.t14 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X64 two_stage_opamp_dummy_magic_0.VD1.t7 VIN-.t0 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X65 two_stage_opamp_dummy_magic_0.V_err_p.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 two_stage_opamp_dummy_magic_0.VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 GNDA.t52 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X68 GNDA.t169 GNDA.t167 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X69 VDDA.t455 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t8 VDDA.t454 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X70 two_stage_opamp_dummy_magic_0.VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 two_stage_opamp_dummy_magic_0.VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 two_stage_opamp_dummy_magic_0.err_amp_out.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 a_9610_5930.t0 GNDA.t307 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 two_stage_opamp_dummy_magic_0.VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 two_stage_opamp_dummy_magic_0.VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 two_stage_opamp_dummy_magic_0.VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 two_stage_opamp_dummy_magic_0.VD1.t19 VIN-.t1 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X77 two_stage_opamp_dummy_magic_0.VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_0.NFET_GATE_10uA.t3 bgr_0.PFET_GATE_10uA.t11 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X79 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 a_9610_5930.t1 GNDA.t306 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X80 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VDDA.t41 bgr_0.PFET_GATE_10uA.t12 bgr_0.TAIL_CUR_MIR_BIAS.t11 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X82 GNDA.t166 GNDA.t164 two_stage_opamp_dummy_magic_0.Y.t2 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X83 two_stage_opamp_dummy_magic_0.VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VDDA.t417 VDDA.t415 bgr_0.NFET_GATE_10uA.t4 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X85 two_stage_opamp_dummy_magic_0.X.t5 GNDA.t161 GNDA.t163 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X86 VDDA.t449 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.VOUT+.t11 VDDA.t448 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X87 VDDA.t35 bgr_0.1st_Vout_1.t14 bgr_0.V_TOP.t0 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X88 GNDA.t160 GNDA.t158 two_stage_opamp_dummy_magic_0.VD1.t4 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X89 two_stage_opamp_dummy_magic_0.VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 two_stage_opamp_dummy_magic_0.VD4.t19 VDDA.t412 VDDA.t414 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X91 two_stage_opamp_dummy_magic_0.VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_0.VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 two_stage_opamp_dummy_magic_0.VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 VDDA.t203 bgr_0.V_mir2.t12 bgr_0.V_mir2.t13 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X95 w_10220_8260.t5 w_10220_8260.t3 a_10480_8490.t1 w_10220_8260.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X96 GNDA.t268 bgr_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t267 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X97 VDDA.t156 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t15 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X98 two_stage_opamp_dummy_magic_0.VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 two_stage_opamp_dummy_magic_0.Vb3.t6 bgr_0.NFET_GATE_10uA.t9 GNDA.t270 GNDA.t269 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X100 GNDA.t157 GNDA.t155 two_stage_opamp_dummy_magic_0.VD1.t3 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X101 VDDA.t213 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t9 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X102 two_stage_opamp_dummy_magic_0.VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 bgr_0.V_TOP.t13 bgr_0.cap_res1.t20 GNDA.t233 sky130_fd_pr__res_high_po_0p35 l=2.05
X104 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 two_stage_opamp_dummy_magic_0.Y.t18 VDDA.t111 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X105 two_stage_opamp_dummy_magic_0.V_p.t37 bgr_0.TAIL_CUR_MIR_BIAS.t15 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X106 a_11220_17410.t0 GNDA.t30 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X107 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 two_stage_opamp_dummy_magic_0.Y.t19 VDDA.t468 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X108 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X109 two_stage_opamp_dummy_magic_0.VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 two_stage_opamp_dummy_magic_0.Vb1.t0 bgr_0.PFET_GATE_10uA.t13 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X111 two_stage_opamp_dummy_magic_0.VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 two_stage_opamp_dummy_magic_0.VOUT-.t6 a_5750_2276.t0 GNDA.t64 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X113 bgr_0.PFET_GATE_10uA.t3 bgr_0.1st_Vout_2.t13 VDDA.t240 VDDA.t239 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X114 two_stage_opamp_dummy_magic_0.VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 GNDA.t55 bgr_0.TAIL_CUR_MIR_BIAS.t16 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X116 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.Vb3.t8 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 two_stage_opamp_dummy_magic_0.VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 two_stage_opamp_dummy_magic_0.VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 two_stage_opamp_dummy_magic_0.VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 two_stage_opamp_dummy_magic_0.VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 two_stage_opamp_dummy_magic_0.VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VDDA.t123 bgr_0.V_mir1.t10 bgr_0.V_mir1.t11 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X123 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 two_stage_opamp_dummy_magic_0.X.t16 VDDA.t30 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X124 two_stage_opamp_dummy_magic_0.VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 two_stage_opamp_dummy_magic_0.VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 a_9610_5930.t7 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X127 two_stage_opamp_dummy_magic_0.VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VDDA.t5 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.Vb3.t9 VDDA.t133 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X131 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t17 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X132 bgr_0.V_TOP.t19 VDDA.t301 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.Vb2.t13 a_8420_8490.t8 w_8160_8260.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X134 two_stage_opamp_dummy_magic_0.VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 two_stage_opamp_dummy_magic_0.VD1.t16 a_10530_5140# two_stage_opamp_dummy_magic_0.Y.t10 GNDA.t247 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X137 two_stage_opamp_dummy_magic_0.VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 a_14640_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA.t78 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X139 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X140 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA.t152 GNDA.t154 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X141 two_stage_opamp_dummy_magic_0.VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 two_stage_opamp_dummy_magic_0.VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 two_stage_opamp_dummy_magic_0.V_p.t5 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X144 two_stage_opamp_dummy_magic_0.VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VDDA.t209 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t5 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X146 two_stage_opamp_dummy_magic_0.VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 two_stage_opamp_dummy_magic_0.VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 a_13730_17020.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t27 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X150 GNDA.t230 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X151 two_stage_opamp_dummy_magic_0.V_p.t16 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X152 two_stage_opamp_dummy_magic_0.VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 bgr_0.V_CUR_REF_REG.t0 VDDA.t409 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X154 a_11220_17410.t1 a_12828_17530.t1 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X155 two_stage_opamp_dummy_magic_0.VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VDDA.t195 two_stage_opamp_dummy_magic_0.X.t19 two_stage_opamp_dummy_magic_0.VOUT-.t13 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X157 two_stage_opamp_dummy_magic_0.VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 bgr_0.TAIL_CUR_MIR_BIAS.t10 bgr_0.PFET_GATE_10uA.t14 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X159 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 two_stage_opamp_dummy_magic_0.Y.t20 VDDA.t70 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X160 two_stage_opamp_dummy_magic_0.VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 two_stage_opamp_dummy_magic_0.VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 two_stage_opamp_dummy_magic_0.V_p.t35 bgr_0.TAIL_CUR_MIR_BIAS.t17 GNDA.t182 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X163 VDDA.t437 bgr_0.PFET_GATE_10uA.t15 bgr_0.V_CUR_REF_REG.t2 VDDA.t436 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X164 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X165 two_stage_opamp_dummy_magic_0.VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 bgr_0.PFET_GATE_10uA.t2 bgr_0.cap_res2.t20 GNDA.t233 sky130_fd_pr__res_high_po_0p35 l=2.05
X167 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.Vb2.t14 a_8420_8490.t7 w_8160_8260.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X168 bgr_0.V_p_1.t9 bgr_0.Vin-.t8 bgr_0.V_mir1.t13 GNDA.t289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X169 VDDA.t459 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t458 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 two_stage_opamp_dummy_magic_0.VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 two_stage_opamp_dummy_magic_0.VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 GNDA.t151 GNDA.t149 two_stage_opamp_dummy_magic_0.X.t4 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X173 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 two_stage_opamp_dummy_magic_0.VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 two_stage_opamp_dummy_magic_0.VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VDDA.t121 bgr_0.1st_Vout_1.t19 bgr_0.V_TOP.t4 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X177 VDDA.t300 bgr_0.V_TOP.t20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X178 two_stage_opamp_dummy_magic_0.VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 GNDA.t220 bgr_0.TAIL_CUR_MIR_BIAS.t18 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X180 two_stage_opamp_dummy_magic_0.VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t3 bgr_0.1st_Vout_2.t9 GNDA.t312 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X182 two_stage_opamp_dummy_magic_0.VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 two_stage_opamp_dummy_magic_0.VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 two_stage_opamp_dummy_magic_0.VOUT-.t12 two_stage_opamp_dummy_magic_0.X.t20 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X185 two_stage_opamp_dummy_magic_0.VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 bgr_0.V_p_1.t8 bgr_0.Vin-.t9 bgr_0.V_mir1.t12 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X187 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 GNDA.t191 bgr_0.TAIL_CUR_MIR_BIAS.t19 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X189 bgr_0.V_TOP.t3 VDDA.t406 VDDA.t408 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X190 two_stage_opamp_dummy_magic_0.VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 bgr_0.Vin-.t2 bgr_0.START_UP.t6 bgr_0.V_TOP.t7 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X192 VDDA.t405 VDDA.t403 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X193 two_stage_opamp_dummy_magic_0.VD1.t15 a_10530_5140# two_stage_opamp_dummy_magic_0.Y.t7 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X194 two_stage_opamp_dummy_magic_0.VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 two_stage_opamp_dummy_magic_0.VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 bgr_0.V_TOP.t21 VDDA.t290 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 two_stage_opamp_dummy_magic_0.err_amp_out.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t6 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X199 two_stage_opamp_dummy_magic_0.VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 two_stage_opamp_dummy_magic_0.VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 VDDA.t425 two_stage_opamp_dummy_magic_0.Vb3.t11 two_stage_opamp_dummy_magic_0.VD4.t20 VDDA.t424 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X202 GNDA.t218 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X203 two_stage_opamp_dummy_magic_0.VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 two_stage_opamp_dummy_magic_0.V_p.t32 bgr_0.TAIL_CUR_MIR_BIAS.t20 GNDA.t196 GNDA.t195 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X205 a_13730_17020.t0 GNDA.t28 GNDA.t27 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X206 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 bgr_0.V_TOP.t22 VDDA.t289 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 w_8160_8260.t5 w_8160_8260.t3 a_8420_8490.t11 w_8160_8260.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X209 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t400 VDDA.t402 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X210 a_11220_17290.t1 a_12828_17650.t1 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X211 VDDA.t248 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD3.t18 VDDA.t247 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X212 two_stage_opamp_dummy_magic_0.VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 two_stage_opamp_dummy_magic_0.VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 two_stage_opamp_dummy_magic_0.VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 two_stage_opamp_dummy_magic_0.VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 bgr_0.V_p_2.t8 bgr_0.V_CUR_REF_REG.t4 bgr_0.1st_Vout_2.t8 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X217 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 bgr_0.PFET_GATE_10uA.t16 VDDA.t95 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X218 two_stage_opamp_dummy_magic_0.VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VDDA.t183 bgr_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X220 two_stage_opamp_dummy_magic_0.V_p.t4 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X221 two_stage_opamp_dummy_magic_0.VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 GNDA.t75 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 two_stage_opamp_dummy_magic_0.VOUT+.t0 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X223 GNDA.t229 two_stage_opamp_dummy_magic_0.X.t21 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X224 a_11220_17290.t0 GNDA.t73 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X225 two_stage_opamp_dummy_magic_0.V_p.t40 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA.t334 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X226 bgr_0.TAIL_CUR_MIR_BIAS.t1 GNDA.t146 GNDA.t148 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X227 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 two_stage_opamp_dummy_magic_0.VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 two_stage_opamp_dummy_magic_0.VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 bgr_0.START_UP.t3 bgr_0.V_TOP.t23 VDDA.t298 VDDA.t297 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X231 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t6 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X232 two_stage_opamp_dummy_magic_0.V_p.t31 bgr_0.TAIL_CUR_MIR_BIAS.t21 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X233 bgr_0.1st_Vout_2.t4 bgr_0.V_mir2.t18 VDDA.t211 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X234 bgr_0.V_TOP.t24 VDDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 two_stage_opamp_dummy_magic_0.VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 two_stage_opamp_dummy_magic_0.VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 two_stage_opamp_dummy_magic_0.VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 two_stage_opamp_dummy_magic_0.VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 VDDA.t244 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD4.t16 VDDA.t243 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X240 VDDA.t457 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t9 VDDA.t456 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X241 two_stage_opamp_dummy_magic_0.VOUT+.t10 two_stage_opamp_dummy_magic_0.Y.t22 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X242 two_stage_opamp_dummy_magic_0.VD2.t12 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t6 GNDA.t204 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X243 two_stage_opamp_dummy_magic_0.VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 two_stage_opamp_dummy_magic_0.VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 GNDA.t202 bgr_0.TAIL_CUR_MIR_BIAS.t22 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X247 bgr_0.V_p_2.t7 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t7 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X248 GNDA.t145 GNDA.t143 two_stage_opamp_dummy_magic_0.VOUT+.t2 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X249 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_0.X.t22 VDDA.t249 GNDA.t266 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X250 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t397 VDDA.t399 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X251 two_stage_opamp_dummy_magic_0.VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X252 two_stage_opamp_dummy_magic_0.VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 VDDA.t223 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.VD3.t15 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X254 two_stage_opamp_dummy_magic_0.VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 two_stage_opamp_dummy_magic_0.VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 two_stage_opamp_dummy_magic_0.VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 bgr_0.V_TOP.t25 VDDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 GNDA.t109 GNDA.t126 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X259 two_stage_opamp_dummy_magic_0.VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 two_stage_opamp_dummy_magic_0.VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 two_stage_opamp_dummy_magic_0.VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 VDDA.t205 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD4.t15 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X263 two_stage_opamp_dummy_magic_0.VOUT-.t15 two_stage_opamp_dummy_magic_0.X.t23 VDDA.t251 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X264 a_8420_8490.t6 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD3.t10 w_8160_8260.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X265 two_stage_opamp_dummy_magic_0.VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 GNDA.t274 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA.t273 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X268 two_stage_opamp_dummy_magic_0.VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDDA.t99 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t14 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X270 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X271 two_stage_opamp_dummy_magic_0.VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 a_14640_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t333 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X273 VDDA.t101 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X274 two_stage_opamp_dummy_magic_0.VD1.t14 a_10530_5140# two_stage_opamp_dummy_magic_0.Y.t5 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X275 two_stage_opamp_dummy_magic_0.VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X277 bgr_0.V_mir2.t11 bgr_0.V_mir2.t10 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X278 VDDA.t294 bgr_0.V_TOP.t26 bgr_0.Vin-.t5 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X279 GNDA.t76 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X280 VDDA.t396 VDDA.t394 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X281 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 bgr_0.PFET_GATE_10uA.t18 VDDA.t228 VDDA.t227 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X282 bgr_0.TAIL_CUR_MIR_BIAS.t2 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X283 two_stage_opamp_dummy_magic_0.V_p.t10 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X284 two_stage_opamp_dummy_magic_0.VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 VDDA.t391 VDDA.t393 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=1.28 ps=7.2 w=3.2 l=0.2
X286 VDDA.t252 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X287 two_stage_opamp_dummy_magic_0.VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 two_stage_opamp_dummy_magic_0.VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 bgr_0.Vin-.t1 a_12828_17650.t0 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X290 two_stage_opamp_dummy_magic_0.VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 two_stage_opamp_dummy_magic_0.VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 two_stage_opamp_dummy_magic_0.VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 GNDA.t101 GNDA.t139 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X294 two_stage_opamp_dummy_magic_0.V_p.t19 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X295 a_8420_8490.t5 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.VD3.t6 w_8160_8260.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X296 VDDA.t447 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.VD4.t21 VDDA.t446 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X297 GNDA.t272 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 VDDA.t253 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X298 two_stage_opamp_dummy_magic_0.VD3.t20 VDDA.t388 VDDA.t390 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X299 GNDA.t40 two_stage_opamp_dummy_magic_0.X.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X300 two_stage_opamp_dummy_magic_0.VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 two_stage_opamp_dummy_magic_0.VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_0.VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 GNDA.t276 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X305 bgr_0.PFET_GATE_10uA.t8 bgr_0.1st_Vout_2.t19 VDDA.t439 VDDA.t438 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X306 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t1 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X307 two_stage_opamp_dummy_magic_0.VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 two_stage_opamp_dummy_magic_0.VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA.t140 GNDA.t142 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X310 GNDA.t138 GNDA.t136 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X311 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t0 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X312 two_stage_opamp_dummy_magic_0.Vb2.t6 bgr_0.NFET_GATE_10uA.t12 GNDA.t198 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X313 bgr_0.START_UP.t5 bgr_0.START_UP.t4 bgr_0.START_UP_NFET1.t0 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X314 two_stage_opamp_dummy_magic_0.VOUT+.t9 two_stage_opamp_dummy_magic_0.Y.t24 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X315 two_stage_opamp_dummy_magic_0.VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 two_stage_opamp_dummy_magic_0.VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_0.VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 two_stage_opamp_dummy_magic_0.VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 two_stage_opamp_dummy_magic_0.VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 two_stage_opamp_dummy_magic_0.VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 two_stage_opamp_dummy_magic_0.VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 two_stage_opamp_dummy_magic_0.VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 GNDA.t200 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X324 bgr_0.V_p_1.t3 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t7 GNDA.t265 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X325 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X326 two_stage_opamp_dummy_magic_0.Vb2.t5 bgr_0.NFET_GATE_10uA.t14 GNDA.t42 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X327 two_stage_opamp_dummy_magic_0.VOUT+.t1 GNDA.t133 GNDA.t135 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X328 two_stage_opamp_dummy_magic_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t15 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X329 two_stage_opamp_dummy_magic_0.VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.Vb2.t17 a_10480_8490.t11 w_10220_8260.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X331 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 two_stage_opamp_dummy_magic_0.VOUT-.t4 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X333 two_stage_opamp_dummy_magic_0.VOUT-.t0 two_stage_opamp_dummy_magic_0.X.t28 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X334 VDDA.t238 two_stage_opamp_dummy_magic_0.Y.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X335 bgr_0.Vin+.t5 bgr_0.V_TOP.t27 VDDA.t292 VDDA.t291 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X336 two_stage_opamp_dummy_magic_0.VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 two_stage_opamp_dummy_magic_0.VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 two_stage_opamp_dummy_magic_0.VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VDDA.t93 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X340 two_stage_opamp_dummy_magic_0.VOUT-.t3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X341 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.Vb3.t17 VDDA.t246 VDDA.t245 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X342 VDDA.t445 bgr_0.PFET_GATE_10uA.t19 bgr_0.TAIL_CUR_MIR_BIAS.t9 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X343 two_stage_opamp_dummy_magic_0.VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 bgr_0.TAIL_CUR_MIR_BIAS.t8 bgr_0.PFET_GATE_10uA.t20 VDDA.t461 VDDA.t460 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X345 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t0 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X346 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 a_9610_5930.t6 GNDA.t304 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X347 two_stage_opamp_dummy_magic_0.VD1.t13 a_10530_5140# two_stage_opamp_dummy_magic_0.Y.t11 GNDA.t244 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X348 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t0 GNDA.t0 sky130_fd_pr__res_high_po_1p41 l=1.41
X349 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_p.t5 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X350 two_stage_opamp_dummy_magic_0.VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GNDA.t330 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X352 two_stage_opamp_dummy_magic_0.VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 two_stage_opamp_dummy_magic_0.VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 two_stage_opamp_dummy_magic_0.VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 bgr_0.V_TOP.t28 VDDA.t288 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 bgr_0.Vin+.t0 a_12828_17530.t0 GNDA.t29 sky130_fd_pr__res_xhigh_po_0p35 l=6
X357 two_stage_opamp_dummy_magic_0.V_p.t12 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X358 two_stage_opamp_dummy_magic_0.VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 GNDA.t132 GNDA.t130 GNDA.t132 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X360 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.Vb3.t18 VDDA.t82 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X361 VDDA.t11 two_stage_opamp_dummy_magic_0.X.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X362 two_stage_opamp_dummy_magic_0.VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA.t127 GNDA.t129 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X365 GNDA.t125 GNDA.t123 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 GNDA.t124 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X366 two_stage_opamp_dummy_magic_0.Vb3.t5 bgr_0.NFET_GATE_10uA.t16 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X367 GNDA.t13 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X368 two_stage_opamp_dummy_magic_0.V_p.t13 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X369 bgr_0.V_mir1.t7 bgr_0.V_mir1.t6 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X370 GNDA.t228 two_stage_opamp_dummy_magic_0.X.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X371 a_5230_5088.t1 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t325 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X372 two_stage_opamp_dummy_magic_0.VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 two_stage_opamp_dummy_magic_0.VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t5 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X375 two_stage_opamp_dummy_magic_0.VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 bgr_0.V_p_2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 bgr_0.V_mir2.t0 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X377 two_stage_opamp_dummy_magic_0.VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VDDA.t178 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.Vb1.t3 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X379 two_stage_opamp_dummy_magic_0.VD2.t14 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.X.t7 GNDA.t206 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X380 two_stage_opamp_dummy_magic_0.VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 two_stage_opamp_dummy_magic_0.VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 two_stage_opamp_dummy_magic_0.VOUT+.t8 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t467 VDDA.t466 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X383 two_stage_opamp_dummy_magic_0.VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t216 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X385 bgr_0.V_p_1.t2 bgr_0.Vin+.t8 bgr_0.1st_Vout_1.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X386 two_stage_opamp_dummy_magic_0.VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t287 bgr_0.V_TOP.t29 bgr_0.START_UP.t2 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X388 two_stage_opamp_dummy_magic_0.V_err_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X389 two_stage_opamp_dummy_magic_0.VOUT+.t3 a_14240_2276.t0 GNDA.t188 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X390 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.Vb2.t18 a_8420_8490.t4 w_8160_8260.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X391 two_stage_opamp_dummy_magic_0.VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t61 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X394 two_stage_opamp_dummy_magic_0.VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 two_stage_opamp_dummy_magic_0.VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 two_stage_opamp_dummy_magic_0.Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X397 a_14520_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t328 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X398 bgr_0.V_p_2.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 bgr_0.V_mir2.t16 GNDA.t282 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X399 two_stage_opamp_dummy_magic_0.VOUT-.t11 two_stage_opamp_dummy_magic_0.X.t31 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X400 two_stage_opamp_dummy_magic_0.VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VDDA.t169 two_stage_opamp_dummy_magic_0.Y.t28 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X402 two_stage_opamp_dummy_magic_0.VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VDDA.t89 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t12 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X405 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_0.V_err_p.t4 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X406 two_stage_opamp_dummy_magic_0.err_amp_out.t0 GNDA.t120 GNDA.t122 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X407 two_stage_opamp_dummy_magic_0.VD1.t12 a_10530_5140# two_stage_opamp_dummy_magic_0.Y.t9 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X408 GNDA.t254 two_stage_opamp_dummy_magic_0.Y.t29 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 VDDA.t225 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X409 two_stage_opamp_dummy_magic_0.VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 two_stage_opamp_dummy_magic_0.VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VDDA.t232 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t231 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0.64 ps=3.6 w=3.2 l=0.2
X412 GNDA.t335 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 VDDA.t462 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X413 two_stage_opamp_dummy_magic_0.VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 two_stage_opamp_dummy_magic_0.V_p.t6 a_11120_2960# GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X415 VDDA.t46 two_stage_opamp_dummy_magic_0.X.t32 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X416 two_stage_opamp_dummy_magic_0.V_p.t3 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t2 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X417 bgr_0.1st_Vout_1.t4 bgr_0.V_mir1.t20 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X418 VDDA.t140 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t11 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X419 VDDA.t47 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X420 GNDA.t298 VDDA.t469 bgr_0.V_TOP.t12 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X421 two_stage_opamp_dummy_magic_0.VD4.t1 two_stage_opamp_dummy_magic_0.Vb3.t21 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X422 two_stage_opamp_dummy_magic_0.VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 a_10480_8490.t0 w_10220_8260.t0 w_10220_8260.t2 w_10220_8260.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X424 a_9610_5930.t3 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t9 GNDA.t303 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X425 two_stage_opamp_dummy_magic_0.VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 two_stage_opamp_dummy_magic_0.VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 bgr_0.1st_Vout_2.t3 bgr_0.V_mir2.t19 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X428 two_stage_opamp_dummy_magic_0.VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 two_stage_opamp_dummy_magic_0.VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 two_stage_opamp_dummy_magic_0.VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_0.VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 GNDA.t264 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 two_stage_opamp_dummy_magic_0.VOUT-.t14 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X435 VDDA.t197 bgr_0.PFET_GATE_10uA.t22 bgr_0.TAIL_CUR_MIR_BIAS.t7 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X436 two_stage_opamp_dummy_magic_0.VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X438 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 two_stage_opamp_dummy_magic_0.VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 bgr_0.V_TOP.t30 VDDA.t285 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t2 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X442 two_stage_opamp_dummy_magic_0.VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 bgr_0.START_UP.t1 bgr_0.V_TOP.t31 VDDA.t284 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X444 two_stage_opamp_dummy_magic_0.VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 two_stage_opamp_dummy_magic_0.VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 two_stage_opamp_dummy_magic_0.VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 two_stage_opamp_dummy_magic_0.VD2.t19 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t10 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X448 two_stage_opamp_dummy_magic_0.VOUT+.t7 two_stage_opamp_dummy_magic_0.Y.t31 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X449 two_stage_opamp_dummy_magic_0.VOUT+.t6 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t465 VDDA.t464 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X450 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 bgr_0.V_mir2.t9 bgr_0.V_mir2.t8 VDDA.t176 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X452 two_stage_opamp_dummy_magic_0.VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 two_stage_opamp_dummy_magic_0.VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 a_10480_8490.t10 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD4.t13 w_10220_8260.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X455 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X457 two_stage_opamp_dummy_magic_0.VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 bgr_0.V_TOP.t10 bgr_0.1st_Vout_1.t27 VDDA.t219 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X459 two_stage_opamp_dummy_magic_0.VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 two_stage_opamp_dummy_magic_0.VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 two_stage_opamp_dummy_magic_0.VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 GNDA.t119 GNDA.t116 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X464 GNDA.t96 GNDA.t114 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X465 bgr_0.V_mir2.t7 bgr_0.V_mir2.t6 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X466 VDDA.t282 bgr_0.V_TOP.t32 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X467 GNDA.t316 bgr_0.TAIL_CUR_MIR_BIAS.t23 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X468 VDDA.t102 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X469 two_stage_opamp_dummy_magic_0.VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 two_stage_opamp_dummy_magic_0.VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 VDDA.t387 VDDA.t385 bgr_0.V_TOP.t6 VDDA.t386 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X472 two_stage_opamp_dummy_magic_0.V_err_gate.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X473 two_stage_opamp_dummy_magic_0.VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VDDA.t146 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X475 two_stage_opamp_dummy_magic_0.VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 bgr_0.V_TOP.t33 VDDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 VDDA.t74 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.VD3.t0 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X478 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 VDDA.t382 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X479 GNDA.t297 VDDA.t379 VDDA.t381 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X480 two_stage_opamp_dummy_magic_0.V_p.t28 bgr_0.TAIL_CUR_MIR_BIAS.t24 GNDA.t19 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X481 two_stage_opamp_dummy_magic_0.VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 two_stage_opamp_dummy_magic_0.VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 two_stage_opamp_dummy_magic_0.VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 GNDA.t109 GNDA.t113 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X485 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 two_stage_opamp_dummy_magic_0.V_p.t7 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X487 bgr_0.V_TOP.t34 VDDA.t279 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 VDDA.t7 two_stage_opamp_dummy_magic_0.X.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X489 two_stage_opamp_dummy_magic_0.VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 two_stage_opamp_dummy_magic_0.V_p.t9 two_stage_opamp_dummy_magic_0.Vb1.t1 two_stage_opamp_dummy_magic_0.Vb1.t2 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=2.9
X491 two_stage_opamp_dummy_magic_0.VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 bgr_0.PFET_GATE_10uA.t9 bgr_0.1st_Vout_2.t26 VDDA.t441 VDDA.t440 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X493 a_13790_17550.t1 bgr_0.V_CUR_REF_REG.t1 GNDA.t178 sky130_fd_pr__res_xhigh_po_0p35 l=6
X494 a_9610_5930.t5 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X495 two_stage_opamp_dummy_magic_0.VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VDDA.t39 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X497 VDDA.t278 bgr_0.V_TOP.t35 bgr_0.Vin+.t4 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X498 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 VDDA.t376 VDDA.t378 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X499 a_5350_5088.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t25 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X500 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 two_stage_opamp_dummy_magic_0.VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 GNDA.t296 VDDA.t470 bgr_0.V_p_2.t5 GNDA.t295 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X503 two_stage_opamp_dummy_magic_0.VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 a_9610_5930.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 GNDA.t301 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X505 two_stage_opamp_dummy_magic_0.Y.t12 a_10530_5140# two_stage_opamp_dummy_magic_0.VD1.t11 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X506 bgr_0.V_p_1.t7 bgr_0.Vin-.t10 bgr_0.V_mir1.t14 GNDA.t287 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X507 VDDA.t117 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD3.t2 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X508 a_10480_8490.t9 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD4.t12 w_10220_8260.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X509 two_stage_opamp_dummy_magic_0.VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 two_stage_opamp_dummy_magic_0.VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 bgr_0.V_TOP.t1 bgr_0.1st_Vout_1.t30 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X512 two_stage_opamp_dummy_magic_0.VOUT+.t17 VDDA.t373 VDDA.t375 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X513 two_stage_opamp_dummy_magic_0.VD2.t1 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.X.t2 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X514 two_stage_opamp_dummy_magic_0.VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 bgr_0.V_TOP.t36 VDDA.t276 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 two_stage_opamp_dummy_magic_0.VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 GNDA.t101 GNDA.t115 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X518 two_stage_opamp_dummy_magic_0.VD1.t6 VIN-.t6 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X519 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_2276.t1 GNDA.t332 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X520 bgr_0.1st_Vout_1.t5 bgr_0.V_mir1.t21 VDDA.t152 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X521 two_stage_opamp_dummy_magic_0.VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 two_stage_opamp_dummy_magic_0.VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 two_stage_opamp_dummy_magic_0.VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 two_stage_opamp_dummy_magic_0.VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 two_stage_opamp_dummy_magic_0.VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 two_stage_opamp_dummy_magic_0.VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 two_stage_opamp_dummy_magic_0.VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 bgr_0.Vin+.t3 bgr_0.V_TOP.t37 VDDA.t275 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X529 bgr_0.V_mir2.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t1 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X530 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X531 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 bgr_0.PFET_GATE_10uA.t4 VDDA.t471 GNDA.t294 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X533 two_stage_opamp_dummy_magic_0.VD1.t18 VIN-.t7 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA.t249 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X534 two_stage_opamp_dummy_magic_0.VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 two_stage_opamp_dummy_magic_0.VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 two_stage_opamp_dummy_magic_0.VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 VDDA.t429 two_stage_opamp_dummy_magic_0.Y.t34 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X539 two_stage_opamp_dummy_magic_0.VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 GNDA.t112 GNDA.t110 bgr_0.NFET_GATE_10uA.t0 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X541 two_stage_opamp_dummy_magic_0.VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 GNDA.t5 bgr_0.TAIL_CUR_MIR_BIAS.t25 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X543 two_stage_opamp_dummy_magic_0.V_err_gate.t8 bgr_0.NFET_GATE_10uA.t18 GNDA.t209 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X544 bgr_0.1st_Vout_1.t1 bgr_0.Vin+.t9 bgr_0.V_p_1.t1 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X545 VDDA.t83 two_stage_opamp_dummy_magic_0.Y.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X546 VDDA.t372 VDDA.t370 VDDA.t372 VDDA.t371 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0 ps=0 w=3.2 l=0.2
X547 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t36 sky130_fd_pr__res_high_po_1p41 l=1.41
X548 bgr_0.V_TOP.t2 bgr_0.1st_Vout_1.t31 VDDA.t80 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X549 two_stage_opamp_dummy_magic_0.VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 two_stage_opamp_dummy_magic_0.VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 bgr_0.PFET_GATE_10uA.t24 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X552 two_stage_opamp_dummy_magic_0.VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_0.VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 bgr_0.Vin-.t6 bgr_0.V_TOP.t38 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X555 VDDA.t443 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 VDDA.t442 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X556 VDDA.t369 VDDA.t367 two_stage_opamp_dummy_magic_0.VD4.t18 VDDA.t368 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X557 two_stage_opamp_dummy_magic_0.VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 two_stage_opamp_dummy_magic_0.V_p.t26 bgr_0.TAIL_CUR_MIR_BIAS.t26 GNDA.t232 GNDA.t231 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X559 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.Vb2.t22 a_10480_8490.t8 w_10220_8260.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X560 two_stage_opamp_dummy_magic_0.VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 a_13790_17550.t0 GNDA.t179 GNDA.t178 sky130_fd_pr__res_xhigh_po_0p35 l=6
X562 two_stage_opamp_dummy_magic_0.VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 two_stage_opamp_dummy_magic_0.VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 bgr_0.V_TOP.t11 VDDA.t364 VDDA.t366 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X565 a_9610_5930.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA.t300 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X566 VDDA.t363 VDDA.t361 two_stage_opamp_dummy_magic_0.VD3.t19 VDDA.t362 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X567 two_stage_opamp_dummy_magic_0.VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 two_stage_opamp_dummy_magic_0.VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 two_stage_opamp_dummy_magic_0.VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 GNDA.t293 VDDA.t358 VDDA.t360 VDDA.t359 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X571 bgr_0.V_TOP.t39 VDDA.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 two_stage_opamp_dummy_magic_0.VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 two_stage_opamp_dummy_magic_0.VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 bgr_0.NFET_GATE_10uA.t19 GNDA.t211 GNDA.t210 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X575 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 bgr_0.NFET_GATE_10uA.t20 GNDA.t215 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X576 two_stage_opamp_dummy_magic_0.VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 two_stage_opamp_dummy_magic_0.VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 VDDA.t54 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t2 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X580 VDDA.t357 VDDA.t355 two_stage_opamp_dummy_magic_0.err_amp_out.t6 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X581 two_stage_opamp_dummy_magic_0.Y.t8 a_10530_5140# two_stage_opamp_dummy_magic_0.VD1.t10 GNDA.t241 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X582 two_stage_opamp_dummy_magic_0.VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 bgr_0.V_TOP.t40 VDDA.t270 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 VDDA.t269 bgr_0.V_TOP.t41 bgr_0.Vin+.t2 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X585 VDDA.t354 VDDA.t352 GNDA.t292 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X586 two_stage_opamp_dummy_magic_0.VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 two_stage_opamp_dummy_magic_0.VD2.t16 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.X.t9 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X588 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.Vb2.t23 a_10480_8490.t7 w_10220_8260.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X589 bgr_0.V_mir1.t3 bgr_0.V_mir1.t2 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X590 two_stage_opamp_dummy_magic_0.VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 bgr_0.NFET_GATE_10uA.t21 GNDA.t217 GNDA.t216 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X592 a_8420_8490.t3 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.VD3.t9 w_8160_8260.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X593 GNDA.t109 GNDA.t108 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X594 bgr_0.V_mir2.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 bgr_0.V_p_2.t0 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X595 bgr_0.PFET_GATE_10uA.t6 VDDA.t349 VDDA.t351 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X596 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_0.X.t35 GNDA.t7 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X597 two_stage_opamp_dummy_magic_0.VD2.t3 VIN+.t7 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X598 two_stage_opamp_dummy_magic_0.VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 two_stage_opamp_dummy_magic_0.VOUT-.t18 VDDA.t346 VDDA.t348 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X600 VDDA.t16 GNDA.t105 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X601 two_stage_opamp_dummy_magic_0.VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 GNDA.t262 bgr_0.TAIL_CUR_MIR_BIAS.t27 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA.t261 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X603 two_stage_opamp_dummy_magic_0.V_err_gate.t10 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X604 two_stage_opamp_dummy_magic_0.VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 VDDA.t345 VDDA.t343 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X606 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t242 VDDA.t241 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X607 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.Vb2.t25 a_10480_8490.t6 w_10220_8260.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X608 two_stage_opamp_dummy_magic_0.VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 bgr_0.V_TOP.t42 VDDA.t267 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 bgr_0.TAIL_CUR_MIR_BIAS.t6 bgr_0.PFET_GATE_10uA.t26 VDDA.t453 VDDA.t452 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X611 two_stage_opamp_dummy_magic_0.VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 two_stage_opamp_dummy_magic_0.VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 two_stage_opamp_dummy_magic_0.X.t12 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA.t336 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X614 VDDA.t342 VDDA.t340 two_stage_opamp_dummy_magic_0.VOUT+.t16 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X615 two_stage_opamp_dummy_magic_0.VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 bgr_0.1st_Vout_2.t1 bgr_0.V_mir2.t21 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X617 two_stage_opamp_dummy_magic_0.VOUT+.t14 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA.t194 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X618 two_stage_opamp_dummy_magic_0.V_p.t24 bgr_0.TAIL_CUR_MIR_BIAS.t28 GNDA.t281 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X619 VDDA.t339 VDDA.t336 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X620 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 a_5350_5088.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA.t331 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X622 GNDA.t101 GNDA.t100 bgr_0.Vin-.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X623 two_stage_opamp_dummy_magic_0.VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 GNDA.t251 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA.t250 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X625 two_stage_opamp_dummy_magic_0.VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_0.VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X627 VDDA.t27 two_stage_opamp_dummy_magic_0.X.t36 two_stage_opamp_dummy_magic_0.VOUT-.t2 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X628 two_stage_opamp_dummy_magic_0.VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 two_stage_opamp_dummy_magic_0.VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 two_stage_opamp_dummy_magic_0.V_p.t23 bgr_0.TAIL_CUR_MIR_BIAS.t29 GNDA.t35 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X631 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 bgr_0.V_TOP.t43 VDDA.t266 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X632 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t333 VDDA.t335 VDDA.t334 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X634 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.Vb2.t26 a_10480_8490.t5 w_10220_8260.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X635 two_stage_opamp_dummy_magic_0.VD3.t21 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t433 VDDA.t432 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X636 two_stage_opamp_dummy_magic_0.V_err_p.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X637 two_stage_opamp_dummy_magic_0.VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 two_stage_opamp_dummy_magic_0.VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 two_stage_opamp_dummy_magic_0.Y.t3 a_10530_5140# two_stage_opamp_dummy_magic_0.VD1.t9 GNDA.t240 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X640 two_stage_opamp_dummy_magic_0.VOUT+.t15 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA.t224 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X641 VDDA.t427 bgr_0.1st_Vout_2.t32 bgr_0.PFET_GATE_10uA.t7 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X642 VDDA.t332 VDDA.t330 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t331 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X643 two_stage_opamp_dummy_magic_0.VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 two_stage_opamp_dummy_magic_0.Vb1.t4 VDDA.t327 VDDA.t329 VDDA.t328 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X645 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X646 two_stage_opamp_dummy_magic_0.VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t36 GNDA.t309 VDDA.t428 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X648 two_stage_opamp_dummy_magic_0.VD2.t10 VIN+.t8 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X649 GNDA.t104 GNDA.t102 bgr_0.TAIL_CUR_MIR_BIAS.t0 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X650 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 two_stage_opamp_dummy_magic_0.VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 two_stage_opamp_dummy_magic_0.VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 two_stage_opamp_dummy_magic_0.VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 two_stage_opamp_dummy_magic_0.VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 bgr_0.V_mir1.t15 bgr_0.Vin-.t11 bgr_0.V_p_1.t6 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X657 two_stage_opamp_dummy_magic_0.VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 two_stage_opamp_dummy_magic_0.VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 two_stage_opamp_dummy_magic_0.VD2.t9 VIN+.t9 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X660 two_stage_opamp_dummy_magic_0.VD4.t0 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t43 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X661 two_stage_opamp_dummy_magic_0.VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 two_stage_opamp_dummy_magic_0.X.t37 GNDA.t15 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X663 VDDA.t326 VDDA.t324 GNDA.t291 VDDA.t325 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X664 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 GNDA.t63 bgr_0.TAIL_CUR_MIR_BIAS.t30 two_stage_opamp_dummy_magic_0.V_p_mir.t2 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X666 two_stage_opamp_dummy_magic_0.V_err_gate.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X667 VDDA.t323 VDDA.t321 two_stage_opamp_dummy_magic_0.Vb2.t10 VDDA.t322 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X668 a_10480_8490.t4 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD4.t8 w_10220_8260.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X669 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X670 VDDA.t431 two_stage_opamp_dummy_magic_0.Y.t37 two_stage_opamp_dummy_magic_0.VOUT+.t5 VDDA.t430 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X671 GNDA.t253 bgr_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X672 VDDA.t264 bgr_0.V_TOP.t44 bgr_0.START_UP.t0 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X673 two_stage_opamp_dummy_magic_0.VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.Vb2.t28 a_8420_8490.t2 w_8160_8260.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X675 two_stage_opamp_dummy_magic_0.VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 two_stage_opamp_dummy_magic_0.V_p.t22 bgr_0.TAIL_CUR_MIR_BIAS.t31 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X677 VDDA.t224 GNDA.t97 GNDA.t99 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X678 two_stage_opamp_dummy_magic_0.VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VDDA.t65 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X680 two_stage_opamp_dummy_magic_0.VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 GNDA.t96 GNDA.t95 bgr_0.Vbe2.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X682 two_stage_opamp_dummy_magic_0.VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 two_stage_opamp_dummy_magic_0.VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 VDDA.t185 two_stage_opamp_dummy_magic_0.X.t38 two_stage_opamp_dummy_magic_0.VOUT-.t10 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X685 VDDA.t320 VDDA.t318 two_stage_opamp_dummy_magic_0.VOUT-.t17 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X686 VDDA.t221 bgr_0.V_mir2.t4 bgr_0.V_mir2.t5 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X687 VDDA.t138 bgr_0.PFET_GATE_10uA.t27 bgr_0.TAIL_CUR_MIR_BIAS.t5 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X688 two_stage_opamp_dummy_magic_0.VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 GNDA.t94 GNDA.t92 VDDA.t128 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X691 bgr_0.TAIL_CUR_MIR_BIAS.t4 bgr_0.PFET_GATE_10uA.t28 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X692 two_stage_opamp_dummy_magic_0.VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 bgr_0.V_TOP.t45 VDDA.t262 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 two_stage_opamp_dummy_magic_0.V_err_p.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X695 bgr_0.1st_Vout_1.t3 bgr_0.V_mir1.t22 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X696 two_stage_opamp_dummy_magic_0.Y.t6 a_10530_5140# two_stage_opamp_dummy_magic_0.VD1.t8 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X697 two_stage_opamp_dummy_magic_0.VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 two_stage_opamp_dummy_magic_0.V_err_p.t19 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 VDDA.t235 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X699 two_stage_opamp_dummy_magic_0.V_err_p.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t2 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X700 two_stage_opamp_dummy_magic_0.VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_0.Y.t38 GNDA.t222 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X702 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 bgr_0.1st_Vout_2.t6 bgr_0.V_CUR_REF_REG.t6 bgr_0.V_p_2.t6 GNDA.t310 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X704 bgr_0.V_TOP.t46 VDDA.t261 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.Vb2.t29 a_8420_8490.t1 w_8160_8260.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X706 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_0.X.t39 VDDA.t186 GNDA.t227 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X707 two_stage_opamp_dummy_magic_0.V_p_mir.t1 VIN-.t8 bgr_0.TAIL_CUR_MIR_BIAS.t3 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X708 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t9 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X709 two_stage_opamp_dummy_magic_0.VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X710 two_stage_opamp_dummy_magic_0.VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 two_stage_opamp_dummy_magic_0.VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 two_stage_opamp_dummy_magic_0.VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 bgr_0.V_p_1.t10 VDDA.t472 GNDA.t290 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X714 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 bgr_0.V_mir1.t16 bgr_0.Vin-.t12 bgr_0.V_p_1.t5 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X716 VDDA.t317 VDDA.t315 bgr_0.PFET_GATE_10uA.t5 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X717 two_stage_opamp_dummy_magic_0.VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 two_stage_opamp_dummy_magic_0.VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 GNDA.t58 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 two_stage_opamp_dummy_magic_0.VOUT-.t5 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X720 two_stage_opamp_dummy_magic_0.VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 two_stage_opamp_dummy_magic_0.VD1.t1 VIN-.t10 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X722 a_10480_8490.t3 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.VD4.t7 w_10220_8260.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X723 bgr_0.V_TOP.t47 VDDA.t260 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X724 VDDA.t234 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD3.t16 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X725 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 two_stage_opamp_dummy_magic_0.X.t40 GNDA.t189 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X726 VDDA.t106 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X727 two_stage_opamp_dummy_magic_0.VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 two_stage_opamp_dummy_magic_0.VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 GNDA.t327 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 two_stage_opamp_dummy_magic_0.VOUT+.t18 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X730 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 bgr_0.V_TOP.t48 VDDA.t259 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X731 bgr_0.V_TOP.t8 bgr_0.START_UP.t7 bgr_0.Vin-.t3 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X732 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t312 VDDA.t314 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X733 two_stage_opamp_dummy_magic_0.VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 bgr_0.1st_Vout_2.t10 bgr_0.V_CUR_REF_REG.t7 bgr_0.V_p_2.t10 GNDA.t318 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X735 two_stage_opamp_dummy_magic_0.V_err_gate.t13 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 VDDA.t450 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X736 two_stage_opamp_dummy_magic_0.VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VDDA.t72 bgr_0.1st_Vout_2.t36 bgr_0.PFET_GATE_10uA.t1 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X738 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t329 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X740 two_stage_opamp_dummy_magic_0.Vb2.t3 two_stage_opamp_dummy_magic_0.Vb2.t2 VDDA.t174 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X741 VDDA.t113 two_stage_opamp_dummy_magic_0.Y.t39 two_stage_opamp_dummy_magic_0.VOUT+.t4 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X742 two_stage_opamp_dummy_magic_0.VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 a_5230_5088.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t24 sky130_fd_pr__res_xhigh_po_0p35 l=1.85
X744 two_stage_opamp_dummy_magic_0.VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 two_stage_opamp_dummy_magic_0.VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 GNDA.t91 GNDA.t89 two_stage_opamp_dummy_magic_0.VOUT-.t7 GNDA.t90 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X747 two_stage_opamp_dummy_magic_0.VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_0.VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 two_stage_opamp_dummy_magic_0.VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 two_stage_opamp_dummy_magic_0.VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VDDA.t25 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t8 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X752 a_8420_8490.t0 w_8160_8260.t0 w_8160_8260.t2 w_8160_8260.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X753 two_stage_opamp_dummy_magic_0.VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_0.VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VDDA.t311 VDDA.t309 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X756 two_stage_opamp_dummy_magic_0.VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 bgr_0.PFET_GATE_10uA.t29 VDDA.t435 VDDA.t434 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X758 a_10480_8490.t2 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD4.t9 w_10220_8260.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X759 two_stage_opamp_dummy_magic_0.VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VDDA.t20 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X761 VDDA.t126 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.VOUT-.t9 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X762 two_stage_opamp_dummy_magic_0.VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 two_stage_opamp_dummy_magic_0.VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_0.Y.t40 VDDA.t463 GNDA.t338 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X765 two_stage_opamp_dummy_magic_0.VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X767 two_stage_opamp_dummy_magic_0.VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t86 GNDA.t88 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X769 two_stage_opamp_dummy_magic_0.V_err_p.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X770 a_9610_5930.t2 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X771 two_stage_opamp_dummy_magic_0.VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 two_stage_opamp_dummy_magic_0.Y.t41 GNDA.t256 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X773 two_stage_opamp_dummy_magic_0.VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 two_stage_opamp_dummy_magic_0.VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 two_stage_opamp_dummy_magic_0.VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 two_stage_opamp_dummy_magic_0.Y.t42 GNDA.t257 VDDA.t237 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X777 two_stage_opamp_dummy_magic_0.VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 bgr_0.V_TOP.t49 VDDA.t257 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 bgr_0.1st_Vout_1.t6 bgr_0.Vin+.t10 bgr_0.V_p_1.t0 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X780 GNDA.t322 two_stage_opamp_dummy_magic_0.err_amp_out.t12 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X781 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t83 GNDA.t85 GNDA.t84 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X782 two_stage_opamp_dummy_magic_0.VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_0.X.t42 VDDA.t119 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X784 GNDA.t82 GNDA.t80 VDDA.t85 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X785 two_stage_opamp_dummy_magic_0.VD2.t18 VIN+.t10 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X786 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5750_2276.t1 GNDA.t323 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X787 bgr_0.Vin+.t1 bgr_0.Vbe2.t8 GNDA.t238 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X788 VDDA.t108 two_stage_opamp_dummy_magic_0.Vb3.t28 two_stage_opamp_dummy_magic_0.VD4.t2 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X789 two_stage_opamp_dummy_magic_0.VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.V_TOP.n0 bgr_0.V_TOP.t43 369.534
R1 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 339.961
R2 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 339.272
R3 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R4 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R5 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R6 bgr_0.V_TOP.n12 bgr_0.V_TOP.n8 334.772
R7 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R8 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R9 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R10 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R11 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R12 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R13 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R14 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R15 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R16 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R17 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R18 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R19 bgr_0.V_TOP bgr_0.V_TOP.t32 214.222
R20 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R21 bgr_0.V_TOP.n7 bgr_0.V_TOP.t13 176.114
R22 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R23 bgr_0.V_TOP.n27 bgr_0.V_TOP.t31 144.601
R24 bgr_0.V_TOP.n26 bgr_0.V_TOP.t44 144.601
R25 bgr_0.V_TOP.n25 bgr_0.V_TOP.t18 144.601
R26 bgr_0.V_TOP.n24 bgr_0.V_TOP.t26 144.601
R27 bgr_0.V_TOP.n23 bgr_0.V_TOP.t37 144.601
R28 bgr_0.V_TOP.n22 bgr_0.V_TOP.t35 144.601
R29 bgr_0.V_TOP.n21 bgr_0.V_TOP.t48 144.601
R30 bgr_0.V_TOP.n20 bgr_0.V_TOP.t20 144.601
R31 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 144.601
R32 bgr_0.V_TOP.n1 bgr_0.V_TOP.t23 144.601
R33 bgr_0.V_TOP.n2 bgr_0.V_TOP.t14 144.601
R34 bgr_0.V_TOP.n3 bgr_0.V_TOP.t38 144.601
R35 bgr_0.V_TOP.n4 bgr_0.V_TOP.t41 144.601
R36 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R37 bgr_0.V_TOP.n18 bgr_0.V_TOP.t12 95.4466
R38 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R39 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R40 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R41 bgr_0.V_TOP.n6 bgr_0.V_TOP.t5 39.4005
R42 bgr_0.V_TOP.n6 bgr_0.V_TOP.t1 39.4005
R43 bgr_0.V_TOP.n8 bgr_0.V_TOP.t0 39.4005
R44 bgr_0.V_TOP.n8 bgr_0.V_TOP.t2 39.4005
R45 bgr_0.V_TOP.n10 bgr_0.V_TOP.t7 39.4005
R46 bgr_0.V_TOP.n10 bgr_0.V_TOP.t3 39.4005
R47 bgr_0.V_TOP.n9 bgr_0.V_TOP.t6 39.4005
R48 bgr_0.V_TOP.n9 bgr_0.V_TOP.t8 39.4005
R49 bgr_0.V_TOP.n14 bgr_0.V_TOP.t4 39.4005
R50 bgr_0.V_TOP.n14 bgr_0.V_TOP.t10 39.4005
R51 bgr_0.V_TOP.n16 bgr_0.V_TOP.t9 39.4005
R52 bgr_0.V_TOP.n16 bgr_0.V_TOP.t11 39.4005
R53 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 8.313
R54 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R55 bgr_0.V_TOP.n28 bgr_0.V_TOP.t49 4.8295
R56 bgr_0.V_TOP.n29 bgr_0.V_TOP.t25 4.8295
R57 bgr_0.V_TOP.n31 bgr_0.V_TOP.t21 4.8295
R58 bgr_0.V_TOP.n32 bgr_0.V_TOP.t34 4.8295
R59 bgr_0.V_TOP.n34 bgr_0.V_TOP.t30 4.8295
R60 bgr_0.V_TOP.n35 bgr_0.V_TOP.t46 4.8295
R61 bgr_0.V_TOP.n37 bgr_0.V_TOP.t24 4.8295
R62 bgr_0.V_TOP.n28 bgr_0.V_TOP.t39 4.5005
R63 bgr_0.V_TOP.n30 bgr_0.V_TOP.t28 4.5005
R64 bgr_0.V_TOP.n29 bgr_0.V_TOP.t33 4.5005
R65 bgr_0.V_TOP.n31 bgr_0.V_TOP.t15 4.5005
R66 bgr_0.V_TOP.n33 bgr_0.V_TOP.t40 4.5005
R67 bgr_0.V_TOP.n32 bgr_0.V_TOP.t45 4.5005
R68 bgr_0.V_TOP.n34 bgr_0.V_TOP.t22 4.5005
R69 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 4.5005
R70 bgr_0.V_TOP.n35 bgr_0.V_TOP.t19 4.5005
R71 bgr_0.V_TOP.n37 bgr_0.V_TOP.t17 4.5005
R72 bgr_0.V_TOP.n38 bgr_0.V_TOP.t42 4.5005
R73 bgr_0.V_TOP.n39 bgr_0.V_TOP.t47 4.5005
R74 bgr_0.V_TOP.n40 bgr_0.V_TOP.t36 4.5005
R75 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R76 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R77 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R78 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R79 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R80 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R81 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R82 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R83 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R84 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R85 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R86 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R87 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R88 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R89 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R90 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R91 bgr_0.Vin-.n21 bgr_0.Vin-.n20 1850.93
R92 bgr_0.Vin-.n9 bgr_0.Vin-.t10 688.859
R93 bgr_0.Vin-.n11 bgr_0.Vin-.n10 514.134
R94 bgr_0.Vin-.n7 bgr_0.Vin-.n6 345.115
R95 bgr_0.Vin-.n13 bgr_0.Vin-.n12 214.713
R96 bgr_0.Vin-.n9 bgr_0.Vin-.t12 174.726
R97 bgr_0.Vin-.n10 bgr_0.Vin-.t8 174.726
R98 bgr_0.Vin-.n11 bgr_0.Vin-.t11 174.726
R99 bgr_0.Vin-.n12 bgr_0.Vin-.t9 174.726
R100 bgr_0.Vin-.n5 bgr_0.Vin-.n3 173.029
R101 bgr_0.Vin-.n5 bgr_0.Vin-.n4 168.654
R102 bgr_0.Vin-.n7 bgr_0.Vin-.t1 162.921
R103 bgr_0.Vin-.n10 bgr_0.Vin-.n9 128.534
R104 bgr_0.Vin-.n12 bgr_0.Vin-.n11 128.534
R105 bgr_0.Vin-.n22 bgr_0.Vin-.n21 84.0884
R106 bgr_0.Vin-.n17 bgr_0.Vin-.n16 83.5719
R107 bgr_0.Vin-.n18 bgr_0.Vin-.n0 83.5719
R108 bgr_0.Vin-.n19 bgr_0.Vin-.n1 83.5719
R109 bgr_0.Vin-.n14 bgr_0.Vin-.t0 65.0299
R110 bgr_0.Vin-.n6 bgr_0.Vin-.t3 39.4005
R111 bgr_0.Vin-.n6 bgr_0.Vin-.t2 39.4005
R112 bgr_0.Vin-.n18 bgr_0.Vin-.n17 26.074
R113 bgr_0.Vin-.n19 bgr_0.Vin-.n18 26.074
R114 bgr_0.Vin-.n21 bgr_0.Vin-.n19 26.074
R115 bgr_0.Vin-.n23 bgr_0.Vin-.n13 17.526
R116 bgr_0.Vin-.n4 bgr_0.Vin-.t4 13.1338
R117 bgr_0.Vin-.n4 bgr_0.Vin-.t6 13.1338
R118 bgr_0.Vin-.n3 bgr_0.Vin-.t5 13.1338
R119 bgr_0.Vin-.n3 bgr_0.Vin-.t7 13.1338
R120 bgr_0.Vin-.n13 bgr_0.Vin-.n8 12.5317
R121 bgr_0.Vin-.n8 bgr_0.Vin-.n7 6.40675
R122 bgr_0.Vin-.n8 bgr_0.Vin-.n5 3.8755
R123 bgr_0.Vin-.n16 bgr_0.Vin-.n14 1.56363
R124 bgr_0.Vin-.n23 bgr_0.Vin-.n22 1.5505
R125 bgr_0.Vin-.n25 bgr_0.Vin-.n24 1.5505
R126 bgr_0.Vin-.n15 bgr_0.Vin-.n2 1.5505
R127 bgr_0.Vin-.n22 bgr_0.Vin-.n1 1.14402
R128 bgr_0.Vin-.n15 bgr_0.Vin-.n0 0.885803
R129 bgr_0.Vin-.n16 bgr_0.Vin-.n15 0.77514
R130 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.756696
R131 bgr_0.Vin-.n25 bgr_0.Vin-.n1 0.701365
R132 bgr_0.Vin-.n14 bgr_0.Vin-.n2 0.537712
R133 bgr_0.Vin-.n17 bgr_0.Vin-.t0 0.290206
R134 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n25 0.203382
R135 bgr_0.Vin-.n24 bgr_0.Vin-.n2 0.0183571
R136 bgr_0.Vin-.n24 bgr_0.Vin-.n23 0.0183571
R137 VDDA.n376 VDDA.n343 6600
R138 VDDA.n378 VDDA.n343 6600
R139 VDDA.n378 VDDA.n344 6570
R140 VDDA.n376 VDDA.n344 6570
R141 VDDA.n331 VDDA.n266 4710
R142 VDDA.n331 VDDA.n267 4710
R143 VDDA.n333 VDDA.n266 4710
R144 VDDA.n333 VDDA.n267 4710
R145 VDDA.n289 VDDA.n288 4710
R146 VDDA.n291 VDDA.n288 4710
R147 VDDA.n289 VDDA.n282 4710
R148 VDDA.n291 VDDA.n282 4710
R149 VDDA.n143 VDDA.n129 4605
R150 VDDA.n145 VDDA.n129 4605
R151 VDDA.n69 VDDA.n65 4605
R152 VDDA.n69 VDDA.n66 4605
R153 VDDA.n179 VDDA.n175 4590
R154 VDDA.n179 VDDA.n176 4590
R155 VDDA.n181 VDDA.n176 4590
R156 VDDA.n181 VDDA.n175 4590
R157 VDDA.n143 VDDA.n130 4575
R158 VDDA.n145 VDDA.n130 4575
R159 VDDA.n71 VDDA.n65 4575
R160 VDDA.n71 VDDA.n66 4575
R161 VDDA.n205 VDDA.n198 4020
R162 VDDA.n207 VDDA.n198 4020
R163 VDDA.n205 VDDA.n204 4020
R164 VDDA.n207 VDDA.n204 4020
R165 VDDA.n93 VDDA.n86 4020
R166 VDDA.n95 VDDA.n86 4020
R167 VDDA.n93 VDDA.n92 4020
R168 VDDA.n95 VDDA.n92 4020
R169 VDDA.n442 VDDA.n410 3420
R170 VDDA.n442 VDDA.n411 3420
R171 VDDA.n122 VDDA.n115 3390
R172 VDDA.n124 VDDA.n115 3390
R173 VDDA.n122 VDDA.n121 3390
R174 VDDA.n124 VDDA.n121 3390
R175 VDDA.n49 VDDA.n42 3390
R176 VDDA.n51 VDDA.n42 3390
R177 VDDA.n49 VDDA.n48 3390
R178 VDDA.n51 VDDA.n48 3390
R179 VDDA.n23 VDDA.n17 2940
R180 VDDA.n25 VDDA.n17 2940
R181 VDDA.n25 VDDA.n22 2940
R182 VDDA.n23 VDDA.n22 2940
R183 VDDA.n31 VDDA.n12 2940
R184 VDDA.n33 VDDA.n12 2940
R185 VDDA.n33 VDDA.n30 2940
R186 VDDA.n31 VDDA.n30 2940
R187 VDDA.n444 VDDA.n410 2760
R188 VDDA.n444 VDDA.n411 2760
R189 VDDA.n235 VDDA.n224 2415
R190 VDDA.n235 VDDA.n225 2370
R191 VDDA.n232 VDDA.n225 2280
R192 VDDA.n232 VDDA.n224 2235
R193 VDDA.n458 VDDA.n404 2145
R194 VDDA.n458 VDDA.n405 2100
R195 VDDA.n455 VDDA.n405 2100
R196 VDDA.n423 VDDA.n416 2100
R197 VDDA.n425 VDDA.n416 2100
R198 VDDA.n425 VDDA.n417 2100
R199 VDDA.n423 VDDA.n417 2100
R200 VDDA.n455 VDDA.n404 2055
R201 VDDA.n391 VDDA.n389 1770
R202 VDDA.n393 VDDA.n389 1770
R203 VDDA.n391 VDDA.n386 1770
R204 VDDA.n393 VDDA.n386 1770
R205 VDDA.n352 VDDA.n350 1770
R206 VDDA.n354 VDDA.n350 1770
R207 VDDA.n352 VDDA.n347 1770
R208 VDDA.n354 VDDA.n347 1770
R209 VDDA.n247 VDDA.n220 1575
R210 VDDA.n246 VDDA.n220 1575
R211 VDDA.n246 VDDA.n219 1545
R212 VDDA.n247 VDDA.n219 1545
R213 VDDA.n140 VDDA.t340 1216.42
R214 VDDA.n148 VDDA.t373 1216.42
R215 VDDA.n63 VDDA.t346 1216.42
R216 VDDA.n74 VDDA.t318 1216.42
R217 VDDA.n375 VDDA.n342 704
R218 VDDA.n379 VDDA.n342 704
R219 VDDA.n19 VDDA.t357 689.4
R220 VDDA.n18 VDDA.t384 689.4
R221 VDDA.n14 VDDA.t423 689.4
R222 VDDA.n13 VDDA.t314 689.4
R223 VDDA.n172 VDDA.t399 663.801
R224 VDDA.n185 VDDA.t405 663.801
R225 VDDA.n201 VDDA.t361 660.109
R226 VDDA.n199 VDDA.t388 660.109
R227 VDDA.n89 VDDA.t367 660.109
R228 VDDA.n87 VDDA.t412 660.109
R229 VDDA.n242 VDDA.t323 647.54
R230 VDDA.n251 VDDA.t339 647.54
R231 VDDA.n216 VDDA.n215 633.361
R232 VDDA.n152 VDDA.n151 626.534
R233 VDDA.n155 VDDA.n154 626.534
R234 VDDA.n157 VDDA.n156 626.534
R235 VDDA.n159 VDDA.n158 626.534
R236 VDDA.n161 VDDA.n160 626.534
R237 VDDA.n163 VDDA.n162 626.534
R238 VDDA.n165 VDDA.n164 626.534
R239 VDDA.n167 VDDA.n166 626.534
R240 VDDA.n169 VDDA.n168 626.534
R241 VDDA.n171 VDDA.n170 626.534
R242 VDDA.n229 VDDA.t370 623.958
R243 VDDA.n238 VDDA.t391 623.958
R244 VDDA.t370 VDDA.n228 615.926
R245 VDDA.n118 VDDA.t352 573.75
R246 VDDA.n116 VDDA.t379 573.75
R247 VDDA.n45 VDDA.t324 573.75
R248 VDDA.n43 VDDA.t358 573.75
R249 VDDA.n374 VDDA.n341 518.4
R250 VDDA.n380 VDDA.n341 518.4
R251 VDDA.n293 VDDA.n292 496
R252 VDDA.n293 VDDA.n281 496
R253 VDDA.n146 VDDA.n128 491.2
R254 VDDA.n142 VDDA.n128 491.2
R255 VDDA.n68 VDDA.n40 491.2
R256 VDDA.n68 VDDA.n67 491.2
R257 VDDA.n178 VDDA.n153 489.601
R258 VDDA.n178 VDDA.n177 489.601
R259 VDDA.n209 VDDA.n208 428.8
R260 VDDA.n209 VDDA.n197 428.8
R261 VDDA.n97 VDDA.n96 428.8
R262 VDDA.n97 VDDA.n85 428.8
R263 VDDA.n387 VDDA.t327 419.108
R264 VDDA.n384 VDDA.t330 419.108
R265 VDDA.n348 VDDA.t406 413.084
R266 VDDA.n345 VDDA.t385 413.084
R267 VDDA.n452 VDDA.t394 409.067
R268 VDDA.n461 VDDA.t333 409.067
R269 VDDA.n439 VDDA.t415 409.067
R270 VDDA.n447 VDDA.t409 409.067
R271 VDDA.n420 VDDA.t309 409.067
R272 VDDA.n428 VDDA.t376 390.322
R273 VDDA.t404 VDDA.n175 389.375
R274 VDDA.t398 VDDA.n176 389.375
R275 VDDA.t422 VDDA.n30 389.375
R276 VDDA.t313 VDDA.n12 389.375
R277 VDDA.n387 VDDA.t329 389.185
R278 VDDA.n384 VDDA.t332 389.185
R279 VDDA.n183 VDDA.n182 387.2
R280 VDDA.n182 VDDA.n174 387.2
R281 VDDA.n439 VDDA.t417 387.051
R282 VDDA.n447 VDDA.t411 387.051
R283 VDDA.n264 VDDA.t351 384.918
R284 VDDA.n268 VDDA.t317 384.918
R285 VDDA.n283 VDDA.t366 384.918
R286 VDDA.n285 VDDA.t420 384.918
R287 VDDA.n348 VDDA.t408 384.918
R288 VDDA.n345 VDDA.t387 384.918
R289 VDDA.t356 VDDA.n22 384.168
R290 VDDA.t383 VDDA.n17 384.168
R291 VDDA.n270 VDDA.n269 384
R292 VDDA.n269 VDDA.n265 384
R293 VDDA.n287 VDDA.n286 384
R294 VDDA.n287 VDDA.n284 384
R295 VDDA.n420 VDDA.t311 370.728
R296 VDDA.n428 VDDA.t378 370.728
R297 VDDA.n452 VDDA.t396 370.3
R298 VDDA.n461 VDDA.t335 370.3
R299 VDDA.n441 VDDA.n409 364.8
R300 VDDA.n373 VDDA.t343 360.868
R301 VDDA.n381 VDDA.t400 360.868
R302 VDDA.n264 VDDA.t349 358.858
R303 VDDA.n268 VDDA.t315 358.858
R304 VDDA.n283 VDDA.t364 358.858
R305 VDDA.n285 VDDA.t418 358.858
R306 VDDA.n126 VDDA.n125 355.2
R307 VDDA.n126 VDDA.n114 355.2
R308 VDDA.n53 VDDA.n52 355.2
R309 VDDA.n53 VDDA.n41 355.2
R310 VDDA.t316 VDDA.n331 351.591
R311 VDDA.n333 VDDA.t350 351.591
R312 VDDA.t419 VDDA.n289 351.591
R313 VDDA.n291 VDDA.t365 351.591
R314 VDDA.t322 VDDA.n246 346.668
R315 VDDA.n247 VDDA.t337 346.668
R316 VDDA.n413 VDDA.n412 345.127
R317 VDDA.n419 VDDA.n418 345.127
R318 VDDA.n401 VDDA.n400 344.7
R319 VDDA.n450 VDDA.n449 344.7
R320 VDDA.t331 VDDA.n391 344.394
R321 VDDA.n393 VDDA.t328 344.394
R322 VDDA.t386 VDDA.n352 344.394
R323 VDDA.n354 VDDA.t407 344.394
R324 VDDA.t395 VDDA.n455 344.394
R325 VDDA.n458 VDDA.t334 344.394
R326 VDDA.n275 VDDA.n273 342.3
R327 VDDA.n303 VDDA.n302 341.675
R328 VDDA.n301 VDDA.n300 341.675
R329 VDDA.n299 VDDA.n298 341.675
R330 VDDA.n297 VDDA.n296 341.675
R331 VDDA.n279 VDDA.n278 341.675
R332 VDDA.n277 VDDA.n276 341.675
R333 VDDA.n275 VDDA.n274 341.675
R334 VDDA.t416 VDDA.n442 340.635
R335 VDDA.n444 VDDA.t410 340.635
R336 VDDA.t310 VDDA.n423 340.635
R337 VDDA.n425 VDDA.t377 340.635
R338 VDDA.n407 VDDA.n406 339.272
R339 VDDA.n431 VDDA.n430 339.272
R340 VDDA.n433 VDDA.n432 339.272
R341 VDDA.n435 VDDA.n434 339.272
R342 VDDA.n437 VDDA.n436 339.272
R343 VDDA.n336 VDDA.n260 337.175
R344 VDDA.n262 VDDA.n261 337.175
R345 VDDA.n312 VDDA.n311 337.175
R346 VDDA.n315 VDDA.n309 337.175
R347 VDDA.n307 VDDA.n306 337.175
R348 VDDA.n319 VDDA.n318 337.175
R349 VDDA.n322 VDDA.n305 337.175
R350 VDDA.n325 VDDA.n324 337.175
R351 VDDA.n328 VDDA.n272 337.175
R352 VDDA.n294 VDDA.n280 337.175
R353 VDDA.n397 VDDA.n383 335.022
R354 VDDA.n173 VDDA.t397 332.75
R355 VDDA.n184 VDDA.t403 332.75
R356 VDDA.n19 VDDA.t355 332.75
R357 VDDA.n18 VDDA.t382 332.75
R358 VDDA.n14 VDDA.t421 332.75
R359 VDDA.n13 VDDA.t312 332.75
R360 VDDA.n243 VDDA.t321 314.274
R361 VDDA.n250 VDDA.t336 314.274
R362 VDDA.n21 VDDA.n16 313.601
R363 VDDA.n28 VDDA.n16 307.2
R364 VDDA.n36 VDDA.n11 307.2
R365 VDDA.n29 VDDA.n11 307.2
R366 VDDA.n445 VDDA.n409 294.401
R367 VDDA.t353 VDDA.n122 285.815
R368 VDDA.n124 VDDA.t380 285.815
R369 VDDA.t325 VDDA.n49 285.815
R370 VDDA.n51 VDDA.t359 285.815
R371 VDDA.t344 VDDA.n376 278.95
R372 VDDA.n378 VDDA.t401 278.95
R373 VDDA.n118 VDDA.t354 277.916
R374 VDDA.n116 VDDA.t381 277.916
R375 VDDA.n45 VDDA.t326 277.916
R376 VDDA.n43 VDDA.t360 277.916
R377 VDDA.n147 VDDA.n146 276.8
R378 VDDA.n142 VDDA.n141 276.8
R379 VDDA.n73 VDDA.n40 276.8
R380 VDDA.n67 VDDA.n64 276.8
R381 VDDA.n373 VDDA.t345 270.705
R382 VDDA.n381 VDDA.t402 270.705
R383 VDDA.n236 VDDA.n223 257.601
R384 VDDA.n440 VDDA.n408 246.4
R385 VDDA.t362 VDDA.n205 239.915
R386 VDDA.n207 VDDA.t389 239.915
R387 VDDA.t368 VDDA.n93 239.915
R388 VDDA.n95 VDDA.t413 239.915
R389 VDDA.n231 VDDA.n223 238.4
R390 VDDA.n203 VDDA.n202 230.4
R391 VDDA.n203 VDDA.n200 230.4
R392 VDDA.n91 VDDA.n90 230.4
R393 VDDA.n91 VDDA.n88 230.4
R394 VDDA.n459 VDDA.n403 228.8
R395 VDDA.n422 VDDA.n415 224
R396 VDDA.n426 VDDA.n415 224
R397 VDDA.n454 VDDA.n403 219.201
R398 VDDA.n120 VDDA.n119 211.201
R399 VDDA.n120 VDDA.n117 211.201
R400 VDDA.n47 VDDA.n46 211.201
R401 VDDA.n47 VDDA.n44 211.201
R402 VDDA.n26 VDDA.n20 211.201
R403 VDDA.n27 VDDA.n26 211.201
R404 VDDA.n35 VDDA.n34 211.201
R405 VDDA.n141 VDDA.n127 204.8
R406 VDDA.n147 VDDA.n127 204.8
R407 VDDA.n73 VDDA.n72 204.8
R408 VDDA.n72 VDDA.n64 204.8
R409 VDDA.n34 VDDA.n15 202.971
R410 VDDA.n208 VDDA.n200 198.4
R411 VDDA.n202 VDDA.n197 198.4
R412 VDDA.n96 VDDA.n88 198.4
R413 VDDA.n90 VDDA.n85 198.4
R414 VDDA.n231 VDDA.n230 192
R415 VDDA.t173 VDDA.t322 190
R416 VDDA.t337 VDDA.t173 190
R417 VDDA.n237 VDDA.n236 188.8
R418 VDDA.n335 VDDA.n334 188.8
R419 VDDA.n330 VDDA.n329 188.8
R420 VDDA.n394 VDDA.n388 188.8
R421 VDDA.n390 VDDA.n388 188.8
R422 VDDA.n355 VDDA.n349 188.8
R423 VDDA.n351 VDDA.n349 188.8
R424 VDDA.t62 VDDA.t404 186.607
R425 VDDA.t100 VDDA.t62 186.607
R426 VDDA.t141 VDDA.t100 186.607
R427 VDDA.t98 VDDA.t141 186.607
R428 VDDA.t22 VDDA.t98 186.607
R429 VDDA.t92 VDDA.t22 186.607
R430 VDDA.t103 VDDA.t92 186.607
R431 VDDA.t88 VDDA.t103 186.607
R432 VDDA.t159 VDDA.t88 186.607
R433 VDDA.t145 VDDA.t159 186.607
R434 VDDA.t157 VDDA.t139 186.607
R435 VDDA.t139 VDDA.t161 186.607
R436 VDDA.t161 VDDA.t64 186.607
R437 VDDA.t64 VDDA.t90 186.607
R438 VDDA.t90 VDDA.t24 186.607
R439 VDDA.t24 VDDA.t86 186.607
R440 VDDA.t86 VDDA.t165 186.607
R441 VDDA.t165 VDDA.t143 186.607
R442 VDDA.t143 VDDA.t155 186.607
R443 VDDA.t155 VDDA.t398 186.607
R444 VDDA.t129 VDDA.t422 186.607
R445 VDDA.t29 VDDA.t129 186.607
R446 VDDA.t450 VDDA.t29 186.607
R447 VDDA.t21 VDDA.t450 186.607
R448 VDDA.t97 VDDA.t21 186.607
R449 VDDA.t84 VDDA.t214 186.607
R450 VDDA.t214 VDDA.t55 186.607
R451 VDDA.t55 VDDA.t76 186.607
R452 VDDA.t76 VDDA.t57 186.607
R453 VDDA.t57 VDDA.t313 186.607
R454 VDDA.t136 VDDA.t356 183.333
R455 VDDA.t75 VDDA.t136 183.333
R456 VDDA.t15 VDDA.t75 183.333
R457 VDDA.t134 VDDA.t15 183.333
R458 VDDA.t56 VDDA.t134 183.333
R459 VDDA.t235 VDDA.t6 183.333
R460 VDDA.t6 VDDA.t135 183.333
R461 VDDA.t135 VDDA.t256 183.333
R462 VDDA.t256 VDDA.t217 183.333
R463 VDDA.t217 VDDA.t383 183.333
R464 VDDA.n375 VDDA.n374 182.4
R465 VDDA.n380 VDDA.n379 182.4
R466 VDDA.n139 VDDA.t342 178.124
R467 VDDA.n149 VDDA.t375 178.124
R468 VDDA.n62 VDDA.t348 178.124
R469 VDDA.n75 VDDA.t320 178.124
R470 VDDA.n446 VDDA.n408 176
R471 VDDA.n226 VDDA.n221 174.393
R472 VDDA.t239 VDDA.t316 172.727
R473 VDDA.t53 VDDA.t239 172.727
R474 VDDA.t210 VDDA.t53 172.727
R475 VDDA.t220 VDDA.t210 172.727
R476 VDDA.t175 VDDA.t220 172.727
R477 VDDA.t426 VDDA.t175 172.727
R478 VDDA.t438 VDDA.t426 172.727
R479 VDDA.t19 VDDA.t438 172.727
R480 VDDA.t51 VDDA.t19 172.727
R481 VDDA.t36 VDDA.t202 172.727
R482 VDDA.t71 VDDA.t36 172.727
R483 VDDA.t440 VDDA.t71 172.727
R484 VDDA.t208 VDDA.t440 172.727
R485 VDDA.t17 VDDA.t208 172.727
R486 VDDA.t114 VDDA.t17 172.727
R487 VDDA.t254 VDDA.t114 172.727
R488 VDDA.t4 VDDA.t254 172.727
R489 VDDA.t350 VDDA.t4 172.727
R490 VDDA.t77 VDDA.t419 172.727
R491 VDDA.t458 VDDA.t77 172.727
R492 VDDA.t32 VDDA.t458 172.727
R493 VDDA.t2 VDDA.t32 172.727
R494 VDDA.t149 VDDA.t2 172.727
R495 VDDA.t34 VDDA.t149 172.727
R496 VDDA.t79 VDDA.t34 172.727
R497 VDDA.t105 VDDA.t79 172.727
R498 VDDA.t60 VDDA.t105 172.727
R499 VDDA.t151 VDDA.t454 172.727
R500 VDDA.t120 VDDA.t151 172.727
R501 VDDA.t218 VDDA.t120 172.727
R502 VDDA.t122 VDDA.t218 172.727
R503 VDDA.t68 VDDA.t122 172.727
R504 VDDA.t456 VDDA.t68 172.727
R505 VDDA.t66 VDDA.t456 172.727
R506 VDDA.t212 VDDA.t66 172.727
R507 VDDA.t365 VDDA.t212 172.727
R508 VDDA.t371 VDDA.n232 172.554
R509 VDDA.n235 VDDA.t392 172.554
R510 VDDA.n340 VDDA.n339 168.435
R511 VDDA.n359 VDDA.n358 168.435
R512 VDDA.n361 VDDA.n360 168.435
R513 VDDA.n363 VDDA.n362 168.435
R514 VDDA.n365 VDDA.n364 168.435
R515 VDDA.n367 VDDA.n366 168.435
R516 VDDA.n369 VDDA.n368 168.435
R517 VDDA.n371 VDDA.n370 168.435
R518 VDDA.n245 VDDA.n218 164.8
R519 VDDA.n248 VDDA.n218 164.8
R520 VDDA.t341 VDDA.n143 161.817
R521 VDDA.n145 VDDA.t374 161.817
R522 VDDA.t319 VDDA.n65 161.817
R523 VDDA.t347 VDDA.n66 161.817
R524 VDDA.n195 VDDA.n193 160.428
R525 VDDA.n192 VDDA.n190 160.428
R526 VDDA.n83 VDDA.n81 160.428
R527 VDDA.n80 VDDA.n78 160.428
R528 VDDA.t265 VDDA.t344 159.814
R529 VDDA.t286 VDDA.t265 159.814
R530 VDDA.t297 VDDA.t286 159.814
R531 VDDA.t307 VDDA.t297 159.814
R532 VDDA.t272 VDDA.t307 159.814
R533 VDDA.t268 VDDA.t272 159.814
R534 VDDA.t291 VDDA.t268 159.814
R535 VDDA.t299 VDDA.t291 159.814
R536 VDDA.t277 VDDA.t258 159.814
R537 VDDA.t274 VDDA.t277 159.814
R538 VDDA.t293 VDDA.t274 159.814
R539 VDDA.t302 VDDA.t293 159.814
R540 VDDA.t263 VDDA.t302 159.814
R541 VDDA.t283 VDDA.t263 159.814
R542 VDDA.t281 VDDA.t283 159.814
R543 VDDA.t401 VDDA.t281 159.814
R544 VDDA.n195 VDDA.n194 159.803
R545 VDDA.n192 VDDA.n191 159.803
R546 VDDA.n83 VDDA.n82 159.803
R547 VDDA.n80 VDDA.n79 159.803
R548 VDDA.t0 VDDA.t331 158.333
R549 VDDA.t328 VDDA.t177 158.333
R550 VDDA.t207 VDDA.t386 158.333
R551 VDDA.t407 VDDA.t206 158.333
R552 VDDA.t163 VDDA.t395 158.333
R553 VDDA.t229 VDDA.t163 158.333
R554 VDDA.t442 VDDA.t227 158.333
R555 VDDA.t334 VDDA.t442 158.333
R556 VDDA.t200 VDDA.t416 155.97
R557 VDDA.t444 VDDA.t200 155.97
R558 VDDA.t452 VDDA.t444 155.97
R559 VDDA.t40 VDDA.t452 155.97
R560 VDDA.t460 VDDA.t40 155.97
R561 VDDA.t137 VDDA.t460 155.97
R562 VDDA.t196 VDDA.t198 155.97
R563 VDDA.t147 VDDA.t196 155.97
R564 VDDA.t436 VDDA.t147 155.97
R565 VDDA.t410 VDDA.t436 155.97
R566 VDDA.t94 VDDA.t310 155.97
R567 VDDA.t38 VDDA.t94 155.97
R568 VDDA.t182 VDDA.t434 155.97
R569 VDDA.t377 VDDA.t182 155.97
R570 VDDA.n201 VDDA.t363 155.125
R571 VDDA.n199 VDDA.t390 155.125
R572 VDDA.n89 VDDA.t369 155.125
R573 VDDA.n87 VDDA.t414 155.125
R574 VDDA.n139 VDDA.n138 151.882
R575 VDDA.n62 VDDA.n61 151.882
R576 VDDA.n150 VDDA.n149 151.321
R577 VDDA.n76 VDDA.n75 151.321
R578 VDDA.n125 VDDA.n117 150.4
R579 VDDA.n119 VDDA.n114 150.4
R580 VDDA.n52 VDDA.n44 150.4
R581 VDDA.n46 VDDA.n41 150.4
R582 VDDA.n211 VDDA.n210 146.002
R583 VDDA.n99 VDDA.n98 146.002
R584 VDDA.n113 VDDA.n112 145.429
R585 VDDA.n132 VDDA.n131 145.429
R586 VDDA.n134 VDDA.n133 145.429
R587 VDDA.n136 VDDA.n135 145.429
R588 VDDA.n138 VDDA.n137 145.429
R589 VDDA.n39 VDDA.n38 145.429
R590 VDDA.n55 VDDA.n54 145.429
R591 VDDA.n57 VDDA.n56 145.429
R592 VDDA.n59 VDDA.n58 145.429
R593 VDDA.n61 VDDA.n60 145.429
R594 VDDA.n149 VDDA.n148 135.387
R595 VDDA.n140 VDDA.n139 135.387
R596 VDDA.n75 VDDA.n74 135.387
R597 VDDA.n63 VDDA.n62 135.387
R598 VDDA.t172 VDDA.t353 121.513
R599 VDDA.t428 VDDA.t172 121.513
R600 VDDA.t96 VDDA.t428 121.513
R601 VDDA.t181 VDDA.t96 121.513
R602 VDDA.t451 VDDA.t181 121.513
R603 VDDA.t462 VDDA.t237 121.513
R604 VDDA.t236 VDDA.t462 121.513
R605 VDDA.t225 VDDA.t236 121.513
R606 VDDA.t127 VDDA.t225 121.513
R607 VDDA.t380 VDDA.t127 121.513
R608 VDDA.t48 VDDA.t325 121.513
R609 VDDA.t124 VDDA.t48 121.513
R610 VDDA.t187 VDDA.t124 121.513
R611 VDDA.t118 VDDA.t187 121.513
R612 VDDA.t193 VDDA.t118 121.513
R613 VDDA.t192 VDDA.t8 121.513
R614 VDDA.t28 VDDA.t192 121.513
R615 VDDA.t253 VDDA.t28 121.513
R616 VDDA.t31 VDDA.t253 121.513
R617 VDDA.t359 VDDA.t31 121.513
R618 VDDA.n334 VDDA.n265 118.4
R619 VDDA.n330 VDDA.n270 118.4
R620 VDDA.n292 VDDA.n284 118.4
R621 VDDA.n286 VDDA.n281 118.4
R622 VDDA.n395 VDDA.n394 118.4
R623 VDDA.n390 VDDA.n385 118.4
R624 VDDA.n356 VDDA.n355 118.4
R625 VDDA.n351 VDDA.n346 118.4
R626 VDDA.n454 VDDA.n453 118.4
R627 VDDA.n460 VDDA.n459 118.4
R628 VDDA.n441 VDDA.n440 118.4
R629 VDDA.n446 VDDA.n445 118.4
R630 VDDA.n422 VDDA.n421 118.4
R631 VDDA.n427 VDDA.n426 118.4
R632 VDDA.n245 VDDA.n244 110.4
R633 VDDA.n249 VDDA.n248 110.4
R634 VDDA.n453 VDDA.n402 105.6
R635 VDDA.n460 VDDA.n402 105.6
R636 VDDA.n421 VDDA.n414 105.6
R637 VDDA.n427 VDDA.n414 105.6
R638 VDDA.t392 VDDA.t231 102.704
R639 VDDA.n183 VDDA.n153 102.4
R640 VDDA.n177 VDDA.n174 102.4
R641 VDDA.n21 VDDA.n20 102.4
R642 VDDA.n240 VDDA.n239 101.267
R643 VDDA.t432 VDDA.t362 98.2764
R644 VDDA.t116 VDDA.t432 98.2764
R645 VDDA.t215 VDDA.t116 98.2764
R646 VDDA.t222 VDDA.t215 98.2764
R647 VDDA.t132 VDDA.t222 98.2764
R648 VDDA.t241 VDDA.t233 98.2764
R649 VDDA.t73 VDDA.t241 98.2764
R650 VDDA.t81 VDDA.t73 98.2764
R651 VDDA.t247 VDDA.t81 98.2764
R652 VDDA.t389 VDDA.t247 98.2764
R653 VDDA.t44 VDDA.t368 98.2764
R654 VDDA.t446 VDDA.t44 98.2764
R655 VDDA.t130 VDDA.t446 98.2764
R656 VDDA.t243 VDDA.t130 98.2764
R657 VDDA.t179 VDDA.t243 98.2764
R658 VDDA.t42 VDDA.t107 98.2764
R659 VDDA.t204 VDDA.t42 98.2764
R660 VDDA.t245 VDDA.t204 98.2764
R661 VDDA.t424 VDDA.t245 98.2764
R662 VDDA.t413 VDDA.t424 98.2764
R663 VDDA.n103 VDDA.n101 97.4034
R664 VDDA.n2 VDDA.n0 97.4034
R665 VDDA.n111 VDDA.n110 96.8409
R666 VDDA.n109 VDDA.n108 96.8409
R667 VDDA.n107 VDDA.n106 96.8409
R668 VDDA.n105 VDDA.n104 96.8409
R669 VDDA.n103 VDDA.n102 96.8409
R670 VDDA.n10 VDDA.n9 96.8409
R671 VDDA.n8 VDDA.n7 96.8409
R672 VDDA.n6 VDDA.n5 96.8409
R673 VDDA.n4 VDDA.n3 96.8409
R674 VDDA.n2 VDDA.n1 96.8409
R675 VDDA.n28 VDDA.n27 96.0005
R676 VDDA.n29 VDDA.n15 96.0005
R677 VDDA.n36 VDDA.n35 96.0005
R678 VDDA.n180 VDDA.t145 93.3041
R679 VDDA.n180 VDDA.t157 93.3041
R680 VDDA.n32 VDDA.t97 93.3041
R681 VDDA.n32 VDDA.t84 93.3041
R682 VDDA.n219 VDDA.n218 92.5005
R683 VDDA.t173 VDDA.n219 92.5005
R684 VDDA.n220 VDDA.n217 92.5005
R685 VDDA.t173 VDDA.n220 92.5005
R686 VDDA.n224 VDDA.n223 92.5005
R687 VDDA.n233 VDDA.n224 92.5005
R688 VDDA.n225 VDDA.n222 92.5005
R689 VDDA.n234 VDDA.n225 92.5005
R690 VDDA.n208 VDDA.n207 92.5005
R691 VDDA.n204 VDDA.n203 92.5005
R692 VDDA.n206 VDDA.n204 92.5005
R693 VDDA.n205 VDDA.n197 92.5005
R694 VDDA.n209 VDDA.n198 92.5005
R695 VDDA.n206 VDDA.n198 92.5005
R696 VDDA.n175 VDDA.n153 92.5005
R697 VDDA.n179 VDDA.n178 92.5005
R698 VDDA.n180 VDDA.n179 92.5005
R699 VDDA.n177 VDDA.n176 92.5005
R700 VDDA.n182 VDDA.n181 92.5005
R701 VDDA.n181 VDDA.n180 92.5005
R702 VDDA.n125 VDDA.n124 92.5005
R703 VDDA.n121 VDDA.n120 92.5005
R704 VDDA.n123 VDDA.n121 92.5005
R705 VDDA.n122 VDDA.n114 92.5005
R706 VDDA.n126 VDDA.n115 92.5005
R707 VDDA.n123 VDDA.n115 92.5005
R708 VDDA.n130 VDDA.n127 92.5005
R709 VDDA.n144 VDDA.n130 92.5005
R710 VDDA.n129 VDDA.n128 92.5005
R711 VDDA.n144 VDDA.n129 92.5005
R712 VDDA.n96 VDDA.n95 92.5005
R713 VDDA.n92 VDDA.n91 92.5005
R714 VDDA.n94 VDDA.n92 92.5005
R715 VDDA.n93 VDDA.n85 92.5005
R716 VDDA.n97 VDDA.n86 92.5005
R717 VDDA.n94 VDDA.n86 92.5005
R718 VDDA.n52 VDDA.n51 92.5005
R719 VDDA.n48 VDDA.n47 92.5005
R720 VDDA.n50 VDDA.n48 92.5005
R721 VDDA.n49 VDDA.n41 92.5005
R722 VDDA.n53 VDDA.n42 92.5005
R723 VDDA.n50 VDDA.n42 92.5005
R724 VDDA.n72 VDDA.n71 92.5005
R725 VDDA.n71 VDDA.n70 92.5005
R726 VDDA.n69 VDDA.n68 92.5005
R727 VDDA.n70 VDDA.n69 92.5005
R728 VDDA.n23 VDDA.n16 92.5005
R729 VDDA.n24 VDDA.n23 92.5005
R730 VDDA.n22 VDDA.n21 92.5005
R731 VDDA.n26 VDDA.n25 92.5005
R732 VDDA.n25 VDDA.n24 92.5005
R733 VDDA.n28 VDDA.n17 92.5005
R734 VDDA.n31 VDDA.n11 92.5005
R735 VDDA.n32 VDDA.n31 92.5005
R736 VDDA.n30 VDDA.n29 92.5005
R737 VDDA.n34 VDDA.n33 92.5005
R738 VDDA.n33 VDDA.n32 92.5005
R739 VDDA.n36 VDDA.n12 92.5005
R740 VDDA.n317 VDDA.n267 92.5005
R741 VDDA.n332 VDDA.n267 92.5005
R742 VDDA.n334 VDDA.n333 92.5005
R743 VDDA.n269 VDDA.n266 92.5005
R744 VDDA.n332 VDDA.n266 92.5005
R745 VDDA.n331 VDDA.n330 92.5005
R746 VDDA.n292 VDDA.n291 92.5005
R747 VDDA.n288 VDDA.n287 92.5005
R748 VDDA.n290 VDDA.n288 92.5005
R749 VDDA.n289 VDDA.n281 92.5005
R750 VDDA.n293 VDDA.n282 92.5005
R751 VDDA.n290 VDDA.n282 92.5005
R752 VDDA.n394 VDDA.n393 92.5005
R753 VDDA.n389 VDDA.n388 92.5005
R754 VDDA.n392 VDDA.n389 92.5005
R755 VDDA.n391 VDDA.n390 92.5005
R756 VDDA.n396 VDDA.n386 92.5005
R757 VDDA.n392 VDDA.n386 92.5005
R758 VDDA.n376 VDDA.n375 92.5005
R759 VDDA.n343 VDDA.n342 92.5005
R760 VDDA.n377 VDDA.n343 92.5005
R761 VDDA.n379 VDDA.n378 92.5005
R762 VDDA.n344 VDDA.n341 92.5005
R763 VDDA.n377 VDDA.n344 92.5005
R764 VDDA.n355 VDDA.n354 92.5005
R765 VDDA.n350 VDDA.n349 92.5005
R766 VDDA.n353 VDDA.n350 92.5005
R767 VDDA.n352 VDDA.n351 92.5005
R768 VDDA.n357 VDDA.n347 92.5005
R769 VDDA.n353 VDDA.n347 92.5005
R770 VDDA.n455 VDDA.n454 92.5005
R771 VDDA.n404 VDDA.n403 92.5005
R772 VDDA.n456 VDDA.n404 92.5005
R773 VDDA.n459 VDDA.n458 92.5005
R774 VDDA.n405 VDDA.n402 92.5005
R775 VDDA.n457 VDDA.n405 92.5005
R776 VDDA.n442 VDDA.n441 92.5005
R777 VDDA.n410 VDDA.n409 92.5005
R778 VDDA.n443 VDDA.n410 92.5005
R779 VDDA.n445 VDDA.n444 92.5005
R780 VDDA.n411 VDDA.n408 92.5005
R781 VDDA.n443 VDDA.n411 92.5005
R782 VDDA.n423 VDDA.n422 92.5005
R783 VDDA.n416 VDDA.n415 92.5005
R784 VDDA.n424 VDDA.n416 92.5005
R785 VDDA.n426 VDDA.n425 92.5005
R786 VDDA.n417 VDDA.n414 92.5005
R787 VDDA.n424 VDDA.n417 92.5005
R788 VDDA.n24 VDDA.t56 91.6672
R789 VDDA.n24 VDDA.t235 91.6672
R790 VDDA.n228 VDDA.n227 87.4672
R791 VDDA.n332 VDDA.t51 86.3641
R792 VDDA.t202 VDDA.n332 86.3641
R793 VDDA.n290 VDDA.t60 86.3641
R794 VDDA.t454 VDDA.n290 86.3641
R795 VDDA.n227 VDDA.t372 85.438
R796 VDDA.n239 VDDA.t393 85.438
R797 VDDA.n233 VDDA.t371 81.3068
R798 VDDA.n239 VDDA.n238 81.0672
R799 VDDA.n229 VDDA.n227 81.0672
R800 VDDA.n377 VDDA.t299 79.907
R801 VDDA.t258 VDDA.n377 79.907
R802 VDDA.n392 VDDA.t0 79.1672
R803 VDDA.t177 VDDA.n392 79.1672
R804 VDDA.n353 VDDA.t207 79.1672
R805 VDDA.t206 VDDA.n353 79.1672
R806 VDDA.t227 VDDA.n457 79.1672
R807 VDDA.n151 VDDA.t63 78.8005
R808 VDDA.n151 VDDA.t101 78.8005
R809 VDDA.n154 VDDA.t142 78.8005
R810 VDDA.n154 VDDA.t99 78.8005
R811 VDDA.n156 VDDA.t23 78.8005
R812 VDDA.n156 VDDA.t93 78.8005
R813 VDDA.n158 VDDA.t104 78.8005
R814 VDDA.n158 VDDA.t89 78.8005
R815 VDDA.n160 VDDA.t160 78.8005
R816 VDDA.n160 VDDA.t146 78.8005
R817 VDDA.n162 VDDA.t158 78.8005
R818 VDDA.n162 VDDA.t140 78.8005
R819 VDDA.n164 VDDA.t162 78.8005
R820 VDDA.n164 VDDA.t65 78.8005
R821 VDDA.n166 VDDA.t91 78.8005
R822 VDDA.n166 VDDA.t25 78.8005
R823 VDDA.n168 VDDA.t87 78.8005
R824 VDDA.n168 VDDA.t166 78.8005
R825 VDDA.n170 VDDA.t144 78.8005
R826 VDDA.n170 VDDA.t156 78.8005
R827 VDDA.n443 VDDA.t137 77.9856
R828 VDDA.t198 VDDA.n443 77.9856
R829 VDDA.n424 VDDA.t38 77.9856
R830 VDDA.t434 VDDA.n424 77.9856
R831 VDDA.n237 VDDA.n222 64.0005
R832 VDDA.n329 VDDA.n271 64.0005
R833 VDDA.n321 VDDA.n271 64.0005
R834 VDDA.n321 VDDA.n320 64.0005
R835 VDDA.n320 VDDA.n317 64.0005
R836 VDDA.n317 VDDA.n316 64.0005
R837 VDDA.n316 VDDA.n308 64.0005
R838 VDDA.n308 VDDA.n263 64.0005
R839 VDDA.n335 VDDA.n263 64.0005
R840 VDDA.n357 VDDA.n356 64.0005
R841 VDDA.n357 VDDA.n346 64.0005
R842 VDDA.t170 VDDA.t341 62.9523
R843 VDDA.t430 VDDA.t170 62.9523
R844 VDDA.t109 VDDA.t430 62.9523
R845 VDDA.t112 VDDA.t109 62.9523
R846 VDDA.t466 VDDA.t112 62.9523
R847 VDDA.t464 VDDA.t167 62.9523
R848 VDDA.t153 VDDA.t464 62.9523
R849 VDDA.t58 VDDA.t153 62.9523
R850 VDDA.t448 VDDA.t58 62.9523
R851 VDDA.t374 VDDA.t448 62.9523
R852 VDDA.t9 VDDA.t319 62.9523
R853 VDDA.t125 VDDA.t9 62.9523
R854 VDDA.t188 VDDA.t125 62.9523
R855 VDDA.t12 VDDA.t188 62.9523
R856 VDDA.t190 VDDA.t12 62.9523
R857 VDDA.t26 VDDA.t250 62.9523
R858 VDDA.t250 VDDA.t184 62.9523
R859 VDDA.t184 VDDA.t49 62.9523
R860 VDDA.t49 VDDA.t194 62.9523
R861 VDDA.t194 VDDA.t347 62.9523
R862 VDDA.n396 VDDA.n395 62.7205
R863 VDDA.n396 VDDA.n385 62.7205
R864 VDDA.n215 VDDA.t174 62.5402
R865 VDDA.n215 VDDA.t338 62.5402
R866 VDDA.n246 VDDA.n245 61.6672
R867 VDDA.n248 VDDA.n247 61.6672
R868 VDDA.n146 VDDA.n145 61.6672
R869 VDDA.n143 VDDA.n142 61.6672
R870 VDDA.n65 VDDA.n40 61.6672
R871 VDDA.n67 VDDA.n66 61.6672
R872 VDDA.n123 VDDA.t451 60.7563
R873 VDDA.t237 VDDA.n123 60.7563
R874 VDDA.n50 VDDA.t193 60.7563
R875 VDDA.t8 VDDA.n50 60.7563
R876 VDDA.n256 VDDA.t471 59.5681
R877 VDDA.n255 VDDA.t469 59.5681
R878 VDDA.n244 VDDA.n217 57.6005
R879 VDDA.n249 VDDA.n217 57.6005
R880 VDDA.n456 VDDA.t229 57.5763
R881 VDDA.n255 VDDA.t472 51.8888
R882 VDDA.n230 VDDA.n222 51.2005
R883 VDDA.n206 VDDA.t132 49.1384
R884 VDDA.t233 VDDA.n206 49.1384
R885 VDDA.n94 VDDA.t179 49.1384
R886 VDDA.t107 VDDA.n94 49.1384
R887 VDDA.n257 VDDA.t470 48.9557
R888 VDDA.n252 VDDA.n251 48.3605
R889 VDDA.n242 VDDA.n241 43.8605
R890 VDDA.n172 VDDA.n171 42.0963
R891 VDDA.n186 VDDA.n185 41.5338
R892 VDDA.n260 VDDA.t255 39.4005
R893 VDDA.n260 VDDA.t5 39.4005
R894 VDDA.n261 VDDA.t18 39.4005
R895 VDDA.n261 VDDA.t115 39.4005
R896 VDDA.n311 VDDA.t441 39.4005
R897 VDDA.n311 VDDA.t209 39.4005
R898 VDDA.n309 VDDA.t37 39.4005
R899 VDDA.n309 VDDA.t72 39.4005
R900 VDDA.n306 VDDA.t52 39.4005
R901 VDDA.n306 VDDA.t203 39.4005
R902 VDDA.n318 VDDA.t439 39.4005
R903 VDDA.n318 VDDA.t20 39.4005
R904 VDDA.n305 VDDA.t176 39.4005
R905 VDDA.n305 VDDA.t427 39.4005
R906 VDDA.n324 VDDA.t211 39.4005
R907 VDDA.n324 VDDA.t221 39.4005
R908 VDDA.n272 VDDA.t240 39.4005
R909 VDDA.n272 VDDA.t54 39.4005
R910 VDDA.n302 VDDA.t67 39.4005
R911 VDDA.n302 VDDA.t213 39.4005
R912 VDDA.n300 VDDA.t69 39.4005
R913 VDDA.n300 VDDA.t457 39.4005
R914 VDDA.n298 VDDA.t219 39.4005
R915 VDDA.n298 VDDA.t123 39.4005
R916 VDDA.n296 VDDA.t152 39.4005
R917 VDDA.n296 VDDA.t121 39.4005
R918 VDDA.n280 VDDA.t61 39.4005
R919 VDDA.n280 VDDA.t455 39.4005
R920 VDDA.n278 VDDA.t80 39.4005
R921 VDDA.n278 VDDA.t106 39.4005
R922 VDDA.n276 VDDA.t150 39.4005
R923 VDDA.n276 VDDA.t35 39.4005
R924 VDDA.n274 VDDA.t33 39.4005
R925 VDDA.n274 VDDA.t3 39.4005
R926 VDDA.n273 VDDA.t78 39.4005
R927 VDDA.n273 VDDA.t459 39.4005
R928 VDDA.n383 VDDA.t1 39.4005
R929 VDDA.n383 VDDA.t178 39.4005
R930 VDDA.n400 VDDA.t228 39.4005
R931 VDDA.n400 VDDA.t443 39.4005
R932 VDDA.n449 VDDA.t164 39.4005
R933 VDDA.n449 VDDA.t230 39.4005
R934 VDDA.n406 VDDA.t148 39.4005
R935 VDDA.n406 VDDA.t437 39.4005
R936 VDDA.n430 VDDA.t199 39.4005
R937 VDDA.n430 VDDA.t197 39.4005
R938 VDDA.n432 VDDA.t461 39.4005
R939 VDDA.n432 VDDA.t138 39.4005
R940 VDDA.n434 VDDA.t453 39.4005
R941 VDDA.n434 VDDA.t41 39.4005
R942 VDDA.n436 VDDA.t201 39.4005
R943 VDDA.n436 VDDA.t445 39.4005
R944 VDDA.n412 VDDA.t435 39.4005
R945 VDDA.n412 VDDA.t183 39.4005
R946 VDDA.n418 VDDA.t95 39.4005
R947 VDDA.n418 VDDA.t39 39.4005
R948 VDDA.n144 VDDA.t466 31.4764
R949 VDDA.t167 VDDA.n144 31.4764
R950 VDDA.n70 VDDA.t190 31.4764
R951 VDDA.n70 VDDA.t26 31.4764
R952 VDDA.n29 VDDA.n28 28.663
R953 VDDA.n251 VDDA.n250 25.6005
R954 VDDA.n243 VDDA.n242 25.6005
R955 VDDA.n185 VDDA.n184 25.6005
R956 VDDA.n173 VDDA.n172 25.6005
R957 VDDA.n258 VDDA.n254 24.7453
R958 VDDA.n250 VDDA.n249 24.5338
R959 VDDA.n244 VDDA.n243 24.5338
R960 VDDA.n238 VDDA.n237 24.5338
R961 VDDA.n230 VDDA.n229 24.5338
R962 VDDA.n457 VDDA.n456 21.5914
R963 VDDA.n254 VDDA.n253 21.5392
R964 VDDA.n202 VDDA.n201 21.3338
R965 VDDA.n200 VDDA.n199 21.3338
R966 VDDA.n184 VDDA.n183 21.3338
R967 VDDA.n174 VDDA.n173 21.3338
R968 VDDA.n119 VDDA.n118 21.3338
R969 VDDA.n117 VDDA.n116 21.3338
R970 VDDA.n148 VDDA.n147 21.3338
R971 VDDA.n141 VDDA.n140 21.3338
R972 VDDA.n90 VDDA.n89 21.3338
R973 VDDA.n88 VDDA.n87 21.3338
R974 VDDA.n46 VDDA.n45 21.3338
R975 VDDA.n44 VDDA.n43 21.3338
R976 VDDA.n74 VDDA.n73 21.3338
R977 VDDA.n64 VDDA.n63 21.3338
R978 VDDA.n20 VDDA.n19 21.3338
R979 VDDA.n27 VDDA.n18 21.3338
R980 VDDA.n15 VDDA.n14 21.3338
R981 VDDA.n35 VDDA.n13 21.3338
R982 VDDA.n265 VDDA.n264 21.3338
R983 VDDA.n270 VDDA.n268 21.3338
R984 VDDA.n284 VDDA.n283 21.3338
R985 VDDA.n286 VDDA.n285 21.3338
R986 VDDA.n395 VDDA.n387 21.3338
R987 VDDA.n385 VDDA.n384 21.3338
R988 VDDA.n356 VDDA.n348 21.3338
R989 VDDA.n346 VDDA.n345 21.3338
R990 VDDA.n37 VDDA.n36 19.5505
R991 VDDA.n127 VDDA.n126 19.538
R992 VDDA.n72 VDDA.n53 19.538
R993 VDDA.n211 VDDA.n209 19.2005
R994 VDDA.n99 VDDA.n97 19.2005
R995 VDDA.n381 VDDA.n380 19.2005
R996 VDDA.n374 VDDA.n373 19.2005
R997 VDDA.n461 VDDA.n460 19.2005
R998 VDDA.n453 VDDA.n452 19.2005
R999 VDDA.n447 VDDA.n446 19.2005
R1000 VDDA.n440 VDDA.n439 19.2005
R1001 VDDA.n428 VDDA.n427 19.2005
R1002 VDDA.n421 VDDA.n420 19.2005
R1003 VDDA.n232 VDDA.n231 18.5005
R1004 VDDA.n236 VDDA.n235 18.5005
R1005 VDDA.t231 VDDA.n234 17.1176
R1006 VDDA.n188 VDDA.n111 16.8443
R1007 VDDA.n372 VDDA.n357 16.363
R1008 VDDA.n468 VDDA.t267 15.0181
R1009 VDDA.n420 VDDA.n419 14.363
R1010 VDDA.n228 VDDA.n221 14.0505
R1011 VDDA.n373 VDDA.n372 13.8005
R1012 VDDA.n382 VDDA.n381 13.8005
R1013 VDDA.n452 VDDA.n451 13.8005
R1014 VDDA.n439 VDDA.n438 13.8005
R1015 VDDA.n429 VDDA.n428 13.8005
R1016 VDDA.n448 VDDA.n447 13.8005
R1017 VDDA.n462 VDDA.n461 13.8005
R1018 VDDA.n37 VDDA.n10 13.6255
R1019 VDDA.n213 VDDA.n189 13.563
R1020 VDDA.n339 VDDA.t284 13.1338
R1021 VDDA.n339 VDDA.t282 13.1338
R1022 VDDA.n358 VDDA.t303 13.1338
R1023 VDDA.n358 VDDA.t264 13.1338
R1024 VDDA.n360 VDDA.t275 13.1338
R1025 VDDA.n360 VDDA.t294 13.1338
R1026 VDDA.n362 VDDA.t259 13.1338
R1027 VDDA.n362 VDDA.t278 13.1338
R1028 VDDA.n364 VDDA.t292 13.1338
R1029 VDDA.n364 VDDA.t300 13.1338
R1030 VDDA.n366 VDDA.t273 13.1338
R1031 VDDA.n366 VDDA.t269 13.1338
R1032 VDDA.n368 VDDA.t298 13.1338
R1033 VDDA.n368 VDDA.t308 13.1338
R1034 VDDA.n370 VDDA.t266 13.1338
R1035 VDDA.n370 VDDA.t287 13.1338
R1036 VDDA.t372 VDDA.n226 12.313
R1037 VDDA.n226 VDDA.t232 12.313
R1038 VDDA.n210 VDDA.t133 11.2576
R1039 VDDA.n210 VDDA.t234 11.2576
R1040 VDDA.n194 VDDA.t242 11.2576
R1041 VDDA.n194 VDDA.t74 11.2576
R1042 VDDA.n193 VDDA.t82 11.2576
R1043 VDDA.n193 VDDA.t248 11.2576
R1044 VDDA.n191 VDDA.t216 11.2576
R1045 VDDA.n191 VDDA.t223 11.2576
R1046 VDDA.n190 VDDA.t433 11.2576
R1047 VDDA.n190 VDDA.t117 11.2576
R1048 VDDA.n98 VDDA.t180 11.2576
R1049 VDDA.n98 VDDA.t108 11.2576
R1050 VDDA.n82 VDDA.t43 11.2576
R1051 VDDA.n82 VDDA.t205 11.2576
R1052 VDDA.n81 VDDA.t246 11.2576
R1053 VDDA.n81 VDDA.t425 11.2576
R1054 VDDA.n79 VDDA.t131 11.2576
R1055 VDDA.n79 VDDA.t244 11.2576
R1056 VDDA.n78 VDDA.t45 11.2576
R1057 VDDA.n78 VDDA.t447 11.2576
R1058 VDDA.n189 VDDA.n188 9.5005
R1059 VDDA.n212 VDDA.n211 9.3005
R1060 VDDA.n100 VDDA.n99 9.3005
R1061 VDDA.n325 VDDA.n271 9.3005
R1062 VDDA.n322 VDDA.n321 9.3005
R1063 VDDA.n320 VDDA.n319 9.3005
R1064 VDDA.n317 VDDA.n307 9.3005
R1065 VDDA.n316 VDDA.n315 9.3005
R1066 VDDA.n312 VDDA.n308 9.3005
R1067 VDDA.n263 VDDA.n262 9.3005
R1068 VDDA.n336 VDDA.n335 9.3005
R1069 VDDA.n329 VDDA.n328 9.3005
R1070 VDDA.n294 VDDA.n293 9.3005
R1071 VDDA.n397 VDDA.n396 9.3005
R1072 VDDA.n241 VDDA.n240 8.938
R1073 VDDA.n258 VDDA.n257 8.03219
R1074 VDDA.n110 VDDA.t70 8.0005
R1075 VDDA.n110 VDDA.t16 8.0005
R1076 VDDA.n108 VDDA.t111 8.0005
R1077 VDDA.n108 VDDA.t429 8.0005
R1078 VDDA.n106 VDDA.t468 8.0005
R1079 VDDA.n106 VDDA.t83 8.0005
R1080 VDDA.n104 VDDA.t226 8.0005
R1081 VDDA.n104 VDDA.t102 8.0005
R1082 VDDA.n102 VDDA.t463 8.0005
R1083 VDDA.n102 VDDA.t169 8.0005
R1084 VDDA.n101 VDDA.t128 8.0005
R1085 VDDA.n101 VDDA.t238 8.0005
R1086 VDDA.n9 VDDA.t85 8.0005
R1087 VDDA.n9 VDDA.t47 8.0005
R1088 VDDA.n7 VDDA.t14 8.0005
R1089 VDDA.n7 VDDA.t7 8.0005
R1090 VDDA.n5 VDDA.t30 8.0005
R1091 VDDA.n5 VDDA.t252 8.0005
R1092 VDDA.n3 VDDA.t186 8.0005
R1093 VDDA.n3 VDDA.t11 8.0005
R1094 VDDA.n1 VDDA.t119 8.0005
R1095 VDDA.n1 VDDA.t46 8.0005
R1096 VDDA.n0 VDDA.t249 8.0005
R1097 VDDA.n0 VDDA.t224 8.0005
R1098 VDDA.n213 VDDA.n212 7.8755
R1099 VDDA.n189 VDDA.n100 7.8755
R1100 VDDA.n463 VDDA.n462 7.44175
R1101 VDDA.n253 VDDA.n252 6.6255
R1102 VDDA.n112 VDDA.t59 6.56717
R1103 VDDA.n112 VDDA.t449 6.56717
R1104 VDDA.n131 VDDA.t465 6.56717
R1105 VDDA.n131 VDDA.t154 6.56717
R1106 VDDA.n133 VDDA.t467 6.56717
R1107 VDDA.n133 VDDA.t168 6.56717
R1108 VDDA.n135 VDDA.t110 6.56717
R1109 VDDA.n135 VDDA.t113 6.56717
R1110 VDDA.n137 VDDA.t171 6.56717
R1111 VDDA.n137 VDDA.t431 6.56717
R1112 VDDA.n38 VDDA.t10 6.56717
R1113 VDDA.n38 VDDA.t126 6.56717
R1114 VDDA.n54 VDDA.t189 6.56717
R1115 VDDA.n54 VDDA.t13 6.56717
R1116 VDDA.n56 VDDA.t191 6.56717
R1117 VDDA.n56 VDDA.t27 6.56717
R1118 VDDA.n58 VDDA.t251 6.56717
R1119 VDDA.n58 VDDA.t185 6.56717
R1120 VDDA.n60 VDDA.t50 6.56717
R1121 VDDA.n60 VDDA.t195 6.56717
R1122 VDDA.n399 VDDA.n398 6.13371
R1123 VDDA.n338 VDDA.n337 6.098
R1124 VDDA.n77 VDDA.n76 5.438
R1125 VDDA.n241 VDDA.n216 5.1255
R1126 VDDA.n214 VDDA.n77 5.0005
R1127 VDDA.n212 VDDA.n196 4.5005
R1128 VDDA.n188 VDDA.n187 4.5005
R1129 VDDA.n100 VDDA.n84 4.5005
R1130 VDDA.n214 VDDA.n213 4.5005
R1131 VDDA.n295 VDDA.n294 4.5005
R1132 VDDA.n328 VDDA.n327 4.5005
R1133 VDDA.n326 VDDA.n325 4.5005
R1134 VDDA.n323 VDDA.n322 4.5005
R1135 VDDA.n319 VDDA.n304 4.5005
R1136 VDDA.n310 VDDA.n307 4.5005
R1137 VDDA.n315 VDDA.n314 4.5005
R1138 VDDA.n313 VDDA.n312 4.5005
R1139 VDDA.n262 VDDA.n259 4.5005
R1140 VDDA.n337 VDDA.n336 4.5005
R1141 VDDA.n398 VDDA.n397 4.5005
R1142 VDDA.n234 VDDA.n233 4.27978
R1143 VDDA.n256 VDDA.n255 4.12334
R1144 VDDA.n469 VDDA 4.08025
R1145 VDDA.n327 VDDA.n303 3.3755
R1146 VDDA.n77 VDDA.n37 3.09425
R1147 VDDA.n187 VDDA.n186 2.938
R1148 VDDA.n257 VDDA.n256 2.93377
R1149 VDDA.n451 VDDA.n448 2.5005
R1150 VDDA.n398 VDDA.n382 2.47371
R1151 VDDA.n253 VDDA.n214 1.938
R1152 VDDA.n438 VDDA.n429 1.813
R1153 VDDA VDDA.n469 1.20605
R1154 VDDA VDDA.n468 1.0815
R1155 VDDA.n372 VDDA.n371 1.0005
R1156 VDDA.n371 VDDA.n369 1.0005
R1157 VDDA.n369 VDDA.n367 1.0005
R1158 VDDA.n367 VDDA.n365 1.0005
R1159 VDDA.n365 VDDA.n363 1.0005
R1160 VDDA.n363 VDDA.n361 1.0005
R1161 VDDA.n361 VDDA.n359 1.0005
R1162 VDDA.n359 VDDA.n340 1.0005
R1163 VDDA.n382 VDDA.n340 1.0005
R1164 VDDA.n187 VDDA.n150 0.938
R1165 VDDA.n338 VDDA.n258 0.840625
R1166 VDDA.n469 VDDA.n254 0.7948
R1167 VDDA.n399 VDDA.n338 0.74075
R1168 VDDA.n240 VDDA.n221 0.6255
R1169 VDDA.n196 VDDA.n195 0.6255
R1170 VDDA.n196 VDDA.n192 0.6255
R1171 VDDA.n84 VDDA.n83 0.6255
R1172 VDDA.n84 VDDA.n80 0.6255
R1173 VDDA.n277 VDDA.n275 0.6255
R1174 VDDA.n279 VDDA.n277 0.6255
R1175 VDDA.n295 VDDA.n279 0.6255
R1176 VDDA.n297 VDDA.n295 0.6255
R1177 VDDA.n299 VDDA.n297 0.6255
R1178 VDDA.n301 VDDA.n299 0.6255
R1179 VDDA.n303 VDDA.n301 0.6255
R1180 VDDA.n327 VDDA.n326 0.6255
R1181 VDDA.n326 VDDA.n323 0.6255
R1182 VDDA.n323 VDDA.n304 0.6255
R1183 VDDA.n310 VDDA.n304 0.6255
R1184 VDDA.n314 VDDA.n310 0.6255
R1185 VDDA.n314 VDDA.n313 0.6255
R1186 VDDA.n313 VDDA.n259 0.6255
R1187 VDDA.n337 VDDA.n259 0.6255
R1188 VDDA.n171 VDDA.n169 0.563
R1189 VDDA.n169 VDDA.n167 0.563
R1190 VDDA.n167 VDDA.n165 0.563
R1191 VDDA.n165 VDDA.n163 0.563
R1192 VDDA.n163 VDDA.n161 0.563
R1193 VDDA.n161 VDDA.n159 0.563
R1194 VDDA.n159 VDDA.n157 0.563
R1195 VDDA.n157 VDDA.n155 0.563
R1196 VDDA.n155 VDDA.n152 0.563
R1197 VDDA.n186 VDDA.n152 0.563
R1198 VDDA.n138 VDDA.n136 0.563
R1199 VDDA.n136 VDDA.n134 0.563
R1200 VDDA.n134 VDDA.n132 0.563
R1201 VDDA.n132 VDDA.n113 0.563
R1202 VDDA.n150 VDDA.n113 0.563
R1203 VDDA.n105 VDDA.n103 0.563
R1204 VDDA.n107 VDDA.n105 0.563
R1205 VDDA.n109 VDDA.n107 0.563
R1206 VDDA.n111 VDDA.n109 0.563
R1207 VDDA.n61 VDDA.n59 0.563
R1208 VDDA.n59 VDDA.n57 0.563
R1209 VDDA.n57 VDDA.n55 0.563
R1210 VDDA.n55 VDDA.n39 0.563
R1211 VDDA.n76 VDDA.n39 0.563
R1212 VDDA.n4 VDDA.n2 0.563
R1213 VDDA.n6 VDDA.n4 0.563
R1214 VDDA.n8 VDDA.n6 0.563
R1215 VDDA.n10 VDDA.n8 0.563
R1216 VDDA.n419 VDDA.n413 0.563
R1217 VDDA.n429 VDDA.n413 0.563
R1218 VDDA.n438 VDDA.n437 0.563
R1219 VDDA.n437 VDDA.n435 0.563
R1220 VDDA.n435 VDDA.n433 0.563
R1221 VDDA.n433 VDDA.n431 0.563
R1222 VDDA.n431 VDDA.n407 0.563
R1223 VDDA.n448 VDDA.n407 0.563
R1224 VDDA.n451 VDDA.n450 0.563
R1225 VDDA.n450 VDDA.n401 0.563
R1226 VDDA.n462 VDDA.n401 0.563
R1227 VDDA.n463 VDDA.n399 0.546875
R1228 VDDA.n468 VDDA.n463 0.370625
R1229 VDDA.n252 VDDA.n216 0.2505
R1230 VDDA.t260 VDDA.t276 0.1603
R1231 VDDA.t304 VDDA.t296 0.1603
R1232 VDDA.t301 VDDA.t261 0.1603
R1233 VDDA.t289 VDDA.t285 0.1603
R1234 VDDA.t262 VDDA.t279 0.1603
R1235 VDDA.t306 VDDA.t290 0.1603
R1236 VDDA.t280 VDDA.t295 0.1603
R1237 VDDA.t271 VDDA.t257 0.1603
R1238 VDDA.n465 VDDA.t288 0.159278
R1239 VDDA.n466 VDDA.t270 0.159278
R1240 VDDA.n467 VDDA.t305 0.159278
R1241 VDDA.n467 VDDA.t260 0.1368
R1242 VDDA.n467 VDDA.t304 0.1368
R1243 VDDA.n466 VDDA.t301 0.1368
R1244 VDDA.n466 VDDA.t289 0.1368
R1245 VDDA.n465 VDDA.t262 0.1368
R1246 VDDA.n465 VDDA.t306 0.1368
R1247 VDDA.n464 VDDA.t280 0.1368
R1248 VDDA.n464 VDDA.t271 0.1368
R1249 VDDA.t288 VDDA.n464 0.00152174
R1250 VDDA.t270 VDDA.n465 0.00152174
R1251 VDDA.t305 VDDA.n466 0.00152174
R1252 VDDA.t267 VDDA.n467 0.00152174
R1253 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 628.034
R1254 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 626.784
R1255 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 622.284
R1256 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 289.2
R1257 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 289.2
R1258 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 227.252
R1259 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 212.733
R1260 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 212.733
R1261 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 176.733
R1262 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 176.733
R1263 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R1264 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 176.733
R1265 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 176.733
R1266 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 152
R1267 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 152
R1268 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 112.468
R1269 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 112.468
R1270 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R1271 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R1272 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 112.468
R1273 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R1274 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R1275 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 112.468
R1276 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 78.8005
R1277 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 78.8005
R1278 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R1279 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R1280 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R1281 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 78.8005
R1282 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 48.0005
R1283 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 48.0005
R1284 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R1285 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R1286 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 48.0005
R1287 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 48.0005
R1288 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R1289 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 45.5227
R1290 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 45.5227
R1291 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 45.5227
R1292 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 15.488
R1293 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 14.238
R1294 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 6.1255
R1295 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 5.7505
R1296 a_9610_5930.n2 a_9610_5930.n0 227.096
R1297 a_9610_5930.n7 a_9610_5930.n6 227.096
R1298 a_9610_5930.n6 a_9610_5930.n5 226.534
R1299 a_9610_5930.n4 a_9610_5930.n3 226.534
R1300 a_9610_5930.n2 a_9610_5930.n1 226.534
R1301 a_9610_5930.n5 a_9610_5930.t0 48.0005
R1302 a_9610_5930.n5 a_9610_5930.t5 48.0005
R1303 a_9610_5930.n3 a_9610_5930.t7 48.0005
R1304 a_9610_5930.n3 a_9610_5930.t9 48.0005
R1305 a_9610_5930.n1 a_9610_5930.t1 48.0005
R1306 a_9610_5930.n1 a_9610_5930.t4 48.0005
R1307 a_9610_5930.n0 a_9610_5930.t6 48.0005
R1308 a_9610_5930.n0 a_9610_5930.t2 48.0005
R1309 a_9610_5930.t8 a_9610_5930.n7 48.0005
R1310 a_9610_5930.n7 a_9610_5930.t3 48.0005
R1311 a_9610_5930.n4 a_9610_5930.n2 0.563
R1312 a_9610_5930.n6 a_9610_5930.n4 0.563
R1313 GNDA.n384 GNDA.n30 227083
R1314 GNDA.n1682 GNDA.n1681 33145.9
R1315 GNDA.n2465 GNDA.n57 30529.2
R1316 GNDA.n387 GNDA.n327 29344.6
R1317 GNDA.n1613 GNDA.n83 28608.1
R1318 GNDA.n2465 GNDA.n56 28430.8
R1319 GNDA.n385 GNDA.n327 28430.8
R1320 GNDA.n386 GNDA.n384 26656.2
R1321 GNDA.n1680 GNDA.n1613 26648.4
R1322 GNDA.n385 GNDA.n79 23523.1
R1323 GNDA.n79 GNDA.n56 23523.1
R1324 GNDA.n1681 GNDA.n82 21442.2
R1325 GNDA.n2446 GNDA.n2445 21037.5
R1326 GNDA.n1681 GNDA.n83 19885.8
R1327 GNDA.n2448 GNDA.n79 19630.8
R1328 GNDA.n2447 GNDA.n80 19055.4
R1329 GNDA.n385 GNDA.n80 17609.2
R1330 GNDA.n2450 GNDA.n56 17609.2
R1331 GNDA.n1684 GNDA.n1680 17265.8
R1332 GNDA.n2448 GNDA.n2447 15992.3
R1333 GNDA.n1682 GNDA.n1680 15861.4
R1334 GNDA.n1686 GNDA.n1615 12361.8
R1335 GNDA.n1690 GNDA.n1615 12312.5
R1336 GNDA.n384 GNDA.n56 11934.7
R1337 GNDA.n1686 GNDA.n1616 11918.5
R1338 GNDA.n1690 GNDA.n1616 11869.2
R1339 GNDA.n490 GNDA.n80 10910.2
R1340 GNDA.n2449 GNDA.n2448 10879.5
R1341 GNDA.n469 GNDA.n363 10441
R1342 GNDA.n459 GNDA.n363 10441
R1343 GNDA.n469 GNDA.n364 10441
R1344 GNDA.n459 GNDA.n364 10441
R1345 GNDA.n1730 GNDA.n1613 10371.4
R1346 GNDA.n2484 GNDA.n31 9259
R1347 GNDA.n1693 GNDA.n1642 9062
R1348 GNDA.n2484 GNDA.n32 8914.25
R1349 GNDA.n106 GNDA.n102 8175.5
R1350 GNDA.n2430 GNDA.n102 8126.25
R1351 GNDA.n1697 GNDA.n1637 7880
R1352 GNDA.n1697 GNDA.n1638 7880
R1353 GNDA.n1736 GNDA.n1610 7880
R1354 GNDA.n1732 GNDA.n1610 7880
R1355 GNDA.n1640 GNDA.n1637 7830.75
R1356 GNDA.n1640 GNDA.n1638 7830.75
R1357 GNDA.n1736 GNDA.n1611 7830.75
R1358 GNDA.n1732 GNDA.n1611 7830.75
R1359 GNDA.n106 GNDA.n100 7732.25
R1360 GNDA.n2472 GNDA.n40 7732.25
R1361 GNDA.n2472 GNDA.n41 7732.25
R1362 GNDA.n2474 GNDA.n40 7732.25
R1363 GNDA.n2474 GNDA.n41 7732.25
R1364 GNDA.n480 GNDA.n328 7732.25
R1365 GNDA.n472 GNDA.n328 7732.25
R1366 GNDA.n480 GNDA.n329 7732.25
R1367 GNDA.n472 GNDA.n329 7732.25
R1368 GNDA.n2430 GNDA.n100 7683
R1369 GNDA.n2177 GNDA.n313 6845.75
R1370 GNDA.n2181 GNDA.n313 6845.75
R1371 GNDA.n2177 GNDA.n312 6796.5
R1372 GNDA.n2181 GNDA.n312 6796.5
R1373 GNDA.n2175 GNDA.n492 6698
R1374 GNDA.n2170 GNDA.n492 6698
R1375 GNDA.n2175 GNDA.n491 6648.75
R1376 GNDA.n2170 GNDA.n491 6648.75
R1377 GNDA.n455 GNDA.n54 6057.75
R1378 GNDA.n2467 GNDA.n54 6057.75
R1379 GNDA.n455 GNDA.n47 6057.75
R1380 GNDA.n2467 GNDA.n47 6057.75
R1381 GNDA.n483 GNDA.n325 6057.75
R1382 GNDA.n465 GNDA.n325 6057.75
R1383 GNDA.n483 GNDA.n326 6057.75
R1384 GNDA.n465 GNDA.n326 6057.75
R1385 GNDA.n388 GNDA.n31 5713
R1386 GNDA.n391 GNDA.n32 5713
R1387 GNDA.n387 GNDA.n386 5446.53
R1388 GNDA.n343 GNDA.n317 5368.25
R1389 GNDA.n73 GNDA.n71 5368.25
R1390 GNDA.n343 GNDA.n318 5319
R1391 GNDA.n445 GNDA.n442 5319
R1392 GNDA.n424 GNDA.n423 5319
R1393 GNDA.n2452 GNDA.n71 5319
R1394 GNDA.n74 GNDA.n73 5319
R1395 GNDA.n488 GNDA.n318 5269.75
R1396 GNDA.n2452 GNDA.n74 5269.75
R1397 GNDA.n354 GNDA.n334 5171.25
R1398 GNDA.n2464 GNDA.n58 5171.25
R1399 GNDA.n2447 GNDA.n2446 5144.1
R1400 GNDA.n488 GNDA.n317 5122
R1401 GNDA.n336 GNDA.n334 5122
R1402 GNDA.n2460 GNDA.n58 5122
R1403 GNDA.n1695 GNDA.n1642 4974.25
R1404 GNDA.n1714 GNDA.n1628 4974.25
R1405 GNDA.n1718 GNDA.n1628 4974.25
R1406 GNDA.n354 GNDA.n353 4944.7
R1407 GNDA.n2464 GNDA.n59 4944.7
R1408 GNDA.n439 GNDA.n430 4925
R1409 GNDA.n439 GNDA.n431 4925
R1410 GNDA.n353 GNDA.n336 4895.45
R1411 GNDA.n2460 GNDA.n59 4895.45
R1412 GNDA.n430 GNDA.n378 4728
R1413 GNDA.n431 GNDA.n378 4728
R1414 GNDA.n2434 GNDA.n95 4678.75
R1415 GNDA.n2434 GNDA.n94 4629.5
R1416 GNDA.n166 GNDA.n95 4629.5
R1417 GNDA.n2444 GNDA.n83 4598.65
R1418 GNDA.n2156 GNDA.n506 4580.25
R1419 GNDA.n2156 GNDA.n507 4580.25
R1420 GNDA.n166 GNDA.n94 4580.25
R1421 GNDA.n2152 GNDA.n505 4580.25
R1422 GNDA.n515 GNDA.n505 4580.25
R1423 GNDA.n1729 GNDA.n1617 4531
R1424 GNDA.n1729 GNDA.n1618 4531
R1425 GNDA.n1617 GNDA.n1614 4531
R1426 GNDA.n1618 GNDA.n1614 4531
R1427 GNDA.n1714 GNDA.n1627 4531
R1428 GNDA.n1718 GNDA.n1627 4531
R1429 GNDA.n2123 GNDA.n506 4481.75
R1430 GNDA.n2123 GNDA.n507 4481.75
R1431 GNDA.n2152 GNDA.n512 4481.75
R1432 GNDA.n515 GNDA.n512 4481.75
R1433 GNDA.n490 GNDA.n489 4275.41
R1434 GNDA.n2445 GNDA.n2444 4159.38
R1435 GNDA.n386 GNDA.n385 3964.58
R1436 GNDA.n420 GNDA.n388 3595.25
R1437 GNDA.n2487 GNDA.n27 3349
R1438 GNDA.n427 GNDA.n27 3299.75
R1439 GNDA.n1685 GNDA.n1684 3287.9
R1440 GNDA.n420 GNDA.n391 3250.5
R1441 GNDA.n2487 GNDA.n28 3250.5
R1442 GNDA.n427 GNDA.n28 3201.25
R1443 GNDA.n1683 GNDA.n1682 3156.82
R1444 GNDA.n340 GNDA.n337 2326.02
R1445 GNDA.n350 GNDA.n337 2326.02
R1446 GNDA.n66 GNDA.n63 2326.02
R1447 GNDA.n76 GNDA.n63 2326.02
R1448 GNDA.n1678 GNDA.n1648 2142.38
R1449 GNDA.n1711 GNDA.n1626 2142.38
R1450 GNDA.n1648 GNDA.n1647 1846.88
R1451 GNDA.n1722 GNDA.n1626 1846.88
R1452 GNDA.n1683 GNDA.n78 1749.05
R1453 GNDA.n1847 GNDA.n602 1672.5
R1454 GNDA.n1684 GNDA.n1683 1226.55
R1455 GNDA.n422 GNDA.n387 1184.62
R1456 GNDA.n2449 GNDA.n78 1163.28
R1457 GNDA.n347 GNDA.n337 1114.8
R1458 GNDA.n2457 GNDA.n63 1114.8
R1459 GNDA.n746 GNDA.n619 1064.42
R1460 GNDA.n1444 GNDA.n592 1064.42
R1461 GNDA.n1426 GNDA.n619 1041.66
R1462 GNDA.n1871 GNDA.n592 1041.66
R1463 GNDA.n1675 GNDA.n1648 991.841
R1464 GNDA.n1706 GNDA.n1626 991.841
R1465 GNDA.n2176 GNDA.n316 991.54
R1466 GNDA.n2451 GNDA.n2450 971.551
R1467 GNDA.n2450 GNDA.n2449 890.324
R1468 GNDA.n82 GNDA.n78 831.111
R1469 GNDA.n1687 GNDA.n1631 803.201
R1470 GNDA.n1689 GNDA.n1631 800
R1471 GNDA.n1688 GNDA.n1687 774.4
R1472 GNDA.n1689 GNDA.n1688 771.201
R1473 GNDA.n462 GNDA.t105 734.418
R1474 GNDA.n322 GNDA.t92 734.418
R1475 GNDA.n48 GNDA.t97 734.418
R1476 GNDA.n51 GNDA.t80 734.418
R1477 GNDA.n447 GNDA.n446 691.201
R1478 GNDA.n383 GNDA.n375 691.201
R1479 GNDA.n2481 GNDA.t116 682.201
R1480 GNDA.n461 GNDA.n460 678.4
R1481 GNDA.n468 GNDA.n461 672
R1482 GNDA.n2075 GNDA.n548 669.307
R1483 GNDA.n416 GNDA.t130 666.134
R1484 GNDA.n2061 GNDA.n2060 662.155
R1485 GNDA.n2334 GNDA.n144 662.155
R1486 GNDA.n349 GNDA.n338 617.601
R1487 GNDA.n68 GNDA.n67 617.601
R1488 GNDA.n2483 GNDA.n33 601.601
R1489 GNDA.n422 GNDA.t165 592.308
R1490 GNDA.t162 GNDA.n57 592.308
R1491 GNDA.n2076 GNDA.n549 585
R1492 GNDA.n2078 GNDA.n2077 585
R1493 GNDA.n2079 GNDA.n2078 585
R1494 GNDA.n561 GNDA.n560 585
R1495 GNDA.n2062 GNDA.n561 585
R1496 GNDA.n2065 GNDA.n2064 585
R1497 GNDA.n2064 GNDA.n2063 585
R1498 GNDA.n2066 GNDA.n559 585
R1499 GNDA.n559 GNDA.n558 585
R1500 GNDA.n2068 GNDA.n2067 585
R1501 GNDA.n2069 GNDA.n2068 585
R1502 GNDA.n557 GNDA.n556 585
R1503 GNDA.n2070 GNDA.n557 585
R1504 GNDA.n2073 GNDA.n2072 585
R1505 GNDA.n2072 GNDA.n2071 585
R1506 GNDA.n547 GNDA.n546 585
R1507 GNDA.n2080 GNDA.n547 585
R1508 GNDA.n2083 GNDA.n2082 585
R1509 GNDA.n2082 GNDA.n2081 585
R1510 GNDA.n2084 GNDA.n545 585
R1511 GNDA.n545 GNDA.n544 585
R1512 GNDA.n2087 GNDA.n2086 585
R1513 GNDA.n2088 GNDA.n2087 585
R1514 GNDA.n2085 GNDA.n541 585
R1515 GNDA.n2089 GNDA.n541 585
R1516 GNDA.n2091 GNDA.n543 585
R1517 GNDA.n2091 GNDA.n2090 585
R1518 GNDA.n898 GNDA.n735 585
R1519 GNDA.n735 GNDA.n734 585
R1520 GNDA.n900 GNDA.n899 585
R1521 GNDA.n901 GNDA.n900 585
R1522 GNDA.n733 GNDA.n732 585
R1523 GNDA.n902 GNDA.n733 585
R1524 GNDA.n906 GNDA.n905 585
R1525 GNDA.n905 GNDA.n904 585
R1526 GNDA.n907 GNDA.n731 585
R1527 GNDA.n903 GNDA.n731 585
R1528 GNDA.n909 GNDA.n908 585
R1529 GNDA.n909 GNDA.n615 585
R1530 GNDA.n910 GNDA.n730 585
R1531 GNDA.n910 GNDA.n616 585
R1532 GNDA.n913 GNDA.n912 585
R1533 GNDA.n912 GNDA.n911 585
R1534 GNDA.n914 GNDA.n729 585
R1535 GNDA.n729 GNDA.n728 585
R1536 GNDA.n917 GNDA.n916 585
R1537 GNDA.n918 GNDA.n917 585
R1538 GNDA.n915 GNDA.n725 585
R1539 GNDA.n919 GNDA.n725 585
R1540 GNDA.n921 GNDA.n727 585
R1541 GNDA.n921 GNDA.n920 585
R1542 GNDA.n922 GNDA.n724 585
R1543 GNDA.n922 GNDA.n562 585
R1544 GNDA.n745 GNDA.n744 585
R1545 GNDA.n878 GNDA.n745 585
R1546 GNDA.n881 GNDA.n880 585
R1547 GNDA.n880 GNDA.n879 585
R1548 GNDA.n882 GNDA.n743 585
R1549 GNDA.n743 GNDA.n742 585
R1550 GNDA.n884 GNDA.n883 585
R1551 GNDA.n885 GNDA.n884 585
R1552 GNDA.n741 GNDA.n740 585
R1553 GNDA.n886 GNDA.n741 585
R1554 GNDA.n889 GNDA.n888 585
R1555 GNDA.n888 GNDA.n887 585
R1556 GNDA.n890 GNDA.n739 585
R1557 GNDA.n739 GNDA.n738 585
R1558 GNDA.n892 GNDA.n891 585
R1559 GNDA.n893 GNDA.n892 585
R1560 GNDA.n737 GNDA.n736 585
R1561 GNDA.n894 GNDA.n737 585
R1562 GNDA.n897 GNDA.n896 585
R1563 GNDA.n896 GNDA.n895 585
R1564 GNDA.n1417 GNDA.n1416 585
R1565 GNDA.n1443 GNDA.n1417 585
R1566 GNDA.n1441 GNDA.n1440 585
R1567 GNDA.n1442 GNDA.n1441 585
R1568 GNDA.n1439 GNDA.n1419 585
R1569 GNDA.n1419 GNDA.n1418 585
R1570 GNDA.n1438 GNDA.n1437 585
R1571 GNDA.n1437 GNDA.n1436 585
R1572 GNDA.n1421 GNDA.n1420 585
R1573 GNDA.n1435 GNDA.n1421 585
R1574 GNDA.n1433 GNDA.n1432 585
R1575 GNDA.n1434 GNDA.n1433 585
R1576 GNDA.n1431 GNDA.n1423 585
R1577 GNDA.n1423 GNDA.n1422 585
R1578 GNDA.n1430 GNDA.n1429 585
R1579 GNDA.n1429 GNDA.n1428 585
R1580 GNDA.n1425 GNDA.n1424 585
R1581 GNDA.n1427 GNDA.n1425 585
R1582 GNDA.n627 GNDA.n626 585
R1583 GNDA.n1426 GNDA.n626 585
R1584 GNDA.n1872 GNDA.n590 585
R1585 GNDA.n1872 GNDA.n1871 585
R1586 GNDA.n595 GNDA.n591 585
R1587 GNDA.n1870 GNDA.n591 585
R1588 GNDA.n1868 GNDA.n1867 585
R1589 GNDA.n1869 GNDA.n1868 585
R1590 GNDA.n1866 GNDA.n594 585
R1591 GNDA.n594 GNDA.n593 585
R1592 GNDA.n1865 GNDA.n1864 585
R1593 GNDA.n1864 GNDA.n1863 585
R1594 GNDA.n597 GNDA.n596 585
R1595 GNDA.n1862 GNDA.n597 585
R1596 GNDA.n1860 GNDA.n1859 585
R1597 GNDA.n1861 GNDA.n1860 585
R1598 GNDA.n1858 GNDA.n599 585
R1599 GNDA.n599 GNDA.n598 585
R1600 GNDA.n1857 GNDA.n1856 585
R1601 GNDA.n1856 GNDA.n1855 585
R1602 GNDA.n601 GNDA.n600 585
R1603 GNDA.n1854 GNDA.n601 585
R1604 GNDA.n1853 GNDA.n1852 585
R1605 GNDA.n603 GNDA.n602 585
R1606 GNDA.n1875 GNDA.n1874 585
R1607 GNDA.n1876 GNDA.n589 585
R1608 GNDA.n1878 GNDA.n1877 585
R1609 GNDA.n1880 GNDA.n588 585
R1610 GNDA.n1883 GNDA.n1882 585
R1611 GNDA.n1884 GNDA.n587 585
R1612 GNDA.n1886 GNDA.n1885 585
R1613 GNDA.n1888 GNDA.n586 585
R1614 GNDA.n1891 GNDA.n1890 585
R1615 GNDA.n1892 GNDA.n585 585
R1616 GNDA.n1894 GNDA.n1893 585
R1617 GNDA.n1896 GNDA.n583 585
R1618 GNDA.n1596 GNDA.n1595 585
R1619 GNDA.n1594 GNDA.n625 585
R1620 GNDA.n1593 GNDA.n1592 585
R1621 GNDA.n1591 GNDA.n1590 585
R1622 GNDA.n1589 GNDA.n1588 585
R1623 GNDA.n1587 GNDA.n1586 585
R1624 GNDA.n1585 GNDA.n1584 585
R1625 GNDA.n1583 GNDA.n1582 585
R1626 GNDA.n1581 GNDA.n1580 585
R1627 GNDA.n1579 GNDA.n1578 585
R1628 GNDA.n1577 GNDA.n1576 585
R1629 GNDA.n1575 GNDA.n1574 585
R1630 GNDA.n953 GNDA.n952 585
R1631 GNDA.n941 GNDA.n714 585
R1632 GNDA.n942 GNDA.n717 585
R1633 GNDA.n945 GNDA.n944 585
R1634 GNDA.n940 GNDA.n719 585
R1635 GNDA.n938 GNDA.n937 585
R1636 GNDA.n721 GNDA.n720 585
R1637 GNDA.n931 GNDA.n930 585
R1638 GNDA.n928 GNDA.n723 585
R1639 GNDA.n926 GNDA.n925 585
R1640 GNDA.n1555 GNDA.n649 585
R1641 GNDA.n1556 GNDA.n647 585
R1642 GNDA.n1557 GNDA.n646 585
R1643 GNDA.n644 GNDA.n642 585
R1644 GNDA.n1563 GNDA.n641 585
R1645 GNDA.n1564 GNDA.n639 585
R1646 GNDA.n1565 GNDA.n638 585
R1647 GNDA.n636 GNDA.n634 585
R1648 GNDA.n1570 GNDA.n633 585
R1649 GNDA.n1571 GNDA.n631 585
R1650 GNDA.n567 GNDA.n564 585
R1651 GNDA.n1927 GNDA.n1926 585
R1652 GNDA.n571 GNDA.n570 585
R1653 GNDA.n1917 GNDA.n573 585
R1654 GNDA.n1919 GNDA.n1918 585
R1655 GNDA.n1914 GNDA.n575 585
R1656 GNDA.n1913 GNDA.n1912 585
R1657 GNDA.n1904 GNDA.n577 585
R1658 GNDA.n1906 GNDA.n1905 585
R1659 GNDA.n1902 GNDA.n579 585
R1660 GNDA.n1901 GNDA.n1900 585
R1661 GNDA.n1901 GNDA.n564 585
R1662 GNDA.n925 GNDA.n924 585
R1663 GNDA.n723 GNDA.n722 585
R1664 GNDA.n932 GNDA.n931 585
R1665 GNDA.n934 GNDA.n721 585
R1666 GNDA.n937 GNDA.n936 585
R1667 GNDA.n719 GNDA.n718 585
R1668 GNDA.n946 GNDA.n945 585
R1669 GNDA.n948 GNDA.n717 585
R1670 GNDA.n949 GNDA.n714 585
R1671 GNDA.n952 GNDA.n951 585
R1672 GNDA.n1573 GNDA.n629 585
R1673 GNDA.n1573 GNDA.n582 585
R1674 GNDA.n1572 GNDA.n1571 585
R1675 GNDA.n1570 GNDA.n1569 585
R1676 GNDA.n1568 GNDA.n634 585
R1677 GNDA.n1566 GNDA.n1565 585
R1678 GNDA.n1564 GNDA.n635 585
R1679 GNDA.n1563 GNDA.n1562 585
R1680 GNDA.n1560 GNDA.n642 585
R1681 GNDA.n1558 GNDA.n1557 585
R1682 GNDA.n1556 GNDA.n643 585
R1683 GNDA.n1555 GNDA.n1554 585
R1684 GNDA.n1897 GNDA.n581 585
R1685 GNDA.n1897 GNDA.n582 585
R1686 GNDA.n1900 GNDA.n1899 585
R1687 GNDA.n579 GNDA.n578 585
R1688 GNDA.n1907 GNDA.n1906 585
R1689 GNDA.n1909 GNDA.n577 585
R1690 GNDA.n1912 GNDA.n1911 585
R1691 GNDA.n575 GNDA.n574 585
R1692 GNDA.n1920 GNDA.n1919 585
R1693 GNDA.n1922 GNDA.n573 585
R1694 GNDA.n1923 GNDA.n571 585
R1695 GNDA.n1926 GNDA.n1925 585
R1696 GNDA.n572 GNDA.n563 585
R1697 GNDA.n1814 GNDA.n563 585
R1698 GNDA.n1215 GNDA.n580 585
R1699 GNDA.n1266 GNDA.n1265 585
R1700 GNDA.n1264 GNDA.n1214 585
R1701 GNDA.n1263 GNDA.n1262 585
R1702 GNDA.n1261 GNDA.n1260 585
R1703 GNDA.n1259 GNDA.n1258 585
R1704 GNDA.n1257 GNDA.n1256 585
R1705 GNDA.n1255 GNDA.n1254 585
R1706 GNDA.n1253 GNDA.n1252 585
R1707 GNDA.n1251 GNDA.n1250 585
R1708 GNDA.n1249 GNDA.n1248 585
R1709 GNDA.n1247 GNDA.n1246 585
R1710 GNDA.n683 GNDA.n682 585
R1711 GNDA.n681 GNDA.n660 585
R1712 GNDA.n680 GNDA.n679 585
R1713 GNDA.n678 GNDA.n677 585
R1714 GNDA.n676 GNDA.n675 585
R1715 GNDA.n674 GNDA.n673 585
R1716 GNDA.n672 GNDA.n671 585
R1717 GNDA.n670 GNDA.n669 585
R1718 GNDA.n668 GNDA.n667 585
R1719 GNDA.n666 GNDA.n665 585
R1720 GNDA.n664 GNDA.n663 585
R1721 GNDA.n662 GNDA.n661 585
R1722 GNDA.n2327 GNDA.n145 585
R1723 GNDA.n1226 GNDA.n147 585
R1724 GNDA.n1227 GNDA.n1224 585
R1725 GNDA.n1230 GNDA.n1223 585
R1726 GNDA.n1231 GNDA.n1222 585
R1727 GNDA.n1234 GNDA.n1221 585
R1728 GNDA.n1235 GNDA.n1220 585
R1729 GNDA.n1238 GNDA.n1219 585
R1730 GNDA.n1239 GNDA.n1218 585
R1731 GNDA.n1242 GNDA.n1217 585
R1732 GNDA.n1243 GNDA.n160 585
R1733 GNDA.n2327 GNDA.n160 585
R1734 GNDA.n1245 GNDA.n1216 585
R1735 GNDA.n1245 GNDA.n186 585
R1736 GNDA.n1244 GNDA.n1243 585
R1737 GNDA.n1242 GNDA.n1241 585
R1738 GNDA.n1240 GNDA.n1239 585
R1739 GNDA.n1238 GNDA.n1237 585
R1740 GNDA.n1236 GNDA.n1235 585
R1741 GNDA.n1234 GNDA.n1233 585
R1742 GNDA.n1232 GNDA.n1231 585
R1743 GNDA.n1230 GNDA.n1229 585
R1744 GNDA.n1228 GNDA.n1227 585
R1745 GNDA.n1226 GNDA.n1225 585
R1746 GNDA.n2296 GNDA.n198 585
R1747 GNDA.n2296 GNDA.n204 585
R1748 GNDA.n1199 GNDA.n1075 585
R1749 GNDA.n1073 GNDA.n1070 585
R1750 GNDA.n1069 GNDA.n1068 585
R1751 GNDA.n1067 GNDA.n1064 585
R1752 GNDA.n1063 GNDA.n1062 585
R1753 GNDA.n1061 GNDA.n1058 585
R1754 GNDA.n1057 GNDA.n1056 585
R1755 GNDA.n1055 GNDA.n1052 585
R1756 GNDA.n1051 GNDA.n539 585
R1757 GNDA.n2095 GNDA.n2094 585
R1758 GNDA.n2092 GNDA.n538 585
R1759 GNDA.n2092 GNDA.n540 585
R1760 GNDA.n2094 GNDA.n2093 585
R1761 GNDA.n1053 GNDA.n539 585
R1762 GNDA.n1055 GNDA.n1054 585
R1763 GNDA.n1059 GNDA.n1056 585
R1764 GNDA.n1061 GNDA.n1060 585
R1765 GNDA.n1065 GNDA.n1062 585
R1766 GNDA.n1067 GNDA.n1066 585
R1767 GNDA.n1071 GNDA.n1068 585
R1768 GNDA.n1073 GNDA.n1072 585
R1769 GNDA.n1075 GNDA.n1074 585
R1770 GNDA.n2096 GNDA.n537 585
R1771 GNDA.n2097 GNDA.n2096 585
R1772 GNDA.n2100 GNDA.n2099 585
R1773 GNDA.n2099 GNDA.n2098 585
R1774 GNDA.n2101 GNDA.n536 585
R1775 GNDA.n536 GNDA.n535 585
R1776 GNDA.n2103 GNDA.n2102 585
R1777 GNDA.n2104 GNDA.n2103 585
R1778 GNDA.n534 GNDA.n533 585
R1779 GNDA.n2105 GNDA.n534 585
R1780 GNDA.n2108 GNDA.n2107 585
R1781 GNDA.n2107 GNDA.n2106 585
R1782 GNDA.n2109 GNDA.n532 585
R1783 GNDA.n532 GNDA.n531 585
R1784 GNDA.n2111 GNDA.n2110 585
R1785 GNDA.n2112 GNDA.n2111 585
R1786 GNDA.n530 GNDA.n529 585
R1787 GNDA.n2113 GNDA.n530 585
R1788 GNDA.n2117 GNDA.n2116 585
R1789 GNDA.n2116 GNDA.n2115 585
R1790 GNDA.n2118 GNDA.n528 585
R1791 GNDA.n2114 GNDA.n528 585
R1792 GNDA.n2120 GNDA.n2119 585
R1793 GNDA.n2120 GNDA.n316 585
R1794 GNDA.n1201 GNDA.n1076 585
R1795 GNDA.n1201 GNDA.n1200 585
R1796 GNDA.n1102 GNDA.n1101 585
R1797 GNDA.n1097 GNDA.n1096 585
R1798 GNDA.n1173 GNDA.n1172 585
R1799 GNDA.n1176 GNDA.n1175 585
R1800 GNDA.n1095 GNDA.n1092 585
R1801 GNDA.n1088 GNDA.n1087 585
R1802 GNDA.n1184 GNDA.n1183 585
R1803 GNDA.n1187 GNDA.n1186 585
R1804 GNDA.n1086 GNDA.n1083 585
R1805 GNDA.n1079 GNDA.n1078 585
R1806 GNDA.n1195 GNDA.n1194 585
R1807 GNDA.n1198 GNDA.n1197 585
R1808 GNDA.n956 GNDA.n564 585
R1809 GNDA.n954 GNDA.n564 585
R1810 GNDA.n1206 GNDA.n1205 585
R1811 GNDA.n1048 GNDA.n691 585
R1812 GNDA.n695 GNDA.n694 585
R1813 GNDA.n972 GNDA.n971 585
R1814 GNDA.n974 GNDA.n973 585
R1815 GNDA.n978 GNDA.n977 585
R1816 GNDA.n976 GNDA.n962 585
R1817 GNDA.n985 GNDA.n984 585
R1818 GNDA.n987 GNDA.n986 585
R1819 GNDA.n991 GNDA.n990 585
R1820 GNDA.n989 GNDA.n960 585
R1821 GNDA.n958 GNDA.n957 585
R1822 GNDA.n1204 GNDA.n692 585
R1823 GNDA.n692 GNDA.n186 585
R1824 GNDA.n2296 GNDA.n192 585
R1825 GNDA.n2296 GNDA.n205 585
R1826 GNDA.n874 GNDA.n746 585
R1827 GNDA.n877 GNDA.n876 585
R1828 GNDA.n778 GNDA.n777 585
R1829 GNDA.n769 GNDA.n768 585
R1830 GNDA.n849 GNDA.n848 585
R1831 GNDA.n852 GNDA.n851 585
R1832 GNDA.n767 GNDA.n764 585
R1833 GNDA.n760 GNDA.n759 585
R1834 GNDA.n860 GNDA.n859 585
R1835 GNDA.n863 GNDA.n862 585
R1836 GNDA.n758 GNDA.n755 585
R1837 GNDA.n751 GNDA.n749 585
R1838 GNDA.n871 GNDA.n870 585
R1839 GNDA.n873 GNDA.n748 585
R1840 GNDA.n776 GNDA.n771 585
R1841 GNDA.n776 GNDA.n582 585
R1842 GNDA.n716 GNDA.n563 585
R1843 GNDA.n775 GNDA.n563 585
R1844 GNDA.n2289 GNDA.n280 585
R1845 GNDA.n278 GNDA.n275 585
R1846 GNDA.n274 GNDA.n273 585
R1847 GNDA.n272 GNDA.n269 585
R1848 GNDA.n268 GNDA.n267 585
R1849 GNDA.n266 GNDA.n263 585
R1850 GNDA.n262 GNDA.n261 585
R1851 GNDA.n260 GNDA.n258 585
R1852 GNDA.n257 GNDA.n183 585
R1853 GNDA.n2300 GNDA.n2299 585
R1854 GNDA.n184 GNDA.n182 585
R1855 GNDA.n186 GNDA.n184 585
R1856 GNDA.n2299 GNDA.n2298 585
R1857 GNDA.n185 GNDA.n183 585
R1858 GNDA.n260 GNDA.n259 585
R1859 GNDA.n264 GNDA.n261 585
R1860 GNDA.n266 GNDA.n265 585
R1861 GNDA.n270 GNDA.n267 585
R1862 GNDA.n272 GNDA.n271 585
R1863 GNDA.n276 GNDA.n273 585
R1864 GNDA.n278 GNDA.n277 585
R1865 GNDA.n280 GNDA.n279 585
R1866 GNDA.n2303 GNDA.n2302 585
R1867 GNDA.n2304 GNDA.n180 585
R1868 GNDA.n2306 GNDA.n2305 585
R1869 GNDA.n2308 GNDA.n179 585
R1870 GNDA.n2311 GNDA.n2310 585
R1871 GNDA.n2312 GNDA.n178 585
R1872 GNDA.n2314 GNDA.n2313 585
R1873 GNDA.n2316 GNDA.n177 585
R1874 GNDA.n2319 GNDA.n2318 585
R1875 GNDA.n2320 GNDA.n176 585
R1876 GNDA.n2322 GNDA.n2321 585
R1877 GNDA.n2324 GNDA.n175 585
R1878 GNDA.n2291 GNDA.n281 585
R1879 GNDA.n2291 GNDA.n2290 585
R1880 GNDA.n654 GNDA.n564 585
R1881 GNDA.n651 GNDA.n564 585
R1882 GNDA.n1293 GNDA.n1292 585
R1883 GNDA.n1289 GNDA.n1288 585
R1884 GNDA.n1364 GNDA.n1363 585
R1885 GNDA.n1367 GNDA.n1366 585
R1886 GNDA.n1287 GNDA.n1284 585
R1887 GNDA.n1280 GNDA.n1279 585
R1888 GNDA.n1375 GNDA.n1374 585
R1889 GNDA.n1378 GNDA.n1377 585
R1890 GNDA.n1278 GNDA.n1275 585
R1891 GNDA.n1271 GNDA.n1270 585
R1892 GNDA.n1386 GNDA.n1385 585
R1893 GNDA.n1389 GNDA.n1388 585
R1894 GNDA.n207 GNDA.n206 585
R1895 GNDA.n206 GNDA.n186 585
R1896 GNDA.n2296 GNDA.n187 585
R1897 GNDA.n2296 GNDA.n2295 585
R1898 GNDA.n1444 GNDA.n1415 585
R1899 GNDA.n1446 GNDA.n1445 585
R1900 GNDA.n1547 GNDA.n1393 585
R1901 GNDA.n1545 GNDA.n1544 585
R1902 GNDA.n1466 GNDA.n1394 585
R1903 GNDA.n1464 GNDA.n1463 585
R1904 GNDA.n1473 GNDA.n1472 585
R1905 GNDA.n1476 GNDA.n1475 585
R1906 GNDA.n1461 GNDA.n1458 585
R1907 GNDA.n1454 GNDA.n1453 585
R1908 GNDA.n1484 GNDA.n1483 585
R1909 GNDA.n1487 GNDA.n1486 585
R1910 GNDA.n1452 GNDA.n1413 585
R1911 GNDA.n1450 GNDA.n1449 585
R1912 GNDA.n1549 GNDA.n1548 585
R1913 GNDA.n1548 GNDA.n582 585
R1914 GNDA.n1552 GNDA.n563 585
R1915 GNDA.n1392 GNDA.n563 585
R1916 GNDA.n2192 GNDA.n2191 585
R1917 GNDA.n302 GNDA.n301 585
R1918 GNDA.n2263 GNDA.n2262 585
R1919 GNDA.n2266 GNDA.n2265 585
R1920 GNDA.n300 GNDA.n297 585
R1921 GNDA.n293 GNDA.n292 585
R1922 GNDA.n2274 GNDA.n2273 585
R1923 GNDA.n2277 GNDA.n2276 585
R1924 GNDA.n291 GNDA.n288 585
R1925 GNDA.n284 GNDA.n283 585
R1926 GNDA.n2285 GNDA.n2284 585
R1927 GNDA.n2288 GNDA.n2287 585
R1928 GNDA.n255 GNDA.n254 585
R1929 GNDA.n252 GNDA.n208 585
R1930 GNDA.n251 GNDA.n250 585
R1931 GNDA.n249 GNDA.n248 585
R1932 GNDA.n247 GNDA.n210 585
R1933 GNDA.n245 GNDA.n244 585
R1934 GNDA.n243 GNDA.n211 585
R1935 GNDA.n242 GNDA.n241 585
R1936 GNDA.n239 GNDA.n212 585
R1937 GNDA.n237 GNDA.n236 585
R1938 GNDA.n235 GNDA.n213 585
R1939 GNDA.n234 GNDA.n233 585
R1940 GNDA.n1099 GNDA.n519 585
R1941 GNDA.n1099 GNDA.n171 585
R1942 GNDA.n2121 GNDA.n527 585
R1943 GNDA.n2122 GNDA.n2121 585
R1944 GNDA.n2127 GNDA.n2126 585
R1945 GNDA.n2126 GNDA.n2125 585
R1946 GNDA.n2128 GNDA.n526 585
R1947 GNDA.n526 GNDA.n525 585
R1948 GNDA.n2130 GNDA.n2129 585
R1949 GNDA.n2131 GNDA.n2130 585
R1950 GNDA.n524 GNDA.n523 585
R1951 GNDA.n2132 GNDA.n524 585
R1952 GNDA.n2136 GNDA.n2135 585
R1953 GNDA.n2135 GNDA.n2134 585
R1954 GNDA.n2137 GNDA.n522 585
R1955 GNDA.n2133 GNDA.n522 585
R1956 GNDA.n2139 GNDA.n2138 585
R1957 GNDA.n2140 GNDA.n2139 585
R1958 GNDA.n521 GNDA.n520 585
R1959 GNDA.n2141 GNDA.n521 585
R1960 GNDA.n2144 GNDA.n2143 585
R1961 GNDA.n2143 GNDA.n2142 585
R1962 GNDA.n2145 GNDA.n517 585
R1963 GNDA.n517 GNDA.n513 585
R1964 GNDA.n2149 GNDA.n2148 585
R1965 GNDA.n518 GNDA.n516 585
R1966 GNDA.n2190 GNDA.n304 585
R1967 GNDA.n2190 GNDA.n168 585
R1968 GNDA.n2325 GNDA.n173 585
R1969 GNDA.n2326 GNDA.n2325 585
R1970 GNDA.n500 GNDA.n174 585
R1971 GNDA.n174 GNDA.n172 585
R1972 GNDA.n501 GNDA.n499 585
R1973 GNDA.n499 GNDA.n498 585
R1974 GNDA.n503 GNDA.n502 585
R1975 GNDA.n504 GNDA.n503 585
R1976 GNDA.n497 GNDA.n496 585
R1977 GNDA.n2158 GNDA.n497 585
R1978 GNDA.n2162 GNDA.n2161 585
R1979 GNDA.n2161 GNDA.n2160 585
R1980 GNDA.n2163 GNDA.n494 585
R1981 GNDA.n2159 GNDA.n494 585
R1982 GNDA.n2167 GNDA.n2166 585
R1983 GNDA.n2168 GNDA.n2167 585
R1984 GNDA.n2165 GNDA.n495 585
R1985 GNDA.n495 GNDA.n311 585
R1986 GNDA.n2164 GNDA.n308 585
R1987 GNDA.n2183 GNDA.n308 585
R1988 GNDA.n2185 GNDA.n310 585
R1989 GNDA.n2185 GNDA.n2184 585
R1990 GNDA.n2187 GNDA.n2186 585
R1991 GNDA.n2189 GNDA.n2188 585
R1992 GNDA.n2438 GNDA.n2437 585
R1993 GNDA.n2437 GNDA.n2436 585
R1994 GNDA.n231 GNDA.n214 585
R1995 GNDA.n231 GNDA.n215 585
R1996 GNDA.n230 GNDA.n217 585
R1997 GNDA.n230 GNDA.n229 585
R1998 GNDA.n220 GNDA.n216 585
R1999 GNDA.n228 GNDA.n216 585
R2000 GNDA.n226 GNDA.n225 585
R2001 GNDA.n227 GNDA.n226 585
R2002 GNDA.n224 GNDA.n219 585
R2003 GNDA.n219 GNDA.n218 585
R2004 GNDA.n223 GNDA.n222 585
R2005 GNDA.n222 GNDA.n221 585
R2006 GNDA.n114 GNDA.n113 585
R2007 GNDA.n116 GNDA.n114 585
R2008 GNDA.n2423 GNDA.n2422 585
R2009 GNDA.n2422 GNDA.n2421 585
R2010 GNDA.n2424 GNDA.n108 585
R2011 GNDA.n108 GNDA.n103 585
R2012 GNDA.n2427 GNDA.n2426 585
R2013 GNDA.n2428 GNDA.n2427 585
R2014 GNDA.n2425 GNDA.n112 585
R2015 GNDA.n112 GNDA.n107 585
R2016 GNDA.n111 GNDA.n110 585
R2017 GNDA.n92 GNDA.n91 585
R2018 GNDA.n2439 GNDA.n87 585
R2019 GNDA.n87 GNDA.n85 585
R2020 GNDA.n2442 GNDA.n2441 585
R2021 GNDA.n2443 GNDA.n2442 585
R2022 GNDA.n2408 GNDA.n86 585
R2023 GNDA.n86 GNDA.n84 585
R2024 GNDA.n2412 GNDA.n2411 585
R2025 GNDA.n2411 GNDA.n2410 585
R2026 GNDA.n123 GNDA.n121 585
R2027 GNDA.n121 GNDA.n119 585
R2028 GNDA.n2419 GNDA.n2418 585
R2029 GNDA.n2420 GNDA.n2419 585
R2030 GNDA.n2338 GNDA.n120 585
R2031 GNDA.n120 GNDA.n118 585
R2032 GNDA.n2345 GNDA.n2344 585
R2033 GNDA.n2346 GNDA.n2345 585
R2034 GNDA.n2336 GNDA.n143 585
R2035 GNDA.n2347 GNDA.n143 585
R2036 GNDA.n2350 GNDA.n2349 585
R2037 GNDA.n2349 GNDA.n2348 585
R2038 GNDA.n142 GNDA.n140 585
R2039 GNDA.n2335 GNDA.n142 585
R2040 GNDA.n2333 GNDA.n2332 585
R2041 GNDA.n2334 GNDA.n2333 585
R2042 GNDA.n2026 GNDA.n1951 585
R2043 GNDA.n1951 GNDA.n1950 585
R2044 GNDA.n2029 GNDA.n2028 585
R2045 GNDA.n2030 GNDA.n2029 585
R2046 GNDA.n1952 GNDA.n1947 585
R2047 GNDA.n2031 GNDA.n1947 585
R2048 GNDA.n2034 GNDA.n2033 585
R2049 GNDA.n2033 GNDA.n2032 585
R2050 GNDA.n1946 GNDA.n1944 585
R2051 GNDA.n1949 GNDA.n1946 585
R2052 GNDA.n1940 GNDA.n1939 585
R2053 GNDA.n1948 GNDA.n1939 585
R2054 GNDA.n2042 GNDA.n2041 585
R2055 GNDA.n2046 GNDA.n2042 585
R2056 GNDA.n2049 GNDA.n2048 585
R2057 GNDA.n2048 GNDA.n2047 585
R2058 GNDA.n1938 GNDA.n1936 585
R2059 GNDA.n2045 GNDA.n1938 585
R2060 GNDA.n2043 GNDA.n1932 585
R2061 GNDA.n2044 GNDA.n2043 585
R2062 GNDA.n2056 GNDA.n568 585
R2063 GNDA.n568 GNDA.n566 585
R2064 GNDA.n2059 GNDA.n2058 585
R2065 GNDA.n2060 GNDA.n2059 585
R2066 GNDA.n2025 GNDA.n2024 585
R2067 GNDA.n2024 GNDA.n2023 585
R2068 GNDA.n1817 GNDA.n1740 585
R2069 GNDA.n1740 GNDA.n1739 585
R2070 GNDA.n1820 GNDA.n1819 585
R2071 GNDA.n1821 GNDA.n1820 585
R2072 GNDA.n1741 GNDA.n1608 585
R2073 GNDA.n1822 GNDA.n1608 585
R2074 GNDA.n1825 GNDA.n1824 585
R2075 GNDA.n1824 GNDA.n1823 585
R2076 GNDA.n1603 GNDA.n1600 585
R2077 GNDA.n1600 GNDA.n1599 585
R2078 GNDA.n1832 GNDA.n1831 585
R2079 GNDA.n1833 GNDA.n1832 585
R2080 GNDA.n1601 GNDA.n614 585
R2081 GNDA.n1834 GNDA.n614 585
R2082 GNDA.n1837 GNDA.n1836 585
R2083 GNDA.n1836 GNDA.n1835 585
R2084 GNDA.n610 GNDA.n607 585
R2085 GNDA.n607 GNDA.n606 585
R2086 GNDA.n1844 GNDA.n1843 585
R2087 GNDA.n1845 GNDA.n1844 585
R2088 GNDA.n608 GNDA.n605 585
R2089 GNDA.n1846 GNDA.n605 585
R2090 GNDA.n1849 GNDA.n1848 585
R2091 GNDA.n1848 GNDA.n1847 585
R2092 GNDA.n1816 GNDA.n1815 585
R2093 GNDA.n1815 GNDA.n565 585
R2094 GNDA.n1738 GNDA.n1737 556.322
R2095 GNDA.n357 GNDA.t133 535.191
R2096 GNDA.n330 GNDA.t143 535.191
R2097 GNDA.n44 GNDA.t170 535.191
R2098 GNDA.n42 GNDA.t89 535.191
R2099 GNDA.n895 GNDA.n734 534.218
R2100 GNDA.n105 GNDA.n99 531.201
R2101 GNDA.n2431 GNDA.n99 528
R2102 GNDA.n895 GNDA.n894 512.29
R2103 GNDA.n894 GNDA.n893 512.29
R2104 GNDA.n893 GNDA.n738 512.29
R2105 GNDA.n887 GNDA.n738 512.29
R2106 GNDA.n887 GNDA.n886 512.29
R2107 GNDA.n885 GNDA.n742 512.29
R2108 GNDA.n879 GNDA.n742 512.29
R2109 GNDA.n879 GNDA.n878 512.29
R2110 GNDA.n878 GNDA.n877 512.29
R2111 GNDA.n877 GNDA.n746 512.29
R2112 GNDA.n1427 GNDA.n1426 512.29
R2113 GNDA.n1428 GNDA.n1427 512.29
R2114 GNDA.n1428 GNDA.n1422 512.29
R2115 GNDA.n1434 GNDA.n1422 512.29
R2116 GNDA.n1435 GNDA.n1434 512.29
R2117 GNDA.n1436 GNDA.n1418 512.29
R2118 GNDA.n1442 GNDA.n1418 512.29
R2119 GNDA.n1443 GNDA.n1442 512.29
R2120 GNDA.n1445 GNDA.n1443 512.29
R2121 GNDA.n1445 GNDA.n1444 512.29
R2122 GNDA.n1871 GNDA.n1870 512.29
R2123 GNDA.n1870 GNDA.n1869 512.29
R2124 GNDA.n1869 GNDA.n593 512.29
R2125 GNDA.n1863 GNDA.n593 512.29
R2126 GNDA.n1863 GNDA.n1862 512.29
R2127 GNDA.n1861 GNDA.n598 512.29
R2128 GNDA.n1855 GNDA.n598 512.29
R2129 GNDA.n1855 GNDA.n1854 512.29
R2130 GNDA.n1854 GNDA.n1853 512.29
R2131 GNDA.n1853 GNDA.n602 512.29
R2132 GNDA.n1698 GNDA.n1635 512
R2133 GNDA.n1698 GNDA.n1636 512
R2134 GNDA.n1733 GNDA.n1612 512
R2135 GNDA.n1735 GNDA.n1612 512
R2136 GNDA.n1639 GNDA.n1635 508.8
R2137 GNDA.n1639 GNDA.n1636 508.8
R2138 GNDA.n1734 GNDA.n1733 508.8
R2139 GNDA.n1735 GNDA.n1734 508.8
R2140 GNDA.n105 GNDA.n104 499.2
R2141 GNDA.t96 GNDA.n117 496.098
R2142 GNDA.n478 GNDA.n473 496
R2143 GNDA.n2475 GNDA.n38 496
R2144 GNDA.n443 GNDA.t161 493.418
R2145 GNDA.n376 GNDA.t149 493.418
R2146 GNDA.n380 GNDA.t86 493.418
R2147 GNDA.n379 GNDA.t164 493.418
R2148 GNDA.n370 GNDA.t102 493.418
R2149 GNDA.n371 GNDA.t83 493.418
R2150 GNDA.n365 GNDA.t158 493.418
R2151 GNDA.n367 GNDA.t174 493.418
R2152 GNDA.n368 GNDA.t155 493.418
R2153 GNDA.n369 GNDA.t146 493.418
R2154 GNDA.n479 GNDA.n478 489.601
R2155 GNDA.n2475 GNDA.n39 489.601
R2156 GNDA.n2446 GNDA.n81 488.889
R2157 GNDA.n2431 GNDA.n98 486.401
R2158 GNDA.n471 GNDA.n470 463.603
R2159 GNDA.n458 GNDA.n457 463.603
R2160 GNDA.n2179 GNDA.n2178 444.8
R2161 GNDA.n2180 GNDA.n2179 444.8
R2162 GNDA.n2180 GNDA.n314 441.601
R2163 GNDA.n2178 GNDA.n315 438.401
R2164 GNDA.n2174 GNDA.n2173 435.2
R2165 GNDA.n2061 GNDA.n565 434.906
R2166 GNDA.n2023 GNDA.n144 434.906
R2167 GNDA.n2482 GNDA.n34 428.8
R2168 GNDA.n2174 GNDA.n493 425.601
R2169 GNDA.n2172 GNDA.n2171 422.401
R2170 GNDA.n444 GNDA.n377 422.401
R2171 GNDA.n382 GNDA.n381 422.401
R2172 GNDA.n372 GNDA.n366 422.401
R2173 GNDA.n453 GNDA.n452 422.401
R2174 GNDA.n2171 GNDA.n493 419.2
R2175 GNDA.n1649 GNDA.t140 413.084
R2176 GNDA.n1650 GNDA.t136 413.084
R2177 GNDA.n1621 GNDA.t127 413.084
R2178 GNDA.n1619 GNDA.t110 413.084
R2179 GNDA.n1623 GNDA.t152 413.084
R2180 GNDA.n1708 GNDA.t167 413.084
R2181 GNDA.n2469 GNDA.n46 387.2
R2182 GNDA.n1694 GNDA.n1693 383.118
R2183 GNDA.n484 GNDA.n324 380.8
R2184 GNDA.n2469 GNDA.n2468 380.8
R2185 GNDA.t165 GNDA.t242 372.308
R2186 GNDA.t241 GNDA.t247 372.308
R2187 GNDA.t243 GNDA.t241 372.308
R2188 GNDA.t243 GNDA.t248 372.308
R2189 GNDA.t248 GNDA.t246 372.308
R2190 GNDA.t246 GNDA.t240 372.308
R2191 GNDA.t302 GNDA.t305 372.308
R2192 GNDA.t300 GNDA.t306 372.308
R2193 GNDA.t26 GNDA.t234 372.308
R2194 GNDA.t234 GNDA.t236 372.308
R2195 GNDA.t329 GNDA.t206 372.308
R2196 GNDA.t206 GNDA.t23 372.308
R2197 GNDA.t23 GNDA.t324 372.308
R2198 GNDA.n392 GNDA.n33 371.2
R2199 GNDA.n417 GNDA.n34 371.2
R2200 GNDA.n592 GNDA.n584 370.214
R2201 GNDA.n1598 GNDA.n619 370.214
R2202 GNDA.n617 GNDA.n592 365.957
R2203 GNDA.n619 GNDA.n618 365.957
R2204 GNDA.n429 GNDA.t245 355.385
R2205 GNDA.t307 GNDA.n425 355.385
R2206 GNDA.n441 GNDA.t301 355.385
R2207 GNDA.t37 GNDA.n29 355.385
R2208 GNDA.t236 GNDA.n30 355.385
R2209 GNDA.n1713 GNDA.n1609 354.024
R2210 GNDA.n1847 GNDA.n1846 352.627
R2211 GNDA.n1846 GNDA.n1845 352.627
R2212 GNDA.n1845 GNDA.n606 352.627
R2213 GNDA.n1835 GNDA.n606 352.627
R2214 GNDA.n1835 GNDA.n1834 352.627
R2215 GNDA.n1833 GNDA.n1599 352.627
R2216 GNDA.n1823 GNDA.n1599 352.627
R2217 GNDA.n1823 GNDA.n1822 352.627
R2218 GNDA.n1822 GNDA.n1821 352.627
R2219 GNDA.n1739 GNDA.n565 352.627
R2220 GNDA.n2060 GNDA.n566 352.627
R2221 GNDA.n2044 GNDA.n566 352.627
R2222 GNDA.n2045 GNDA.n2044 352.627
R2223 GNDA.n2047 GNDA.n2045 352.627
R2224 GNDA.n2047 GNDA.n2046 352.627
R2225 GNDA.n1949 GNDA.n1948 352.627
R2226 GNDA.n2032 GNDA.n1949 352.627
R2227 GNDA.n2032 GNDA.n2031 352.627
R2228 GNDA.n2031 GNDA.n2030 352.627
R2229 GNDA.n2030 GNDA.n1950 352.627
R2230 GNDA.n2023 GNDA.n1950 352.627
R2231 GNDA.n2335 GNDA.n2334 352.627
R2232 GNDA.n2348 GNDA.n2335 352.627
R2233 GNDA.n2348 GNDA.n2347 352.627
R2234 GNDA.n2347 GNDA.n2346 352.627
R2235 GNDA.n2346 GNDA.n118 352.627
R2236 GNDA.n2420 GNDA.n119 352.627
R2237 GNDA.n321 GNDA.n320 348.8
R2238 GNDA.n72 GNDA.n69 348.8
R2239 GNDA.n2410 GNDA.n84 343.452
R2240 GNDA.n2443 GNDA.n85 343.452
R2241 GNDA.n487 GNDA.n486 342.401
R2242 GNDA.n2453 GNDA.n70 342.401
R2243 GNDA.n1692 GNDA.n1691 341.38
R2244 GNDA.n335 GNDA.n332 332.8
R2245 GNDA.n2461 GNDA.n61 332.8
R2246 GNDA.n435 GNDA.t120 332.75
R2247 GNDA.n432 GNDA.t123 332.75
R2248 GNDA.t96 GNDA.n165 172.876
R2249 GNDA.t109 GNDA.n617 327.661
R2250 GNDA.t109 GNDA.n618 327.661
R2251 GNDA.n1269 GNDA.t101 172.876
R2252 GNDA.n1208 GNDA.t101 172.876
R2253 GNDA.t96 GNDA.n169 172.876
R2254 GNDA.t96 GNDA.n170 172.615
R2255 GNDA.t109 GNDA.n584 323.404
R2256 GNDA.t109 GNDA.n1598 323.404
R2257 GNDA.n1268 GNDA.t101 172.615
R2258 GNDA.n685 GNDA.t101 172.615
R2259 GNDA.t96 GNDA.n115 172.615
R2260 GNDA.n1716 GNDA.n1715 323.2
R2261 GNDA.n1695 GNDA.n1694 322.861
R2262 GNDA.n355 GNDA.n333 321.281
R2263 GNDA.n2463 GNDA.n2462 321.281
R2264 GNDA.n487 GNDA.n319 320
R2265 GNDA.n2454 GNDA.n2453 320
R2266 GNDA.n335 GNDA.n333 318.08
R2267 GNDA.n2462 GNDA.n2461 318.08
R2268 GNDA.n1717 GNDA.n1716 316.8
R2269 GNDA.n473 GNDA.n360 310.401
R2270 GNDA.n43 GNDA.n38 310.401
R2271 GNDA.n467 GNDA.n324 307.2
R2272 GNDA.n2433 GNDA.n2432 304
R2273 GNDA.n479 GNDA.n331 304
R2274 GNDA.n45 GNDA.n39 304
R2275 GNDA.n2410 GNDA.n117 301.474
R2276 GNDA.n2432 GNDA.n97 300.8
R2277 GNDA.n2433 GNDA.n96 300.8
R2278 GNDA.n356 GNDA.n332 300.8
R2279 GNDA.n436 GNDA.n374 300.8
R2280 GNDA.n433 GNDA.n374 300.8
R2281 GNDA.n61 GNDA.n60 300.8
R2282 GNDA.n2155 GNDA.n508 297.601
R2283 GNDA.n2155 GNDA.n2154 297.601
R2284 GNDA.n97 GNDA.n96 297.601
R2285 GNDA.n2153 GNDA.n511 297.601
R2286 GNDA.n514 GNDA.n511 297.601
R2287 GNDA.n349 GNDA.n348 296
R2288 GNDA.n2456 GNDA.n67 296
R2289 GNDA.n1726 GNDA.n1725 294.401
R2290 GNDA.n1725 GNDA.n1724 294.401
R2291 GNDA.n1715 GNDA.n1629 294.401
R2292 GNDA.n2461 GNDA.n2460 292.5
R2293 GNDA.n2460 GNDA.n2459 292.5
R2294 GNDA.n2462 GNDA.n59 292.5
R2295 GNDA.n64 GNDA.n59 292.5
R2296 GNDA.n61 GNDA.n58 292.5
R2297 GNDA.n64 GNDA.n58 292.5
R2298 GNDA.n2453 GNDA.n2452 292.5
R2299 GNDA.n2452 GNDA.n2451 292.5
R2300 GNDA.n74 GNDA.n70 292.5
R2301 GNDA.n75 GNDA.n74 292.5
R2302 GNDA.n73 GNDA.n72 292.5
R2303 GNDA.n73 GNDA.n62 292.5
R2304 GNDA.n71 GNDA.n69 292.5
R2305 GNDA.n75 GNDA.n71 292.5
R2306 GNDA.n2457 GNDA.n2456 292.5
R2307 GNDA.n2458 GNDA.n2457 292.5
R2308 GNDA.n424 GNDA.n375 292.5
R2309 GNDA.n425 GNDA.n424 292.5
R2310 GNDA.n423 GNDA.n383 292.5
R2311 GNDA.n423 GNDA.n422 292.5
R2312 GNDA.n446 GNDA.n445 292.5
R2313 GNDA.n445 GNDA.n57 292.5
R2314 GNDA.n447 GNDA.n442 292.5
R2315 GNDA.n442 GNDA.n441 292.5
R2316 GNDA.n436 GNDA.n431 292.5
R2317 GNDA.n431 GNDA.n29 292.5
R2318 GNDA.n378 GNDA.n374 292.5
R2319 GNDA.n440 GNDA.n378 292.5
R2320 GNDA.n433 GNDA.n430 292.5
R2321 GNDA.n430 GNDA.n429 292.5
R2322 GNDA.n439 GNDA.n438 292.5
R2323 GNDA.n440 GNDA.n439 292.5
R2324 GNDA.n2488 GNDA.n2487 292.5
R2325 GNDA.n2487 GNDA.n2486 292.5
R2326 GNDA.n28 GNDA.n25 292.5
R2327 GNDA.n440 GNDA.n28 292.5
R2328 GNDA.n427 GNDA.n426 292.5
R2329 GNDA.n428 GNDA.n427 292.5
R2330 GNDA.n27 GNDA.n26 292.5
R2331 GNDA.n440 GNDA.n27 292.5
R2332 GNDA.n2484 GNDA.n2483 292.5
R2333 GNDA.n2485 GNDA.n2484 292.5
R2334 GNDA.n34 GNDA.n32 292.5
R2335 GNDA.n440 GNDA.n32 292.5
R2336 GNDA.n417 GNDA.n391 292.5
R2337 GNDA.n391 GNDA.n390 292.5
R2338 GNDA.n420 GNDA.n419 292.5
R2339 GNDA.n421 GNDA.n420 292.5
R2340 GNDA.n392 GNDA.n388 292.5
R2341 GNDA.n390 GNDA.n388 292.5
R2342 GNDA.n33 GNDA.n31 292.5
R2343 GNDA.n440 GNDA.n31 292.5
R2344 GNDA.n473 GNDA.n472 292.5
R2345 GNDA.n472 GNDA.n471 292.5
R2346 GNDA.n478 GNDA.n329 292.5
R2347 GNDA.n361 GNDA.n329 292.5
R2348 GNDA.n480 GNDA.n479 292.5
R2349 GNDA.n481 GNDA.n480 292.5
R2350 GNDA.n359 GNDA.n328 292.5
R2351 GNDA.n361 GNDA.n328 292.5
R2352 GNDA.n2464 GNDA.n2463 292.5
R2353 GNDA.n2465 GNDA.n2464 292.5
R2354 GNDA.n41 GNDA.n39 292.5
R2355 GNDA.n55 GNDA.n41 292.5
R2356 GNDA.n2475 GNDA.n2474 292.5
R2357 GNDA.n2474 GNDA.n2473 292.5
R2358 GNDA.n40 GNDA.n38 292.5
R2359 GNDA.n457 GNDA.n40 292.5
R2360 GNDA.n2472 GNDA.n2471 292.5
R2361 GNDA.n2473 GNDA.n2472 292.5
R2362 GNDA.n460 GNDA.n459 292.5
R2363 GNDA.n459 GNDA.n458 292.5
R2364 GNDA.n461 GNDA.n364 292.5
R2365 GNDA.n440 GNDA.n364 292.5
R2366 GNDA.n469 GNDA.n468 292.5
R2367 GNDA.n470 GNDA.n469 292.5
R2368 GNDA.n450 GNDA.n363 292.5
R2369 GNDA.n440 GNDA.n363 292.5
R2370 GNDA.n466 GNDA.n465 292.5
R2371 GNDA.n465 GNDA.n362 292.5
R2372 GNDA.n326 GNDA.n324 292.5
R2373 GNDA.t74 GNDA.n326 292.5
R2374 GNDA.n484 GNDA.n483 292.5
R2375 GNDA.n483 GNDA.n482 292.5
R2376 GNDA.n463 GNDA.n325 292.5
R2377 GNDA.t74 GNDA.n325 292.5
R2378 GNDA.n2468 GNDA.n2467 292.5
R2379 GNDA.n2467 GNDA.n2466 292.5
R2380 GNDA.n2469 GNDA.n47 292.5
R2381 GNDA.t279 GNDA.n47 292.5
R2382 GNDA.n455 GNDA.n46 292.5
R2383 GNDA.n456 GNDA.n455 292.5
R2384 GNDA.n54 GNDA.n53 292.5
R2385 GNDA.t279 GNDA.n54 292.5
R2386 GNDA.n355 GNDA.n354 292.5
R2387 GNDA.n354 GNDA.n327 292.5
R2388 GNDA.n353 GNDA.n333 292.5
R2389 GNDA.n353 GNDA.n352 292.5
R2390 GNDA.n336 GNDA.n335 292.5
R2391 GNDA.n345 GNDA.n336 292.5
R2392 GNDA.n334 GNDA.n332 292.5
R2393 GNDA.n352 GNDA.n334 292.5
R2394 GNDA.n320 GNDA.n317 292.5
R2395 GNDA.n342 GNDA.n317 292.5
R2396 GNDA.n343 GNDA.n321 292.5
R2397 GNDA.n344 GNDA.n343 292.5
R2398 GNDA.n486 GNDA.n318 292.5
R2399 GNDA.n342 GNDA.n318 292.5
R2400 GNDA.n488 GNDA.n487 292.5
R2401 GNDA.n489 GNDA.n488 292.5
R2402 GNDA.n348 GNDA.n347 292.5
R2403 GNDA.n347 GNDA.n346 292.5
R2404 GNDA.n2181 GNDA.n2180 292.5
R2405 GNDA.n2182 GNDA.n2181 292.5
R2406 GNDA.n2179 GNDA.n313 292.5
R2407 GNDA.n2150 GNDA.n313 292.5
R2408 GNDA.n2178 GNDA.n2177 292.5
R2409 GNDA.n2177 GNDA.n2176 292.5
R2410 GNDA.n314 GNDA.n312 292.5
R2411 GNDA.n2150 GNDA.n312 292.5
R2412 GNDA.n2171 GNDA.n2170 292.5
R2413 GNDA.n2170 GNDA.n2169 292.5
R2414 GNDA.n2173 GNDA.n492 292.5
R2415 GNDA.n2151 GNDA.n492 292.5
R2416 GNDA.n2175 GNDA.n2174 292.5
R2417 GNDA.n2176 GNDA.n2175 292.5
R2418 GNDA.n493 GNDA.n491 292.5
R2419 GNDA.n2151 GNDA.n491 292.5
R2420 GNDA.n102 GNDA.n99 292.5
R2421 GNDA.n102 GNDA.n101 292.5
R2422 GNDA.n106 GNDA.n105 292.5
R2423 GNDA.n2429 GNDA.n106 292.5
R2424 GNDA.n104 GNDA.n100 292.5
R2425 GNDA.n307 GNDA.n100 292.5
R2426 GNDA.n2431 GNDA.n2430 292.5
R2427 GNDA.n2430 GNDA.n2429 292.5
R2428 GNDA.n511 GNDA.n505 292.5
R2429 GNDA.n2157 GNDA.n505 292.5
R2430 GNDA.n515 GNDA.n514 292.5
R2431 GNDA.n2151 GNDA.n515 292.5
R2432 GNDA.n512 GNDA.n510 292.5
R2433 GNDA.n2124 GNDA.n512 292.5
R2434 GNDA.n2153 GNDA.n2152 292.5
R2435 GNDA.n2152 GNDA.n2151 292.5
R2436 GNDA.n2434 GNDA.n2433 292.5
R2437 GNDA.n2435 GNDA.n2434 292.5
R2438 GNDA.n2432 GNDA.n95 292.5
R2439 GNDA.n2429 GNDA.n95 292.5
R2440 GNDA.n166 GNDA.n97 292.5
R2441 GNDA.n167 GNDA.n166 292.5
R2442 GNDA.n96 GNDA.n94 292.5
R2443 GNDA.n2429 GNDA.n94 292.5
R2444 GNDA.n2156 GNDA.n2155 292.5
R2445 GNDA.n2157 GNDA.n2156 292.5
R2446 GNDA.n2154 GNDA.n507 292.5
R2447 GNDA.n2151 GNDA.n507 292.5
R2448 GNDA.n2123 GNDA.n509 292.5
R2449 GNDA.n2124 GNDA.n2123 292.5
R2450 GNDA.n508 GNDA.n506 292.5
R2451 GNDA.n2151 GNDA.n506 292.5
R2452 GNDA.n1718 GNDA.n1717 292.5
R2453 GNDA.n1719 GNDA.n1718 292.5
R2454 GNDA.n1716 GNDA.n1628 292.5
R2455 GNDA.n1705 GNDA.n1628 292.5
R2456 GNDA.n1715 GNDA.n1714 292.5
R2457 GNDA.n1714 GNDA.n1713 292.5
R2458 GNDA.n1629 GNDA.n1627 292.5
R2459 GNDA.n1705 GNDA.n1627 292.5
R2460 GNDA.n1693 GNDA.n1692 292.5
R2461 GNDA.n1696 GNDA.n1695 292.5
R2462 GNDA.n1642 GNDA.n1630 292.5
R2463 GNDA.n1644 GNDA.n1642 292.5
R2464 GNDA.n1638 GNDA.n1636 292.5
R2465 GNDA.n1685 GNDA.n1638 292.5
R2466 GNDA.n1640 GNDA.n1639 292.5
R2467 GNDA.n1696 GNDA.n1640 292.5
R2468 GNDA.n1637 GNDA.n1635 292.5
R2469 GNDA.n1643 GNDA.n1637 292.5
R2470 GNDA.n1698 GNDA.n1697 292.5
R2471 GNDA.n1697 GNDA.n1696 292.5
R2472 GNDA.n1690 GNDA.n1689 292.5
R2473 GNDA.n1691 GNDA.n1690 292.5
R2474 GNDA.n1631 GNDA.n1615 292.5
R2475 GNDA.n1730 GNDA.n1615 292.5
R2476 GNDA.n1687 GNDA.n1686 292.5
R2477 GNDA.n1686 GNDA.n1609 292.5
R2478 GNDA.n1688 GNDA.n1616 292.5
R2479 GNDA.n1730 GNDA.n1616 292.5
R2480 GNDA.n1723 GNDA.n1722 292.5
R2481 GNDA.n1722 GNDA.n1721 292.5
R2482 GNDA.n1706 GNDA.n1625 292.5
R2483 GNDA.n1707 GNDA.n1706 292.5
R2484 GNDA.n1711 GNDA.n1710 292.5
R2485 GNDA.n1712 GNDA.n1711 292.5
R2486 GNDA.n1726 GNDA.n1618 292.5
R2487 GNDA.n1645 GNDA.n1618 292.5
R2488 GNDA.n1725 GNDA.n1614 292.5
R2489 GNDA.n1730 GNDA.n1614 292.5
R2490 GNDA.n1724 GNDA.n1617 292.5
R2491 GNDA.n1720 GNDA.n1617 292.5
R2492 GNDA.n1729 GNDA.n1728 292.5
R2493 GNDA.n1730 GNDA.n1729 292.5
R2494 GNDA.n1678 GNDA.n1677 292.5
R2495 GNDA.n1679 GNDA.n1678 292.5
R2496 GNDA.n1676 GNDA.n1675 292.5
R2497 GNDA.n1675 GNDA.n1641 292.5
R2498 GNDA.n1647 GNDA.n1622 292.5
R2499 GNDA.n1647 GNDA.n1646 292.5
R2500 GNDA.n1733 GNDA.n1732 292.5
R2501 GNDA.n1732 GNDA.n1731 292.5
R2502 GNDA.n1734 GNDA.n1611 292.5
R2503 GNDA.n1705 GNDA.n1611 292.5
R2504 GNDA.n1736 GNDA.n1735 292.5
R2505 GNDA.n1737 GNDA.n1736 292.5
R2506 GNDA.n1612 GNDA.n1610 292.5
R2507 GNDA.n1705 GNDA.n1610 292.5
R2508 GNDA.n509 GNDA.n508 291.2
R2509 GNDA.n2154 GNDA.n509 291.2
R2510 GNDA.n2153 GNDA.n510 291.2
R2511 GNDA.n514 GNDA.n510 291.2
R2512 GNDA.n1717 GNDA.n1629 288
R2513 GNDA.n1652 GNDA.n1651 281.601
R2514 GNDA.n1709 GNDA.n1624 281.601
R2515 GNDA.n1677 GNDA.n1676 278.401
R2516 GNDA.n1710 GNDA.n1625 278.401
R2517 GNDA.n886 GNDA.t109 267.529
R2518 GNDA.t109 GNDA.n1435 267.529
R2519 GNDA.n1862 GNDA.t109 267.529
R2520 GNDA.n1691 GNDA.n1685 265.517
R2521 GNDA.n2287 GNDA.n281 259.416
R2522 GNDA.n2333 GNDA.n145 259.416
R2523 GNDA.n2059 GNDA.n567 259.416
R2524 GNDA.n1388 GNDA.n654 259.416
R2525 GNDA.n1848 GNDA.n603 259.416
R2526 GNDA.n1450 GNDA.n1415 259.416
R2527 GNDA.n874 GNDA.n873 259.416
R2528 GNDA.n957 GNDA.n956 259.416
R2529 GNDA.n1197 GNDA.n1076 259.416
R2530 GNDA.n435 GNDA.t122 258.601
R2531 GNDA.n432 GNDA.t125 258.601
R2532 GNDA.n1851 GNDA.n1850 254.494
R2533 GNDA.n875 GNDA.n747 254.392
R2534 GNDA.n1448 GNDA.n1447 254.392
R2535 GNDA.n1873 GNDA.n584 254.34
R2536 GNDA.n1879 GNDA.n584 254.34
R2537 GNDA.n1881 GNDA.n584 254.34
R2538 GNDA.n1887 GNDA.n584 254.34
R2539 GNDA.n1889 GNDA.n584 254.34
R2540 GNDA.n1895 GNDA.n584 254.34
R2541 GNDA.n1598 GNDA.n1597 254.34
R2542 GNDA.n1598 GNDA.n624 254.34
R2543 GNDA.n1598 GNDA.n623 254.34
R2544 GNDA.n1598 GNDA.n622 254.34
R2545 GNDA.n1598 GNDA.n621 254.34
R2546 GNDA.n1598 GNDA.n620 254.34
R2547 GNDA.n713 GNDA.n564 254.34
R2548 GNDA.n943 GNDA.n564 254.34
R2549 GNDA.n939 GNDA.n564 254.34
R2550 GNDA.n929 GNDA.n564 254.34
R2551 GNDA.n927 GNDA.n564 254.34
R2552 GNDA.n648 GNDA.n564 254.34
R2553 GNDA.n645 GNDA.n564 254.34
R2554 GNDA.n640 GNDA.n564 254.34
R2555 GNDA.n637 GNDA.n564 254.34
R2556 GNDA.n632 GNDA.n564 254.34
R2557 GNDA.n1930 GNDA.n1929 254.34
R2558 GNDA.n1928 GNDA.n564 254.34
R2559 GNDA.n1916 GNDA.n564 254.34
R2560 GNDA.n1915 GNDA.n564 254.34
R2561 GNDA.n576 GNDA.n564 254.34
R2562 GNDA.n1903 GNDA.n564 254.34
R2563 GNDA.n923 GNDA.n563 254.34
R2564 GNDA.n933 GNDA.n563 254.34
R2565 GNDA.n935 GNDA.n563 254.34
R2566 GNDA.n947 GNDA.n563 254.34
R2567 GNDA.n950 GNDA.n563 254.34
R2568 GNDA.n630 GNDA.n563 254.34
R2569 GNDA.n1567 GNDA.n563 254.34
R2570 GNDA.n1561 GNDA.n563 254.34
R2571 GNDA.n1559 GNDA.n563 254.34
R2572 GNDA.n1553 GNDA.n563 254.34
R2573 GNDA.n1898 GNDA.n563 254.34
R2574 GNDA.n1908 GNDA.n563 254.34
R2575 GNDA.n1910 GNDA.n563 254.34
R2576 GNDA.n1921 GNDA.n563 254.34
R2577 GNDA.n1924 GNDA.n563 254.34
R2578 GNDA.n1813 GNDA.n1812 254.34
R2579 GNDA.n1268 GNDA.n1267 254.34
R2580 GNDA.n1268 GNDA.n1213 254.34
R2581 GNDA.n1268 GNDA.n1212 254.34
R2582 GNDA.n1268 GNDA.n1211 254.34
R2583 GNDA.n1268 GNDA.n1210 254.34
R2584 GNDA.n1268 GNDA.n1209 254.34
R2585 GNDA.n685 GNDA.n684 254.34
R2586 GNDA.n685 GNDA.n659 254.34
R2587 GNDA.n685 GNDA.n658 254.34
R2588 GNDA.n685 GNDA.n657 254.34
R2589 GNDA.n685 GNDA.n656 254.34
R2590 GNDA.n685 GNDA.n655 254.34
R2591 GNDA.n2330 GNDA.n2329 254.34
R2592 GNDA.n2328 GNDA.n2327 254.34
R2593 GNDA.n2327 GNDA.n164 254.34
R2594 GNDA.n2327 GNDA.n163 254.34
R2595 GNDA.n2327 GNDA.n162 254.34
R2596 GNDA.n2327 GNDA.n161 254.34
R2597 GNDA.n2296 GNDA.n203 254.34
R2598 GNDA.n2296 GNDA.n202 254.34
R2599 GNDA.n2296 GNDA.n201 254.34
R2600 GNDA.n2296 GNDA.n200 254.34
R2601 GNDA.n2296 GNDA.n199 254.34
R2602 GNDA.n2022 GNDA.n2021 254.34
R2603 GNDA.n2327 GNDA.n159 254.34
R2604 GNDA.n2327 GNDA.n158 254.34
R2605 GNDA.n2327 GNDA.n157 254.34
R2606 GNDA.n2327 GNDA.n156 254.34
R2607 GNDA.n2327 GNDA.n155 254.34
R2608 GNDA.n2296 GNDA.n197 254.34
R2609 GNDA.n2296 GNDA.n196 254.34
R2610 GNDA.n2296 GNDA.n195 254.34
R2611 GNDA.n2296 GNDA.n194 254.34
R2612 GNDA.n2296 GNDA.n193 254.34
R2613 GNDA.n2327 GNDA.n154 254.34
R2614 GNDA.n1100 GNDA.n165 254.34
R2615 GNDA.n1174 GNDA.n165 254.34
R2616 GNDA.n1094 GNDA.n165 254.34
R2617 GNDA.n1185 GNDA.n165 254.34
R2618 GNDA.n1085 GNDA.n165 254.34
R2619 GNDA.n1196 GNDA.n165 254.34
R2620 GNDA.n955 GNDA.n712 254.34
R2621 GNDA.n1208 GNDA.n1207 254.34
R2622 GNDA.n1208 GNDA.n690 254.34
R2623 GNDA.n1208 GNDA.n689 254.34
R2624 GNDA.n1208 GNDA.n688 254.34
R2625 GNDA.n1208 GNDA.n687 254.34
R2626 GNDA.n1208 GNDA.n686 254.34
R2627 GNDA.n1203 GNDA.n1050 254.34
R2628 GNDA.n772 GNDA.n618 254.34
R2629 GNDA.n850 GNDA.n618 254.34
R2630 GNDA.n766 GNDA.n618 254.34
R2631 GNDA.n861 GNDA.n618 254.34
R2632 GNDA.n757 GNDA.n618 254.34
R2633 GNDA.n872 GNDA.n618 254.34
R2634 GNDA.n774 GNDA.n773 254.34
R2635 GNDA.n2327 GNDA.n153 254.34
R2636 GNDA.n2327 GNDA.n152 254.34
R2637 GNDA.n2327 GNDA.n151 254.34
R2638 GNDA.n2327 GNDA.n150 254.34
R2639 GNDA.n2327 GNDA.n149 254.34
R2640 GNDA.n2297 GNDA.n2296 254.34
R2641 GNDA.n2296 GNDA.n191 254.34
R2642 GNDA.n2296 GNDA.n190 254.34
R2643 GNDA.n2296 GNDA.n189 254.34
R2644 GNDA.n2296 GNDA.n188 254.34
R2645 GNDA.n2301 GNDA.n170 254.34
R2646 GNDA.n2307 GNDA.n170 254.34
R2647 GNDA.n2309 GNDA.n170 254.34
R2648 GNDA.n2315 GNDA.n170 254.34
R2649 GNDA.n2317 GNDA.n170 254.34
R2650 GNDA.n2323 GNDA.n170 254.34
R2651 GNDA.n2327 GNDA.n148 254.34
R2652 GNDA.n1390 GNDA.n652 254.34
R2653 GNDA.n1291 GNDA.n1269 254.34
R2654 GNDA.n1365 GNDA.n1269 254.34
R2655 GNDA.n1286 GNDA.n1269 254.34
R2656 GNDA.n1376 GNDA.n1269 254.34
R2657 GNDA.n1277 GNDA.n1269 254.34
R2658 GNDA.n1387 GNDA.n1269 254.34
R2659 GNDA.n2294 GNDA.n2293 254.34
R2660 GNDA.n1546 GNDA.n617 254.34
R2661 GNDA.n1462 GNDA.n617 254.34
R2662 GNDA.n1474 GNDA.n617 254.34
R2663 GNDA.n1460 GNDA.n617 254.34
R2664 GNDA.n1485 GNDA.n617 254.34
R2665 GNDA.n1451 GNDA.n617 254.34
R2666 GNDA.n1551 GNDA.n1550 254.34
R2667 GNDA.n305 GNDA.n169 254.34
R2668 GNDA.n2264 GNDA.n169 254.34
R2669 GNDA.n299 GNDA.n169 254.34
R2670 GNDA.n2275 GNDA.n169 254.34
R2671 GNDA.n290 GNDA.n169 254.34
R2672 GNDA.n2286 GNDA.n169 254.34
R2673 GNDA.n253 GNDA.n115 254.34
R2674 GNDA.n209 GNDA.n115 254.34
R2675 GNDA.n246 GNDA.n115 254.34
R2676 GNDA.n240 GNDA.n115 254.34
R2677 GNDA.n238 GNDA.n115 254.34
R2678 GNDA.n232 GNDA.n115 254.34
R2679 GNDA.n2147 GNDA.n2146 254.34
R2680 GNDA.n309 GNDA.n306 254.34
R2681 GNDA.n109 GNDA.n90 254.34
R2682 GNDA.n1737 GNDA.n1609 252.875
R2683 GNDA.n2079 GNDA.n548 250.349
R2684 GNDA.n2302 GNDA.n2300 249.663
R2685 GNDA.n254 GNDA.n160 249.663
R2686 GNDA.n1901 GNDA.n580 249.663
R2687 GNDA.n683 GNDA.n631 249.663
R2688 GNDA.n1874 GNDA.n1872 249.663
R2689 GNDA.n1596 GNDA.n626 249.663
R2690 GNDA.n896 GNDA.n735 249.663
R2691 GNDA.n926 GNDA.n561 249.663
R2692 GNDA.n2096 GNDA.n2095 249.663
R2693 GNDA.n2444 GNDA.n2443 248.049
R2694 GNDA.n486 GNDA.n485 246.4
R2695 GNDA.n70 GNDA.n50 246.4
R2696 GNDA.t109 GNDA.n885 244.762
R2697 GNDA.n1436 GNDA.t109 244.762
R2698 GNDA.t109 GNDA.n1861 244.762
R2699 GNDA.n2445 GNDA.n82 241.291
R2700 GNDA.n1676 GNDA.n1622 240
R2701 GNDA.n1723 GNDA.n1625 240
R2702 GNDA.n1834 GNDA.t109 239.004
R2703 GNDA.n1821 GNDA.n1738 239.004
R2704 GNDA.n2046 GNDA.t101 239.004
R2705 GNDA.t96 GNDA.n118 239.004
R2706 GNDA.n339 GNDA.n338 238.4
R2707 GNDA.n2455 GNDA.n68 238.4
R2708 GNDA.t245 GNDA.t124 236.923
R2709 GNDA.t239 GNDA.t308 236.923
R2710 GNDA.t244 GNDA.t303 236.923
R2711 GNDA.t87 GNDA.t307 236.923
R2712 GNDA.t301 GNDA.t150 236.923
R2713 GNDA.t304 GNDA.t336 236.923
R2714 GNDA.t204 GNDA.t299 236.923
R2715 GNDA.t37 GNDA.t121 236.923
R2716 GNDA.n419 GNDA.n392 233.601
R2717 GNDA.n357 GNDA.t135 224.525
R2718 GNDA.n330 GNDA.t145 224.525
R2719 GNDA.n44 GNDA.t172 224.525
R2720 GNDA.n42 GNDA.t91 224.525
R2721 GNDA.n1527 GNDA.n1402 221.667
R2722 GNDA.n1344 GNDA.n1343 221.667
R2723 GNDA.n2243 GNDA.n2242 221.667
R2724 GNDA.n829 GNDA.n828 221.667
R2725 GNDA.n1029 GNDA.n1028 221.667
R2726 GNDA.n1153 GNDA.n1152 221.667
R2727 GNDA.n1796 GNDA.n1750 221.667
R2728 GNDA.n2005 GNDA.n1961 221.667
R2729 GNDA.n2388 GNDA.n2387 221.667
R2730 GNDA.n2488 GNDA.n26 217.601
R2731 GNDA.n426 GNDA.n26 214.4
R2732 GNDA.n438 GNDA.n434 211.201
R2733 GNDA.n438 GNDA.n437 211.201
R2734 GNDA.n463 GNDA.n323 211.201
R2735 GNDA.n464 GNDA.n463 211.201
R2736 GNDA.n53 GNDA.n52 211.201
R2737 GNDA.n53 GNDA.n49 211.201
R2738 GNDA.n15 GNDA.n13 206.052
R2739 GNDA.n4 GNDA.n2 206.052
R2740 GNDA.n23 GNDA.n22 205.488
R2741 GNDA.n21 GNDA.n20 205.488
R2742 GNDA.n19 GNDA.n18 205.488
R2743 GNDA.n17 GNDA.n16 205.488
R2744 GNDA.n15 GNDA.n14 205.488
R2745 GNDA.n12 GNDA.n11 205.488
R2746 GNDA.n10 GNDA.n9 205.488
R2747 GNDA.n8 GNDA.n7 205.488
R2748 GNDA.n6 GNDA.n5 205.488
R2749 GNDA.n4 GNDA.n3 205.488
R2750 GNDA.n426 GNDA.n25 203.201
R2751 GNDA.n2489 GNDA.n2488 201.601
R2752 GNDA.n2436 GNDA.n2435 200.225
R2753 GNDA.n2190 GNDA.n2189 197
R2754 GNDA.n2437 GNDA.n91 197
R2755 GNDA.n2024 GNDA.n204 197
R2756 GNDA.n2295 GNDA.n206 197
R2757 GNDA.n1815 GNDA.n1814 197
R2758 GNDA.n1548 GNDA.n1392 197
R2759 GNDA.n776 GNDA.n775 197
R2760 GNDA.n692 GNDA.n205 197
R2761 GNDA.n2078 GNDA.n549 197
R2762 GNDA.n1099 GNDA.n518 197
R2763 GNDA.n76 GNDA.n68 195
R2764 GNDA.n77 GNDA.n76 195
R2765 GNDA.n67 GNDA.n66 195
R2766 GNDA.n66 GNDA.n65 195
R2767 GNDA.n350 GNDA.n349 195
R2768 GNDA.n351 GNDA.n350 195
R2769 GNDA.n340 GNDA.n338 195
R2770 GNDA.n341 GNDA.n340 195
R2771 GNDA.n360 GNDA.n359 192
R2772 GNDA.n2471 GNDA.n43 192
R2773 GNDA.n2325 GNDA.n174 187.249
R2774 GNDA.n231 GNDA.n230 187.249
R2775 GNDA.n1245 GNDA.n1244 187.249
R2776 GNDA.n2298 GNDA.n184 187.249
R2777 GNDA.n1899 GNDA.n1897 187.249
R2778 GNDA.n1573 GNDA.n1572 187.249
R2779 GNDA.n924 GNDA.n922 187.249
R2780 GNDA.n2093 GNDA.n2092 187.249
R2781 GNDA.n2126 GNDA.n2121 187.249
R2782 GNDA.n440 GNDA.t305 186.155
R2783 GNDA.n440 GNDA.t300 186.155
R2784 GNDA.n1492 GNDA.n1491 185
R2785 GNDA.n1493 GNDA.n1410 185
R2786 GNDA.n1410 GNDA.t108 185
R2787 GNDA.n1495 GNDA.n1494 185
R2788 GNDA.n1497 GNDA.n1409 185
R2789 GNDA.n1500 GNDA.n1499 185
R2790 GNDA.n1501 GNDA.n1408 185
R2791 GNDA.n1503 GNDA.n1502 185
R2792 GNDA.n1505 GNDA.n1407 185
R2793 GNDA.n1508 GNDA.n1507 185
R2794 GNDA.n1509 GNDA.n1406 185
R2795 GNDA.n1511 GNDA.n1510 185
R2796 GNDA.n1513 GNDA.n1405 185
R2797 GNDA.n1516 GNDA.n1515 185
R2798 GNDA.n1517 GNDA.n1404 185
R2799 GNDA.n1519 GNDA.n1518 185
R2800 GNDA.n1521 GNDA.n1403 185
R2801 GNDA.n1524 GNDA.n1523 185
R2802 GNDA.n1525 GNDA.n1402 185
R2803 GNDA.n1542 GNDA.n1541 185
R2804 GNDA.n1539 GNDA.n1396 185
R2805 GNDA.n1538 GNDA.n1398 185
R2806 GNDA.n1536 GNDA.n1535 185
R2807 GNDA.n1534 GNDA.n1399 185
R2808 GNDA.n1533 GNDA.n1532 185
R2809 GNDA.n1530 GNDA.n1400 185
R2810 GNDA.n1530 GNDA.t108 185
R2811 GNDA.n1529 GNDA.n1401 185
R2812 GNDA.n1527 GNDA.n1526 185
R2813 GNDA.n1310 GNDA.n1309 185
R2814 GNDA.n1311 GNDA.n1308 185
R2815 GNDA.n1311 GNDA.t100 185
R2816 GNDA.n1314 GNDA.n1313 185
R2817 GNDA.n1315 GNDA.n1307 185
R2818 GNDA.n1317 GNDA.n1316 185
R2819 GNDA.n1319 GNDA.n1306 185
R2820 GNDA.n1322 GNDA.n1321 185
R2821 GNDA.n1323 GNDA.n1305 185
R2822 GNDA.n1325 GNDA.n1324 185
R2823 GNDA.n1327 GNDA.n1304 185
R2824 GNDA.n1330 GNDA.n1329 185
R2825 GNDA.n1331 GNDA.n1303 185
R2826 GNDA.n1333 GNDA.n1332 185
R2827 GNDA.n1335 GNDA.n1302 185
R2828 GNDA.n1338 GNDA.n1337 185
R2829 GNDA.n1339 GNDA.n1301 185
R2830 GNDA.n1341 GNDA.n1340 185
R2831 GNDA.n1343 GNDA.n1300 185
R2832 GNDA.n1360 GNDA.n1295 185
R2833 GNDA.n1358 GNDA.n1357 185
R2834 GNDA.n1356 GNDA.n1296 185
R2835 GNDA.n1355 GNDA.n1354 185
R2836 GNDA.n1352 GNDA.n1297 185
R2837 GNDA.n1350 GNDA.n1349 185
R2838 GNDA.n1348 GNDA.n1298 185
R2839 GNDA.n1298 GNDA.t100 185
R2840 GNDA.n1347 GNDA.n1346 185
R2841 GNDA.n1344 GNDA.n1299 185
R2842 GNDA.n2209 GNDA.n2208 185
R2843 GNDA.n2210 GNDA.n2207 185
R2844 GNDA.n2210 GNDA.t173 185
R2845 GNDA.n2213 GNDA.n2212 185
R2846 GNDA.n2214 GNDA.n2206 185
R2847 GNDA.n2216 GNDA.n2215 185
R2848 GNDA.n2218 GNDA.n2205 185
R2849 GNDA.n2221 GNDA.n2220 185
R2850 GNDA.n2222 GNDA.n2204 185
R2851 GNDA.n2224 GNDA.n2223 185
R2852 GNDA.n2226 GNDA.n2203 185
R2853 GNDA.n2229 GNDA.n2228 185
R2854 GNDA.n2230 GNDA.n2202 185
R2855 GNDA.n2232 GNDA.n2231 185
R2856 GNDA.n2234 GNDA.n2201 185
R2857 GNDA.n2237 GNDA.n2236 185
R2858 GNDA.n2238 GNDA.n2200 185
R2859 GNDA.n2240 GNDA.n2239 185
R2860 GNDA.n2242 GNDA.n2199 185
R2861 GNDA.n2259 GNDA.n2194 185
R2862 GNDA.n2257 GNDA.n2256 185
R2863 GNDA.n2255 GNDA.n2195 185
R2864 GNDA.n2254 GNDA.n2253 185
R2865 GNDA.n2251 GNDA.n2196 185
R2866 GNDA.n2249 GNDA.n2248 185
R2867 GNDA.n2247 GNDA.n2197 185
R2868 GNDA.n2197 GNDA.t173 185
R2869 GNDA.n2246 GNDA.n2245 185
R2870 GNDA.n2243 GNDA.n2198 185
R2871 GNDA.n795 GNDA.n794 185
R2872 GNDA.n796 GNDA.n793 185
R2873 GNDA.n796 GNDA.t126 185
R2874 GNDA.n799 GNDA.n798 185
R2875 GNDA.n800 GNDA.n792 185
R2876 GNDA.n802 GNDA.n801 185
R2877 GNDA.n804 GNDA.n791 185
R2878 GNDA.n807 GNDA.n806 185
R2879 GNDA.n808 GNDA.n790 185
R2880 GNDA.n810 GNDA.n809 185
R2881 GNDA.n812 GNDA.n789 185
R2882 GNDA.n815 GNDA.n814 185
R2883 GNDA.n816 GNDA.n788 185
R2884 GNDA.n818 GNDA.n817 185
R2885 GNDA.n820 GNDA.n787 185
R2886 GNDA.n823 GNDA.n822 185
R2887 GNDA.n824 GNDA.n786 185
R2888 GNDA.n826 GNDA.n825 185
R2889 GNDA.n828 GNDA.n785 185
R2890 GNDA.n845 GNDA.n780 185
R2891 GNDA.n843 GNDA.n842 185
R2892 GNDA.n841 GNDA.n781 185
R2893 GNDA.n840 GNDA.n839 185
R2894 GNDA.n837 GNDA.n782 185
R2895 GNDA.n835 GNDA.n834 185
R2896 GNDA.n833 GNDA.n783 185
R2897 GNDA.n783 GNDA.t126 185
R2898 GNDA.n832 GNDA.n831 185
R2899 GNDA.n829 GNDA.n784 185
R2900 GNDA.n995 GNDA.n710 185
R2901 GNDA.n996 GNDA.n709 185
R2902 GNDA.n996 GNDA.t139 185
R2903 GNDA.n999 GNDA.n998 185
R2904 GNDA.n1000 GNDA.n708 185
R2905 GNDA.n1002 GNDA.n1001 185
R2906 GNDA.n1004 GNDA.n707 185
R2907 GNDA.n1007 GNDA.n1006 185
R2908 GNDA.n1008 GNDA.n706 185
R2909 GNDA.n1010 GNDA.n1009 185
R2910 GNDA.n1012 GNDA.n705 185
R2911 GNDA.n1015 GNDA.n1014 185
R2912 GNDA.n1016 GNDA.n704 185
R2913 GNDA.n1018 GNDA.n1017 185
R2914 GNDA.n1020 GNDA.n703 185
R2915 GNDA.n1023 GNDA.n1022 185
R2916 GNDA.n1024 GNDA.n702 185
R2917 GNDA.n1026 GNDA.n1025 185
R2918 GNDA.n1028 GNDA.n701 185
R2919 GNDA.n1045 GNDA.n693 185
R2920 GNDA.n1043 GNDA.n1042 185
R2921 GNDA.n1041 GNDA.n697 185
R2922 GNDA.n1040 GNDA.n1039 185
R2923 GNDA.n1037 GNDA.n698 185
R2924 GNDA.n1035 GNDA.n1034 185
R2925 GNDA.n1033 GNDA.n699 185
R2926 GNDA.n699 GNDA.t139 185
R2927 GNDA.n1032 GNDA.n1031 185
R2928 GNDA.n1029 GNDA.n700 185
R2929 GNDA.n1119 GNDA.n1118 185
R2930 GNDA.n1120 GNDA.n1117 185
R2931 GNDA.n1120 GNDA.t114 185
R2932 GNDA.n1123 GNDA.n1122 185
R2933 GNDA.n1124 GNDA.n1116 185
R2934 GNDA.n1126 GNDA.n1125 185
R2935 GNDA.n1128 GNDA.n1115 185
R2936 GNDA.n1131 GNDA.n1130 185
R2937 GNDA.n1132 GNDA.n1114 185
R2938 GNDA.n1134 GNDA.n1133 185
R2939 GNDA.n1136 GNDA.n1113 185
R2940 GNDA.n1139 GNDA.n1138 185
R2941 GNDA.n1140 GNDA.n1112 185
R2942 GNDA.n1142 GNDA.n1141 185
R2943 GNDA.n1144 GNDA.n1111 185
R2944 GNDA.n1147 GNDA.n1146 185
R2945 GNDA.n1148 GNDA.n1110 185
R2946 GNDA.n1150 GNDA.n1149 185
R2947 GNDA.n1152 GNDA.n1109 185
R2948 GNDA.n1169 GNDA.n1104 185
R2949 GNDA.n1167 GNDA.n1166 185
R2950 GNDA.n1165 GNDA.n1105 185
R2951 GNDA.n1164 GNDA.n1163 185
R2952 GNDA.n1161 GNDA.n1106 185
R2953 GNDA.n1159 GNDA.n1158 185
R2954 GNDA.n1157 GNDA.n1107 185
R2955 GNDA.n1107 GNDA.t114 185
R2956 GNDA.n1156 GNDA.n1155 185
R2957 GNDA.n1153 GNDA.n1108 185
R2958 GNDA.n1761 GNDA.n1760 185
R2959 GNDA.n1762 GNDA.n1758 185
R2960 GNDA.n1758 GNDA.t113 185
R2961 GNDA.n1764 GNDA.n1763 185
R2962 GNDA.n1766 GNDA.n1757 185
R2963 GNDA.n1769 GNDA.n1768 185
R2964 GNDA.n1770 GNDA.n1756 185
R2965 GNDA.n1772 GNDA.n1771 185
R2966 GNDA.n1774 GNDA.n1755 185
R2967 GNDA.n1777 GNDA.n1776 185
R2968 GNDA.n1778 GNDA.n1754 185
R2969 GNDA.n1780 GNDA.n1779 185
R2970 GNDA.n1782 GNDA.n1753 185
R2971 GNDA.n1785 GNDA.n1784 185
R2972 GNDA.n1786 GNDA.n1752 185
R2973 GNDA.n1788 GNDA.n1787 185
R2974 GNDA.n1790 GNDA.n1751 185
R2975 GNDA.n1793 GNDA.n1792 185
R2976 GNDA.n1794 GNDA.n1750 185
R2977 GNDA.n1811 GNDA.n1810 185
R2978 GNDA.n1808 GNDA.n1743 185
R2979 GNDA.n1807 GNDA.n1746 185
R2980 GNDA.n1805 GNDA.n1804 185
R2981 GNDA.n1803 GNDA.n1747 185
R2982 GNDA.n1802 GNDA.n1801 185
R2983 GNDA.n1799 GNDA.n1748 185
R2984 GNDA.n1799 GNDA.t113 185
R2985 GNDA.n1798 GNDA.n1749 185
R2986 GNDA.n1796 GNDA.n1795 185
R2987 GNDA.n1969 GNDA.n1931 185
R2988 GNDA.n1971 GNDA.n1970 185
R2989 GNDA.n1970 GNDA.t115 185
R2990 GNDA.n1973 GNDA.n1972 185
R2991 GNDA.n1975 GNDA.n1968 185
R2992 GNDA.n1978 GNDA.n1977 185
R2993 GNDA.n1979 GNDA.n1967 185
R2994 GNDA.n1981 GNDA.n1980 185
R2995 GNDA.n1983 GNDA.n1966 185
R2996 GNDA.n1986 GNDA.n1985 185
R2997 GNDA.n1987 GNDA.n1965 185
R2998 GNDA.n1989 GNDA.n1988 185
R2999 GNDA.n1991 GNDA.n1964 185
R3000 GNDA.n1994 GNDA.n1993 185
R3001 GNDA.n1995 GNDA.n1963 185
R3002 GNDA.n1997 GNDA.n1996 185
R3003 GNDA.n1999 GNDA.n1962 185
R3004 GNDA.n2002 GNDA.n2001 185
R3005 GNDA.n2003 GNDA.n1961 185
R3006 GNDA.n2020 GNDA.n2019 185
R3007 GNDA.n2017 GNDA.n1954 185
R3008 GNDA.n2016 GNDA.n1957 185
R3009 GNDA.n2014 GNDA.n2013 185
R3010 GNDA.n2012 GNDA.n1958 185
R3011 GNDA.n2011 GNDA.n2010 185
R3012 GNDA.n2008 GNDA.n1959 185
R3013 GNDA.n2008 GNDA.t115 185
R3014 GNDA.n2007 GNDA.n1960 185
R3015 GNDA.n2005 GNDA.n2004 185
R3016 GNDA.n2354 GNDA.n138 185
R3017 GNDA.n2355 GNDA.n137 185
R3018 GNDA.n2355 GNDA.t95 185
R3019 GNDA.n2358 GNDA.n2357 185
R3020 GNDA.n2359 GNDA.n136 185
R3021 GNDA.n2361 GNDA.n2360 185
R3022 GNDA.n2363 GNDA.n135 185
R3023 GNDA.n2366 GNDA.n2365 185
R3024 GNDA.n2367 GNDA.n134 185
R3025 GNDA.n2369 GNDA.n2368 185
R3026 GNDA.n2371 GNDA.n133 185
R3027 GNDA.n2374 GNDA.n2373 185
R3028 GNDA.n2375 GNDA.n132 185
R3029 GNDA.n2377 GNDA.n2376 185
R3030 GNDA.n2379 GNDA.n131 185
R3031 GNDA.n2382 GNDA.n2381 185
R3032 GNDA.n2383 GNDA.n130 185
R3033 GNDA.n2385 GNDA.n2384 185
R3034 GNDA.n2387 GNDA.n129 185
R3035 GNDA.n2404 GNDA.n89 185
R3036 GNDA.n2402 GNDA.n2401 185
R3037 GNDA.n2400 GNDA.n125 185
R3038 GNDA.n2399 GNDA.n2398 185
R3039 GNDA.n2396 GNDA.n126 185
R3040 GNDA.n2394 GNDA.n2393 185
R3041 GNDA.n2392 GNDA.n127 185
R3042 GNDA.n127 GNDA.t95 185
R3043 GNDA.n2391 GNDA.n2390 185
R3044 GNDA.n2388 GNDA.n128 185
R3045 GNDA.n2405 GNDA.n88 185
R3046 GNDA.n2409 GNDA.n2407 185
R3047 GNDA.n2414 GNDA.n2413 185
R3048 GNDA.n2417 GNDA.n2416 185
R3049 GNDA.n124 GNDA.n122 185
R3050 GNDA.n2343 GNDA.n2342 185
R3051 GNDA.n2340 GNDA.n2337 185
R3052 GNDA.n141 GNDA.n139 185
R3053 GNDA.n2352 GNDA.n2351 185
R3054 GNDA.n1956 GNDA.n1953 185
R3055 GNDA.n1945 GNDA.n1943 185
R3056 GNDA.n2036 GNDA.n2035 185
R3057 GNDA.n2038 GNDA.n1942 185
R3058 GNDA.n2040 GNDA.n2039 185
R3059 GNDA.n1937 GNDA.n1935 185
R3060 GNDA.n2051 GNDA.n2050 185
R3061 GNDA.n2053 GNDA.n1934 185
R3062 GNDA.n2055 GNDA.n2054 185
R3063 GNDA.n1745 GNDA.n1742 185
R3064 GNDA.n1607 GNDA.n1606 185
R3065 GNDA.n1827 GNDA.n1826 185
R3066 GNDA.n1830 GNDA.n1829 185
R3067 GNDA.n1605 GNDA.n1602 185
R3068 GNDA.n613 GNDA.n612 185
R3069 GNDA.n1839 GNDA.n1838 185
R3070 GNDA.n1842 GNDA.n1841 185
R3071 GNDA.n611 GNDA.n609 185
R3072 GNDA.n1171 GNDA.n1170 185
R3073 GNDA.n1093 GNDA.n1091 185
R3074 GNDA.n1178 GNDA.n1177 185
R3075 GNDA.n1180 GNDA.n1090 185
R3076 GNDA.n1182 GNDA.n1181 185
R3077 GNDA.n1084 GNDA.n1082 185
R3078 GNDA.n1189 GNDA.n1188 185
R3079 GNDA.n1191 GNDA.n1081 185
R3080 GNDA.n1193 GNDA.n1192 185
R3081 GNDA.n1047 GNDA.n1046 185
R3082 GNDA.n970 GNDA.n969 185
R3083 GNDA.n968 GNDA.n966 185
R3084 GNDA.n975 GNDA.n965 185
R3085 GNDA.n980 GNDA.n979 185
R3086 GNDA.n983 GNDA.n982 185
R3087 GNDA.n964 GNDA.n961 185
R3088 GNDA.n988 GNDA.n711 185
R3089 GNDA.n993 GNDA.n992 185
R3090 GNDA.n847 GNDA.n846 185
R3091 GNDA.n765 GNDA.n763 185
R3092 GNDA.n854 GNDA.n853 185
R3093 GNDA.n856 GNDA.n762 185
R3094 GNDA.n858 GNDA.n857 185
R3095 GNDA.n756 GNDA.n754 185
R3096 GNDA.n865 GNDA.n864 185
R3097 GNDA.n867 GNDA.n753 185
R3098 GNDA.n869 GNDA.n868 185
R3099 GNDA.n2261 GNDA.n2260 185
R3100 GNDA.n298 GNDA.n296 185
R3101 GNDA.n2268 GNDA.n2267 185
R3102 GNDA.n2270 GNDA.n295 185
R3103 GNDA.n2272 GNDA.n2271 185
R3104 GNDA.n289 GNDA.n287 185
R3105 GNDA.n2279 GNDA.n2278 185
R3106 GNDA.n2281 GNDA.n286 185
R3107 GNDA.n2283 GNDA.n2282 185
R3108 GNDA.n1362 GNDA.n1361 185
R3109 GNDA.n1285 GNDA.n1283 185
R3110 GNDA.n1369 GNDA.n1368 185
R3111 GNDA.n1371 GNDA.n1282 185
R3112 GNDA.n1373 GNDA.n1372 185
R3113 GNDA.n1276 GNDA.n1274 185
R3114 GNDA.n1380 GNDA.n1379 185
R3115 GNDA.n1382 GNDA.n1273 185
R3116 GNDA.n1384 GNDA.n1383 185
R3117 GNDA.n1397 GNDA.n1395 185
R3118 GNDA.n1469 GNDA.n1467 185
R3119 GNDA.n1471 GNDA.n1470 185
R3120 GNDA.n1459 GNDA.n1457 185
R3121 GNDA.n1478 GNDA.n1477 185
R3122 GNDA.n1480 GNDA.n1456 185
R3123 GNDA.n1482 GNDA.n1481 185
R3124 GNDA.n1414 GNDA.n1412 185
R3125 GNDA.n1489 GNDA.n1488 185
R3126 GNDA.n466 GNDA.n464 182.4
R3127 GNDA.n52 GNDA.n46 182.4
R3128 GNDA.n2062 GNDA.n2061 181.233
R3129 GNDA.n2097 GNDA.n144 181.233
R3130 GNDA.n1694 GNDA.n1630 179.917
R3131 GNDA.n1728 GNDA.n1620 176
R3132 GNDA.n1728 GNDA.n1727 176
R3133 GNDA.n484 GNDA.n323 176
R3134 GNDA.n2468 GNDA.n49 176
R3135 GNDA.n2285 GNDA.n283 175.546
R3136 GNDA.n2276 GNDA.n291 175.546
R3137 GNDA.n2274 GNDA.n292 175.546
R3138 GNDA.n2265 GNDA.n300 175.546
R3139 GNDA.n2263 GNDA.n301 175.546
R3140 GNDA.n499 GNDA.n174 175.546
R3141 GNDA.n503 GNDA.n499 175.546
R3142 GNDA.n503 GNDA.n497 175.546
R3143 GNDA.n2161 GNDA.n497 175.546
R3144 GNDA.n2161 GNDA.n494 175.546
R3145 GNDA.n2167 GNDA.n494 175.546
R3146 GNDA.n2167 GNDA.n495 175.546
R3147 GNDA.n495 GNDA.n308 175.546
R3148 GNDA.n2185 GNDA.n308 175.546
R3149 GNDA.n2186 GNDA.n2185 175.546
R3150 GNDA.n2306 GNDA.n180 175.546
R3151 GNDA.n2310 GNDA.n2308 175.546
R3152 GNDA.n2314 GNDA.n178 175.546
R3153 GNDA.n2318 GNDA.n2316 175.546
R3154 GNDA.n2322 GNDA.n176 175.546
R3155 GNDA.n258 GNDA.n257 175.546
R3156 GNDA.n263 GNDA.n262 175.546
R3157 GNDA.n269 GNDA.n268 175.546
R3158 GNDA.n275 GNDA.n274 175.546
R3159 GNDA.n2290 GNDA.n2289 175.546
R3160 GNDA.n2333 GNDA.n142 175.546
R3161 GNDA.n2349 GNDA.n142 175.546
R3162 GNDA.n2349 GNDA.n143 175.546
R3163 GNDA.n2345 GNDA.n143 175.546
R3164 GNDA.n2345 GNDA.n120 175.546
R3165 GNDA.n2419 GNDA.n120 175.546
R3166 GNDA.n2419 GNDA.n121 175.546
R3167 GNDA.n2411 GNDA.n121 175.546
R3168 GNDA.n2411 GNDA.n86 175.546
R3169 GNDA.n2442 GNDA.n86 175.546
R3170 GNDA.n2442 GNDA.n87 175.546
R3171 GNDA.n230 GNDA.n216 175.546
R3172 GNDA.n226 GNDA.n216 175.546
R3173 GNDA.n226 GNDA.n219 175.546
R3174 GNDA.n222 GNDA.n219 175.546
R3175 GNDA.n222 GNDA.n114 175.546
R3176 GNDA.n2422 GNDA.n114 175.546
R3177 GNDA.n2422 GNDA.n108 175.546
R3178 GNDA.n2427 GNDA.n108 175.546
R3179 GNDA.n2427 GNDA.n112 175.546
R3180 GNDA.n112 GNDA.n111 175.546
R3181 GNDA.n252 GNDA.n251 175.546
R3182 GNDA.n248 GNDA.n247 175.546
R3183 GNDA.n245 GNDA.n211 175.546
R3184 GNDA.n241 GNDA.n239 175.546
R3185 GNDA.n237 GNDA.n213 175.546
R3186 GNDA.n1217 GNDA.n160 175.546
R3187 GNDA.n1219 GNDA.n1218 175.546
R3188 GNDA.n1221 GNDA.n1220 175.546
R3189 GNDA.n1223 GNDA.n1222 175.546
R3190 GNDA.n1224 GNDA.n147 175.546
R3191 GNDA.n2059 GNDA.n568 175.546
R3192 GNDA.n2043 GNDA.n568 175.546
R3193 GNDA.n2043 GNDA.n1938 175.546
R3194 GNDA.n2048 GNDA.n1938 175.546
R3195 GNDA.n2048 GNDA.n2042 175.546
R3196 GNDA.n2042 GNDA.n1939 175.546
R3197 GNDA.n1946 GNDA.n1939 175.546
R3198 GNDA.n2033 GNDA.n1946 175.546
R3199 GNDA.n2033 GNDA.n1947 175.546
R3200 GNDA.n2029 GNDA.n1947 175.546
R3201 GNDA.n2029 GNDA.n1951 175.546
R3202 GNDA.n1241 GNDA.n1240 175.546
R3203 GNDA.n1237 GNDA.n1236 175.546
R3204 GNDA.n1233 GNDA.n1232 175.546
R3205 GNDA.n1229 GNDA.n1228 175.546
R3206 GNDA.n1225 GNDA.n198 175.546
R3207 GNDA.n1266 GNDA.n1214 175.546
R3208 GNDA.n1262 GNDA.n1261 175.546
R3209 GNDA.n1258 GNDA.n1257 175.546
R3210 GNDA.n1254 GNDA.n1253 175.546
R3211 GNDA.n1250 GNDA.n1249 175.546
R3212 GNDA.n1902 GNDA.n1901 175.546
R3213 GNDA.n1905 GNDA.n1904 175.546
R3214 GNDA.n1914 GNDA.n1913 175.546
R3215 GNDA.n1918 GNDA.n1917 175.546
R3216 GNDA.n1927 GNDA.n570 175.546
R3217 GNDA.n1386 GNDA.n1270 175.546
R3218 GNDA.n1377 GNDA.n1278 175.546
R3219 GNDA.n1375 GNDA.n1279 175.546
R3220 GNDA.n1366 GNDA.n1287 175.546
R3221 GNDA.n1364 GNDA.n1288 175.546
R3222 GNDA.n259 GNDA.n185 175.546
R3223 GNDA.n265 GNDA.n264 175.546
R3224 GNDA.n271 GNDA.n270 175.546
R3225 GNDA.n277 GNDA.n276 175.546
R3226 GNDA.n279 GNDA.n187 175.546
R3227 GNDA.n679 GNDA.n660 175.546
R3228 GNDA.n677 GNDA.n676 175.546
R3229 GNDA.n673 GNDA.n672 175.546
R3230 GNDA.n669 GNDA.n668 175.546
R3231 GNDA.n665 GNDA.n664 175.546
R3232 GNDA.n636 GNDA.n633 175.546
R3233 GNDA.n639 GNDA.n638 175.546
R3234 GNDA.n644 GNDA.n641 175.546
R3235 GNDA.n647 GNDA.n646 175.546
R3236 GNDA.n651 GNDA.n649 175.546
R3237 GNDA.n1848 GNDA.n605 175.546
R3238 GNDA.n1844 GNDA.n605 175.546
R3239 GNDA.n1844 GNDA.n607 175.546
R3240 GNDA.n1836 GNDA.n607 175.546
R3241 GNDA.n1836 GNDA.n614 175.546
R3242 GNDA.n1832 GNDA.n614 175.546
R3243 GNDA.n1832 GNDA.n1600 175.546
R3244 GNDA.n1824 GNDA.n1600 175.546
R3245 GNDA.n1824 GNDA.n1608 175.546
R3246 GNDA.n1820 GNDA.n1608 175.546
R3247 GNDA.n1820 GNDA.n1740 175.546
R3248 GNDA.n1907 GNDA.n578 175.546
R3249 GNDA.n1911 GNDA.n1909 175.546
R3250 GNDA.n1920 GNDA.n574 175.546
R3251 GNDA.n1923 GNDA.n1922 175.546
R3252 GNDA.n1925 GNDA.n572 175.546
R3253 GNDA.n1878 GNDA.n589 175.546
R3254 GNDA.n1882 GNDA.n1880 175.546
R3255 GNDA.n1886 GNDA.n587 175.546
R3256 GNDA.n1890 GNDA.n1888 175.546
R3257 GNDA.n1894 GNDA.n585 175.546
R3258 GNDA.n1872 GNDA.n591 175.546
R3259 GNDA.n1868 GNDA.n591 175.546
R3260 GNDA.n1868 GNDA.n594 175.546
R3261 GNDA.n1864 GNDA.n594 175.546
R3262 GNDA.n1864 GNDA.n597 175.546
R3263 GNDA.n1860 GNDA.n597 175.546
R3264 GNDA.n1860 GNDA.n599 175.546
R3265 GNDA.n1856 GNDA.n599 175.546
R3266 GNDA.n1856 GNDA.n601 175.546
R3267 GNDA.n1852 GNDA.n601 175.546
R3268 GNDA.n1486 GNDA.n1452 175.546
R3269 GNDA.n1484 GNDA.n1453 175.546
R3270 GNDA.n1475 GNDA.n1461 175.546
R3271 GNDA.n1473 GNDA.n1463 175.546
R3272 GNDA.n1545 GNDA.n1394 175.546
R3273 GNDA.n1569 GNDA.n1568 175.546
R3274 GNDA.n1566 GNDA.n635 175.546
R3275 GNDA.n1562 GNDA.n1560 175.546
R3276 GNDA.n1558 GNDA.n643 175.546
R3277 GNDA.n1554 GNDA.n1552 175.546
R3278 GNDA.n1592 GNDA.n625 175.546
R3279 GNDA.n1590 GNDA.n1589 175.546
R3280 GNDA.n1586 GNDA.n1585 175.546
R3281 GNDA.n1582 GNDA.n1581 175.546
R3282 GNDA.n1578 GNDA.n1577 175.546
R3283 GNDA.n1425 GNDA.n626 175.546
R3284 GNDA.n1429 GNDA.n1425 175.546
R3285 GNDA.n1429 GNDA.n1423 175.546
R3286 GNDA.n1433 GNDA.n1423 175.546
R3287 GNDA.n1433 GNDA.n1421 175.546
R3288 GNDA.n1437 GNDA.n1421 175.546
R3289 GNDA.n1437 GNDA.n1419 175.546
R3290 GNDA.n1441 GNDA.n1419 175.546
R3291 GNDA.n1441 GNDA.n1417 175.546
R3292 GNDA.n1446 GNDA.n1417 175.546
R3293 GNDA.n871 GNDA.n749 175.546
R3294 GNDA.n862 GNDA.n758 175.546
R3295 GNDA.n860 GNDA.n759 175.546
R3296 GNDA.n851 GNDA.n767 175.546
R3297 GNDA.n849 GNDA.n768 175.546
R3298 GNDA.n896 GNDA.n737 175.546
R3299 GNDA.n892 GNDA.n737 175.546
R3300 GNDA.n892 GNDA.n739 175.546
R3301 GNDA.n888 GNDA.n739 175.546
R3302 GNDA.n888 GNDA.n741 175.546
R3303 GNDA.n884 GNDA.n741 175.546
R3304 GNDA.n884 GNDA.n743 175.546
R3305 GNDA.n880 GNDA.n743 175.546
R3306 GNDA.n880 GNDA.n745 175.546
R3307 GNDA.n876 GNDA.n745 175.546
R3308 GNDA.n932 GNDA.n722 175.546
R3309 GNDA.n936 GNDA.n934 175.546
R3310 GNDA.n946 GNDA.n718 175.546
R3311 GNDA.n949 GNDA.n948 175.546
R3312 GNDA.n951 GNDA.n716 175.546
R3313 GNDA.n900 GNDA.n735 175.546
R3314 GNDA.n900 GNDA.n733 175.546
R3315 GNDA.n905 GNDA.n733 175.546
R3316 GNDA.n905 GNDA.n731 175.546
R3317 GNDA.n909 GNDA.n731 175.546
R3318 GNDA.n910 GNDA.n909 175.546
R3319 GNDA.n912 GNDA.n910 175.546
R3320 GNDA.n912 GNDA.n729 175.546
R3321 GNDA.n917 GNDA.n729 175.546
R3322 GNDA.n917 GNDA.n725 175.546
R3323 GNDA.n921 GNDA.n725 175.546
R3324 GNDA.n990 GNDA.n989 175.546
R3325 GNDA.n986 GNDA.n985 175.546
R3326 GNDA.n977 GNDA.n976 175.546
R3327 GNDA.n973 GNDA.n972 175.546
R3328 GNDA.n694 GNDA.n691 175.546
R3329 GNDA.n930 GNDA.n928 175.546
R3330 GNDA.n938 GNDA.n720 175.546
R3331 GNDA.n944 GNDA.n940 175.546
R3332 GNDA.n942 GNDA.n941 175.546
R3333 GNDA.n954 GNDA.n953 175.546
R3334 GNDA.n1054 GNDA.n1053 175.546
R3335 GNDA.n1060 GNDA.n1059 175.546
R3336 GNDA.n1066 GNDA.n1065 175.546
R3337 GNDA.n1072 GNDA.n1071 175.546
R3338 GNDA.n1074 GNDA.n192 175.546
R3339 GNDA.n2064 GNDA.n561 175.546
R3340 GNDA.n2064 GNDA.n559 175.546
R3341 GNDA.n2068 GNDA.n559 175.546
R3342 GNDA.n2068 GNDA.n557 175.546
R3343 GNDA.n2072 GNDA.n557 175.546
R3344 GNDA.n2072 GNDA.n547 175.546
R3345 GNDA.n2082 GNDA.n547 175.546
R3346 GNDA.n2082 GNDA.n545 175.546
R3347 GNDA.n2087 GNDA.n545 175.546
R3348 GNDA.n2087 GNDA.n541 175.546
R3349 GNDA.n2091 GNDA.n541 175.546
R3350 GNDA.n1195 GNDA.n1078 175.546
R3351 GNDA.n1186 GNDA.n1086 175.546
R3352 GNDA.n1184 GNDA.n1087 175.546
R3353 GNDA.n1175 GNDA.n1095 175.546
R3354 GNDA.n1173 GNDA.n1096 175.546
R3355 GNDA.n2126 GNDA.n526 175.546
R3356 GNDA.n2130 GNDA.n526 175.546
R3357 GNDA.n2130 GNDA.n524 175.546
R3358 GNDA.n2135 GNDA.n524 175.546
R3359 GNDA.n2135 GNDA.n522 175.546
R3360 GNDA.n2139 GNDA.n522 175.546
R3361 GNDA.n2139 GNDA.n521 175.546
R3362 GNDA.n2143 GNDA.n521 175.546
R3363 GNDA.n2143 GNDA.n517 175.546
R3364 GNDA.n2148 GNDA.n517 175.546
R3365 GNDA.n2099 GNDA.n2096 175.546
R3366 GNDA.n2099 GNDA.n536 175.546
R3367 GNDA.n2103 GNDA.n536 175.546
R3368 GNDA.n2103 GNDA.n534 175.546
R3369 GNDA.n2107 GNDA.n534 175.546
R3370 GNDA.n2107 GNDA.n532 175.546
R3371 GNDA.n2111 GNDA.n532 175.546
R3372 GNDA.n2111 GNDA.n530 175.546
R3373 GNDA.n2116 GNDA.n530 175.546
R3374 GNDA.n2116 GNDA.n528 175.546
R3375 GNDA.n2120 GNDA.n528 175.546
R3376 GNDA.n1052 GNDA.n1051 175.546
R3377 GNDA.n1058 GNDA.n1057 175.546
R3378 GNDA.n1064 GNDA.n1063 175.546
R3379 GNDA.n1070 GNDA.n1069 175.546
R3380 GNDA.n1200 GNDA.n1199 175.546
R3381 GNDA.n1720 GNDA.n1719 164.369
R3382 GNDA.n1645 GNDA.n1644 164.369
R3383 GNDA.n1541 GNDA.n1397 163.333
R3384 GNDA.n1361 GNDA.n1360 163.333
R3385 GNDA.n2260 GNDA.n2259 163.333
R3386 GNDA.n846 GNDA.n845 163.333
R3387 GNDA.n1046 GNDA.n1045 163.333
R3388 GNDA.n1170 GNDA.n1169 163.333
R3389 GNDA.n1810 GNDA.n1745 163.333
R3390 GNDA.n2019 GNDA.n1956 163.333
R3391 GNDA.n2405 GNDA.n2404 163.333
R3392 GNDA.n1649 GNDA.t142 160.725
R3393 GNDA.n1650 GNDA.t138 160.725
R3394 GNDA.n1621 GNDA.t129 160.725
R3395 GNDA.n1619 GNDA.t112 160.725
R3396 GNDA.n1623 GNDA.t154 160.725
R3397 GNDA.n1708 GNDA.t169 160.725
R3398 GNDA.n553 GNDA.t179 157.555
R3399 GNDA.n552 GNDA.t28 157.555
R3400 GNDA.n419 GNDA.n418 156.8
R3401 GNDA.n358 GNDA.n331 153.601
R3402 GNDA.n2470 GNDA.n45 153.601
R3403 GNDA.n1653 GNDA.t2 153.294
R3404 GNDA.n462 GNDA.t107 152.994
R3405 GNDA.n322 GNDA.t94 152.994
R3406 GNDA.n48 GNDA.t99 152.994
R3407 GNDA.n51 GNDA.t82 152.994
R3408 GNDA.n2329 GNDA.n2328 152.643
R3409 GNDA.n1929 GNDA.n1928 152.643
R3410 GNDA.n101 GNDA.n93 150.988
R3411 GNDA.n2483 GNDA.n2482 150.4
R3412 GNDA.n1489 GNDA.n1412 150
R3413 GNDA.n1481 GNDA.n1480 150
R3414 GNDA.n1478 GNDA.n1457 150
R3415 GNDA.n1470 GNDA.n1469 150
R3416 GNDA.n1530 GNDA.n1529 150
R3417 GNDA.n1532 GNDA.n1530 150
R3418 GNDA.n1536 GNDA.n1399 150
R3419 GNDA.n1539 GNDA.n1538 150
R3420 GNDA.n1511 GNDA.n1406 150
R3421 GNDA.n1515 GNDA.n1513 150
R3422 GNDA.n1519 GNDA.n1404 150
R3423 GNDA.n1523 GNDA.n1521 150
R3424 GNDA.n1507 GNDA.n1505 150
R3425 GNDA.n1503 GNDA.n1408 150
R3426 GNDA.n1499 GNDA.n1497 150
R3427 GNDA.n1495 GNDA.n1410 150
R3428 GNDA.n1491 GNDA.n1410 150
R3429 GNDA.n1383 GNDA.n1382 150
R3430 GNDA.n1380 GNDA.n1274 150
R3431 GNDA.n1372 GNDA.n1371 150
R3432 GNDA.n1369 GNDA.n1283 150
R3433 GNDA.n1346 GNDA.n1298 150
R3434 GNDA.n1350 GNDA.n1298 150
R3435 GNDA.n1354 GNDA.n1352 150
R3436 GNDA.n1358 GNDA.n1296 150
R3437 GNDA.n1329 GNDA.n1327 150
R3438 GNDA.n1333 GNDA.n1303 150
R3439 GNDA.n1337 GNDA.n1335 150
R3440 GNDA.n1341 GNDA.n1301 150
R3441 GNDA.n1325 GNDA.n1305 150
R3442 GNDA.n1321 GNDA.n1319 150
R3443 GNDA.n1317 GNDA.n1307 150
R3444 GNDA.n1313 GNDA.n1311 150
R3445 GNDA.n1311 GNDA.n1310 150
R3446 GNDA.n2282 GNDA.n2281 150
R3447 GNDA.n2279 GNDA.n287 150
R3448 GNDA.n2271 GNDA.n2270 150
R3449 GNDA.n2268 GNDA.n296 150
R3450 GNDA.n2245 GNDA.n2197 150
R3451 GNDA.n2249 GNDA.n2197 150
R3452 GNDA.n2253 GNDA.n2251 150
R3453 GNDA.n2257 GNDA.n2195 150
R3454 GNDA.n2228 GNDA.n2226 150
R3455 GNDA.n2232 GNDA.n2202 150
R3456 GNDA.n2236 GNDA.n2234 150
R3457 GNDA.n2240 GNDA.n2200 150
R3458 GNDA.n2224 GNDA.n2204 150
R3459 GNDA.n2220 GNDA.n2218 150
R3460 GNDA.n2216 GNDA.n2206 150
R3461 GNDA.n2212 GNDA.n2210 150
R3462 GNDA.n2210 GNDA.n2209 150
R3463 GNDA.n868 GNDA.n867 150
R3464 GNDA.n865 GNDA.n754 150
R3465 GNDA.n857 GNDA.n856 150
R3466 GNDA.n854 GNDA.n763 150
R3467 GNDA.n831 GNDA.n783 150
R3468 GNDA.n835 GNDA.n783 150
R3469 GNDA.n839 GNDA.n837 150
R3470 GNDA.n843 GNDA.n781 150
R3471 GNDA.n814 GNDA.n812 150
R3472 GNDA.n818 GNDA.n788 150
R3473 GNDA.n822 GNDA.n820 150
R3474 GNDA.n826 GNDA.n786 150
R3475 GNDA.n810 GNDA.n790 150
R3476 GNDA.n806 GNDA.n804 150
R3477 GNDA.n802 GNDA.n792 150
R3478 GNDA.n798 GNDA.n796 150
R3479 GNDA.n796 GNDA.n795 150
R3480 GNDA.n993 GNDA.n711 150
R3481 GNDA.n982 GNDA.n964 150
R3482 GNDA.n980 GNDA.n965 150
R3483 GNDA.n969 GNDA.n968 150
R3484 GNDA.n1031 GNDA.n699 150
R3485 GNDA.n1035 GNDA.n699 150
R3486 GNDA.n1039 GNDA.n1037 150
R3487 GNDA.n1043 GNDA.n697 150
R3488 GNDA.n1014 GNDA.n1012 150
R3489 GNDA.n1018 GNDA.n704 150
R3490 GNDA.n1022 GNDA.n1020 150
R3491 GNDA.n1026 GNDA.n702 150
R3492 GNDA.n1010 GNDA.n706 150
R3493 GNDA.n1006 GNDA.n1004 150
R3494 GNDA.n1002 GNDA.n708 150
R3495 GNDA.n998 GNDA.n996 150
R3496 GNDA.n996 GNDA.n995 150
R3497 GNDA.n1192 GNDA.n1191 150
R3498 GNDA.n1189 GNDA.n1082 150
R3499 GNDA.n1181 GNDA.n1180 150
R3500 GNDA.n1178 GNDA.n1091 150
R3501 GNDA.n1155 GNDA.n1107 150
R3502 GNDA.n1159 GNDA.n1107 150
R3503 GNDA.n1163 GNDA.n1161 150
R3504 GNDA.n1167 GNDA.n1105 150
R3505 GNDA.n1138 GNDA.n1136 150
R3506 GNDA.n1142 GNDA.n1112 150
R3507 GNDA.n1146 GNDA.n1144 150
R3508 GNDA.n1150 GNDA.n1110 150
R3509 GNDA.n1134 GNDA.n1114 150
R3510 GNDA.n1130 GNDA.n1128 150
R3511 GNDA.n1126 GNDA.n1116 150
R3512 GNDA.n1122 GNDA.n1120 150
R3513 GNDA.n1120 GNDA.n1119 150
R3514 GNDA.n1841 GNDA.n611 150
R3515 GNDA.n1839 GNDA.n612 150
R3516 GNDA.n1829 GNDA.n1605 150
R3517 GNDA.n1827 GNDA.n1606 150
R3518 GNDA.n1799 GNDA.n1798 150
R3519 GNDA.n1801 GNDA.n1799 150
R3520 GNDA.n1805 GNDA.n1747 150
R3521 GNDA.n1808 GNDA.n1807 150
R3522 GNDA.n1780 GNDA.n1754 150
R3523 GNDA.n1784 GNDA.n1782 150
R3524 GNDA.n1788 GNDA.n1752 150
R3525 GNDA.n1792 GNDA.n1790 150
R3526 GNDA.n1776 GNDA.n1774 150
R3527 GNDA.n1772 GNDA.n1756 150
R3528 GNDA.n1768 GNDA.n1766 150
R3529 GNDA.n1764 GNDA.n1758 150
R3530 GNDA.n1760 GNDA.n1758 150
R3531 GNDA.n2054 GNDA.n2053 150
R3532 GNDA.n2051 GNDA.n1935 150
R3533 GNDA.n2039 GNDA.n2038 150
R3534 GNDA.n2036 GNDA.n1943 150
R3535 GNDA.n2008 GNDA.n2007 150
R3536 GNDA.n2010 GNDA.n2008 150
R3537 GNDA.n2014 GNDA.n1958 150
R3538 GNDA.n2017 GNDA.n2016 150
R3539 GNDA.n1989 GNDA.n1965 150
R3540 GNDA.n1993 GNDA.n1991 150
R3541 GNDA.n1997 GNDA.n1963 150
R3542 GNDA.n2001 GNDA.n1999 150
R3543 GNDA.n1985 GNDA.n1983 150
R3544 GNDA.n1981 GNDA.n1967 150
R3545 GNDA.n1977 GNDA.n1975 150
R3546 GNDA.n1973 GNDA.n1970 150
R3547 GNDA.n1970 GNDA.n1969 150
R3548 GNDA.n2352 GNDA.n139 150
R3549 GNDA.n2342 GNDA.n2340 150
R3550 GNDA.n2416 GNDA.n124 150
R3551 GNDA.n2414 GNDA.n2407 150
R3552 GNDA.n2390 GNDA.n127 150
R3553 GNDA.n2394 GNDA.n127 150
R3554 GNDA.n2398 GNDA.n2396 150
R3555 GNDA.n2402 GNDA.n125 150
R3556 GNDA.n2373 GNDA.n2371 150
R3557 GNDA.n2377 GNDA.n132 150
R3558 GNDA.n2381 GNDA.n2379 150
R3559 GNDA.n2385 GNDA.n130 150
R3560 GNDA.n2369 GNDA.n134 150
R3561 GNDA.n2365 GNDA.n2363 150
R3562 GNDA.n2361 GNDA.n136 150
R3563 GNDA.n2357 GNDA.n2355 150
R3564 GNDA.n2355 GNDA.n2354 150
R3565 GNDA.n550 GNDA.t30 148.906
R3566 GNDA.n550 GNDA.t73 148.653
R3567 GNDA.n362 GNDA.t106 147.511
R3568 GNDA.n470 GNDA.t159 147.511
R3569 GNDA.n458 GNDA.t175 147.511
R3570 GNDA.n456 GNDA.t81 147.511
R3571 GNDA.t153 GNDA.t337 145.403
R3572 GNDA.t312 GNDA.t137 145.403
R3573 GNDA.n93 GNDA.n85 145.013
R3574 GNDA.n1656 GNDA.n1654 139.638
R3575 GNDA.t111 GNDA.t277 139.081
R3576 GNDA.t277 GNDA.t273 139.081
R3577 GNDA.t273 GNDA.t208 139.081
R3578 GNDA.t269 GNDA.t250 139.081
R3579 GNDA.t12 GNDA.t269 139.081
R3580 GNDA.t128 GNDA.t12 139.081
R3581 GNDA.n1672 GNDA.n1671 139.077
R3582 GNDA.n1670 GNDA.n1669 139.077
R3583 GNDA.n1668 GNDA.n1667 139.077
R3584 GNDA.n1666 GNDA.n1665 139.077
R3585 GNDA.n1664 GNDA.n1663 139.077
R3586 GNDA.n1662 GNDA.n1661 139.077
R3587 GNDA.n1660 GNDA.n1659 139.077
R3588 GNDA.n1658 GNDA.n1657 139.077
R3589 GNDA.n1656 GNDA.n1655 139.077
R3590 GNDA.t239 GNDA.t124 135.386
R3591 GNDA.t244 GNDA.t308 135.386
R3592 GNDA.t87 GNDA.t303 135.386
R3593 GNDA.t150 GNDA.t304 135.386
R3594 GNDA.t299 GNDA.t336 135.386
R3595 GNDA.t204 GNDA.t121 135.386
R3596 GNDA.n482 GNDA.n481 134.867
R3597 GNDA.n2466 GNDA.n55 134.867
R3598 GNDA.n447 GNDA.n377 134.4
R3599 GNDA.n446 GNDA.n444 134.4
R3600 GNDA.n383 GNDA.n382 134.4
R3601 GNDA.n381 GNDA.n375 134.4
R3602 GNDA.n460 GNDA.n453 134.4
R3603 GNDA.n1731 GNDA.t208 132.76
R3604 GNDA.t250 GNDA.n1643 132.76
R3605 GNDA.n468 GNDA.n366 128
R3606 GNDA.n1712 GNDA.t32 126.438
R3607 GNDA.n1679 GNDA.t295 126.438
R3608 GNDA.n2191 GNDA.n2190 124.832
R3609 GNDA.n2325 GNDA.n2324 124.832
R3610 GNDA.n2437 GNDA.n87 124.832
R3611 GNDA.n233 GNDA.n231 124.832
R3612 GNDA.n2024 GNDA.n1951 124.832
R3613 GNDA.n1246 GNDA.n1245 124.832
R3614 GNDA.n1292 GNDA.n206 124.832
R3615 GNDA.n661 GNDA.n184 124.832
R3616 GNDA.n1815 GNDA.n1740 124.832
R3617 GNDA.n1897 GNDA.n1896 124.832
R3618 GNDA.n1548 GNDA.n1547 124.832
R3619 GNDA.n1574 GNDA.n1573 124.832
R3620 GNDA.n777 GNDA.n776 124.832
R3621 GNDA.n922 GNDA.n921 124.832
R3622 GNDA.n1206 GNDA.n692 124.832
R3623 GNDA.n2092 GNDA.n2091 124.832
R3624 GNDA.n1101 GNDA.n1099 124.832
R3625 GNDA.n2121 GNDA.n2120 124.832
R3626 GNDA.t41 GNDA.t285 120.115
R3627 GNDA.t282 GNDA.t49 120.115
R3628 GNDA.n2061 GNDA.n562 119.035
R3629 GNDA.n540 GNDA.n144 119.035
R3630 GNDA.n1651 GNDA.n1622 118.4
R3631 GNDA.n1677 GNDA.n1652 118.4
R3632 GNDA.n1724 GNDA.n1620 118.4
R3633 GNDA.n1727 GNDA.n1726 118.4
R3634 GNDA.n1710 GNDA.n1709 118.4
R3635 GNDA.n1723 GNDA.n1624 118.4
R3636 GNDA.n443 GNDA.t163 113.974
R3637 GNDA.n376 GNDA.t151 113.974
R3638 GNDA.n380 GNDA.t88 113.974
R3639 GNDA.n379 GNDA.t166 113.974
R3640 GNDA.n370 GNDA.t104 113.974
R3641 GNDA.n371 GNDA.t85 113.974
R3642 GNDA.n365 GNDA.t160 113.974
R3643 GNDA.n367 GNDA.t176 113.974
R3644 GNDA.n368 GNDA.t157 113.974
R3645 GNDA.n369 GNDA.t148 113.974
R3646 GNDA.t109 GNDA.n1833 113.624
R3647 GNDA.n1739 GNDA.n1738 113.624
R3648 GNDA.n1948 GNDA.t101 113.624
R3649 GNDA.t96 GNDA.n2420 113.624
R3650 GNDA.n437 GNDA.n436 108.8
R3651 GNDA.n434 GNDA.n433 108.8
R3652 GNDA.n2061 GNDA.n563 103.144
R3653 GNDA.n2296 GNDA.n144 103.144
R3654 GNDA.n1713 GNDA.n1712 101.15
R3655 GNDA.t320 GNDA.t33 101.15
R3656 GNDA.t318 GNDA.t1 101.15
R3657 GNDA.n1692 GNDA.n1679 101.15
R3658 GNDA.n2061 GNDA.n564 99.6276
R3659 GNDA.n2327 GNDA.n144 99.6276
R3660 GNDA.n414 GNDA.n413 99.0842
R3661 GNDA.n412 GNDA.n411 99.0842
R3662 GNDA.n410 GNDA.n409 99.0842
R3663 GNDA.n408 GNDA.n407 99.0842
R3664 GNDA.n406 GNDA.n405 99.0842
R3665 GNDA.n404 GNDA.n403 99.0842
R3666 GNDA.n402 GNDA.n401 99.0842
R3667 GNDA.n400 GNDA.n399 99.0842
R3668 GNDA.n398 GNDA.n397 99.0842
R3669 GNDA.n396 GNDA.n395 99.0842
R3670 GNDA.n394 GNDA.n393 99.0842
R3671 GNDA.n36 GNDA.n35 99.0842
R3672 GNDA.n2444 GNDA.n81 98.4712
R3673 GNDA.n901 GNDA.n734 96.5152
R3674 GNDA.n902 GNDA.n901 96.5152
R3675 GNDA.n904 GNDA.n902 96.5152
R3676 GNDA.n904 GNDA.n903 96.5152
R3677 GNDA.n903 GNDA.n615 96.5152
R3678 GNDA.n911 GNDA.n616 96.5152
R3679 GNDA.n911 GNDA.n728 96.5152
R3680 GNDA.n918 GNDA.n728 96.5152
R3681 GNDA.n919 GNDA.n918 96.5152
R3682 GNDA.n920 GNDA.n919 96.5152
R3683 GNDA.n920 GNDA.n562 96.5152
R3684 GNDA.n2063 GNDA.n2062 96.5152
R3685 GNDA.n2063 GNDA.n558 96.5152
R3686 GNDA.n2069 GNDA.n558 96.5152
R3687 GNDA.n2070 GNDA.n2069 96.5152
R3688 GNDA.n2071 GNDA.n2070 96.5152
R3689 GNDA.n2081 GNDA.n2080 96.5152
R3690 GNDA.n2081 GNDA.n544 96.5152
R3691 GNDA.n2088 GNDA.n544 96.5152
R3692 GNDA.n2089 GNDA.n2088 96.5152
R3693 GNDA.n2090 GNDA.n2089 96.5152
R3694 GNDA.n2090 GNDA.n540 96.5152
R3695 GNDA.n2098 GNDA.n2097 96.5152
R3696 GNDA.n2098 GNDA.n535 96.5152
R3697 GNDA.n2104 GNDA.n535 96.5152
R3698 GNDA.n2105 GNDA.n2104 96.5152
R3699 GNDA.n2106 GNDA.n2105 96.5152
R3700 GNDA.n2112 GNDA.n531 96.5152
R3701 GNDA.n2113 GNDA.n2112 96.5152
R3702 GNDA.n2115 GNDA.n2113 96.5152
R3703 GNDA.n2115 GNDA.n2114 96.5152
R3704 GNDA.n2114 GNDA.n316 96.5152
R3705 GNDA.n2176 GNDA.n490 95.7359
R3706 GNDA.n2444 GNDA.n84 95.4038
R3707 GNDA.n2476 GNDA.n37 95.101
R3708 GNDA.n477 GNDA.n474 95.101
R3709 GNDA.n2481 GNDA.t119 94.8842
R3710 GNDA.n416 GNDA.t132 94.8842
R3711 GNDA.t32 GNDA.t168 94.8281
R3712 GNDA.t216 GNDA.t235 94.8281
R3713 GNDA.t275 GNDA.t311 94.8281
R3714 GNDA.t295 GNDA.t141 94.8281
R3715 GNDA.n2478 GNDA.n2477 94.601
R3716 GNDA.n476 GNDA.n475 94.601
R3717 GNDA.t258 GNDA.t93 92.7208
R3718 GNDA.t207 GNDA.t338 92.7208
R3719 GNDA.t77 GNDA.t255 92.7208
R3720 GNDA.t317 GNDA.t183 92.7208
R3721 GNDA.t219 GNDA.t103 92.7208
R3722 GNDA.t103 GNDA.t201 92.7208
R3723 GNDA.t147 GNDA.t212 92.7208
R3724 GNDA.t34 GNDA.t147 92.7208
R3725 GNDA.t9 GNDA.t6 92.7208
R3726 GNDA.t8 GNDA.t227 92.7208
R3727 GNDA.t38 GNDA.t186 92.7208
R3728 GNDA.t98 GNDA.t266 92.7208
R3729 GNDA.t101 GNDA.n564 91.423
R3730 GNDA.n2327 GNDA.t96 91.423
R3731 GNDA.t134 GNDA.t59 88.5063
R3732 GNDA.t90 GNDA.t39 88.5063
R3733 GNDA.n485 GNDA.n321 86.4005
R3734 GNDA.n72 GNDA.n50 86.4005
R3735 GNDA.n1700 GNDA.n1699 85.2845
R3736 GNDA.n1633 GNDA.n1632 85.2845
R3737 GNDA.n549 GNDA.n548 84.306
R3738 GNDA.t288 GNDA.t43 82.1844
R3739 GNDA.t199 GNDA.t265 82.1844
R3740 GNDA.t210 GNDA.t310 82.1844
R3741 GNDA.t203 GNDA.t283 82.1844
R3742 GNDA.t144 GNDA.t258 80.0771
R3743 GNDA.t59 GNDA.t326 80.0771
R3744 GNDA.t39 GNDA.t21 80.0771
R3745 GNDA.t266 GNDA.t171 80.0771
R3746 GNDA.n467 GNDA.n466 80.0005
R3747 GNDA.n2286 GNDA.n2285 76.3222
R3748 GNDA.n291 GNDA.n290 76.3222
R3749 GNDA.n2275 GNDA.n2274 76.3222
R3750 GNDA.n300 GNDA.n299 76.3222
R3751 GNDA.n2264 GNDA.n2263 76.3222
R3752 GNDA.n2191 GNDA.n305 76.3222
R3753 GNDA.n2186 GNDA.n306 76.3222
R3754 GNDA.n2302 GNDA.n2301 76.3222
R3755 GNDA.n2307 GNDA.n2306 76.3222
R3756 GNDA.n2310 GNDA.n2309 76.3222
R3757 GNDA.n2315 GNDA.n2314 76.3222
R3758 GNDA.n2318 GNDA.n2317 76.3222
R3759 GNDA.n2323 GNDA.n2322 76.3222
R3760 GNDA.n2300 GNDA.n149 76.3222
R3761 GNDA.n258 GNDA.n150 76.3222
R3762 GNDA.n263 GNDA.n151 76.3222
R3763 GNDA.n269 GNDA.n152 76.3222
R3764 GNDA.n2289 GNDA.n153 76.3222
R3765 GNDA.n2290 GNDA.n148 76.3222
R3766 GNDA.n111 GNDA.n109 76.3222
R3767 GNDA.n254 GNDA.n253 76.3222
R3768 GNDA.n251 GNDA.n209 76.3222
R3769 GNDA.n247 GNDA.n246 76.3222
R3770 GNDA.n240 GNDA.n211 76.3222
R3771 GNDA.n239 GNDA.n238 76.3222
R3772 GNDA.n232 GNDA.n213 76.3222
R3773 GNDA.n1218 GNDA.n161 76.3222
R3774 GNDA.n1220 GNDA.n162 76.3222
R3775 GNDA.n1222 GNDA.n163 76.3222
R3776 GNDA.n1224 GNDA.n164 76.3222
R3777 GNDA.n2329 GNDA.n145 76.3222
R3778 GNDA.n1244 GNDA.n203 76.3222
R3779 GNDA.n1240 GNDA.n202 76.3222
R3780 GNDA.n1236 GNDA.n201 76.3222
R3781 GNDA.n1232 GNDA.n200 76.3222
R3782 GNDA.n1228 GNDA.n199 76.3222
R3783 GNDA.n2021 GNDA.n198 76.3222
R3784 GNDA.n1267 GNDA.n580 76.3222
R3785 GNDA.n1214 GNDA.n1213 76.3222
R3786 GNDA.n1261 GNDA.n1212 76.3222
R3787 GNDA.n1257 GNDA.n1211 76.3222
R3788 GNDA.n1253 GNDA.n1210 76.3222
R3789 GNDA.n1249 GNDA.n1209 76.3222
R3790 GNDA.n1905 GNDA.n1903 76.3222
R3791 GNDA.n1913 GNDA.n576 76.3222
R3792 GNDA.n1918 GNDA.n1915 76.3222
R3793 GNDA.n1916 GNDA.n570 76.3222
R3794 GNDA.n1929 GNDA.n567 76.3222
R3795 GNDA.n1387 GNDA.n1386 76.3222
R3796 GNDA.n1278 GNDA.n1277 76.3222
R3797 GNDA.n1376 GNDA.n1375 76.3222
R3798 GNDA.n1287 GNDA.n1286 76.3222
R3799 GNDA.n1365 GNDA.n1364 76.3222
R3800 GNDA.n1292 GNDA.n1291 76.3222
R3801 GNDA.n2298 GNDA.n2297 76.3222
R3802 GNDA.n259 GNDA.n191 76.3222
R3803 GNDA.n265 GNDA.n190 76.3222
R3804 GNDA.n271 GNDA.n189 76.3222
R3805 GNDA.n277 GNDA.n188 76.3222
R3806 GNDA.n2294 GNDA.n187 76.3222
R3807 GNDA.n684 GNDA.n683 76.3222
R3808 GNDA.n679 GNDA.n659 76.3222
R3809 GNDA.n676 GNDA.n658 76.3222
R3810 GNDA.n672 GNDA.n657 76.3222
R3811 GNDA.n668 GNDA.n656 76.3222
R3812 GNDA.n664 GNDA.n655 76.3222
R3813 GNDA.n633 GNDA.n632 76.3222
R3814 GNDA.n638 GNDA.n637 76.3222
R3815 GNDA.n641 GNDA.n640 76.3222
R3816 GNDA.n646 GNDA.n645 76.3222
R3817 GNDA.n649 GNDA.n648 76.3222
R3818 GNDA.n654 GNDA.n652 76.3222
R3819 GNDA.n1899 GNDA.n1898 76.3222
R3820 GNDA.n1908 GNDA.n1907 76.3222
R3821 GNDA.n1911 GNDA.n1910 76.3222
R3822 GNDA.n1921 GNDA.n1920 76.3222
R3823 GNDA.n1924 GNDA.n1923 76.3222
R3824 GNDA.n1813 GNDA.n572 76.3222
R3825 GNDA.n1874 GNDA.n1873 76.3222
R3826 GNDA.n1879 GNDA.n1878 76.3222
R3827 GNDA.n1882 GNDA.n1881 76.3222
R3828 GNDA.n1887 GNDA.n1886 76.3222
R3829 GNDA.n1890 GNDA.n1889 76.3222
R3830 GNDA.n1895 GNDA.n1894 76.3222
R3831 GNDA.n1852 GNDA.n1851 76.3222
R3832 GNDA.n1452 GNDA.n1451 76.3222
R3833 GNDA.n1485 GNDA.n1484 76.3222
R3834 GNDA.n1461 GNDA.n1460 76.3222
R3835 GNDA.n1474 GNDA.n1473 76.3222
R3836 GNDA.n1462 GNDA.n1394 76.3222
R3837 GNDA.n1547 GNDA.n1546 76.3222
R3838 GNDA.n1572 GNDA.n630 76.3222
R3839 GNDA.n1568 GNDA.n1567 76.3222
R3840 GNDA.n1561 GNDA.n635 76.3222
R3841 GNDA.n1560 GNDA.n1559 76.3222
R3842 GNDA.n1553 GNDA.n643 76.3222
R3843 GNDA.n1552 GNDA.n1551 76.3222
R3844 GNDA.n1597 GNDA.n1596 76.3222
R3845 GNDA.n1592 GNDA.n624 76.3222
R3846 GNDA.n1589 GNDA.n623 76.3222
R3847 GNDA.n1585 GNDA.n622 76.3222
R3848 GNDA.n1581 GNDA.n621 76.3222
R3849 GNDA.n1577 GNDA.n620 76.3222
R3850 GNDA.n1447 GNDA.n1415 76.3222
R3851 GNDA.n872 GNDA.n871 76.3222
R3852 GNDA.n758 GNDA.n757 76.3222
R3853 GNDA.n861 GNDA.n860 76.3222
R3854 GNDA.n767 GNDA.n766 76.3222
R3855 GNDA.n850 GNDA.n849 76.3222
R3856 GNDA.n777 GNDA.n772 76.3222
R3857 GNDA.n875 GNDA.n874 76.3222
R3858 GNDA.n924 GNDA.n923 76.3222
R3859 GNDA.n933 GNDA.n932 76.3222
R3860 GNDA.n936 GNDA.n935 76.3222
R3861 GNDA.n947 GNDA.n946 76.3222
R3862 GNDA.n950 GNDA.n949 76.3222
R3863 GNDA.n774 GNDA.n716 76.3222
R3864 GNDA.n989 GNDA.n686 76.3222
R3865 GNDA.n986 GNDA.n687 76.3222
R3866 GNDA.n976 GNDA.n688 76.3222
R3867 GNDA.n973 GNDA.n689 76.3222
R3868 GNDA.n694 GNDA.n690 76.3222
R3869 GNDA.n1207 GNDA.n1206 76.3222
R3870 GNDA.n928 GNDA.n927 76.3222
R3871 GNDA.n929 GNDA.n720 76.3222
R3872 GNDA.n940 GNDA.n939 76.3222
R3873 GNDA.n943 GNDA.n942 76.3222
R3874 GNDA.n953 GNDA.n713 76.3222
R3875 GNDA.n956 GNDA.n955 76.3222
R3876 GNDA.n2093 GNDA.n197 76.3222
R3877 GNDA.n1054 GNDA.n196 76.3222
R3878 GNDA.n1060 GNDA.n195 76.3222
R3879 GNDA.n1066 GNDA.n194 76.3222
R3880 GNDA.n1072 GNDA.n193 76.3222
R3881 GNDA.n1050 GNDA.n192 76.3222
R3882 GNDA.n1851 GNDA.n603 76.3222
R3883 GNDA.n1873 GNDA.n589 76.3222
R3884 GNDA.n1880 GNDA.n1879 76.3222
R3885 GNDA.n1881 GNDA.n587 76.3222
R3886 GNDA.n1888 GNDA.n1887 76.3222
R3887 GNDA.n1889 GNDA.n585 76.3222
R3888 GNDA.n1896 GNDA.n1895 76.3222
R3889 GNDA.n1597 GNDA.n625 76.3222
R3890 GNDA.n1590 GNDA.n624 76.3222
R3891 GNDA.n1586 GNDA.n623 76.3222
R3892 GNDA.n1582 GNDA.n622 76.3222
R3893 GNDA.n1578 GNDA.n621 76.3222
R3894 GNDA.n1574 GNDA.n620 76.3222
R3895 GNDA.n941 GNDA.n713 76.3222
R3896 GNDA.n944 GNDA.n943 76.3222
R3897 GNDA.n939 GNDA.n938 76.3222
R3898 GNDA.n930 GNDA.n929 76.3222
R3899 GNDA.n927 GNDA.n926 76.3222
R3900 GNDA.n648 GNDA.n647 76.3222
R3901 GNDA.n645 GNDA.n644 76.3222
R3902 GNDA.n640 GNDA.n639 76.3222
R3903 GNDA.n637 GNDA.n636 76.3222
R3904 GNDA.n632 GNDA.n631 76.3222
R3905 GNDA.n1928 GNDA.n1927 76.3222
R3906 GNDA.n1917 GNDA.n1916 76.3222
R3907 GNDA.n1915 GNDA.n1914 76.3222
R3908 GNDA.n1904 GNDA.n576 76.3222
R3909 GNDA.n1903 GNDA.n1902 76.3222
R3910 GNDA.n923 GNDA.n722 76.3222
R3911 GNDA.n934 GNDA.n933 76.3222
R3912 GNDA.n935 GNDA.n718 76.3222
R3913 GNDA.n948 GNDA.n947 76.3222
R3914 GNDA.n951 GNDA.n950 76.3222
R3915 GNDA.n1569 GNDA.n630 76.3222
R3916 GNDA.n1567 GNDA.n1566 76.3222
R3917 GNDA.n1562 GNDA.n1561 76.3222
R3918 GNDA.n1559 GNDA.n1558 76.3222
R3919 GNDA.n1554 GNDA.n1553 76.3222
R3920 GNDA.n1898 GNDA.n578 76.3222
R3921 GNDA.n1909 GNDA.n1908 76.3222
R3922 GNDA.n1910 GNDA.n574 76.3222
R3923 GNDA.n1922 GNDA.n1921 76.3222
R3924 GNDA.n1925 GNDA.n1924 76.3222
R3925 GNDA.n1814 GNDA.n1813 76.3222
R3926 GNDA.n1267 GNDA.n1266 76.3222
R3927 GNDA.n1262 GNDA.n1213 76.3222
R3928 GNDA.n1258 GNDA.n1212 76.3222
R3929 GNDA.n1254 GNDA.n1211 76.3222
R3930 GNDA.n1250 GNDA.n1210 76.3222
R3931 GNDA.n1246 GNDA.n1209 76.3222
R3932 GNDA.n684 GNDA.n660 76.3222
R3933 GNDA.n677 GNDA.n659 76.3222
R3934 GNDA.n673 GNDA.n658 76.3222
R3935 GNDA.n669 GNDA.n657 76.3222
R3936 GNDA.n665 GNDA.n656 76.3222
R3937 GNDA.n661 GNDA.n655 76.3222
R3938 GNDA.n2328 GNDA.n147 76.3222
R3939 GNDA.n1223 GNDA.n164 76.3222
R3940 GNDA.n1221 GNDA.n163 76.3222
R3941 GNDA.n1219 GNDA.n162 76.3222
R3942 GNDA.n1217 GNDA.n161 76.3222
R3943 GNDA.n1241 GNDA.n203 76.3222
R3944 GNDA.n1237 GNDA.n202 76.3222
R3945 GNDA.n1233 GNDA.n201 76.3222
R3946 GNDA.n1229 GNDA.n200 76.3222
R3947 GNDA.n1225 GNDA.n199 76.3222
R3948 GNDA.n2021 GNDA.n204 76.3222
R3949 GNDA.n1197 GNDA.n1196 76.3222
R3950 GNDA.n1085 GNDA.n1078 76.3222
R3951 GNDA.n1186 GNDA.n1185 76.3222
R3952 GNDA.n1094 GNDA.n1087 76.3222
R3953 GNDA.n1175 GNDA.n1174 76.3222
R3954 GNDA.n1100 GNDA.n1096 76.3222
R3955 GNDA.n2148 GNDA.n2147 76.3222
R3956 GNDA.n2095 GNDA.n155 76.3222
R3957 GNDA.n1052 GNDA.n156 76.3222
R3958 GNDA.n1058 GNDA.n157 76.3222
R3959 GNDA.n1064 GNDA.n158 76.3222
R3960 GNDA.n1070 GNDA.n159 76.3222
R3961 GNDA.n1200 GNDA.n154 76.3222
R3962 GNDA.n1199 GNDA.n159 76.3222
R3963 GNDA.n1069 GNDA.n158 76.3222
R3964 GNDA.n1063 GNDA.n157 76.3222
R3965 GNDA.n1057 GNDA.n156 76.3222
R3966 GNDA.n1051 GNDA.n155 76.3222
R3967 GNDA.n1053 GNDA.n197 76.3222
R3968 GNDA.n1059 GNDA.n196 76.3222
R3969 GNDA.n1065 GNDA.n195 76.3222
R3970 GNDA.n1071 GNDA.n194 76.3222
R3971 GNDA.n1074 GNDA.n193 76.3222
R3972 GNDA.n1076 GNDA.n154 76.3222
R3973 GNDA.n1101 GNDA.n1100 76.3222
R3974 GNDA.n1174 GNDA.n1173 76.3222
R3975 GNDA.n1095 GNDA.n1094 76.3222
R3976 GNDA.n1185 GNDA.n1184 76.3222
R3977 GNDA.n1086 GNDA.n1085 76.3222
R3978 GNDA.n1196 GNDA.n1195 76.3222
R3979 GNDA.n955 GNDA.n954 76.3222
R3980 GNDA.n1207 GNDA.n691 76.3222
R3981 GNDA.n972 GNDA.n690 76.3222
R3982 GNDA.n977 GNDA.n689 76.3222
R3983 GNDA.n985 GNDA.n688 76.3222
R3984 GNDA.n990 GNDA.n687 76.3222
R3985 GNDA.n957 GNDA.n686 76.3222
R3986 GNDA.n1050 GNDA.n205 76.3222
R3987 GNDA.n876 GNDA.n875 76.3222
R3988 GNDA.n772 GNDA.n768 76.3222
R3989 GNDA.n851 GNDA.n850 76.3222
R3990 GNDA.n766 GNDA.n759 76.3222
R3991 GNDA.n862 GNDA.n861 76.3222
R3992 GNDA.n757 GNDA.n749 76.3222
R3993 GNDA.n873 GNDA.n872 76.3222
R3994 GNDA.n775 GNDA.n774 76.3222
R3995 GNDA.n275 GNDA.n153 76.3222
R3996 GNDA.n274 GNDA.n152 76.3222
R3997 GNDA.n268 GNDA.n151 76.3222
R3998 GNDA.n262 GNDA.n150 76.3222
R3999 GNDA.n257 GNDA.n149 76.3222
R4000 GNDA.n2297 GNDA.n185 76.3222
R4001 GNDA.n264 GNDA.n191 76.3222
R4002 GNDA.n270 GNDA.n190 76.3222
R4003 GNDA.n276 GNDA.n189 76.3222
R4004 GNDA.n279 GNDA.n188 76.3222
R4005 GNDA.n2301 GNDA.n180 76.3222
R4006 GNDA.n2308 GNDA.n2307 76.3222
R4007 GNDA.n2309 GNDA.n178 76.3222
R4008 GNDA.n2316 GNDA.n2315 76.3222
R4009 GNDA.n2317 GNDA.n176 76.3222
R4010 GNDA.n2324 GNDA.n2323 76.3222
R4011 GNDA.n281 GNDA.n148 76.3222
R4012 GNDA.n652 GNDA.n651 76.3222
R4013 GNDA.n1291 GNDA.n1288 76.3222
R4014 GNDA.n1366 GNDA.n1365 76.3222
R4015 GNDA.n1286 GNDA.n1279 76.3222
R4016 GNDA.n1377 GNDA.n1376 76.3222
R4017 GNDA.n1277 GNDA.n1270 76.3222
R4018 GNDA.n1388 GNDA.n1387 76.3222
R4019 GNDA.n2295 GNDA.n2294 76.3222
R4020 GNDA.n1447 GNDA.n1446 76.3222
R4021 GNDA.n1546 GNDA.n1545 76.3222
R4022 GNDA.n1463 GNDA.n1462 76.3222
R4023 GNDA.n1475 GNDA.n1474 76.3222
R4024 GNDA.n1460 GNDA.n1453 76.3222
R4025 GNDA.n1486 GNDA.n1485 76.3222
R4026 GNDA.n1451 GNDA.n1450 76.3222
R4027 GNDA.n1551 GNDA.n1392 76.3222
R4028 GNDA.n305 GNDA.n301 76.3222
R4029 GNDA.n2265 GNDA.n2264 76.3222
R4030 GNDA.n299 GNDA.n292 76.3222
R4031 GNDA.n2276 GNDA.n2275 76.3222
R4032 GNDA.n290 GNDA.n283 76.3222
R4033 GNDA.n2287 GNDA.n2286 76.3222
R4034 GNDA.n253 GNDA.n252 76.3222
R4035 GNDA.n248 GNDA.n209 76.3222
R4036 GNDA.n246 GNDA.n245 76.3222
R4037 GNDA.n241 GNDA.n240 76.3222
R4038 GNDA.n238 GNDA.n237 76.3222
R4039 GNDA.n233 GNDA.n232 76.3222
R4040 GNDA.n2147 GNDA.n518 76.3222
R4041 GNDA.n2189 GNDA.n306 76.3222
R4042 GNDA.n109 GNDA.n91 76.3222
R4043 GNDA.n1506 GNDA.n1406 76.062
R4044 GNDA.n1507 GNDA.n1506 76.062
R4045 GNDA.n1327 GNDA.n1326 76.062
R4046 GNDA.n1326 GNDA.n1325 76.062
R4047 GNDA.n2226 GNDA.n2225 76.062
R4048 GNDA.n2225 GNDA.n2224 76.062
R4049 GNDA.n812 GNDA.n811 76.062
R4050 GNDA.n811 GNDA.n810 76.062
R4051 GNDA.n1012 GNDA.n1011 76.062
R4052 GNDA.n1011 GNDA.n1010 76.062
R4053 GNDA.n1136 GNDA.n1135 76.062
R4054 GNDA.n1135 GNDA.n1134 76.062
R4055 GNDA.n1775 GNDA.n1754 76.062
R4056 GNDA.n1776 GNDA.n1775 76.062
R4057 GNDA.n1984 GNDA.n1965 76.062
R4058 GNDA.n1985 GNDA.n1984 76.062
R4059 GNDA.n2371 GNDA.n2370 76.062
R4060 GNDA.n2370 GNDA.n2369 76.062
R4061 GNDA.t165 GNDA.t159 75.8626
R4062 GNDA.t23 GNDA.t31 75.8626
R4063 GNDA.t175 GNDA.t162 75.8626
R4064 GNDA.n1705 GNDA.t289 75.8626
R4065 GNDA.n1721 GNDA.t337 75.8626
R4066 GNDA.n1721 GNDA.t287 75.8626
R4067 GNDA.n1646 GNDA.t192 75.8626
R4068 GNDA.n1646 GNDA.t312 75.8626
R4069 GNDA.n1696 GNDA.t65 75.8626
R4070 GNDA.n1490 GNDA.n1489 74.5978
R4071 GNDA.n1491 GNDA.n1490 74.5978
R4072 GNDA.n1383 GNDA.n1272 74.5978
R4073 GNDA.n1310 GNDA.n1272 74.5978
R4074 GNDA.n2282 GNDA.n285 74.5978
R4075 GNDA.n2209 GNDA.n285 74.5978
R4076 GNDA.n868 GNDA.n752 74.5978
R4077 GNDA.n795 GNDA.n752 74.5978
R4078 GNDA.n994 GNDA.n993 74.5978
R4079 GNDA.n995 GNDA.n994 74.5978
R4080 GNDA.n1192 GNDA.n1080 74.5978
R4081 GNDA.n1119 GNDA.n1080 74.5978
R4082 GNDA.n1759 GNDA.n611 74.5978
R4083 GNDA.n1760 GNDA.n1759 74.5978
R4084 GNDA.n2054 GNDA.n1933 74.5978
R4085 GNDA.n1969 GNDA.n1933 74.5978
R4086 GNDA.n2353 GNDA.n2352 74.5978
R4087 GNDA.n2354 GNDA.n2353 74.5978
R4088 GNDA.n2435 GNDA.n93 73.3065
R4089 GNDA.n2465 GNDA.t64 72.3996
R4090 GNDA.n2451 GNDA.t325 72.3996
R4091 GNDA.n489 GNDA.t328 72.3996
R4092 GNDA.t188 GNDA.n327 72.3996
R4093 GNDA.t225 GNDA.n421 71.648
R4094 GNDA.n2459 GNDA.n62 70.0642
R4095 GNDA.n345 GNDA.n344 70.0642
R4096 GNDA.t43 GNDA.t286 69.5407
R4097 GNDA.t286 GNDA.t199 69.5407
R4098 GNDA.t267 GNDA.n1730 69.5407
R4099 GNDA.n1730 GNDA.t10 69.5407
R4100 GNDA.t14 GNDA.t210 69.5407
R4101 GNDA.t283 GNDA.t14 69.5407
R4102 GNDA.n1496 GNDA.t108 65.8183
R4103 GNDA.n1498 GNDA.t108 65.8183
R4104 GNDA.n1504 GNDA.t108 65.8183
R4105 GNDA.n1512 GNDA.t108 65.8183
R4106 GNDA.n1514 GNDA.t108 65.8183
R4107 GNDA.n1520 GNDA.t108 65.8183
R4108 GNDA.n1522 GNDA.t108 65.8183
R4109 GNDA.n1540 GNDA.t108 65.8183
R4110 GNDA.n1537 GNDA.t108 65.8183
R4111 GNDA.n1531 GNDA.t108 65.8183
R4112 GNDA.n1528 GNDA.t108 65.8183
R4113 GNDA.n1312 GNDA.t100 65.8183
R4114 GNDA.n1318 GNDA.t100 65.8183
R4115 GNDA.n1320 GNDA.t100 65.8183
R4116 GNDA.n1328 GNDA.t100 65.8183
R4117 GNDA.n1334 GNDA.t100 65.8183
R4118 GNDA.n1336 GNDA.t100 65.8183
R4119 GNDA.n1342 GNDA.t100 65.8183
R4120 GNDA.n1359 GNDA.t100 65.8183
R4121 GNDA.n1353 GNDA.t100 65.8183
R4122 GNDA.n1351 GNDA.t100 65.8183
R4123 GNDA.n1345 GNDA.t100 65.8183
R4124 GNDA.n2211 GNDA.t173 65.8183
R4125 GNDA.n2217 GNDA.t173 65.8183
R4126 GNDA.n2219 GNDA.t173 65.8183
R4127 GNDA.n2227 GNDA.t173 65.8183
R4128 GNDA.n2233 GNDA.t173 65.8183
R4129 GNDA.n2235 GNDA.t173 65.8183
R4130 GNDA.n2241 GNDA.t173 65.8183
R4131 GNDA.n2258 GNDA.t173 65.8183
R4132 GNDA.n2252 GNDA.t173 65.8183
R4133 GNDA.n2250 GNDA.t173 65.8183
R4134 GNDA.n2244 GNDA.t173 65.8183
R4135 GNDA.n797 GNDA.t126 65.8183
R4136 GNDA.n803 GNDA.t126 65.8183
R4137 GNDA.n805 GNDA.t126 65.8183
R4138 GNDA.n813 GNDA.t126 65.8183
R4139 GNDA.n819 GNDA.t126 65.8183
R4140 GNDA.n821 GNDA.t126 65.8183
R4141 GNDA.n827 GNDA.t126 65.8183
R4142 GNDA.n844 GNDA.t126 65.8183
R4143 GNDA.n838 GNDA.t126 65.8183
R4144 GNDA.n836 GNDA.t126 65.8183
R4145 GNDA.n830 GNDA.t126 65.8183
R4146 GNDA.n997 GNDA.t139 65.8183
R4147 GNDA.n1003 GNDA.t139 65.8183
R4148 GNDA.n1005 GNDA.t139 65.8183
R4149 GNDA.n1013 GNDA.t139 65.8183
R4150 GNDA.n1019 GNDA.t139 65.8183
R4151 GNDA.n1021 GNDA.t139 65.8183
R4152 GNDA.n1027 GNDA.t139 65.8183
R4153 GNDA.n1044 GNDA.t139 65.8183
R4154 GNDA.n1038 GNDA.t139 65.8183
R4155 GNDA.n1036 GNDA.t139 65.8183
R4156 GNDA.n1030 GNDA.t139 65.8183
R4157 GNDA.n1121 GNDA.t114 65.8183
R4158 GNDA.n1127 GNDA.t114 65.8183
R4159 GNDA.n1129 GNDA.t114 65.8183
R4160 GNDA.n1137 GNDA.t114 65.8183
R4161 GNDA.n1143 GNDA.t114 65.8183
R4162 GNDA.n1145 GNDA.t114 65.8183
R4163 GNDA.n1151 GNDA.t114 65.8183
R4164 GNDA.n1168 GNDA.t114 65.8183
R4165 GNDA.n1162 GNDA.t114 65.8183
R4166 GNDA.n1160 GNDA.t114 65.8183
R4167 GNDA.n1154 GNDA.t114 65.8183
R4168 GNDA.n1765 GNDA.t113 65.8183
R4169 GNDA.n1767 GNDA.t113 65.8183
R4170 GNDA.n1773 GNDA.t113 65.8183
R4171 GNDA.n1781 GNDA.t113 65.8183
R4172 GNDA.n1783 GNDA.t113 65.8183
R4173 GNDA.n1789 GNDA.t113 65.8183
R4174 GNDA.n1791 GNDA.t113 65.8183
R4175 GNDA.n1809 GNDA.t113 65.8183
R4176 GNDA.n1806 GNDA.t113 65.8183
R4177 GNDA.n1800 GNDA.t113 65.8183
R4178 GNDA.n1797 GNDA.t113 65.8183
R4179 GNDA.n1974 GNDA.t115 65.8183
R4180 GNDA.n1976 GNDA.t115 65.8183
R4181 GNDA.n1982 GNDA.t115 65.8183
R4182 GNDA.n1990 GNDA.t115 65.8183
R4183 GNDA.n1992 GNDA.t115 65.8183
R4184 GNDA.n1998 GNDA.t115 65.8183
R4185 GNDA.n2000 GNDA.t115 65.8183
R4186 GNDA.n2018 GNDA.t115 65.8183
R4187 GNDA.n2015 GNDA.t115 65.8183
R4188 GNDA.n2009 GNDA.t115 65.8183
R4189 GNDA.n2006 GNDA.t115 65.8183
R4190 GNDA.n2356 GNDA.t95 65.8183
R4191 GNDA.n2362 GNDA.t95 65.8183
R4192 GNDA.n2364 GNDA.t95 65.8183
R4193 GNDA.n2372 GNDA.t95 65.8183
R4194 GNDA.n2378 GNDA.t95 65.8183
R4195 GNDA.n2380 GNDA.t95 65.8183
R4196 GNDA.n2386 GNDA.t95 65.8183
R4197 GNDA.n2403 GNDA.t95 65.8183
R4198 GNDA.n2397 GNDA.t95 65.8183
R4199 GNDA.n2395 GNDA.t95 65.8183
R4200 GNDA.n2389 GNDA.t95 65.8183
R4201 GNDA.n2406 GNDA.t95 65.8183
R4202 GNDA.n2415 GNDA.t95 65.8183
R4203 GNDA.n2341 GNDA.t95 65.8183
R4204 GNDA.n2339 GNDA.t95 65.8183
R4205 GNDA.n1955 GNDA.t115 65.8183
R4206 GNDA.n2037 GNDA.t115 65.8183
R4207 GNDA.n1941 GNDA.t115 65.8183
R4208 GNDA.n2052 GNDA.t115 65.8183
R4209 GNDA.n1744 GNDA.t113 65.8183
R4210 GNDA.n1828 GNDA.t113 65.8183
R4211 GNDA.n1604 GNDA.t113 65.8183
R4212 GNDA.n1840 GNDA.t113 65.8183
R4213 GNDA.n1098 GNDA.t114 65.8183
R4214 GNDA.n1179 GNDA.t114 65.8183
R4215 GNDA.n1089 GNDA.t114 65.8183
R4216 GNDA.n1190 GNDA.t114 65.8183
R4217 GNDA.t139 GNDA.n696 65.8183
R4218 GNDA.n967 GNDA.t139 65.8183
R4219 GNDA.n981 GNDA.t139 65.8183
R4220 GNDA.n963 GNDA.t139 65.8183
R4221 GNDA.n770 GNDA.t126 65.8183
R4222 GNDA.n855 GNDA.t126 65.8183
R4223 GNDA.n761 GNDA.t126 65.8183
R4224 GNDA.n866 GNDA.t126 65.8183
R4225 GNDA.n303 GNDA.t173 65.8183
R4226 GNDA.n2269 GNDA.t173 65.8183
R4227 GNDA.n294 GNDA.t173 65.8183
R4228 GNDA.n2280 GNDA.t173 65.8183
R4229 GNDA.n1290 GNDA.t100 65.8183
R4230 GNDA.n1370 GNDA.t100 65.8183
R4231 GNDA.n1281 GNDA.t100 65.8183
R4232 GNDA.n1381 GNDA.t100 65.8183
R4233 GNDA.n1468 GNDA.t108 65.8183
R4234 GNDA.n1465 GNDA.t108 65.8183
R4235 GNDA.n1479 GNDA.t108 65.8183
R4236 GNDA.n1455 GNDA.t108 65.8183
R4237 GNDA.n101 GNDA.n81 65.6476
R4238 GNDA.t109 GNDA.n615 65.4161
R4239 GNDA.n2071 GNDA.t101 65.4161
R4240 GNDA.n2106 GNDA.t96 65.4161
R4241 GNDA.n450 GNDA.n373 64.0005
R4242 GNDA.n451 GNDA.n450 64.0005
R4243 GNDA.t223 GNDA.t207 63.2189
R4244 GNDA.t183 GNDA.t193 63.2189
R4245 GNDA.t6 GNDA.t57 63.2189
R4246 GNDA.t186 GNDA.t263 63.2189
R4247 GNDA.t287 GNDA.n1720 63.2189
R4248 GNDA.t192 GNDA.n1645 63.2189
R4249 GNDA.t109 GNDA.n582 60.9488
R4250 GNDA.t101 GNDA.n186 60.9488
R4251 GNDA.n454 GNDA.t324 60.7372
R4252 GNDA.t247 GNDA.n389 60.7372
R4253 GNDA.t87 GNDA.t219 59.0043
R4254 GNDA.t150 GNDA.t34 59.0043
R4255 GNDA.t168 GNDA.t288 56.897
R4256 GNDA.t265 GNDA.t216 56.897
R4257 GNDA.n1719 GNDA.t111 56.897
R4258 GNDA.n1644 GNDA.t128 56.897
R4259 GNDA.t310 GNDA.t275 56.897
R4260 GNDA.t141 GNDA.t203 56.897
R4261 GNDA.n516 GNDA.n171 55.2535
R4262 GNDA.n2188 GNDA.n168 55.2535
R4263 GNDA.n2436 GNDA.n92 55.2535
R4264 GNDA.n2353 GNDA.t95 55.2026
R4265 GNDA.t115 GNDA.n1933 55.2026
R4266 GNDA.n1759 GNDA.t113 55.2026
R4267 GNDA.t114 GNDA.n1080 55.2026
R4268 GNDA.n994 GNDA.t139 55.2026
R4269 GNDA.t126 GNDA.n752 55.2026
R4270 GNDA.t173 GNDA.n285 55.2026
R4271 GNDA.t100 GNDA.n1272 55.2026
R4272 GNDA.n1490 GNDA.t108 55.2026
R4273 GNDA.t70 GNDA.n361 54.7898
R4274 GNDA.n2473 GNDA.t16 54.7898
R4275 GNDA.n1506 GNDA.t108 54.4705
R4276 GNDA.n1326 GNDA.t100 54.4705
R4277 GNDA.n2225 GNDA.t173 54.4705
R4278 GNDA.n811 GNDA.t126 54.4705
R4279 GNDA.n1011 GNDA.t139 54.4705
R4280 GNDA.n1135 GNDA.t114 54.4705
R4281 GNDA.n1775 GNDA.t113 54.4705
R4282 GNDA.n1984 GNDA.t115 54.4705
R4283 GNDA.n2370 GNDA.t95 54.4705
R4284 GNDA.n418 GNDA.n417 54.4005
R4285 GNDA.n1481 GNDA.n1455 53.3664
R4286 GNDA.n1479 GNDA.n1478 53.3664
R4287 GNDA.n1470 GNDA.n1465 53.3664
R4288 GNDA.n1468 GNDA.n1397 53.3664
R4289 GNDA.n1528 GNDA.n1527 53.3664
R4290 GNDA.n1532 GNDA.n1531 53.3664
R4291 GNDA.n1537 GNDA.n1536 53.3664
R4292 GNDA.n1540 GNDA.n1539 53.3664
R4293 GNDA.n1512 GNDA.n1511 53.3664
R4294 GNDA.n1515 GNDA.n1514 53.3664
R4295 GNDA.n1520 GNDA.n1519 53.3664
R4296 GNDA.n1523 GNDA.n1522 53.3664
R4297 GNDA.n1505 GNDA.n1504 53.3664
R4298 GNDA.n1498 GNDA.n1408 53.3664
R4299 GNDA.n1497 GNDA.n1496 53.3664
R4300 GNDA.n1496 GNDA.n1495 53.3664
R4301 GNDA.n1499 GNDA.n1498 53.3664
R4302 GNDA.n1504 GNDA.n1503 53.3664
R4303 GNDA.n1513 GNDA.n1512 53.3664
R4304 GNDA.n1514 GNDA.n1404 53.3664
R4305 GNDA.n1521 GNDA.n1520 53.3664
R4306 GNDA.n1522 GNDA.n1402 53.3664
R4307 GNDA.n1541 GNDA.n1540 53.3664
R4308 GNDA.n1538 GNDA.n1537 53.3664
R4309 GNDA.n1531 GNDA.n1399 53.3664
R4310 GNDA.n1529 GNDA.n1528 53.3664
R4311 GNDA.n1381 GNDA.n1380 53.3664
R4312 GNDA.n1372 GNDA.n1281 53.3664
R4313 GNDA.n1370 GNDA.n1369 53.3664
R4314 GNDA.n1361 GNDA.n1290 53.3664
R4315 GNDA.n1345 GNDA.n1344 53.3664
R4316 GNDA.n1351 GNDA.n1350 53.3664
R4317 GNDA.n1354 GNDA.n1353 53.3664
R4318 GNDA.n1359 GNDA.n1358 53.3664
R4319 GNDA.n1329 GNDA.n1328 53.3664
R4320 GNDA.n1334 GNDA.n1333 53.3664
R4321 GNDA.n1337 GNDA.n1336 53.3664
R4322 GNDA.n1342 GNDA.n1341 53.3664
R4323 GNDA.n1320 GNDA.n1305 53.3664
R4324 GNDA.n1319 GNDA.n1318 53.3664
R4325 GNDA.n1312 GNDA.n1307 53.3664
R4326 GNDA.n1313 GNDA.n1312 53.3664
R4327 GNDA.n1318 GNDA.n1317 53.3664
R4328 GNDA.n1321 GNDA.n1320 53.3664
R4329 GNDA.n1328 GNDA.n1303 53.3664
R4330 GNDA.n1335 GNDA.n1334 53.3664
R4331 GNDA.n1336 GNDA.n1301 53.3664
R4332 GNDA.n1343 GNDA.n1342 53.3664
R4333 GNDA.n1360 GNDA.n1359 53.3664
R4334 GNDA.n1353 GNDA.n1296 53.3664
R4335 GNDA.n1352 GNDA.n1351 53.3664
R4336 GNDA.n1346 GNDA.n1345 53.3664
R4337 GNDA.n2280 GNDA.n2279 53.3664
R4338 GNDA.n2271 GNDA.n294 53.3664
R4339 GNDA.n2269 GNDA.n2268 53.3664
R4340 GNDA.n2260 GNDA.n303 53.3664
R4341 GNDA.n2244 GNDA.n2243 53.3664
R4342 GNDA.n2250 GNDA.n2249 53.3664
R4343 GNDA.n2253 GNDA.n2252 53.3664
R4344 GNDA.n2258 GNDA.n2257 53.3664
R4345 GNDA.n2228 GNDA.n2227 53.3664
R4346 GNDA.n2233 GNDA.n2232 53.3664
R4347 GNDA.n2236 GNDA.n2235 53.3664
R4348 GNDA.n2241 GNDA.n2240 53.3664
R4349 GNDA.n2219 GNDA.n2204 53.3664
R4350 GNDA.n2218 GNDA.n2217 53.3664
R4351 GNDA.n2211 GNDA.n2206 53.3664
R4352 GNDA.n2212 GNDA.n2211 53.3664
R4353 GNDA.n2217 GNDA.n2216 53.3664
R4354 GNDA.n2220 GNDA.n2219 53.3664
R4355 GNDA.n2227 GNDA.n2202 53.3664
R4356 GNDA.n2234 GNDA.n2233 53.3664
R4357 GNDA.n2235 GNDA.n2200 53.3664
R4358 GNDA.n2242 GNDA.n2241 53.3664
R4359 GNDA.n2259 GNDA.n2258 53.3664
R4360 GNDA.n2252 GNDA.n2195 53.3664
R4361 GNDA.n2251 GNDA.n2250 53.3664
R4362 GNDA.n2245 GNDA.n2244 53.3664
R4363 GNDA.n866 GNDA.n865 53.3664
R4364 GNDA.n857 GNDA.n761 53.3664
R4365 GNDA.n855 GNDA.n854 53.3664
R4366 GNDA.n846 GNDA.n770 53.3664
R4367 GNDA.n830 GNDA.n829 53.3664
R4368 GNDA.n836 GNDA.n835 53.3664
R4369 GNDA.n839 GNDA.n838 53.3664
R4370 GNDA.n844 GNDA.n843 53.3664
R4371 GNDA.n814 GNDA.n813 53.3664
R4372 GNDA.n819 GNDA.n818 53.3664
R4373 GNDA.n822 GNDA.n821 53.3664
R4374 GNDA.n827 GNDA.n826 53.3664
R4375 GNDA.n805 GNDA.n790 53.3664
R4376 GNDA.n804 GNDA.n803 53.3664
R4377 GNDA.n797 GNDA.n792 53.3664
R4378 GNDA.n798 GNDA.n797 53.3664
R4379 GNDA.n803 GNDA.n802 53.3664
R4380 GNDA.n806 GNDA.n805 53.3664
R4381 GNDA.n813 GNDA.n788 53.3664
R4382 GNDA.n820 GNDA.n819 53.3664
R4383 GNDA.n821 GNDA.n786 53.3664
R4384 GNDA.n828 GNDA.n827 53.3664
R4385 GNDA.n845 GNDA.n844 53.3664
R4386 GNDA.n838 GNDA.n781 53.3664
R4387 GNDA.n837 GNDA.n836 53.3664
R4388 GNDA.n831 GNDA.n830 53.3664
R4389 GNDA.n964 GNDA.n963 53.3664
R4390 GNDA.n981 GNDA.n980 53.3664
R4391 GNDA.n968 GNDA.n967 53.3664
R4392 GNDA.n1046 GNDA.n696 53.3664
R4393 GNDA.n1030 GNDA.n1029 53.3664
R4394 GNDA.n1036 GNDA.n1035 53.3664
R4395 GNDA.n1039 GNDA.n1038 53.3664
R4396 GNDA.n1044 GNDA.n1043 53.3664
R4397 GNDA.n1014 GNDA.n1013 53.3664
R4398 GNDA.n1019 GNDA.n1018 53.3664
R4399 GNDA.n1022 GNDA.n1021 53.3664
R4400 GNDA.n1027 GNDA.n1026 53.3664
R4401 GNDA.n1005 GNDA.n706 53.3664
R4402 GNDA.n1004 GNDA.n1003 53.3664
R4403 GNDA.n997 GNDA.n708 53.3664
R4404 GNDA.n998 GNDA.n997 53.3664
R4405 GNDA.n1003 GNDA.n1002 53.3664
R4406 GNDA.n1006 GNDA.n1005 53.3664
R4407 GNDA.n1013 GNDA.n704 53.3664
R4408 GNDA.n1020 GNDA.n1019 53.3664
R4409 GNDA.n1021 GNDA.n702 53.3664
R4410 GNDA.n1028 GNDA.n1027 53.3664
R4411 GNDA.n1045 GNDA.n1044 53.3664
R4412 GNDA.n1038 GNDA.n697 53.3664
R4413 GNDA.n1037 GNDA.n1036 53.3664
R4414 GNDA.n1031 GNDA.n1030 53.3664
R4415 GNDA.n1190 GNDA.n1189 53.3664
R4416 GNDA.n1181 GNDA.n1089 53.3664
R4417 GNDA.n1179 GNDA.n1178 53.3664
R4418 GNDA.n1170 GNDA.n1098 53.3664
R4419 GNDA.n1154 GNDA.n1153 53.3664
R4420 GNDA.n1160 GNDA.n1159 53.3664
R4421 GNDA.n1163 GNDA.n1162 53.3664
R4422 GNDA.n1168 GNDA.n1167 53.3664
R4423 GNDA.n1138 GNDA.n1137 53.3664
R4424 GNDA.n1143 GNDA.n1142 53.3664
R4425 GNDA.n1146 GNDA.n1145 53.3664
R4426 GNDA.n1151 GNDA.n1150 53.3664
R4427 GNDA.n1129 GNDA.n1114 53.3664
R4428 GNDA.n1128 GNDA.n1127 53.3664
R4429 GNDA.n1121 GNDA.n1116 53.3664
R4430 GNDA.n1122 GNDA.n1121 53.3664
R4431 GNDA.n1127 GNDA.n1126 53.3664
R4432 GNDA.n1130 GNDA.n1129 53.3664
R4433 GNDA.n1137 GNDA.n1112 53.3664
R4434 GNDA.n1144 GNDA.n1143 53.3664
R4435 GNDA.n1145 GNDA.n1110 53.3664
R4436 GNDA.n1152 GNDA.n1151 53.3664
R4437 GNDA.n1169 GNDA.n1168 53.3664
R4438 GNDA.n1162 GNDA.n1105 53.3664
R4439 GNDA.n1161 GNDA.n1160 53.3664
R4440 GNDA.n1155 GNDA.n1154 53.3664
R4441 GNDA.n1840 GNDA.n1839 53.3664
R4442 GNDA.n1605 GNDA.n1604 53.3664
R4443 GNDA.n1828 GNDA.n1827 53.3664
R4444 GNDA.n1745 GNDA.n1744 53.3664
R4445 GNDA.n1797 GNDA.n1796 53.3664
R4446 GNDA.n1801 GNDA.n1800 53.3664
R4447 GNDA.n1806 GNDA.n1805 53.3664
R4448 GNDA.n1809 GNDA.n1808 53.3664
R4449 GNDA.n1781 GNDA.n1780 53.3664
R4450 GNDA.n1784 GNDA.n1783 53.3664
R4451 GNDA.n1789 GNDA.n1788 53.3664
R4452 GNDA.n1792 GNDA.n1791 53.3664
R4453 GNDA.n1774 GNDA.n1773 53.3664
R4454 GNDA.n1767 GNDA.n1756 53.3664
R4455 GNDA.n1766 GNDA.n1765 53.3664
R4456 GNDA.n1765 GNDA.n1764 53.3664
R4457 GNDA.n1768 GNDA.n1767 53.3664
R4458 GNDA.n1773 GNDA.n1772 53.3664
R4459 GNDA.n1782 GNDA.n1781 53.3664
R4460 GNDA.n1783 GNDA.n1752 53.3664
R4461 GNDA.n1790 GNDA.n1789 53.3664
R4462 GNDA.n1791 GNDA.n1750 53.3664
R4463 GNDA.n1810 GNDA.n1809 53.3664
R4464 GNDA.n1807 GNDA.n1806 53.3664
R4465 GNDA.n1800 GNDA.n1747 53.3664
R4466 GNDA.n1798 GNDA.n1797 53.3664
R4467 GNDA.n2052 GNDA.n2051 53.3664
R4468 GNDA.n2039 GNDA.n1941 53.3664
R4469 GNDA.n2037 GNDA.n2036 53.3664
R4470 GNDA.n1956 GNDA.n1955 53.3664
R4471 GNDA.n2006 GNDA.n2005 53.3664
R4472 GNDA.n2010 GNDA.n2009 53.3664
R4473 GNDA.n2015 GNDA.n2014 53.3664
R4474 GNDA.n2018 GNDA.n2017 53.3664
R4475 GNDA.n1990 GNDA.n1989 53.3664
R4476 GNDA.n1993 GNDA.n1992 53.3664
R4477 GNDA.n1998 GNDA.n1997 53.3664
R4478 GNDA.n2001 GNDA.n2000 53.3664
R4479 GNDA.n1983 GNDA.n1982 53.3664
R4480 GNDA.n1976 GNDA.n1967 53.3664
R4481 GNDA.n1975 GNDA.n1974 53.3664
R4482 GNDA.n1974 GNDA.n1973 53.3664
R4483 GNDA.n1977 GNDA.n1976 53.3664
R4484 GNDA.n1982 GNDA.n1981 53.3664
R4485 GNDA.n1991 GNDA.n1990 53.3664
R4486 GNDA.n1992 GNDA.n1963 53.3664
R4487 GNDA.n1999 GNDA.n1998 53.3664
R4488 GNDA.n2000 GNDA.n1961 53.3664
R4489 GNDA.n2019 GNDA.n2018 53.3664
R4490 GNDA.n2016 GNDA.n2015 53.3664
R4491 GNDA.n2009 GNDA.n1958 53.3664
R4492 GNDA.n2007 GNDA.n2006 53.3664
R4493 GNDA.n2340 GNDA.n2339 53.3664
R4494 GNDA.n2341 GNDA.n124 53.3664
R4495 GNDA.n2415 GNDA.n2414 53.3664
R4496 GNDA.n2406 GNDA.n2405 53.3664
R4497 GNDA.n2389 GNDA.n2388 53.3664
R4498 GNDA.n2395 GNDA.n2394 53.3664
R4499 GNDA.n2398 GNDA.n2397 53.3664
R4500 GNDA.n2403 GNDA.n2402 53.3664
R4501 GNDA.n2373 GNDA.n2372 53.3664
R4502 GNDA.n2378 GNDA.n2377 53.3664
R4503 GNDA.n2381 GNDA.n2380 53.3664
R4504 GNDA.n2386 GNDA.n2385 53.3664
R4505 GNDA.n2364 GNDA.n134 53.3664
R4506 GNDA.n2363 GNDA.n2362 53.3664
R4507 GNDA.n2356 GNDA.n136 53.3664
R4508 GNDA.n2357 GNDA.n2356 53.3664
R4509 GNDA.n2362 GNDA.n2361 53.3664
R4510 GNDA.n2365 GNDA.n2364 53.3664
R4511 GNDA.n2372 GNDA.n132 53.3664
R4512 GNDA.n2379 GNDA.n2378 53.3664
R4513 GNDA.n2380 GNDA.n130 53.3664
R4514 GNDA.n2387 GNDA.n2386 53.3664
R4515 GNDA.n2404 GNDA.n2403 53.3664
R4516 GNDA.n2397 GNDA.n125 53.3664
R4517 GNDA.n2396 GNDA.n2395 53.3664
R4518 GNDA.n2390 GNDA.n2389 53.3664
R4519 GNDA.n2407 GNDA.n2406 53.3664
R4520 GNDA.n2416 GNDA.n2415 53.3664
R4521 GNDA.n2342 GNDA.n2341 53.3664
R4522 GNDA.n2339 GNDA.n139 53.3664
R4523 GNDA.n1955 GNDA.n1943 53.3664
R4524 GNDA.n2038 GNDA.n2037 53.3664
R4525 GNDA.n1941 GNDA.n1935 53.3664
R4526 GNDA.n2053 GNDA.n2052 53.3664
R4527 GNDA.n1744 GNDA.n1606 53.3664
R4528 GNDA.n1829 GNDA.n1828 53.3664
R4529 GNDA.n1604 GNDA.n612 53.3664
R4530 GNDA.n1841 GNDA.n1840 53.3664
R4531 GNDA.n1098 GNDA.n1091 53.3664
R4532 GNDA.n1180 GNDA.n1179 53.3664
R4533 GNDA.n1089 GNDA.n1082 53.3664
R4534 GNDA.n1191 GNDA.n1190 53.3664
R4535 GNDA.n969 GNDA.n696 53.3664
R4536 GNDA.n967 GNDA.n965 53.3664
R4537 GNDA.n982 GNDA.n981 53.3664
R4538 GNDA.n963 GNDA.n711 53.3664
R4539 GNDA.n770 GNDA.n763 53.3664
R4540 GNDA.n856 GNDA.n855 53.3664
R4541 GNDA.n761 GNDA.n754 53.3664
R4542 GNDA.n867 GNDA.n866 53.3664
R4543 GNDA.n303 GNDA.n296 53.3664
R4544 GNDA.n2270 GNDA.n2269 53.3664
R4545 GNDA.n294 GNDA.n287 53.3664
R4546 GNDA.n2281 GNDA.n2280 53.3664
R4547 GNDA.n1290 GNDA.n1283 53.3664
R4548 GNDA.n1371 GNDA.n1370 53.3664
R4549 GNDA.n1281 GNDA.n1274 53.3664
R4550 GNDA.n1382 GNDA.n1381 53.3664
R4551 GNDA.n1469 GNDA.n1468 53.3664
R4552 GNDA.n1465 GNDA.n1457 53.3664
R4553 GNDA.n1480 GNDA.n1479 53.3664
R4554 GNDA.n1455 GNDA.n1412 53.3664
R4555 GNDA.n2125 GNDA.n2122 52.5182
R4556 GNDA.n2326 GNDA.n172 52.5182
R4557 GNDA.n229 GNDA.n215 52.5182
R4558 GNDA.n373 GNDA.n372 51.2005
R4559 GNDA.n452 GNDA.n451 51.2005
R4560 GNDA.n482 GNDA.n327 50.5752
R4561 GNDA.n2466 GNDA.n2465 50.5752
R4562 GNDA.n2131 GNDA.n525 49.2359
R4563 GNDA.n2132 GNDA.n2131 49.2359
R4564 GNDA.n2134 GNDA.n2132 49.2359
R4565 GNDA.n2134 GNDA.n2133 49.2359
R4566 GNDA.n2141 GNDA.n2140 49.2359
R4567 GNDA.n2142 GNDA.n2141 49.2359
R4568 GNDA.n2142 GNDA.n513 49.2359
R4569 GNDA.n2149 GNDA.n516 49.2359
R4570 GNDA.n498 GNDA.n172 49.2359
R4571 GNDA.n504 GNDA.n498 49.2359
R4572 GNDA.n2160 GNDA.n2158 49.2359
R4573 GNDA.n2160 GNDA.n2159 49.2359
R4574 GNDA.n2184 GNDA.n2183 49.2359
R4575 GNDA.n2188 GNDA.n2187 49.2359
R4576 GNDA.n229 GNDA.n228 49.2359
R4577 GNDA.n228 GNDA.n227 49.2359
R4578 GNDA.n227 GNDA.n218 49.2359
R4579 GNDA.n221 GNDA.n218 49.2359
R4580 GNDA.n221 GNDA.n116 49.2359
R4581 GNDA.n2421 GNDA.n103 49.2359
R4582 GNDA.n2428 GNDA.n107 49.2359
R4583 GNDA.n110 GNDA.n107 49.2359
R4584 GNDA.n110 GNDA.n92 49.2359
R4585 GNDA.n77 GNDA.t25 49.0451
R4586 GNDA.t333 GNDA.n341 49.0451
R4587 GNDA.t96 GNDA.n2326 47.5947
R4588 GNDA.n2169 GNDA.n2168 47.5947
R4589 GNDA.t96 GNDA.n171 47.0476
R4590 GNDA.t96 GNDA.n168 47.0476
R4591 GNDA.t74 GNDA.t77 46.3607
R4592 GNDA.t339 GNDA.t74 46.3607
R4593 GNDA.n440 GNDA.t201 46.3607
R4594 GNDA.t279 GNDA.t271 46.3607
R4595 GNDA.t227 GNDA.t279 46.3607
R4596 GNDA.n348 GNDA.n339 44.8005
R4597 GNDA.n2456 GNDA.n2455 44.8005
R4598 GNDA.t235 GNDA.t51 44.2534
R4599 GNDA.t311 GNDA.t197 44.2534
R4600 GNDA.n119 GNDA.n117 43.0993
R4601 GNDA.t131 GNDA.t319 42.1461
R4602 GNDA.t226 GNDA.t68 42.1461
R4603 GNDA.t79 GNDA.t313 42.1461
R4604 GNDA.t184 GNDA.t195 42.1461
R4605 GNDA.t71 GNDA.t180 42.1461
R4606 GNDA.t3 GNDA.t18 42.1461
R4607 GNDA.t187 GNDA.t54 42.1461
R4608 GNDA.t84 GNDA.t231 42.1461
R4609 GNDA.t315 GNDA.t156 42.1461
R4610 GNDA.t47 GNDA.t249 42.1461
R4611 GNDA.t4 GNDA.t237 42.1461
R4612 GNDA.t181 GNDA.t53 42.1461
R4613 GNDA.t261 GNDA.t334 42.1461
R4614 GNDA.t60 GNDA.t259 42.1461
R4615 GNDA.t62 GNDA.t66 42.1461
R4616 GNDA.t45 GNDA.t177 42.1461
R4617 GNDA.t117 GNDA.t260 42.1461
R4618 GNDA.n2157 GNDA.n504 42.1241
R4619 GNDA.t24 GNDA.n2458 39.7033
R4620 GNDA.n346 GNDA.t20 39.7033
R4621 GNDA.n361 GNDA.t339 37.9315
R4622 GNDA.n390 GNDA.t56 37.9315
R4623 GNDA.t212 GNDA.t221 37.9315
R4624 GNDA.n2473 GNDA.t271 37.9315
R4625 GNDA.n2184 GNDA.n307 36.6535
R4626 GNDA.n24 GNDA.n23 34.813
R4627 GNDA.n2491 GNDA.n12 34.813
R4628 GNDA.n2122 GNDA.n490 33.9182
R4629 GNDA.n471 GNDA.n362 33.717
R4630 GNDA.t241 GNDA.t131 33.717
R4631 GNDA.t321 GNDA.t243 33.717
R4632 GNDA.t68 GNDA.t248 33.717
R4633 GNDA.t313 GNDA.t246 33.717
R4634 GNDA.t195 GNDA.t240 33.717
R4635 GNDA.t245 GNDA.t71 33.717
R4636 GNDA.t18 GNDA.t239 33.717
R4637 GNDA.t54 GNDA.t244 33.717
R4638 GNDA.t231 GNDA.t87 33.717
R4639 GNDA.t150 GNDA.t315 33.717
R4640 GNDA.t204 GNDA.t4 33.717
R4641 GNDA.t37 GNDA.t181 33.717
R4642 GNDA.t26 GNDA.t261 33.717
R4643 GNDA.t234 GNDA.t60 33.717
R4644 GNDA.t236 GNDA.t62 33.717
R4645 GNDA.t329 GNDA.t45 33.717
R4646 GNDA.t206 GNDA.t117 33.717
R4647 GNDA.n457 GNDA.n456 33.717
R4648 GNDA.t289 GNDA.t41 31.6097
R4649 GNDA.t252 GNDA.t320 31.6097
R4650 GNDA.t1 GNDA.t214 31.6097
R4651 GNDA.t49 GNDA.t65 31.6097
R4652 GNDA.n2125 GNDA.n2124 31.1829
R4653 GNDA.n2182 GNDA.n311 31.1829
R4654 GNDA.n215 GNDA.n167 31.1829
R4655 GNDA.t109 GNDA.n616 31.0997
R4656 GNDA.n531 GNDA.t96 31.0997
R4657 GNDA.n64 GNDA.t64 30.3614
R4658 GNDA.n75 GNDA.t331 30.3614
R4659 GNDA.t78 GNDA.n342 30.3614
R4660 GNDA.n352 GNDA.t188 30.3614
R4661 GNDA.t255 GNDA.t223 29.5024
R4662 GNDA.t193 GNDA.t70 29.5024
R4663 GNDA.n2486 GNDA.t47 29.5024
R4664 GNDA.t57 GNDA.t16 29.5024
R4665 GNDA.t263 GNDA.t8 29.5024
R4666 GNDA.n468 GNDA.n467 29.3193
R4667 GNDA.n485 GNDA.n484 28.413
R4668 GNDA.n2468 GNDA.n50 28.413
R4669 GNDA.n2171 GNDA.n98 28.1318
R4670 GNDA.n479 GNDA.n356 28.038
R4671 GNDA.n60 GNDA.n39 28.038
R4672 GNDA.n1726 GNDA.n1622 27.8193
R4673 GNDA.n1724 GNDA.n1723 27.8193
R4674 GNDA.n1509 GNDA.n1508 27.5561
R4675 GNDA.n1324 GNDA.n1304 27.5561
R4676 GNDA.n2223 GNDA.n2203 27.5561
R4677 GNDA.n809 GNDA.n789 27.5561
R4678 GNDA.n1009 GNDA.n705 27.5561
R4679 GNDA.n1133 GNDA.n1113 27.5561
R4680 GNDA.n1778 GNDA.n1777 27.5561
R4681 GNDA.n1987 GNDA.n1986 27.5561
R4682 GNDA.n2368 GNDA.n133 27.5561
R4683 GNDA.n582 GNDA.n563 26.9584
R4684 GNDA.n2296 GNDA.n186 26.9584
R4685 GNDA.n2133 GNDA.t96 25.7123
R4686 GNDA.n2159 GNDA.t96 25.7123
R4687 GNDA.t96 GNDA.n116 25.7123
R4688 GNDA.t25 GNDA.n75 25.6905
R4689 GNDA.n342 GNDA.t333 25.6905
R4690 GNDA.n359 GNDA.n358 25.6005
R4691 GNDA.n2471 GNDA.n2470 25.6005
R4692 GNDA.n1707 GNDA.n1705 25.2879
R4693 GNDA.n1696 GNDA.n1641 25.2879
R4694 GNDA.n1671 GNDA.t211 24.0005
R4695 GNDA.n1671 GNDA.t284 24.0005
R4696 GNDA.n1669 GNDA.t198 24.0005
R4697 GNDA.n1669 GNDA.t276 24.0005
R4698 GNDA.n1667 GNDA.t215 24.0005
R4699 GNDA.n1667 GNDA.t50 24.0005
R4700 GNDA.n1665 GNDA.t270 24.0005
R4701 GNDA.n1665 GNDA.t13 24.0005
R4702 GNDA.n1663 GNDA.t11 24.0005
R4703 GNDA.n1663 GNDA.t251 24.0005
R4704 GNDA.n1661 GNDA.t209 24.0005
R4705 GNDA.n1661 GNDA.t268 24.0005
R4706 GNDA.n1659 GNDA.t278 24.0005
R4707 GNDA.n1659 GNDA.t274 24.0005
R4708 GNDA.n1657 GNDA.t42 24.0005
R4709 GNDA.n1657 GNDA.t253 24.0005
R4710 GNDA.n1655 GNDA.t217 24.0005
R4711 GNDA.n1655 GNDA.t52 24.0005
R4712 GNDA.n1654 GNDA.t44 24.0005
R4713 GNDA.n1654 GNDA.t200 24.0005
R4714 GNDA.n1526 GNDA.n1525 23.6449
R4715 GNDA.n1300 GNDA.n1299 23.6449
R4716 GNDA.n2199 GNDA.n2198 23.6449
R4717 GNDA.n785 GNDA.n784 23.6449
R4718 GNDA.n701 GNDA.n700 23.6449
R4719 GNDA.n1109 GNDA.n1108 23.6449
R4720 GNDA.n1795 GNDA.n1794 23.6449
R4721 GNDA.n2004 GNDA.n2003 23.6449
R4722 GNDA.n129 GNDA.n128 23.6449
R4723 GNDA.n2140 GNDA.t96 23.5241
R4724 GNDA.n2168 GNDA.t96 23.5241
R4725 GNDA.n2421 GNDA.t96 23.5241
R4726 GNDA.n356 GNDA.n355 22.4005
R4727 GNDA.n418 GNDA.n416 22.4005
R4728 GNDA.n2482 GNDA.n2481 22.4005
R4729 GNDA.n2463 GNDA.n60 22.4005
R4730 GNDA.t238 GNDA.t29 21.8829
R4731 GNDA.n554 GNDA.n493 21.4917
R4732 GNDA.n2079 GNDA.t101 21.4482
R4733 GNDA.n1652 GNDA.n1649 21.3338
R4734 GNDA.n1651 GNDA.n1650 21.3338
R4735 GNDA.n1727 GNDA.n1621 21.3338
R4736 GNDA.n1620 GNDA.n1619 21.3338
R4737 GNDA.n1624 GNDA.n1623 21.3338
R4738 GNDA.n1709 GNDA.n1708 21.3338
R4739 GNDA.n444 GNDA.n443 21.3338
R4740 GNDA.n377 GNDA.n376 21.3338
R4741 GNDA.n381 GNDA.n380 21.3338
R4742 GNDA.n382 GNDA.n379 21.3338
R4743 GNDA.n437 GNDA.n435 21.3338
R4744 GNDA.n434 GNDA.n432 21.3338
R4745 GNDA.n373 GNDA.n370 21.3338
R4746 GNDA.n372 GNDA.n371 21.3338
R4747 GNDA.n366 GNDA.n365 21.3338
R4748 GNDA.n453 GNDA.n367 21.3338
R4749 GNDA.n452 GNDA.n368 21.3338
R4750 GNDA.n451 GNDA.n369 21.3338
R4751 GNDA.n464 GNDA.n462 21.3338
R4752 GNDA.n323 GNDA.n322 21.3338
R4753 GNDA.n360 GNDA.n357 21.3338
R4754 GNDA.n331 GNDA.n330 21.3338
R4755 GNDA.n49 GNDA.n48 21.3338
R4756 GNDA.n52 GNDA.n51 21.3338
R4757 GNDA.n45 GNDA.n44 21.3338
R4758 GNDA.n43 GNDA.n42 21.3338
R4759 GNDA.n1677 GNDA.n1674 21.1792
R4760 GNDA.n339 GNDA.n319 20.6005
R4761 GNDA.n2455 GNDA.n2454 20.6005
R4762 GNDA.n2493 GNDA.n0 19.9817
R4763 GNDA.n22 GNDA.t17 19.7005
R4764 GNDA.n22 GNDA.t293 19.7005
R4765 GNDA.n20 GNDA.t15 19.7005
R4766 GNDA.n20 GNDA.t272 19.7005
R4767 GNDA.n18 GNDA.t7 19.7005
R4768 GNDA.n18 GNDA.t229 19.7005
R4769 GNDA.n16 GNDA.t185 19.7005
R4770 GNDA.n16 GNDA.t230 19.7005
R4771 GNDA.n14 GNDA.t189 19.7005
R4772 GNDA.n14 GNDA.t228 19.7005
R4773 GNDA.n13 GNDA.t291 19.7005
R4774 GNDA.n13 GNDA.t40 19.7005
R4775 GNDA.n11 GNDA.t292 19.7005
R4776 GNDA.n11 GNDA.t218 19.7005
R4777 GNDA.n9 GNDA.t309 19.7005
R4778 GNDA.n9 GNDA.t76 19.7005
R4779 GNDA.n7 GNDA.t222 19.7005
R4780 GNDA.n7 GNDA.t330 19.7005
R4781 GNDA.n5 GNDA.t257 19.7005
R4782 GNDA.n5 GNDA.t335 19.7005
R4783 GNDA.n3 GNDA.t256 19.7005
R4784 GNDA.n3 GNDA.t254 19.7005
R4785 GNDA.n2 GNDA.t190 19.7005
R4786 GNDA.n2 GNDA.t297 19.7005
R4787 GNDA.n551 GNDA.n550 19.4279
R4788 GNDA.n1700 GNDA.n1698 19.2005
R4789 GNDA.n2154 GNDA.n2153 19.2005
R4790 GNDA.n2432 GNDA.n2431 19.2005
R4791 GNDA.n514 GNDA.n493 19.2005
R4792 GNDA.n2172 GNDA.n315 19.2005
R4793 GNDA.n1633 GNDA.n1612 19.2005
R4794 GNDA.n358 GNDA.n324 19.1005
R4795 GNDA.n2470 GNDA.n2469 19.1005
R4796 GNDA.t285 GNDA.t252 18.966
R4797 GNDA.t214 GNDA.t282 18.966
R4798 GNDA.n65 GNDA.n64 18.6842
R4799 GNDA.n352 GNDA.n351 18.6842
R4800 GNDA.n2124 GNDA.n525 18.0535
R4801 GNDA.n2183 GNDA.n2182 18.0535
R4802 GNDA.n1702 GNDA.n1633 17.613
R4803 GNDA.n2493 GNDA.n2492 17.508
R4804 GNDA.n2077 GNDA.n555 17.4917
R4805 GNDA.n2075 GNDA.n2074 16.9605
R4806 GNDA.n1875 GNDA.n590 16.9379
R4807 GNDA.n1595 GNDA.n627 16.9379
R4808 GNDA.n898 GNDA.n897 16.9379
R4809 GNDA.n429 GNDA.t240 16.9236
R4810 GNDA.n425 GNDA.t302 16.9236
R4811 GNDA.n441 GNDA.t306 16.9236
R4812 GNDA.t26 GNDA.n29 16.9236
R4813 GNDA.t329 GNDA.n30 16.9236
R4814 GNDA.t165 GNDA.t225 16.8587
R4815 GNDA.t319 GNDA.t247 16.8587
R4816 GNDA.t241 GNDA.t56 16.8587
R4817 GNDA.t243 GNDA.t226 16.8587
R4818 GNDA.t248 GNDA.t79 16.8587
R4819 GNDA.t246 GNDA.t184 16.8587
R4820 GNDA.t180 GNDA.t240 16.8587
R4821 GNDA.t245 GNDA.t3 16.8587
R4822 GNDA.t239 GNDA.t187 16.8587
R4823 GNDA.t156 GNDA.t336 16.8587
R4824 GNDA.t249 GNDA.t204 16.8587
R4825 GNDA.t237 GNDA.t37 16.8587
R4826 GNDA.t53 GNDA.t26 16.8587
R4827 GNDA.t334 GNDA.t234 16.8587
R4828 GNDA.t259 GNDA.t236 16.8587
R4829 GNDA.t66 GNDA.t329 16.8587
R4830 GNDA.t177 GNDA.t206 16.8587
R4831 GNDA.t260 GNDA.t23 16.8587
R4832 GNDA.t96 GNDA.n167 16.4123
R4833 GNDA.n1508 GNDA.n1407 16.0005
R4834 GNDA.n1502 GNDA.n1407 16.0005
R4835 GNDA.n1502 GNDA.n1501 16.0005
R4836 GNDA.n1501 GNDA.n1500 16.0005
R4837 GNDA.n1500 GNDA.n1409 16.0005
R4838 GNDA.n1494 GNDA.n1409 16.0005
R4839 GNDA.n1494 GNDA.n1493 16.0005
R4840 GNDA.n1493 GNDA.n1492 16.0005
R4841 GNDA.n1510 GNDA.n1509 16.0005
R4842 GNDA.n1510 GNDA.n1405 16.0005
R4843 GNDA.n1516 GNDA.n1405 16.0005
R4844 GNDA.n1517 GNDA.n1516 16.0005
R4845 GNDA.n1518 GNDA.n1517 16.0005
R4846 GNDA.n1518 GNDA.n1403 16.0005
R4847 GNDA.n1524 GNDA.n1403 16.0005
R4848 GNDA.n1525 GNDA.n1524 16.0005
R4849 GNDA.n1526 GNDA.n1401 16.0005
R4850 GNDA.n1401 GNDA.n1400 16.0005
R4851 GNDA.n1533 GNDA.n1400 16.0005
R4852 GNDA.n1534 GNDA.n1533 16.0005
R4853 GNDA.n1535 GNDA.n1398 16.0005
R4854 GNDA.n1398 GNDA.n1396 16.0005
R4855 GNDA.n1542 GNDA.n1396 16.0005
R4856 GNDA.n1324 GNDA.n1323 16.0005
R4857 GNDA.n1323 GNDA.n1322 16.0005
R4858 GNDA.n1322 GNDA.n1306 16.0005
R4859 GNDA.n1316 GNDA.n1306 16.0005
R4860 GNDA.n1316 GNDA.n1315 16.0005
R4861 GNDA.n1315 GNDA.n1314 16.0005
R4862 GNDA.n1314 GNDA.n1308 16.0005
R4863 GNDA.n1309 GNDA.n1308 16.0005
R4864 GNDA.n1330 GNDA.n1304 16.0005
R4865 GNDA.n1331 GNDA.n1330 16.0005
R4866 GNDA.n1332 GNDA.n1331 16.0005
R4867 GNDA.n1332 GNDA.n1302 16.0005
R4868 GNDA.n1338 GNDA.n1302 16.0005
R4869 GNDA.n1339 GNDA.n1338 16.0005
R4870 GNDA.n1340 GNDA.n1339 16.0005
R4871 GNDA.n1340 GNDA.n1300 16.0005
R4872 GNDA.n1347 GNDA.n1299 16.0005
R4873 GNDA.n1348 GNDA.n1347 16.0005
R4874 GNDA.n1349 GNDA.n1348 16.0005
R4875 GNDA.n1349 GNDA.n1297 16.0005
R4876 GNDA.n1356 GNDA.n1355 16.0005
R4877 GNDA.n1357 GNDA.n1356 16.0005
R4878 GNDA.n1357 GNDA.n1295 16.0005
R4879 GNDA.n2223 GNDA.n2222 16.0005
R4880 GNDA.n2222 GNDA.n2221 16.0005
R4881 GNDA.n2221 GNDA.n2205 16.0005
R4882 GNDA.n2215 GNDA.n2205 16.0005
R4883 GNDA.n2215 GNDA.n2214 16.0005
R4884 GNDA.n2214 GNDA.n2213 16.0005
R4885 GNDA.n2213 GNDA.n2207 16.0005
R4886 GNDA.n2208 GNDA.n2207 16.0005
R4887 GNDA.n2229 GNDA.n2203 16.0005
R4888 GNDA.n2230 GNDA.n2229 16.0005
R4889 GNDA.n2231 GNDA.n2230 16.0005
R4890 GNDA.n2231 GNDA.n2201 16.0005
R4891 GNDA.n2237 GNDA.n2201 16.0005
R4892 GNDA.n2238 GNDA.n2237 16.0005
R4893 GNDA.n2239 GNDA.n2238 16.0005
R4894 GNDA.n2239 GNDA.n2199 16.0005
R4895 GNDA.n2246 GNDA.n2198 16.0005
R4896 GNDA.n2247 GNDA.n2246 16.0005
R4897 GNDA.n2248 GNDA.n2247 16.0005
R4898 GNDA.n2248 GNDA.n2196 16.0005
R4899 GNDA.n2255 GNDA.n2254 16.0005
R4900 GNDA.n2256 GNDA.n2255 16.0005
R4901 GNDA.n2256 GNDA.n2194 16.0005
R4902 GNDA.n809 GNDA.n808 16.0005
R4903 GNDA.n808 GNDA.n807 16.0005
R4904 GNDA.n807 GNDA.n791 16.0005
R4905 GNDA.n801 GNDA.n791 16.0005
R4906 GNDA.n801 GNDA.n800 16.0005
R4907 GNDA.n800 GNDA.n799 16.0005
R4908 GNDA.n799 GNDA.n793 16.0005
R4909 GNDA.n794 GNDA.n793 16.0005
R4910 GNDA.n815 GNDA.n789 16.0005
R4911 GNDA.n816 GNDA.n815 16.0005
R4912 GNDA.n817 GNDA.n816 16.0005
R4913 GNDA.n817 GNDA.n787 16.0005
R4914 GNDA.n823 GNDA.n787 16.0005
R4915 GNDA.n824 GNDA.n823 16.0005
R4916 GNDA.n825 GNDA.n824 16.0005
R4917 GNDA.n825 GNDA.n785 16.0005
R4918 GNDA.n832 GNDA.n784 16.0005
R4919 GNDA.n833 GNDA.n832 16.0005
R4920 GNDA.n834 GNDA.n833 16.0005
R4921 GNDA.n834 GNDA.n782 16.0005
R4922 GNDA.n841 GNDA.n840 16.0005
R4923 GNDA.n842 GNDA.n841 16.0005
R4924 GNDA.n842 GNDA.n780 16.0005
R4925 GNDA.n1009 GNDA.n1008 16.0005
R4926 GNDA.n1008 GNDA.n1007 16.0005
R4927 GNDA.n1007 GNDA.n707 16.0005
R4928 GNDA.n1001 GNDA.n707 16.0005
R4929 GNDA.n1001 GNDA.n1000 16.0005
R4930 GNDA.n1000 GNDA.n999 16.0005
R4931 GNDA.n999 GNDA.n709 16.0005
R4932 GNDA.n710 GNDA.n709 16.0005
R4933 GNDA.n1015 GNDA.n705 16.0005
R4934 GNDA.n1016 GNDA.n1015 16.0005
R4935 GNDA.n1017 GNDA.n1016 16.0005
R4936 GNDA.n1017 GNDA.n703 16.0005
R4937 GNDA.n1023 GNDA.n703 16.0005
R4938 GNDA.n1024 GNDA.n1023 16.0005
R4939 GNDA.n1025 GNDA.n1024 16.0005
R4940 GNDA.n1025 GNDA.n701 16.0005
R4941 GNDA.n1032 GNDA.n700 16.0005
R4942 GNDA.n1033 GNDA.n1032 16.0005
R4943 GNDA.n1034 GNDA.n1033 16.0005
R4944 GNDA.n1034 GNDA.n698 16.0005
R4945 GNDA.n1041 GNDA.n1040 16.0005
R4946 GNDA.n1042 GNDA.n1041 16.0005
R4947 GNDA.n1042 GNDA.n693 16.0005
R4948 GNDA.n1133 GNDA.n1132 16.0005
R4949 GNDA.n1132 GNDA.n1131 16.0005
R4950 GNDA.n1131 GNDA.n1115 16.0005
R4951 GNDA.n1125 GNDA.n1115 16.0005
R4952 GNDA.n1125 GNDA.n1124 16.0005
R4953 GNDA.n1124 GNDA.n1123 16.0005
R4954 GNDA.n1123 GNDA.n1117 16.0005
R4955 GNDA.n1118 GNDA.n1117 16.0005
R4956 GNDA.n1139 GNDA.n1113 16.0005
R4957 GNDA.n1140 GNDA.n1139 16.0005
R4958 GNDA.n1141 GNDA.n1140 16.0005
R4959 GNDA.n1141 GNDA.n1111 16.0005
R4960 GNDA.n1147 GNDA.n1111 16.0005
R4961 GNDA.n1148 GNDA.n1147 16.0005
R4962 GNDA.n1149 GNDA.n1148 16.0005
R4963 GNDA.n1149 GNDA.n1109 16.0005
R4964 GNDA.n1156 GNDA.n1108 16.0005
R4965 GNDA.n1157 GNDA.n1156 16.0005
R4966 GNDA.n1158 GNDA.n1157 16.0005
R4967 GNDA.n1158 GNDA.n1106 16.0005
R4968 GNDA.n1165 GNDA.n1164 16.0005
R4969 GNDA.n1166 GNDA.n1165 16.0005
R4970 GNDA.n1166 GNDA.n1104 16.0005
R4971 GNDA.n1777 GNDA.n1755 16.0005
R4972 GNDA.n1771 GNDA.n1755 16.0005
R4973 GNDA.n1771 GNDA.n1770 16.0005
R4974 GNDA.n1770 GNDA.n1769 16.0005
R4975 GNDA.n1769 GNDA.n1757 16.0005
R4976 GNDA.n1763 GNDA.n1757 16.0005
R4977 GNDA.n1763 GNDA.n1762 16.0005
R4978 GNDA.n1762 GNDA.n1761 16.0005
R4979 GNDA.n1779 GNDA.n1778 16.0005
R4980 GNDA.n1779 GNDA.n1753 16.0005
R4981 GNDA.n1785 GNDA.n1753 16.0005
R4982 GNDA.n1786 GNDA.n1785 16.0005
R4983 GNDA.n1787 GNDA.n1786 16.0005
R4984 GNDA.n1787 GNDA.n1751 16.0005
R4985 GNDA.n1793 GNDA.n1751 16.0005
R4986 GNDA.n1794 GNDA.n1793 16.0005
R4987 GNDA.n1795 GNDA.n1749 16.0005
R4988 GNDA.n1749 GNDA.n1748 16.0005
R4989 GNDA.n1802 GNDA.n1748 16.0005
R4990 GNDA.n1803 GNDA.n1802 16.0005
R4991 GNDA.n1804 GNDA.n1746 16.0005
R4992 GNDA.n1746 GNDA.n1743 16.0005
R4993 GNDA.n1811 GNDA.n1743 16.0005
R4994 GNDA.n1986 GNDA.n1966 16.0005
R4995 GNDA.n1980 GNDA.n1966 16.0005
R4996 GNDA.n1980 GNDA.n1979 16.0005
R4997 GNDA.n1979 GNDA.n1978 16.0005
R4998 GNDA.n1978 GNDA.n1968 16.0005
R4999 GNDA.n1972 GNDA.n1968 16.0005
R5000 GNDA.n1972 GNDA.n1971 16.0005
R5001 GNDA.n1971 GNDA.n1931 16.0005
R5002 GNDA.n1988 GNDA.n1987 16.0005
R5003 GNDA.n1988 GNDA.n1964 16.0005
R5004 GNDA.n1994 GNDA.n1964 16.0005
R5005 GNDA.n1995 GNDA.n1994 16.0005
R5006 GNDA.n1996 GNDA.n1995 16.0005
R5007 GNDA.n1996 GNDA.n1962 16.0005
R5008 GNDA.n2002 GNDA.n1962 16.0005
R5009 GNDA.n2003 GNDA.n2002 16.0005
R5010 GNDA.n2004 GNDA.n1960 16.0005
R5011 GNDA.n1960 GNDA.n1959 16.0005
R5012 GNDA.n2011 GNDA.n1959 16.0005
R5013 GNDA.n2012 GNDA.n2011 16.0005
R5014 GNDA.n2013 GNDA.n1957 16.0005
R5015 GNDA.n1957 GNDA.n1954 16.0005
R5016 GNDA.n2020 GNDA.n1954 16.0005
R5017 GNDA.n2368 GNDA.n2367 16.0005
R5018 GNDA.n2367 GNDA.n2366 16.0005
R5019 GNDA.n2366 GNDA.n135 16.0005
R5020 GNDA.n2360 GNDA.n135 16.0005
R5021 GNDA.n2360 GNDA.n2359 16.0005
R5022 GNDA.n2359 GNDA.n2358 16.0005
R5023 GNDA.n2358 GNDA.n137 16.0005
R5024 GNDA.n138 GNDA.n137 16.0005
R5025 GNDA.n2374 GNDA.n133 16.0005
R5026 GNDA.n2375 GNDA.n2374 16.0005
R5027 GNDA.n2376 GNDA.n2375 16.0005
R5028 GNDA.n2376 GNDA.n131 16.0005
R5029 GNDA.n2382 GNDA.n131 16.0005
R5030 GNDA.n2383 GNDA.n2382 16.0005
R5031 GNDA.n2384 GNDA.n2383 16.0005
R5032 GNDA.n2384 GNDA.n129 16.0005
R5033 GNDA.n2391 GNDA.n128 16.0005
R5034 GNDA.n2392 GNDA.n2391 16.0005
R5035 GNDA.n2393 GNDA.n2392 16.0005
R5036 GNDA.n2393 GNDA.n126 16.0005
R5037 GNDA.n2400 GNDA.n2399 16.0005
R5038 GNDA.n2401 GNDA.n2400 16.0005
R5039 GNDA.n2401 GNDA.n89 16.0005
R5040 GNDA.n2077 GNDA.n2076 16.0005
R5041 GNDA.n2076 GNDA.n2075 16.0005
R5042 GNDA.t331 GNDA.t0 15.8816
R5043 GNDA.t36 GNDA.t78 15.8816
R5044 GNDA.n1704 GNDA.n1630 15.363
R5045 GNDA.n1717 GNDA.n1704 15.363
R5046 GNDA.t27 GNDA.n2149 14.7711
R5047 GNDA.t29 GNDA.n2428 14.7711
R5048 GNDA.n448 GNDA.n447 14.2068
R5049 GNDA.n448 GNDA.n375 14.2068
R5050 GNDA.n478 GNDA.n477 14.0505
R5051 GNDA.n2476 GNDA.n2475 14.0505
R5052 GNDA.n1535 GNDA 14.0449
R5053 GNDA.n1355 GNDA 14.0449
R5054 GNDA.n2254 GNDA 14.0449
R5055 GNDA.n840 GNDA 14.0449
R5056 GNDA.n1040 GNDA 14.0449
R5057 GNDA.n1164 GNDA 14.0449
R5058 GNDA.n1804 GNDA 14.0449
R5059 GNDA.n2013 GNDA 14.0449
R5060 GNDA.n2399 GNDA 14.0449
R5061 GNDA.n2490 GNDA.n2489 14.0193
R5062 GNDA.n2481 GNDA.n2480 13.8005
R5063 GNDA.n416 GNDA.n415 13.8005
R5064 GNDA.n1701 GNDA.n1700 13.8005
R5065 GNDA.n1674 GNDA.n555 13.7706
R5066 GNDA.n389 GNDA.t242 13.4979
R5067 GNDA.t162 GNDA.n454 13.4979
R5068 GNDA.n2292 GNDA.n256 12.9309
R5069 GNDA.n1391 GNDA.n650 12.9309
R5070 GNDA.n715 GNDA.n628 12.9309
R5071 GNDA.n1202 GNDA.n181 12.9309
R5072 GNDA.n320 GNDA.n319 12.8005
R5073 GNDA.n2454 GNDA.n69 12.8005
R5074 GNDA.n481 GNDA.t93 12.6442
R5075 GNDA.t338 GNDA.t144 12.6442
R5076 GNDA.t326 GNDA.t317 12.6442
R5077 GNDA.n428 GNDA.t84 12.6442
R5078 GNDA.t31 GNDA.n2485 12.6442
R5079 GNDA.t21 GNDA.t9 12.6442
R5080 GNDA.t171 GNDA.t38 12.6442
R5081 GNDA.n55 GNDA.t98 12.6442
R5082 GNDA.n2187 GNDA.n307 12.5829
R5083 GNDA.n217 GNDA.n214 12.4126
R5084 GNDA.n2127 GNDA.n527 12.4126
R5085 GNDA.n500 GNDA.n173 12.4126
R5086 GNDA.n1265 GNDA.n1215 11.6369
R5087 GNDA.n1265 GNDA.n1264 11.6369
R5088 GNDA.n1264 GNDA.n1263 11.6369
R5089 GNDA.n1263 GNDA.n1260 11.6369
R5090 GNDA.n1260 GNDA.n1259 11.6369
R5091 GNDA.n1259 GNDA.n1256 11.6369
R5092 GNDA.n1256 GNDA.n1255 11.6369
R5093 GNDA.n1255 GNDA.n1252 11.6369
R5094 GNDA.n1252 GNDA.n1251 11.6369
R5095 GNDA.n1251 GNDA.n1248 11.6369
R5096 GNDA.n1248 GNDA.n1247 11.6369
R5097 GNDA.n255 GNDA.n208 11.6369
R5098 GNDA.n250 GNDA.n208 11.6369
R5099 GNDA.n250 GNDA.n249 11.6369
R5100 GNDA.n249 GNDA.n210 11.6369
R5101 GNDA.n244 GNDA.n210 11.6369
R5102 GNDA.n244 GNDA.n243 11.6369
R5103 GNDA.n243 GNDA.n242 11.6369
R5104 GNDA.n242 GNDA.n212 11.6369
R5105 GNDA.n236 GNDA.n212 11.6369
R5106 GNDA.n236 GNDA.n235 11.6369
R5107 GNDA.n235 GNDA.n234 11.6369
R5108 GNDA.n220 GNDA.n217 11.6369
R5109 GNDA.n225 GNDA.n220 11.6369
R5110 GNDA.n225 GNDA.n224 11.6369
R5111 GNDA.n224 GNDA.n223 11.6369
R5112 GNDA.n223 GNDA.n113 11.6369
R5113 GNDA.n2423 GNDA.n113 11.6369
R5114 GNDA.n2426 GNDA.n2424 11.6369
R5115 GNDA.n2426 GNDA.n2425 11.6369
R5116 GNDA.n1876 GNDA.n1875 11.6369
R5117 GNDA.n1877 GNDA.n1876 11.6369
R5118 GNDA.n1877 GNDA.n588 11.6369
R5119 GNDA.n1883 GNDA.n588 11.6369
R5120 GNDA.n1884 GNDA.n1883 11.6369
R5121 GNDA.n1885 GNDA.n1884 11.6369
R5122 GNDA.n1885 GNDA.n586 11.6369
R5123 GNDA.n1891 GNDA.n586 11.6369
R5124 GNDA.n1892 GNDA.n1891 11.6369
R5125 GNDA.n1893 GNDA.n1892 11.6369
R5126 GNDA.n1893 GNDA.n583 11.6369
R5127 GNDA.n595 GNDA.n590 11.6369
R5128 GNDA.n1867 GNDA.n595 11.6369
R5129 GNDA.n1867 GNDA.n1866 11.6369
R5130 GNDA.n1866 GNDA.n1865 11.6369
R5131 GNDA.n1865 GNDA.n596 11.6369
R5132 GNDA.n1859 GNDA.n596 11.6369
R5133 GNDA.n1859 GNDA.n1858 11.6369
R5134 GNDA.n1858 GNDA.n1857 11.6369
R5135 GNDA.n1857 GNDA.n600 11.6369
R5136 GNDA.n682 GNDA.n681 11.6369
R5137 GNDA.n681 GNDA.n680 11.6369
R5138 GNDA.n680 GNDA.n678 11.6369
R5139 GNDA.n678 GNDA.n675 11.6369
R5140 GNDA.n675 GNDA.n674 11.6369
R5141 GNDA.n674 GNDA.n671 11.6369
R5142 GNDA.n671 GNDA.n670 11.6369
R5143 GNDA.n670 GNDA.n667 11.6369
R5144 GNDA.n667 GNDA.n666 11.6369
R5145 GNDA.n666 GNDA.n663 11.6369
R5146 GNDA.n663 GNDA.n662 11.6369
R5147 GNDA.n1595 GNDA.n1594 11.6369
R5148 GNDA.n1594 GNDA.n1593 11.6369
R5149 GNDA.n1593 GNDA.n1591 11.6369
R5150 GNDA.n1591 GNDA.n1588 11.6369
R5151 GNDA.n1588 GNDA.n1587 11.6369
R5152 GNDA.n1587 GNDA.n1584 11.6369
R5153 GNDA.n1584 GNDA.n1583 11.6369
R5154 GNDA.n1583 GNDA.n1580 11.6369
R5155 GNDA.n1580 GNDA.n1579 11.6369
R5156 GNDA.n1579 GNDA.n1576 11.6369
R5157 GNDA.n1576 GNDA.n1575 11.6369
R5158 GNDA.n1424 GNDA.n627 11.6369
R5159 GNDA.n1430 GNDA.n1424 11.6369
R5160 GNDA.n1431 GNDA.n1430 11.6369
R5161 GNDA.n1432 GNDA.n1431 11.6369
R5162 GNDA.n1432 GNDA.n1420 11.6369
R5163 GNDA.n1438 GNDA.n1420 11.6369
R5164 GNDA.n1439 GNDA.n1438 11.6369
R5165 GNDA.n1440 GNDA.n1439 11.6369
R5166 GNDA.n1440 GNDA.n1416 11.6369
R5167 GNDA.n897 GNDA.n736 11.6369
R5168 GNDA.n891 GNDA.n736 11.6369
R5169 GNDA.n891 GNDA.n890 11.6369
R5170 GNDA.n890 GNDA.n889 11.6369
R5171 GNDA.n889 GNDA.n740 11.6369
R5172 GNDA.n883 GNDA.n740 11.6369
R5173 GNDA.n883 GNDA.n882 11.6369
R5174 GNDA.n882 GNDA.n881 11.6369
R5175 GNDA.n881 GNDA.n744 11.6369
R5176 GNDA.n899 GNDA.n898 11.6369
R5177 GNDA.n899 GNDA.n732 11.6369
R5178 GNDA.n906 GNDA.n732 11.6369
R5179 GNDA.n907 GNDA.n906 11.6369
R5180 GNDA.n908 GNDA.n907 11.6369
R5181 GNDA.n908 GNDA.n730 11.6369
R5182 GNDA.n913 GNDA.n730 11.6369
R5183 GNDA.n914 GNDA.n913 11.6369
R5184 GNDA.n916 GNDA.n914 11.6369
R5185 GNDA.n916 GNDA.n915 11.6369
R5186 GNDA.n915 GNDA.n727 11.6369
R5187 GNDA.n2065 GNDA.n560 11.6369
R5188 GNDA.n2066 GNDA.n2065 11.6369
R5189 GNDA.n2067 GNDA.n2066 11.6369
R5190 GNDA.n2067 GNDA.n556 11.6369
R5191 GNDA.n2073 GNDA.n556 11.6369
R5192 GNDA.n2083 GNDA.n546 11.6369
R5193 GNDA.n2084 GNDA.n2083 11.6369
R5194 GNDA.n2086 GNDA.n2084 11.6369
R5195 GNDA.n2086 GNDA.n2085 11.6369
R5196 GNDA.n2085 GNDA.n543 11.6369
R5197 GNDA.n2100 GNDA.n537 11.6369
R5198 GNDA.n2101 GNDA.n2100 11.6369
R5199 GNDA.n2102 GNDA.n2101 11.6369
R5200 GNDA.n2102 GNDA.n533 11.6369
R5201 GNDA.n2108 GNDA.n533 11.6369
R5202 GNDA.n2109 GNDA.n2108 11.6369
R5203 GNDA.n2110 GNDA.n2109 11.6369
R5204 GNDA.n2110 GNDA.n529 11.6369
R5205 GNDA.n2117 GNDA.n529 11.6369
R5206 GNDA.n2118 GNDA.n2117 11.6369
R5207 GNDA.n2119 GNDA.n2118 11.6369
R5208 GNDA.n2128 GNDA.n2127 11.6369
R5209 GNDA.n2129 GNDA.n2128 11.6369
R5210 GNDA.n2129 GNDA.n523 11.6369
R5211 GNDA.n2136 GNDA.n523 11.6369
R5212 GNDA.n2137 GNDA.n2136 11.6369
R5213 GNDA.n2138 GNDA.n2137 11.6369
R5214 GNDA.n2144 GNDA.n520 11.6369
R5215 GNDA.n2145 GNDA.n2144 11.6369
R5216 GNDA.n2304 GNDA.n2303 11.6369
R5217 GNDA.n2305 GNDA.n2304 11.6369
R5218 GNDA.n2305 GNDA.n179 11.6369
R5219 GNDA.n2311 GNDA.n179 11.6369
R5220 GNDA.n2312 GNDA.n2311 11.6369
R5221 GNDA.n2313 GNDA.n2312 11.6369
R5222 GNDA.n2313 GNDA.n177 11.6369
R5223 GNDA.n2319 GNDA.n177 11.6369
R5224 GNDA.n2320 GNDA.n2319 11.6369
R5225 GNDA.n2321 GNDA.n2320 11.6369
R5226 GNDA.n2321 GNDA.n175 11.6369
R5227 GNDA.n501 GNDA.n500 11.6369
R5228 GNDA.n502 GNDA.n501 11.6369
R5229 GNDA.n502 GNDA.n496 11.6369
R5230 GNDA.n2162 GNDA.n496 11.6369
R5231 GNDA.n2163 GNDA.n2162 11.6369
R5232 GNDA.n2166 GNDA.n2163 11.6369
R5233 GNDA.n2165 GNDA.n2164 11.6369
R5234 GNDA.n2164 GNDA.n310 11.6369
R5235 GNDA.n2424 GNDA 11.5076
R5236 GNDA GNDA.n520 11.5076
R5237 GNDA GNDA.n2165 11.5076
R5238 GNDA.n2425 GNDA.n90 11.4026
R5239 GNDA.n2146 GNDA.n2145 11.4026
R5240 GNDA.n310 GNDA.n309 11.4026
R5241 GNDA.n1850 GNDA.n600 11.249
R5242 GNDA.n1448 GNDA.n1416 11.249
R5243 GNDA.n747 GNDA.n744 11.249
R5244 GNDA.n450 GNDA.n449 11.0505
R5245 GNDA.n449 GNDA.n374 10.488
R5246 GNDA.n2074 GNDA.n2073 10.4732
R5247 GNDA.n1703 GNDA.n1631 9.78488
R5248 GNDA GNDA.n0 9.67325
R5249 GNDA.n2080 GNDA.n2079 9.65197
R5250 GNDA.n1699 GNDA.t294 9.6005
R5251 GNDA.n1699 GNDA.t296 9.6005
R5252 GNDA.n413 GNDA.t132 9.6005
R5253 GNDA.n413 GNDA.t322 9.6005
R5254 GNDA.n411 GNDA.t69 9.6005
R5255 GNDA.n411 GNDA.t314 9.6005
R5256 GNDA.n409 GNDA.t196 9.6005
R5257 GNDA.n409 GNDA.t72 9.6005
R5258 GNDA.n407 GNDA.t19 9.6005
R5259 GNDA.n407 GNDA.t55 9.6005
R5260 GNDA.n405 GNDA.t232 9.6005
R5261 GNDA.n405 GNDA.t220 9.6005
R5262 GNDA.n403 GNDA.t281 9.6005
R5263 GNDA.n403 GNDA.t202 9.6005
R5264 GNDA.n401 GNDA.t213 9.6005
R5265 GNDA.n401 GNDA.t191 9.6005
R5266 GNDA.n399 GNDA.t35 9.6005
R5267 GNDA.n399 GNDA.t316 9.6005
R5268 GNDA.n397 GNDA.t48 9.6005
R5269 GNDA.n397 GNDA.t5 9.6005
R5270 GNDA.n395 GNDA.t182 9.6005
R5271 GNDA.n395 GNDA.t262 9.6005
R5272 GNDA.n393 GNDA.t61 9.6005
R5273 GNDA.n393 GNDA.t63 9.6005
R5274 GNDA.n35 GNDA.t46 9.6005
R5275 GNDA.n35 GNDA.t118 9.6005
R5276 GNDA.n1632 GNDA.t290 9.6005
R5277 GNDA.n1632 GNDA.t298 9.6005
R5278 GNDA.n1701 GNDA.n1634 9.37925
R5279 GNDA.n2151 GNDA.n513 9.30051
R5280 GNDA.n2429 GNDA.n103 9.30051
R5281 GNDA.n2480 GNDA.n2479 9.0005
R5282 GNDA.n415 GNDA.n1 8.96925
R5283 GNDA.n2150 GNDA.t27 8.75345
R5284 GNDA.n234 GNDA.n214 8.66313
R5285 GNDA.n2119 GNDA.n527 8.66313
R5286 GNDA.n175 GNDA.n173 8.66313
R5287 GNDA.n1247 GNDA.n256 8.53383
R5288 GNDA.n650 GNDA.n583 8.53383
R5289 GNDA.n662 GNDA.n181 8.53383
R5290 GNDA.n1575 GNDA.n628 8.53383
R5291 GNDA.n727 GNDA.n726 8.53383
R5292 GNDA.n543 GNDA.n542 8.53383
R5293 GNDA.n1673 GNDA.n1672 8.44175
R5294 GNDA.t221 GNDA.n440 8.42962
R5295 GNDA.n1492 GNDA.n1411 8.35606
R5296 GNDA.n1309 GNDA.n653 8.35606
R5297 GNDA.n2208 GNDA.n282 8.35606
R5298 GNDA.n794 GNDA.n750 8.35606
R5299 GNDA.n959 GNDA.n710 8.35606
R5300 GNDA.n1118 GNDA.n1077 8.35606
R5301 GNDA.n1761 GNDA.n604 8.35606
R5302 GNDA.n2057 GNDA.n1931 8.35606
R5303 GNDA.n2331 GNDA.n138 8.35606
R5304 GNDA.n1704 GNDA.n1703 7.71925
R5305 GNDA.t178 GNDA.n2150 7.65933
R5306 GNDA.n2158 GNDA.n2157 7.11227
R5307 GNDA.n65 GNDA.t323 7.00687
R5308 GNDA.t325 GNDA.n77 7.00687
R5309 GNDA.n341 GNDA.t328 7.00687
R5310 GNDA.n351 GNDA.t332 7.00687
R5311 GNDA.n2491 GNDA.n2490 6.7505
R5312 GNDA.n2490 GNDA.n24 6.688
R5313 GNDA.n476 GNDA.n1 6.563
R5314 GNDA.n2479 GNDA.n2478 6.563
R5315 GNDA.n2173 GNDA.n2172 6.4005
R5316 GNDA.t51 GNDA.n1707 6.32234
R5317 GNDA.t33 GNDA.t153 6.32234
R5318 GNDA.n1731 GNDA.t267 6.32234
R5319 GNDA.n1643 GNDA.t10 6.32234
R5320 GNDA.t137 GNDA.t318 6.32234
R5321 GNDA.t197 GNDA.n1641 6.32234
R5322 GNDA.n2479 GNDA.n24 5.03175
R5323 GNDA.n551 GNDA.n0 5.02613
R5324 GNDA.n2151 GNDA.t233 4.92404
R5325 GNDA GNDA.n2493 4.8321
R5326 GNDA.n1817 GNDA.n1816 4.6085
R5327 GNDA.n2026 GNDA.n2025 4.6085
R5328 GNDA.n2439 GNDA.n2438 4.6085
R5329 GNDA.n778 GNDA.n771 4.6085
R5330 GNDA.n1205 GNDA.n1204 4.6085
R5331 GNDA.n1102 GNDA.n519 4.6085
R5332 GNDA.n1549 GNDA.n1393 4.6085
R5333 GNDA.n1293 GNDA.n207 4.6085
R5334 GNDA.n2192 GNDA.n304 4.6085
R5335 GNDA.n1243 GNDA.n1216 4.55161
R5336 GNDA.n1900 GNDA.n581 4.55161
R5337 GNDA.n1571 GNDA.n629 4.55161
R5338 GNDA.n925 GNDA.n724 4.55161
R5339 GNDA.n2094 GNDA.n538 4.55161
R5340 GNDA.n2299 GNDA.n182 4.55161
R5341 GNDA.n1812 GNDA.n569 4.5061
R5342 GNDA.n2022 GNDA.n146 4.5061
R5343 GNDA.n773 GNDA.n715 4.5061
R5344 GNDA.n1203 GNDA.n1202 4.5061
R5345 GNDA.n1550 GNDA.n1391 4.5061
R5346 GNDA.n2293 GNDA.n2292 4.5061
R5347 GNDA.n449 GNDA.n448 4.5005
R5348 GNDA.n2492 GNDA.n2491 4.5005
R5349 GNDA.n1703 GNDA.n1702 4.5005
R5350 GNDA.n1215 GNDA.n650 4.39646
R5351 GNDA.n256 GNDA.n255 4.39646
R5352 GNDA.n682 GNDA.n628 4.39646
R5353 GNDA.n726 GNDA.n560 4.39646
R5354 GNDA.n542 GNDA.n537 4.39646
R5355 GNDA.n2303 GNDA.n181 4.39646
R5356 GNDA.n1930 GNDA.n569 4.3525
R5357 GNDA.n2330 GNDA.n146 4.3525
R5358 GNDA.n715 GNDA.n712 4.3525
R5359 GNDA.n1202 GNDA.n1201 4.3525
R5360 GNDA.n1391 GNDA.n1390 4.3525
R5361 GNDA.n2292 GNDA.n2291 4.3525
R5362 GNDA.n2058 GNDA.n1930 4.3013
R5363 GNDA.n2332 GNDA.n2330 4.3013
R5364 GNDA.n958 GNDA.n712 4.3013
R5365 GNDA.n1201 GNDA.n1198 4.3013
R5366 GNDA.n1390 GNDA.n1389 4.3013
R5367 GNDA.n2291 GNDA.n2288 4.3013
R5368 GNDA.n1243 GNDA.n1242 4.26717
R5369 GNDA.n1242 GNDA.n1239 4.26717
R5370 GNDA.n1239 GNDA.n1238 4.26717
R5371 GNDA.n1238 GNDA.n1235 4.26717
R5372 GNDA.n1235 GNDA.n1234 4.26717
R5373 GNDA.n1234 GNDA.n1231 4.26717
R5374 GNDA.n1230 GNDA.n1227 4.26717
R5375 GNDA.n1227 GNDA.n1226 4.26717
R5376 GNDA.n1900 GNDA.n579 4.26717
R5377 GNDA.n1906 GNDA.n579 4.26717
R5378 GNDA.n1906 GNDA.n577 4.26717
R5379 GNDA.n1912 GNDA.n577 4.26717
R5380 GNDA.n1912 GNDA.n575 4.26717
R5381 GNDA.n1919 GNDA.n575 4.26717
R5382 GNDA.n573 GNDA.n571 4.26717
R5383 GNDA.n1926 GNDA.n571 4.26717
R5384 GNDA.n1571 GNDA.n1570 4.26717
R5385 GNDA.n1570 GNDA.n634 4.26717
R5386 GNDA.n1565 GNDA.n634 4.26717
R5387 GNDA.n1565 GNDA.n1564 4.26717
R5388 GNDA.n1564 GNDA.n1563 4.26717
R5389 GNDA.n1563 GNDA.n642 4.26717
R5390 GNDA.n1557 GNDA.n1556 4.26717
R5391 GNDA.n1556 GNDA.n1555 4.26717
R5392 GNDA.n925 GNDA.n723 4.26717
R5393 GNDA.n931 GNDA.n723 4.26717
R5394 GNDA.n931 GNDA.n721 4.26717
R5395 GNDA.n937 GNDA.n721 4.26717
R5396 GNDA.n937 GNDA.n719 4.26717
R5397 GNDA.n945 GNDA.n719 4.26717
R5398 GNDA.n717 GNDA.n714 4.26717
R5399 GNDA.n952 GNDA.n714 4.26717
R5400 GNDA.n2094 GNDA.n539 4.26717
R5401 GNDA.n1055 GNDA.n539 4.26717
R5402 GNDA.n1056 GNDA.n1055 4.26717
R5403 GNDA.n1061 GNDA.n1056 4.26717
R5404 GNDA.n1062 GNDA.n1061 4.26717
R5405 GNDA.n1067 GNDA.n1062 4.26717
R5406 GNDA.n1073 GNDA.n1068 4.26717
R5407 GNDA.n1075 GNDA.n1073 4.26717
R5408 GNDA.n2299 GNDA.n183 4.26717
R5409 GNDA.n260 GNDA.n183 4.26717
R5410 GNDA.n261 GNDA.n260 4.26717
R5411 GNDA.n266 GNDA.n261 4.26717
R5412 GNDA.n267 GNDA.n266 4.26717
R5413 GNDA.n272 GNDA.n267 4.26717
R5414 GNDA.n278 GNDA.n273 4.26717
R5415 GNDA.n280 GNDA.n278 4.26717
R5416 GNDA.n748 GNDA.n747 4.2501
R5417 GNDA.n1449 GNDA.n1448 4.2501
R5418 GNDA GNDA.n1230 4.21976
R5419 GNDA GNDA.n573 4.21976
R5420 GNDA.n1557 GNDA 4.21976
R5421 GNDA GNDA.n717 4.21976
R5422 GNDA.n1068 GNDA 4.21976
R5423 GNDA.n273 GNDA 4.21976
R5424 GNDA.t106 GNDA.t134 4.21506
R5425 GNDA.n421 GNDA.t242 4.21506
R5426 GNDA.n390 GNDA.t321 4.21506
R5427 GNDA.t244 GNDA.n428 4.21506
R5428 GNDA.n2486 GNDA.t336 4.21506
R5429 GNDA.n2485 GNDA.t324 4.21506
R5430 GNDA.t81 GNDA.t90 4.21506
R5431 GNDA.n1850 GNDA.n1849 4.1477
R5432 GNDA.n1226 GNDA.n146 4.12494
R5433 GNDA.n1926 GNDA.n569 4.12494
R5434 GNDA.n1555 GNDA.n1391 4.12494
R5435 GNDA.n952 GNDA.n715 4.12494
R5436 GNDA.n1202 GNDA.n1075 4.12494
R5437 GNDA.n2292 GNDA.n280 4.12494
R5438 GNDA.t233 GNDA.t178 3.82992
R5439 GNDA.n1702 GNDA.n1701 3.813
R5440 GNDA.n1634 GNDA 3.68412
R5441 GNDA.n609 GNDA.n608 3.5845
R5442 GNDA.n1843 GNDA.n1842 3.5845
R5443 GNDA.n1838 GNDA.n610 3.5845
R5444 GNDA.n1837 GNDA.n613 3.5845
R5445 GNDA.n1602 GNDA.n1601 3.5845
R5446 GNDA.n1831 GNDA.n1830 3.5845
R5447 GNDA.n1826 GNDA.n1603 3.5845
R5448 GNDA.n1825 GNDA.n1607 3.5845
R5449 GNDA.n1742 GNDA.n1741 3.5845
R5450 GNDA.n2056 GNDA.n2055 3.5845
R5451 GNDA.n1934 GNDA.n1932 3.5845
R5452 GNDA.n2050 GNDA.n1936 3.5845
R5453 GNDA.n2049 GNDA.n1937 3.5845
R5454 GNDA.n2041 GNDA.n2040 3.5845
R5455 GNDA.n1942 GNDA.n1940 3.5845
R5456 GNDA.n2035 GNDA.n1944 3.5845
R5457 GNDA.n2034 GNDA.n1945 3.5845
R5458 GNDA.n1953 GNDA.n1952 3.5845
R5459 GNDA.n2351 GNDA.n140 3.5845
R5460 GNDA.n2350 GNDA.n141 3.5845
R5461 GNDA.n2337 GNDA.n2336 3.5845
R5462 GNDA.n2344 GNDA.n2343 3.5845
R5463 GNDA.n2338 GNDA.n122 3.5845
R5464 GNDA.n2418 GNDA.n2417 3.5845
R5465 GNDA.n2413 GNDA.n123 3.5845
R5466 GNDA.n2412 GNDA.n2409 3.5845
R5467 GNDA.n2408 GNDA.n88 3.5845
R5468 GNDA.n870 GNDA.n869 3.5845
R5469 GNDA.n753 GNDA.n751 3.5845
R5470 GNDA.n864 GNDA.n755 3.5845
R5471 GNDA.n863 GNDA.n756 3.5845
R5472 GNDA.n859 GNDA.n858 3.5845
R5473 GNDA.n762 GNDA.n760 3.5845
R5474 GNDA.n853 GNDA.n764 3.5845
R5475 GNDA.n852 GNDA.n765 3.5845
R5476 GNDA.n848 GNDA.n847 3.5845
R5477 GNDA.n992 GNDA.n960 3.5845
R5478 GNDA.n991 GNDA.n988 3.5845
R5479 GNDA.n987 GNDA.n961 3.5845
R5480 GNDA.n984 GNDA.n983 3.5845
R5481 GNDA.n979 GNDA.n962 3.5845
R5482 GNDA.n978 GNDA.n975 3.5845
R5483 GNDA.n974 GNDA.n966 3.5845
R5484 GNDA.n971 GNDA.n970 3.5845
R5485 GNDA.n1047 GNDA.n695 3.5845
R5486 GNDA.n1194 GNDA.n1193 3.5845
R5487 GNDA.n1081 GNDA.n1079 3.5845
R5488 GNDA.n1188 GNDA.n1083 3.5845
R5489 GNDA.n1187 GNDA.n1084 3.5845
R5490 GNDA.n1183 GNDA.n1182 3.5845
R5491 GNDA.n1090 GNDA.n1088 3.5845
R5492 GNDA.n1177 GNDA.n1092 3.5845
R5493 GNDA.n1176 GNDA.n1093 3.5845
R5494 GNDA.n1172 GNDA.n1171 3.5845
R5495 GNDA.n1488 GNDA.n1413 3.5845
R5496 GNDA.n1487 GNDA.n1414 3.5845
R5497 GNDA.n1483 GNDA.n1482 3.5845
R5498 GNDA.n1456 GNDA.n1454 3.5845
R5499 GNDA.n1477 GNDA.n1458 3.5845
R5500 GNDA.n1476 GNDA.n1459 3.5845
R5501 GNDA.n1472 GNDA.n1471 3.5845
R5502 GNDA.n1467 GNDA.n1464 3.5845
R5503 GNDA.n1466 GNDA.n1395 3.5845
R5504 GNDA.n1385 GNDA.n1384 3.5845
R5505 GNDA.n1273 GNDA.n1271 3.5845
R5506 GNDA.n1379 GNDA.n1275 3.5845
R5507 GNDA.n1378 GNDA.n1276 3.5845
R5508 GNDA.n1374 GNDA.n1373 3.5845
R5509 GNDA.n1282 GNDA.n1280 3.5845
R5510 GNDA.n1368 GNDA.n1284 3.5845
R5511 GNDA.n1367 GNDA.n1285 3.5845
R5512 GNDA.n1363 GNDA.n1362 3.5845
R5513 GNDA.n2284 GNDA.n2283 3.5845
R5514 GNDA.n286 GNDA.n284 3.5845
R5515 GNDA.n2278 GNDA.n288 3.5845
R5516 GNDA.n2277 GNDA.n289 3.5845
R5517 GNDA.n2273 GNDA.n2272 3.5845
R5518 GNDA.n295 GNDA.n293 3.5845
R5519 GNDA.n2267 GNDA.n297 3.5845
R5520 GNDA.n2266 GNDA.n298 3.5845
R5521 GNDA.n2262 GNDA.n2261 3.5845
R5522 GNDA.n37 GNDA.t280 3.42907
R5523 GNDA.n37 GNDA.t264 3.42907
R5524 GNDA.n2477 GNDA.t22 3.42907
R5525 GNDA.n2477 GNDA.t58 3.42907
R5526 GNDA.n475 GNDA.t194 3.42907
R5527 GNDA.n475 GNDA.t327 3.42907
R5528 GNDA.n474 GNDA.t224 3.42907
R5529 GNDA.n474 GNDA.t75 3.42907
R5530 GNDA.n1849 GNDA.n604 3.3797
R5531 GNDA.n2058 GNDA.n2057 3.3797
R5532 GNDA.n2332 GNDA.n2331 3.3797
R5533 GNDA.n750 GNDA.n748 3.3797
R5534 GNDA.n959 GNDA.n958 3.3797
R5535 GNDA.n1198 GNDA.n1077 3.3797
R5536 GNDA.n1449 GNDA.n1411 3.3797
R5537 GNDA.n1389 GNDA.n653 3.3797
R5538 GNDA.n2288 GNDA.n282 3.3797
R5539 GNDA.n2429 GNDA.t238 3.28286
R5540 GNDA.n104 GNDA.n98 3.2005
R5541 GNDA.n315 GNDA.n314 3.2005
R5542 GNDA.n1819 GNDA.n1818 2.8677
R5543 GNDA.n2028 GNDA.n2027 2.8677
R5544 GNDA.n2441 GNDA.n2440 2.8677
R5545 GNDA.n779 GNDA.n769 2.8677
R5546 GNDA.n1049 GNDA.n1048 2.8677
R5547 GNDA.n1103 GNDA.n1097 2.8677
R5548 GNDA.n1544 GNDA.n1543 2.8677
R5549 GNDA.n1294 GNDA.n1289 2.8677
R5550 GNDA.n2193 GNDA.n302 2.8677
R5551 GNDA.n389 GNDA.t67 2.75116
R5552 GNDA.n454 GNDA.t205 2.75116
R5553 GNDA.n1660 GNDA.n1658 2.34425
R5554 GNDA.n1668 GNDA.n1666 2.34425
R5555 GNDA.t323 GNDA.n62 2.33596
R5556 GNDA.n2459 GNDA.t24 2.33596
R5557 GNDA.t20 GNDA.n345 2.33596
R5558 GNDA.n344 GNDA.t332 2.33596
R5559 GNDA.n1543 GNDA.n1542 2.31161
R5560 GNDA.n1295 GNDA.n1294 2.31161
R5561 GNDA.n2194 GNDA.n2193 2.31161
R5562 GNDA.n780 GNDA.n779 2.31161
R5563 GNDA.n1049 GNDA.n693 2.31161
R5564 GNDA.n1104 GNDA.n1103 2.31161
R5565 GNDA.n1818 GNDA.n1811 2.31161
R5566 GNDA.n2027 GNDA.n2020 2.31161
R5567 GNDA.n2440 GNDA.n89 2.31161
R5568 GNDA GNDA.n1534 1.95606
R5569 GNDA.n1297 GNDA 1.95606
R5570 GNDA.n2196 GNDA 1.95606
R5571 GNDA.n782 GNDA 1.95606
R5572 GNDA.n698 GNDA 1.95606
R5573 GNDA.n1106 GNDA 1.95606
R5574 GNDA GNDA.n1803 1.95606
R5575 GNDA GNDA.n2012 1.95606
R5576 GNDA.n126 GNDA 1.95606
R5577 GNDA.n1818 GNDA.n1817 1.7413
R5578 GNDA.n2027 GNDA.n2026 1.7413
R5579 GNDA.n2440 GNDA.n2439 1.7413
R5580 GNDA.n779 GNDA.n778 1.7413
R5581 GNDA.n1205 GNDA.n1049 1.7413
R5582 GNDA.n1103 GNDA.n1102 1.7413
R5583 GNDA.n1543 GNDA.n1393 1.7413
R5584 GNDA.n1294 GNDA.n1293 1.7413
R5585 GNDA.n2193 GNDA.n2192 1.7413
R5586 GNDA.n555 GNDA.n554 1.73362
R5587 GNDA.n2169 GNDA.n311 1.64168
R5588 GNDA.n2489 GNDA.n25 1.6005
R5589 GNDA.n608 GNDA.n604 1.2293
R5590 GNDA.n2057 GNDA.n2056 1.2293
R5591 GNDA.n2331 GNDA.n140 1.2293
R5592 GNDA.n870 GNDA.n750 1.2293
R5593 GNDA.n960 GNDA.n959 1.2293
R5594 GNDA.n1194 GNDA.n1077 1.2293
R5595 GNDA.n1413 GNDA.n1411 1.2293
R5596 GNDA.n1385 GNDA.n653 1.2293
R5597 GNDA.n2284 GNDA.n282 1.2293
R5598 GNDA.n1816 GNDA.n1812 1.1781
R5599 GNDA.n2025 GNDA.n2022 1.1781
R5600 GNDA.n2438 GNDA.n90 1.1781
R5601 GNDA.n773 GNDA.n771 1.1781
R5602 GNDA.n1204 GNDA.n1203 1.1781
R5603 GNDA.n2146 GNDA.n519 1.1781
R5604 GNDA.n1550 GNDA.n1549 1.1781
R5605 GNDA.n2293 GNDA.n207 1.1781
R5606 GNDA.n309 GNDA.n304 1.1781
R5607 GNDA.n2074 GNDA.n546 1.16414
R5608 GNDA.n1843 GNDA.n609 1.0245
R5609 GNDA.n1842 GNDA.n610 1.0245
R5610 GNDA.n1838 GNDA.n1837 1.0245
R5611 GNDA.n1601 GNDA.n613 1.0245
R5612 GNDA.n1831 GNDA.n1602 1.0245
R5613 GNDA.n1830 GNDA.n1603 1.0245
R5614 GNDA.n1826 GNDA.n1825 1.0245
R5615 GNDA.n1741 GNDA.n1607 1.0245
R5616 GNDA.n1819 GNDA.n1742 1.0245
R5617 GNDA.n2055 GNDA.n1932 1.0245
R5618 GNDA.n1936 GNDA.n1934 1.0245
R5619 GNDA.n2050 GNDA.n2049 1.0245
R5620 GNDA.n2041 GNDA.n1937 1.0245
R5621 GNDA.n2040 GNDA.n1940 1.0245
R5622 GNDA.n1944 GNDA.n1942 1.0245
R5623 GNDA.n2035 GNDA.n2034 1.0245
R5624 GNDA.n1952 GNDA.n1945 1.0245
R5625 GNDA.n2028 GNDA.n1953 1.0245
R5626 GNDA.n2351 GNDA.n2350 1.0245
R5627 GNDA.n2336 GNDA.n141 1.0245
R5628 GNDA.n2344 GNDA.n2337 1.0245
R5629 GNDA.n2343 GNDA.n2338 1.0245
R5630 GNDA.n2418 GNDA.n122 1.0245
R5631 GNDA.n2417 GNDA.n123 1.0245
R5632 GNDA.n2413 GNDA.n2412 1.0245
R5633 GNDA.n2409 GNDA.n2408 1.0245
R5634 GNDA.n2441 GNDA.n88 1.0245
R5635 GNDA.n869 GNDA.n751 1.0245
R5636 GNDA.n755 GNDA.n753 1.0245
R5637 GNDA.n864 GNDA.n863 1.0245
R5638 GNDA.n859 GNDA.n756 1.0245
R5639 GNDA.n858 GNDA.n760 1.0245
R5640 GNDA.n764 GNDA.n762 1.0245
R5641 GNDA.n853 GNDA.n852 1.0245
R5642 GNDA.n848 GNDA.n765 1.0245
R5643 GNDA.n847 GNDA.n769 1.0245
R5644 GNDA.n992 GNDA.n991 1.0245
R5645 GNDA.n988 GNDA.n987 1.0245
R5646 GNDA.n984 GNDA.n961 1.0245
R5647 GNDA.n983 GNDA.n962 1.0245
R5648 GNDA.n979 GNDA.n978 1.0245
R5649 GNDA.n975 GNDA.n974 1.0245
R5650 GNDA.n971 GNDA.n966 1.0245
R5651 GNDA.n970 GNDA.n695 1.0245
R5652 GNDA.n1048 GNDA.n1047 1.0245
R5653 GNDA.n1193 GNDA.n1079 1.0245
R5654 GNDA.n1083 GNDA.n1081 1.0245
R5655 GNDA.n1188 GNDA.n1187 1.0245
R5656 GNDA.n1183 GNDA.n1084 1.0245
R5657 GNDA.n1182 GNDA.n1088 1.0245
R5658 GNDA.n1092 GNDA.n1090 1.0245
R5659 GNDA.n1177 GNDA.n1176 1.0245
R5660 GNDA.n1172 GNDA.n1093 1.0245
R5661 GNDA.n1171 GNDA.n1097 1.0245
R5662 GNDA.n1488 GNDA.n1487 1.0245
R5663 GNDA.n1483 GNDA.n1414 1.0245
R5664 GNDA.n1482 GNDA.n1454 1.0245
R5665 GNDA.n1458 GNDA.n1456 1.0245
R5666 GNDA.n1477 GNDA.n1476 1.0245
R5667 GNDA.n1472 GNDA.n1459 1.0245
R5668 GNDA.n1471 GNDA.n1464 1.0245
R5669 GNDA.n1467 GNDA.n1466 1.0245
R5670 GNDA.n1544 GNDA.n1395 1.0245
R5671 GNDA.n1384 GNDA.n1271 1.0245
R5672 GNDA.n1275 GNDA.n1273 1.0245
R5673 GNDA.n1379 GNDA.n1378 1.0245
R5674 GNDA.n1374 GNDA.n1276 1.0245
R5675 GNDA.n1373 GNDA.n1280 1.0245
R5676 GNDA.n1284 GNDA.n1282 1.0245
R5677 GNDA.n1368 GNDA.n1367 1.0245
R5678 GNDA.n1363 GNDA.n1285 1.0245
R5679 GNDA.n1362 GNDA.n1289 1.0245
R5680 GNDA.n2283 GNDA.n284 1.0245
R5681 GNDA.n288 GNDA.n286 1.0245
R5682 GNDA.n2278 GNDA.n2277 1.0245
R5683 GNDA.n2273 GNDA.n289 1.0245
R5684 GNDA.n2272 GNDA.n293 1.0245
R5685 GNDA.n297 GNDA.n295 1.0245
R5686 GNDA.n2267 GNDA.n2266 1.0245
R5687 GNDA.n2262 GNDA.n298 1.0245
R5688 GNDA.n2261 GNDA.n302 1.0245
R5689 GNDA.n1658 GNDA.n1656 0.563
R5690 GNDA.n1662 GNDA.n1660 0.563
R5691 GNDA.n1664 GNDA.n1662 0.563
R5692 GNDA.n1666 GNDA.n1664 0.563
R5693 GNDA.n1670 GNDA.n1668 0.563
R5694 GNDA.n1672 GNDA.n1670 0.563
R5695 GNDA.n17 GNDA.n15 0.563
R5696 GNDA.n19 GNDA.n17 0.563
R5697 GNDA.n21 GNDA.n19 0.563
R5698 GNDA.n23 GNDA.n21 0.563
R5699 GNDA.n394 GNDA.n36 0.563
R5700 GNDA.n396 GNDA.n394 0.563
R5701 GNDA.n398 GNDA.n396 0.563
R5702 GNDA.n400 GNDA.n398 0.563
R5703 GNDA.n402 GNDA.n400 0.563
R5704 GNDA.n404 GNDA.n402 0.563
R5705 GNDA.n406 GNDA.n404 0.563
R5706 GNDA.n408 GNDA.n406 0.563
R5707 GNDA.n410 GNDA.n408 0.563
R5708 GNDA.n412 GNDA.n410 0.563
R5709 GNDA.n414 GNDA.n412 0.563
R5710 GNDA.n6 GNDA.n4 0.563
R5711 GNDA.n8 GNDA.n6 0.563
R5712 GNDA.n10 GNDA.n8 0.563
R5713 GNDA.n12 GNDA.n10 0.563
R5714 GNDA.n2492 GNDA.n1 0.53175
R5715 GNDA.n477 GNDA.n476 0.5005
R5716 GNDA.n2478 GNDA.n2476 0.5005
R5717 GNDA.n2458 GNDA.t0 0.467591
R5718 GNDA.n346 GNDA.t36 0.467591
R5719 GNDA.n552 GNDA.n551 0.41175
R5720 GNDA.n553 GNDA.n552 0.311875
R5721 GNDA.n2480 GNDA.n36 0.28175
R5722 GNDA.n1653 GNDA.n1634 0.276625
R5723 GNDA.n415 GNDA.n414 0.2505
R5724 GNDA.n1673 GNDA.n1653 0.22375
R5725 GNDA GNDA.n2423 0.129793
R5726 GNDA.n2138 GNDA 0.129793
R5727 GNDA.n2166 GNDA 0.129793
R5728 GNDA.n1674 GNDA.n1673 0.100375
R5729 GNDA.n554 GNDA.n553 0.076875
R5730 GNDA.n1216 GNDA.n256 0.0479074
R5731 GNDA.n1231 GNDA 0.0479074
R5732 GNDA.n650 GNDA.n581 0.0479074
R5733 GNDA.n1919 GNDA 0.0479074
R5734 GNDA.n629 GNDA.n628 0.0479074
R5735 GNDA GNDA.n642 0.0479074
R5736 GNDA.n726 GNDA.n724 0.0479074
R5737 GNDA.n945 GNDA 0.0479074
R5738 GNDA.n542 GNDA.n538 0.0479074
R5739 GNDA GNDA.n1067 0.0479074
R5740 GNDA.n182 GNDA.n181 0.0479074
R5741 GNDA GNDA.n272 0.0479074
R5742 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t15 354.854
R5743 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t30 346.8
R5744 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n4 339.522
R5745 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 339.522
R5746 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n9 335.022
R5747 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t1 275.909
R5748 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 227.909
R5749 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 222.034
R5750 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t31 184.097
R5751 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t14 184.097
R5752 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t27 184.097
R5753 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t19 184.097
R5754 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 166.05
R5755 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 166.05
R5756 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t7 48.0005
R5757 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t6 48.0005
R5758 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t2 48.0005
R5759 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t10 48.0005
R5760 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t8 39.4005
R5761 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t5 39.4005
R5762 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t9 39.4005
R5763 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t3 39.4005
R5764 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t0 39.4005
R5765 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t4 39.4005
R5766 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n2 33.1711
R5767 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n0 5.6255
R5768 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 5.28175
R5769 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R5770 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t29 4.8295
R5771 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t25 4.8295
R5772 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t35 4.8295
R5773 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t33 4.8295
R5774 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t17 4.8295
R5775 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t28 4.8295
R5776 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n7 4.5005
R5777 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t11 4.5005
R5778 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t32 4.5005
R5779 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t34 4.5005
R5780 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t21 4.5005
R5781 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t12 4.5005
R5782 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t16 4.5005
R5783 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t26 4.5005
R5784 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t22 4.5005
R5785 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.5005
R5786 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.5005
R5787 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t13 4.5005
R5788 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t18 4.5005
R5789 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t36 4.5005
R5790 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.8075
R5791 bgr_0.cap_res1.t20 bgr_0.cap_res1.t17 178.633
R5792 bgr_0.cap_res1.t14 bgr_0.cap_res1.t0 0.1603
R5793 bgr_0.cap_res1.t10 bgr_0.cap_res1.t6 0.1603
R5794 bgr_0.cap_res1.t9 bgr_0.cap_res1.t15 0.1603
R5795 bgr_0.cap_res1.t7 bgr_0.cap_res1.t3 0.1603
R5796 bgr_0.cap_res1.t16 bgr_0.cap_res1.t1 0.1603
R5797 bgr_0.cap_res1.t12 bgr_0.cap_res1.t8 0.1603
R5798 bgr_0.cap_res1.t2 bgr_0.cap_res1.t5 0.1603
R5799 bgr_0.cap_res1.t19 bgr_0.cap_res1.t13 0.1603
R5800 bgr_0.cap_res1.n1 bgr_0.cap_res1.t4 0.159278
R5801 bgr_0.cap_res1.n2 bgr_0.cap_res1.t18 0.159278
R5802 bgr_0.cap_res1.n3 bgr_0.cap_res1.t11 0.159278
R5803 bgr_0.cap_res1.n3 bgr_0.cap_res1.t14 0.1368
R5804 bgr_0.cap_res1.n3 bgr_0.cap_res1.t10 0.1368
R5805 bgr_0.cap_res1.n2 bgr_0.cap_res1.t9 0.1368
R5806 bgr_0.cap_res1.n2 bgr_0.cap_res1.t7 0.1368
R5807 bgr_0.cap_res1.n1 bgr_0.cap_res1.t16 0.1368
R5808 bgr_0.cap_res1.n1 bgr_0.cap_res1.t12 0.1368
R5809 bgr_0.cap_res1.n0 bgr_0.cap_res1.t2 0.1368
R5810 bgr_0.cap_res1.n0 bgr_0.cap_res1.t19 0.1368
R5811 bgr_0.cap_res1.t4 bgr_0.cap_res1.n0 0.00152174
R5812 bgr_0.cap_res1.t18 bgr_0.cap_res1.n1 0.00152174
R5813 bgr_0.cap_res1.t11 bgr_0.cap_res1.n2 0.00152174
R5814 bgr_0.cap_res1.t17 bgr_0.cap_res1.n3 0.00152174
R5815 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.n7 114.719
R5816 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5817 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5818 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.n8 114.156
R5819 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5820 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5821 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5822 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5823 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5824 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5825 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5826 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5827 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5828 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5829 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5830 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5831 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5832 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5833 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5834 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5835 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5836 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5837 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5838 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t17 16.0005
R5839 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5840 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5841 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5842 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5843 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5844 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5845 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5846 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5847 two_stage_opamp_dummy_magic_0.VD2.t8 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5848 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5849 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5850 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5851 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5852 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5853 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5854 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 0.563
R5855 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5856 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.n5 145.989
R5857 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n6 145.989
R5858 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n11 145.427
R5859 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n9 145.427
R5860 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n7 145.427
R5861 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n14 140.927
R5862 two_stage_opamp_dummy_magic_0.VOUT-.t6 two_stage_opamp_dummy_magic_0.VOUT-.n96 113.192
R5863 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n0 95.7303
R5864 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n3 94.6053
R5865 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n1 94.6053
R5866 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.n15 20.688
R5867 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.n94 11.7059
R5868 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n95 10.438
R5869 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t9 6.56717
R5870 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t11 6.56717
R5871 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t1 6.56717
R5872 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t12 6.56717
R5873 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t2 6.56717
R5874 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t15 6.56717
R5875 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t10 6.56717
R5876 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t4 6.56717
R5877 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.t13 6.56717
R5878 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.t18 6.56717
R5879 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t17 6.56717
R5880 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t0 6.56717
R5881 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t85 4.8295
R5882 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t131 4.8295
R5883 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t31 4.8295
R5884 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t62 4.8295
R5885 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t114 4.8295
R5886 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t40 4.8295
R5887 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t34 4.8295
R5888 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t136 4.8295
R5889 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t70 4.8295
R5890 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t36 4.8295
R5891 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.t95 4.8295
R5892 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t66 4.8295
R5893 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.t55 4.8295
R5894 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t29 4.8295
R5895 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.t91 4.8295
R5896 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t58 4.8295
R5897 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.t49 4.8295
R5898 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t20 4.8295
R5899 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.t148 4.8295
R5900 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t122 4.8295
R5901 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.t44 4.8295
R5902 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t152 4.8295
R5903 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.t142 4.8295
R5904 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t116 4.8295
R5905 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t108 4.8295
R5906 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t28 4.8295
R5907 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t24 4.8295
R5908 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t129 4.8295
R5909 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t61 4.8295
R5910 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t32 4.8295
R5911 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t100 4.8295
R5912 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t71 4.8295
R5913 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t69 4.8295
R5914 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t35 4.8295
R5915 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t77 4.8295
R5916 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t26 4.8154
R5917 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t59 4.8154
R5918 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t37 4.8154
R5919 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t81 4.8154
R5920 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t132 4.806
R5921 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t115 4.806
R5922 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t146 4.806
R5923 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.t46 4.806
R5924 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t87 4.806
R5925 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t65 4.806
R5926 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t102 4.806
R5927 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t134 4.806
R5928 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t120 4.806
R5929 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t155 4.806
R5930 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t48 4.806
R5931 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t92 4.806
R5932 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t42 4.806
R5933 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t130 4.806
R5934 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t84 4.806
R5935 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t125 4.806
R5936 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t74 4.806
R5937 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t23 4.806
R5938 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t64 4.806
R5939 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t150 4.806
R5940 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.t96 4.5005
R5941 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t57 4.5005
R5942 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t104 4.5005
R5943 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.t73 4.5005
R5944 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t138 4.5005
R5945 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.t107 4.5005
R5946 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t41 4.5005
R5947 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.t143 4.5005
R5948 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t21 4.5005
R5949 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.t126 4.5005
R5950 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t119 4.5005
R5951 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t82 4.5005
R5952 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t97 4.5005
R5953 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t63 4.5005
R5954 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t27 4.5005
R5955 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t45 4.5005
R5956 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.t144 4.5005
R5957 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t112 4.5005
R5958 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t76 4.5005
R5959 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t93 4.5005
R5960 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.t56 4.5005
R5961 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t19 4.5005
R5962 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t52 4.5005
R5963 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.t156 4.5005
R5964 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t121 4.5005
R5965 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t89 4.5005
R5966 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.t50 4.5005
R5967 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t151 4.5005
R5968 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.t43 4.5005
R5969 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.t145 4.5005
R5970 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t118 4.5005
R5971 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.t141 4.5005
R5972 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.t111 4.5005
R5973 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t80 4.5005
R5974 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.t39 4.5005
R5975 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.t139 4.5005
R5976 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t109 4.5005
R5977 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.t135 4.5005
R5978 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.t103 4.5005
R5979 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t72 4.5005
R5980 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.t99 4.5005
R5981 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.t68 4.5005
R5982 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t33 4.5005
R5983 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.t133 4.5005
R5984 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.t98 4.5005
R5985 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t67 4.5005
R5986 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.t94 4.5005
R5987 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.t60 4.5005
R5988 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t30 4.5005
R5989 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.t101 4.5005
R5990 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t149 4.5005
R5991 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t88 4.5005
R5992 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t51 4.5005
R5993 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t137 4.5005
R5994 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t106 4.5005
R5995 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t75 4.5005
R5996 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t25 4.5005
R5997 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t128 4.5005
R5998 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t90 4.5005
R5999 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t54 4.5005
R6000 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t140 4.5005
R6001 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.t110 4.5005
R6002 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t79 4.5005
R6003 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t113 4.5005
R6004 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.t78 4.5005
R6005 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t38 4.5005
R6006 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t147 4.5005
R6007 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.t117 4.5005
R6008 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t83 4.5005
R6009 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t47 4.5005
R6010 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.t153 4.5005
R6011 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t123 4.5005
R6012 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t154 4.5005
R6013 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.t124 4.5005
R6014 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t86 4.5005
R6015 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.t105 4.5005
R6016 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.t53 4.5005
R6017 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.t22 4.5005
R6018 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t127 4.5005
R6019 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n13 4.5005
R6020 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t14 3.42907
R6021 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t8 3.42907
R6022 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t5 3.42907
R6023 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t16 3.42907
R6024 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t7 3.42907
R6025 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t3 3.42907
R6026 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n4 2.03175
R6027 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n2 1.1255
R6028 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n8 0.563
R6029 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n10 0.563
R6030 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.n12 0.563
R6031 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.n42 0.3295
R6032 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.n44 0.3295
R6033 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.n46 0.3295
R6034 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.n48 0.3295
R6035 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.n50 0.3295
R6036 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.n52 0.3295
R6037 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.n53 0.3295
R6038 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.n54 0.3295
R6039 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.n55 0.3295
R6040 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.n56 0.3295
R6041 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n57 0.3295
R6042 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.n58 0.3295
R6043 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.n59 0.3295
R6044 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.n60 0.3295
R6045 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n61 0.3295
R6046 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n62 0.3295
R6047 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n64 0.3295
R6048 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n65 0.3295
R6049 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.n67 0.3295
R6050 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.n68 0.3295
R6051 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.n70 0.3295
R6052 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.n71 0.3295
R6053 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.n73 0.3295
R6054 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.n74 0.3295
R6055 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.n76 0.3295
R6056 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.n77 0.3295
R6057 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.n79 0.3295
R6058 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.n80 0.3295
R6059 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.n82 0.3295
R6060 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.n83 0.3295
R6061 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n85 0.3295
R6062 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n86 0.3295
R6063 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n88 0.3295
R6064 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n89 0.3295
R6065 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.n16 0.3295
R6066 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.n18 0.3295
R6067 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.n19 0.3295
R6068 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.n20 0.3295
R6069 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.n21 0.3295
R6070 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.n22 0.3295
R6071 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.n23 0.3295
R6072 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.n24 0.3295
R6073 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.n25 0.3295
R6074 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.n26 0.3295
R6075 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n27 0.3295
R6076 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n28 0.3295
R6077 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n30 0.3295
R6078 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n31 0.3295
R6079 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n33 0.3295
R6080 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n34 0.3295
R6081 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n36 0.3295
R6082 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n37 0.3295
R6083 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n39 0.3295
R6084 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n40 0.3295
R6085 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.n93 0.3295
R6086 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.n92 0.3295
R6087 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.n91 0.3295
R6088 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.n45 0.306
R6089 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n47 0.306
R6090 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.n49 0.306
R6091 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.n51 0.306
R6092 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.n43 0.2825
R6093 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.n63 0.2825
R6094 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.n66 0.2825
R6095 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.n69 0.2825
R6096 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.n72 0.2825
R6097 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.n75 0.2825
R6098 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.n78 0.2825
R6099 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.n81 0.2825
R6100 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n84 0.2825
R6101 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n87 0.2825
R6102 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.n17 0.2825
R6103 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.n29 0.2825
R6104 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.n32 0.2825
R6105 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n35 0.2825
R6106 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n38 0.2825
R6107 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.n41 0.2825
R6108 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.n90 0.2825
R6109 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t0 49.083
R6110 two_stage_opamp_dummy_magic_0.cap_res_X two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.922875
R6111 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1603
R6112 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.1603
R6113 two_stage_opamp_dummy_magic_0.cap_res_X.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R6114 two_stage_opamp_dummy_magic_0.cap_res_X.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R6115 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.1603
R6116 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1603
R6117 two_stage_opamp_dummy_magic_0.cap_res_X.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R6118 two_stage_opamp_dummy_magic_0.cap_res_X.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.1603
R6119 two_stage_opamp_dummy_magic_0.cap_res_X.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R6120 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.1603
R6121 two_stage_opamp_dummy_magic_0.cap_res_X.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.1603
R6122 two_stage_opamp_dummy_magic_0.cap_res_X.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R6123 two_stage_opamp_dummy_magic_0.cap_res_X.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R6124 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1603
R6125 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.1603
R6126 two_stage_opamp_dummy_magic_0.cap_res_X.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1603
R6127 two_stage_opamp_dummy_magic_0.cap_res_X.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.1603
R6128 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R6129 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.1603
R6130 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1603
R6131 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.1603
R6132 two_stage_opamp_dummy_magic_0.cap_res_X.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.1603
R6133 two_stage_opamp_dummy_magic_0.cap_res_X.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.1603
R6134 two_stage_opamp_dummy_magic_0.cap_res_X.t3 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.1603
R6135 two_stage_opamp_dummy_magic_0.cap_res_X.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1603
R6136 two_stage_opamp_dummy_magic_0.cap_res_X.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1603
R6137 two_stage_opamp_dummy_magic_0.cap_res_X.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.1603
R6138 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.1603
R6139 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1603
R6140 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.1603
R6141 two_stage_opamp_dummy_magic_0.cap_res_X.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1603
R6142 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.1603
R6143 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R6144 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1603
R6145 two_stage_opamp_dummy_magic_0.cap_res_X.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R6146 two_stage_opamp_dummy_magic_0.cap_res_X.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.1603
R6147 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1603
R6148 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1603
R6149 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1603
R6150 two_stage_opamp_dummy_magic_0.cap_res_X.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1603
R6151 two_stage_opamp_dummy_magic_0.cap_res_X.t17 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1603
R6152 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1603
R6153 two_stage_opamp_dummy_magic_0.cap_res_X.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.1603
R6154 two_stage_opamp_dummy_magic_0.cap_res_X.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R6155 two_stage_opamp_dummy_magic_0.cap_res_X.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1603
R6156 two_stage_opamp_dummy_magic_0.cap_res_X.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1603
R6157 two_stage_opamp_dummy_magic_0.cap_res_X.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1603
R6158 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R6159 two_stage_opamp_dummy_magic_0.cap_res_X.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.1603
R6160 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.1603
R6161 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R6162 two_stage_opamp_dummy_magic_0.cap_res_X.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1603
R6163 two_stage_opamp_dummy_magic_0.cap_res_X.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R6164 two_stage_opamp_dummy_magic_0.cap_res_X.t14 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1603
R6165 two_stage_opamp_dummy_magic_0.cap_res_X.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R6166 two_stage_opamp_dummy_magic_0.cap_res_X.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.1603
R6167 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R6168 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.1603
R6169 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.159278
R6170 two_stage_opamp_dummy_magic_0.cap_res_X.t47 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R6171 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R6172 two_stage_opamp_dummy_magic_0.cap_res_X.t40 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R6173 two_stage_opamp_dummy_magic_0.cap_res_X.t4 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R6174 two_stage_opamp_dummy_magic_0.cap_res_X.t33 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R6175 two_stage_opamp_dummy_magic_0.cap_res_X.t135 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R6176 two_stage_opamp_dummy_magic_0.cap_res_X.t97 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R6177 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R6178 two_stage_opamp_dummy_magic_0.cap_res_X.t89 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R6179 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R6180 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.159278
R6181 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.159278
R6182 two_stage_opamp_dummy_magic_0.cap_res_X.t12 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.159278
R6183 two_stage_opamp_dummy_magic_0.cap_res_X.t107 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.159278
R6184 two_stage_opamp_dummy_magic_0.cap_res_X.t1 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.159278
R6185 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.159278
R6186 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.159278
R6187 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.159278
R6188 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.159278
R6189 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.159278
R6190 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.159278
R6191 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.159278
R6192 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.159278
R6193 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.159278
R6194 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.159278
R6195 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.159278
R6196 two_stage_opamp_dummy_magic_0.cap_res_X.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.137822
R6197 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.1368
R6198 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1368
R6199 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1368
R6200 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t6 0.1368
R6201 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R6202 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1368
R6203 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1368
R6204 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1368
R6205 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R6206 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1368
R6207 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1368
R6208 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1368
R6209 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R6210 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R6211 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1368
R6212 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1368
R6213 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.1368
R6214 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R6215 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.1368
R6216 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.1368
R6217 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.1368
R6218 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.1368
R6219 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1368
R6220 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.1368
R6221 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.1368
R6222 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1368
R6223 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.1368
R6224 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R6225 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.1368
R6226 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1368
R6227 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.1368
R6228 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.114322
R6229 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R6230 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R6231 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R6232 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.1133
R6233 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.1133
R6234 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.1133
R6235 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.1133
R6236 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.1133
R6237 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.1133
R6238 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R6239 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R6240 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R6241 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R6242 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R6243 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R6244 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R6245 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R6246 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R6247 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R6248 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.00152174
R6249 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.00152174
R6250 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.00152174
R6251 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R6252 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.00152174
R6253 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R6254 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.00152174
R6255 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.00152174
R6256 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.00152174
R6257 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.00152174
R6258 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.00152174
R6259 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.00152174
R6260 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.00152174
R6261 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.00152174
R6262 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.00152174
R6263 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.00152174
R6264 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.00152174
R6265 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.00152174
R6266 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.00152174
R6267 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.00152174
R6268 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R6269 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R6270 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.00152174
R6271 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.00152174
R6272 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.00152174
R6273 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.00152174
R6274 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.00152174
R6275 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.00152174
R6276 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.00152174
R6277 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.00152174
R6278 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.00152174
R6279 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R6280 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.00152174
R6281 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.00152174
R6282 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.00152174
R6283 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R6284 bgr_0.Vbe2.n145 bgr_0.Vbe2.n144 413.99
R6285 bgr_0.Vbe2.n136 bgr_0.Vbe2.t8 162.458
R6286 bgr_0.Vbe2.n146 bgr_0.Vbe2.n145 84.0884
R6287 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 83.5719
R6288 bgr_0.Vbe2.n55 bgr_0.Vbe2.n48 83.5719
R6289 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 83.5719
R6290 bgr_0.Vbe2.n127 bgr_0.Vbe2.n6 83.5719
R6291 bgr_0.Vbe2.n122 bgr_0.Vbe2.n7 83.5719
R6292 bgr_0.Vbe2.n45 bgr_0.Vbe2.n44 83.5719
R6293 bgr_0.Vbe2.n43 bgr_0.Vbe2.n42 83.5719
R6294 bgr_0.Vbe2.n41 bgr_0.Vbe2.n40 83.5719
R6295 bgr_0.Vbe2.n78 bgr_0.Vbe2.n77 83.5719
R6296 bgr_0.Vbe2.n76 bgr_0.Vbe2.n75 83.5719
R6297 bgr_0.Vbe2.n27 bgr_0.Vbe2.n26 83.5719
R6298 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 83.5719
R6299 bgr_0.Vbe2.n22 bgr_0.Vbe2.n20 83.5719
R6300 bgr_0.Vbe2.n91 bgr_0.Vbe2.n19 83.5719
R6301 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 83.5719
R6302 bgr_0.Vbe2.n17 bgr_0.Vbe2.n16 83.5719
R6303 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 83.5719
R6304 bgr_0.Vbe2.n112 bgr_0.Vbe2.n111 83.5719
R6305 bgr_0.Vbe2.n110 bgr_0.Vbe2.n109 83.5719
R6306 bgr_0.Vbe2.n143 bgr_0.Vbe2.n1 83.5719
R6307 bgr_0.Vbe2.n142 bgr_0.Vbe2.n0 83.5719
R6308 bgr_0.Vbe2.n141 bgr_0.Vbe2.n140 83.5719
R6309 bgr_0.Vbe2.n132 bgr_0.Vbe2.n4 83.5719
R6310 bgr_0.Vbe2.n72 bgr_0.Vbe2.n26 73.8495
R6311 bgr_0.Vbe2.n59 bgr_0.Vbe2.n58 73.3165
R6312 bgr_0.Vbe2.n129 bgr_0.Vbe2.n6 73.3165
R6313 bgr_0.Vbe2.n44 bgr_0.Vbe2.n36 73.3165
R6314 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 73.3165
R6315 bgr_0.Vbe2.n98 bgr_0.Vbe2.n97 73.3165
R6316 bgr_0.Vbe2.n115 bgr_0.Vbe2.n114 73.3165
R6317 bgr_0.Vbe2.n54 bgr_0.Vbe2.n49 73.19
R6318 bgr_0.Vbe2.n41 bgr_0.Vbe2.n39 73.19
R6319 bgr_0.Vbe2.n77 bgr_0.Vbe2.n23 73.19
R6320 bgr_0.Vbe2.n93 bgr_0.Vbe2.n19 73.19
R6321 bgr_0.Vbe2.n110 bgr_0.Vbe2.n13 73.19
R6322 bgr_0.Vbe2.n133 bgr_0.Vbe2.n132 73.19
R6323 bgr_0.Vbe2.n123 bgr_0.Vbe2.t4 65.0299
R6324 bgr_0.Vbe2.t6 bgr_0.Vbe2.n14 65.0299
R6325 bgr_0.Vbe2.n59 bgr_0.Vbe2.n55 26.074
R6326 bgr_0.Vbe2.n122 bgr_0.Vbe2.n6 26.074
R6327 bgr_0.Vbe2.n44 bgr_0.Vbe2.n43 26.074
R6328 bgr_0.Vbe2.n76 bgr_0.Vbe2.n26 26.074
R6329 bgr_0.Vbe2.n85 bgr_0.Vbe2.n22 26.074
R6330 bgr_0.Vbe2.n98 bgr_0.Vbe2.n17 26.074
R6331 bgr_0.Vbe2.n114 bgr_0.Vbe2.n112 26.074
R6332 bgr_0.Vbe2.n142 bgr_0.Vbe2.n141 26.074
R6333 bgr_0.Vbe2.n143 bgr_0.Vbe2.n142 26.074
R6334 bgr_0.Vbe2.n145 bgr_0.Vbe2.n143 26.074
R6335 bgr_0.Vbe2.t0 bgr_0.Vbe2.n54 25.7843
R6336 bgr_0.Vbe2.t2 bgr_0.Vbe2.n41 25.7843
R6337 bgr_0.Vbe2.n77 bgr_0.Vbe2.t3 25.7843
R6338 bgr_0.Vbe2.t1 bgr_0.Vbe2.n19 25.7843
R6339 bgr_0.Vbe2.t5 bgr_0.Vbe2.n110 25.7843
R6340 bgr_0.Vbe2.n132 bgr_0.Vbe2.t7 25.7843
R6341 bgr_0.Vbe2.n116 bgr_0.Vbe2.n104 9.3005
R6342 bgr_0.Vbe2.n104 bgr_0.Vbe2.n11 9.3005
R6343 bgr_0.Vbe2.n104 bgr_0.Vbe2.n12 9.3005
R6344 bgr_0.Vbe2.n120 bgr_0.Vbe2.n104 9.3005
R6345 bgr_0.Vbe2.n106 bgr_0.Vbe2.n11 9.3005
R6346 bgr_0.Vbe2.n106 bgr_0.Vbe2.n12 9.3005
R6347 bgr_0.Vbe2.n106 bgr_0.Vbe2.n9 9.3005
R6348 bgr_0.Vbe2.n120 bgr_0.Vbe2.n106 9.3005
R6349 bgr_0.Vbe2.n121 bgr_0.Vbe2.n11 9.3005
R6350 bgr_0.Vbe2.n121 bgr_0.Vbe2.n10 9.3005
R6351 bgr_0.Vbe2.n121 bgr_0.Vbe2.n12 9.3005
R6352 bgr_0.Vbe2.n121 bgr_0.Vbe2.n9 9.3005
R6353 bgr_0.Vbe2.n121 bgr_0.Vbe2.n120 9.3005
R6354 bgr_0.Vbe2.n120 bgr_0.Vbe2.n108 9.3005
R6355 bgr_0.Vbe2.n108 bgr_0.Vbe2.n9 9.3005
R6356 bgr_0.Vbe2.n108 bgr_0.Vbe2.n12 9.3005
R6357 bgr_0.Vbe2.n108 bgr_0.Vbe2.n10 9.3005
R6358 bgr_0.Vbe2.n120 bgr_0.Vbe2.n103 9.3005
R6359 bgr_0.Vbe2.n103 bgr_0.Vbe2.n9 9.3005
R6360 bgr_0.Vbe2.n103 bgr_0.Vbe2.n12 9.3005
R6361 bgr_0.Vbe2.n103 bgr_0.Vbe2.n10 9.3005
R6362 bgr_0.Vbe2.n116 bgr_0.Vbe2.n103 9.3005
R6363 bgr_0.Vbe2.n119 bgr_0.Vbe2.n11 9.3005
R6364 bgr_0.Vbe2.n119 bgr_0.Vbe2.n10 9.3005
R6365 bgr_0.Vbe2.n119 bgr_0.Vbe2.n12 9.3005
R6366 bgr_0.Vbe2.n120 bgr_0.Vbe2.n119 9.3005
R6367 bgr_0.Vbe2.n69 bgr_0.Vbe2.n68 9.3005
R6368 bgr_0.Vbe2.n68 bgr_0.Vbe2.n67 9.3005
R6369 bgr_0.Vbe2.n68 bgr_0.Vbe2.n29 9.3005
R6370 bgr_0.Vbe2.n68 bgr_0.Vbe2.n30 9.3005
R6371 bgr_0.Vbe2.n67 bgr_0.Vbe2.n65 9.3005
R6372 bgr_0.Vbe2.n65 bgr_0.Vbe2.n29 9.3005
R6373 bgr_0.Vbe2.n65 bgr_0.Vbe2.n31 9.3005
R6374 bgr_0.Vbe2.n65 bgr_0.Vbe2.n30 9.3005
R6375 bgr_0.Vbe2.n67 bgr_0.Vbe2.n64 9.3005
R6376 bgr_0.Vbe2.n64 bgr_0.Vbe2.n32 9.3005
R6377 bgr_0.Vbe2.n64 bgr_0.Vbe2.n29 9.3005
R6378 bgr_0.Vbe2.n64 bgr_0.Vbe2.n31 9.3005
R6379 bgr_0.Vbe2.n64 bgr_0.Vbe2.n30 9.3005
R6380 bgr_0.Vbe2.n33 bgr_0.Vbe2.n30 9.3005
R6381 bgr_0.Vbe2.n33 bgr_0.Vbe2.n31 9.3005
R6382 bgr_0.Vbe2.n33 bgr_0.Vbe2.n29 9.3005
R6383 bgr_0.Vbe2.n33 bgr_0.Vbe2.n32 9.3005
R6384 bgr_0.Vbe2.n70 bgr_0.Vbe2.n30 9.3005
R6385 bgr_0.Vbe2.n70 bgr_0.Vbe2.n31 9.3005
R6386 bgr_0.Vbe2.n70 bgr_0.Vbe2.n29 9.3005
R6387 bgr_0.Vbe2.n70 bgr_0.Vbe2.n32 9.3005
R6388 bgr_0.Vbe2.n70 bgr_0.Vbe2.n69 9.3005
R6389 bgr_0.Vbe2.n67 bgr_0.Vbe2.n66 9.3005
R6390 bgr_0.Vbe2.n66 bgr_0.Vbe2.n32 9.3005
R6391 bgr_0.Vbe2.n66 bgr_0.Vbe2.n29 9.3005
R6392 bgr_0.Vbe2.n66 bgr_0.Vbe2.n30 9.3005
R6393 bgr_0.Vbe2.n118 bgr_0.Vbe2.n9 4.64654
R6394 bgr_0.Vbe2.n105 bgr_0.Vbe2.n10 4.64654
R6395 bgr_0.Vbe2.n116 bgr_0.Vbe2.n8 4.64654
R6396 bgr_0.Vbe2.n107 bgr_0.Vbe2.n11 4.64654
R6397 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 4.64654
R6398 bgr_0.Vbe2.n37 bgr_0.Vbe2.n31 4.64654
R6399 bgr_0.Vbe2.n38 bgr_0.Vbe2.n32 4.64654
R6400 bgr_0.Vbe2.n69 bgr_0.Vbe2.n35 4.64654
R6401 bgr_0.Vbe2.n67 bgr_0.Vbe2.n28 4.64654
R6402 bgr_0.Vbe2.n69 bgr_0.Vbe2.n34 4.64654
R6403 bgr_0.Vbe2.n49 bgr_0.Vbe2.n3 2.36206
R6404 bgr_0.Vbe2.n81 bgr_0.Vbe2.n23 2.36206
R6405 bgr_0.Vbe2.n94 bgr_0.Vbe2.n93 2.36206
R6406 bgr_0.Vbe2.n133 bgr_0.Vbe2.n131 2.36206
R6407 bgr_0.Vbe2.n58 bgr_0.Vbe2.n56 2.19742
R6408 bgr_0.Vbe2.n130 bgr_0.Vbe2.n129 2.19742
R6409 bgr_0.Vbe2.n84 bgr_0.Vbe2.n82 2.19742
R6410 bgr_0.Vbe2.n97 bgr_0.Vbe2.n95 2.19742
R6411 bgr_0.Vbe2.n123 bgr_0.Vbe2.n7 1.56363
R6412 bgr_0.Vbe2.n16 bgr_0.Vbe2.n14 1.56363
R6413 bgr_0.Vbe2.n96 bgr_0.Vbe2.n15 1.5505
R6414 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 1.5505
R6415 bgr_0.Vbe2.n83 bgr_0.Vbe2.n21 1.5505
R6416 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 1.5505
R6417 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 1.5505
R6418 bgr_0.Vbe2.n92 bgr_0.Vbe2.n18 1.5505
R6419 bgr_0.Vbe2.n74 bgr_0.Vbe2.n73 1.5505
R6420 bgr_0.Vbe2.n80 bgr_0.Vbe2.n79 1.5505
R6421 bgr_0.Vbe2.n25 bgr_0.Vbe2.n24 1.5505
R6422 bgr_0.Vbe2.n128 bgr_0.Vbe2.n5 1.5505
R6423 bgr_0.Vbe2.n126 bgr_0.Vbe2.n125 1.5505
R6424 bgr_0.Vbe2.n57 bgr_0.Vbe2.n47 1.5505
R6425 bgr_0.Vbe2.n62 bgr_0.Vbe2.n61 1.5505
R6426 bgr_0.Vbe2.n52 bgr_0.Vbe2.n46 1.5505
R6427 bgr_0.Vbe2.n51 bgr_0.Vbe2.n50 1.5505
R6428 bgr_0.Vbe2.n147 bgr_0.Vbe2.n146 1.5505
R6429 bgr_0.Vbe2.n149 bgr_0.Vbe2.n148 1.5505
R6430 bgr_0.Vbe2.n139 bgr_0.Vbe2.n2 1.5505
R6431 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 1.5505
R6432 bgr_0.Vbe2.n135 bgr_0.Vbe2.n134 1.5505
R6433 bgr_0.Vbe2.n53 bgr_0.Vbe2.n51 1.25468
R6434 bgr_0.Vbe2.n40 bgr_0.Vbe2.n31 1.25468
R6435 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 1.25468
R6436 bgr_0.Vbe2.n92 bgr_0.Vbe2.n91 1.25468
R6437 bgr_0.Vbe2.n109 bgr_0.Vbe2.n9 1.25468
R6438 bgr_0.Vbe2.n134 bgr_0.Vbe2.n4 1.25468
R6439 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 1.19225
R6440 bgr_0.Vbe2.n129 bgr_0.Vbe2.n128 1.19225
R6441 bgr_0.Vbe2.n67 bgr_0.Vbe2.n36 1.19225
R6442 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 1.19225
R6443 bgr_0.Vbe2.n97 bgr_0.Vbe2.n96 1.19225
R6444 bgr_0.Vbe2.n115 bgr_0.Vbe2.n11 1.19225
R6445 bgr_0.Vbe2.n146 bgr_0.Vbe2.n1 1.14402
R6446 bgr_0.Vbe2.n52 bgr_0.Vbe2.n48 1.07024
R6447 bgr_0.Vbe2.n42 bgr_0.Vbe2.n29 1.07024
R6448 bgr_0.Vbe2.n75 bgr_0.Vbe2.n25 1.07024
R6449 bgr_0.Vbe2.n90 bgr_0.Vbe2.n20 1.07024
R6450 bgr_0.Vbe2.n111 bgr_0.Vbe2.n12 1.07024
R6451 bgr_0.Vbe2.n140 bgr_0.Vbe2.n138 1.07024
R6452 bgr_0.Vbe2.n51 bgr_0.Vbe2.n49 1.0237
R6453 bgr_0.Vbe2.n39 bgr_0.Vbe2.n31 1.0237
R6454 bgr_0.Vbe2.n79 bgr_0.Vbe2.n23 1.0237
R6455 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 1.0237
R6456 bgr_0.Vbe2.n13 bgr_0.Vbe2.n9 1.0237
R6457 bgr_0.Vbe2.n134 bgr_0.Vbe2.n133 1.0237
R6458 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 0.885803
R6459 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 0.885803
R6460 bgr_0.Vbe2.n45 bgr_0.Vbe2.n32 0.885803
R6461 bgr_0.Vbe2.n74 bgr_0.Vbe2.n27 0.885803
R6462 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 0.885803
R6463 bgr_0.Vbe2.n100 bgr_0.Vbe2.n99 0.885803
R6464 bgr_0.Vbe2.n113 bgr_0.Vbe2.n10 0.885803
R6465 bgr_0.Vbe2.n139 bgr_0.Vbe2.n0 0.885803
R6466 bgr_0.Vbe2.n39 bgr_0.Vbe2.n30 0.812055
R6467 bgr_0.Vbe2.n120 bgr_0.Vbe2.n13 0.812055
R6468 bgr_0.Vbe2.n61 bgr_0.Vbe2.n48 0.77514
R6469 bgr_0.Vbe2.n126 bgr_0.Vbe2.n7 0.77514
R6470 bgr_0.Vbe2.n42 bgr_0.Vbe2.n32 0.77514
R6471 bgr_0.Vbe2.n75 bgr_0.Vbe2.n74 0.77514
R6472 bgr_0.Vbe2.n87 bgr_0.Vbe2.n20 0.77514
R6473 bgr_0.Vbe2.n100 bgr_0.Vbe2.n16 0.77514
R6474 bgr_0.Vbe2.n111 bgr_0.Vbe2.n10 0.77514
R6475 bgr_0.Vbe2.n140 bgr_0.Vbe2.n139 0.77514
R6476 bgr_0.Vbe2.n60 bgr_0.Vbe2 0.756696
R6477 bgr_0.Vbe2 bgr_0.Vbe2.n127 0.756696
R6478 bgr_0.Vbe2 bgr_0.Vbe2.n45 0.756696
R6479 bgr_0.Vbe2 bgr_0.Vbe2.n27 0.756696
R6480 bgr_0.Vbe2.n86 bgr_0.Vbe2 0.756696
R6481 bgr_0.Vbe2.n99 bgr_0.Vbe2 0.756696
R6482 bgr_0.Vbe2.n113 bgr_0.Vbe2 0.756696
R6483 bgr_0.Vbe2 bgr_0.Vbe2.n0 0.756696
R6484 bgr_0.Vbe2.n73 bgr_0.Vbe2.n72 0.711459
R6485 bgr_0.Vbe2.n149 bgr_0.Vbe2.n1 0.701365
R6486 bgr_0.Vbe2.n69 bgr_0.Vbe2.n36 0.647417
R6487 bgr_0.Vbe2.n116 bgr_0.Vbe2.n115 0.647417
R6488 bgr_0.Vbe2.n53 bgr_0.Vbe2.n52 0.590702
R6489 bgr_0.Vbe2.n40 bgr_0.Vbe2.n29 0.590702
R6490 bgr_0.Vbe2.n78 bgr_0.Vbe2.n25 0.590702
R6491 bgr_0.Vbe2.n91 bgr_0.Vbe2.n90 0.590702
R6492 bgr_0.Vbe2.n109 bgr_0.Vbe2.n12 0.590702
R6493 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 0.590702
R6494 bgr_0.Vbe2.n72 bgr_0.Vbe2 0.576566
R6495 bgr_0.Vbe2.n102 bgr_0.Vbe2.n14 0.530034
R6496 bgr_0.Vbe2.n124 bgr_0.Vbe2.n123 0.530034
R6497 bgr_0.Vbe2.n55 bgr_0.Vbe2.t0 0.290206
R6498 bgr_0.Vbe2.t4 bgr_0.Vbe2.n122 0.290206
R6499 bgr_0.Vbe2.n43 bgr_0.Vbe2.t2 0.290206
R6500 bgr_0.Vbe2.t3 bgr_0.Vbe2.n76 0.290206
R6501 bgr_0.Vbe2.n22 bgr_0.Vbe2.t1 0.290206
R6502 bgr_0.Vbe2.n17 bgr_0.Vbe2.t6 0.290206
R6503 bgr_0.Vbe2.n112 bgr_0.Vbe2.t5 0.290206
R6504 bgr_0.Vbe2.n141 bgr_0.Vbe2.t7 0.290206
R6505 bgr_0.Vbe2.n57 bgr_0.Vbe2 0.203382
R6506 bgr_0.Vbe2.n128 bgr_0.Vbe2 0.203382
R6507 bgr_0.Vbe2.n67 bgr_0.Vbe2 0.203382
R6508 bgr_0.Vbe2.n83 bgr_0.Vbe2 0.203382
R6509 bgr_0.Vbe2.n96 bgr_0.Vbe2 0.203382
R6510 bgr_0.Vbe2 bgr_0.Vbe2.n11 0.203382
R6511 bgr_0.Vbe2 bgr_0.Vbe2.n149 0.203382
R6512 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.154071
R6513 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 0.154071
R6514 bgr_0.Vbe2.n131 bgr_0.Vbe2.n130 0.154071
R6515 bgr_0.Vbe2.n147 bgr_0.Vbe2.n3 0.154071
R6516 bgr_0.Vbe2.n124 bgr_0.Vbe2.n121 0.137464
R6517 bgr_0.Vbe2.n64 bgr_0.Vbe2.n63 0.137464
R6518 bgr_0.Vbe2.n103 bgr_0.Vbe2.n102 0.134964
R6519 bgr_0.Vbe2.n71 bgr_0.Vbe2.n70 0.134964
R6520 bgr_0.Vbe2.n56 bgr_0.Vbe2 0.0196071
R6521 bgr_0.Vbe2.n101 bgr_0.Vbe2.n15 0.0183571
R6522 bgr_0.Vbe2.n95 bgr_0.Vbe2.n15 0.0183571
R6523 bgr_0.Vbe2.n94 bgr_0.Vbe2.n18 0.0183571
R6524 bgr_0.Vbe2.n89 bgr_0.Vbe2.n18 0.0183571
R6525 bgr_0.Vbe2.n89 bgr_0.Vbe2.n88 0.0183571
R6526 bgr_0.Vbe2.n88 bgr_0.Vbe2.n21 0.0183571
R6527 bgr_0.Vbe2.n82 bgr_0.Vbe2.n21 0.0183571
R6528 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 0.0183571
R6529 bgr_0.Vbe2.n80 bgr_0.Vbe2.n24 0.0183571
R6530 bgr_0.Vbe2.n125 bgr_0.Vbe2.n5 0.0183571
R6531 bgr_0.Vbe2.n130 bgr_0.Vbe2.n5 0.0183571
R6532 bgr_0.Vbe2.n135 bgr_0.Vbe2.n131 0.0183571
R6533 bgr_0.Vbe2.n137 bgr_0.Vbe2.n135 0.0183571
R6534 bgr_0.Vbe2.n148 bgr_0.Vbe2.n2 0.0183571
R6535 bgr_0.Vbe2.n148 bgr_0.Vbe2.n147 0.0183571
R6536 bgr_0.Vbe2.n50 bgr_0.Vbe2.n3 0.0183571
R6537 bgr_0.Vbe2.n50 bgr_0.Vbe2.n46 0.0183571
R6538 bgr_0.Vbe2.n62 bgr_0.Vbe2.n47 0.0183571
R6539 bgr_0.Vbe2.n56 bgr_0.Vbe2.n47 0.0183571
R6540 bgr_0.Vbe2.n71 bgr_0.Vbe2.n24 0.0106786
R6541 bgr_0.Vbe2.n63 bgr_0.Vbe2.n46 0.0106786
R6542 bgr_0.Vbe2.n136 bgr_0.Vbe2.n2 0.00996429
R6543 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 0.00992001
R6544 bgr_0.Vbe2.n119 bgr_0.Vbe2.n117 0.00992001
R6545 bgr_0.Vbe2.n118 bgr_0.Vbe2.n104 0.00992001
R6546 bgr_0.Vbe2.n106 bgr_0.Vbe2.n105 0.00992001
R6547 bgr_0.Vbe2.n121 bgr_0.Vbe2.n8 0.00992001
R6548 bgr_0.Vbe2.n105 bgr_0.Vbe2.n104 0.00992001
R6549 bgr_0.Vbe2.n106 bgr_0.Vbe2.n8 0.00992001
R6550 bgr_0.Vbe2.n117 bgr_0.Vbe2.n108 0.00992001
R6551 bgr_0.Vbe2.n107 bgr_0.Vbe2.n103 0.00992001
R6552 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 0.00992001
R6553 bgr_0.Vbe2.n33 bgr_0.Vbe2.n28 0.00992001
R6554 bgr_0.Vbe2.n66 bgr_0.Vbe2.n34 0.00992001
R6555 bgr_0.Vbe2.n68 bgr_0.Vbe2.n37 0.00992001
R6556 bgr_0.Vbe2.n65 bgr_0.Vbe2.n38 0.00992001
R6557 bgr_0.Vbe2.n64 bgr_0.Vbe2.n35 0.00992001
R6558 bgr_0.Vbe2.n68 bgr_0.Vbe2.n38 0.00992001
R6559 bgr_0.Vbe2.n65 bgr_0.Vbe2.n35 0.00992001
R6560 bgr_0.Vbe2.n34 bgr_0.Vbe2.n33 0.00992001
R6561 bgr_0.Vbe2.n70 bgr_0.Vbe2.n28 0.00992001
R6562 bgr_0.Vbe2.n66 bgr_0.Vbe2.n37 0.00992001
R6563 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 0.00889286
R6564 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 0.00817857
R6565 bgr_0.Vbe2.n73 bgr_0.Vbe2.n71 0.00817857
R6566 bgr_0.Vbe2.n125 bgr_0.Vbe2.n124 0.00817857
R6567 bgr_0.Vbe2.n63 bgr_0.Vbe2.n62 0.00817857
R6568 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t19 1172.87
R6569 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.t28 1172.87
R6570 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t38 996.134
R6571 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t27 996.134
R6572 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.t41 996.134
R6573 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t31 996.134
R6574 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t14 996.134
R6575 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t20 996.134
R6576 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t36 996.134
R6577 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t23 996.134
R6578 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t22 690.867
R6579 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t33 690.867
R6580 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t17 530.201
R6581 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t26 530.201
R6582 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t32 514.134
R6583 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t42 514.134
R6584 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.t29 514.134
R6585 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t39 514.134
R6586 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.t24 514.134
R6587 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t16 514.134
R6588 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.t34 514.134
R6589 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t15 514.134
R6590 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t30 353.467
R6591 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.t13 353.467
R6592 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t18 353.467
R6593 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.t35 353.467
R6594 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t21 353.467
R6595 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t37 353.467
R6596 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t25 353.467
R6597 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t40 353.467
R6598 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R6599 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.n31 176.733
R6600 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 176.733
R6601 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R6602 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R6603 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R6604 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n17 176.733
R6605 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 176.733
R6606 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.n15 176.733
R6607 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 176.733
R6608 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n13 176.733
R6609 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.n12 176.733
R6610 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 176.733
R6611 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.n25 176.733
R6612 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 176.733
R6613 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.n23 176.733
R6614 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 176.733
R6615 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.n21 176.733
R6616 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 166.436
R6617 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n19 161.843
R6618 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 161.718
R6619 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n8 114.689
R6620 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.n1 114.689
R6621 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.n6 114.126
R6622 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.n4 114.126
R6623 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.n2 114.126
R6624 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n0 109.626
R6625 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n38 51.9494
R6626 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.n36 51.9494
R6627 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 51.9494
R6628 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n11 51.9494
R6629 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n27 51.9494
R6630 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.n20 51.9494
R6631 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.X.n40 49.3036
R6632 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n29 18.4693
R6633 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.t10 16.0005
R6634 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.t5 16.0005
R6635 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.t9 16.0005
R6636 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.t11 16.0005
R6637 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.t2 16.0005
R6638 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.t8 16.0005
R6639 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t6 16.0005
R6640 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t3 16.0005
R6641 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t4 16.0005
R6642 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t12 16.0005
R6643 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t7 16.0005
R6644 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t1 16.0005
R6645 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.n10 9.28175
R6646 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 4.5005
R6647 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n30 3.40675
R6648 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.n3 0.563
R6649 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.n5 0.563
R6650 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n7 0.563
R6651 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R6652 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R6653 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R6654 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 206.052
R6655 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 205.488
R6656 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 205.488
R6657 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 205.488
R6658 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 205.488
R6659 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 122.504
R6660 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 71.2813
R6661 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 54.5005
R6662 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R6663 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 39.4005
R6664 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 39.4005
R6665 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 39.4005
R6666 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R6667 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 39.4005
R6668 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R6669 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R6670 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R6671 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R6672 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 19.7005
R6673 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R6674 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R6675 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R6676 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R6677 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R6678 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 19.7005
R6679 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 6.09425
R6680 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 1.15675
R6681 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R6682 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R6683 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R6684 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t1 384.967
R6685 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t5 369.534
R6686 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t20 369.534
R6687 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t23 369.534
R6688 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t15 369.534
R6689 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t17 369.534
R6690 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.n18 369.534
R6691 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 365.491
R6692 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t12 192.8
R6693 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t11 192.8
R6694 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t19 192.8
R6695 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t6 192.8
R6696 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t14 192.8
R6697 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t13 192.8
R6698 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t21 192.8
R6699 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t7 192.8
R6700 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t16 192.8
R6701 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t22 192.8
R6702 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t9 192.8
R6703 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t10 192.8
R6704 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t18 192.8
R6705 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t8 192.8
R6706 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R6707 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R6708 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R6709 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R6710 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R6711 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R6712 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R6713 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R6714 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R6715 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R6716 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R6717 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R6718 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R6719 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R6720 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R6721 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R6722 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R6723 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R6724 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 39.4005
R6725 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t3 39.4005
R6726 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 28.6755
R6727 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t0 24.0005
R6728 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t2 24.0005
R6729 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R6730 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R6731 bgr_0.V_mir2.n4 bgr_0.V_mir2.n3 325.473
R6732 bgr_0.V_mir2.n16 bgr_0.V_mir2.t17 310.488
R6733 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R6734 bgr_0.V_mir2.n0 bgr_0.V_mir2.t20 310.488
R6735 bgr_0.V_mir2.n7 bgr_0.V_mir2.t2 278.312
R6736 bgr_0.V_mir2.n7 bgr_0.V_mir2.n6 228.939
R6737 bgr_0.V_mir2.n8 bgr_0.V_mir2.n5 224.439
R6738 bgr_0.V_mir2.n18 bgr_0.V_mir2.t6 184.097
R6739 bgr_0.V_mir2.n11 bgr_0.V_mir2.t10 184.097
R6740 bgr_0.V_mir2.n2 bgr_0.V_mir2.t8 184.097
R6741 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R6742 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R6743 bgr_0.V_mir2.n1 bgr_0.V_mir2.n0 167.094
R6744 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R6745 bgr_0.V_mir2.n4 bgr_0.V_mir2.n2 152
R6746 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R6747 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 120.501
R6748 bgr_0.V_mir2.n17 bgr_0.V_mir2.t14 120.501
R6749 bgr_0.V_mir2.n9 bgr_0.V_mir2.t19 120.501
R6750 bgr_0.V_mir2.n10 bgr_0.V_mir2.t12 120.501
R6751 bgr_0.V_mir2.n0 bgr_0.V_mir2.t18 120.501
R6752 bgr_0.V_mir2.n1 bgr_0.V_mir2.t4 120.501
R6753 bgr_0.V_mir2.n6 bgr_0.V_mir2.t16 48.0005
R6754 bgr_0.V_mir2.n6 bgr_0.V_mir2.t1 48.0005
R6755 bgr_0.V_mir2.n5 bgr_0.V_mir2.t0 48.0005
R6756 bgr_0.V_mir2.n5 bgr_0.V_mir2.t3 48.0005
R6757 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R6758 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R6759 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 40.7027
R6760 bgr_0.V_mir2.n12 bgr_0.V_mir2.t13 39.4005
R6761 bgr_0.V_mir2.n12 bgr_0.V_mir2.t11 39.4005
R6762 bgr_0.V_mir2.n3 bgr_0.V_mir2.t5 39.4005
R6763 bgr_0.V_mir2.n3 bgr_0.V_mir2.t9 39.4005
R6764 bgr_0.V_mir2.t15 bgr_0.V_mir2.n20 39.4005
R6765 bgr_0.V_mir2.n20 bgr_0.V_mir2.t7 39.4005
R6766 bgr_0.V_mir2.n15 bgr_0.V_mir2.n4 15.8005
R6767 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 15.8005
R6768 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 9.3005
R6769 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 5.8755
R6770 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R6771 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 0.78175
R6772 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6773 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 514.134
R6774 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 323.491
R6775 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 322.692
R6776 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6777 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6778 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 270.591
R6779 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 270.591
R6780 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 233.374
R6781 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 233.374
R6782 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 233.374
R6783 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 233.374
R6784 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 208.838
R6785 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 197.964
R6786 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 174.726
R6787 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 174.726
R6788 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 174.726
R6789 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6790 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 169.216
R6791 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 169.216
R6792 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 169.216
R6793 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 129.24
R6794 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 129.24
R6795 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6796 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6797 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 128.534
R6798 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 128.534
R6799 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 16.8443
R6800 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6801 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6802 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6803 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6804 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6805 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6806 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 4.3755
R6807 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 4.3755
R6808 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 3.688
R6809 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 3.1255
R6810 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 2.0005
R6811 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 1.2755
R6812 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 1.2755
R6813 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 0.8005
R6814 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 632.186
R6815 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 630.264
R6816 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6817 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6818 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 628.003
R6819 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 628.003
R6820 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 626.753
R6821 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 626.753
R6822 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 625.756
R6823 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 622.231
R6824 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6825 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6826 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6827 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6828 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6829 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6830 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6831 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6832 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6833 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6834 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6835 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6836 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6837 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6838 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6839 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6840 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6841 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6842 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6843 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6844 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 8.22272
R6845 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 6.188
R6846 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 630.264
R6847 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n2 627.316
R6848 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 626.784
R6849 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n3 626.784
R6850 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 626.784
R6851 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.n24 585
R6852 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6853 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6854 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.n21 176.733
R6855 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R6856 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6857 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6858 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6859 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6860 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6861 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6862 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6863 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6864 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6865 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6866 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6867 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6868 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6869 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6870 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n23 162.494
R6871 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 135.81
R6872 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n1 131.392
R6873 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6874 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6875 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6876 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6877 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6878 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6879 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6880 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6881 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6882 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6883 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6884 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6885 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6886 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6887 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6888 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6889 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6890 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6891 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6892 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6893 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R6894 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6895 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6896 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6897 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6898 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6899 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6900 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6901 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R6902 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t7 78.8005
R6903 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 49.8072
R6904 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n20 49.8072
R6905 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n25 41.7838
R6906 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6907 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t9 24.0005
R6908 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t8 24.0005
R6909 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 2.313
R6910 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t19 673.034
R6911 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 619.134
R6912 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t28 611.739
R6913 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t16 611.739
R6914 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R6915 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t31 611.739
R6916 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R6917 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R6918 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R6919 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t18 421.75
R6920 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R6921 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t12 421.75
R6922 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R6923 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t24 421.75
R6924 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t27 421.75
R6925 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R6926 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R6927 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R6928 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R6929 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R6930 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R6931 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R6932 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t2 288.166
R6933 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n10 169.311
R6934 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 168.936
R6935 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R6936 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R6937 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R6938 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R6939 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R6940 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R6941 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R6942 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R6943 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R6944 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R6945 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.n3 167.094
R6946 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R6947 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n23 140.547
R6948 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n26 140.546
R6949 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 139.297
R6950 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.n24 139.297
R6951 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n22 109.312
R6952 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t10 62.5402
R6953 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t3 62.5402
R6954 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n18 47.1294
R6955 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n14 47.1294
R6956 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 47.1294
R6957 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n5 47.1294
R6958 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t8 24.0005
R6959 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R6960 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R6961 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R6962 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t1 24.0005
R6963 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R6964 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R6965 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t0 24.0005
R6966 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n1 18.0505
R6967 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 13.0943
R6968 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 5.6255
R6969 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 4.34425
R6970 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n25 3.71925
R6971 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 3.71925
R6972 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n0 160.428
R6973 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n9 160.427
R6974 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 159.803
R6975 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 159.803
R6976 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n3 159.803
R6977 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.n1 159.803
R6978 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n10 159.802
R6979 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n12 159.802
R6980 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n14 159.802
R6981 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n16 159.802
R6982 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 159.802
R6983 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.t0 11.2576
R6984 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R6985 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t16 11.2576
R6986 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R6987 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R6988 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R6989 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t2 11.2576
R6990 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t14 11.2576
R6991 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t19 11.2576
R6992 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R6993 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R6994 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.t8 11.2576
R6995 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t10 11.2576
R6996 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.t12 11.2576
R6997 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R6998 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R6999 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R7000 two_stage_opamp_dummy_magic_0.VD3.n1 two_stage_opamp_dummy_magic_0.VD3.t4 11.2576
R7001 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t6 11.2576
R7002 two_stage_opamp_dummy_magic_0.VD3.n0 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R7003 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t18 11.2576
R7004 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R7005 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n19 8.3755
R7006 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.VD3.n8 6.063
R7007 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.n2 0.6255
R7008 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n4 0.6255
R7009 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n17 0.6255
R7010 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 0.6255
R7011 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n13 0.6255
R7012 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.n11 0.6255
R7013 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n6 0.5005
R7014 a_8420_8490.n8 a_8420_8490.n7 160.427
R7015 a_8420_8490.n2 a_8420_8490.n0 160.427
R7016 a_8420_8490.n6 a_8420_8490.n5 159.802
R7017 a_8420_8490.n4 a_8420_8490.n3 159.802
R7018 a_8420_8490.n2 a_8420_8490.n1 159.802
R7019 a_8420_8490.n9 a_8420_8490.n8 159.798
R7020 a_8420_8490.n7 a_8420_8490.t2 11.2576
R7021 a_8420_8490.n7 a_8420_8490.t0 11.2576
R7022 a_8420_8490.n5 a_8420_8490.t4 11.2576
R7023 a_8420_8490.n5 a_8420_8490.t6 11.2576
R7024 a_8420_8490.n3 a_8420_8490.t1 11.2576
R7025 a_8420_8490.n3 a_8420_8490.t3 11.2576
R7026 a_8420_8490.n1 a_8420_8490.t7 11.2576
R7027 a_8420_8490.n1 a_8420_8490.t9 11.2576
R7028 a_8420_8490.n0 a_8420_8490.t11 11.2576
R7029 a_8420_8490.n0 a_8420_8490.t5 11.2576
R7030 a_8420_8490.n9 a_8420_8490.t8 11.2576
R7031 a_8420_8490.t10 a_8420_8490.n9 11.2576
R7032 a_8420_8490.n4 a_8420_8490.n2 0.6255
R7033 a_8420_8490.n6 a_8420_8490.n4 0.6255
R7034 a_8420_8490.n8 a_8420_8490.n6 0.6255
R7035 w_8160_8260.n6 w_8160_8260.n0 4020
R7036 w_8160_8260.n12 w_8160_8260.n0 4020
R7037 w_8160_8260.n6 w_8160_8260.n1 4020
R7038 w_8160_8260.n12 w_8160_8260.n1 4020
R7039 w_8160_8260.n4 w_8160_8260.t3 660.109
R7040 w_8160_8260.n3 w_8160_8260.t0 660.109
R7041 w_8160_8260.n7 w_8160_8260.n2 428.8
R7042 w_8160_8260.n11 w_8160_8260.n2 428.8
R7043 w_8160_8260.n6 w_8160_8260.t4 239.915
R7044 w_8160_8260.n9 w_8160_8260.n8 230.4
R7045 w_8160_8260.n10 w_8160_8260.n9 230.4
R7046 w_8160_8260.n8 w_8160_8260.n7 198.4
R7047 w_8160_8260.n11 w_8160_8260.n10 198.4
R7048 w_8160_8260.n4 w_8160_8260.t5 155.125
R7049 w_8160_8260.n3 w_8160_8260.t2 155.125
R7050 w_8160_8260.n13 w_8160_8260.t1 147.415
R7051 w_8160_8260.t4 w_8160_8260.t10 98.2764
R7052 w_8160_8260.t10 w_8160_8260.t12 98.2764
R7053 w_8160_8260.t12 w_8160_8260.t14 98.2764
R7054 w_8160_8260.t14 w_8160_8260.t6 98.2764
R7055 w_8160_8260.t6 w_8160_8260.t8 98.2764
R7056 w_8160_8260.t9 w_8160_8260.t11 98.2764
R7057 w_8160_8260.t11 w_8160_8260.t13 98.2764
R7058 w_8160_8260.t13 w_8160_8260.t15 98.2764
R7059 w_8160_8260.t15 w_8160_8260.t7 98.2764
R7060 w_8160_8260.t7 w_8160_8260.t1 98.2764
R7061 w_8160_8260.n12 w_8160_8260.n11 92.5005
R7062 w_8160_8260.n13 w_8160_8260.n12 92.5005
R7063 w_8160_8260.n9 w_8160_8260.n1 92.5005
R7064 w_8160_8260.n5 w_8160_8260.n1 92.5005
R7065 w_8160_8260.n7 w_8160_8260.n6 92.5005
R7066 w_8160_8260.n2 w_8160_8260.n0 92.5005
R7067 w_8160_8260.n5 w_8160_8260.n0 92.5005
R7068 w_8160_8260.t8 w_8160_8260.n5 49.1384
R7069 w_8160_8260.n5 w_8160_8260.t9 49.1384
R7070 w_8160_8260.n14 w_8160_8260.n13 49.1384
R7071 w_8160_8260.n8 w_8160_8260.n4 21.3338
R7072 w_8160_8260.n10 w_8160_8260.n3 21.3338
R7073 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t17 1172.87
R7074 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t22 1172.87
R7075 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t39 996.134
R7076 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.t27 996.134
R7077 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t14 996.134
R7078 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R7079 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t13 996.134
R7080 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.t31 996.134
R7081 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t37 996.134
R7082 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t24 996.134
R7083 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t20 690.867
R7084 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.t25 690.867
R7085 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t16 530.201
R7086 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.t21 530.201
R7087 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t34 514.134
R7088 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t18 514.134
R7089 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t35 514.134
R7090 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t19 514.134
R7091 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t33 514.134
R7092 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t15 514.134
R7093 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t28 514.134
R7094 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.t40 514.134
R7095 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t29 353.467
R7096 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.t36 353.467
R7097 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t23 353.467
R7098 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t38 353.467
R7099 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t26 353.467
R7100 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t42 353.467
R7101 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t30 353.467
R7102 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t41 353.467
R7103 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.n17 176.733
R7104 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 176.733
R7105 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.n15 176.733
R7106 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 176.733
R7107 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.n13 176.733
R7108 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.n11 176.733
R7109 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.n21 176.733
R7110 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.n22 176.733
R7111 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R7112 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R7113 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R7114 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R7115 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.n30 176.733
R7116 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.n31 176.733
R7117 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R7118 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R7119 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R7120 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R7121 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.n19 166.436
R7122 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n29 161.843
R7123 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 161.718
R7124 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n2 114.689
R7125 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n1 114.689
R7126 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n7 114.126
R7127 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n5 114.126
R7128 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.n3 114.126
R7129 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n0 109.626
R7130 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 51.9494
R7131 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n12 51.9494
R7132 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n28 51.9494
R7133 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n27 51.9494
R7134 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 51.9494
R7135 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n36 51.9494
R7136 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t0 49.3037
R7137 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 18.3443
R7138 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R7139 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.t4 16.0005
R7140 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t7 16.0005
R7141 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.t3 16.0005
R7142 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R7143 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R7144 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R7145 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R7146 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t2 16.0005
R7147 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t12 16.0005
R7148 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t10 16.0005
R7149 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t8 16.0005
R7150 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 7.6255
R7151 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 4.5005
R7152 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n20 3.28175
R7153 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n10 1.71925
R7154 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.n4 0.563
R7155 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.n6 0.563
R7156 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n8 0.563
R7157 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.Y.n41 0.063
R7158 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n0 145.989
R7159 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n7 145.989
R7160 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.n5 145.427
R7161 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n3 145.427
R7162 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n1 145.427
R7163 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n9 140.927
R7164 two_stage_opamp_dummy_magic_0.VOUT+.t3 two_stage_opamp_dummy_magic_0.VOUT+.n96 113.192
R7165 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.n91 95.7303
R7166 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.n94 94.6053
R7167 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.n92 94.6053
R7168 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n10 20.688
R7169 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n89 11.7059
R7170 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.n90 10.438
R7171 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t13 6.56717
R7172 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t7 6.56717
R7173 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t11 6.56717
R7174 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t17 6.56717
R7175 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t12 6.56717
R7176 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t6 6.56717
R7177 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t4 6.56717
R7178 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t8 6.56717
R7179 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t5 6.56717
R7180 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t9 6.56717
R7181 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t16 6.56717
R7182 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t10 6.56717
R7183 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t108 4.8295
R7184 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t65 4.8295
R7185 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t118 4.8295
R7186 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t151 4.8295
R7187 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t44 4.8295
R7188 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t67 4.8295
R7189 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t27 4.8295
R7190 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t76 4.8295
R7191 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t62 4.8295
R7192 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t112 4.8295
R7193 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t114 4.8295
R7194 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t99 4.8295
R7195 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t74 4.8295
R7196 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t55 4.8295
R7197 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t109 4.8295
R7198 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t91 4.8295
R7199 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t68 4.8295
R7200 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t52 4.8295
R7201 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t29 4.8295
R7202 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t153 4.8295
R7203 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t63 4.8295
R7204 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t46 4.8295
R7205 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t22 4.8295
R7206 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t146 4.8295
R7207 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t117 4.8295
R7208 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.t72 4.8295
R7209 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t37 4.8295
R7210 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t20 4.8295
R7211 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t79 4.8295
R7212 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t60 4.8295
R7213 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t121 4.8295
R7214 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t104 4.8295
R7215 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t84 4.8295
R7216 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t66 4.8295
R7217 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t123 4.8295
R7218 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t95 4.8154
R7219 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t70 4.8154
R7220 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t110 4.8154
R7221 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t145 4.8154
R7222 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t32 4.806
R7223 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t150 4.806
R7224 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t50 4.806
R7225 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t87 4.806
R7226 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t125 4.806
R7227 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t105 4.806
R7228 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t140 4.806
R7229 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t36 4.806
R7230 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t156 4.806
R7231 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t53 4.806
R7232 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t73 4.806
R7233 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.t116 4.806
R7234 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t64 4.806
R7235 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t154 4.806
R7236 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t106 4.806
R7237 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t143 4.806
R7238 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t96 4.806
R7239 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t42 4.806
R7240 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t86 4.806
R7241 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t34 4.806
R7242 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t69 4.5005
R7243 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.t90 4.5005
R7244 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t80 4.5005
R7245 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.t43 4.5005
R7246 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t56 4.5005
R7247 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.t21 4.5005
R7248 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t98 4.5005
R7249 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.t59 4.5005
R7250 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t136 4.5005
R7251 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.t101 4.5005
R7252 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t30 4.5005
R7253 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.t51 4.5005
R7254 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t155 4.5005
R7255 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t119 4.5005
R7256 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t139 4.5005
R7257 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t102 4.5005
R7258 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t61 4.5005
R7259 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t85 4.5005
R7260 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t45 4.5005
R7261 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t147 4.5005
R7262 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t111 4.5005
R7263 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t134 4.5005
R7264 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t130 4.5005
R7265 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.t152 4.5005
R7266 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t115 4.5005
R7267 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t23 4.5005
R7268 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.t47 4.5005
R7269 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t148 4.5005
R7270 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t78 4.5005
R7271 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.t26 4.5005
R7272 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t132 4.5005
R7273 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t39 4.5005
R7274 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.t128 4.5005
R7275 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t92 4.5005
R7276 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t71 4.5005
R7277 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.t19 4.5005
R7278 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t126 4.5005
R7279 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t33 4.5005
R7280 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.t122 4.5005
R7281 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t88 4.5005
R7282 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t135 4.5005
R7283 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.t82 4.5005
R7284 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t48 4.5005
R7285 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t28 4.5005
R7286 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.t120 4.5005
R7287 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t81 4.5005
R7288 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t129 4.5005
R7289 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.t77 4.5005
R7290 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t40 4.5005
R7291 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t25 4.5005
R7292 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.t124 4.5005
R7293 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.t38 4.5005
R7294 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.t127 4.5005
R7295 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t94 4.5005
R7296 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t54 4.5005
R7297 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t144 4.5005
R7298 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t113 4.5005
R7299 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t75 4.5005
R7300 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t24 4.5005
R7301 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t131 4.5005
R7302 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t97 4.5005
R7303 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.t58 4.5005
R7304 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t149 4.5005
R7305 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t142 4.5005
R7306 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.t93 4.5005
R7307 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t57 4.5005
R7308 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t41 4.5005
R7309 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.t133 4.5005
R7310 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t100 4.5005
R7311 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t83 4.5005
R7312 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.t31 4.5005
R7313 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t137 4.5005
R7314 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t49 4.5005
R7315 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.t138 4.5005
R7316 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t103 4.5005
R7317 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t89 4.5005
R7318 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.t35 4.5005
R7319 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.t141 4.5005
R7320 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.t107 4.5005
R7321 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n8 4.5005
R7322 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.t2 3.42907
R7323 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.t15 3.42907
R7324 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.t0 3.42907
R7325 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.t14 3.42907
R7326 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t18 3.42907
R7327 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t1 3.42907
R7328 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.n95 2.03175
R7329 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.n93 1.1255
R7330 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n2 0.563
R7331 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.n4 0.563
R7332 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n6 0.563
R7333 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.n37 0.3295
R7334 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.n46 0.3295
R7335 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.n44 0.3295
R7336 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.n42 0.3295
R7337 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.n40 0.3295
R7338 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n39 0.3295
R7339 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n57 0.3295
R7340 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.n56 0.3295
R7341 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.n55 0.3295
R7342 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.n54 0.3295
R7343 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.n53 0.3295
R7344 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.n52 0.3295
R7345 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.n51 0.3295
R7346 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.n50 0.3295
R7347 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.n49 0.3295
R7348 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.n48 0.3295
R7349 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n59 0.3295
R7350 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n60 0.3295
R7351 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n62 0.3295
R7352 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n63 0.3295
R7353 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.n65 0.3295
R7354 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.n66 0.3295
R7355 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.n68 0.3295
R7356 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.n69 0.3295
R7357 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.n71 0.3295
R7358 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.n72 0.3295
R7359 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.n74 0.3295
R7360 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.n75 0.3295
R7361 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.n77 0.3295
R7362 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.n78 0.3295
R7363 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.n80 0.3295
R7364 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.n81 0.3295
R7365 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.n83 0.3295
R7366 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.n84 0.3295
R7367 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.n11 0.3295
R7368 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n13 0.3295
R7369 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n23 0.3295
R7370 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.n22 0.3295
R7371 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.n21 0.3295
R7372 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.n20 0.3295
R7373 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.n19 0.3295
R7374 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.n18 0.3295
R7375 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.n17 0.3295
R7376 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.n16 0.3295
R7377 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.n15 0.3295
R7378 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.n14 0.3295
R7379 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n25 0.3295
R7380 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n26 0.3295
R7381 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n28 0.3295
R7382 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n29 0.3295
R7383 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n31 0.3295
R7384 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n32 0.3295
R7385 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n34 0.3295
R7386 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n35 0.3295
R7387 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n86 0.3295
R7388 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.n87 0.3295
R7389 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.n88 0.3295
R7390 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.n47 0.306
R7391 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.n45 0.306
R7392 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.n43 0.306
R7393 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.n41 0.306
R7394 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n38 0.2825
R7395 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n58 0.2825
R7396 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.n61 0.2825
R7397 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.n64 0.2825
R7398 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.n67 0.2825
R7399 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.n70 0.2825
R7400 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.n73 0.2825
R7401 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.n76 0.2825
R7402 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.n79 0.2825
R7403 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.n82 0.2825
R7404 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n12 0.2825
R7405 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n24 0.2825
R7406 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.n27 0.2825
R7407 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.n30 0.2825
R7408 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.n33 0.2825
R7409 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n36 0.2825
R7410 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n85 0.2825
R7411 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t10 449.868
R7412 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7413 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R7414 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R7415 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7416 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7417 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7418 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7419 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7420 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7421 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t14 273.134
R7422 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7423 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t2 184.625
R7424 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n11 182.972
R7425 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R7426 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R7427 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R7428 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R7429 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R7430 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7431 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n13 99.2817
R7432 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t1 61.1914
R7433 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 56.2338
R7434 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n6 56.2338
R7435 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t3 39.4005
R7436 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t4 39.4005
R7437 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7438 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7439 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 14.3735
R7440 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 4.46925
R7441 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t25 369.534
R7442 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t24 369.534
R7443 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t15 369.534
R7444 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t11 369.534
R7445 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t17 369.534
R7446 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t16 369.534
R7447 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7448 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7449 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7450 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7451 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t21 238.322
R7452 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t13 238.322
R7453 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t2 194.895
R7454 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t18 192.8
R7455 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t10 192.8
R7456 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t14 192.8
R7457 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t22 192.8
R7458 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t28 192.8
R7459 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t19 192.8
R7460 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t26 192.8
R7461 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t12 192.8
R7462 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t20 192.8
R7463 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t27 192.8
R7464 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t29 192.8
R7465 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t23 192.8
R7466 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7467 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7468 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7469 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7470 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7471 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7472 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7473 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 169.394
R7474 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7475 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7476 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t4 100.635
R7477 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7478 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7479 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7480 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7481 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7482 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7483 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t5 39.4005
R7484 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t3 39.4005
R7485 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t7 39.4005
R7486 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t8 39.4005
R7487 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t1 39.4005
R7488 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t9 39.4005
R7489 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t0 39.4005
R7490 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t6 39.4005
R7491 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 26.9067
R7492 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 5.15675
R7493 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7494 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n14 4.188
R7495 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 3.03175
R7496 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7497 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7498 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R7499 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 344.7
R7500 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R7501 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 206.052
R7502 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 205.488
R7503 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 205.488
R7504 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 205.488
R7505 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 205.488
R7506 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 122.474
R7507 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 83.3443
R7508 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 39.4005
R7509 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 39.4005
R7510 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 39.4005
R7511 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R7512 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 39.4005
R7513 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R7514 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R7515 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R7516 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R7517 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 19.7005
R7518 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R7519 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 19.7005
R7520 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R7521 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 19.7005
R7522 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R7523 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R7524 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 6.15675
R7525 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 6.1255
R7526 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R7527 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R7528 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R7529 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R7530 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 0.21925
R7531 a_14520_5068.t0 a_14520_5068.t1 294.339
R7532 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 144.827
R7533 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 134.577
R7534 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 120.629
R7535 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 114.501
R7536 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 97.4009
R7537 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 96.8384
R7538 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 96.8384
R7539 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 96.8384
R7540 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 96.8384
R7541 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R7542 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 24.0005
R7543 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R7544 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 24.0005
R7545 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R7546 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 8.0005
R7547 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R7548 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 8.0005
R7549 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R7550 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R7551 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 8.0005
R7552 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R7553 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R7554 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R7555 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 5.84425
R7556 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 1.46925
R7557 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 0.563
R7558 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 0.563
R7559 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 0.563
R7560 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7561 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7562 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7563 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 310.488
R7564 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7565 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7566 bgr_0.V_mir1.n7 bgr_0.V_mir1.t14 278.312
R7567 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7568 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7569 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R7570 bgr_0.V_mir1.n11 bgr_0.V_mir1.t0 184.097
R7571 bgr_0.V_mir1.n2 bgr_0.V_mir1.t8 184.097
R7572 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7573 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7574 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7575 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7576 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7577 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7578 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 120.501
R7579 bgr_0.V_mir1.n17 bgr_0.V_mir1.t2 120.501
R7580 bgr_0.V_mir1.n9 bgr_0.V_mir1.t18 120.501
R7581 bgr_0.V_mir1.n10 bgr_0.V_mir1.t4 120.501
R7582 bgr_0.V_mir1.n0 bgr_0.V_mir1.t17 120.501
R7583 bgr_0.V_mir1.n1 bgr_0.V_mir1.t6 120.501
R7584 bgr_0.V_mir1.n6 bgr_0.V_mir1.t13 48.0005
R7585 bgr_0.V_mir1.n6 bgr_0.V_mir1.t16 48.0005
R7586 bgr_0.V_mir1.n5 bgr_0.V_mir1.t12 48.0005
R7587 bgr_0.V_mir1.n5 bgr_0.V_mir1.t15 48.0005
R7588 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7589 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7590 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7591 bgr_0.V_mir1.n12 bgr_0.V_mir1.t1 39.4005
R7592 bgr_0.V_mir1.n12 bgr_0.V_mir1.t5 39.4005
R7593 bgr_0.V_mir1.n3 bgr_0.V_mir1.t9 39.4005
R7594 bgr_0.V_mir1.n3 bgr_0.V_mir1.t7 39.4005
R7595 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7596 bgr_0.V_mir1.n20 bgr_0.V_mir1.t3 39.4005
R7597 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7598 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7599 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7600 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7601 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7602 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7603 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 50.0055
R7604 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1603
R7605 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R7606 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.1603
R7607 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.1603
R7608 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.1603
R7609 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1603
R7610 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1603
R7611 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1603
R7612 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.1603
R7613 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R7614 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1603
R7615 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R7616 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.1603
R7617 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.1603
R7618 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.1603
R7619 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R7620 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1603
R7621 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1603
R7622 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.1603
R7623 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R7624 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1603
R7625 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1603
R7626 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.1603
R7627 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.1603
R7628 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.1603
R7629 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R7630 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.1603
R7631 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.1603
R7632 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.1603
R7633 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.1603
R7634 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R7635 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1603
R7636 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R7637 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1603
R7638 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1603
R7639 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1603
R7640 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.1603
R7641 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1603
R7642 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R7643 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R7644 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R7645 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1603
R7646 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R7647 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1603
R7648 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.1603
R7649 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R7650 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.1603
R7651 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R7652 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1603
R7653 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1603
R7654 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1603
R7655 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.1603
R7656 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R7657 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1603
R7658 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.1603
R7659 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.1603
R7660 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1603
R7661 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.1603
R7662 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.159278
R7663 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.159278
R7664 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.159278
R7665 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.159278
R7666 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.159278
R7667 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.159278
R7668 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.159278
R7669 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.159278
R7670 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.159278
R7671 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.159278
R7672 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.159278
R7673 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.159278
R7674 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.159278
R7675 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R7676 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R7677 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R7678 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R7679 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R7680 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R7681 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R7682 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R7683 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R7684 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R7685 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.159278
R7686 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.159278
R7687 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.159278
R7688 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.159278
R7689 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.137822
R7690 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1368
R7691 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.1368
R7692 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1368
R7693 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1368
R7694 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1368
R7695 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.1368
R7696 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.1368
R7697 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1368
R7698 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R7699 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1368
R7700 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1368
R7701 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.1368
R7702 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1368
R7703 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1368
R7704 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.1368
R7705 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1368
R7706 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1368
R7707 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1368
R7708 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.1368
R7709 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.1368
R7710 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1368
R7711 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.1368
R7712 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1368
R7713 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.1368
R7714 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.1368
R7715 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1368
R7716 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1368
R7717 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.1368
R7718 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1368
R7719 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1368
R7720 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.1368
R7721 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.114322
R7722 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.1133
R7723 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.1133
R7724 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R7725 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R7726 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R7727 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R7728 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R7729 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R7730 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R7731 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R7732 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R7733 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R7734 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R7735 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R7736 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.1133
R7737 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.1133
R7738 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.1133
R7739 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.1133
R7740 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R7741 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.00152174
R7742 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R7743 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.00152174
R7744 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.00152174
R7745 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.00152174
R7746 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.00152174
R7747 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.00152174
R7748 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R7749 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.00152174
R7750 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.00152174
R7751 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.00152174
R7752 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.00152174
R7753 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.00152174
R7754 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.00152174
R7755 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.00152174
R7756 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.00152174
R7757 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.00152174
R7758 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.00152174
R7759 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.00152174
R7760 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.00152174
R7761 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.00152174
R7762 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.00152174
R7763 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.00152174
R7764 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.00152174
R7765 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.00152174
R7766 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.00152174
R7767 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.00152174
R7768 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R7769 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.00152174
R7770 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.00152174
R7771 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.00152174
R7772 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R7773 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.00152174
R7774 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R7775 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R7776 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R7777 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R7778 bgr_0.TAIL_CUR_MIR_BIAS.n17 bgr_0.TAIL_CUR_MIR_BIAS.t12 610.534
R7779 bgr_0.TAIL_CUR_MIR_BIAS.n8 bgr_0.TAIL_CUR_MIR_BIAS.t14 610.534
R7780 bgr_0.TAIL_CUR_MIR_BIAS.n17 bgr_0.TAIL_CUR_MIR_BIAS.t30 433.8
R7781 bgr_0.TAIL_CUR_MIR_BIAS.n18 bgr_0.TAIL_CUR_MIR_BIAS.t21 433.8
R7782 bgr_0.TAIL_CUR_MIR_BIAS.n19 bgr_0.TAIL_CUR_MIR_BIAS.t27 433.8
R7783 bgr_0.TAIL_CUR_MIR_BIAS.n20 bgr_0.TAIL_CUR_MIR_BIAS.t17 433.8
R7784 bgr_0.TAIL_CUR_MIR_BIAS.n21 bgr_0.TAIL_CUR_MIR_BIAS.t25 433.8
R7785 bgr_0.TAIL_CUR_MIR_BIAS.n22 bgr_0.TAIL_CUR_MIR_BIAS.t15 433.8
R7786 bgr_0.TAIL_CUR_MIR_BIAS.n23 bgr_0.TAIL_CUR_MIR_BIAS.t23 433.8
R7787 bgr_0.TAIL_CUR_MIR_BIAS.n24 bgr_0.TAIL_CUR_MIR_BIAS.t29 433.8
R7788 bgr_0.TAIL_CUR_MIR_BIAS.n25 bgr_0.TAIL_CUR_MIR_BIAS.t19 433.8
R7789 bgr_0.TAIL_CUR_MIR_BIAS.n16 bgr_0.TAIL_CUR_MIR_BIAS.t31 433.8
R7790 bgr_0.TAIL_CUR_MIR_BIAS.n15 bgr_0.TAIL_CUR_MIR_BIAS.t22 433.8
R7791 bgr_0.TAIL_CUR_MIR_BIAS.n14 bgr_0.TAIL_CUR_MIR_BIAS.t28 433.8
R7792 bgr_0.TAIL_CUR_MIR_BIAS.n13 bgr_0.TAIL_CUR_MIR_BIAS.t18 433.8
R7793 bgr_0.TAIL_CUR_MIR_BIAS.n12 bgr_0.TAIL_CUR_MIR_BIAS.t26 433.8
R7794 bgr_0.TAIL_CUR_MIR_BIAS.n11 bgr_0.TAIL_CUR_MIR_BIAS.t16 433.8
R7795 bgr_0.TAIL_CUR_MIR_BIAS.n10 bgr_0.TAIL_CUR_MIR_BIAS.t24 433.8
R7796 bgr_0.TAIL_CUR_MIR_BIAS.n9 bgr_0.TAIL_CUR_MIR_BIAS.t13 433.8
R7797 bgr_0.TAIL_CUR_MIR_BIAS.n8 bgr_0.TAIL_CUR_MIR_BIAS.t20 433.8
R7798 bgr_0.TAIL_CUR_MIR_BIAS.n3 bgr_0.TAIL_CUR_MIR_BIAS.n1 339.836
R7799 bgr_0.TAIL_CUR_MIR_BIAS.n5 bgr_0.TAIL_CUR_MIR_BIAS.n4 339.834
R7800 bgr_0.TAIL_CUR_MIR_BIAS.n3 bgr_0.TAIL_CUR_MIR_BIAS.n2 339.272
R7801 bgr_0.TAIL_CUR_MIR_BIAS.n6 bgr_0.TAIL_CUR_MIR_BIAS.n0 334.772
R7802 bgr_0.TAIL_CUR_MIR_BIAS.n28 bgr_0.TAIL_CUR_MIR_BIAS.n26 221.293
R7803 bgr_0.TAIL_CUR_MIR_BIAS.n25 bgr_0.TAIL_CUR_MIR_BIAS.n24 176.733
R7804 bgr_0.TAIL_CUR_MIR_BIAS.n24 bgr_0.TAIL_CUR_MIR_BIAS.n23 176.733
R7805 bgr_0.TAIL_CUR_MIR_BIAS.n23 bgr_0.TAIL_CUR_MIR_BIAS.n22 176.733
R7806 bgr_0.TAIL_CUR_MIR_BIAS.n22 bgr_0.TAIL_CUR_MIR_BIAS.n21 176.733
R7807 bgr_0.TAIL_CUR_MIR_BIAS.n21 bgr_0.TAIL_CUR_MIR_BIAS.n20 176.733
R7808 bgr_0.TAIL_CUR_MIR_BIAS.n20 bgr_0.TAIL_CUR_MIR_BIAS.n19 176.733
R7809 bgr_0.TAIL_CUR_MIR_BIAS.n19 bgr_0.TAIL_CUR_MIR_BIAS.n18 176.733
R7810 bgr_0.TAIL_CUR_MIR_BIAS.n18 bgr_0.TAIL_CUR_MIR_BIAS.n17 176.733
R7811 bgr_0.TAIL_CUR_MIR_BIAS.n9 bgr_0.TAIL_CUR_MIR_BIAS.n8 176.733
R7812 bgr_0.TAIL_CUR_MIR_BIAS.n10 bgr_0.TAIL_CUR_MIR_BIAS.n9 176.733
R7813 bgr_0.TAIL_CUR_MIR_BIAS.n11 bgr_0.TAIL_CUR_MIR_BIAS.n10 176.733
R7814 bgr_0.TAIL_CUR_MIR_BIAS.n12 bgr_0.TAIL_CUR_MIR_BIAS.n11 176.733
R7815 bgr_0.TAIL_CUR_MIR_BIAS.n13 bgr_0.TAIL_CUR_MIR_BIAS.n12 176.733
R7816 bgr_0.TAIL_CUR_MIR_BIAS.n14 bgr_0.TAIL_CUR_MIR_BIAS.n13 176.733
R7817 bgr_0.TAIL_CUR_MIR_BIAS.n15 bgr_0.TAIL_CUR_MIR_BIAS.n14 176.733
R7818 bgr_0.TAIL_CUR_MIR_BIAS.n16 bgr_0.TAIL_CUR_MIR_BIAS.n15 176.733
R7819 bgr_0.TAIL_CUR_MIR_BIAS.n29 bgr_0.TAIL_CUR_MIR_BIAS.n7 118.45
R7820 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.TAIL_CUR_MIR_BIAS.n29 86.7036
R7821 bgr_0.TAIL_CUR_MIR_BIAS.n29 bgr_0.TAIL_CUR_MIR_BIAS.n28 64.5795
R7822 bgr_0.TAIL_CUR_MIR_BIAS.n26 bgr_0.TAIL_CUR_MIR_BIAS.n25 56.2338
R7823 bgr_0.TAIL_CUR_MIR_BIAS.n26 bgr_0.TAIL_CUR_MIR_BIAS.n16 56.2338
R7824 bgr_0.TAIL_CUR_MIR_BIAS.n28 bgr_0.TAIL_CUR_MIR_BIAS.n27 53.2453
R7825 bgr_0.TAIL_CUR_MIR_BIAS.n0 bgr_0.TAIL_CUR_MIR_BIAS.t5 39.4005
R7826 bgr_0.TAIL_CUR_MIR_BIAS.n0 bgr_0.TAIL_CUR_MIR_BIAS.t10 39.4005
R7827 bgr_0.TAIL_CUR_MIR_BIAS.n4 bgr_0.TAIL_CUR_MIR_BIAS.t7 39.4005
R7828 bgr_0.TAIL_CUR_MIR_BIAS.n4 bgr_0.TAIL_CUR_MIR_BIAS.t4 39.4005
R7829 bgr_0.TAIL_CUR_MIR_BIAS.n1 bgr_0.TAIL_CUR_MIR_BIAS.t9 39.4005
R7830 bgr_0.TAIL_CUR_MIR_BIAS.n1 bgr_0.TAIL_CUR_MIR_BIAS.t6 39.4005
R7831 bgr_0.TAIL_CUR_MIR_BIAS.n2 bgr_0.TAIL_CUR_MIR_BIAS.t11 39.4005
R7832 bgr_0.TAIL_CUR_MIR_BIAS.n2 bgr_0.TAIL_CUR_MIR_BIAS.t8 39.4005
R7833 bgr_0.TAIL_CUR_MIR_BIAS bgr_0.TAIL_CUR_MIR_BIAS.n6 18.3599
R7834 bgr_0.TAIL_CUR_MIR_BIAS.n27 bgr_0.TAIL_CUR_MIR_BIAS.t3 16.0005
R7835 bgr_0.TAIL_CUR_MIR_BIAS.n27 bgr_0.TAIL_CUR_MIR_BIAS.t1 16.0005
R7836 bgr_0.TAIL_CUR_MIR_BIAS.n7 bgr_0.TAIL_CUR_MIR_BIAS.t0 16.0005
R7837 bgr_0.TAIL_CUR_MIR_BIAS.n7 bgr_0.TAIL_CUR_MIR_BIAS.t2 16.0005
R7838 bgr_0.TAIL_CUR_MIR_BIAS.n6 bgr_0.TAIL_CUR_MIR_BIAS.n5 4.5005
R7839 bgr_0.TAIL_CUR_MIR_BIAS.n5 bgr_0.TAIL_CUR_MIR_BIAS.n3 0.563
R7840 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 219.928
R7841 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R7842 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t1 16.0005
R7843 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R7844 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t3 9.6005
R7845 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 229.562
R7846 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7847 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7848 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7849 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7850 bgr_0.V_p_2.n1 bgr_0.V_p_2.t5 98.2279
R7851 bgr_0.V_p_2.n5 bgr_0.V_p_2.t6 48.0005
R7852 bgr_0.V_p_2.n5 bgr_0.V_p_2.t3 48.0005
R7853 bgr_0.V_p_2.n4 bgr_0.V_p_2.t0 48.0005
R7854 bgr_0.V_p_2.n4 bgr_0.V_p_2.t7 48.0005
R7855 bgr_0.V_p_2.n3 bgr_0.V_p_2.t10 48.0005
R7856 bgr_0.V_p_2.n3 bgr_0.V_p_2.t2 48.0005
R7857 bgr_0.V_p_2.n2 bgr_0.V_p_2.t1 48.0005
R7858 bgr_0.V_p_2.n2 bgr_0.V_p_2.t9 48.0005
R7859 bgr_0.V_p_2.t4 bgr_0.V_p_2.n6 48.0005
R7860 bgr_0.V_p_2.n6 bgr_0.V_p_2.t8 48.0005
R7861 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7862 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7863 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7864 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7865 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7866 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7867 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7868 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7869 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7870 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7871 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7872 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7873 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7874 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7875 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7876 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7877 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7878 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7879 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7880 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7881 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7882 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7883 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7884 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t19 78.8005
R7885 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7886 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7887 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7888 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7889 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7890 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7891 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7892 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7893 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7894 two_stage_opamp_dummy_magic_0.V_err_p.t17 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7895 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7896 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7897 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.60845
R7898 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R7899 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R7900 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R7901 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7902 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7903 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R7904 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R7905 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R7906 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R7907 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 167.05
R7908 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R7909 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R7910 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R7911 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R7912 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R7913 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R7914 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R7915 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R7916 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R7917 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 117.591
R7918 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 117.591
R7919 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t1 108.424
R7920 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t2 108.424
R7921 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 35.9871
R7922 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n0 35.9246
R7923 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 10.6255
R7924 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 1.8755
R7925 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n4 1.31612
R7926 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.26612
R7927 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 1.15363
R7928 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 114.719
R7929 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7930 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7931 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n7 114.156
R7932 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7933 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7934 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7935 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7936 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7937 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7938 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7939 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7940 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7941 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7942 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7943 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7944 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7945 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7946 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7947 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7948 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7949 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7950 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7951 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7952 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7953 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7954 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7955 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7956 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7957 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7958 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7959 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7960 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7961 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7962 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7963 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7964 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7965 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7966 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7967 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n8 0.563
R7968 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7969 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7970 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 525.38
R7971 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 525.38
R7972 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 366.856
R7973 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 366.856
R7974 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 281.168
R7975 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 281.168
R7976 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 281.168
R7977 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 281.168
R7978 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7979 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7980 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7981 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7982 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7983 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7984 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7985 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7986 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 17.688
R7987 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R7988 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R7989 bgr_0.Vin+.n0 bgr_0.Vin+.t6 303.259
R7990 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R7991 bgr_0.Vin+.n0 bgr_0.Vin+.t8 174.726
R7992 bgr_0.Vin+.n1 bgr_0.Vin+.t10 174.726
R7993 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R7994 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R7995 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R7996 bgr_0.Vin+.n8 bgr_0.Vin+.t1 158.796
R7997 bgr_0.Vin+.t0 bgr_0.Vin+.n8 147.981
R7998 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R7999 bgr_0.Vin+.n3 bgr_0.Vin+.t9 96.4005
R8000 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R8001 bgr_0.Vin+.n5 bgr_0.Vin+.t2 13.1338
R8002 bgr_0.Vin+.n5 bgr_0.Vin+.t5 13.1338
R8003 bgr_0.Vin+.n4 bgr_0.Vin+.t4 13.1338
R8004 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R8005 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R8006 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 229.562
R8007 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R8008 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R8009 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R8010 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R8011 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.2279
R8012 bgr_0.V_p_1.n5 bgr_0.V_p_1.t5 48.0005
R8013 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R8014 bgr_0.V_p_1.n4 bgr_0.V_p_1.t0 48.0005
R8015 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8016 bgr_0.V_p_1.n3 bgr_0.V_p_1.t6 48.0005
R8017 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R8018 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R8019 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R8020 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8021 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R8022 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R8023 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t13 355.293
R8024 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.t14 346.8
R8025 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.n20 339.522
R8026 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 339.522
R8027 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n14 335.022
R8028 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t8 275.909
R8029 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 227.909
R8030 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 222.034
R8031 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t26 184.097
R8032 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t36 184.097
R8033 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t19 184.097
R8034 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t32 184.097
R8035 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n17 166.05
R8036 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n8 166.05
R8037 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n4 57.7228
R8038 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t7 48.0005
R8039 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t6 48.0005
R8040 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t9 48.0005
R8041 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t10 48.0005
R8042 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t0 39.4005
R8043 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t3 39.4005
R8044 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t2 39.4005
R8045 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t4 39.4005
R8046 bgr_0.1st_Vout_2.t5 bgr_0.1st_Vout_2.n21 39.4005
R8047 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.t1 39.4005
R8048 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t17 4.8295
R8049 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t16 4.8295
R8050 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t27 4.8295
R8051 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t23 4.8295
R8052 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t35 4.8295
R8053 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t34 4.8295
R8054 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t28 4.8295
R8055 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R8056 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t15 4.5005
R8057 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t12 4.5005
R8058 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t30 4.5005
R8059 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t22 4.5005
R8060 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t18 4.5005
R8061 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t11 4.5005
R8062 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R8063 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t29 4.5005
R8064 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.5005
R8065 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t24 4.5005
R8066 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R8067 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.5005
R8068 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n11 4.5005
R8069 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n15 4.5005
R8070 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n7 1.3755
R8071 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n16 1.3755
R8072 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 1.188
R8073 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 0.9405
R8074 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n0 0.8935
R8075 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n13 0.78175
R8076 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 0.6585
R8077 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n3 0.6585
R8078 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n1 0.6585
R8079 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n9 0.6255
R8080 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n18 0.6255
R8081 bgr_0.cap_res2 bgr_0.cap_res2.t20 188.315
R8082 bgr_0.cap_res2 bgr_0.cap_res2.t9 0.259
R8083 bgr_0.cap_res2.t13 bgr_0.cap_res2.t8 0.1603
R8084 bgr_0.cap_res2.t2 bgr_0.cap_res2.t6 0.1603
R8085 bgr_0.cap_res2.t5 bgr_0.cap_res2.t1 0.1603
R8086 bgr_0.cap_res2.t19 bgr_0.cap_res2.t0 0.1603
R8087 bgr_0.cap_res2.t14 bgr_0.cap_res2.t10 0.1603
R8088 bgr_0.cap_res2.t4 bgr_0.cap_res2.t7 0.1603
R8089 bgr_0.cap_res2.t18 bgr_0.cap_res2.t16 0.1603
R8090 bgr_0.cap_res2.t12 bgr_0.cap_res2.t15 0.1603
R8091 bgr_0.cap_res2.n1 bgr_0.cap_res2.t17 0.159278
R8092 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.159278
R8093 bgr_0.cap_res2.n3 bgr_0.cap_res2.t3 0.159278
R8094 bgr_0.cap_res2.n3 bgr_0.cap_res2.t13 0.1368
R8095 bgr_0.cap_res2.n3 bgr_0.cap_res2.t2 0.1368
R8096 bgr_0.cap_res2.n2 bgr_0.cap_res2.t5 0.1368
R8097 bgr_0.cap_res2.n2 bgr_0.cap_res2.t19 0.1368
R8098 bgr_0.cap_res2.n1 bgr_0.cap_res2.t14 0.1368
R8099 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R8100 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R8101 bgr_0.cap_res2.n0 bgr_0.cap_res2.t12 0.1368
R8102 bgr_0.cap_res2.t17 bgr_0.cap_res2.n0 0.00152174
R8103 bgr_0.cap_res2.t11 bgr_0.cap_res2.n1 0.00152174
R8104 bgr_0.cap_res2.t3 bgr_0.cap_res2.n2 0.00152174
R8105 bgr_0.cap_res2.t9 bgr_0.cap_res2.n3 0.00152174
R8106 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.t9 206.407
R8107 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n26 118.168
R8108 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n19 117.831
R8109 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n33 117.269
R8110 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n31 117.269
R8111 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n29 117.269
R8112 two_stage_opamp_dummy_magic_0.V_p.n28 two_stage_opamp_dummy_magic_0.V_p.n27 117.269
R8113 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n24 117.269
R8114 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n22 117.269
R8115 two_stage_opamp_dummy_magic_0.V_p.n21 two_stage_opamp_dummy_magic_0.V_p.n20 117.269
R8116 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n18 113.136
R8117 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n3 99.647
R8118 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n0 99.5532
R8119 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n15 99.0845
R8120 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.n13 99.0845
R8121 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.n11 99.0845
R8122 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n6 99.0845
R8123 two_stage_opamp_dummy_magic_0.V_p.n5 two_stage_opamp_dummy_magic_0.V_p.n4 99.0845
R8124 two_stage_opamp_dummy_magic_0.V_p.n2 two_stage_opamp_dummy_magic_0.V_p.n1 99.0845
R8125 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.n37 94.5857
R8126 two_stage_opamp_dummy_magic_0.V_p.n9 two_stage_opamp_dummy_magic_0.V_p.n8 94.5845
R8127 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.t17 16.0005
R8128 two_stage_opamp_dummy_magic_0.V_p.n33 two_stage_opamp_dummy_magic_0.V_p.t16 16.0005
R8129 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t2 16.0005
R8130 two_stage_opamp_dummy_magic_0.V_p.n31 two_stage_opamp_dummy_magic_0.V_p.t40 16.0005
R8131 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t18 16.0005
R8132 two_stage_opamp_dummy_magic_0.V_p.n29 two_stage_opamp_dummy_magic_0.V_p.t4 16.0005
R8133 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t8 16.0005
R8134 two_stage_opamp_dummy_magic_0.V_p.n27 two_stage_opamp_dummy_magic_0.V_p.t19 16.0005
R8135 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t1 16.0005
R8136 two_stage_opamp_dummy_magic_0.V_p.n26 two_stage_opamp_dummy_magic_0.V_p.t13 16.0005
R8137 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t11 16.0005
R8138 two_stage_opamp_dummy_magic_0.V_p.n24 two_stage_opamp_dummy_magic_0.V_p.t10 16.0005
R8139 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t15 16.0005
R8140 two_stage_opamp_dummy_magic_0.V_p.n22 two_stage_opamp_dummy_magic_0.V_p.t7 16.0005
R8141 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t20 16.0005
R8142 two_stage_opamp_dummy_magic_0.V_p.n20 two_stage_opamp_dummy_magic_0.V_p.t3 16.0005
R8143 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t14 16.0005
R8144 two_stage_opamp_dummy_magic_0.V_p.n19 two_stage_opamp_dummy_magic_0.V_p.t5 16.0005
R8145 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.t0 16.0005
R8146 two_stage_opamp_dummy_magic_0.V_p.n18 two_stage_opamp_dummy_magic_0.V_p.t12 16.0005
R8147 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t36 9.6005
R8148 two_stage_opamp_dummy_magic_0.V_p.n15 two_stage_opamp_dummy_magic_0.V_p.t26 9.6005
R8149 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t34 9.6005
R8150 two_stage_opamp_dummy_magic_0.V_p.n13 two_stage_opamp_dummy_magic_0.V_p.t24 9.6005
R8151 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.t30 9.6005
R8152 two_stage_opamp_dummy_magic_0.V_p.n11 two_stage_opamp_dummy_magic_0.V_p.t22 9.6005
R8153 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t33 9.6005
R8154 two_stage_opamp_dummy_magic_0.V_p.n8 two_stage_opamp_dummy_magic_0.V_p.t23 9.6005
R8155 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t29 9.6005
R8156 two_stage_opamp_dummy_magic_0.V_p.n6 two_stage_opamp_dummy_magic_0.V_p.t37 9.6005
R8157 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t27 9.6005
R8158 two_stage_opamp_dummy_magic_0.V_p.n4 two_stage_opamp_dummy_magic_0.V_p.t35 9.6005
R8159 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t25 9.6005
R8160 two_stage_opamp_dummy_magic_0.V_p.n3 two_stage_opamp_dummy_magic_0.V_p.t31 9.6005
R8161 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t38 9.6005
R8162 two_stage_opamp_dummy_magic_0.V_p.n1 two_stage_opamp_dummy_magic_0.V_p.t32 9.6005
R8163 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t21 9.6005
R8164 two_stage_opamp_dummy_magic_0.V_p.n0 two_stage_opamp_dummy_magic_0.V_p.t6 9.6005
R8165 two_stage_opamp_dummy_magic_0.V_p.t39 two_stage_opamp_dummy_magic_0.V_p.n38 9.6005
R8166 two_stage_opamp_dummy_magic_0.V_p.n38 two_stage_opamp_dummy_magic_0.V_p.t28 9.6005
R8167 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.n9 4.5005
R8168 two_stage_opamp_dummy_magic_0.V_p.n36 two_stage_opamp_dummy_magic_0.V_p.n35 4.5005
R8169 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n17 4.5005
R8170 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.n34 3.65675
R8171 two_stage_opamp_dummy_magic_0.V_p.n37 two_stage_opamp_dummy_magic_0.V_p.n36 1.28175
R8172 two_stage_opamp_dummy_magic_0.V_p.n7 two_stage_opamp_dummy_magic_0.V_p.n5 0.563
R8173 two_stage_opamp_dummy_magic_0.V_p.n10 two_stage_opamp_dummy_magic_0.V_p.n7 0.563
R8174 two_stage_opamp_dummy_magic_0.V_p.n12 two_stage_opamp_dummy_magic_0.V_p.n10 0.563
R8175 two_stage_opamp_dummy_magic_0.V_p.n14 two_stage_opamp_dummy_magic_0.V_p.n12 0.563
R8176 two_stage_opamp_dummy_magic_0.V_p.n16 two_stage_opamp_dummy_magic_0.V_p.n14 0.563
R8177 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n16 0.563
R8178 two_stage_opamp_dummy_magic_0.V_p.n17 two_stage_opamp_dummy_magic_0.V_p.n2 0.563
R8179 two_stage_opamp_dummy_magic_0.V_p.n30 two_stage_opamp_dummy_magic_0.V_p.n28 0.563
R8180 two_stage_opamp_dummy_magic_0.V_p.n32 two_stage_opamp_dummy_magic_0.V_p.n30 0.563
R8181 two_stage_opamp_dummy_magic_0.V_p.n34 two_stage_opamp_dummy_magic_0.V_p.n32 0.563
R8182 two_stage_opamp_dummy_magic_0.V_p.n23 two_stage_opamp_dummy_magic_0.V_p.n21 0.563
R8183 two_stage_opamp_dummy_magic_0.V_p.n25 two_stage_opamp_dummy_magic_0.V_p.n23 0.563
R8184 two_stage_opamp_dummy_magic_0.V_p.n35 two_stage_opamp_dummy_magic_0.V_p.n25 0.53175
R8185 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 144.827
R8186 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 134.577
R8187 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 120.66
R8188 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 98.063
R8189 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 97.4009
R8190 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 96.8384
R8191 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 96.8384
R8192 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 96.8384
R8193 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 96.8384
R8194 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 24.0005
R8195 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 24.0005
R8196 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 24.0005
R8197 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 24.0005
R8198 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R8199 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 8.0005
R8200 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R8201 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R8202 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 8.0005
R8203 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R8204 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R8205 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 8.0005
R8206 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R8207 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 8.0005
R8208 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 5.813
R8209 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 1.46925
R8210 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 0.563
R8211 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 0.563
R8212 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 0.563
R8213 VIN-.n4 VIN-.t8 485.021
R8214 VIN-.n1 VIN-.t6 484.159
R8215 VIN-.n5 VIN-.t7 483.358
R8216 VIN-.n8 VIN-.t10 431.536
R8217 VIN-.n2 VIN-.t9 431.536
R8218 VIN-.n6 VIN-.t1 431.257
R8219 VIN-.n0 VIN-.t0 431.257
R8220 VIN-.n6 VIN-.t2 289.908
R8221 VIN-.n0 VIN-.t5 289.908
R8222 VIN-.n8 VIN-.t4 279.183
R8223 VIN-.n2 VIN-.t3 279.183
R8224 VIN-.n7 VIN-.n6 233.374
R8225 VIN-.n1 VIN-.n0 233.374
R8226 VIN-.n9 VIN-.n8 188.989
R8227 VIN-.n3 VIN-.n2 188.989
R8228 VIN-.n4 VIN-.n3 2.463
R8229 VIN- VIN-.n9 1.78175
R8230 VIN-.n5 VIN-.n4 1.563
R8231 VIN-.n3 VIN-.n1 1.2755
R8232 VIN-.n9 VIN-.n7 1.2755
R8233 VIN-.n7 VIN-.n5 0.8005
R8234 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t12 668.604
R8235 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 631.982
R8236 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n3 627.128
R8237 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 627.128
R8238 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 226.534
R8239 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 226.534
R8240 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n4 222.034
R8241 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R8242 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R8243 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R8244 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t4 78.8005
R8245 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t6 78.8005
R8246 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t5 78.8005
R8247 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R8248 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t10 48.0005
R8249 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R8250 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t0 48.0005
R8251 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R8252 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t11 48.0005
R8253 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 8.938
R8254 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 5.7505
R8255 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.313
R8256 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 1.2505
R8257 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n9 160.428
R8258 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n0 160.427
R8259 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 159.803
R8260 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n14 159.803
R8261 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n12 159.803
R8262 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 159.803
R8263 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 159.802
R8264 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 159.802
R8265 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.n3 159.802
R8266 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n1 159.802
R8267 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.n18 159.798
R8268 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n17 14.438
R8269 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t9 11.2576
R8270 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t11 11.2576
R8271 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t12 11.2576
R8272 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.t4 11.2576
R8273 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.t13 11.2576
R8274 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R8275 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t7 11.2576
R8276 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R8277 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R8278 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.t5 11.2576
R8279 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t15 11.2576
R8280 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t17 11.2576
R8281 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t2 11.2576
R8282 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R8283 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.t16 11.2576
R8284 two_stage_opamp_dummy_magic_0.VD4.n3 two_stage_opamp_dummy_magic_0.VD4.t14 11.2576
R8285 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R8286 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t3 11.2576
R8287 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t18 11.2576
R8288 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t1 11.2576
R8289 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t20 11.2576
R8290 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.n19 11.2576
R8291 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n11 0.6255
R8292 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n13 0.6255
R8293 two_stage_opamp_dummy_magic_0.VD4.n4 two_stage_opamp_dummy_magic_0.VD4.n2 0.6255
R8294 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n4 0.6255
R8295 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n6 0.6255
R8296 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n8 0.6255
R8297 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 0.5005
R8298 w_10220_8260.n7 w_10220_8260.n2 4020
R8299 w_10220_8260.n9 w_10220_8260.n2 4020
R8300 w_10220_8260.n9 w_10220_8260.n3 4020
R8301 w_10220_8260.n7 w_10220_8260.n3 4020
R8302 w_10220_8260.n12 w_10220_8260.t0 660.109
R8303 w_10220_8260.n4 w_10220_8260.t3 660.109
R8304 w_10220_8260.n6 w_10220_8260.n1 428.8
R8305 w_10220_8260.n10 w_10220_8260.n1 428.8
R8306 w_10220_8260.t4 w_10220_8260.n7 239.915
R8307 w_10220_8260.n9 w_10220_8260.t1 239.915
R8308 w_10220_8260.n5 w_10220_8260.n0 230.4
R8309 w_10220_8260.n11 w_10220_8260.n0 230.4
R8310 w_10220_8260.n6 w_10220_8260.n5 198.4
R8311 w_10220_8260.n11 w_10220_8260.n10 198.4
R8312 w_10220_8260.n4 w_10220_8260.t5 155.125
R8313 w_10220_8260.t2 w_10220_8260.n12 155.125
R8314 w_10220_8260.t6 w_10220_8260.t4 98.2764
R8315 w_10220_8260.t9 w_10220_8260.t6 98.2764
R8316 w_10220_8260.t13 w_10220_8260.t9 98.2764
R8317 w_10220_8260.t11 w_10220_8260.t13 98.2764
R8318 w_10220_8260.t14 w_10220_8260.t11 98.2764
R8319 w_10220_8260.t7 w_10220_8260.t15 98.2764
R8320 w_10220_8260.t10 w_10220_8260.t7 98.2764
R8321 w_10220_8260.t8 w_10220_8260.t10 98.2764
R8322 w_10220_8260.t12 w_10220_8260.t8 98.2764
R8323 w_10220_8260.t1 w_10220_8260.t12 98.2764
R8324 w_10220_8260.n7 w_10220_8260.n6 92.5005
R8325 w_10220_8260.n2 w_10220_8260.n1 92.5005
R8326 w_10220_8260.n8 w_10220_8260.n2 92.5005
R8327 w_10220_8260.n10 w_10220_8260.n9 92.5005
R8328 w_10220_8260.n3 w_10220_8260.n0 92.5005
R8329 w_10220_8260.n8 w_10220_8260.n3 92.5005
R8330 w_10220_8260.n8 w_10220_8260.t14 49.1384
R8331 w_10220_8260.t15 w_10220_8260.n8 49.1384
R8332 w_10220_8260.n5 w_10220_8260.n4 21.3338
R8333 w_10220_8260.n12 w_10220_8260.n11 21.3338
R8334 a_10480_8490.n5 a_10480_8490.n3 160.427
R8335 a_10480_8490.n2 a_10480_8490.n0 160.427
R8336 a_10480_8490.n7 a_10480_8490.n6 159.802
R8337 a_10480_8490.n5 a_10480_8490.n4 159.802
R8338 a_10480_8490.n2 a_10480_8490.n1 159.802
R8339 a_10480_8490.n9 a_10480_8490.n8 159.798
R8340 a_10480_8490.n6 a_10480_8490.t11 11.2576
R8341 a_10480_8490.n6 a_10480_8490.t3 11.2576
R8342 a_10480_8490.n4 a_10480_8490.t6 11.2576
R8343 a_10480_8490.n4 a_10480_8490.t4 11.2576
R8344 a_10480_8490.n3 a_10480_8490.t8 11.2576
R8345 a_10480_8490.n3 a_10480_8490.t0 11.2576
R8346 a_10480_8490.n1 a_10480_8490.t5 11.2576
R8347 a_10480_8490.n1 a_10480_8490.t9 11.2576
R8348 a_10480_8490.n0 a_10480_8490.t1 11.2576
R8349 a_10480_8490.n0 a_10480_8490.t2 11.2576
R8350 a_10480_8490.n9 a_10480_8490.t7 11.2576
R8351 a_10480_8490.t10 a_10480_8490.n9 11.2576
R8352 a_10480_8490.n7 a_10480_8490.n5 0.6255
R8353 a_10480_8490.n8 a_10480_8490.n7 0.6255
R8354 a_10480_8490.n8 a_10480_8490.n2 0.6255
R8355 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.t20 619.201
R8356 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t12 611.739
R8357 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t25 611.739
R8358 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R8359 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t21 611.739
R8360 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R8361 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R8362 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R8363 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R8364 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R8365 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R8366 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R8367 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R8368 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R8369 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R8370 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t26 421.75
R8371 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R8372 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R8373 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R8374 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R8375 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R8376 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 176.155
R8377 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n13 175.79
R8378 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 172.667
R8379 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R8380 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R8381 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R8382 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R8383 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R8384 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R8385 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R8386 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R8387 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R8388 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R8389 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R8390 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R8391 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n1 139.639
R8392 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 139.638
R8393 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n0 134.577
R8394 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 106.891
R8395 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 47.1294
R8396 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n17 47.1294
R8397 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 47.1294
R8398 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n8 47.1294
R8399 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R8400 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t6 24.0005
R8401 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R8402 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t0 24.0005
R8403 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R8404 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R8405 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t1 10.9449
R8406 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t2 10.9449
R8407 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 9.5005
R8408 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n24 8.79738
R8409 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 4.5005
R8410 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 0.96925
R8411 a_11220_17410.t0 a_11220_17410.t1 258.591
R8412 a_5750_2276.t0 a_5750_2276.t1 169.905
R8413 a_14640_5068.t0 a_14640_5068.t1 169.905
R8414 VIN+.n9 VIN+.t5 485.127
R8415 VIN+.n4 VIN+.t3 485.127
R8416 VIN+.n3 VIN+.t4 485.127
R8417 VIN+.n7 VIN+.t9 318.656
R8418 VIN+.n7 VIN+.t2 318.656
R8419 VIN+.n5 VIN+.t7 318.656
R8420 VIN+.n5 VIN+.t1 318.656
R8421 VIN+.n1 VIN+.t8 318.656
R8422 VIN+.n1 VIN+.t6 318.656
R8423 VIN+.n0 VIN+.t10 318.656
R8424 VIN+.n0 VIN+.t0 318.656
R8425 VIN+.n2 VIN+.n0 167.05
R8426 VIN+.n8 VIN+.n7 165.8
R8427 VIN+.n6 VIN+.n5 165.8
R8428 VIN+.n2 VIN+.n1 165.8
R8429 VIN+.n6 VIN+.n4 2.34425
R8430 VIN+.n4 VIN+.n3 1.3005
R8431 VIN+.n8 VIN+.n6 1.2505
R8432 VIN+.n3 VIN+.n2 1.15675
R8433 VIN+.n9 VIN+.n8 1.15675
R8434 VIN+ VIN+.n9 0.963
R8435 a_13730_17020.t0 a_13730_17020.t1 258.591
R8436 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R8437 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R8438 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t3 303.259
R8439 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R8440 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R8441 bgr_0.V_CUR_REF_REG.t1 bgr_0.V_CUR_REF_REG.n5 245.284
R8442 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t7 174.726
R8443 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 174.726
R8444 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R8445 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R8446 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 96.4005
R8447 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t2 39.4005
R8448 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t0 39.4005
R8449 a_12828_17530.t0 a_12828_17530.t1 376.99
R8450 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8451 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8452 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8453 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8454 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8455 bgr_0.START_UP.n0 bgr_0.START_UP.t5 130.001
R8456 bgr_0.START_UP.n0 bgr_0.START_UP.t4 81.7074
R8457 bgr_0.START_UP bgr_0.START_UP.n0 38.2614
R8458 bgr_0.START_UP bgr_0.START_UP.n5 14.7817
R8459 bgr_0.START_UP.n1 bgr_0.START_UP.t0 13.1338
R8460 bgr_0.START_UP.n1 bgr_0.START_UP.t1 13.1338
R8461 bgr_0.START_UP.n2 bgr_0.START_UP.t2 13.1338
R8462 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8463 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8464 a_11220_17290.t0 a_11220_17290.t1 376.99
R8465 a_12828_17650.t0 a_12828_17650.t1 258.591
R8466 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8467 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2595
R8468 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2280
R8469 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2250
R8470 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 672.159
R8471 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 672.159
R8472 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 276.8
R8473 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 240
R8474 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 206.4
R8475 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 204.8
R8476 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 180.904
R8477 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 170.3
R8478 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 160.517
R8479 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 160.517
R8480 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 110.425
R8481 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 110.05
R8482 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 95.7988
R8483 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8484 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8485 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8486 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8487 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8488 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8489 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 76.8005
R8490 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 75.9449
R8491 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 75.9449
R8492 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 47.8997
R8493 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 47.8997
R8494 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 38.4005
R8495 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 24.5338
R8496 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 24.5338
R8497 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 16.8187
R8498 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 16.8187
R8499 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 12.313
R8500 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 12.313
R8501 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 10.9449
R8502 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 10.9449
R8503 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8504 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8505 a_5230_5088.t0 a_5230_5088.t1 294.339
R8506 a_14240_2276.t0 a_14240_2276.t1 169.905
R8507 a_13790_17550.t0 a_13790_17550.t1 258.591
R8508 a_5350_5088.t0 a_5350_5088.t1 169.905
C0 two_stage_opamp_dummy_magic_0.V_err_gate bgr_0.TAIL_CUR_MIR_BIAS 0.039198f
C1 bgr_0.PFET_GATE_10uA bgr_0.1st_Vout_1 0.035393f
C2 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.err_amp_out 0.425326f
C3 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.cap_res_X 0.790473f
C4 VDDA two_stage_opamp_dummy_magic_0.err_amp_out 1.20093f
C5 VIN+ two_stage_opamp_dummy_magic_0.VD1 0.058217f
C6 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.err_amp_out 0.253351f
C7 two_stage_opamp_dummy_magic_0.Vb2_Vb3 VDDA 0.875085f
C8 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.Vb2_Vb3 0.065464f
C9 VDDA two_stage_opamp_dummy_magic_0.Y 3.97699f
C10 bgr_0.cap_res2 VDDA 0.58582f
C11 bgr_0.1st_Vout_1 m2_8540_19780# 0.075543f
C12 bgr_0.NFET_GATE_10uA VDDA 1.04958f
C13 two_stage_opamp_dummy_magic_0.V_err_gate bgr_0.NFET_GATE_10uA 0.136183f
C14 two_stage_opamp_dummy_magic_0.V_err_gate VDDA 5.0275f
C15 bgr_0.START_UP bgr_0.NFET_GATE_10uA 0.518732f
C16 bgr_0.TAIL_CUR_MIR_BIAS VIN- 0.306616f
C17 bgr_0.START_UP VDDA 1.37392f
C18 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 2.47368f
C19 two_stage_opamp_dummy_magic_0.Y a_10530_5140# 0.829736f
C20 bgr_0.PFET_GATE_10uA m2_7180_19780# 0.012f
C21 bgr_0.Vbe2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.014154f
C22 bgr_0.PFET_GATE_10uA bgr_0.TAIL_CUR_MIR_BIAS 0.213841f
C23 bgr_0.cap_res2 li_10610_16720# 0.020538f
C24 bgr_0.TAIL_CUR_MIR_BIAS VIN+ 0.111541f
C25 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.1st_Vout_1 0.477103f
C26 bgr_0.V_TOP m2_8540_19780# 0.012f
C27 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.VD3 0.363482f
C28 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.cap_res_X 0.442088f
C29 bgr_0.PFET_GATE_10uA bgr_0.cap_res2 0.018633f
C30 bgr_0.PFET_GATE_10uA bgr_0.NFET_GATE_10uA 0.050552f
C31 bgr_0.PFET_GATE_10uA VDDA 10.3925f
C32 VDDA li_7110_16510# 0.021911f
C33 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.13839f
C34 bgr_0.START_UP bgr_0.PFET_GATE_10uA 0.166283f
C35 bgr_0.TAIL_CUR_MIR_BIAS a_11120_2960# 0.012f
C36 VDDA two_stage_opamp_dummy_magic_0.VD3 3.95386f
C37 bgr_0.cap_res2 two_stage_opamp_dummy_magic_0.cap_res_X 0.048779f
C38 VDDA m2_8540_19780# 0.010446f
C39 VDDA two_stage_opamp_dummy_magic_0.cap_res_X 0.921518f
C40 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.TAIL_CUR_MIR_BIAS 3.74826f
C41 bgr_0.Vbe2 bgr_0.V_TOP 0.285619f
C42 two_stage_opamp_dummy_magic_0.err_amp_out a_11120_2960# 0.012f
C43 bgr_0.V_TOP bgr_0.1st_Vout_1 0.925484f
C44 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.err_amp_out 0.528215f
C45 VIN- VIN+ 0.562828f
C46 bgr_0.V_TOP li_5710_16610# 0.020062f
C47 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.cap_res2 0.551434f
C48 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.VD1 0.92136f
C49 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.NFET_GATE_10uA 0.559544f
C50 bgr_0.START_UP_NFET1 bgr_0.NFET_GATE_10uA 0.318695f
C51 two_stage_opamp_dummy_magic_0.V_err_amp_ref VDDA 4.37237f
C52 bgr_0.START_UP_NFET1 VDDA 0.150608f
C53 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.37399f
C54 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.09763f
C55 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C56 bgr_0.Vbe2 bgr_0.NFET_GATE_10uA 0.021455f
C57 bgr_0.Vbe2 VDDA 0.016701f
C58 bgr_0.1st_Vout_1 bgr_0.cap_res2 0.822981f
C59 bgr_0.NFET_GATE_10uA bgr_0.1st_Vout_1 1.02268f
C60 two_stage_opamp_dummy_magic_0.Y two_stage_opamp_dummy_magic_0.VD1 1.05325f
C61 bgr_0.1st_Vout_1 VDDA 2.06087f
C62 bgr_0.START_UP bgr_0.Vbe2 0.193132f
C63 bgr_0.V_TOP bgr_0.TAIL_CUR_MIR_BIAS 0.036996f
C64 bgr_0.START_UP bgr_0.1st_Vout_1 0.030647f
C65 two_stage_opamp_dummy_magic_0.VD3 two_stage_opamp_dummy_magic_0.cap_res_X 0.033524f
C66 a_10530_5140# two_stage_opamp_dummy_magic_0.VD1 0.349817f
C67 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.err_amp_out 0.010868f
C68 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.46518f
C69 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.080353f
C70 bgr_0.V_TOP VDDA 16.1354f
C71 VDDA m2_7180_19780# 0.010446f
C72 VIN- two_stage_opamp_dummy_magic_0.VD1 0.881216f
C73 bgr_0.1st_Vout_1 li_12710_16610# 0.020439f
C74 bgr_0.Vbe2 bgr_0.PFET_GATE_10uA 0.242909f
C75 bgr_0.START_UP bgr_0.V_TOP 0.815644f
C76 bgr_0.NFET_GATE_10uA bgr_0.TAIL_CUR_MIR_BIAS 0.064423f
C77 bgr_0.TAIL_CUR_MIR_BIAS VDDA 5.87048f
C78 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.VD3 0.102485f
C79 VOUT+ GNDA 0.038145f
C80 VOUT- GNDA 0.038151f
C81 VIN+ GNDA 2.062944f
C82 VIN- GNDA 2.127458f
C83 VDDA GNDA 0.151107p
C84 li_7110_16510# GNDA 0.050654f $ **FLOATING
C85 li_14110_16610# GNDA 0.050514f $ **FLOATING
C86 li_12710_16610# GNDA 0.049721f $ **FLOATING
C87 li_5710_16610# GNDA 0.047034f $ **FLOATING
C88 li_10610_16720# GNDA 0.049096f $ **FLOATING
C89 li_9210_16720# GNDA 0.043891f $ **FLOATING
C90 a_11120_2960# GNDA 0.110549f
C91 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.43445f
C92 a_10530_5140# GNDA 1.24614f
C93 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.373356f
C94 two_stage_opamp_dummy_magic_0.Y GNDA 5.133595f
C95 two_stage_opamp_dummy_magic_0.cap_res_X GNDA 33.15933f
C96 two_stage_opamp_dummy_magic_0.VD3 GNDA 0.365122f
C97 bgr_0.cap_res2 GNDA 7.936877f
C98 bgr_0.TAIL_CUR_MIR_BIAS GNDA 10.97818f
C99 bgr_0.1st_Vout_1 GNDA 4.986571f
C100 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 15.217911f
C101 bgr_0.V_TOP GNDA 6.838887f
C102 bgr_0.PFET_GATE_10uA GNDA 5.13254f
C103 bgr_0.Vbe2 GNDA 17.0659f
C104 bgr_0.START_UP GNDA 7.190383f
C105 bgr_0.START_UP_NFET1 GNDA 5.28339f
C106 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 15.080791f
C107 bgr_0.NFET_GATE_10uA GNDA 7.08898f
C108 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.6041f
C109 bgr_0.START_UP.t4 GNDA 1.6623f
C110 bgr_0.START_UP.t5 GNDA 0.043697f
C111 bgr_0.START_UP.n0 GNDA 1.12862f
C112 bgr_0.START_UP.t0 GNDA 0.041701f
C113 bgr_0.START_UP.t1 GNDA 0.041701f
C114 bgr_0.START_UP.n1 GNDA 0.151283f
C115 bgr_0.START_UP.t2 GNDA 0.041701f
C116 bgr_0.START_UP.t3 GNDA 0.041701f
C117 bgr_0.START_UP.n2 GNDA 0.139173f
C118 bgr_0.START_UP.n3 GNDA 0.720787f
C119 bgr_0.START_UP.t7 GNDA 0.01567f
C120 bgr_0.START_UP.t6 GNDA 0.01567f
C121 bgr_0.START_UP.n4 GNDA 0.044238f
C122 bgr_0.START_UP.n5 GNDA 0.445182f
C123 bgr_0.V_CUR_REF_REG.t3 GNDA 0.014208f
C124 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C125 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C126 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C127 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C128 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C129 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C130 bgr_0.V_CUR_REF_REG.t1 GNDA 0.42777f
C131 VIN+.t0 GNDA 0.042021f
C132 VIN+.t10 GNDA 0.042021f
C133 VIN+.n0 GNDA 0.086842f
C134 VIN+.t6 GNDA 0.042021f
C135 VIN+.t8 GNDA 0.042021f
C136 VIN+.n1 GNDA 0.085639f
C137 VIN+.n2 GNDA 0.361638f
C138 VIN+.t4 GNDA 0.059118f
C139 VIN+.n3 GNDA 0.216459f
C140 VIN+.t3 GNDA 0.059118f
C141 VIN+.n4 GNDA 0.263959f
C142 VIN+.t1 GNDA 0.042021f
C143 VIN+.t7 GNDA 0.042021f
C144 VIN+.n5 GNDA 0.085639f
C145 VIN+.n6 GNDA 0.249653f
C146 VIN+.t2 GNDA 0.042021f
C147 VIN+.t9 GNDA 0.042021f
C148 VIN+.n7 GNDA 0.085639f
C149 VIN+.n8 GNDA 0.202005f
C150 VIN+.t5 GNDA 0.059118f
C151 VIN+.n9 GNDA 0.202625f
C152 bgr_0.VB3_CUR_BIAS GNDA 4.60549f
C153 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.031172f
C154 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.031172f
C155 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.094152f
C156 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.031172f
C157 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.031172f
C158 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.100408f
C159 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.031172f
C160 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.031172f
C161 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.100408f
C162 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.553544f
C163 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.206656f
C164 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.177535f
C165 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.154301f
C166 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.154301f
C167 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.154301f
C168 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.154301f
C169 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.178062f
C170 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.144567f
C171 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.08884f
C172 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.08884f
C173 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.083186f
C174 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.154301f
C175 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.154301f
C176 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.154301f
C177 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.154301f
C178 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.178062f
C179 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.144567f
C180 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.08884f
C181 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.08884f
C182 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.083186f
C183 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.086286f
C184 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.154301f
C185 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.154301f
C186 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.154301f
C187 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.154301f
C188 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.178062f
C189 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.144567f
C190 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.08884f
C191 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.08884f
C192 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.083186f
C193 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.154301f
C194 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.154301f
C195 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.154301f
C196 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.154301f
C197 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.178062f
C198 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.144567f
C199 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.08884f
C200 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.08884f
C201 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.083186f
C202 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.089524f
C203 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 2.44739f
C204 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.682611f
C205 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.112219f
C206 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.112219f
C207 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.401639f
C208 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 4.9401f
C209 a_10480_8490.t7 GNDA 0.043655f
C210 a_10480_8490.t1 GNDA 0.043655f
C211 a_10480_8490.t2 GNDA 0.043655f
C212 a_10480_8490.n0 GNDA 0.151823f
C213 a_10480_8490.t5 GNDA 0.043655f
C214 a_10480_8490.t9 GNDA 0.043655f
C215 a_10480_8490.n1 GNDA 0.151285f
C216 a_10480_8490.n2 GNDA 0.285611f
C217 a_10480_8490.t8 GNDA 0.043655f
C218 a_10480_8490.t0 GNDA 0.043655f
C219 a_10480_8490.n3 GNDA 0.151823f
C220 a_10480_8490.t6 GNDA 0.043655f
C221 a_10480_8490.t4 GNDA 0.043655f
C222 a_10480_8490.n4 GNDA 0.151285f
C223 a_10480_8490.n5 GNDA 0.285612f
C224 a_10480_8490.t11 GNDA 0.043655f
C225 a_10480_8490.t3 GNDA 0.043655f
C226 a_10480_8490.n6 GNDA 0.151285f
C227 a_10480_8490.n7 GNDA 0.148064f
C228 a_10480_8490.n8 GNDA 0.148064f
C229 a_10480_8490.n9 GNDA 0.151285f
C230 a_10480_8490.t10 GNDA 0.043655f
C231 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.061318f
C232 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.061318f
C233 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.061318f
C234 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.213252f
C235 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.061318f
C236 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.061318f
C237 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.212496f
C238 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.401171f
C239 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.061318f
C240 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.061318f
C241 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.212496f
C242 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.207971f
C243 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.061318f
C244 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.061318f
C245 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.212496f
C246 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.207971f
C247 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.061318f
C248 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.061318f
C249 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.212496f
C250 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.207971f
C251 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.061318f
C252 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.061318f
C253 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.213251f
C254 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.061318f
C255 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.061318f
C256 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.212496f
C257 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.401172f
C258 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.061318f
C259 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.061318f
C260 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.212496f
C261 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.207971f
C262 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.061318f
C263 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.061318f
C264 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.212496f
C265 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.200964f
C266 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.061318f
C267 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.061318f
C268 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.212496f
C269 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.381399f
C270 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.395445f
C271 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.212496f
C272 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.061318f
C273 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.017507f
C274 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.017316f
C275 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.345034f
C276 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.017316f
C277 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.019333f
C278 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.068944f
C279 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 0.020653f
C280 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 1.01255f
C281 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.020653f
C282 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.181418f
C283 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.176738f
C284 VIN-.t6 GNDA 0.050911f
C285 VIN-.t5 GNDA 0.03359f
C286 VIN-.t0 GNDA 0.04147f
C287 VIN-.n0 GNDA 0.05959f
C288 VIN-.n1 GNDA 0.281971f
C289 VIN-.t3 GNDA 0.033038f
C290 VIN-.t9 GNDA 0.041485f
C291 VIN-.n2 GNDA 0.065237f
C292 VIN-.n3 GNDA 0.201948f
C293 VIN-.t8 GNDA 0.050345f
C294 VIN-.n4 GNDA 0.237498f
C295 VIN-.t7 GNDA 0.050694f
C296 VIN-.n5 GNDA 0.181582f
C297 VIN-.t2 GNDA 0.03359f
C298 VIN-.t1 GNDA 0.04147f
C299 VIN-.n6 GNDA 0.05959f
C300 VIN-.n7 GNDA 0.150425f
C301 VIN-.t4 GNDA 0.033038f
C302 VIN-.t10 GNDA 0.041485f
C303 VIN-.n8 GNDA 0.065237f
C304 VIN-.n9 GNDA 0.178598f
C305 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.425414f
C306 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.102505f
C307 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.102505f
C308 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.423897f
C309 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.102505f
C310 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.102505f
C311 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.422271f
C312 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.585479f
C313 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.102505f
C314 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.102505f
C315 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.422271f
C316 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.305512f
C317 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.102505f
C318 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.102505f
C319 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.422271f
C320 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.305512f
C321 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.102505f
C322 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.102505f
C323 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.422271f
C324 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.439098f
C325 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 5.50033f
C326 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.034168f
C327 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.034168f
C328 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.124192f
C329 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.034168f
C330 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.034168f
C331 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.103202f
C332 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.645167f
C333 bgr_0.V_CMFB_S2 GNDA 4.4914f
C334 two_stage_opamp_dummy_magic_0.V_p.t28 GNDA 0.024537f
C335 two_stage_opamp_dummy_magic_0.V_p.t21 GNDA 0.024537f
C336 two_stage_opamp_dummy_magic_0.V_p.t6 GNDA 0.024537f
C337 two_stage_opamp_dummy_magic_0.V_p.n0 GNDA 0.097795f
C338 two_stage_opamp_dummy_magic_0.V_p.t38 GNDA 0.024537f
C339 two_stage_opamp_dummy_magic_0.V_p.t32 GNDA 0.024537f
C340 two_stage_opamp_dummy_magic_0.V_p.n1 GNDA 0.097424f
C341 two_stage_opamp_dummy_magic_0.V_p.n2 GNDA 0.164007f
C342 two_stage_opamp_dummy_magic_0.V_p.t25 GNDA 0.024537f
C343 two_stage_opamp_dummy_magic_0.V_p.t31 GNDA 0.024537f
C344 two_stage_opamp_dummy_magic_0.V_p.n3 GNDA 0.097877f
C345 two_stage_opamp_dummy_magic_0.V_p.t27 GNDA 0.024537f
C346 two_stage_opamp_dummy_magic_0.V_p.t35 GNDA 0.024537f
C347 two_stage_opamp_dummy_magic_0.V_p.n4 GNDA 0.097424f
C348 two_stage_opamp_dummy_magic_0.V_p.n5 GNDA 0.166869f
C349 two_stage_opamp_dummy_magic_0.V_p.t29 GNDA 0.024537f
C350 two_stage_opamp_dummy_magic_0.V_p.t37 GNDA 0.024537f
C351 two_stage_opamp_dummy_magic_0.V_p.n6 GNDA 0.097424f
C352 two_stage_opamp_dummy_magic_0.V_p.n7 GNDA 0.087096f
C353 two_stage_opamp_dummy_magic_0.V_p.t9 GNDA 0.102522f
C354 two_stage_opamp_dummy_magic_0.V_p.t33 GNDA 0.024537f
C355 two_stage_opamp_dummy_magic_0.V_p.t23 GNDA 0.024537f
C356 two_stage_opamp_dummy_magic_0.V_p.n8 GNDA 0.094681f
C357 two_stage_opamp_dummy_magic_0.V_p.n9 GNDA 0.675343f
C358 two_stage_opamp_dummy_magic_0.V_p.n10 GNDA 0.029445f
C359 two_stage_opamp_dummy_magic_0.V_p.t30 GNDA 0.024537f
C360 two_stage_opamp_dummy_magic_0.V_p.t22 GNDA 0.024537f
C361 two_stage_opamp_dummy_magic_0.V_p.n11 GNDA 0.097424f
C362 two_stage_opamp_dummy_magic_0.V_p.n12 GNDA 0.087096f
C363 two_stage_opamp_dummy_magic_0.V_p.t34 GNDA 0.024537f
C364 two_stage_opamp_dummy_magic_0.V_p.t24 GNDA 0.024537f
C365 two_stage_opamp_dummy_magic_0.V_p.n13 GNDA 0.097424f
C366 two_stage_opamp_dummy_magic_0.V_p.n14 GNDA 0.087096f
C367 two_stage_opamp_dummy_magic_0.V_p.t36 GNDA 0.024537f
C368 two_stage_opamp_dummy_magic_0.V_p.t26 GNDA 0.024537f
C369 two_stage_opamp_dummy_magic_0.V_p.n15 GNDA 0.097424f
C370 two_stage_opamp_dummy_magic_0.V_p.n16 GNDA 0.087096f
C371 two_stage_opamp_dummy_magic_0.V_p.n17 GNDA 0.029445f
C372 two_stage_opamp_dummy_magic_0.V_p.t0 GNDA 0.014722f
C373 two_stage_opamp_dummy_magic_0.V_p.t12 GNDA 0.014722f
C374 two_stage_opamp_dummy_magic_0.V_p.n18 GNDA 0.050019f
C375 two_stage_opamp_dummy_magic_0.V_p.t14 GNDA 0.014722f
C376 two_stage_opamp_dummy_magic_0.V_p.t5 GNDA 0.014722f
C377 two_stage_opamp_dummy_magic_0.V_p.n19 GNDA 0.052892f
C378 two_stage_opamp_dummy_magic_0.V_p.t20 GNDA 0.014722f
C379 two_stage_opamp_dummy_magic_0.V_p.t3 GNDA 0.014722f
C380 two_stage_opamp_dummy_magic_0.V_p.n20 GNDA 0.052484f
C381 two_stage_opamp_dummy_magic_0.V_p.n21 GNDA 0.17749f
C382 two_stage_opamp_dummy_magic_0.V_p.t15 GNDA 0.014722f
C383 two_stage_opamp_dummy_magic_0.V_p.t7 GNDA 0.014722f
C384 two_stage_opamp_dummy_magic_0.V_p.n22 GNDA 0.052484f
C385 two_stage_opamp_dummy_magic_0.V_p.n23 GNDA 0.092385f
C386 two_stage_opamp_dummy_magic_0.V_p.t11 GNDA 0.014722f
C387 two_stage_opamp_dummy_magic_0.V_p.t10 GNDA 0.014722f
C388 two_stage_opamp_dummy_magic_0.V_p.n24 GNDA 0.052484f
C389 two_stage_opamp_dummy_magic_0.V_p.n25 GNDA 0.091894f
C390 two_stage_opamp_dummy_magic_0.V_p.t1 GNDA 0.014722f
C391 two_stage_opamp_dummy_magic_0.V_p.t13 GNDA 0.014722f
C392 two_stage_opamp_dummy_magic_0.V_p.n26 GNDA 0.052869f
C393 two_stage_opamp_dummy_magic_0.V_p.t8 GNDA 0.014722f
C394 two_stage_opamp_dummy_magic_0.V_p.t19 GNDA 0.014722f
C395 two_stage_opamp_dummy_magic_0.V_p.n27 GNDA 0.052484f
C396 two_stage_opamp_dummy_magic_0.V_p.n28 GNDA 0.175746f
C397 two_stage_opamp_dummy_magic_0.V_p.t18 GNDA 0.014722f
C398 two_stage_opamp_dummy_magic_0.V_p.t4 GNDA 0.014722f
C399 two_stage_opamp_dummy_magic_0.V_p.n29 GNDA 0.052484f
C400 two_stage_opamp_dummy_magic_0.V_p.n30 GNDA 0.092385f
C401 two_stage_opamp_dummy_magic_0.V_p.t2 GNDA 0.014722f
C402 two_stage_opamp_dummy_magic_0.V_p.t40 GNDA 0.014722f
C403 two_stage_opamp_dummy_magic_0.V_p.n31 GNDA 0.052484f
C404 two_stage_opamp_dummy_magic_0.V_p.n32 GNDA 0.092385f
C405 two_stage_opamp_dummy_magic_0.V_p.t17 GNDA 0.014722f
C406 two_stage_opamp_dummy_magic_0.V_p.t16 GNDA 0.014722f
C407 two_stage_opamp_dummy_magic_0.V_p.n33 GNDA 0.052484f
C408 two_stage_opamp_dummy_magic_0.V_p.n34 GNDA 0.140968f
C409 two_stage_opamp_dummy_magic_0.V_p.n35 GNDA 0.077538f
C410 two_stage_opamp_dummy_magic_0.V_p.n36 GNDA 0.082969f
C411 two_stage_opamp_dummy_magic_0.V_p.n37 GNDA 0.082287f
C412 two_stage_opamp_dummy_magic_0.V_p.n38 GNDA 0.094681f
C413 two_stage_opamp_dummy_magic_0.V_p.t39 GNDA 0.024537f
C414 bgr_0.cap_res2.t6 GNDA 0.406156f
C415 bgr_0.cap_res2.t2 GNDA 0.407628f
C416 bgr_0.cap_res2.t8 GNDA 0.406156f
C417 bgr_0.cap_res2.t13 GNDA 0.407628f
C418 bgr_0.cap_res2.t0 GNDA 0.406156f
C419 bgr_0.cap_res2.t19 GNDA 0.407628f
C420 bgr_0.cap_res2.t1 GNDA 0.406156f
C421 bgr_0.cap_res2.t5 GNDA 0.407628f
C422 bgr_0.cap_res2.t7 GNDA 0.406156f
C423 bgr_0.cap_res2.t4 GNDA 0.407628f
C424 bgr_0.cap_res2.t10 GNDA 0.406156f
C425 bgr_0.cap_res2.t14 GNDA 0.407628f
C426 bgr_0.cap_res2.t15 GNDA 0.406156f
C427 bgr_0.cap_res2.t12 GNDA 0.407628f
C428 bgr_0.cap_res2.t16 GNDA 0.406156f
C429 bgr_0.cap_res2.t18 GNDA 0.407628f
C430 bgr_0.cap_res2.n0 GNDA 0.272247f
C431 bgr_0.cap_res2.t17 GNDA 0.216805f
C432 bgr_0.cap_res2.n1 GNDA 0.295394f
C433 bgr_0.cap_res2.t11 GNDA 0.216805f
C434 bgr_0.cap_res2.n2 GNDA 0.295394f
C435 bgr_0.cap_res2.t3 GNDA 0.216805f
C436 bgr_0.cap_res2.n3 GNDA 0.295394f
C437 bgr_0.cap_res2.t9 GNDA 0.214043f
C438 bgr_0.cap_res2.t20 GNDA 0.133038f
C439 bgr_0.1st_Vout_2.n0 GNDA 0.995956f
C440 bgr_0.1st_Vout_2.n1 GNDA 0.240335f
C441 bgr_0.1st_Vout_2.n2 GNDA 0.995956f
C442 bgr_0.1st_Vout_2.n3 GNDA 0.240335f
C443 bgr_0.1st_Vout_2.n4 GNDA 0.805677f
C444 bgr_0.1st_Vout_2.n5 GNDA 0.240335f
C445 bgr_0.1st_Vout_2.t13 GNDA 0.021508f
C446 bgr_0.1st_Vout_2.n6 GNDA 0.02259f
C447 bgr_0.1st_Vout_2.n7 GNDA 0.171874f
C448 bgr_0.1st_Vout_2.t32 GNDA 0.013652f
C449 bgr_0.1st_Vout_2.t19 GNDA 0.013652f
C450 bgr_0.1st_Vout_2.n8 GNDA 0.03037f
C451 bgr_0.1st_Vout_2.n9 GNDA 0.083918f
C452 bgr_0.1st_Vout_2.n10 GNDA 0.012945f
C453 bgr_0.1st_Vout_2.t8 GNDA 0.018875f
C454 bgr_0.1st_Vout_2.n11 GNDA 0.195802f
C455 bgr_0.1st_Vout_2.n12 GNDA 0.011712f
C456 bgr_0.1st_Vout_2.n13 GNDA 0.049674f
C457 bgr_0.1st_Vout_2.n14 GNDA 0.021654f
C458 bgr_0.1st_Vout_2.n15 GNDA 0.080059f
C459 bgr_0.1st_Vout_2.n16 GNDA 0.03943f
C460 bgr_0.1st_Vout_2.t36 GNDA 0.013652f
C461 bgr_0.1st_Vout_2.t26 GNDA 0.013652f
C462 bgr_0.1st_Vout_2.n17 GNDA 0.03037f
C463 bgr_0.1st_Vout_2.n18 GNDA 0.083918f
C464 bgr_0.1st_Vout_2.t17 GNDA 0.364565f
C465 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C466 bgr_0.1st_Vout_2.t15 GNDA 0.358459f
C467 bgr_0.1st_Vout_2.t16 GNDA 0.364565f
C468 bgr_0.1st_Vout_2.t12 GNDA 0.358459f
C469 bgr_0.1st_Vout_2.t27 GNDA 0.364565f
C470 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C471 bgr_0.1st_Vout_2.t22 GNDA 0.358459f
C472 bgr_0.1st_Vout_2.t23 GNDA 0.364565f
C473 bgr_0.1st_Vout_2.t18 GNDA 0.358459f
C474 bgr_0.1st_Vout_2.t35 GNDA 0.364565f
C475 bgr_0.1st_Vout_2.t11 GNDA 0.358459f
C476 bgr_0.1st_Vout_2.t31 GNDA 0.358459f
C477 bgr_0.1st_Vout_2.t34 GNDA 0.364565f
C478 bgr_0.1st_Vout_2.t29 GNDA 0.358459f
C479 bgr_0.1st_Vout_2.t28 GNDA 0.364565f
C480 bgr_0.1st_Vout_2.t33 GNDA 0.358459f
C481 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C482 bgr_0.1st_Vout_2.t20 GNDA 0.358459f
C483 bgr_0.1st_Vout_2.t25 GNDA 0.358459f
C484 bgr_0.1st_Vout_2.t14 GNDA 0.023417f
C485 bgr_0.1st_Vout_2.n19 GNDA 0.516024f
C486 bgr_0.1st_Vout_2.n20 GNDA 0.106455f
C487 bgr_0.1st_Vout_2.n21 GNDA 0.02259f
C488 bgr_0.Vin+.t6 GNDA 0.020459f
C489 bgr_0.Vin+.t8 GNDA 0.013299f
C490 bgr_0.Vin+.n0 GNDA 0.04388f
C491 bgr_0.Vin+.t10 GNDA 0.013299f
C492 bgr_0.Vin+.n1 GNDA 0.034146f
C493 bgr_0.Vin+.t7 GNDA 0.013299f
C494 bgr_0.Vin+.n2 GNDA 0.034607f
C495 bgr_0.Vin+.n3 GNDA 0.074523f
C496 bgr_0.Vin+.t4 GNDA 0.043132f
C497 bgr_0.Vin+.t3 GNDA 0.043132f
C498 bgr_0.Vin+.n4 GNDA 0.144858f
C499 bgr_0.Vin+.t2 GNDA 0.043132f
C500 bgr_0.Vin+.t5 GNDA 0.043132f
C501 bgr_0.Vin+.n5 GNDA 0.142495f
C502 bgr_0.Vin+.n6 GNDA 0.656763f
C503 bgr_0.Vin+.n7 GNDA 0.71769f
C504 bgr_0.Vin+.t1 GNDA 0.137433f
C505 bgr_0.Vin+.n8 GNDA 0.446219f
C506 bgr_0.Vin+.t0 GNDA 0.125873f
C507 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.174475f
C508 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.435852f
C509 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.435852f
C510 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.517289f
C511 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.273228f
C512 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.17292f
C513 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.475244f
C514 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.159805f
C515 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.805343f
C516 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.475244f
C517 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.435852f
C518 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.435852f
C519 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.517289f
C520 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.273228f
C521 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.17292f
C522 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.159805f
C523 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.805323f
C524 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.174475f
C525 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.175672f
C526 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.187134f
C527 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.175672f
C528 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.867065f
C529 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.041343f
C530 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.040593f
C531 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.225382f
C532 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.021075f
C533 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.123074f
C534 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.021216f
C535 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.034546f
C536 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.202018f
C537 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.040593f
C538 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.144283f
C539 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.160783f
C540 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 1.41037f
C541 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.867885f
C542 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.187155f
C543 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.021118f
C544 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020212f
C545 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020262f
C546 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021093f
C547 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.020966f
C548 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.297859f
C549 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.020966f
C550 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.155369f
C551 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.020966f
C552 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.189616f
C553 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.160506f
C554 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.14076f
C555 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.241198f
C556 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.021118f
C557 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020826f
C558 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.326026f
C559 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020826f
C560 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.179554f
C561 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.179554f
C562 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020826f
C563 bgr_0.TAIL_CUR_MIR_BIAS.t5 GNDA 0.03008f
C564 bgr_0.TAIL_CUR_MIR_BIAS.t10 GNDA 0.03008f
C565 bgr_0.TAIL_CUR_MIR_BIAS.n0 GNDA 0.072545f
C566 bgr_0.TAIL_CUR_MIR_BIAS.t9 GNDA 0.03008f
C567 bgr_0.TAIL_CUR_MIR_BIAS.t6 GNDA 0.03008f
C568 bgr_0.TAIL_CUR_MIR_BIAS.n1 GNDA 0.075298f
C569 bgr_0.TAIL_CUR_MIR_BIAS.t11 GNDA 0.03008f
C570 bgr_0.TAIL_CUR_MIR_BIAS.t8 GNDA 0.03008f
C571 bgr_0.TAIL_CUR_MIR_BIAS.n2 GNDA 0.074895f
C572 bgr_0.TAIL_CUR_MIR_BIAS.n3 GNDA 0.50855f
C573 bgr_0.TAIL_CUR_MIR_BIAS.t7 GNDA 0.03008f
C574 bgr_0.TAIL_CUR_MIR_BIAS.t4 GNDA 0.03008f
C575 bgr_0.TAIL_CUR_MIR_BIAS.n4 GNDA 0.075298f
C576 bgr_0.TAIL_CUR_MIR_BIAS.n5 GNDA 0.333784f
C577 bgr_0.TAIL_CUR_MIR_BIAS.n6 GNDA 0.774051f
C578 bgr_0.TAIL_CUR_MIR_BIAS.t0 GNDA 0.045119f
C579 bgr_0.TAIL_CUR_MIR_BIAS.t2 GNDA 0.045119f
C580 bgr_0.TAIL_CUR_MIR_BIAS.n7 GNDA 0.163283f
C581 bgr_0.TAIL_CUR_MIR_BIAS.t31 GNDA 0.080087f
C582 bgr_0.TAIL_CUR_MIR_BIAS.t22 GNDA 0.080087f
C583 bgr_0.TAIL_CUR_MIR_BIAS.t28 GNDA 0.080087f
C584 bgr_0.TAIL_CUR_MIR_BIAS.t18 GNDA 0.080087f
C585 bgr_0.TAIL_CUR_MIR_BIAS.t26 GNDA 0.080087f
C586 bgr_0.TAIL_CUR_MIR_BIAS.t16 GNDA 0.080087f
C587 bgr_0.TAIL_CUR_MIR_BIAS.t24 GNDA 0.080087f
C588 bgr_0.TAIL_CUR_MIR_BIAS.t13 GNDA 0.080087f
C589 bgr_0.TAIL_CUR_MIR_BIAS.t20 GNDA 0.080087f
C590 bgr_0.TAIL_CUR_MIR_BIAS.t14 GNDA 0.093474f
C591 bgr_0.TAIL_CUR_MIR_BIAS.n8 GNDA 0.088131f
C592 bgr_0.TAIL_CUR_MIR_BIAS.n9 GNDA 0.055271f
C593 bgr_0.TAIL_CUR_MIR_BIAS.n10 GNDA 0.055271f
C594 bgr_0.TAIL_CUR_MIR_BIAS.n11 GNDA 0.055271f
C595 bgr_0.TAIL_CUR_MIR_BIAS.n12 GNDA 0.055271f
C596 bgr_0.TAIL_CUR_MIR_BIAS.n13 GNDA 0.055271f
C597 bgr_0.TAIL_CUR_MIR_BIAS.n14 GNDA 0.055271f
C598 bgr_0.TAIL_CUR_MIR_BIAS.n15 GNDA 0.055271f
C599 bgr_0.TAIL_CUR_MIR_BIAS.n16 GNDA 0.04939f
C600 bgr_0.TAIL_CUR_MIR_BIAS.t19 GNDA 0.080087f
C601 bgr_0.TAIL_CUR_MIR_BIAS.t29 GNDA 0.080087f
C602 bgr_0.TAIL_CUR_MIR_BIAS.t23 GNDA 0.080087f
C603 bgr_0.TAIL_CUR_MIR_BIAS.t15 GNDA 0.080087f
C604 bgr_0.TAIL_CUR_MIR_BIAS.t25 GNDA 0.080087f
C605 bgr_0.TAIL_CUR_MIR_BIAS.t17 GNDA 0.080087f
C606 bgr_0.TAIL_CUR_MIR_BIAS.t27 GNDA 0.080087f
C607 bgr_0.TAIL_CUR_MIR_BIAS.t21 GNDA 0.080087f
C608 bgr_0.TAIL_CUR_MIR_BIAS.t30 GNDA 0.080087f
C609 bgr_0.TAIL_CUR_MIR_BIAS.t12 GNDA 0.093474f
C610 bgr_0.TAIL_CUR_MIR_BIAS.n17 GNDA 0.088131f
C611 bgr_0.TAIL_CUR_MIR_BIAS.n18 GNDA 0.055271f
C612 bgr_0.TAIL_CUR_MIR_BIAS.n19 GNDA 0.055271f
C613 bgr_0.TAIL_CUR_MIR_BIAS.n20 GNDA 0.055271f
C614 bgr_0.TAIL_CUR_MIR_BIAS.n21 GNDA 0.055271f
C615 bgr_0.TAIL_CUR_MIR_BIAS.n22 GNDA 0.055271f
C616 bgr_0.TAIL_CUR_MIR_BIAS.n23 GNDA 0.055271f
C617 bgr_0.TAIL_CUR_MIR_BIAS.n24 GNDA 0.055271f
C618 bgr_0.TAIL_CUR_MIR_BIAS.n25 GNDA 0.04939f
C619 bgr_0.TAIL_CUR_MIR_BIAS.n26 GNDA 0.12343f
C620 bgr_0.TAIL_CUR_MIR_BIAS.t3 GNDA 0.045119f
C621 bgr_0.TAIL_CUR_MIR_BIAS.t1 GNDA 0.045119f
C622 bgr_0.TAIL_CUR_MIR_BIAS.n27 GNDA 0.090239f
C623 bgr_0.TAIL_CUR_MIR_BIAS.n28 GNDA 0.349784f
C624 bgr_0.TAIL_CUR_MIR_BIAS.n29 GNDA 3.57484f
C625 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.344645f
C626 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.345894f
C627 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.344645f
C628 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.347347f
C629 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.37779f
C630 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.344645f
C631 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.345894f
C632 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.344645f
C633 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.345894f
C634 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.344645f
C635 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.345894f
C636 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.344645f
C637 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.345894f
C638 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.344645f
C639 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.345894f
C640 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.344645f
C641 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.345894f
C642 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.344645f
C643 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.345894f
C644 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.344645f
C645 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.345894f
C646 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.344645f
C647 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.345894f
C648 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.344645f
C649 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.345894f
C650 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.344645f
C651 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.345894f
C652 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.344645f
C653 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.345894f
C654 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.344645f
C655 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.345894f
C656 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.344645f
C657 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.345894f
C658 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.344645f
C659 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.345894f
C660 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.344645f
C661 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.345894f
C662 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.344645f
C663 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.345894f
C664 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.344645f
C665 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.345894f
C666 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.344645f
C667 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.345894f
C668 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.344645f
C669 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.345894f
C670 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.344645f
C671 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.345894f
C672 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.344645f
C673 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.345894f
C674 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.344645f
C675 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.345894f
C676 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.344645f
C677 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.345894f
C678 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.344645f
C679 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.345894f
C680 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.344645f
C681 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.345894f
C682 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.344645f
C683 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.345894f
C684 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.344645f
C685 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.345894f
C686 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.344645f
C687 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.345894f
C688 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.344645f
C689 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.361543f
C690 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.344645f
C691 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.185116f
C692 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.19812f
C693 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.344645f
C694 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.185116f
C695 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.196522f
C696 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.344645f
C697 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.185116f
C698 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.196522f
C699 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.344645f
C700 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.185116f
C701 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.196522f
C702 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.344645f
C703 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.185116f
C704 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.196522f
C705 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.344645f
C706 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.185116f
C707 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.196522f
C708 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.344645f
C709 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.185116f
C710 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.196522f
C711 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.344645f
C712 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.185116f
C713 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196522f
C714 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.344645f
C715 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.185116f
C716 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196522f
C717 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.344645f
C718 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.345894f
C719 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.166619f
C720 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.214914f
C721 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.18397f
C722 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.23341f
C723 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.18397f
C724 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.250658f
C725 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.18397f
C726 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.250658f
C727 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.18397f
C728 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.250658f
C729 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.18397f
C730 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.250658f
C731 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.18397f
C732 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.250658f
C733 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.18397f
C734 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.250658f
C735 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.18397f
C736 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250658f
C737 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.18397f
C738 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250658f
C739 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.18397f
C740 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250658f
C741 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.18397f
C742 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250658f
C743 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.18397f
C744 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250658f
C745 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.18397f
C746 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250658f
C747 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.18397f
C748 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250658f
C749 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.18397f
C750 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250658f
C751 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.18397f
C752 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.23341f
C753 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.343499f
C754 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.166619f
C755 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.216163f
C756 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.343499f
C757 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.166619f
C758 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.216163f
C759 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.343499f
C760 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.344645f
C761 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.363141f
C762 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.363141f
C763 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.185116f
C764 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.216163f
C765 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.343499f
C766 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.344645f
C767 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.185116f
C768 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.197667f
C769 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.343499f
C770 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.344645f
C771 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.185116f
C772 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.216163f
C773 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.343499f
C774 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.344645f
C775 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.185116f
C776 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.216163f
C777 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.343499f
C778 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.344645f
C779 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.185116f
C780 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216163f
C781 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.343499f
C782 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.344645f
C783 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.363141f
C784 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.363141f
C785 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.185116f
C786 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216163f
C787 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.343499f
C788 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.344645f
C789 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.363141f
C790 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.363141f
C791 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.185116f
C792 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216163f
C793 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.343499f
C794 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216163f
C795 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.185116f
C796 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.363141f
C797 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.363141f
C798 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.764814f
C799 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.3034f
C800 bgr_0.V_mir1.t8 GNDA 0.053881f
C801 bgr_0.V_mir1.t6 GNDA 0.042444f
C802 bgr_0.V_mir1.t17 GNDA 0.042444f
C803 bgr_0.V_mir1.t20 GNDA 0.06851f
C804 bgr_0.V_mir1.n0 GNDA 0.076506f
C805 bgr_0.V_mir1.n1 GNDA 0.052264f
C806 bgr_0.V_mir1.n2 GNDA 0.081315f
C807 bgr_0.V_mir1.t9 GNDA 0.03537f
C808 bgr_0.V_mir1.t7 GNDA 0.03537f
C809 bgr_0.V_mir1.n3 GNDA 0.08097f
C810 bgr_0.V_mir1.n4 GNDA 0.203577f
C811 bgr_0.V_mir1.t12 GNDA 0.017685f
C812 bgr_0.V_mir1.t15 GNDA 0.017685f
C813 bgr_0.V_mir1.n5 GNDA 0.046242f
C814 bgr_0.V_mir1.t14 GNDA 0.075466f
C815 bgr_0.V_mir1.t13 GNDA 0.017685f
C816 bgr_0.V_mir1.t16 GNDA 0.017685f
C817 bgr_0.V_mir1.n6 GNDA 0.050199f
C818 bgr_0.V_mir1.n7 GNDA 0.827814f
C819 bgr_0.V_mir1.n8 GNDA 0.268286f
C820 bgr_0.V_mir1.t0 GNDA 0.053881f
C821 bgr_0.V_mir1.t4 GNDA 0.042444f
C822 bgr_0.V_mir1.t18 GNDA 0.042444f
C823 bgr_0.V_mir1.t21 GNDA 0.06851f
C824 bgr_0.V_mir1.n9 GNDA 0.076506f
C825 bgr_0.V_mir1.n10 GNDA 0.052264f
C826 bgr_0.V_mir1.n11 GNDA 0.081315f
C827 bgr_0.V_mir1.t1 GNDA 0.03537f
C828 bgr_0.V_mir1.t5 GNDA 0.03537f
C829 bgr_0.V_mir1.n12 GNDA 0.08097f
C830 bgr_0.V_mir1.n13 GNDA 0.156007f
C831 bgr_0.V_mir1.n14 GNDA 0.09373f
C832 bgr_0.V_mir1.n15 GNDA 0.699157f
C833 bgr_0.V_mir1.t10 GNDA 0.053881f
C834 bgr_0.V_mir1.t2 GNDA 0.042444f
C835 bgr_0.V_mir1.t19 GNDA 0.042444f
C836 bgr_0.V_mir1.t22 GNDA 0.06851f
C837 bgr_0.V_mir1.n16 GNDA 0.076506f
C838 bgr_0.V_mir1.n17 GNDA 0.052264f
C839 bgr_0.V_mir1.n18 GNDA 0.081315f
C840 bgr_0.V_mir1.n19 GNDA 0.201563f
C841 bgr_0.V_mir1.t3 GNDA 0.03537f
C842 bgr_0.V_mir1.n20 GNDA 0.08097f
C843 bgr_0.V_mir1.t11 GNDA 0.03537f
C844 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.477162f
C845 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.115051f
C846 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.115051f
C847 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.47578f
C848 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.115051f
C849 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.115051f
C850 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.473954f
C851 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.657138f
C852 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.115051f
C853 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.115051f
C854 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.473954f
C855 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.342904f
C856 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.115051f
C857 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.115051f
C858 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.473954f
C859 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.342904f
C860 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.115051f
C861 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.115051f
C862 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.473954f
C863 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.49568f
C864 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 7.289f
C865 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.03835f
C866 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.03835f
C867 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.139392f
C868 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.03835f
C869 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.03835f
C870 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.115834f
C871 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.724132f
C872 bgr_0.V_CMFB_S4 GNDA 5.94035f
C873 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.033671f
C874 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.033671f
C875 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.084438f
C876 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.033671f
C877 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.033671f
C878 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.083993f
C879 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.568968f
C880 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.033671f
C881 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.033671f
C882 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.083993f
C883 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.597848f
C884 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.430908f
C885 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.067342f
C886 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.067342f
C887 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.19758f
C888 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.067342f
C889 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.067342f
C890 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.196683f
C891 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.679849f
C892 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.067342f
C893 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.067342f
C894 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.196683f
C895 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.352158f
C896 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.067342f
C897 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.067342f
C898 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.196683f
C899 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.352158f
C900 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.067342f
C901 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.067342f
C902 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.196683f
C903 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.508351f
C904 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 5.05557f
C905 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 GNDA 4.02733f
C906 bgr_0.V_CMFB_S3 GNDA 0.014671f
C907 bgr_0.PFET_GATE_10uA.t23 GNDA 0.039179f
C908 bgr_0.PFET_GATE_10uA.t16 GNDA 0.057916f
C909 bgr_0.PFET_GATE_10uA.n0 GNDA 0.063817f
C910 bgr_0.PFET_GATE_10uA.t29 GNDA 0.039179f
C911 bgr_0.PFET_GATE_10uA.t17 GNDA 0.057916f
C912 bgr_0.PFET_GATE_10uA.n1 GNDA 0.063817f
C913 bgr_0.PFET_GATE_10uA.n2 GNDA 0.076791f
C914 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039179f
C915 bgr_0.PFET_GATE_10uA.t24 GNDA 0.057916f
C916 bgr_0.PFET_GATE_10uA.n3 GNDA 0.063817f
C917 bgr_0.PFET_GATE_10uA.t18 GNDA 0.039179f
C918 bgr_0.PFET_GATE_10uA.t25 GNDA 0.057916f
C919 bgr_0.PFET_GATE_10uA.n4 GNDA 0.063817f
C920 bgr_0.PFET_GATE_10uA.n5 GNDA 0.064022f
C921 bgr_0.PFET_GATE_10uA.t2 GNDA 0.781422f
C922 bgr_0.PFET_GATE_10uA.t4 GNDA 0.586977f
C923 bgr_0.PFET_GATE_10uA.t0 GNDA 0.040183f
C924 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040183f
C925 bgr_0.PFET_GATE_10uA.n6 GNDA 0.102705f
C926 bgr_0.PFET_GATE_10uA.t1 GNDA 0.040183f
C927 bgr_0.PFET_GATE_10uA.t9 GNDA 0.040183f
C928 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100051f
C929 bgr_0.PFET_GATE_10uA.n8 GNDA 0.978629f
C930 bgr_0.PFET_GATE_10uA.t7 GNDA 0.040183f
C931 bgr_0.PFET_GATE_10uA.t8 GNDA 0.040183f
C932 bgr_0.PFET_GATE_10uA.n9 GNDA 0.100051f
C933 bgr_0.PFET_GATE_10uA.n10 GNDA 0.554934f
C934 bgr_0.PFET_GATE_10uA.n11 GNDA 1.13286f
C935 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040183f
C936 bgr_0.PFET_GATE_10uA.t3 GNDA 0.040183f
C937 bgr_0.PFET_GATE_10uA.n12 GNDA 0.096913f
C938 bgr_0.PFET_GATE_10uA.n13 GNDA 0.356682f
C939 bgr_0.PFET_GATE_10uA.n14 GNDA 3.84996f
C940 bgr_0.PFET_GATE_10uA.t13 GNDA 0.045299f
C941 bgr_0.PFET_GATE_10uA.t21 GNDA 0.045299f
C942 bgr_0.PFET_GATE_10uA.n15 GNDA 0.137138f
C943 bgr_0.PFET_GATE_10uA.n16 GNDA 1.78858f
C944 bgr_0.PFET_GATE_10uA.n17 GNDA 1.41725f
C945 bgr_0.PFET_GATE_10uA.t27 GNDA 0.039179f
C946 bgr_0.PFET_GATE_10uA.t20 GNDA 0.039179f
C947 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039179f
C948 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039179f
C949 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039179f
C950 bgr_0.PFET_GATE_10uA.t11 GNDA 0.057916f
C951 bgr_0.PFET_GATE_10uA.n18 GNDA 0.071675f
C952 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051234f
C953 bgr_0.PFET_GATE_10uA.n20 GNDA 0.051234f
C954 bgr_0.PFET_GATE_10uA.n21 GNDA 0.051234f
C955 bgr_0.PFET_GATE_10uA.n22 GNDA 0.043376f
C956 bgr_0.PFET_GATE_10uA.t14 GNDA 0.039179f
C957 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039179f
C958 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039179f
C959 bgr_0.PFET_GATE_10uA.t15 GNDA 0.057916f
C960 bgr_0.PFET_GATE_10uA.n23 GNDA 0.071675f
C961 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051234f
C962 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043376f
C963 bgr_0.PFET_GATE_10uA.n26 GNDA 0.05954f
C964 two_stage_opamp_dummy_magic_0.VOUT+.t16 GNDA 0.043632f
C965 two_stage_opamp_dummy_magic_0.VOUT+.t10 GNDA 0.043632f
C966 two_stage_opamp_dummy_magic_0.VOUT+.n0 GNDA 0.175369f
C967 two_stage_opamp_dummy_magic_0.VOUT+.t5 GNDA 0.043632f
C968 two_stage_opamp_dummy_magic_0.VOUT+.t9 GNDA 0.043632f
C969 two_stage_opamp_dummy_magic_0.VOUT+.n1 GNDA 0.175046f
C970 two_stage_opamp_dummy_magic_0.VOUT+.n2 GNDA 0.17244f
C971 two_stage_opamp_dummy_magic_0.VOUT+.t4 GNDA 0.043632f
C972 two_stage_opamp_dummy_magic_0.VOUT+.t8 GNDA 0.043632f
C973 two_stage_opamp_dummy_magic_0.VOUT+.n3 GNDA 0.175046f
C974 two_stage_opamp_dummy_magic_0.VOUT+.n4 GNDA 0.088927f
C975 two_stage_opamp_dummy_magic_0.VOUT+.t12 GNDA 0.043632f
C976 two_stage_opamp_dummy_magic_0.VOUT+.t6 GNDA 0.043632f
C977 two_stage_opamp_dummy_magic_0.VOUT+.n5 GNDA 0.175046f
C978 two_stage_opamp_dummy_magic_0.VOUT+.n6 GNDA 0.088927f
C979 two_stage_opamp_dummy_magic_0.VOUT+.t11 GNDA 0.043632f
C980 two_stage_opamp_dummy_magic_0.VOUT+.t17 GNDA 0.043632f
C981 two_stage_opamp_dummy_magic_0.VOUT+.n7 GNDA 0.175368f
C982 two_stage_opamp_dummy_magic_0.VOUT+.n8 GNDA 0.10533f
C983 two_stage_opamp_dummy_magic_0.VOUT+.t13 GNDA 0.043632f
C984 two_stage_opamp_dummy_magic_0.VOUT+.t7 GNDA 0.043632f
C985 two_stage_opamp_dummy_magic_0.VOUT+.n9 GNDA 0.172903f
C986 two_stage_opamp_dummy_magic_0.VOUT+.n10 GNDA 0.212302f
C987 two_stage_opamp_dummy_magic_0.VOUT+.t117 GNDA 0.295834f
C988 two_stage_opamp_dummy_magic_0.VOUT+.t25 GNDA 0.290879f
C989 two_stage_opamp_dummy_magic_0.VOUT+.n11 GNDA 0.195025f
C990 two_stage_opamp_dummy_magic_0.VOUT+.t124 GNDA 0.290879f
C991 two_stage_opamp_dummy_magic_0.VOUT+.n12 GNDA 0.12726f
C992 two_stage_opamp_dummy_magic_0.VOUT+.t72 GNDA 0.295834f
C993 two_stage_opamp_dummy_magic_0.VOUT+.t38 GNDA 0.290879f
C994 two_stage_opamp_dummy_magic_0.VOUT+.n13 GNDA 0.195025f
C995 two_stage_opamp_dummy_magic_0.VOUT+.t127 GNDA 0.290879f
C996 two_stage_opamp_dummy_magic_0.VOUT+.t34 GNDA 0.295213f
C997 two_stage_opamp_dummy_magic_0.VOUT+.t86 GNDA 0.295213f
C998 two_stage_opamp_dummy_magic_0.VOUT+.t42 GNDA 0.295213f
C999 two_stage_opamp_dummy_magic_0.VOUT+.t96 GNDA 0.295213f
C1000 two_stage_opamp_dummy_magic_0.VOUT+.t143 GNDA 0.295213f
C1001 two_stage_opamp_dummy_magic_0.VOUT+.t106 GNDA 0.295213f
C1002 two_stage_opamp_dummy_magic_0.VOUT+.t154 GNDA 0.295213f
C1003 two_stage_opamp_dummy_magic_0.VOUT+.t64 GNDA 0.295213f
C1004 two_stage_opamp_dummy_magic_0.VOUT+.t116 GNDA 0.295213f
C1005 two_stage_opamp_dummy_magic_0.VOUT+.t73 GNDA 0.295213f
C1006 two_stage_opamp_dummy_magic_0.VOUT+.t149 GNDA 0.290879f
C1007 two_stage_opamp_dummy_magic_0.VOUT+.n14 GNDA 0.195645f
C1008 two_stage_opamp_dummy_magic_0.VOUT+.t58 GNDA 0.290879f
C1009 two_stage_opamp_dummy_magic_0.VOUT+.n15 GNDA 0.250185f
C1010 two_stage_opamp_dummy_magic_0.VOUT+.t97 GNDA 0.290879f
C1011 two_stage_opamp_dummy_magic_0.VOUT+.n16 GNDA 0.250185f
C1012 two_stage_opamp_dummy_magic_0.VOUT+.t131 GNDA 0.290879f
C1013 two_stage_opamp_dummy_magic_0.VOUT+.n17 GNDA 0.250185f
C1014 two_stage_opamp_dummy_magic_0.VOUT+.t24 GNDA 0.290879f
C1015 two_stage_opamp_dummy_magic_0.VOUT+.n18 GNDA 0.250185f
C1016 two_stage_opamp_dummy_magic_0.VOUT+.t75 GNDA 0.290879f
C1017 two_stage_opamp_dummy_magic_0.VOUT+.n19 GNDA 0.250185f
C1018 two_stage_opamp_dummy_magic_0.VOUT+.t113 GNDA 0.290879f
C1019 two_stage_opamp_dummy_magic_0.VOUT+.n20 GNDA 0.250185f
C1020 two_stage_opamp_dummy_magic_0.VOUT+.t144 GNDA 0.290879f
C1021 two_stage_opamp_dummy_magic_0.VOUT+.n21 GNDA 0.250185f
C1022 two_stage_opamp_dummy_magic_0.VOUT+.t54 GNDA 0.290879f
C1023 two_stage_opamp_dummy_magic_0.VOUT+.n22 GNDA 0.250185f
C1024 two_stage_opamp_dummy_magic_0.VOUT+.t94 GNDA 0.290879f
C1025 two_stage_opamp_dummy_magic_0.VOUT+.n23 GNDA 0.250185f
C1026 two_stage_opamp_dummy_magic_0.VOUT+.n24 GNDA 0.236339f
C1027 two_stage_opamp_dummy_magic_0.VOUT+.t37 GNDA 0.295834f
C1028 two_stage_opamp_dummy_magic_0.VOUT+.t142 GNDA 0.290879f
C1029 two_stage_opamp_dummy_magic_0.VOUT+.n25 GNDA 0.195025f
C1030 two_stage_opamp_dummy_magic_0.VOUT+.t93 GNDA 0.290879f
C1031 two_stage_opamp_dummy_magic_0.VOUT+.t20 GNDA 0.295834f
C1032 two_stage_opamp_dummy_magic_0.VOUT+.t57 GNDA 0.290879f
C1033 two_stage_opamp_dummy_magic_0.VOUT+.n26 GNDA 0.195025f
C1034 two_stage_opamp_dummy_magic_0.VOUT+.n27 GNDA 0.236339f
C1035 two_stage_opamp_dummy_magic_0.VOUT+.t79 GNDA 0.295834f
C1036 two_stage_opamp_dummy_magic_0.VOUT+.t41 GNDA 0.290879f
C1037 two_stage_opamp_dummy_magic_0.VOUT+.n28 GNDA 0.195025f
C1038 two_stage_opamp_dummy_magic_0.VOUT+.t133 GNDA 0.290879f
C1039 two_stage_opamp_dummy_magic_0.VOUT+.t60 GNDA 0.295834f
C1040 two_stage_opamp_dummy_magic_0.VOUT+.t100 GNDA 0.290879f
C1041 two_stage_opamp_dummy_magic_0.VOUT+.n29 GNDA 0.195025f
C1042 two_stage_opamp_dummy_magic_0.VOUT+.n30 GNDA 0.236339f
C1043 two_stage_opamp_dummy_magic_0.VOUT+.t121 GNDA 0.295834f
C1044 two_stage_opamp_dummy_magic_0.VOUT+.t83 GNDA 0.290879f
C1045 two_stage_opamp_dummy_magic_0.VOUT+.n31 GNDA 0.195025f
C1046 two_stage_opamp_dummy_magic_0.VOUT+.t31 GNDA 0.290879f
C1047 two_stage_opamp_dummy_magic_0.VOUT+.t104 GNDA 0.295834f
C1048 two_stage_opamp_dummy_magic_0.VOUT+.t137 GNDA 0.290879f
C1049 two_stage_opamp_dummy_magic_0.VOUT+.n32 GNDA 0.195025f
C1050 two_stage_opamp_dummy_magic_0.VOUT+.n33 GNDA 0.236339f
C1051 two_stage_opamp_dummy_magic_0.VOUT+.t84 GNDA 0.295834f
C1052 two_stage_opamp_dummy_magic_0.VOUT+.t49 GNDA 0.290879f
C1053 two_stage_opamp_dummy_magic_0.VOUT+.n34 GNDA 0.195025f
C1054 two_stage_opamp_dummy_magic_0.VOUT+.t138 GNDA 0.290879f
C1055 two_stage_opamp_dummy_magic_0.VOUT+.t66 GNDA 0.295834f
C1056 two_stage_opamp_dummy_magic_0.VOUT+.t103 GNDA 0.290879f
C1057 two_stage_opamp_dummy_magic_0.VOUT+.n35 GNDA 0.195025f
C1058 two_stage_opamp_dummy_magic_0.VOUT+.n36 GNDA 0.236339f
C1059 two_stage_opamp_dummy_magic_0.VOUT+.t108 GNDA 0.295834f
C1060 two_stage_opamp_dummy_magic_0.VOUT+.t69 GNDA 0.290879f
C1061 two_stage_opamp_dummy_magic_0.VOUT+.n37 GNDA 0.195025f
C1062 two_stage_opamp_dummy_magic_0.VOUT+.t90 GNDA 0.290879f
C1063 two_stage_opamp_dummy_magic_0.VOUT+.n38 GNDA 0.12726f
C1064 two_stage_opamp_dummy_magic_0.VOUT+.t67 GNDA 0.295834f
C1065 two_stage_opamp_dummy_magic_0.VOUT+.t30 GNDA 0.290879f
C1066 two_stage_opamp_dummy_magic_0.VOUT+.n39 GNDA 0.195025f
C1067 two_stage_opamp_dummy_magic_0.VOUT+.t51 GNDA 0.290879f
C1068 two_stage_opamp_dummy_magic_0.VOUT+.t53 GNDA 0.295213f
C1069 two_stage_opamp_dummy_magic_0.VOUT+.t156 GNDA 0.295213f
C1070 two_stage_opamp_dummy_magic_0.VOUT+.t44 GNDA 0.295834f
C1071 two_stage_opamp_dummy_magic_0.VOUT+.t136 GNDA 0.290879f
C1072 two_stage_opamp_dummy_magic_0.VOUT+.n40 GNDA 0.195025f
C1073 two_stage_opamp_dummy_magic_0.VOUT+.t101 GNDA 0.290879f
C1074 two_stage_opamp_dummy_magic_0.VOUT+.n41 GNDA 0.122715f
C1075 two_stage_opamp_dummy_magic_0.VOUT+.t36 GNDA 0.295213f
C1076 two_stage_opamp_dummy_magic_0.VOUT+.t151 GNDA 0.295834f
C1077 two_stage_opamp_dummy_magic_0.VOUT+.t98 GNDA 0.290879f
C1078 two_stage_opamp_dummy_magic_0.VOUT+.n42 GNDA 0.195025f
C1079 two_stage_opamp_dummy_magic_0.VOUT+.t59 GNDA 0.290879f
C1080 two_stage_opamp_dummy_magic_0.VOUT+.n43 GNDA 0.122715f
C1081 two_stage_opamp_dummy_magic_0.VOUT+.t140 GNDA 0.295213f
C1082 two_stage_opamp_dummy_magic_0.VOUT+.t118 GNDA 0.295834f
C1083 two_stage_opamp_dummy_magic_0.VOUT+.t56 GNDA 0.290879f
C1084 two_stage_opamp_dummy_magic_0.VOUT+.n44 GNDA 0.195025f
C1085 two_stage_opamp_dummy_magic_0.VOUT+.t21 GNDA 0.290879f
C1086 two_stage_opamp_dummy_magic_0.VOUT+.n45 GNDA 0.122715f
C1087 two_stage_opamp_dummy_magic_0.VOUT+.t105 GNDA 0.295213f
C1088 two_stage_opamp_dummy_magic_0.VOUT+.t65 GNDA 0.295834f
C1089 two_stage_opamp_dummy_magic_0.VOUT+.t80 GNDA 0.290879f
C1090 two_stage_opamp_dummy_magic_0.VOUT+.n46 GNDA 0.195025f
C1091 two_stage_opamp_dummy_magic_0.VOUT+.t43 GNDA 0.290879f
C1092 two_stage_opamp_dummy_magic_0.VOUT+.n47 GNDA 0.122715f
C1093 two_stage_opamp_dummy_magic_0.VOUT+.t125 GNDA 0.295213f
C1094 two_stage_opamp_dummy_magic_0.VOUT+.t145 GNDA 0.295457f
C1095 two_stage_opamp_dummy_magic_0.VOUT+.t87 GNDA 0.295213f
C1096 two_stage_opamp_dummy_magic_0.VOUT+.t110 GNDA 0.295457f
C1097 two_stage_opamp_dummy_magic_0.VOUT+.t50 GNDA 0.295213f
C1098 two_stage_opamp_dummy_magic_0.VOUT+.t70 GNDA 0.295457f
C1099 two_stage_opamp_dummy_magic_0.VOUT+.t150 GNDA 0.295213f
C1100 two_stage_opamp_dummy_magic_0.VOUT+.t95 GNDA 0.295457f
C1101 two_stage_opamp_dummy_magic_0.VOUT+.t32 GNDA 0.295213f
C1102 two_stage_opamp_dummy_magic_0.VOUT+.t134 GNDA 0.290879f
C1103 two_stage_opamp_dummy_magic_0.VOUT+.n48 GNDA 0.321963f
C1104 two_stage_opamp_dummy_magic_0.VOUT+.t111 GNDA 0.290879f
C1105 two_stage_opamp_dummy_magic_0.VOUT+.n49 GNDA 0.376503f
C1106 two_stage_opamp_dummy_magic_0.VOUT+.t147 GNDA 0.290879f
C1107 two_stage_opamp_dummy_magic_0.VOUT+.n50 GNDA 0.376503f
C1108 two_stage_opamp_dummy_magic_0.VOUT+.t45 GNDA 0.290879f
C1109 two_stage_opamp_dummy_magic_0.VOUT+.n51 GNDA 0.376503f
C1110 two_stage_opamp_dummy_magic_0.VOUT+.t85 GNDA 0.290879f
C1111 two_stage_opamp_dummy_magic_0.VOUT+.n52 GNDA 0.30927f
C1112 two_stage_opamp_dummy_magic_0.VOUT+.t61 GNDA 0.290879f
C1113 two_stage_opamp_dummy_magic_0.VOUT+.n53 GNDA 0.30927f
C1114 two_stage_opamp_dummy_magic_0.VOUT+.t102 GNDA 0.290879f
C1115 two_stage_opamp_dummy_magic_0.VOUT+.n54 GNDA 0.30927f
C1116 two_stage_opamp_dummy_magic_0.VOUT+.t139 GNDA 0.290879f
C1117 two_stage_opamp_dummy_magic_0.VOUT+.n55 GNDA 0.30927f
C1118 two_stage_opamp_dummy_magic_0.VOUT+.t119 GNDA 0.290879f
C1119 two_stage_opamp_dummy_magic_0.VOUT+.n56 GNDA 0.250185f
C1120 two_stage_opamp_dummy_magic_0.VOUT+.t155 GNDA 0.290879f
C1121 two_stage_opamp_dummy_magic_0.VOUT+.n57 GNDA 0.250185f
C1122 two_stage_opamp_dummy_magic_0.VOUT+.n58 GNDA 0.236339f
C1123 two_stage_opamp_dummy_magic_0.VOUT+.t27 GNDA 0.295834f
C1124 two_stage_opamp_dummy_magic_0.VOUT+.t130 GNDA 0.290879f
C1125 two_stage_opamp_dummy_magic_0.VOUT+.n59 GNDA 0.195025f
C1126 two_stage_opamp_dummy_magic_0.VOUT+.t152 GNDA 0.290879f
C1127 two_stage_opamp_dummy_magic_0.VOUT+.t76 GNDA 0.295834f
C1128 two_stage_opamp_dummy_magic_0.VOUT+.t115 GNDA 0.290879f
C1129 two_stage_opamp_dummy_magic_0.VOUT+.n60 GNDA 0.195025f
C1130 two_stage_opamp_dummy_magic_0.VOUT+.n61 GNDA 0.236339f
C1131 two_stage_opamp_dummy_magic_0.VOUT+.t62 GNDA 0.295834f
C1132 two_stage_opamp_dummy_magic_0.VOUT+.t23 GNDA 0.290879f
C1133 two_stage_opamp_dummy_magic_0.VOUT+.n62 GNDA 0.195025f
C1134 two_stage_opamp_dummy_magic_0.VOUT+.t47 GNDA 0.290879f
C1135 two_stage_opamp_dummy_magic_0.VOUT+.t112 GNDA 0.295834f
C1136 two_stage_opamp_dummy_magic_0.VOUT+.t148 GNDA 0.290879f
C1137 two_stage_opamp_dummy_magic_0.VOUT+.n63 GNDA 0.195025f
C1138 two_stage_opamp_dummy_magic_0.VOUT+.n64 GNDA 0.236339f
C1139 two_stage_opamp_dummy_magic_0.VOUT+.t114 GNDA 0.295834f
C1140 two_stage_opamp_dummy_magic_0.VOUT+.t78 GNDA 0.290879f
C1141 two_stage_opamp_dummy_magic_0.VOUT+.n65 GNDA 0.195025f
C1142 two_stage_opamp_dummy_magic_0.VOUT+.t26 GNDA 0.290879f
C1143 two_stage_opamp_dummy_magic_0.VOUT+.t99 GNDA 0.295834f
C1144 two_stage_opamp_dummy_magic_0.VOUT+.t132 GNDA 0.290879f
C1145 two_stage_opamp_dummy_magic_0.VOUT+.n66 GNDA 0.195025f
C1146 two_stage_opamp_dummy_magic_0.VOUT+.n67 GNDA 0.236339f
C1147 two_stage_opamp_dummy_magic_0.VOUT+.t74 GNDA 0.295834f
C1148 two_stage_opamp_dummy_magic_0.VOUT+.t39 GNDA 0.290879f
C1149 two_stage_opamp_dummy_magic_0.VOUT+.n68 GNDA 0.195025f
C1150 two_stage_opamp_dummy_magic_0.VOUT+.t128 GNDA 0.290879f
C1151 two_stage_opamp_dummy_magic_0.VOUT+.t55 GNDA 0.295834f
C1152 two_stage_opamp_dummy_magic_0.VOUT+.t92 GNDA 0.290879f
C1153 two_stage_opamp_dummy_magic_0.VOUT+.n69 GNDA 0.195025f
C1154 two_stage_opamp_dummy_magic_0.VOUT+.n70 GNDA 0.236339f
C1155 two_stage_opamp_dummy_magic_0.VOUT+.t109 GNDA 0.295834f
C1156 two_stage_opamp_dummy_magic_0.VOUT+.t71 GNDA 0.290879f
C1157 two_stage_opamp_dummy_magic_0.VOUT+.n71 GNDA 0.195025f
C1158 two_stage_opamp_dummy_magic_0.VOUT+.t19 GNDA 0.290879f
C1159 two_stage_opamp_dummy_magic_0.VOUT+.t91 GNDA 0.295834f
C1160 two_stage_opamp_dummy_magic_0.VOUT+.t126 GNDA 0.290879f
C1161 two_stage_opamp_dummy_magic_0.VOUT+.n72 GNDA 0.195025f
C1162 two_stage_opamp_dummy_magic_0.VOUT+.n73 GNDA 0.236339f
C1163 two_stage_opamp_dummy_magic_0.VOUT+.t68 GNDA 0.295834f
C1164 two_stage_opamp_dummy_magic_0.VOUT+.t33 GNDA 0.290879f
C1165 two_stage_opamp_dummy_magic_0.VOUT+.n74 GNDA 0.195025f
C1166 two_stage_opamp_dummy_magic_0.VOUT+.t122 GNDA 0.290879f
C1167 two_stage_opamp_dummy_magic_0.VOUT+.t52 GNDA 0.295834f
C1168 two_stage_opamp_dummy_magic_0.VOUT+.t88 GNDA 0.290879f
C1169 two_stage_opamp_dummy_magic_0.VOUT+.n75 GNDA 0.195025f
C1170 two_stage_opamp_dummy_magic_0.VOUT+.n76 GNDA 0.236339f
C1171 two_stage_opamp_dummy_magic_0.VOUT+.t29 GNDA 0.295834f
C1172 two_stage_opamp_dummy_magic_0.VOUT+.t135 GNDA 0.290879f
C1173 two_stage_opamp_dummy_magic_0.VOUT+.n77 GNDA 0.195025f
C1174 two_stage_opamp_dummy_magic_0.VOUT+.t82 GNDA 0.290879f
C1175 two_stage_opamp_dummy_magic_0.VOUT+.t153 GNDA 0.295834f
C1176 two_stage_opamp_dummy_magic_0.VOUT+.t48 GNDA 0.290879f
C1177 two_stage_opamp_dummy_magic_0.VOUT+.n78 GNDA 0.195025f
C1178 two_stage_opamp_dummy_magic_0.VOUT+.n79 GNDA 0.236339f
C1179 two_stage_opamp_dummy_magic_0.VOUT+.t63 GNDA 0.295834f
C1180 two_stage_opamp_dummy_magic_0.VOUT+.t28 GNDA 0.290879f
C1181 two_stage_opamp_dummy_magic_0.VOUT+.n80 GNDA 0.195025f
C1182 two_stage_opamp_dummy_magic_0.VOUT+.t120 GNDA 0.290879f
C1183 two_stage_opamp_dummy_magic_0.VOUT+.t46 GNDA 0.295834f
C1184 two_stage_opamp_dummy_magic_0.VOUT+.t81 GNDA 0.290879f
C1185 two_stage_opamp_dummy_magic_0.VOUT+.n81 GNDA 0.195025f
C1186 two_stage_opamp_dummy_magic_0.VOUT+.n82 GNDA 0.236339f
C1187 two_stage_opamp_dummy_magic_0.VOUT+.t22 GNDA 0.295834f
C1188 two_stage_opamp_dummy_magic_0.VOUT+.t129 GNDA 0.290879f
C1189 two_stage_opamp_dummy_magic_0.VOUT+.n83 GNDA 0.195025f
C1190 two_stage_opamp_dummy_magic_0.VOUT+.t77 GNDA 0.290879f
C1191 two_stage_opamp_dummy_magic_0.VOUT+.t146 GNDA 0.295834f
C1192 two_stage_opamp_dummy_magic_0.VOUT+.t40 GNDA 0.290879f
C1193 two_stage_opamp_dummy_magic_0.VOUT+.n84 GNDA 0.195025f
C1194 two_stage_opamp_dummy_magic_0.VOUT+.n85 GNDA 0.236339f
C1195 two_stage_opamp_dummy_magic_0.VOUT+.t123 GNDA 0.295834f
C1196 two_stage_opamp_dummy_magic_0.VOUT+.t89 GNDA 0.290879f
C1197 two_stage_opamp_dummy_magic_0.VOUT+.n86 GNDA 0.195025f
C1198 two_stage_opamp_dummy_magic_0.VOUT+.t35 GNDA 0.290879f
C1199 two_stage_opamp_dummy_magic_0.VOUT+.n87 GNDA 0.236339f
C1200 two_stage_opamp_dummy_magic_0.VOUT+.t141 GNDA 0.290879f
C1201 two_stage_opamp_dummy_magic_0.VOUT+.n88 GNDA 0.12726f
C1202 two_stage_opamp_dummy_magic_0.VOUT+.t107 GNDA 0.290879f
C1203 two_stage_opamp_dummy_magic_0.VOUT+.n89 GNDA 0.238316f
C1204 two_stage_opamp_dummy_magic_0.VOUT+.n90 GNDA 0.291354f
C1205 two_stage_opamp_dummy_magic_0.VOUT+.t18 GNDA 0.050904f
C1206 two_stage_opamp_dummy_magic_0.VOUT+.t1 GNDA 0.050904f
C1207 two_stage_opamp_dummy_magic_0.VOUT+.n91 GNDA 0.235484f
C1208 two_stage_opamp_dummy_magic_0.VOUT+.t0 GNDA 0.050904f
C1209 two_stage_opamp_dummy_magic_0.VOUT+.t14 GNDA 0.050904f
C1210 two_stage_opamp_dummy_magic_0.VOUT+.n92 GNDA 0.234695f
C1211 two_stage_opamp_dummy_magic_0.VOUT+.n93 GNDA 0.14503f
C1212 two_stage_opamp_dummy_magic_0.VOUT+.t2 GNDA 0.050904f
C1213 two_stage_opamp_dummy_magic_0.VOUT+.t15 GNDA 0.050904f
C1214 two_stage_opamp_dummy_magic_0.VOUT+.n94 GNDA 0.234695f
C1215 two_stage_opamp_dummy_magic_0.VOUT+.n95 GNDA 0.089271f
C1216 two_stage_opamp_dummy_magic_0.VOUT+.n96 GNDA 0.165389f
C1217 two_stage_opamp_dummy_magic_0.VOUT+.t3 GNDA 0.084162f
C1218 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.019819f
C1219 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.019819f
C1220 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.066913f
C1221 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.019819f
C1222 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.019819f
C1223 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.071516f
C1224 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.019819f
C1225 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.019819f
C1226 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.071516f
C1227 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.019819f
C1228 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.019819f
C1229 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.070891f
C1230 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.26322f
C1231 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.019819f
C1232 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.019819f
C1233 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.070891f
C1234 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.136547f
C1235 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.019819f
C1236 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.019819f
C1237 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.070891f
C1238 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.136547f
C1239 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.166311f
C1240 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.134435f
C1241 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.645498f
C1242 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.087203f
C1243 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.087203f
C1244 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.092877f
C1245 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.073601f
C1246 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.039346f
C1247 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.087203f
C1248 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.087203f
C1249 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.087203f
C1250 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.087203f
C1251 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.087203f
C1252 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.087203f
C1253 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.092877f
C1254 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.073601f
C1255 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.04162f
C1256 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.04162f
C1257 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.04162f
C1258 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.04162f
C1259 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.039346f
C1260 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.02132f
C1261 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.765352f
C1262 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.027747f
C1263 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.027747f
C1264 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.027747f
C1265 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.027747f
C1266 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.027747f
C1267 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.027747f
C1268 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.027747f
C1269 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.033692f
C1270 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.033692f
C1271 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.021801f
C1272 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.021801f
C1273 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.021801f
C1274 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.021801f
C1275 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.021801f
C1276 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.019527f
C1277 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.027747f
C1278 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.033692f
C1279 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.031419f
C1280 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.019205f
C1281 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.042611f
C1282 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.042611f
C1283 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.042611f
C1284 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.042611f
C1285 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.042611f
C1286 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.042611f
C1287 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.042611f
C1288 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.048441f
C1289 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.043717f
C1290 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.026756f
C1291 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.026756f
C1292 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.026756f
C1293 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.026756f
C1294 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.026756f
C1295 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.024482f
C1296 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.042611f
C1297 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.048441f
C1298 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.041443f
C1299 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.019165f
C1300 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.251975f
C1301 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.347762f
C1302 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.08699f
C1303 a_8420_8490.t8 GNDA 0.043655f
C1304 a_8420_8490.t11 GNDA 0.043655f
C1305 a_8420_8490.t5 GNDA 0.043655f
C1306 a_8420_8490.n0 GNDA 0.151823f
C1307 a_8420_8490.t7 GNDA 0.043655f
C1308 a_8420_8490.t9 GNDA 0.043655f
C1309 a_8420_8490.n1 GNDA 0.151285f
C1310 a_8420_8490.n2 GNDA 0.285611f
C1311 a_8420_8490.t1 GNDA 0.043655f
C1312 a_8420_8490.t3 GNDA 0.043655f
C1313 a_8420_8490.n3 GNDA 0.151285f
C1314 a_8420_8490.n4 GNDA 0.148064f
C1315 a_8420_8490.t4 GNDA 0.043655f
C1316 a_8420_8490.t6 GNDA 0.043655f
C1317 a_8420_8490.n5 GNDA 0.151285f
C1318 a_8420_8490.n6 GNDA 0.148064f
C1319 a_8420_8490.t2 GNDA 0.043655f
C1320 a_8420_8490.t0 GNDA 0.043655f
C1321 a_8420_8490.n7 GNDA 0.151823f
C1322 a_8420_8490.n8 GNDA 0.285612f
C1323 a_8420_8490.n9 GNDA 0.151285f
C1324 a_8420_8490.t10 GNDA 0.043655f
C1325 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.061318f
C1326 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.061318f
C1327 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.213251f
C1328 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.061318f
C1329 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.061318f
C1330 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.212496f
C1331 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.401172f
C1332 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.061318f
C1333 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.061318f
C1334 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.212496f
C1335 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.207971f
C1336 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.061318f
C1337 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.061318f
C1338 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.212496f
C1339 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.200964f
C1340 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.061318f
C1341 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.061318f
C1342 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.212496f
C1343 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.270572f
C1344 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.061318f
C1345 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.061318f
C1346 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.213251f
C1347 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.061318f
C1348 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.061318f
C1349 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.212496f
C1350 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.401172f
C1351 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.061318f
C1352 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.061318f
C1353 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.212496f
C1354 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.207971f
C1355 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.061318f
C1356 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.061318f
C1357 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.212496f
C1358 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.207971f
C1359 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.061318f
C1360 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.061318f
C1361 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.212496f
C1362 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.207971f
C1363 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.061318f
C1364 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.061318f
C1365 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.212496f
C1366 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.315219f
C1367 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.012583f
C1368 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.012583f
C1369 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.027269f
C1370 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.03908f
C1371 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.168132f
C1372 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.09887f
C1373 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.09887f
C1374 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.09887f
C1375 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.09887f
C1376 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.114095f
C1377 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.092633f
C1378 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.056925f
C1379 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.056925f
C1380 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.053303f
C1381 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.09887f
C1382 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.09887f
C1383 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.09887f
C1384 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.09887f
C1385 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.114095f
C1386 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.092633f
C1387 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.056925f
C1388 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.056925f
C1389 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.053303f
C1390 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.036003f
C1391 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.09887f
C1392 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.09887f
C1393 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.09887f
C1394 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.09887f
C1395 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.114095f
C1396 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.092633f
C1397 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.056925f
C1398 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.056925f
C1399 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.053303f
C1400 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.09887f
C1401 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.09887f
C1402 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.09887f
C1403 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.09887f
C1404 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.114095f
C1405 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.092633f
C1406 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.056925f
C1407 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.056925f
C1408 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.053303f
C1409 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.035316f
C1410 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.802639f
C1411 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.604613f
C1412 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.119293f
C1413 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 3.15867f
C1414 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.019974f
C1415 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.019974f
C1416 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.066969f
C1417 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.019974f
C1418 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.019974f
C1419 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.065132f
C1420 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.526032f
C1421 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.019974f
C1422 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.019974f
C1423 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.066969f
C1424 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.019974f
C1425 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.019974f
C1426 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.065132f
C1427 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.526032f
C1428 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.274372f
C1429 bgr_0.VB2_CUR_BIAS GNDA 3.05596f
C1430 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.7726f
C1431 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 8.91394f
C1432 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.024917f
C1433 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.024917f
C1434 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.058161f
C1435 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.024917f
C1436 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.024917f
C1437 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.057785f
C1438 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.024917f
C1439 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.024917f
C1440 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.057785f
C1441 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.020556f
C1442 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.020556f
C1443 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.020556f
C1444 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.020556f
C1445 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.020556f
C1446 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.020556f
C1447 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.020556f
C1448 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.020556f
C1449 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.020556f
C1450 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.020556f
C1451 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.020556f
C1452 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.020556f
C1453 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.020556f
C1454 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.020556f
C1455 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.020556f
C1456 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.020556f
C1457 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.044539f
C1458 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.069456f
C1459 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.054194f
C1460 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.054194f
C1461 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.054194f
C1462 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.054194f
C1463 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.054194f
C1464 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.054194f
C1465 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.054194f
C1466 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.054194f
C1467 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.054194f
C1468 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.054194f
C1469 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.054194f
C1470 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.054194f
C1471 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.054194f
C1472 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.054194f
C1473 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.046376f
C1474 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.020556f
C1475 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.020556f
C1476 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.044539f
C1477 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.069456f
C1478 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.046376f
C1479 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.075239f
C1480 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.024917f
C1481 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.024917f
C1482 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.049834f
C1483 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.148444f
C1484 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.024917f
C1485 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.024917f
C1486 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.057785f
C1487 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.024917f
C1488 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.024917f
C1489 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.057355f
C1490 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.049834f
C1491 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.049834f
C1492 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.153708f
C1493 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.074255f
C1494 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.027767f
C1495 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.087091f
C1496 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.027767f
C1497 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.071293f
C1498 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.027767f
C1499 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.071293f
C1500 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.027767f
C1501 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.109376f
C1502 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.709082f
C1503 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.090054f
C1504 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.090054f
C1505 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.301772f
C1506 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 3.40029f
C1507 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.090054f
C1508 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.090054f
C1509 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.301772f
C1510 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.814897f
C1511 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.090054f
C1512 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.090054f
C1513 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.301772f
C1514 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 1.16504f
C1515 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 1.01344f
C1516 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.043395f
C1517 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.013631f
C1518 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.025436f
C1519 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.060728f
C1520 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.379723f
C1521 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.013631f
C1522 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.025436f
C1523 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.060728f
C1524 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.350774f
C1525 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.042979f
C1526 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.341551f
C1527 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.013631f
C1528 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.025436f
C1529 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.060728f
C1530 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.212091f
C1531 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.013631f
C1532 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.025436f
C1533 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.060728f
C1534 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.269546f
C1535 bgr_0.V_mir2.t4 GNDA 0.042444f
C1536 bgr_0.V_mir2.t18 GNDA 0.042444f
C1537 bgr_0.V_mir2.t20 GNDA 0.06851f
C1538 bgr_0.V_mir2.n0 GNDA 0.076506f
C1539 bgr_0.V_mir2.n1 GNDA 0.052264f
C1540 bgr_0.V_mir2.t8 GNDA 0.053881f
C1541 bgr_0.V_mir2.n2 GNDA 0.081315f
C1542 bgr_0.V_mir2.t5 GNDA 0.03537f
C1543 bgr_0.V_mir2.t9 GNDA 0.03537f
C1544 bgr_0.V_mir2.n3 GNDA 0.08097f
C1545 bgr_0.V_mir2.n4 GNDA 0.201563f
C1546 bgr_0.V_mir2.t0 GNDA 0.017685f
C1547 bgr_0.V_mir2.t3 GNDA 0.017685f
C1548 bgr_0.V_mir2.n5 GNDA 0.046242f
C1549 bgr_0.V_mir2.t2 GNDA 0.075466f
C1550 bgr_0.V_mir2.t16 GNDA 0.017685f
C1551 bgr_0.V_mir2.t1 GNDA 0.017685f
C1552 bgr_0.V_mir2.n6 GNDA 0.050199f
C1553 bgr_0.V_mir2.n7 GNDA 0.827814f
C1554 bgr_0.V_mir2.n8 GNDA 0.268286f
C1555 bgr_0.V_mir2.t12 GNDA 0.042444f
C1556 bgr_0.V_mir2.t19 GNDA 0.042444f
C1557 bgr_0.V_mir2.t22 GNDA 0.06851f
C1558 bgr_0.V_mir2.n9 GNDA 0.076506f
C1559 bgr_0.V_mir2.n10 GNDA 0.052264f
C1560 bgr_0.V_mir2.t10 GNDA 0.053881f
C1561 bgr_0.V_mir2.n11 GNDA 0.081315f
C1562 bgr_0.V_mir2.t13 GNDA 0.03537f
C1563 bgr_0.V_mir2.t11 GNDA 0.03537f
C1564 bgr_0.V_mir2.n12 GNDA 0.08097f
C1565 bgr_0.V_mir2.n13 GNDA 0.156007f
C1566 bgr_0.V_mir2.n14 GNDA 0.09373f
C1567 bgr_0.V_mir2.n15 GNDA 0.699157f
C1568 bgr_0.V_mir2.t14 GNDA 0.042444f
C1569 bgr_0.V_mir2.t21 GNDA 0.042444f
C1570 bgr_0.V_mir2.t17 GNDA 0.06851f
C1571 bgr_0.V_mir2.n16 GNDA 0.076506f
C1572 bgr_0.V_mir2.n17 GNDA 0.052264f
C1573 bgr_0.V_mir2.t6 GNDA 0.053881f
C1574 bgr_0.V_mir2.n18 GNDA 0.081315f
C1575 bgr_0.V_mir2.n19 GNDA 0.203577f
C1576 bgr_0.V_mir2.t7 GNDA 0.03537f
C1577 bgr_0.V_mir2.n20 GNDA 0.08097f
C1578 bgr_0.V_mir2.t15 GNDA 0.03537f
C1579 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.03109f
C1580 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.03109f
C1581 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.077932f
C1582 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.03109f
C1583 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.03109f
C1584 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.077521f
C1585 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.689005f
C1586 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.03109f
C1587 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.03109f
C1588 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.06218f
C1589 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.347514f
C1590 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.398172f
C1591 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.06218f
C1592 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.06218f
C1593 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.182434f
C1594 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.06218f
C1595 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.06218f
C1596 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.181606f
C1597 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.627735f
C1598 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.06218f
C1599 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.06218f
C1600 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.181606f
C1601 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.325163f
C1602 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.06218f
C1603 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.06218f
C1604 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.181606f
C1605 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.325163f
C1606 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.06218f
C1607 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.06218f
C1608 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.181606f
C1609 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.467149f
C1610 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 3.26646f
C1611 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 3.56079f
C1612 bgr_0.V_CMFB_S1 GNDA 0.058021f
C1613 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.020126f
C1614 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.020126f
C1615 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.067951f
C1616 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.020126f
C1617 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.020126f
C1618 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.072625f
C1619 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.020126f
C1620 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.020126f
C1621 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.071991f
C1622 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.267304f
C1623 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.020126f
C1624 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.020126f
C1625 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.071991f
C1626 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.138665f
C1627 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.020126f
C1628 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.020126f
C1629 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.071991f
C1630 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.138665f
C1631 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.020126f
C1632 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.020126f
C1633 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.072625f
C1634 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.168892f
C1635 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.210979f
C1636 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.028177f
C1637 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.034215f
C1638 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.031906f
C1639 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.028177f
C1640 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.028177f
C1641 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.028177f
C1642 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.028177f
C1643 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.028177f
C1644 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.028177f
C1645 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.028177f
C1646 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.034215f
C1647 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.034215f
C1648 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.022139f
C1649 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.022139f
C1650 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.022139f
C1651 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.022139f
C1652 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.022139f
C1653 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.01983f
C1654 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.019503f
C1655 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.043272f
C1656 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.049193f
C1657 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.042086f
C1658 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.043272f
C1659 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.043272f
C1660 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.043272f
C1661 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.043272f
C1662 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.043272f
C1663 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.043272f
C1664 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.043272f
C1665 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.049193f
C1666 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.044395f
C1667 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.027171f
C1668 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.027171f
C1669 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.027171f
C1670 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.027171f
C1671 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.027171f
C1672 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.024862f
C1673 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.019462f
C1674 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.259144f
C1675 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.37183f
C1676 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.088556f
C1677 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.088556f
C1678 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.088556f
C1679 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.088556f
C1680 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.088556f
C1681 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.088556f
C1682 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.094318f
C1683 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.074743f
C1684 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.042265f
C1685 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.042265f
C1686 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.042265f
C1687 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.042265f
C1688 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.039957f
C1689 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.088556f
C1690 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.088556f
C1691 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.094318f
C1692 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.074743f
C1693 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.039957f
C1694 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.021651f
C1695 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.77991f
C1696 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.655511f
C1697 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.343499f
C1698 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.344645f
C1699 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.185116f
C1700 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.197667f
C1701 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.343499f
C1702 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.344645f
C1703 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.185116f
C1704 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.216163f
C1705 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.343499f
C1706 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.344645f
C1707 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.185116f
C1708 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.216163f
C1709 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.343499f
C1710 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.344645f
C1711 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.185116f
C1712 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.216163f
C1713 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.343499f
C1714 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C1715 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.363141f
C1716 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.363141f
C1717 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.185116f
C1718 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.216163f
C1719 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.343499f
C1720 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.344645f
C1721 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.363141f
C1722 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.363141f
C1723 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.185116f
C1724 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.216163f
C1725 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.344645f
C1726 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.345894f
C1727 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.344645f
C1728 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.347347f
C1729 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.377789f
C1730 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.344645f
C1731 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.345894f
C1732 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.344645f
C1733 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.345894f
C1734 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.344645f
C1735 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345894f
C1736 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.344645f
C1737 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.345894f
C1738 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.344645f
C1739 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.345894f
C1740 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.344645f
C1741 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.345894f
C1742 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.344645f
C1743 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.345894f
C1744 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.344645f
C1745 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.345894f
C1746 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.344645f
C1747 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345894f
C1748 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.344645f
C1749 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.345894f
C1750 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.344645f
C1751 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.345894f
C1752 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.344645f
C1753 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.345894f
C1754 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.344645f
C1755 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.345894f
C1756 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.344645f
C1757 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.345894f
C1758 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.344645f
C1759 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.345894f
C1760 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.344645f
C1761 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.345894f
C1762 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.344645f
C1763 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.345894f
C1764 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.344645f
C1765 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.345894f
C1766 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.344645f
C1767 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.345894f
C1768 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.344645f
C1769 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.345894f
C1770 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.344645f
C1771 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.345894f
C1772 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.344645f
C1773 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.345894f
C1774 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.344645f
C1775 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.345894f
C1776 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.344645f
C1777 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.345894f
C1778 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.344645f
C1779 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.345894f
C1780 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.344645f
C1781 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345894f
C1782 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.344645f
C1783 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.345894f
C1784 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.344645f
C1785 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.345894f
C1786 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.344645f
C1787 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.361543f
C1788 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.344645f
C1789 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.185116f
C1790 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.19812f
C1791 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.344645f
C1792 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.185116f
C1793 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.196521f
C1794 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.344645f
C1795 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.185116f
C1796 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.196521f
C1797 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.344645f
C1798 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.185116f
C1799 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.196521f
C1800 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.344645f
C1801 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.185116f
C1802 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.196521f
C1803 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.344645f
C1804 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.185116f
C1805 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.196521f
C1806 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.344645f
C1807 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.185116f
C1808 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.196521f
C1809 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.344645f
C1810 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.185116f
C1811 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.196521f
C1812 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.344645f
C1813 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.185116f
C1814 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.196521f
C1815 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.344645f
C1816 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.345894f
C1817 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.344645f
C1818 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.345894f
C1819 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.166619f
C1820 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.214914f
C1821 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.18397f
C1822 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.23341f
C1823 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.18397f
C1824 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.250658f
C1825 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.18397f
C1826 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.250658f
C1827 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.18397f
C1828 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.250658f
C1829 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.18397f
C1830 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.250658f
C1831 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.18397f
C1832 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.250658f
C1833 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.18397f
C1834 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.250658f
C1835 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.18397f
C1836 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.250658f
C1837 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.18397f
C1838 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.250658f
C1839 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.18397f
C1840 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.250658f
C1841 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.18397f
C1842 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.250658f
C1843 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.18397f
C1844 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.250658f
C1845 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.18397f
C1846 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.250658f
C1847 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.18397f
C1848 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.250658f
C1849 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.18397f
C1850 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.250658f
C1851 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.18397f
C1852 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.23341f
C1853 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.343499f
C1854 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.166619f
C1855 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216163f
C1856 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.343499f
C1857 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.166619f
C1858 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216163f
C1859 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.343499f
C1860 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.344645f
C1861 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.363141f
C1862 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.363141f
C1863 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.185116f
C1864 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216163f
C1865 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.343499f
C1866 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216163f
C1867 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185116f
C1868 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.363141f
C1869 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.363141f
C1870 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.434494f
C1871 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.297192f
C1872 two_stage_opamp_dummy_magic_0.VOUT-.t7 GNDA 0.050904f
C1873 two_stage_opamp_dummy_magic_0.VOUT-.t3 GNDA 0.050904f
C1874 two_stage_opamp_dummy_magic_0.VOUT-.n0 GNDA 0.235484f
C1875 two_stage_opamp_dummy_magic_0.VOUT-.t5 GNDA 0.050904f
C1876 two_stage_opamp_dummy_magic_0.VOUT-.t16 GNDA 0.050904f
C1877 two_stage_opamp_dummy_magic_0.VOUT-.n1 GNDA 0.234695f
C1878 two_stage_opamp_dummy_magic_0.VOUT-.n2 GNDA 0.14503f
C1879 two_stage_opamp_dummy_magic_0.VOUT-.t14 GNDA 0.050904f
C1880 two_stage_opamp_dummy_magic_0.VOUT-.t8 GNDA 0.050904f
C1881 two_stage_opamp_dummy_magic_0.VOUT-.n3 GNDA 0.234695f
C1882 two_stage_opamp_dummy_magic_0.VOUT-.n4 GNDA 0.089271f
C1883 two_stage_opamp_dummy_magic_0.VOUT-.t17 GNDA 0.043632f
C1884 two_stage_opamp_dummy_magic_0.VOUT-.t0 GNDA 0.043632f
C1885 two_stage_opamp_dummy_magic_0.VOUT-.n5 GNDA 0.175369f
C1886 two_stage_opamp_dummy_magic_0.VOUT-.t13 GNDA 0.043632f
C1887 two_stage_opamp_dummy_magic_0.VOUT-.t18 GNDA 0.043632f
C1888 two_stage_opamp_dummy_magic_0.VOUT-.n6 GNDA 0.175368f
C1889 two_stage_opamp_dummy_magic_0.VOUT-.t10 GNDA 0.043632f
C1890 two_stage_opamp_dummy_magic_0.VOUT-.t4 GNDA 0.043632f
C1891 two_stage_opamp_dummy_magic_0.VOUT-.n7 GNDA 0.175046f
C1892 two_stage_opamp_dummy_magic_0.VOUT-.n8 GNDA 0.172441f
C1893 two_stage_opamp_dummy_magic_0.VOUT-.t2 GNDA 0.043632f
C1894 two_stage_opamp_dummy_magic_0.VOUT-.t15 GNDA 0.043632f
C1895 two_stage_opamp_dummy_magic_0.VOUT-.n9 GNDA 0.175046f
C1896 two_stage_opamp_dummy_magic_0.VOUT-.n10 GNDA 0.088927f
C1897 two_stage_opamp_dummy_magic_0.VOUT-.t1 GNDA 0.043632f
C1898 two_stage_opamp_dummy_magic_0.VOUT-.t12 GNDA 0.043632f
C1899 two_stage_opamp_dummy_magic_0.VOUT-.n11 GNDA 0.175046f
C1900 two_stage_opamp_dummy_magic_0.VOUT-.n12 GNDA 0.088927f
C1901 two_stage_opamp_dummy_magic_0.VOUT-.n13 GNDA 0.105329f
C1902 two_stage_opamp_dummy_magic_0.VOUT-.t9 GNDA 0.043632f
C1903 two_stage_opamp_dummy_magic_0.VOUT-.t11 GNDA 0.043632f
C1904 two_stage_opamp_dummy_magic_0.VOUT-.n14 GNDA 0.172903f
C1905 two_stage_opamp_dummy_magic_0.VOUT-.n15 GNDA 0.212301f
C1906 two_stage_opamp_dummy_magic_0.VOUT-.t101 GNDA 0.290879f
C1907 two_stage_opamp_dummy_magic_0.VOUT-.t108 GNDA 0.295834f
C1908 two_stage_opamp_dummy_magic_0.VOUT-.t149 GNDA 0.290879f
C1909 two_stage_opamp_dummy_magic_0.VOUT-.n16 GNDA 0.195025f
C1910 two_stage_opamp_dummy_magic_0.VOUT-.n17 GNDA 0.12726f
C1911 two_stage_opamp_dummy_magic_0.VOUT-.t48 GNDA 0.295213f
C1912 two_stage_opamp_dummy_magic_0.VOUT-.t92 GNDA 0.295213f
C1913 two_stage_opamp_dummy_magic_0.VOUT-.t42 GNDA 0.295213f
C1914 two_stage_opamp_dummy_magic_0.VOUT-.t130 GNDA 0.295213f
C1915 two_stage_opamp_dummy_magic_0.VOUT-.t84 GNDA 0.295213f
C1916 two_stage_opamp_dummy_magic_0.VOUT-.t125 GNDA 0.295213f
C1917 two_stage_opamp_dummy_magic_0.VOUT-.t74 GNDA 0.295213f
C1918 two_stage_opamp_dummy_magic_0.VOUT-.t23 GNDA 0.295213f
C1919 two_stage_opamp_dummy_magic_0.VOUT-.t64 GNDA 0.295213f
C1920 two_stage_opamp_dummy_magic_0.VOUT-.t150 GNDA 0.295213f
C1921 two_stage_opamp_dummy_magic_0.VOUT-.t88 GNDA 0.290879f
C1922 two_stage_opamp_dummy_magic_0.VOUT-.n18 GNDA 0.195645f
C1923 two_stage_opamp_dummy_magic_0.VOUT-.t51 GNDA 0.290879f
C1924 two_stage_opamp_dummy_magic_0.VOUT-.n19 GNDA 0.250185f
C1925 two_stage_opamp_dummy_magic_0.VOUT-.t137 GNDA 0.290879f
C1926 two_stage_opamp_dummy_magic_0.VOUT-.n20 GNDA 0.250185f
C1927 two_stage_opamp_dummy_magic_0.VOUT-.t106 GNDA 0.290879f
C1928 two_stage_opamp_dummy_magic_0.VOUT-.n21 GNDA 0.250185f
C1929 two_stage_opamp_dummy_magic_0.VOUT-.t75 GNDA 0.290879f
C1930 two_stage_opamp_dummy_magic_0.VOUT-.n22 GNDA 0.250185f
C1931 two_stage_opamp_dummy_magic_0.VOUT-.t25 GNDA 0.290879f
C1932 two_stage_opamp_dummy_magic_0.VOUT-.n23 GNDA 0.250185f
C1933 two_stage_opamp_dummy_magic_0.VOUT-.t128 GNDA 0.290879f
C1934 two_stage_opamp_dummy_magic_0.VOUT-.n24 GNDA 0.250185f
C1935 two_stage_opamp_dummy_magic_0.VOUT-.t90 GNDA 0.290879f
C1936 two_stage_opamp_dummy_magic_0.VOUT-.n25 GNDA 0.250185f
C1937 two_stage_opamp_dummy_magic_0.VOUT-.t54 GNDA 0.290879f
C1938 two_stage_opamp_dummy_magic_0.VOUT-.n26 GNDA 0.250185f
C1939 two_stage_opamp_dummy_magic_0.VOUT-.t140 GNDA 0.290879f
C1940 two_stage_opamp_dummy_magic_0.VOUT-.n27 GNDA 0.250185f
C1941 two_stage_opamp_dummy_magic_0.VOUT-.t110 GNDA 0.290879f
C1942 two_stage_opamp_dummy_magic_0.VOUT-.t28 GNDA 0.295834f
C1943 two_stage_opamp_dummy_magic_0.VOUT-.t79 GNDA 0.290879f
C1944 two_stage_opamp_dummy_magic_0.VOUT-.n28 GNDA 0.195025f
C1945 two_stage_opamp_dummy_magic_0.VOUT-.n29 GNDA 0.236339f
C1946 two_stage_opamp_dummy_magic_0.VOUT-.t24 GNDA 0.295834f
C1947 two_stage_opamp_dummy_magic_0.VOUT-.t113 GNDA 0.290879f
C1948 two_stage_opamp_dummy_magic_0.VOUT-.n30 GNDA 0.195025f
C1949 two_stage_opamp_dummy_magic_0.VOUT-.t78 GNDA 0.290879f
C1950 two_stage_opamp_dummy_magic_0.VOUT-.t129 GNDA 0.295834f
C1951 two_stage_opamp_dummy_magic_0.VOUT-.t38 GNDA 0.290879f
C1952 two_stage_opamp_dummy_magic_0.VOUT-.n31 GNDA 0.195025f
C1953 two_stage_opamp_dummy_magic_0.VOUT-.n32 GNDA 0.236339f
C1954 two_stage_opamp_dummy_magic_0.VOUT-.t61 GNDA 0.295834f
C1955 two_stage_opamp_dummy_magic_0.VOUT-.t147 GNDA 0.290879f
C1956 two_stage_opamp_dummy_magic_0.VOUT-.n33 GNDA 0.195025f
C1957 two_stage_opamp_dummy_magic_0.VOUT-.t117 GNDA 0.290879f
C1958 two_stage_opamp_dummy_magic_0.VOUT-.t32 GNDA 0.295834f
C1959 two_stage_opamp_dummy_magic_0.VOUT-.t83 GNDA 0.290879f
C1960 two_stage_opamp_dummy_magic_0.VOUT-.n34 GNDA 0.195025f
C1961 two_stage_opamp_dummy_magic_0.VOUT-.n35 GNDA 0.236339f
C1962 two_stage_opamp_dummy_magic_0.VOUT-.t100 GNDA 0.295834f
C1963 two_stage_opamp_dummy_magic_0.VOUT-.t47 GNDA 0.290879f
C1964 two_stage_opamp_dummy_magic_0.VOUT-.n36 GNDA 0.195025f
C1965 two_stage_opamp_dummy_magic_0.VOUT-.t153 GNDA 0.290879f
C1966 two_stage_opamp_dummy_magic_0.VOUT-.t71 GNDA 0.295834f
C1967 two_stage_opamp_dummy_magic_0.VOUT-.t123 GNDA 0.290879f
C1968 two_stage_opamp_dummy_magic_0.VOUT-.n37 GNDA 0.195025f
C1969 two_stage_opamp_dummy_magic_0.VOUT-.n38 GNDA 0.236339f
C1970 two_stage_opamp_dummy_magic_0.VOUT-.t69 GNDA 0.295834f
C1971 two_stage_opamp_dummy_magic_0.VOUT-.t154 GNDA 0.290879f
C1972 two_stage_opamp_dummy_magic_0.VOUT-.n39 GNDA 0.195025f
C1973 two_stage_opamp_dummy_magic_0.VOUT-.t124 GNDA 0.290879f
C1974 two_stage_opamp_dummy_magic_0.VOUT-.t35 GNDA 0.295834f
C1975 two_stage_opamp_dummy_magic_0.VOUT-.t86 GNDA 0.290879f
C1976 two_stage_opamp_dummy_magic_0.VOUT-.n40 GNDA 0.195025f
C1977 two_stage_opamp_dummy_magic_0.VOUT-.n41 GNDA 0.236339f
C1978 two_stage_opamp_dummy_magic_0.VOUT-.t96 GNDA 0.290879f
C1979 two_stage_opamp_dummy_magic_0.VOUT-.t85 GNDA 0.295834f
C1980 two_stage_opamp_dummy_magic_0.VOUT-.t57 GNDA 0.290879f
C1981 two_stage_opamp_dummy_magic_0.VOUT-.n42 GNDA 0.195025f
C1982 two_stage_opamp_dummy_magic_0.VOUT-.n43 GNDA 0.12726f
C1983 two_stage_opamp_dummy_magic_0.VOUT-.t132 GNDA 0.295213f
C1984 two_stage_opamp_dummy_magic_0.VOUT-.t115 GNDA 0.295213f
C1985 two_stage_opamp_dummy_magic_0.VOUT-.t131 GNDA 0.295834f
C1986 two_stage_opamp_dummy_magic_0.VOUT-.t104 GNDA 0.290879f
C1987 two_stage_opamp_dummy_magic_0.VOUT-.n44 GNDA 0.195025f
C1988 two_stage_opamp_dummy_magic_0.VOUT-.t73 GNDA 0.290879f
C1989 two_stage_opamp_dummy_magic_0.VOUT-.n45 GNDA 0.122715f
C1990 two_stage_opamp_dummy_magic_0.VOUT-.t146 GNDA 0.295213f
C1991 two_stage_opamp_dummy_magic_0.VOUT-.t31 GNDA 0.295834f
C1992 two_stage_opamp_dummy_magic_0.VOUT-.t138 GNDA 0.290879f
C1993 two_stage_opamp_dummy_magic_0.VOUT-.n46 GNDA 0.195025f
C1994 two_stage_opamp_dummy_magic_0.VOUT-.t107 GNDA 0.290879f
C1995 two_stage_opamp_dummy_magic_0.VOUT-.n47 GNDA 0.122715f
C1996 two_stage_opamp_dummy_magic_0.VOUT-.t46 GNDA 0.295213f
C1997 two_stage_opamp_dummy_magic_0.VOUT-.t62 GNDA 0.295834f
C1998 two_stage_opamp_dummy_magic_0.VOUT-.t41 GNDA 0.290879f
C1999 two_stage_opamp_dummy_magic_0.VOUT-.n48 GNDA 0.195025f
C2000 two_stage_opamp_dummy_magic_0.VOUT-.t143 GNDA 0.290879f
C2001 two_stage_opamp_dummy_magic_0.VOUT-.n49 GNDA 0.122715f
C2002 two_stage_opamp_dummy_magic_0.VOUT-.t87 GNDA 0.295213f
C2003 two_stage_opamp_dummy_magic_0.VOUT-.t114 GNDA 0.295834f
C2004 two_stage_opamp_dummy_magic_0.VOUT-.t21 GNDA 0.290879f
C2005 two_stage_opamp_dummy_magic_0.VOUT-.n50 GNDA 0.195025f
C2006 two_stage_opamp_dummy_magic_0.VOUT-.t126 GNDA 0.290879f
C2007 two_stage_opamp_dummy_magic_0.VOUT-.n51 GNDA 0.122715f
C2008 two_stage_opamp_dummy_magic_0.VOUT-.t65 GNDA 0.295213f
C2009 two_stage_opamp_dummy_magic_0.VOUT-.t26 GNDA 0.295457f
C2010 two_stage_opamp_dummy_magic_0.VOUT-.t102 GNDA 0.295213f
C2011 two_stage_opamp_dummy_magic_0.VOUT-.t59 GNDA 0.295457f
C2012 two_stage_opamp_dummy_magic_0.VOUT-.t134 GNDA 0.295213f
C2013 two_stage_opamp_dummy_magic_0.VOUT-.t37 GNDA 0.295457f
C2014 two_stage_opamp_dummy_magic_0.VOUT-.t120 GNDA 0.295213f
C2015 two_stage_opamp_dummy_magic_0.VOUT-.t81 GNDA 0.295457f
C2016 two_stage_opamp_dummy_magic_0.VOUT-.t155 GNDA 0.295213f
C2017 two_stage_opamp_dummy_magic_0.VOUT-.t119 GNDA 0.290879f
C2018 two_stage_opamp_dummy_magic_0.VOUT-.n52 GNDA 0.321963f
C2019 two_stage_opamp_dummy_magic_0.VOUT-.t82 GNDA 0.290879f
C2020 two_stage_opamp_dummy_magic_0.VOUT-.n53 GNDA 0.376503f
C2021 two_stage_opamp_dummy_magic_0.VOUT-.t97 GNDA 0.290879f
C2022 two_stage_opamp_dummy_magic_0.VOUT-.n54 GNDA 0.376503f
C2023 two_stage_opamp_dummy_magic_0.VOUT-.t63 GNDA 0.290879f
C2024 two_stage_opamp_dummy_magic_0.VOUT-.n55 GNDA 0.376503f
C2025 two_stage_opamp_dummy_magic_0.VOUT-.t27 GNDA 0.290879f
C2026 two_stage_opamp_dummy_magic_0.VOUT-.n56 GNDA 0.30927f
C2027 two_stage_opamp_dummy_magic_0.VOUT-.t45 GNDA 0.290879f
C2028 two_stage_opamp_dummy_magic_0.VOUT-.n57 GNDA 0.30927f
C2029 two_stage_opamp_dummy_magic_0.VOUT-.t144 GNDA 0.290879f
C2030 two_stage_opamp_dummy_magic_0.VOUT-.n58 GNDA 0.30927f
C2031 two_stage_opamp_dummy_magic_0.VOUT-.t112 GNDA 0.290879f
C2032 two_stage_opamp_dummy_magic_0.VOUT-.n59 GNDA 0.30927f
C2033 two_stage_opamp_dummy_magic_0.VOUT-.t76 GNDA 0.290879f
C2034 two_stage_opamp_dummy_magic_0.VOUT-.n60 GNDA 0.250185f
C2035 two_stage_opamp_dummy_magic_0.VOUT-.t93 GNDA 0.290879f
C2036 two_stage_opamp_dummy_magic_0.VOUT-.n61 GNDA 0.250185f
C2037 two_stage_opamp_dummy_magic_0.VOUT-.t56 GNDA 0.290879f
C2038 two_stage_opamp_dummy_magic_0.VOUT-.t40 GNDA 0.295834f
C2039 two_stage_opamp_dummy_magic_0.VOUT-.t19 GNDA 0.290879f
C2040 two_stage_opamp_dummy_magic_0.VOUT-.n62 GNDA 0.195025f
C2041 two_stage_opamp_dummy_magic_0.VOUT-.n63 GNDA 0.236339f
C2042 two_stage_opamp_dummy_magic_0.VOUT-.t34 GNDA 0.295834f
C2043 two_stage_opamp_dummy_magic_0.VOUT-.t52 GNDA 0.290879f
C2044 two_stage_opamp_dummy_magic_0.VOUT-.n64 GNDA 0.195025f
C2045 two_stage_opamp_dummy_magic_0.VOUT-.t156 GNDA 0.290879f
C2046 two_stage_opamp_dummy_magic_0.VOUT-.t136 GNDA 0.295834f
C2047 two_stage_opamp_dummy_magic_0.VOUT-.t121 GNDA 0.290879f
C2048 two_stage_opamp_dummy_magic_0.VOUT-.n65 GNDA 0.195025f
C2049 two_stage_opamp_dummy_magic_0.VOUT-.n66 GNDA 0.236339f
C2050 two_stage_opamp_dummy_magic_0.VOUT-.t70 GNDA 0.295834f
C2051 two_stage_opamp_dummy_magic_0.VOUT-.t89 GNDA 0.290879f
C2052 two_stage_opamp_dummy_magic_0.VOUT-.n67 GNDA 0.195025f
C2053 two_stage_opamp_dummy_magic_0.VOUT-.t50 GNDA 0.290879f
C2054 two_stage_opamp_dummy_magic_0.VOUT-.t36 GNDA 0.295834f
C2055 two_stage_opamp_dummy_magic_0.VOUT-.t151 GNDA 0.290879f
C2056 two_stage_opamp_dummy_magic_0.VOUT-.n68 GNDA 0.195025f
C2057 two_stage_opamp_dummy_magic_0.VOUT-.n69 GNDA 0.236339f
C2058 two_stage_opamp_dummy_magic_0.VOUT-.t95 GNDA 0.295834f
C2059 two_stage_opamp_dummy_magic_0.VOUT-.t43 GNDA 0.290879f
C2060 two_stage_opamp_dummy_magic_0.VOUT-.n70 GNDA 0.195025f
C2061 two_stage_opamp_dummy_magic_0.VOUT-.t145 GNDA 0.290879f
C2062 two_stage_opamp_dummy_magic_0.VOUT-.t66 GNDA 0.295834f
C2063 two_stage_opamp_dummy_magic_0.VOUT-.t118 GNDA 0.290879f
C2064 two_stage_opamp_dummy_magic_0.VOUT-.n71 GNDA 0.195025f
C2065 two_stage_opamp_dummy_magic_0.VOUT-.n72 GNDA 0.236339f
C2066 two_stage_opamp_dummy_magic_0.VOUT-.t55 GNDA 0.295834f
C2067 two_stage_opamp_dummy_magic_0.VOUT-.t141 GNDA 0.290879f
C2068 two_stage_opamp_dummy_magic_0.VOUT-.n73 GNDA 0.195025f
C2069 two_stage_opamp_dummy_magic_0.VOUT-.t111 GNDA 0.290879f
C2070 two_stage_opamp_dummy_magic_0.VOUT-.t29 GNDA 0.295834f
C2071 two_stage_opamp_dummy_magic_0.VOUT-.t80 GNDA 0.290879f
C2072 two_stage_opamp_dummy_magic_0.VOUT-.n74 GNDA 0.195025f
C2073 two_stage_opamp_dummy_magic_0.VOUT-.n75 GNDA 0.236339f
C2074 two_stage_opamp_dummy_magic_0.VOUT-.t91 GNDA 0.295834f
C2075 two_stage_opamp_dummy_magic_0.VOUT-.t39 GNDA 0.290879f
C2076 two_stage_opamp_dummy_magic_0.VOUT-.n76 GNDA 0.195025f
C2077 two_stage_opamp_dummy_magic_0.VOUT-.t139 GNDA 0.290879f
C2078 two_stage_opamp_dummy_magic_0.VOUT-.t58 GNDA 0.295834f
C2079 two_stage_opamp_dummy_magic_0.VOUT-.t109 GNDA 0.290879f
C2080 two_stage_opamp_dummy_magic_0.VOUT-.n77 GNDA 0.195025f
C2081 two_stage_opamp_dummy_magic_0.VOUT-.n78 GNDA 0.236339f
C2082 two_stage_opamp_dummy_magic_0.VOUT-.t49 GNDA 0.295834f
C2083 two_stage_opamp_dummy_magic_0.VOUT-.t135 GNDA 0.290879f
C2084 two_stage_opamp_dummy_magic_0.VOUT-.n79 GNDA 0.195025f
C2085 two_stage_opamp_dummy_magic_0.VOUT-.t103 GNDA 0.290879f
C2086 two_stage_opamp_dummy_magic_0.VOUT-.t20 GNDA 0.295834f
C2087 two_stage_opamp_dummy_magic_0.VOUT-.t72 GNDA 0.290879f
C2088 two_stage_opamp_dummy_magic_0.VOUT-.n80 GNDA 0.195025f
C2089 two_stage_opamp_dummy_magic_0.VOUT-.n81 GNDA 0.236339f
C2090 two_stage_opamp_dummy_magic_0.VOUT-.t148 GNDA 0.295834f
C2091 two_stage_opamp_dummy_magic_0.VOUT-.t99 GNDA 0.290879f
C2092 two_stage_opamp_dummy_magic_0.VOUT-.n82 GNDA 0.195025f
C2093 two_stage_opamp_dummy_magic_0.VOUT-.t68 GNDA 0.290879f
C2094 two_stage_opamp_dummy_magic_0.VOUT-.t122 GNDA 0.295834f
C2095 two_stage_opamp_dummy_magic_0.VOUT-.t33 GNDA 0.290879f
C2096 two_stage_opamp_dummy_magic_0.VOUT-.n83 GNDA 0.195025f
C2097 two_stage_opamp_dummy_magic_0.VOUT-.n84 GNDA 0.236339f
C2098 two_stage_opamp_dummy_magic_0.VOUT-.t44 GNDA 0.295834f
C2099 two_stage_opamp_dummy_magic_0.VOUT-.t133 GNDA 0.290879f
C2100 two_stage_opamp_dummy_magic_0.VOUT-.n85 GNDA 0.195025f
C2101 two_stage_opamp_dummy_magic_0.VOUT-.t98 GNDA 0.290879f
C2102 two_stage_opamp_dummy_magic_0.VOUT-.t152 GNDA 0.295834f
C2103 two_stage_opamp_dummy_magic_0.VOUT-.t67 GNDA 0.290879f
C2104 two_stage_opamp_dummy_magic_0.VOUT-.n86 GNDA 0.195025f
C2105 two_stage_opamp_dummy_magic_0.VOUT-.n87 GNDA 0.236339f
C2106 two_stage_opamp_dummy_magic_0.VOUT-.t142 GNDA 0.295834f
C2107 two_stage_opamp_dummy_magic_0.VOUT-.t94 GNDA 0.290879f
C2108 two_stage_opamp_dummy_magic_0.VOUT-.n88 GNDA 0.195025f
C2109 two_stage_opamp_dummy_magic_0.VOUT-.t60 GNDA 0.290879f
C2110 two_stage_opamp_dummy_magic_0.VOUT-.t116 GNDA 0.295834f
C2111 two_stage_opamp_dummy_magic_0.VOUT-.t30 GNDA 0.290879f
C2112 two_stage_opamp_dummy_magic_0.VOUT-.n89 GNDA 0.195025f
C2113 two_stage_opamp_dummy_magic_0.VOUT-.n90 GNDA 0.236339f
C2114 two_stage_opamp_dummy_magic_0.VOUT-.t77 GNDA 0.295834f
C2115 two_stage_opamp_dummy_magic_0.VOUT-.t127 GNDA 0.290879f
C2116 two_stage_opamp_dummy_magic_0.VOUT-.n91 GNDA 0.195025f
C2117 two_stage_opamp_dummy_magic_0.VOUT-.t22 GNDA 0.290879f
C2118 two_stage_opamp_dummy_magic_0.VOUT-.n92 GNDA 0.236339f
C2119 two_stage_opamp_dummy_magic_0.VOUT-.t53 GNDA 0.290879f
C2120 two_stage_opamp_dummy_magic_0.VOUT-.n93 GNDA 0.12726f
C2121 two_stage_opamp_dummy_magic_0.VOUT-.t105 GNDA 0.290879f
C2122 two_stage_opamp_dummy_magic_0.VOUT-.n94 GNDA 0.238316f
C2123 two_stage_opamp_dummy_magic_0.VOUT-.n95 GNDA 0.291354f
C2124 two_stage_opamp_dummy_magic_0.VOUT-.n96 GNDA 0.165389f
C2125 two_stage_opamp_dummy_magic_0.VOUT-.t6 GNDA 0.084162f
C2126 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2127 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2128 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2129 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2130 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2131 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2132 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2133 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2134 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2135 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2136 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2137 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2138 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2139 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2140 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2141 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2142 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2143 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2144 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2145 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2146 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.050131f
C2147 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2148 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2149 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.04969f
C2150 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.186051f
C2151 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2152 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2153 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2154 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.096484f
C2155 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.117322f
C2156 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2157 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2158 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2159 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2160 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2161 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2162 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2163 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2164 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2165 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2166 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2167 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2168 bgr_0.cap_res1.t6 GNDA 0.417173f
C2169 bgr_0.cap_res1.t10 GNDA 0.418684f
C2170 bgr_0.cap_res1.t0 GNDA 0.417173f
C2171 bgr_0.cap_res1.t14 GNDA 0.418684f
C2172 bgr_0.cap_res1.t3 GNDA 0.417173f
C2173 bgr_0.cap_res1.t7 GNDA 0.418684f
C2174 bgr_0.cap_res1.t15 GNDA 0.417173f
C2175 bgr_0.cap_res1.t9 GNDA 0.418684f
C2176 bgr_0.cap_res1.t8 GNDA 0.417173f
C2177 bgr_0.cap_res1.t12 GNDA 0.418684f
C2178 bgr_0.cap_res1.t1 GNDA 0.417173f
C2179 bgr_0.cap_res1.t16 GNDA 0.418684f
C2180 bgr_0.cap_res1.t13 GNDA 0.417173f
C2181 bgr_0.cap_res1.t19 GNDA 0.418684f
C2182 bgr_0.cap_res1.t5 GNDA 0.417173f
C2183 bgr_0.cap_res1.t2 GNDA 0.418684f
C2184 bgr_0.cap_res1.n0 GNDA 0.279631f
C2185 bgr_0.cap_res1.t4 GNDA 0.222685f
C2186 bgr_0.cap_res1.n1 GNDA 0.303406f
C2187 bgr_0.cap_res1.t18 GNDA 0.222685f
C2188 bgr_0.cap_res1.n2 GNDA 0.303406f
C2189 bgr_0.cap_res1.t11 GNDA 0.222685f
C2190 bgr_0.cap_res1.n3 GNDA 0.303406f
C2191 bgr_0.cap_res1.t17 GNDA 0.649059f
C2192 bgr_0.cap_res1.t20 GNDA 0.10618f
C2193 bgr_0.1st_Vout_1.n0 GNDA 0.573726f
C2194 bgr_0.1st_Vout_1.n1 GNDA 1.42916f
C2195 bgr_0.1st_Vout_1.n2 GNDA 1.78489f
C2196 bgr_0.1st_Vout_1.n3 GNDA 0.125562f
C2197 bgr_0.1st_Vout_1.t20 GNDA 0.352846f
C2198 bgr_0.1st_Vout_1.t11 GNDA 0.346937f
C2199 bgr_0.1st_Vout_1.t32 GNDA 0.346937f
C2200 bgr_0.1st_Vout_1.t29 GNDA 0.352846f
C2201 bgr_0.1st_Vout_1.t34 GNDA 0.346937f
C2202 bgr_0.1st_Vout_1.t25 GNDA 0.352846f
C2203 bgr_0.1st_Vout_1.t21 GNDA 0.346937f
C2204 bgr_0.1st_Vout_1.t12 GNDA 0.346937f
C2205 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C2206 bgr_0.1st_Vout_1.t16 GNDA 0.346937f
C2207 bgr_0.1st_Vout_1.t33 GNDA 0.352846f
C2208 bgr_0.1st_Vout_1.t26 GNDA 0.346937f
C2209 bgr_0.1st_Vout_1.t22 GNDA 0.346937f
C2210 bgr_0.1st_Vout_1.t17 GNDA 0.352846f
C2211 bgr_0.1st_Vout_1.t24 GNDA 0.346937f
C2212 bgr_0.1st_Vout_1.t28 GNDA 0.352846f
C2213 bgr_0.1st_Vout_1.t23 GNDA 0.346937f
C2214 bgr_0.1st_Vout_1.t13 GNDA 0.346937f
C2215 bgr_0.1st_Vout_1.t18 GNDA 0.346937f
C2216 bgr_0.1st_Vout_1.t36 GNDA 0.346937f
C2217 bgr_0.1st_Vout_1.t30 GNDA 0.022665f
C2218 bgr_0.1st_Vout_1.n4 GNDA 0.021864f
C2219 bgr_0.1st_Vout_1.t14 GNDA 0.013213f
C2220 bgr_0.1st_Vout_1.t31 GNDA 0.013213f
C2221 bgr_0.1st_Vout_1.n5 GNDA 0.029393f
C2222 bgr_0.1st_Vout_1.t1 GNDA 0.018268f
C2223 bgr_0.1st_Vout_1.n6 GNDA 0.012529f
C2224 bgr_0.1st_Vout_1.n7 GNDA 0.189508f
C2225 bgr_0.1st_Vout_1.n8 GNDA 0.011336f
C2226 bgr_0.1st_Vout_1.n9 GNDA 0.020958f
C2227 bgr_0.1st_Vout_1.t19 GNDA 0.013213f
C2228 bgr_0.1st_Vout_1.t27 GNDA 0.013213f
C2229 bgr_0.1st_Vout_1.n10 GNDA 0.029393f
C2230 bgr_0.1st_Vout_1.n11 GNDA 0.021864f
C2231 bgr_0.1st_Vout_1.t15 GNDA 0.020738f
C2232 VDDA.t249 GNDA 0.020007f
C2233 VDDA.t224 GNDA 0.020007f
C2234 VDDA.n0 GNDA 0.082739f
C2235 VDDA.t119 GNDA 0.020007f
C2236 VDDA.t46 GNDA 0.020007f
C2237 VDDA.n1 GNDA 0.082421f
C2238 VDDA.n2 GNDA 0.114273f
C2239 VDDA.t186 GNDA 0.020007f
C2240 VDDA.t11 GNDA 0.020007f
C2241 VDDA.n3 GNDA 0.082421f
C2242 VDDA.n4 GNDA 0.059629f
C2243 VDDA.t30 GNDA 0.020007f
C2244 VDDA.t252 GNDA 0.020007f
C2245 VDDA.n5 GNDA 0.082421f
C2246 VDDA.n6 GNDA 0.059629f
C2247 VDDA.t14 GNDA 0.020007f
C2248 VDDA.t7 GNDA 0.020007f
C2249 VDDA.n7 GNDA 0.082421f
C2250 VDDA.n8 GNDA 0.059629f
C2251 VDDA.t85 GNDA 0.020007f
C2252 VDDA.t47 GNDA 0.020007f
C2253 VDDA.n9 GNDA 0.082421f
C2254 VDDA.n10 GNDA 0.141701f
C2255 VDDA.n11 GNDA 0.064606f
C2256 VDDA.n12 GNDA 0.17248f
C2257 VDDA.t314 GNDA 0.012566f
C2258 VDDA.n13 GNDA 0.026738f
C2259 VDDA.t423 GNDA 0.012566f
C2260 VDDA.n14 GNDA 0.026738f
C2261 VDDA.n15 GNDA 0.038823f
C2262 VDDA.n16 GNDA 0.065254f
C2263 VDDA.n17 GNDA 0.173903f
C2264 VDDA.t384 GNDA 0.012566f
C2265 VDDA.n18 GNDA 0.026738f
C2266 VDDA.t357 GNDA 0.012566f
C2267 VDDA.n19 GNDA 0.026738f
C2268 VDDA.n20 GNDA 0.03618f
C2269 VDDA.n21 GNDA 0.044911f
C2270 VDDA.n22 GNDA 0.173903f
C2271 VDDA.t356 GNDA 0.169175f
C2272 VDDA.t136 GNDA 0.104537f
C2273 VDDA.t75 GNDA 0.104537f
C2274 VDDA.t15 GNDA 0.104537f
C2275 VDDA.t134 GNDA 0.104537f
C2276 VDDA.t56 GNDA 0.078403f
C2277 VDDA.t383 GNDA 0.169175f
C2278 VDDA.t217 GNDA 0.104537f
C2279 VDDA.t256 GNDA 0.104537f
C2280 VDDA.t135 GNDA 0.104537f
C2281 VDDA.t6 GNDA 0.104537f
C2282 VDDA.t235 GNDA 0.078403f
C2283 VDDA.n23 GNDA 0.065901f
C2284 VDDA.n24 GNDA 0.052269f
C2285 VDDA.n25 GNDA 0.065901f
C2286 VDDA.n26 GNDA 0.044016f
C2287 VDDA.n27 GNDA 0.035613f
C2288 VDDA.n28 GNDA 0.082804f
C2289 VDDA.n29 GNDA 0.082804f
C2290 VDDA.n30 GNDA 0.17248f
C2291 VDDA.t422 GNDA 0.165763f
C2292 VDDA.t129 GNDA 0.102703f
C2293 VDDA.t29 GNDA 0.102703f
C2294 VDDA.t450 GNDA 0.102703f
C2295 VDDA.t21 GNDA 0.102703f
C2296 VDDA.t97 GNDA 0.077027f
C2297 VDDA.t313 GNDA 0.165763f
C2298 VDDA.t57 GNDA 0.102703f
C2299 VDDA.t76 GNDA 0.102703f
C2300 VDDA.t55 GNDA 0.102703f
C2301 VDDA.t214 GNDA 0.102703f
C2302 VDDA.t84 GNDA 0.077027f
C2303 VDDA.n31 GNDA 0.065901f
C2304 VDDA.n32 GNDA 0.051352f
C2305 VDDA.n33 GNDA 0.065901f
C2306 VDDA.n34 GNDA 0.043806f
C2307 VDDA.n35 GNDA 0.035613f
C2308 VDDA.n36 GNDA 0.068943f
C2309 VDDA.n37 GNDA 0.204887f
C2310 VDDA.t10 GNDA 0.040014f
C2311 VDDA.t126 GNDA 0.040014f
C2312 VDDA.n38 GNDA 0.160532f
C2313 VDDA.n39 GNDA 0.081554f
C2314 VDDA.t320 GNDA 0.039861f
C2315 VDDA.n40 GNDA 0.080891f
C2316 VDDA.n41 GNDA 0.053975f
C2317 VDDA.n42 GNDA 0.076186f
C2318 VDDA.t360 GNDA 0.04427f
C2319 VDDA.t358 GNDA 0.019386f
C2320 VDDA.n43 GNDA 0.070225f
C2321 VDDA.n44 GNDA 0.041341f
C2322 VDDA.t326 GNDA 0.04427f
C2323 VDDA.t324 GNDA 0.019386f
C2324 VDDA.n45 GNDA 0.070225f
C2325 VDDA.n46 GNDA 0.041341f
C2326 VDDA.n47 GNDA 0.044016f
C2327 VDDA.n48 GNDA 0.076186f
C2328 VDDA.n49 GNDA 0.220247f
C2329 VDDA.t325 GNDA 0.272769f
C2330 VDDA.t48 GNDA 0.157723f
C2331 VDDA.t124 GNDA 0.157723f
C2332 VDDA.t187 GNDA 0.157723f
C2333 VDDA.t118 GNDA 0.157723f
C2334 VDDA.t193 GNDA 0.118292f
C2335 VDDA.n50 GNDA 0.078861f
C2336 VDDA.t8 GNDA 0.118292f
C2337 VDDA.t192 GNDA 0.157723f
C2338 VDDA.t28 GNDA 0.157723f
C2339 VDDA.t253 GNDA 0.157723f
C2340 VDDA.t31 GNDA 0.157723f
C2341 VDDA.t359 GNDA 0.272769f
C2342 VDDA.n51 GNDA 0.220247f
C2343 VDDA.n52 GNDA 0.053975f
C2344 VDDA.n53 GNDA 0.102138f
C2345 VDDA.t348 GNDA 0.039861f
C2346 VDDA.t189 GNDA 0.040014f
C2347 VDDA.t13 GNDA 0.040014f
C2348 VDDA.n54 GNDA 0.160532f
C2349 VDDA.n55 GNDA 0.081554f
C2350 VDDA.t191 GNDA 0.040014f
C2351 VDDA.t27 GNDA 0.040014f
C2352 VDDA.n56 GNDA 0.160532f
C2353 VDDA.n57 GNDA 0.081554f
C2354 VDDA.t251 GNDA 0.040014f
C2355 VDDA.t185 GNDA 0.040014f
C2356 VDDA.n58 GNDA 0.160532f
C2357 VDDA.n59 GNDA 0.081554f
C2358 VDDA.t50 GNDA 0.040014f
C2359 VDDA.t195 GNDA 0.040014f
C2360 VDDA.n60 GNDA 0.160532f
C2361 VDDA.n61 GNDA 0.171374f
C2362 VDDA.n62 GNDA 0.129391f
C2363 VDDA.t346 GNDA 0.048365f
C2364 VDDA.n63 GNDA 0.092538f
C2365 VDDA.n64 GNDA 0.054063f
C2366 VDDA.n65 GNDA 0.356054f
C2367 VDDA.n66 GNDA 0.356054f
C2368 VDDA.t319 GNDA 0.549961f
C2369 VDDA.t9 GNDA 0.304442f
C2370 VDDA.t125 GNDA 0.304442f
C2371 VDDA.t188 GNDA 0.304442f
C2372 VDDA.t12 GNDA 0.304442f
C2373 VDDA.t190 GNDA 0.228331f
C2374 VDDA.n67 GNDA 0.080891f
C2375 VDDA.n68 GNDA 0.103682f
C2376 VDDA.n69 GNDA 0.103682f
C2377 VDDA.t347 GNDA 0.549961f
C2378 VDDA.t194 GNDA 0.304442f
C2379 VDDA.t49 GNDA 0.304442f
C2380 VDDA.t184 GNDA 0.304442f
C2381 VDDA.t250 GNDA 0.304442f
C2382 VDDA.t26 GNDA 0.228331f
C2383 VDDA.n70 GNDA 0.152221f
C2384 VDDA.n71 GNDA 0.103006f
C2385 VDDA.n72 GNDA 0.0699f
C2386 VDDA.n73 GNDA 0.054063f
C2387 VDDA.t318 GNDA 0.048365f
C2388 VDDA.n74 GNDA 0.092538f
C2389 VDDA.n75 GNDA 0.129057f
C2390 VDDA.n76 GNDA 0.114829f
C2391 VDDA.n77 GNDA 0.097701f
C2392 VDDA.t45 GNDA 0.023342f
C2393 VDDA.t447 GNDA 0.023342f
C2394 VDDA.n78 GNDA 0.081177f
C2395 VDDA.t131 GNDA 0.023342f
C2396 VDDA.t244 GNDA 0.023342f
C2397 VDDA.n79 GNDA 0.08089f
C2398 VDDA.n80 GNDA 0.152712f
C2399 VDDA.t246 GNDA 0.023342f
C2400 VDDA.t425 GNDA 0.023342f
C2401 VDDA.n81 GNDA 0.081177f
C2402 VDDA.t43 GNDA 0.023342f
C2403 VDDA.t205 GNDA 0.023342f
C2404 VDDA.n82 GNDA 0.08089f
C2405 VDDA.n83 GNDA 0.152712f
C2406 VDDA.n84 GNDA 0.021341f
C2407 VDDA.n85 GNDA 0.066451f
C2408 VDDA.n86 GNDA 0.09036f
C2409 VDDA.t414 GNDA 0.115149f
C2410 VDDA.t412 GNDA 0.040646f
C2411 VDDA.n87 GNDA 0.07512f
C2412 VDDA.n88 GNDA 0.048426f
C2413 VDDA.t369 GNDA 0.115149f
C2414 VDDA.t367 GNDA 0.040646f
C2415 VDDA.n89 GNDA 0.07512f
C2416 VDDA.n90 GNDA 0.048426f
C2417 VDDA.n91 GNDA 0.048017f
C2418 VDDA.n92 GNDA 0.09036f
C2419 VDDA.n93 GNDA 0.26929f
C2420 VDDA.t368 GNDA 0.401954f
C2421 VDDA.t44 GNDA 0.232082f
C2422 VDDA.t446 GNDA 0.232082f
C2423 VDDA.t130 GNDA 0.232082f
C2424 VDDA.t243 GNDA 0.232082f
C2425 VDDA.t179 GNDA 0.174062f
C2426 VDDA.n94 GNDA 0.116041f
C2427 VDDA.t107 GNDA 0.174062f
C2428 VDDA.t42 GNDA 0.232082f
C2429 VDDA.t204 GNDA 0.232082f
C2430 VDDA.t245 GNDA 0.232082f
C2431 VDDA.t424 GNDA 0.232082f
C2432 VDDA.t413 GNDA 0.401954f
C2433 VDDA.n95 GNDA 0.26929f
C2434 VDDA.n96 GNDA 0.066451f
C2435 VDDA.n97 GNDA 0.093028f
C2436 VDDA.t180 GNDA 0.023342f
C2437 VDDA.t108 GNDA 0.023342f
C2438 VDDA.n98 GNDA 0.076104f
C2439 VDDA.n99 GNDA 0.051942f
C2440 VDDA.n100 GNDA 0.043635f
C2441 VDDA.t128 GNDA 0.020007f
C2442 VDDA.t238 GNDA 0.020007f
C2443 VDDA.n101 GNDA 0.082739f
C2444 VDDA.t463 GNDA 0.020007f
C2445 VDDA.t169 GNDA 0.020007f
C2446 VDDA.n102 GNDA 0.082421f
C2447 VDDA.n103 GNDA 0.114273f
C2448 VDDA.t226 GNDA 0.020007f
C2449 VDDA.t102 GNDA 0.020007f
C2450 VDDA.n104 GNDA 0.082421f
C2451 VDDA.n105 GNDA 0.059629f
C2452 VDDA.t468 GNDA 0.020007f
C2453 VDDA.t83 GNDA 0.020007f
C2454 VDDA.n106 GNDA 0.082421f
C2455 VDDA.n107 GNDA 0.059629f
C2456 VDDA.t111 GNDA 0.020007f
C2457 VDDA.t429 GNDA 0.020007f
C2458 VDDA.n108 GNDA 0.082421f
C2459 VDDA.n109 GNDA 0.059629f
C2460 VDDA.t70 GNDA 0.020007f
C2461 VDDA.t16 GNDA 0.020007f
C2462 VDDA.n110 GNDA 0.082421f
C2463 VDDA.n111 GNDA 0.172215f
C2464 VDDA.t59 GNDA 0.040014f
C2465 VDDA.t449 GNDA 0.040014f
C2466 VDDA.n112 GNDA 0.160532f
C2467 VDDA.n113 GNDA 0.081554f
C2468 VDDA.t375 GNDA 0.039861f
C2469 VDDA.n114 GNDA 0.053975f
C2470 VDDA.n115 GNDA 0.076186f
C2471 VDDA.t381 GNDA 0.04427f
C2472 VDDA.t379 GNDA 0.019386f
C2473 VDDA.n116 GNDA 0.070225f
C2474 VDDA.n117 GNDA 0.041341f
C2475 VDDA.t354 GNDA 0.04427f
C2476 VDDA.t352 GNDA 0.019386f
C2477 VDDA.n118 GNDA 0.070225f
C2478 VDDA.n119 GNDA 0.041341f
C2479 VDDA.n120 GNDA 0.044016f
C2480 VDDA.n121 GNDA 0.076186f
C2481 VDDA.n122 GNDA 0.220247f
C2482 VDDA.t353 GNDA 0.272769f
C2483 VDDA.t172 GNDA 0.157723f
C2484 VDDA.t428 GNDA 0.157723f
C2485 VDDA.t96 GNDA 0.157723f
C2486 VDDA.t181 GNDA 0.157723f
C2487 VDDA.t451 GNDA 0.118292f
C2488 VDDA.n123 GNDA 0.078861f
C2489 VDDA.t237 GNDA 0.118292f
C2490 VDDA.t462 GNDA 0.157723f
C2491 VDDA.t236 GNDA 0.157723f
C2492 VDDA.t225 GNDA 0.157723f
C2493 VDDA.t127 GNDA 0.157723f
C2494 VDDA.t380 GNDA 0.272769f
C2495 VDDA.n124 GNDA 0.220247f
C2496 VDDA.n125 GNDA 0.053975f
C2497 VDDA.n126 GNDA 0.102138f
C2498 VDDA.n127 GNDA 0.0699f
C2499 VDDA.n128 GNDA 0.103682f
C2500 VDDA.n129 GNDA 0.103682f
C2501 VDDA.n130 GNDA 0.103006f
C2502 VDDA.t342 GNDA 0.039861f
C2503 VDDA.t465 GNDA 0.040014f
C2504 VDDA.t154 GNDA 0.040014f
C2505 VDDA.n131 GNDA 0.160532f
C2506 VDDA.n132 GNDA 0.081554f
C2507 VDDA.t467 GNDA 0.040014f
C2508 VDDA.t168 GNDA 0.040014f
C2509 VDDA.n133 GNDA 0.160532f
C2510 VDDA.n134 GNDA 0.081554f
C2511 VDDA.t110 GNDA 0.040014f
C2512 VDDA.t113 GNDA 0.040014f
C2513 VDDA.n135 GNDA 0.160532f
C2514 VDDA.n136 GNDA 0.081554f
C2515 VDDA.t171 GNDA 0.040014f
C2516 VDDA.t431 GNDA 0.040014f
C2517 VDDA.n137 GNDA 0.160532f
C2518 VDDA.n138 GNDA 0.171374f
C2519 VDDA.n139 GNDA 0.129391f
C2520 VDDA.t340 GNDA 0.048365f
C2521 VDDA.n140 GNDA 0.092538f
C2522 VDDA.n141 GNDA 0.054063f
C2523 VDDA.n142 GNDA 0.080891f
C2524 VDDA.n143 GNDA 0.356054f
C2525 VDDA.t341 GNDA 0.549961f
C2526 VDDA.t170 GNDA 0.304442f
C2527 VDDA.t430 GNDA 0.304442f
C2528 VDDA.t109 GNDA 0.304442f
C2529 VDDA.t112 GNDA 0.304442f
C2530 VDDA.t466 GNDA 0.228331f
C2531 VDDA.n144 GNDA 0.152221f
C2532 VDDA.t167 GNDA 0.228331f
C2533 VDDA.t464 GNDA 0.304442f
C2534 VDDA.t153 GNDA 0.304442f
C2535 VDDA.t58 GNDA 0.304442f
C2536 VDDA.t448 GNDA 0.304442f
C2537 VDDA.t374 GNDA 0.549961f
C2538 VDDA.n145 GNDA 0.356054f
C2539 VDDA.n146 GNDA 0.080891f
C2540 VDDA.n147 GNDA 0.054063f
C2541 VDDA.t373 GNDA 0.048365f
C2542 VDDA.n148 GNDA 0.092538f
C2543 VDDA.n149 GNDA 0.129057f
C2544 VDDA.n150 GNDA 0.098824f
C2545 VDDA.n152 GNDA 0.051063f
C2546 VDDA.n153 GNDA 0.063348f
C2547 VDDA.n155 GNDA 0.051063f
C2548 VDDA.n157 GNDA 0.051063f
C2549 VDDA.n159 GNDA 0.051063f
C2550 VDDA.n161 GNDA 0.051063f
C2551 VDDA.n163 GNDA 0.051063f
C2552 VDDA.n165 GNDA 0.051063f
C2553 VDDA.n167 GNDA 0.051063f
C2554 VDDA.n169 GNDA 0.051063f
C2555 VDDA.n171 GNDA 0.08356f
C2556 VDDA.t399 GNDA 0.012151f
C2557 VDDA.n172 GNDA 0.018041f
C2558 VDDA.n173 GNDA 0.015963f
C2559 VDDA.n174 GNDA 0.054519f
C2560 VDDA.n175 GNDA 0.209355f
C2561 VDDA.n176 GNDA 0.209355f
C2562 VDDA.t404 GNDA 0.165763f
C2563 VDDA.t62 GNDA 0.102703f
C2564 VDDA.t100 GNDA 0.102703f
C2565 VDDA.t141 GNDA 0.102703f
C2566 VDDA.t98 GNDA 0.102703f
C2567 VDDA.t22 GNDA 0.102703f
C2568 VDDA.t92 GNDA 0.102703f
C2569 VDDA.t103 GNDA 0.102703f
C2570 VDDA.t88 GNDA 0.102703f
C2571 VDDA.t159 GNDA 0.102703f
C2572 VDDA.t145 GNDA 0.077027f
C2573 VDDA.t398 GNDA 0.165763f
C2574 VDDA.t155 GNDA 0.102703f
C2575 VDDA.t143 GNDA 0.102703f
C2576 VDDA.t165 GNDA 0.102703f
C2577 VDDA.t86 GNDA 0.102703f
C2578 VDDA.t24 GNDA 0.102703f
C2579 VDDA.t90 GNDA 0.102703f
C2580 VDDA.t64 GNDA 0.102703f
C2581 VDDA.t161 GNDA 0.102703f
C2582 VDDA.t139 GNDA 0.102703f
C2583 VDDA.t157 GNDA 0.077027f
C2584 VDDA.n177 GNDA 0.063348f
C2585 VDDA.n178 GNDA 0.102385f
C2586 VDDA.n179 GNDA 0.102385f
C2587 VDDA.n180 GNDA 0.051352f
C2588 VDDA.n181 GNDA 0.102385f
C2589 VDDA.n182 GNDA 0.080695f
C2590 VDDA.n183 GNDA 0.054519f
C2591 VDDA.n184 GNDA 0.015963f
C2592 VDDA.t405 GNDA 0.012151f
C2593 VDDA.n185 GNDA 0.017601f
C2594 VDDA.n186 GNDA 0.062948f
C2595 VDDA.n187 GNDA 0.049351f
C2596 VDDA.n188 GNDA 0.254562f
C2597 VDDA.n189 GNDA 0.242116f
C2598 VDDA.t433 GNDA 0.023342f
C2599 VDDA.t117 GNDA 0.023342f
C2600 VDDA.n190 GNDA 0.081177f
C2601 VDDA.t216 GNDA 0.023342f
C2602 VDDA.t223 GNDA 0.023342f
C2603 VDDA.n191 GNDA 0.08089f
C2604 VDDA.n192 GNDA 0.152712f
C2605 VDDA.t82 GNDA 0.023342f
C2606 VDDA.t248 GNDA 0.023342f
C2607 VDDA.n193 GNDA 0.081177f
C2608 VDDA.t242 GNDA 0.023342f
C2609 VDDA.t74 GNDA 0.023342f
C2610 VDDA.n194 GNDA 0.08089f
C2611 VDDA.n195 GNDA 0.152712f
C2612 VDDA.n196 GNDA 0.021341f
C2613 VDDA.n197 GNDA 0.066451f
C2614 VDDA.n198 GNDA 0.09036f
C2615 VDDA.t390 GNDA 0.115149f
C2616 VDDA.t388 GNDA 0.040646f
C2617 VDDA.n199 GNDA 0.07512f
C2618 VDDA.n200 GNDA 0.048426f
C2619 VDDA.t363 GNDA 0.115149f
C2620 VDDA.t361 GNDA 0.040646f
C2621 VDDA.n201 GNDA 0.07512f
C2622 VDDA.n202 GNDA 0.048426f
C2623 VDDA.n203 GNDA 0.048017f
C2624 VDDA.n204 GNDA 0.09036f
C2625 VDDA.n205 GNDA 0.26929f
C2626 VDDA.t362 GNDA 0.401954f
C2627 VDDA.t432 GNDA 0.232082f
C2628 VDDA.t116 GNDA 0.232082f
C2629 VDDA.t215 GNDA 0.232082f
C2630 VDDA.t222 GNDA 0.232082f
C2631 VDDA.t132 GNDA 0.174062f
C2632 VDDA.n206 GNDA 0.116041f
C2633 VDDA.t233 GNDA 0.174062f
C2634 VDDA.t241 GNDA 0.232082f
C2635 VDDA.t73 GNDA 0.232082f
C2636 VDDA.t81 GNDA 0.232082f
C2637 VDDA.t247 GNDA 0.232082f
C2638 VDDA.t389 GNDA 0.401954f
C2639 VDDA.n207 GNDA 0.26929f
C2640 VDDA.n208 GNDA 0.066451f
C2641 VDDA.n209 GNDA 0.093028f
C2642 VDDA.t133 GNDA 0.023342f
C2643 VDDA.t234 GNDA 0.023342f
C2644 VDDA.n210 GNDA 0.076104f
C2645 VDDA.n211 GNDA 0.051942f
C2646 VDDA.n212 GNDA 0.043635f
C2647 VDDA.n213 GNDA 0.209122f
C2648 VDDA.n214 GNDA 0.082029f
C2649 VDDA.n216 GNDA 0.065075f
C2650 VDDA.n217 GNDA 0.012004f
C2651 VDDA.n218 GNDA 0.035459f
C2652 VDDA.n219 GNDA 0.035459f
C2653 VDDA.n220 GNDA 0.036156f
C2654 VDDA.n221 GNDA 0.09085f
C2655 VDDA.n222 GNDA 0.012004f
C2656 VDDA.n223 GNDA 0.053322f
C2657 VDDA.n224 GNDA 0.053322f
C2658 VDDA.n225 GNDA 0.053321f
C2659 VDDA.t232 GNDA 0.021341f
C2660 VDDA.n226 GNDA 0.074056f
C2661 VDDA.t372 GNDA 0.097478f
C2662 VDDA.n227 GNDA 0.048338f
C2663 VDDA.n228 GNDA 0.046404f
C2664 VDDA.t370 GNDA 0.037039f
C2665 VDDA.n229 GNDA 0.039214f
C2666 VDDA.n230 GNDA 0.029353f
C2667 VDDA.n231 GNDA 0.045608f
C2668 VDDA.n232 GNDA 0.299005f
C2669 VDDA.t371 GNDA 0.284228f
C2670 VDDA.n233 GNDA 0.092533f
C2671 VDDA.n234 GNDA 0.023133f
C2672 VDDA.t231 GNDA 0.129546f
C2673 VDDA.t392 GNDA 0.307361f
C2674 VDDA.n235 GNDA 0.302101f
C2675 VDDA.n236 GNDA 0.047326f
C2676 VDDA.n237 GNDA 0.030348f
C2677 VDDA.t391 GNDA 0.037705f
C2678 VDDA.n238 GNDA 0.039214f
C2679 VDDA.t393 GNDA 0.076137f
C2680 VDDA.n239 GNDA 0.052252f
C2681 VDDA.n240 GNDA 0.109851f
C2682 VDDA.n241 GNDA 0.071975f
C2683 VDDA.t323 GNDA 0.015589f
C2684 VDDA.n242 GNDA 0.016935f
C2685 VDDA.t321 GNDA 0.013078f
C2686 VDDA.n243 GNDA 0.016557f
C2687 VDDA.n244 GNDA 0.021319f
C2688 VDDA.n245 GNDA 0.029918f
C2689 VDDA.n246 GNDA 0.159579f
C2690 VDDA.t322 GNDA 0.176746f
C2691 VDDA.t173 GNDA 0.120043f
C2692 VDDA.t337 GNDA 0.176746f
C2693 VDDA.n247 GNDA 0.159579f
C2694 VDDA.n248 GNDA 0.029918f
C2695 VDDA.n249 GNDA 0.021319f
C2696 VDDA.t336 GNDA 0.013078f
C2697 VDDA.n250 GNDA 0.016557f
C2698 VDDA.t339 GNDA 0.015589f
C2699 VDDA.n251 GNDA 0.018904f
C2700 VDDA.n252 GNDA 0.074281f
C2701 VDDA.n253 GNDA 0.216216f
C2702 VDDA.n254 GNDA 4.41322f
C2703 VDDA.t470 GNDA 0.73729f
C2704 VDDA.t471 GNDA 0.78581f
C2705 VDDA.t469 GNDA 0.78581f
C2706 VDDA.t472 GNDA 0.75352f
C2707 VDDA.n255 GNDA 0.526732f
C2708 VDDA.n256 GNDA 0.255726f
C2709 VDDA.n257 GNDA 0.327858f
C2710 VDDA.n258 GNDA 2.34238f
C2711 VDDA.n259 GNDA 0.021341f
C2712 VDDA.n260 GNDA 0.016152f
C2713 VDDA.n261 GNDA 0.016152f
C2714 VDDA.n262 GNDA 0.047203f
C2715 VDDA.n263 GNDA 0.021341f
C2716 VDDA.t351 GNDA 0.025053f
C2717 VDDA.t349 GNDA 0.016508f
C2718 VDDA.n264 GNDA 0.039301f
C2719 VDDA.n265 GNDA 0.055921f
C2720 VDDA.n266 GNDA 0.105129f
C2721 VDDA.n267 GNDA 0.105129f
C2722 VDDA.t317 GNDA 0.025053f
C2723 VDDA.t315 GNDA 0.016508f
C2724 VDDA.n268 GNDA 0.039301f
C2725 VDDA.n269 GNDA 0.080028f
C2726 VDDA.n270 GNDA 0.055921f
C2727 VDDA.n271 GNDA 0.021341f
C2728 VDDA.n272 GNDA 0.016152f
C2729 VDDA.n273 GNDA 0.016888f
C2730 VDDA.n274 GNDA 0.016774f
C2731 VDDA.n275 GNDA 0.130396f
C2732 VDDA.n276 GNDA 0.016774f
C2733 VDDA.n277 GNDA 0.067923f
C2734 VDDA.n278 GNDA 0.016774f
C2735 VDDA.n279 GNDA 0.067923f
C2736 VDDA.n280 GNDA 0.016152f
C2737 VDDA.n281 GNDA 0.0656f
C2738 VDDA.n282 GNDA 0.105129f
C2739 VDDA.t366 GNDA 0.025053f
C2740 VDDA.t364 GNDA 0.016508f
C2741 VDDA.n283 GNDA 0.039301f
C2742 VDDA.n284 GNDA 0.055921f
C2743 VDDA.t420 GNDA 0.025053f
C2744 VDDA.t418 GNDA 0.016508f
C2745 VDDA.n285 GNDA 0.039301f
C2746 VDDA.n286 GNDA 0.055921f
C2747 VDDA.n287 GNDA 0.080028f
C2748 VDDA.n288 GNDA 0.105129f
C2749 VDDA.n289 GNDA 0.22858f
C2750 VDDA.t419 GNDA 0.208484f
C2751 VDDA.t77 GNDA 0.132047f
C2752 VDDA.t458 GNDA 0.132047f
C2753 VDDA.t32 GNDA 0.132047f
C2754 VDDA.t2 GNDA 0.132047f
C2755 VDDA.t149 GNDA 0.132047f
C2756 VDDA.t34 GNDA 0.132047f
C2757 VDDA.t79 GNDA 0.132047f
C2758 VDDA.t105 GNDA 0.132047f
C2759 VDDA.t60 GNDA 0.099035f
C2760 VDDA.n290 GNDA 0.066023f
C2761 VDDA.t454 GNDA 0.099035f
C2762 VDDA.t151 GNDA 0.132047f
C2763 VDDA.t120 GNDA 0.132047f
C2764 VDDA.t218 GNDA 0.132047f
C2765 VDDA.t122 GNDA 0.132047f
C2766 VDDA.t68 GNDA 0.132047f
C2767 VDDA.t456 GNDA 0.132047f
C2768 VDDA.t66 GNDA 0.132047f
C2769 VDDA.t212 GNDA 0.132047f
C2770 VDDA.t365 GNDA 0.208484f
C2771 VDDA.n291 GNDA 0.22858f
C2772 VDDA.n292 GNDA 0.0656f
C2773 VDDA.n293 GNDA 0.111752f
C2774 VDDA.n294 GNDA 0.047203f
C2775 VDDA.n295 GNDA 0.021341f
C2776 VDDA.n296 GNDA 0.016774f
C2777 VDDA.n297 GNDA 0.067923f
C2778 VDDA.n298 GNDA 0.016774f
C2779 VDDA.n299 GNDA 0.067923f
C2780 VDDA.n300 GNDA 0.016774f
C2781 VDDA.n301 GNDA 0.067923f
C2782 VDDA.n302 GNDA 0.016774f
C2783 VDDA.n303 GNDA 0.097267f
C2784 VDDA.n304 GNDA 0.021341f
C2785 VDDA.n305 GNDA 0.016152f
C2786 VDDA.n306 GNDA 0.016152f
C2787 VDDA.n307 GNDA 0.047203f
C2788 VDDA.n308 GNDA 0.021341f
C2789 VDDA.n309 GNDA 0.016152f
C2790 VDDA.n310 GNDA 0.021341f
C2791 VDDA.n311 GNDA 0.016152f
C2792 VDDA.n312 GNDA 0.047203f
C2793 VDDA.n313 GNDA 0.021341f
C2794 VDDA.n314 GNDA 0.021341f
C2795 VDDA.n315 GNDA 0.047203f
C2796 VDDA.n316 GNDA 0.021341f
C2797 VDDA.n317 GNDA 0.021341f
C2798 VDDA.n318 GNDA 0.016152f
C2799 VDDA.n319 GNDA 0.047203f
C2800 VDDA.n320 GNDA 0.021341f
C2801 VDDA.n321 GNDA 0.021341f
C2802 VDDA.n322 GNDA 0.047203f
C2803 VDDA.n323 GNDA 0.021341f
C2804 VDDA.n324 GNDA 0.016152f
C2805 VDDA.n325 GNDA 0.047203f
C2806 VDDA.n326 GNDA 0.021341f
C2807 VDDA.n327 GNDA 0.050685f
C2808 VDDA.n328 GNDA 0.047203f
C2809 VDDA.n329 GNDA 0.034843f
C2810 VDDA.n330 GNDA 0.03328f
C2811 VDDA.n331 GNDA 0.22858f
C2812 VDDA.t316 GNDA 0.208484f
C2813 VDDA.t239 GNDA 0.132047f
C2814 VDDA.t53 GNDA 0.132047f
C2815 VDDA.t210 GNDA 0.132047f
C2816 VDDA.t220 GNDA 0.132047f
C2817 VDDA.t175 GNDA 0.132047f
C2818 VDDA.t426 GNDA 0.132047f
C2819 VDDA.t438 GNDA 0.132047f
C2820 VDDA.t19 GNDA 0.132047f
C2821 VDDA.t51 GNDA 0.099035f
C2822 VDDA.n332 GNDA 0.066023f
C2823 VDDA.t202 GNDA 0.099035f
C2824 VDDA.t36 GNDA 0.132047f
C2825 VDDA.t71 GNDA 0.132047f
C2826 VDDA.t440 GNDA 0.132047f
C2827 VDDA.t208 GNDA 0.132047f
C2828 VDDA.t17 GNDA 0.132047f
C2829 VDDA.t114 GNDA 0.132047f
C2830 VDDA.t254 GNDA 0.132047f
C2831 VDDA.t4 GNDA 0.132047f
C2832 VDDA.t350 GNDA 0.208484f
C2833 VDDA.n333 GNDA 0.22858f
C2834 VDDA.n334 GNDA 0.03328f
C2835 VDDA.n335 GNDA 0.034843f
C2836 VDDA.n336 GNDA 0.047203f
C2837 VDDA.n337 GNDA 0.064608f
C2838 VDDA.n338 GNDA 0.196152f
C2839 VDDA.t284 GNDA 0.020007f
C2840 VDDA.t282 GNDA 0.020007f
C2841 VDDA.n339 GNDA 0.066097f
C2842 VDDA.n340 GNDA 0.08529f
C2843 VDDA.t402 GNDA 0.061313f
C2844 VDDA.n341 GNDA 0.108038f
C2845 VDDA.n342 GNDA 0.147277f
C2846 VDDA.n343 GNDA 0.147277f
C2847 VDDA.n344 GNDA 0.1466f
C2848 VDDA.t345 GNDA 0.061313f
C2849 VDDA.t343 GNDA 0.095402f
C2850 VDDA.t387 GNDA 0.025053f
C2851 VDDA.t385 GNDA 0.012643f
C2852 VDDA.n345 GNDA 0.039499f
C2853 VDDA.n346 GNDA 0.022776f
C2854 VDDA.n347 GNDA 0.040478f
C2855 VDDA.t408 GNDA 0.025053f
C2856 VDDA.t406 GNDA 0.012643f
C2857 VDDA.n348 GNDA 0.039499f
C2858 VDDA.n349 GNDA 0.040478f
C2859 VDDA.n350 GNDA 0.040478f
C2860 VDDA.n351 GNDA 0.033213f
C2861 VDDA.n352 GNDA 0.159598f
C2862 VDDA.t386 GNDA 0.2004f
C2863 VDDA.t207 GNDA 0.090782f
C2864 VDDA.n353 GNDA 0.060521f
C2865 VDDA.t206 GNDA 0.090782f
C2866 VDDA.t407 GNDA 0.203355f
C2867 VDDA.n354 GNDA 0.167647f
C2868 VDDA.n355 GNDA 0.033213f
C2869 VDDA.n356 GNDA 0.022776f
C2870 VDDA.n357 GNDA 0.031997f
C2871 VDDA.t303 GNDA 0.020007f
C2872 VDDA.t264 GNDA 0.020007f
C2873 VDDA.n358 GNDA 0.066097f
C2874 VDDA.n359 GNDA 0.08529f
C2875 VDDA.t275 GNDA 0.020007f
C2876 VDDA.t294 GNDA 0.020007f
C2877 VDDA.n360 GNDA 0.066097f
C2878 VDDA.n361 GNDA 0.08529f
C2879 VDDA.t259 GNDA 0.020007f
C2880 VDDA.t278 GNDA 0.020007f
C2881 VDDA.n362 GNDA 0.066097f
C2882 VDDA.n363 GNDA 0.08529f
C2883 VDDA.t292 GNDA 0.020007f
C2884 VDDA.t300 GNDA 0.020007f
C2885 VDDA.n364 GNDA 0.066097f
C2886 VDDA.n365 GNDA 0.08529f
C2887 VDDA.t273 GNDA 0.020007f
C2888 VDDA.t269 GNDA 0.020007f
C2889 VDDA.n366 GNDA 0.066097f
C2890 VDDA.n367 GNDA 0.08529f
C2891 VDDA.t298 GNDA 0.020007f
C2892 VDDA.t308 GNDA 0.020007f
C2893 VDDA.n368 GNDA 0.066097f
C2894 VDDA.n369 GNDA 0.08529f
C2895 VDDA.t266 GNDA 0.020007f
C2896 VDDA.t287 GNDA 0.020007f
C2897 VDDA.n370 GNDA 0.066097f
C2898 VDDA.n371 GNDA 0.08529f
C2899 VDDA.n372 GNDA 0.09417f
C2900 VDDA.n373 GNDA 0.113859f
C2901 VDDA.n374 GNDA 0.076747f
C2902 VDDA.n375 GNDA 0.093702f
C2903 VDDA.n376 GNDA 0.345246f
C2904 VDDA.t344 GNDA 0.445482f
C2905 VDDA.t265 GNDA 0.321114f
C2906 VDDA.t286 GNDA 0.321114f
C2907 VDDA.t297 GNDA 0.321114f
C2908 VDDA.t307 GNDA 0.321114f
C2909 VDDA.t272 GNDA 0.321114f
C2910 VDDA.t268 GNDA 0.321114f
C2911 VDDA.t291 GNDA 0.321114f
C2912 VDDA.t299 GNDA 0.240836f
C2913 VDDA.n377 GNDA 0.160557f
C2914 VDDA.t258 GNDA 0.240836f
C2915 VDDA.t277 GNDA 0.321114f
C2916 VDDA.t274 GNDA 0.321114f
C2917 VDDA.t293 GNDA 0.321114f
C2918 VDDA.t302 GNDA 0.321114f
C2919 VDDA.t263 GNDA 0.321114f
C2920 VDDA.t283 GNDA 0.321114f
C2921 VDDA.t281 GNDA 0.321114f
C2922 VDDA.t401 GNDA 0.445482f
C2923 VDDA.n378 GNDA 0.345246f
C2924 VDDA.n379 GNDA 0.093702f
C2925 VDDA.n380 GNDA 0.076747f
C2926 VDDA.t400 GNDA 0.095402f
C2927 VDDA.n381 GNDA 0.113859f
C2928 VDDA.n382 GNDA 0.052266f
C2929 VDDA.n383 GNDA 0.016107f
C2930 VDDA.t332 GNDA 0.025239f
C2931 VDDA.t330 GNDA 0.012316f
C2932 VDDA.n384 GNDA 0.037806f
C2933 VDDA.n385 GNDA 0.022671f
C2934 VDDA.n386 GNDA 0.040478f
C2935 VDDA.t329 GNDA 0.025239f
C2936 VDDA.t327 GNDA 0.012316f
C2937 VDDA.n387 GNDA 0.037806f
C2938 VDDA.n388 GNDA 0.040478f
C2939 VDDA.n389 GNDA 0.040478f
C2940 VDDA.n390 GNDA 0.033213f
C2941 VDDA.n391 GNDA 0.159598f
C2942 VDDA.t331 GNDA 0.2004f
C2943 VDDA.t0 GNDA 0.090782f
C2944 VDDA.n392 GNDA 0.060521f
C2945 VDDA.t177 GNDA 0.090782f
C2946 VDDA.t328 GNDA 0.2004f
C2947 VDDA.n393 GNDA 0.159598f
C2948 VDDA.n394 GNDA 0.033213f
C2949 VDDA.n395 GNDA 0.022671f
C2950 VDDA.n396 GNDA 0.023818f
C2951 VDDA.n397 GNDA 0.044582f
C2952 VDDA.n398 GNDA 0.093928f
C2953 VDDA.n399 GNDA 0.163104f
C2954 VDDA.n400 GNDA 0.016636f
C2955 VDDA.n401 GNDA 0.058724f
C2956 VDDA.t335 GNDA 0.02632f
C2957 VDDA.n402 GNDA 0.022008f
C2958 VDDA.n403 GNDA 0.047636f
C2959 VDDA.n404 GNDA 0.047636f
C2960 VDDA.n405 GNDA 0.047636f
C2961 VDDA.t396 GNDA 0.02632f
C2962 VDDA.t394 GNDA 0.013134f
C2963 VDDA.n406 GNDA 0.016605f
C2964 VDDA.n407 GNDA 0.058755f
C2965 VDDA.t411 GNDA 0.025117f
C2966 VDDA.n408 GNDA 0.044016f
C2967 VDDA.n409 GNDA 0.069346f
C2968 VDDA.n410 GNDA 0.069346f
C2969 VDDA.n411 GNDA 0.069346f
C2970 VDDA.t417 GNDA 0.025117f
C2971 VDDA.t415 GNDA 0.013134f
C2972 VDDA.n412 GNDA 0.016643f
C2973 VDDA.n413 GNDA 0.058717f
C2974 VDDA.t378 GNDA 0.02633f
C2975 VDDA.n414 GNDA 0.022008f
C2976 VDDA.n415 GNDA 0.047636f
C2977 VDDA.n416 GNDA 0.047636f
C2978 VDDA.n417 GNDA 0.047636f
C2979 VDDA.t311 GNDA 0.02633f
C2980 VDDA.t309 GNDA 0.013134f
C2981 VDDA.n418 GNDA 0.016643f
C2982 VDDA.n419 GNDA 0.080365f
C2983 VDDA.n420 GNDA 0.045093f
C2984 VDDA.n421 GNDA 0.026911f
C2985 VDDA.n422 GNDA 0.036969f
C2986 VDDA.n423 GNDA 0.168422f
C2987 VDDA.t310 GNDA 0.203924f
C2988 VDDA.t94 GNDA 0.122877f
C2989 VDDA.t38 GNDA 0.092158f
C2990 VDDA.n424 GNDA 0.061439f
C2991 VDDA.t434 GNDA 0.092158f
C2992 VDDA.t182 GNDA 0.122877f
C2993 VDDA.t377 GNDA 0.203924f
C2994 VDDA.n425 GNDA 0.168422f
C2995 VDDA.n426 GNDA 0.036969f
C2996 VDDA.n427 GNDA 0.026911f
C2997 VDDA.t376 GNDA 0.01355f
C2998 VDDA.n428 GNDA 0.044628f
C2999 VDDA.n429 GNDA 0.040536f
C3000 VDDA.n430 GNDA 0.016605f
C3001 VDDA.n431 GNDA 0.058755f
C3002 VDDA.n432 GNDA 0.016605f
C3003 VDDA.n433 GNDA 0.058755f
C3004 VDDA.n434 GNDA 0.016605f
C3005 VDDA.n435 GNDA 0.058755f
C3006 VDDA.n436 GNDA 0.016605f
C3007 VDDA.n437 GNDA 0.058755f
C3008 VDDA.n438 GNDA 0.040536f
C3009 VDDA.n439 GNDA 0.045424f
C3010 VDDA.n440 GNDA 0.041582f
C3011 VDDA.n441 GNDA 0.051825f
C3012 VDDA.n442 GNDA 0.198134f
C3013 VDDA.t416 GNDA 0.203924f
C3014 VDDA.t200 GNDA 0.122877f
C3015 VDDA.t444 GNDA 0.122877f
C3016 VDDA.t452 GNDA 0.122877f
C3017 VDDA.t40 GNDA 0.122877f
C3018 VDDA.t460 GNDA 0.122877f
C3019 VDDA.t137 GNDA 0.092158f
C3020 VDDA.n443 GNDA 0.061439f
C3021 VDDA.t198 GNDA 0.092158f
C3022 VDDA.t196 GNDA 0.122877f
C3023 VDDA.t147 GNDA 0.122877f
C3024 VDDA.t436 GNDA 0.122877f
C3025 VDDA.t410 GNDA 0.203924f
C3026 VDDA.n444 GNDA 0.183322f
C3027 VDDA.n445 GNDA 0.044419f
C3028 VDDA.n446 GNDA 0.034246f
C3029 VDDA.t409 GNDA 0.013134f
C3030 VDDA.n447 GNDA 0.045424f
C3031 VDDA.n448 GNDA 0.047872f
C3032 VDDA.n449 GNDA 0.016636f
C3033 VDDA.n450 GNDA 0.058724f
C3034 VDDA.n451 GNDA 0.047872f
C3035 VDDA.n452 GNDA 0.044221f
C3036 VDDA.n453 GNDA 0.026911f
C3037 VDDA.n454 GNDA 0.036459f
C3038 VDDA.n455 GNDA 0.166601f
C3039 VDDA.t395 GNDA 0.2004f
C3040 VDDA.t163 GNDA 0.121043f
C3041 VDDA.t229 GNDA 0.082529f
C3042 VDDA.n456 GNDA 0.030261f
C3043 VDDA.n457 GNDA 0.038514f
C3044 VDDA.t227 GNDA 0.090782f
C3045 VDDA.t442 GNDA 0.121043f
C3046 VDDA.t334 GNDA 0.2004f
C3047 VDDA.n458 GNDA 0.167622f
C3048 VDDA.n459 GNDA 0.03748f
C3049 VDDA.n460 GNDA 0.026911f
C3050 VDDA.t333 GNDA 0.013134f
C3051 VDDA.n461 GNDA 0.044221f
C3052 VDDA.n462 GNDA 0.088202f
C3053 VDDA.n463 GNDA 0.132398f
C3054 VDDA.t296 GNDA 0.372799f
C3055 VDDA.t304 GNDA 0.37415f
C3056 VDDA.t276 GNDA 0.372799f
C3057 VDDA.t260 GNDA 0.37415f
C3058 VDDA.t285 GNDA 0.372799f
C3059 VDDA.t289 GNDA 0.37415f
C3060 VDDA.t261 GNDA 0.372799f
C3061 VDDA.t301 GNDA 0.37415f
C3062 VDDA.t290 GNDA 0.372799f
C3063 VDDA.t306 GNDA 0.37415f
C3064 VDDA.t279 GNDA 0.372799f
C3065 VDDA.t262 GNDA 0.37415f
C3066 VDDA.t257 GNDA 0.372799f
C3067 VDDA.t271 GNDA 0.37415f
C3068 VDDA.t295 GNDA 0.372799f
C3069 VDDA.t280 GNDA 0.37415f
C3070 VDDA.n464 GNDA 0.249888f
C3071 VDDA.t288 GNDA 0.198999f
C3072 VDDA.n465 GNDA 0.271134f
C3073 VDDA.t270 GNDA 0.198999f
C3074 VDDA.n466 GNDA 0.271134f
C3075 VDDA.t305 GNDA 0.198999f
C3076 VDDA.n467 GNDA 0.271134f
C3077 VDDA.t267 GNDA 0.296946f
C3078 VDDA.n468 GNDA 0.258751f
C3079 VDDA.n469 GNDA 0.804137f
C3080 bgr_0.Vin-.n0 GNDA 0.073641f
C3081 bgr_0.Vin-.n1 GNDA 0.082742f
C3082 bgr_0.Vin-.n2 GNDA 0.998979f
C3083 bgr_0.Vin-.t5 GNDA 0.028614f
C3084 bgr_0.Vin-.t7 GNDA 0.028614f
C3085 bgr_0.Vin-.n3 GNDA 0.099613f
C3086 bgr_0.Vin-.t4 GNDA 0.028614f
C3087 bgr_0.Vin-.t6 GNDA 0.028614f
C3088 bgr_0.Vin-.n4 GNDA 0.095121f
C3089 bgr_0.Vin-.n5 GNDA 0.408067f
C3090 bgr_0.Vin-.t1 GNDA 0.098662f
C3091 bgr_0.Vin-.n6 GNDA 0.025702f
C3092 bgr_0.Vin-.n7 GNDA 0.469862f
C3093 bgr_0.Vin-.n8 GNDA 0.222852f
C3094 bgr_0.Vin-.t10 GNDA 0.023594f
C3095 bgr_0.Vin-.n9 GNDA 0.027673f
C3096 bgr_0.Vin-.n10 GNDA 0.022653f
C3097 bgr_0.Vin-.n11 GNDA 0.022653f
C3098 bgr_0.Vin-.n12 GNDA 0.040466f
C3099 bgr_0.Vin-.n13 GNDA 0.524007f
C3100 bgr_0.Vin-.t0 GNDA 0.276208f
C3101 bgr_0.Vin-.n14 GNDA 0.510829f
C3102 bgr_0.Vin-.n15 GNDA 0.074468f
C3103 bgr_0.Vin-.n16 GNDA 0.126176f
C3104 bgr_0.Vin-.n17 GNDA 0.073776f
C3105 bgr_0.Vin-.n18 GNDA 0.145931f
C3106 bgr_0.Vin-.n19 GNDA 0.145931f
C3107 bgr_0.Vin-.n20 GNDA -5.06787f
C3108 bgr_0.Vin-.n21 GNDA 5.25363f
C3109 bgr_0.Vin-.n22 GNDA 0.222489f
C3110 bgr_0.Vin-.n23 GNDA 0.382836f
C3111 bgr_0.Vin-.n24 GNDA 0.166915f
C3112 bgr_0.Vin-.n25 GNDA 0.040544f
C3113 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.043026f
C3114 bgr_0.V_TOP.t31 GNDA 0.115045f
C3115 bgr_0.V_TOP.t44 GNDA 0.115045f
C3116 bgr_0.V_TOP.t18 GNDA 0.115045f
C3117 bgr_0.V_TOP.t26 GNDA 0.115045f
C3118 bgr_0.V_TOP.t37 GNDA 0.115045f
C3119 bgr_0.V_TOP.t35 GNDA 0.115045f
C3120 bgr_0.V_TOP.t48 GNDA 0.115045f
C3121 bgr_0.V_TOP.t20 GNDA 0.115045f
C3122 bgr_0.V_TOP.t27 GNDA 0.115045f
C3123 bgr_0.V_TOP.t41 GNDA 0.115045f
C3124 bgr_0.V_TOP.t38 GNDA 0.115045f
C3125 bgr_0.V_TOP.t14 GNDA 0.115045f
C3126 bgr_0.V_TOP.t23 GNDA 0.115045f
C3127 bgr_0.V_TOP.t29 GNDA 0.115045f
C3128 bgr_0.V_TOP.t43 GNDA 0.150392f
C3129 bgr_0.V_TOP.n0 GNDA 0.084081f
C3130 bgr_0.V_TOP.n1 GNDA 0.061357f
C3131 bgr_0.V_TOP.n2 GNDA 0.061357f
C3132 bgr_0.V_TOP.n3 GNDA 0.061357f
C3133 bgr_0.V_TOP.n4 GNDA 0.061357f
C3134 bgr_0.V_TOP.n5 GNDA 0.057217f
C3135 bgr_0.V_TOP.t12 GNDA 0.147947f
C3136 bgr_0.V_TOP.t13 GNDA 0.155772f
C3137 bgr_0.V_TOP.t5 GNDA 0.010957f
C3138 bgr_0.V_TOP.t1 GNDA 0.010957f
C3139 bgr_0.V_TOP.n6 GNDA 0.027281f
C3140 bgr_0.V_TOP.n7 GNDA 0.726844f
C3141 bgr_0.V_TOP.t0 GNDA 0.010957f
C3142 bgr_0.V_TOP.t2 GNDA 0.010957f
C3143 bgr_0.V_TOP.n8 GNDA 0.026425f
C3144 bgr_0.V_TOP.t6 GNDA 0.010957f
C3145 bgr_0.V_TOP.t8 GNDA 0.010957f
C3146 bgr_0.V_TOP.n9 GNDA 0.027465f
C3147 bgr_0.V_TOP.t7 GNDA 0.010957f
C3148 bgr_0.V_TOP.t3 GNDA 0.010957f
C3149 bgr_0.V_TOP.n10 GNDA 0.027281f
C3150 bgr_0.V_TOP.n11 GNDA 0.252824f
C3151 bgr_0.V_TOP.n12 GNDA 0.153577f
C3152 bgr_0.V_TOP.n13 GNDA 0.087653f
C3153 bgr_0.V_TOP.t4 GNDA 0.010957f
C3154 bgr_0.V_TOP.t10 GNDA 0.010957f
C3155 bgr_0.V_TOP.n14 GNDA 0.027281f
C3156 bgr_0.V_TOP.n15 GNDA 0.151313f
C3157 bgr_0.V_TOP.t9 GNDA 0.010957f
C3158 bgr_0.V_TOP.t11 GNDA 0.010957f
C3159 bgr_0.V_TOP.n16 GNDA 0.027281f
C3160 bgr_0.V_TOP.n17 GNDA 0.149874f
C3161 bgr_0.V_TOP.n18 GNDA 0.329448f
C3162 bgr_0.V_TOP.n19 GNDA 0.023183f
C3163 bgr_0.V_TOP.n20 GNDA 0.057217f
C3164 bgr_0.V_TOP.n21 GNDA 0.061357f
C3165 bgr_0.V_TOP.n22 GNDA 0.061357f
C3166 bgr_0.V_TOP.n23 GNDA 0.061357f
C3167 bgr_0.V_TOP.n24 GNDA 0.061357f
C3168 bgr_0.V_TOP.n25 GNDA 0.061357f
C3169 bgr_0.V_TOP.n26 GNDA 0.061357f
C3170 bgr_0.V_TOP.n27 GNDA 0.057217f
C3171 bgr_0.V_TOP.t32 GNDA 0.132572f
C3172 bgr_0.V_TOP.t49 GNDA 0.445732f
C3173 bgr_0.V_TOP.t39 GNDA 0.438267f
C3174 bgr_0.V_TOP.n28 GNDA 0.293844f
C3175 bgr_0.V_TOP.t28 GNDA 0.438267f
C3176 bgr_0.V_TOP.t25 GNDA 0.445732f
C3177 bgr_0.V_TOP.t33 GNDA 0.438267f
C3178 bgr_0.V_TOP.n29 GNDA 0.293844f
C3179 bgr_0.V_TOP.n30 GNDA 0.273917f
C3180 bgr_0.V_TOP.t21 GNDA 0.445732f
C3181 bgr_0.V_TOP.t15 GNDA 0.438267f
C3182 bgr_0.V_TOP.n31 GNDA 0.293844f
C3183 bgr_0.V_TOP.t40 GNDA 0.438267f
C3184 bgr_0.V_TOP.t34 GNDA 0.445732f
C3185 bgr_0.V_TOP.t45 GNDA 0.438267f
C3186 bgr_0.V_TOP.n32 GNDA 0.293844f
C3187 bgr_0.V_TOP.n33 GNDA 0.356092f
C3188 bgr_0.V_TOP.t30 GNDA 0.445732f
C3189 bgr_0.V_TOP.t22 GNDA 0.438267f
C3190 bgr_0.V_TOP.n34 GNDA 0.293844f
C3191 bgr_0.V_TOP.t16 GNDA 0.438267f
C3192 bgr_0.V_TOP.t46 GNDA 0.445732f
C3193 bgr_0.V_TOP.t19 GNDA 0.438267f
C3194 bgr_0.V_TOP.n35 GNDA 0.293844f
C3195 bgr_0.V_TOP.n36 GNDA 0.356092f
C3196 bgr_0.V_TOP.t24 GNDA 0.445732f
C3197 bgr_0.V_TOP.t17 GNDA 0.438267f
C3198 bgr_0.V_TOP.n37 GNDA 0.293844f
C3199 bgr_0.V_TOP.t42 GNDA 0.438267f
C3200 bgr_0.V_TOP.n38 GNDA 0.273917f
C3201 bgr_0.V_TOP.t47 GNDA 0.438267f
C3202 bgr_0.V_TOP.n39 GNDA 0.191742f
C3203 bgr_0.V_TOP.t36 GNDA 0.438267f
C3204 bgr_0.V_TOP.n40 GNDA 0.893239f
.ends

