* PEX produced on Tue Aug 26 07:38:37 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr.ext - technology: sky130A

.subckt bgr VDDA CURRENT_OUTPUT GNDA
X0 V_CUR_REF_REG.t12 V2.t10 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X1 1st_Vout_1.t7 cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 CURRENT_OUTPUT.t11 V2.t11 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X3 Vin+.t5 V_TOP.t14 VDDA.t25 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X4 GNDA.t26 START_UP_NFET1.t0 START_UP_NFET1.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X5 1st_Vout_2.t6 a_36200_n1130.t13 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X6 1st_Vout_1.t5 V_mir1.t13 VDDA.t95 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X7 1st_Vout_2.t7 cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 V_CUR_REF_REG.t0 GNDA.t1 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1
X9 1st_Vout_2.t8 cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 1st_Vout_2.t9 cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 VDDA.t69 V_TOP.t15 Vin-.t7 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X12 VDDA.t201 1st_Vout_1.t8 V_TOP.t13 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X13 Vin-.t2 START_UP.t6 V_TOP.t1 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X14 V2.t6 VDDA.t129 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X15 1st_Vout_2.t10 cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 1st_Vout_2.t11 cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 V_CUR_REF_REG.t11 V2.t12 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X18 1st_Vout_1.t9 cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VDDA.t40 V_mir1.t14 1st_Vout_1.t3 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X20 1st_Vout_2.t12 cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 CURRENT_OUTPUT.t10 V2.t13 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X22 V1.t6 V_TOP.t16 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X23 V_TOP.t6 VDDA.t126 VDDA.t128 VDDA.t127 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X24 1st_Vout_2.t13 cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 1st_Vout_1.t10 cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 VDDA.t191 V2.t14 V_CUR_REF_REG.t10 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X27 1st_Vout_1.t11 cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 V_TOP.t17 VDDA.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 VDDA.t125 VDDA.t123 V2.t7 VDDA.t124 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X30 1st_Vout_1.t12 cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 VDDA.t189 V2.t15 CURRENT_OUTPUT.t9 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X32 1st_Vout_2.t5 a_36200_n1130.t14 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X33 1st_Vout_1.t13 cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 V_TOP.t18 VDDA.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 V_CUR_REF_REG.t9 V2.t16 VDDA.t187 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X36 VDDA.t122 VDDA.t120 V_TOP.t5 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X37 V_TOP.t19 VDDA.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 1st_Vout_2.t14 cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 V_TOP.t20 VDDA.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 VDDA.t36 a_36200_n1130.t11 a_36200_n1130.t12 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X41 CURRENT_OUTPUT.t1 VDDA.t117 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X42 a_38370_n6700.t0 a_38490_n7778.t1 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X43 V_p_2.t1 VDDA.t202 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X44 VDDA.t185 V2.t17 V_CUR_REF_REG.t8 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X45 VDDA.t138 a_36200_n1130.t15 1st_Vout_2.t4 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X46 VDDA.t23 V_mir1.t15 1st_Vout_1.t1 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X47 VDDA.t15 V_mir1.t11 V_mir1.t12 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X48 VDDA.t150 V_mir1.t9 V_mir1.t10 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X49 VDDA.t46 a_36200_n1130.t9 a_36200_n1130.t10 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 VDDA.t66 1st_Vout_1.t14 V_TOP.t12 VDDA.t65 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X51 VDDA.t116 VDDA.t114 CURRENT_OUTPUT.t0 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X52 1st_Vout_2.t15 cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 V_p_2.t2 V_CUR_REF_REG.t13 1st_Vout_2.t0 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X54 VDDA.t11 a_36200_n1130.t16 1st_Vout_2.t3 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X55 1st_Vout_2.t16 cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 Vin+.t1 a_38040_n7928.t0 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=6
X57 V_TOP.t2 cap_res1.t0 GNDA.t13 sky130_fd_pr__res_high_po_0p35 l=2.05
X58 1st_Vout_2.t17 cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 1st_Vout_2.t18 cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 VDDA.t82 1st_Vout_2.t19 V2.t4 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X61 V1.t2 VDDA.t111 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X62 VDDA.t17 V_mir1.t7 V_mir1.t8 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X63 V_p_1.t0 Vin-.t8 V_mir1.t0 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X64 VDDA.t110 VDDA.t108 V_CUR_REF_REG.t2 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X65 1st_Vout_2.t20 cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 1st_Vout_1.t15 cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 VDDA.t44 1st_Vout_2.t21 V2.t2 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X68 Vin+.t0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 GNDA.t10 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X69 1st_Vout_1.t16 cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VDDA.t183 V2.t18 CURRENT_OUTPUT.t8 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X71 1st_Vout_2.t22 cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 V_TOP.t11 1st_Vout_1.t17 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X73 1st_Vout_1.t18 cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 V_TOP.t21 VDDA.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VDDA.t74 V_TOP.t22 Vin+.t4 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X76 VDDA.t60 a_36200_n1130.t7 a_36200_n1130.t8 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X77 V_TOP.t23 VDDA.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 VDDA.t133 1st_Vout_1.t19 V_TOP.t10 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 1st_Vout_1.t20 cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 V_TOP.t24 VDDA.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 V_TOP.t25 VDDA.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 1st_Vout_2.t23 cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 Vin+.t3 V_TOP.t26 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X84 VDDA.t38 V_mir1.t16 1st_Vout_1.t2 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X85 V_TOP.t27 VDDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 VDDA.t181 V2.t19 CURRENT_OUTPUT.t7 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X87 GNDA.t32 VDDA.t203 V2.t5 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X88 VDDA.t152 V_TOP.t28 V1.t5 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X89 V_TOP.t7 VDDA.t204 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X90 GNDA.t16 GNDA.t15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X91 V_TOP.t0 START_UP.t7 Vin-.t1 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X92 V_TOP.t29 VDDA.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 Vin-.t0 a_32970_n7928.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=6
X94 GNDA.t16 GNDA.t21 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X95 VDDA.t179 V2.t20 V_CUR_REF_REG.t7 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X96 VDDA.t107 VDDA.t105 V1.t1 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X97 GNDA.t16 GNDA.t20 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X98 VDDA.t177 V2.t21 CURRENT_OUTPUT.t6 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X99 VDDA.t48 a_36200_n1130.t17 1st_Vout_2.t2 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X100 V_TOP.t30 VDDA.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 Vin-.t6 V_TOP.t31 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X102 a_33090_n6320.t0 GNDA.t7 GNDA.t6 sky130_fd_pr__res_xhigh_po_0p35 l=6
X103 V_TOP.t32 VDDA.t153 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VDDA.t52 1st_Vout_2.t24 V2.t3 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X105 CURRENT_OUTPUT.t5 V2.t22 VDDA.t175 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X106 V_TOP.t33 VDDA.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 1st_Vout_2.t25 cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 a_37920_n6320.t0 GNDA.t12 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=6
X109 VDDA.t173 V2.t23 V_CUR_REF_REG.t6 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X110 VDDA.t136 V_TOP.t34 Vin+.t2 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X111 V_TOP.t35 VDDA.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 a_36200_n1130.t6 a_36200_n1130.t5 VDDA.t157 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X113 V_TOP.t9 1st_Vout_1.t21 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X114 1st_Vout_1.t22 cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VDDA.t171 V2.t24 CURRENT_OUTPUT.t4 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X116 1st_Vout_2.t26 cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 V_CUR_REF_REG.t5 V2.t25 VDDA.t169 VDDA.t168 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X118 1st_Vout_1.t23 cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 START_UP.t5 V_TOP.t36 VDDA.t42 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X120 1st_Vout_1.t0 V_mir1.t17 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X121 V_TOP.t37 VDDA.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 START_UP_NFET1.t1 START_UP.t0 START_UP.t1 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X123 1st_Vout_1.t24 cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 GNDA.t28 VDDA.t205 V_p_1.t1 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X125 1st_Vout_1.t25 cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 V2.t8 1st_Vout_2.t27 VDDA.t146 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X127 VDDA.t167 V2.t26 V_CUR_REF_REG.t4 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X128 VDDA.t93 V_TOP.t38 Vin-.t5 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X129 V_mir1.t6 V_mir1.t5 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X130 1st_Vout_1.t26 cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 a_36200_n1130.t0 V1.t7 V_p_2.t0 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X132 V1.t4 V_TOP.t39 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X133 a_36200_n1130.t4 a_36200_n1130.t3 VDDA.t159 VDDA.t158 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X134 V2.t1 cap_res2.t0 GNDA.t5 sky130_fd_pr__res_high_po_0p35 l=2.05
X135 a_38370_n6700.t1 GNDA.t9 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X136 1st_Vout_2.t1 a_36200_n1130.t18 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X137 V_TOP.t40 VDDA.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 1st_Vout_1.t6 Vin+.t6 V_p_1.t2 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X139 GNDA.t16 GNDA.t19 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X140 1st_Vout_1.t4 V_mir1.t18 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X141 GNDA.t16 GNDA.t18 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X142 VDDA.t86 V_TOP.t41 START_UP.t4 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X143 V_mir1.t4 V_mir1.t3 VDDA.t140 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X144 a_33090_n6320.t1 a_32970_n7928.t1 GNDA.t14 sky130_fd_pr__res_xhigh_po_0p35 l=6
X145 GNDA.t16 GNDA.t24 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X146 V2.t9 1st_Vout_2.t28 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X147 START_UP.t3 V_TOP.t42 VDDA.t64 VDDA.t63 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X148 V_mir1.t2 V_mir1.t1 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X149 CURRENT_OUTPUT.t3 V2.t27 VDDA.t165 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X150 V_TOP.t43 VDDA.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 1st_Vout_1.t27 cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 V_TOP.t4 VDDA.t102 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X153 V_TOP.t8 1st_Vout_1.t28 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X154 V_TOP.t44 VDDA.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VDDA.t9 V_TOP.t45 V1.t3 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X156 V_TOP.t46 VDDA.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 1st_Vout_2.t29 cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 1st_Vout_2.t30 cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 V_CUR_REF_REG.t1 VDDA.t99 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X160 V_CUR_REF_REG.t3 V2.t28 VDDA.t163 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X161 V_TOP.t47 VDDA.t144 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 GNDA.t16 GNDA.t17 Vin-.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X163 Vin-.t4 V_TOP.t48 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X164 1st_Vout_2.t31 cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 1st_Vout_1.t29 cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 a_37920_n6320.t1 a_38040_n7928.t1 GNDA.t11 sky130_fd_pr__res_xhigh_po_0p35 l=6
X167 GNDA.t16 GNDA.t23 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X168 CURRENT_OUTPUT.t2 V2.t29 VDDA.t161 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X169 V2.t0 1st_Vout_2.t32 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 1st_Vout_1.t30 cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 V1.t0 a_38490_n7778.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=3.35
X172 VDDA.t98 VDDA.t96 V_TOP.t3 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.2 ps=1.4 w=1 l=0.15
X173 1st_Vout_1.t31 cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 GNDA.t16 GNDA.t22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X175 VDDA.t80 V_TOP.t49 START_UP.t2 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X176 1st_Vout_1.t32 cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 a_36200_n1130.t2 a_36200_n1130.t1 VDDA.t84 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 V2.n0 V2.t24 403.952
R1 V2.n0 V2.t13 403.755
R2 V2.n1 V2.t21 403.755
R3 V2.n2 V2.t11 403.755
R4 V2.n3 V2.t19 403.755
R5 V2.n4 V2.t29 403.755
R6 V2.n5 V2.t15 403.755
R7 V2.n6 V2.t22 403.755
R8 V2.n7 V2.t18 403.755
R9 V2.n8 V2.t27 403.755
R10 V2.n9 V2.t26 403.755
R11 V2.n10 V2.t16 403.755
R12 V2.n11 V2.t23 403.755
R13 V2.n12 V2.t12 403.755
R14 V2.n13 V2.t20 403.755
R15 V2.n14 V2.t10 403.755
R16 V2.n15 V2.t17 403.755
R17 V2.n16 V2.t25 403.755
R18 V2.n17 V2.t14 403.755
R19 V2.n18 V2.t28 403.755
R20 V2.n20 V2.n19 301.933
R21 V2.n22 V2.n21 301.933
R22 V2.n24 V2.n23 301.933
R23 V2.n26 V2.n25 301.933
R24 V2.t1 V2.n27 117.322
R25 V2.n20 V2.t5 104.245
R26 V2.n19 V2.t2 39.4005
R27 V2.n19 V2.t6 39.4005
R28 V2.n21 V2.t3 39.4005
R29 V2.n21 V2.t9 39.4005
R30 V2.n23 V2.t4 39.4005
R31 V2.n23 V2.t0 39.4005
R32 V2.n25 V2.t7 39.4005
R33 V2.n25 V2.t8 39.4005
R34 V2.n27 V2.n18 10.78
R35 V2.n27 V2.n26 5.70362
R36 V2.n9 V2.n8 1.6255
R37 V2.n26 V2.n24 1.1255
R38 V2.n24 V2.n22 1.1255
R39 V2.n22 V2.n20 1.1255
R40 V2.n18 V2.n17 0.196929
R41 V2.n17 V2.n16 0.196929
R42 V2.n16 V2.n15 0.196929
R43 V2.n15 V2.n14 0.196929
R44 V2.n14 V2.n13 0.196929
R45 V2.n13 V2.n12 0.196929
R46 V2.n12 V2.n11 0.196929
R47 V2.n11 V2.n10 0.196929
R48 V2.n10 V2.n9 0.196929
R49 V2.n8 V2.n7 0.196929
R50 V2.n7 V2.n6 0.196929
R51 V2.n6 V2.n5 0.196929
R52 V2.n5 V2.n4 0.196929
R53 V2.n4 V2.n3 0.196929
R54 V2.n3 V2.n2 0.196929
R55 V2.n2 V2.n1 0.196929
R56 V2.n1 V2.n0 0.196929
R57 VDDA.n47 VDDA.t116 708.125
R58 VDDA.t116 VDDA.n13 708.125
R59 VDDA.n29 VDDA.t110 708.125
R60 VDDA.t110 VDDA.n18 708.125
R61 VDDA.n126 VDDA.t104 708.125
R62 VDDA.t104 VDDA.n119 708.125
R63 VDDA.n188 VDDA.t122 708.125
R64 VDDA.t122 VDDA.n139 708.125
R65 VDDA.n191 VDDA.t128 708.125
R66 VDDA.t128 VDDA.n138 708.125
R67 VDDA.n162 VDDA.t125 708.125
R68 VDDA.t125 VDDA.n143 708.125
R69 VDDA.n165 VDDA.t131 708.125
R70 VDDA.t131 VDDA.n142 708.125
R71 VDDA.n123 VDDA.t98 694.444
R72 VDDA.t98 VDDA.n120 694.444
R73 VDDA.t97 VDDA.n124 674.87
R74 VDDA.t121 VDDA.n189 657.76
R75 VDDA.t124 VDDA.n163 657.76
R76 VDDA.t115 VDDA.n48 640.794
R77 VDDA.t109 VDDA.n30 640.794
R78 VDDA.n80 VDDA.n78 587.407
R79 VDDA.n84 VDDA.n81 587.407
R80 VDDA.n110 VDDA.n57 587.407
R81 VDDA.n109 VDDA.n108 587.407
R82 VDDA.n111 VDDA.n110 585
R83 VDDA.n109 VDDA.n102 585
R84 VDDA.n91 VDDA.n80 585
R85 VDDA.n88 VDDA.n81 585
R86 VDDA.n190 VDDA.t127 540.818
R87 VDDA.n164 VDDA.t130 540.818
R88 VDDA.n49 VDDA.t118 523.855
R89 VDDA.n31 VDDA.t100 523.855
R90 VDDA.n125 VDDA.t103 523.855
R91 VDDA.n121 VDDA.t96 422.384
R92 VDDA.n128 VDDA.t102 422.384
R93 VDDA.n45 VDDA.t114 418.368
R94 VDDA.n52 VDDA.t117 418.368
R95 VDDA.n27 VDDA.t108 418.368
R96 VDDA.n34 VDDA.t99 418.368
R97 VDDA.t1 VDDA.t121 407.144
R98 VDDA.t39 VDDA.t1 407.144
R99 VDDA.t12 VDDA.t39 407.144
R100 VDDA.t14 VDDA.t12 407.144
R101 VDDA.t139 VDDA.t14 407.144
R102 VDDA.t200 VDDA.t139 407.144
R103 VDDA.t88 VDDA.t200 407.144
R104 VDDA.t22 VDDA.t88 407.144
R105 VDDA.t71 VDDA.t22 407.144
R106 VDDA.t16 VDDA.t71 407.144
R107 VDDA.t29 VDDA.t16 407.144
R108 VDDA.t65 VDDA.t29 407.144
R109 VDDA.t55 VDDA.t65 407.144
R110 VDDA.t37 VDDA.t55 407.144
R111 VDDA.t94 VDDA.t37 407.144
R112 VDDA.t149 VDDA.t94 407.144
R113 VDDA.t31 VDDA.t149 407.144
R114 VDDA.t132 VDDA.t31 407.144
R115 VDDA.t127 VDDA.t132 407.144
R116 VDDA.t145 VDDA.t124 407.144
R117 VDDA.t45 VDDA.t145 407.144
R118 VDDA.t156 VDDA.t45 407.144
R119 VDDA.t137 VDDA.t156 407.144
R120 VDDA.t18 VDDA.t137 407.144
R121 VDDA.t81 VDDA.t18 407.144
R122 VDDA.t3 VDDA.t81 407.144
R123 VDDA.t35 VDDA.t3 407.144
R124 VDDA.t158 VDDA.t35 407.144
R125 VDDA.t10 VDDA.t158 407.144
R126 VDDA.t147 VDDA.t10 407.144
R127 VDDA.t51 VDDA.t147 407.144
R128 VDDA.t154 VDDA.t51 407.144
R129 VDDA.t59 VDDA.t154 407.144
R130 VDDA.t83 VDDA.t59 407.144
R131 VDDA.t47 VDDA.t83 407.144
R132 VDDA.t53 VDDA.t47 407.144
R133 VDDA.t43 VDDA.t53 407.144
R134 VDDA.t130 VDDA.t43 407.144
R135 VDDA.t164 VDDA.t115 373.214
R136 VDDA.t182 VDDA.t164 373.214
R137 VDDA.t174 VDDA.t182 373.214
R138 VDDA.t188 VDDA.t174 373.214
R139 VDDA.t160 VDDA.t188 373.214
R140 VDDA.t180 VDDA.t160 373.214
R141 VDDA.t196 VDDA.t180 373.214
R142 VDDA.t176 VDDA.t196 373.214
R143 VDDA.t192 VDDA.t176 373.214
R144 VDDA.t170 VDDA.t192 373.214
R145 VDDA.t118 VDDA.t170 373.214
R146 VDDA.t162 VDDA.t109 373.214
R147 VDDA.t190 VDDA.t162 373.214
R148 VDDA.t168 VDDA.t190 373.214
R149 VDDA.t184 VDDA.t168 373.214
R150 VDDA.t198 VDDA.t184 373.214
R151 VDDA.t178 VDDA.t198 373.214
R152 VDDA.t194 VDDA.t178 373.214
R153 VDDA.t172 VDDA.t194 373.214
R154 VDDA.t186 VDDA.t172 373.214
R155 VDDA.t166 VDDA.t186 373.214
R156 VDDA.t100 VDDA.t166 373.214
R157 VDDA.t33 VDDA.t97 373.214
R158 VDDA.t87 VDDA.t33 373.214
R159 VDDA.t103 VDDA.t87 373.214
R160 VDDA.n186 VDDA.t120 370.168
R161 VDDA.n193 VDDA.t126 370.168
R162 VDDA.n160 VDDA.t123 370.168
R163 VDDA.n167 VDDA.t129 370.168
R164 VDDA.n77 VDDA.t105 360.868
R165 VDDA.n116 VDDA.t111 360.868
R166 VDDA.n12 VDDA.t119 351.793
R167 VDDA.n17 VDDA.t101 351.793
R168 VDDA.n10 VDDA.n9 301.933
R169 VDDA.n37 VDDA.n36 301.933
R170 VDDA.n39 VDDA.n38 301.933
R171 VDDA.n41 VDDA.n40 301.933
R172 VDDA.n43 VDDA.n42 301.933
R173 VDDA.n15 VDDA.n14 301.933
R174 VDDA.n20 VDDA.n19 301.933
R175 VDDA.n22 VDDA.n21 301.933
R176 VDDA.n24 VDDA.n23 301.933
R177 VDDA.n26 VDDA.n25 301.933
R178 VDDA.n137 VDDA.n136 299.231
R179 VDDA.n170 VDDA.n169 299.231
R180 VDDA.n172 VDDA.n171 299.231
R181 VDDA.n174 VDDA.n173 299.231
R182 VDDA.n176 VDDA.n175 299.231
R183 VDDA.n178 VDDA.n177 299.231
R184 VDDA.n180 VDDA.n179 299.231
R185 VDDA.n182 VDDA.n181 299.231
R186 VDDA.n184 VDDA.n183 299.231
R187 VDDA.n141 VDDA.n140 299.231
R188 VDDA.n145 VDDA.n144 299.231
R189 VDDA.n147 VDDA.n146 299.231
R190 VDDA.n149 VDDA.n148 299.231
R191 VDDA.n151 VDDA.n150 299.231
R192 VDDA.n153 VDDA.n152 299.231
R193 VDDA.n155 VDDA.n154 299.231
R194 VDDA.n157 VDDA.n156 299.231
R195 VDDA.n159 VDDA.n158 299.231
R196 VDDA.t20 VDDA.t106 251.471
R197 VDDA.t79 VDDA.t20 251.471
R198 VDDA.t63 VDDA.t79 251.471
R199 VDDA.t92 VDDA.t63 251.471
R200 VDDA.t5 VDDA.t92 251.471
R201 VDDA.t73 VDDA.t5 251.471
R202 VDDA.t24 VDDA.t73 251.471
R203 VDDA.t8 VDDA.t24 251.471
R204 VDDA.t75 VDDA.t8 251.471
R205 VDDA.t135 VDDA.t75 251.471
R206 VDDA.t141 VDDA.t135 251.471
R207 VDDA.t68 VDDA.t141 251.471
R208 VDDA.t77 VDDA.t68 251.471
R209 VDDA.t85 VDDA.t77 251.471
R210 VDDA.t41 VDDA.t85 251.471
R211 VDDA.t151 VDDA.t41 251.471
R212 VDDA.t112 VDDA.t151 251.471
R213 VDDA.n50 VDDA.n49 238.367
R214 VDDA.n49 VDDA.n11 238.367
R215 VDDA.n32 VDDA.n31 238.367
R216 VDDA.n31 VDDA.n16 238.367
R217 VDDA.n115 VDDA.n114 238.367
R218 VDDA.n126 VDDA.n125 238.367
R219 VDDA.n125 VDDA.n119 238.367
R220 VDDA.n191 VDDA.n190 238.367
R221 VDDA.n190 VDDA.n138 238.367
R222 VDDA.n165 VDDA.n164 238.367
R223 VDDA.n164 VDDA.n142 238.367
R224 VDDA.t106 VDDA.n96 237.5
R225 VDDA.n113 VDDA.t112 237.5
R226 VDDA.n100 VDDA.n58 185
R227 VDDA.n112 VDDA.n111 185
R228 VDDA.n113 VDDA.n112 185
R229 VDDA.n102 VDDA.n99 185
R230 VDDA.n107 VDDA.n106 185
R231 VDDA.n103 VDDA.n98 185
R232 VDDA.n113 VDDA.n98 185
R233 VDDA.n95 VDDA.n94 185
R234 VDDA.n96 VDDA.n95 185
R235 VDDA.n92 VDDA.n62 185
R236 VDDA.n91 VDDA.n90 185
R237 VDDA.n89 VDDA.n88 185
R238 VDDA.n83 VDDA.n82 185
R239 VDDA.n85 VDDA.n61 185
R240 VDDA.n96 VDDA.n61 185
R241 VDDA.n112 VDDA.n58 150
R242 VDDA.n112 VDDA.n99 150
R243 VDDA.n106 VDDA.n98 150
R244 VDDA.n95 VDDA.n62 150
R245 VDDA.n90 VDDA.n89 150
R246 VDDA.n82 VDDA.n61 150
R247 VDDA.n76 VDDA.n75 141.712
R248 VDDA.n74 VDDA.n73 141.712
R249 VDDA.n72 VDDA.n71 141.712
R250 VDDA.n70 VDDA.n69 141.712
R251 VDDA.n68 VDDA.n67 141.712
R252 VDDA.n66 VDDA.n65 141.712
R253 VDDA.n64 VDDA.n63 141.712
R254 VDDA.n55 VDDA.n54 141.712
R255 VDDA.t107 VDDA.n80 123.126
R256 VDDA.n81 VDDA.t107 123.126
R257 VDDA.n110 VDDA.t113 123.126
R258 VDDA.t113 VDDA.n109 123.126
R259 VDDA.n114 VDDA.n113 65.8183
R260 VDDA.n113 VDDA.n97 65.8183
R261 VDDA.n96 VDDA.n59 65.8183
R262 VDDA.n96 VDDA.n60 65.8183
R263 VDDA.n201 VDDA.t203 58.8003
R264 VDDA.n202 VDDA.t204 58.8003
R265 VDDA.n99 VDDA.n97 53.3664
R266 VDDA.n114 VDDA.n58 53.3664
R267 VDDA.n106 VDDA.n97 53.3664
R268 VDDA.n62 VDDA.n59 53.3664
R269 VDDA.n89 VDDA.n60 53.3664
R270 VDDA.n90 VDDA.n59 53.3664
R271 VDDA.n82 VDDA.n60 53.3664
R272 VDDA.n201 VDDA.t202 49.164
R273 VDDA.n203 VDDA.t205 48.516
R274 VDDA.n9 VDDA.t193 39.4005
R275 VDDA.n9 VDDA.t171 39.4005
R276 VDDA.n36 VDDA.t197 39.4005
R277 VDDA.n36 VDDA.t177 39.4005
R278 VDDA.n38 VDDA.t161 39.4005
R279 VDDA.n38 VDDA.t181 39.4005
R280 VDDA.n40 VDDA.t175 39.4005
R281 VDDA.n40 VDDA.t189 39.4005
R282 VDDA.n42 VDDA.t165 39.4005
R283 VDDA.n42 VDDA.t183 39.4005
R284 VDDA.n14 VDDA.t187 39.4005
R285 VDDA.n14 VDDA.t167 39.4005
R286 VDDA.n19 VDDA.t195 39.4005
R287 VDDA.n19 VDDA.t173 39.4005
R288 VDDA.n21 VDDA.t199 39.4005
R289 VDDA.n21 VDDA.t179 39.4005
R290 VDDA.n23 VDDA.t169 39.4005
R291 VDDA.n23 VDDA.t185 39.4005
R292 VDDA.n25 VDDA.t163 39.4005
R293 VDDA.n25 VDDA.t191 39.4005
R294 VDDA.n136 VDDA.t32 39.4005
R295 VDDA.n136 VDDA.t133 39.4005
R296 VDDA.n169 VDDA.t95 39.4005
R297 VDDA.n169 VDDA.t150 39.4005
R298 VDDA.n171 VDDA.t56 39.4005
R299 VDDA.n171 VDDA.t38 39.4005
R300 VDDA.n173 VDDA.t30 39.4005
R301 VDDA.n173 VDDA.t66 39.4005
R302 VDDA.n175 VDDA.t72 39.4005
R303 VDDA.n175 VDDA.t17 39.4005
R304 VDDA.n177 VDDA.t89 39.4005
R305 VDDA.n177 VDDA.t23 39.4005
R306 VDDA.n179 VDDA.t140 39.4005
R307 VDDA.n179 VDDA.t201 39.4005
R308 VDDA.n181 VDDA.t13 39.4005
R309 VDDA.n181 VDDA.t15 39.4005
R310 VDDA.n183 VDDA.t2 39.4005
R311 VDDA.n183 VDDA.t40 39.4005
R312 VDDA.n140 VDDA.t54 39.4005
R313 VDDA.n140 VDDA.t44 39.4005
R314 VDDA.n144 VDDA.t84 39.4005
R315 VDDA.n144 VDDA.t48 39.4005
R316 VDDA.n146 VDDA.t155 39.4005
R317 VDDA.n146 VDDA.t60 39.4005
R318 VDDA.n148 VDDA.t148 39.4005
R319 VDDA.n148 VDDA.t52 39.4005
R320 VDDA.n150 VDDA.t159 39.4005
R321 VDDA.n150 VDDA.t11 39.4005
R322 VDDA.n152 VDDA.t4 39.4005
R323 VDDA.n152 VDDA.t36 39.4005
R324 VDDA.n154 VDDA.t19 39.4005
R325 VDDA.n154 VDDA.t82 39.4005
R326 VDDA.n156 VDDA.t157 39.4005
R327 VDDA.n156 VDDA.t138 39.4005
R328 VDDA.n158 VDDA.t146 39.4005
R329 VDDA.n158 VDDA.t46 39.4005
R330 VDDA.n116 VDDA.n115 22.8576
R331 VDDA.n94 VDDA.n77 22.8576
R332 VDDA.n54 VDDA.t42 13.1338
R333 VDDA.n54 VDDA.t152 13.1338
R334 VDDA.n63 VDDA.t78 13.1338
R335 VDDA.n63 VDDA.t86 13.1338
R336 VDDA.n65 VDDA.t142 13.1338
R337 VDDA.n65 VDDA.t69 13.1338
R338 VDDA.n67 VDDA.t76 13.1338
R339 VDDA.n67 VDDA.t136 13.1338
R340 VDDA.n69 VDDA.t25 13.1338
R341 VDDA.n69 VDDA.t9 13.1338
R342 VDDA.n71 VDDA.t6 13.1338
R343 VDDA.n71 VDDA.t74 13.1338
R344 VDDA.n73 VDDA.t64 13.1338
R345 VDDA.n73 VDDA.t93 13.1338
R346 VDDA.n75 VDDA.t21 13.1338
R347 VDDA.n75 VDDA.t80 13.1338
R348 VDDA VDDA.t57 12.8011
R349 VDDA.n77 VDDA.n76 11.0571
R350 VDDA.n117 VDDA.n116 10.869
R351 VDDA.n94 VDDA.n93 9.50883
R352 VDDA.n86 VDDA.n85 9.50883
R353 VDDA.n115 VDDA.n56 9.50883
R354 VDDA.n105 VDDA.n103 9.50883
R355 VDDA.n122 VDDA.n120 9.50883
R356 VDDA.n187 VDDA.n139 9.50883
R357 VDDA.n161 VDDA.n143 9.50883
R358 VDDA.n100 VDDA.n56 9.3005
R359 VDDA.n111 VDDA.n101 9.3005
R360 VDDA.n104 VDDA.n102 9.3005
R361 VDDA.n107 VDDA.n105 9.3005
R362 VDDA.n93 VDDA.n92 9.3005
R363 VDDA.n91 VDDA.n79 9.3005
R364 VDDA.n88 VDDA.n87 9.3005
R365 VDDA.n86 VDDA.n83 9.3005
R366 VDDA.n123 VDDA.n122 9.3005
R367 VDDA.n188 VDDA.n187 9.3005
R368 VDDA.n162 VDDA.n161 9.3005
R369 VDDA.n111 VDDA.n100 9.14336
R370 VDDA.n111 VDDA.n102 9.14336
R371 VDDA.n107 VDDA.n102 9.14336
R372 VDDA.n92 VDDA.n91 9.14336
R373 VDDA.n91 VDDA.n88 9.14336
R374 VDDA.n88 VDDA.n83 9.14336
R375 VDDA.n132 VDDA.n53 5.58881
R376 VDDA.n115 VDDA.n57 5.33286
R377 VDDA.n108 VDDA.n103 5.33286
R378 VDDA.n94 VDDA.n78 5.33286
R379 VDDA.n85 VDDA.n84 5.33286
R380 VDDA.n27 VDDA.n26 4.84425
R381 VDDA.n51 VDDA.n11 4.73979
R382 VDDA.n46 VDDA.n13 4.73979
R383 VDDA.n33 VDDA.n16 4.73979
R384 VDDA.n28 VDDA.n18 4.73979
R385 VDDA.n51 VDDA.n50 4.6505
R386 VDDA.n47 VDDA.n46 4.6505
R387 VDDA.n33 VDDA.n32 4.6505
R388 VDDA.n29 VDDA.n28 4.6505
R389 VDDA.n12 VDDA.n11 4.54311
R390 VDDA.n50 VDDA.n12 4.54311
R391 VDDA.n17 VDDA.n16 4.54311
R392 VDDA.n32 VDDA.n17 4.54311
R393 VDDA.n35 VDDA.n34 4.5005
R394 VDDA.n45 VDDA.n44 4.5005
R395 VDDA.n53 VDDA.n52 4.5005
R396 VDDA.n48 VDDA.n13 4.48641
R397 VDDA.n48 VDDA.n47 4.48641
R398 VDDA.n30 VDDA.n18 4.48641
R399 VDDA.n30 VDDA.n29 4.48641
R400 VDDA.n189 VDDA.n139 4.48641
R401 VDDA.n189 VDDA.n188 4.48641
R402 VDDA.n163 VDDA.n143 4.48641
R403 VDDA.n163 VDDA.n162 4.48641
R404 VDDA.n124 VDDA.n120 4.19264
R405 VDDA.n124 VDDA.n123 4.19264
R406 VDDA.n100 VDDA.n57 3.75335
R407 VDDA.n108 VDDA.n107 3.75335
R408 VDDA.n92 VDDA.n78 3.75335
R409 VDDA.n84 VDDA.n83 3.75335
R410 VDDA.n193 VDDA.n192 3.41464
R411 VDDA.n167 VDDA.n166 3.41464
R412 VDDA.n2 VDDA.n1 3.4105
R413 VDDA.n5 VDDA.n4 3.4105
R414 VDDA.n8 VDDA.n7 3.4105
R415 VDDA.n128 VDDA.n127 3.39381
R416 VDDA.n127 VDDA.n119 3.11118
R417 VDDA.n192 VDDA.n138 3.11118
R418 VDDA.n166 VDDA.n142 3.11118
R419 VDDA.n127 VDDA.n126 3.04304
R420 VDDA.n192 VDDA.n191 3.04304
R421 VDDA.n166 VDDA.n165 3.04304
R422 VDDA.n129 VDDA.n128 1.94319
R423 VDDA.n121 VDDA.n118 1.94319
R424 VDDA.n160 VDDA.n159 1.90152
R425 VDDA.n194 VDDA.n193 1.77652
R426 VDDA.n186 VDDA.n185 1.77652
R427 VDDA.n168 VDDA.n167 1.77652
R428 VDDA.n134 VDDA.n133 1.72394
R429 VDDA.n199 VDDA.n198 1.72394
R430 VDDA.n208 VDDA.n207 1.72394
R431 VDDA.n204 VDDA.n0 1.70194
R432 VDDA.n195 VDDA.n3 1.70194
R433 VDDA.n130 VDDA.n6 1.70194
R434 VDDA.n206 VDDA.n205 1.69525
R435 VDDA.n197 VDDA.n196 1.69525
R436 VDDA.n132 VDDA.n131 1.69525
R437 VDDA.n209 VDDA.n208 1.69525
R438 VDDA.n200 VDDA.n199 1.69525
R439 VDDA.n135 VDDA.n134 1.69525
R440 VDDA.n204 VDDA.n203 1.2502
R441 VDDA.n44 VDDA.n35 0.90675
R442 VDDA.n130 VDDA.n129 0.868689
R443 VDDA.n195 VDDA.n194 0.853064
R444 VDDA.n202 VDDA.n201 0.75233
R445 VDDA.n203 VDDA.n202 0.648391
R446 VDDA VDDA.n209 0.447
R447 VDDA.n26 VDDA.n24 0.34425
R448 VDDA.n24 VDDA.n22 0.34425
R449 VDDA.n22 VDDA.n20 0.34425
R450 VDDA.n20 VDDA.n15 0.34425
R451 VDDA.n35 VDDA.n15 0.34425
R452 VDDA.n44 VDDA.n43 0.34425
R453 VDDA.n43 VDDA.n41 0.34425
R454 VDDA.n41 VDDA.n39 0.34425
R455 VDDA.n39 VDDA.n37 0.34425
R456 VDDA.n37 VDDA.n10 0.34425
R457 VDDA.n53 VDDA.n10 0.34425
R458 VDDA.n185 VDDA.n168 0.333833
R459 VDDA.n118 VDDA.n117 0.328625
R460 VDDA.n206 VDDA.n200 0.304192
R461 VDDA.n187 VDDA.n186 0.2505
R462 VDDA.n161 VDDA.n160 0.2505
R463 VDDA.n197 VDDA.n135 0.230077
R464 VDDA.n122 VDDA.n121 0.229667
R465 VDDA.n129 VDDA.n118 0.229667
R466 VDDA.n93 VDDA.n79 0.208833
R467 VDDA.n87 VDDA.n79 0.208833
R468 VDDA.n87 VDDA.n86 0.208833
R469 VDDA.n101 VDDA.n56 0.208833
R470 VDDA.n104 VDDA.n101 0.208833
R471 VDDA.n105 VDDA.n104 0.208833
R472 VDDA.n76 VDDA.n74 0.188
R473 VDDA.n74 VDDA.n72 0.188
R474 VDDA.n72 VDDA.n70 0.188
R475 VDDA.n70 VDDA.n68 0.188
R476 VDDA.n68 VDDA.n66 0.188
R477 VDDA.n66 VDDA.n64 0.188
R478 VDDA.n64 VDDA.n55 0.188
R479 VDDA.n117 VDDA.n55 0.188
R480 VDDA.n46 VDDA.n45 0.182048
R481 VDDA.n28 VDDA.n27 0.182048
R482 VDDA.n52 VDDA.n51 0.182048
R483 VDDA.n34 VDDA.n33 0.182048
R484 VDDA.t34 VDDA.t91 0.1603
R485 VDDA.t70 VDDA.t26 0.1603
R486 VDDA.t7 VDDA.t90 0.1603
R487 VDDA.t0 VDDA.t67 0.1603
R488 VDDA.t143 VDDA.t61 0.1603
R489 VDDA.n211 VDDA.t62 0.159278
R490 VDDA.n212 VDDA.t58 0.159278
R491 VDDA.n213 VDDA.t49 0.159278
R492 VDDA.n214 VDDA.t134 0.159278
R493 VDDA.n214 VDDA.t34 0.1368
R494 VDDA.n214 VDDA.t50 0.1368
R495 VDDA.n213 VDDA.t70 0.1368
R496 VDDA.n213 VDDA.t153 0.1368
R497 VDDA.n212 VDDA.t7 0.1368
R498 VDDA.n212 VDDA.t28 0.1368
R499 VDDA.n211 VDDA.t0 0.1368
R500 VDDA.n211 VDDA.t27 0.1368
R501 VDDA.n210 VDDA.t143 0.1368
R502 VDDA.n210 VDDA.t144 0.1368
R503 VDDA.n159 VDDA.n157 0.1255
R504 VDDA.n157 VDDA.n155 0.1255
R505 VDDA.n155 VDDA.n153 0.1255
R506 VDDA.n153 VDDA.n151 0.1255
R507 VDDA.n151 VDDA.n149 0.1255
R508 VDDA.n149 VDDA.n147 0.1255
R509 VDDA.n147 VDDA.n145 0.1255
R510 VDDA.n145 VDDA.n141 0.1255
R511 VDDA.n168 VDDA.n141 0.1255
R512 VDDA.n185 VDDA.n184 0.1255
R513 VDDA.n184 VDDA.n182 0.1255
R514 VDDA.n182 VDDA.n180 0.1255
R515 VDDA.n180 VDDA.n178 0.1255
R516 VDDA.n178 VDDA.n176 0.1255
R517 VDDA.n176 VDDA.n174 0.1255
R518 VDDA.n174 VDDA.n172 0.1255
R519 VDDA.n172 VDDA.n170 0.1255
R520 VDDA.n170 VDDA.n137 0.1255
R521 VDDA.n194 VDDA.n137 0.1255
R522 VDDA.n131 VDDA.n7 0.0224982
R523 VDDA.n196 VDDA.n4 0.0224982
R524 VDDA.n205 VDDA.n1 0.0224982
R525 VDDA.n205 VDDA.n204 0.0224982
R526 VDDA.n196 VDDA.n195 0.0224982
R527 VDDA.n131 VDDA.n130 0.0224982
R528 VDDA.n208 VDDA.n1 0.0224982
R529 VDDA.n199 VDDA.n4 0.0224982
R530 VDDA.n134 VDDA.n7 0.0224982
R531 VDDA.n133 VDDA.n8 0.00911526
R532 VDDA.n198 VDDA.n5 0.00911526
R533 VDDA.n207 VDDA.n2 0.00911526
R534 VDDA.n207 VDDA.n206 0.00911526
R535 VDDA.n198 VDDA.n197 0.00911526
R536 VDDA.n133 VDDA.n132 0.00911526
R537 VDDA.n8 VDDA.n6 0.00911526
R538 VDDA.n5 VDDA.n3 0.00911526
R539 VDDA.n2 VDDA.n0 0.00911526
R540 VDDA.n209 VDDA.n0 0.00911526
R541 VDDA.n200 VDDA.n3 0.00911526
R542 VDDA.n135 VDDA.n6 0.00911526
R543 VDDA.t62 VDDA.n210 0.00152174
R544 VDDA.t58 VDDA.n211 0.00152174
R545 VDDA.t49 VDDA.n212 0.00152174
R546 VDDA.t134 VDDA.n213 0.00152174
R547 VDDA.t57 VDDA.n214 0.00152174
R548 V_CUR_REF_REG V_CUR_REF_REG.t13 701.501
R549 V_CUR_REF_REG.n2 V_CUR_REF_REG.n0 302.507
R550 V_CUR_REF_REG.n2 V_CUR_REF_REG.n1 302.163
R551 V_CUR_REF_REG.n4 V_CUR_REF_REG.n3 302.163
R552 V_CUR_REF_REG.n6 V_CUR_REF_REG.n5 302.163
R553 V_CUR_REF_REG.n8 V_CUR_REF_REG.n7 302.163
R554 V_CUR_REF_REG.n10 V_CUR_REF_REG.n9 302.163
R555 V_CUR_REF_REG.n11 V_CUR_REF_REG.t0 133.911
R556 V_CUR_REF_REG.n0 V_CUR_REF_REG.t4 39.4005
R557 V_CUR_REF_REG.n0 V_CUR_REF_REG.t1 39.4005
R558 V_CUR_REF_REG.n1 V_CUR_REF_REG.t6 39.4005
R559 V_CUR_REF_REG.n1 V_CUR_REF_REG.t9 39.4005
R560 V_CUR_REF_REG.n3 V_CUR_REF_REG.t7 39.4005
R561 V_CUR_REF_REG.n3 V_CUR_REF_REG.t11 39.4005
R562 V_CUR_REF_REG.n5 V_CUR_REF_REG.t8 39.4005
R563 V_CUR_REF_REG.n5 V_CUR_REF_REG.t12 39.4005
R564 V_CUR_REF_REG.n7 V_CUR_REF_REG.t10 39.4005
R565 V_CUR_REF_REG.n7 V_CUR_REF_REG.t5 39.4005
R566 V_CUR_REF_REG.n9 V_CUR_REF_REG.t2 39.4005
R567 V_CUR_REF_REG.n9 V_CUR_REF_REG.t3 39.4005
R568 V_CUR_REF_REG.n11 V_CUR_REF_REG.n10 12.3599
R569 V_CUR_REF_REG V_CUR_REF_REG.n11 5.48488
R570 V_CUR_REF_REG.n10 V_CUR_REF_REG.n8 0.34425
R571 V_CUR_REF_REG.n8 V_CUR_REF_REG.n6 0.34425
R572 V_CUR_REF_REG.n6 V_CUR_REF_REG.n4 0.34425
R573 V_CUR_REF_REG.n4 V_CUR_REF_REG.n2 0.34425
R574 1st_Vout_1.n3 1st_Vout_1.t19 363.911
R575 1st_Vout_1.n4 1st_Vout_1.t17 351.976
R576 1st_Vout_1.n4 1st_Vout_1.n5 299.252
R577 1st_Vout_1.n3 1st_Vout_1.n7 299.252
R578 1st_Vout_1.n10 1st_Vout_1.n9 297.805
R579 1st_Vout_1.n8 1st_Vout_1.t28 194.809
R580 1st_Vout_1.n8 1st_Vout_1.t14 194.809
R581 1st_Vout_1.n6 1st_Vout_1.t21 194.809
R582 1st_Vout_1.n6 1st_Vout_1.t8 194.809
R583 1st_Vout_1.n3 1st_Vout_1.n8 163.1
R584 1st_Vout_1.n4 1st_Vout_1.n6 163.1
R585 1st_Vout_1.t6 1st_Vout_1.n10 49.4489
R586 1st_Vout_1.n7 1st_Vout_1.t2 39.4005
R587 1st_Vout_1.n7 1st_Vout_1.t5 39.4005
R588 1st_Vout_1.n5 1st_Vout_1.t3 39.4005
R589 1st_Vout_1.n5 1st_Vout_1.t0 39.4005
R590 1st_Vout_1.n9 1st_Vout_1.t1 39.4005
R591 1st_Vout_1.n9 1st_Vout_1.t4 39.4005
R592 1st_Vout_1.n1 1st_Vout_1.t20 4.8295
R593 1st_Vout_1.n1 1st_Vout_1.t31 4.8295
R594 1st_Vout_1.n2 1st_Vout_1.t13 4.8295
R595 1st_Vout_1.n2 1st_Vout_1.t24 4.8295
R596 1st_Vout_1.n2 1st_Vout_1.t16 4.8295
R597 1st_Vout_1.n2 1st_Vout_1.t29 4.8295
R598 1st_Vout_1.n0 1st_Vout_1.t10 4.8295
R599 1st_Vout_1.n0 1st_Vout_1.t22 4.8295
R600 1st_Vout_1.n0 1st_Vout_1.t26 4.8295
R601 1st_Vout_1.n1 1st_Vout_1.t18 4.5005
R602 1st_Vout_1.n1 1st_Vout_1.t32 4.5005
R603 1st_Vout_1.n2 1st_Vout_1.t11 4.5005
R604 1st_Vout_1.n2 1st_Vout_1.t25 4.5005
R605 1st_Vout_1.n2 1st_Vout_1.t15 4.5005
R606 1st_Vout_1.n2 1st_Vout_1.t30 4.5005
R607 1st_Vout_1.n0 1st_Vout_1.t9 4.5005
R608 1st_Vout_1.n0 1st_Vout_1.t23 4.5005
R609 1st_Vout_1.n0 1st_Vout_1.t12 4.5005
R610 1st_Vout_1.n0 1st_Vout_1.t27 4.5005
R611 1st_Vout_1.n0 1st_Vout_1.t7 4.5005
R612 1st_Vout_1.n3 1st_Vout_1.n0 8.9477
R613 1st_Vout_1.n0 1st_Vout_1.n2 2.2095
R614 1st_Vout_1.n10 1st_Vout_1.n4 1.44719
R615 1st_Vout_1.n4 1st_Vout_1.n3 0.96925
R616 1st_Vout_1.n2 1st_Vout_1.n1 0.8935
R617 cap_res1 cap_res1.t0 114.728
R618 cap_res1 cap_res1.t20 3.8015
R619 cap_res1.t5 cap_res1.t16 0.1603
R620 cap_res1.t19 cap_res1.t18 0.1603
R621 cap_res1.t14 cap_res1.t13 0.1603
R622 cap_res1.t17 cap_res1.t15 0.1603
R623 cap_res1.t12 cap_res1.t11 0.1603
R624 cap_res1.n1 cap_res1.t1 0.159278
R625 cap_res1.n2 cap_res1.t7 0.159278
R626 cap_res1.n3 cap_res1.t3 0.159278
R627 cap_res1.n4 cap_res1.t9 0.159278
R628 cap_res1.n4 cap_res1.t6 0.1368
R629 cap_res1.n4 cap_res1.t5 0.1368
R630 cap_res1.n3 cap_res1.t10 0.1368
R631 cap_res1.n3 cap_res1.t19 0.1368
R632 cap_res1.n2 cap_res1.t4 0.1368
R633 cap_res1.n2 cap_res1.t14 0.1368
R634 cap_res1.n1 cap_res1.t8 0.1368
R635 cap_res1.n1 cap_res1.t17 0.1368
R636 cap_res1.n0 cap_res1.t2 0.1368
R637 cap_res1.n0 cap_res1.t12 0.1368
R638 cap_res1.t1 cap_res1.n0 0.00152174
R639 cap_res1.t7 cap_res1.n1 0.00152174
R640 cap_res1.t3 cap_res1.n2 0.00152174
R641 cap_res1.t9 cap_res1.n3 0.00152174
R642 cap_res1.t20 cap_res1.n4 0.00152174
R643 CURRENT_OUTPUT.n3 CURRENT_OUTPUT.n1 302.507
R644 CURRENT_OUTPUT.n8 CURRENT_OUTPUT.n7 302.163
R645 CURRENT_OUTPUT.n10 CURRENT_OUTPUT.n9 302.163
R646 CURRENT_OUTPUT.n3 CURRENT_OUTPUT.n2 302.163
R647 CURRENT_OUTPUT.n12 CURRENT_OUTPUT.n0 297.663
R648 CURRENT_OUTPUT.n6 CURRENT_OUTPUT.n4 297.599
R649 CURRENT_OUTPUT.n4 CURRENT_OUTPUT.t4 39.4005
R650 CURRENT_OUTPUT.n4 CURRENT_OUTPUT.t1 39.4005
R651 CURRENT_OUTPUT.n7 CURRENT_OUTPUT.t6 39.4005
R652 CURRENT_OUTPUT.n7 CURRENT_OUTPUT.t10 39.4005
R653 CURRENT_OUTPUT.n9 CURRENT_OUTPUT.t7 39.4005
R654 CURRENT_OUTPUT.n9 CURRENT_OUTPUT.t11 39.4005
R655 CURRENT_OUTPUT.n0 CURRENT_OUTPUT.t9 39.4005
R656 CURRENT_OUTPUT.n0 CURRENT_OUTPUT.t2 39.4005
R657 CURRENT_OUTPUT.n2 CURRENT_OUTPUT.t8 39.4005
R658 CURRENT_OUTPUT.n2 CURRENT_OUTPUT.t5 39.4005
R659 CURRENT_OUTPUT.n1 CURRENT_OUTPUT.t0 39.4005
R660 CURRENT_OUTPUT.n1 CURRENT_OUTPUT.t3 39.4005
R661 CURRENT_OUTPUT.n8 CURRENT_OUTPUT.n6 4.84425
R662 CURRENT_OUTPUT.n12 CURRENT_OUTPUT.n11 4.5005
R663 CURRENT_OUTPUT CURRENT_OUTPUT.n12 0.78175
R664 CURRENT_OUTPUT.n11 CURRENT_OUTPUT.n3 0.34425
R665 CURRENT_OUTPUT.n11 CURRENT_OUTPUT.n10 0.34425
R666 CURRENT_OUTPUT.n10 CURRENT_OUTPUT.n8 0.34425
R667 CURRENT_OUTPUT.n6 CURRENT_OUTPUT.n5 0.153278
R668 V_TOP.n1 V_TOP.t28 312.798
R669 V_TOP V_TOP.t16 312.639
R670 V_TOP.n36 V_TOP.t45 312.5
R671 V_TOP.n1 V_TOP.t36 310.401
R672 V_TOP.n2 V_TOP.t41 310.401
R673 V_TOP.n3 V_TOP.t48 310.401
R674 V_TOP.n4 V_TOP.t15 310.401
R675 V_TOP.n5 V_TOP.t26 310.401
R676 V_TOP.n37 V_TOP.t14 310.401
R677 V_TOP.n38 V_TOP.t22 310.401
R678 V_TOP.n39 V_TOP.t31 310.401
R679 V_TOP.n40 V_TOP.t38 310.401
R680 V_TOP.n41 V_TOP.t42 310.401
R681 V_TOP.n42 V_TOP.t49 310.401
R682 V_TOP.n34 V_TOP.t39 308
R683 V_TOP.n22 V_TOP.n21 306.808
R684 V_TOP.n7 V_TOP.t34 305.901
R685 V_TOP.n27 V_TOP.n26 301.933
R686 V_TOP.n29 V_TOP.n28 301.933
R687 V_TOP.n31 V_TOP.n30 301.933
R688 V_TOP.n22 V_TOP.n20 297.433
R689 V_TOP.n24 V_TOP.n23 297.433
R690 V_TOP.n19 V_TOP.t2 108.424
R691 V_TOP.n32 V_TOP.t7 99.3386
R692 V_TOP.n21 V_TOP.t3 39.4005
R693 V_TOP.n21 V_TOP.t0 39.4005
R694 V_TOP.n20 V_TOP.t1 39.4005
R695 V_TOP.n20 V_TOP.t4 39.4005
R696 V_TOP.n23 V_TOP.t10 39.4005
R697 V_TOP.n23 V_TOP.t6 39.4005
R698 V_TOP.n26 V_TOP.t12 39.4005
R699 V_TOP.n26 V_TOP.t8 39.4005
R700 V_TOP.n28 V_TOP.t13 39.4005
R701 V_TOP.n28 V_TOP.t9 39.4005
R702 V_TOP.n30 V_TOP.t5 39.4005
R703 V_TOP.n30 V_TOP.t11 39.4005
R704 V_TOP.n19 V_TOP.n18 28.0324
R705 V_TOP.n25 V_TOP.n19 14.5688
R706 V_TOP.n32 V_TOP.n31 4.90675
R707 V_TOP.n9 V_TOP.t47 4.8295
R708 V_TOP.n8 V_TOP.t25 4.8295
R709 V_TOP.n11 V_TOP.t35 4.8295
R710 V_TOP.n10 V_TOP.t19 4.8295
R711 V_TOP.n13 V_TOP.t44 4.8295
R712 V_TOP.n12 V_TOP.t23 4.8295
R713 V_TOP.n15 V_TOP.t32 4.8295
R714 V_TOP.n14 V_TOP.t17 4.8295
R715 V_TOP.n16 V_TOP.t40 4.8295
R716 V_TOP.n9 V_TOP.t46 4.5005
R717 V_TOP.n8 V_TOP.t27 4.5005
R718 V_TOP.n11 V_TOP.t33 4.5005
R719 V_TOP.n10 V_TOP.t20 4.5005
R720 V_TOP.n13 V_TOP.t43 4.5005
R721 V_TOP.n12 V_TOP.t24 4.5005
R722 V_TOP.n15 V_TOP.t30 4.5005
R723 V_TOP.n14 V_TOP.t18 4.5005
R724 V_TOP.n16 V_TOP.t29 4.5005
R725 V_TOP.n17 V_TOP.t37 4.5005
R726 V_TOP.n18 V_TOP.t21 4.5005
R727 V_TOP.n35 V_TOP.n34 4.5005
R728 V_TOP.n33 V_TOP.n0 4.5005
R729 V_TOP.n7 V_TOP.n6 4.5005
R730 V_TOP.n25 V_TOP.n24 4.5005
R731 V_TOP.n24 V_TOP.n22 1.59425
R732 V_TOP.n33 V_TOP.n32 1.21925
R733 V_TOP.n31 V_TOP.n29 1.1255
R734 V_TOP.n29 V_TOP.n27 1.1255
R735 V_TOP.n27 V_TOP.n25 1.1255
R736 V_TOP.n9 V_TOP.n8 0.3295
R737 V_TOP.n11 V_TOP.n10 0.3295
R738 V_TOP.n13 V_TOP.n12 0.3295
R739 V_TOP.n15 V_TOP.n14 0.3295
R740 V_TOP.n17 V_TOP.n16 0.3295
R741 V_TOP.n18 V_TOP.n17 0.3295
R742 V_TOP.n11 V_TOP.n9 0.2825
R743 V_TOP.n13 V_TOP.n11 0.2825
R744 V_TOP.n15 V_TOP.n13 0.2825
R745 V_TOP.n16 V_TOP.n15 0.2825
R746 V_TOP.n42 V_TOP.n41 0.28175
R747 V_TOP.n41 V_TOP.n40 0.28175
R748 V_TOP.n40 V_TOP.n39 0.28175
R749 V_TOP.n39 V_TOP.n38 0.28175
R750 V_TOP.n38 V_TOP.n37 0.28175
R751 V_TOP.n37 V_TOP.n36 0.28175
R752 V_TOP.n36 V_TOP.n35 0.28175
R753 V_TOP.n6 V_TOP.n5 0.28175
R754 V_TOP.n5 V_TOP.n4 0.28175
R755 V_TOP.n4 V_TOP.n3 0.28175
R756 V_TOP.n3 V_TOP.n2 0.28175
R757 V_TOP.n2 V_TOP.n1 0.28175
R758 V_TOP V_TOP.n42 0.141125
R759 V_TOP.n35 V_TOP.n0 0.141125
R760 V_TOP.n6 V_TOP.n0 0.141125
R761 V_TOP.n34 V_TOP.n33 0.141125
R762 V_TOP.n33 V_TOP.n7 0.141125
R763 Vin+ Vin+.t6 529.879
R764 Vin+.n3 Vin+.t0 148.653
R765 Vin+.n3 Vin+.t1 125.418
R766 Vin+.n2 Vin+.n0 105.609
R767 Vin+.n2 Vin+.n1 104.484
R768 Vin+.n4 Vin+.n3 21.4871
R769 Vin+.n4 Vin+.n2 14.8911
R770 Vin+.n1 Vin+.t2 13.1338
R771 Vin+.n1 Vin+.t3 13.1338
R772 Vin+.n0 Vin+.t4 13.1338
R773 Vin+.n0 Vin+.t5 13.1338
R774 Vin+ Vin+.n4 6.53175
R775 START_UP_NFET1.t1 START_UP_NFET1.t0 178.194
R776 GNDA.n2054 GNDA.n2053 14052.5
R777 GNDA.n2054 GNDA.n19 10589.3
R778 GNDA.t16 GNDA.n2054 4573.59
R779 GNDA.n2053 GNDA.t27 1721.74
R780 GNDA.n1405 GNDA.n1249 1141.35
R781 GNDA.n1543 GNDA.n19 1109.84
R782 GNDA.n1854 GNDA.n1853 686.717
R783 GNDA.n1632 GNDA.n1631 686.717
R784 GNDA.n1542 GNDA.n1541 686.717
R785 GNDA.n1542 GNDA.n223 686.717
R786 GNDA.n1628 GNDA.n1617 686.717
R787 GNDA.n1846 GNDA.n182 686.717
R788 GNDA.n1816 GNDA.n1815 669.307
R789 GNDA.n1826 GNDA.n1824 669.307
R790 GNDA.n253 GNDA.n249 654.447
R791 GNDA.n977 GNDA.n23 585
R792 GNDA.n1001 GNDA.n850 585
R793 GNDA.n999 GNDA.n998 585
R794 GNDA.n997 GNDA.n852 585
R795 GNDA.n996 GNDA.n995 585
R796 GNDA.n993 GNDA.n853 585
R797 GNDA.n991 GNDA.n990 585
R798 GNDA.n989 GNDA.n854 585
R799 GNDA.n988 GNDA.n987 585
R800 GNDA.n985 GNDA.n855 585
R801 GNDA.n983 GNDA.n982 585
R802 GNDA.n981 GNDA.n856 585
R803 GNDA.n2031 GNDA.n2030 585
R804 GNDA.n2032 GNDA.n30 585
R805 GNDA.n2034 GNDA.n2033 585
R806 GNDA.n2036 GNDA.n28 585
R807 GNDA.n2038 GNDA.n2037 585
R808 GNDA.n2039 GNDA.n27 585
R809 GNDA.n2041 GNDA.n2040 585
R810 GNDA.n2043 GNDA.n25 585
R811 GNDA.n2045 GNDA.n2044 585
R812 GNDA.n2046 GNDA.n24 585
R813 GNDA.n2048 GNDA.n2047 585
R814 GNDA.n1384 GNDA.n1383 585
R815 GNDA.n1383 GNDA.n1382 585
R816 GNDA.n1384 GNDA.n1260 585
R817 GNDA.n1260 GNDA.n1259 585
R818 GNDA.n1386 GNDA.n1385 585
R819 GNDA.n1387 GNDA.n1386 585
R820 GNDA.n1258 GNDA.n1257 585
R821 GNDA.n1388 GNDA.n1258 585
R822 GNDA.n1392 GNDA.n1391 585
R823 GNDA.n1391 GNDA.n1390 585
R824 GNDA.n1393 GNDA.n1256 585
R825 GNDA.n1389 GNDA.n1256 585
R826 GNDA.n1395 GNDA.n1394 585
R827 GNDA.n1395 GNDA.n1243 585
R828 GNDA.n1396 GNDA.n1255 585
R829 GNDA.n1396 GNDA.n1244 585
R830 GNDA.n1399 GNDA.n1398 585
R831 GNDA.n1398 GNDA.n1397 585
R832 GNDA.n1400 GNDA.n1254 585
R833 GNDA.n1254 GNDA.n1253 585
R834 GNDA.n1402 GNDA.n1401 585
R835 GNDA.n1403 GNDA.n1402 585
R836 GNDA.n1252 GNDA.n1251 585
R837 GNDA.n1404 GNDA.n1252 585
R838 GNDA.n1407 GNDA.n1406 585
R839 GNDA.n1406 GNDA.n1405 585
R840 GNDA.n571 GNDA.n570 585
R841 GNDA.n570 GNDA.n52 585
R842 GNDA.n571 GNDA.n569 585
R843 GNDA.n569 GNDA.n568 585
R844 GNDA.n509 GNDA.n508 585
R845 GNDA.n567 GNDA.n509 585
R846 GNDA.n565 GNDA.n564 585
R847 GNDA.n566 GNDA.n565 585
R848 GNDA.n563 GNDA.n511 585
R849 GNDA.n511 GNDA.n510 585
R850 GNDA.n562 GNDA.n561 585
R851 GNDA.n561 GNDA.n560 585
R852 GNDA.n559 GNDA.n512 585
R853 GNDA.n559 GNDA.n59 585
R854 GNDA.n558 GNDA.n557 585
R855 GNDA.n558 GNDA.n60 585
R856 GNDA.n556 GNDA.n513 585
R857 GNDA.n516 GNDA.n513 585
R858 GNDA.n555 GNDA.n554 585
R859 GNDA.n554 GNDA.n553 585
R860 GNDA.n515 GNDA.n514 585
R861 GNDA.n552 GNDA.n515 585
R862 GNDA.n550 GNDA.n549 585
R863 GNDA.n551 GNDA.n550 585
R864 GNDA.n548 GNDA.n518 585
R865 GNDA.n518 GNDA.n517 585
R866 GNDA.n1548 GNDA.n1546 585
R867 GNDA.n1600 GNDA.n1548 585
R868 GNDA.n1598 GNDA.n1597 585
R869 GNDA.n1599 GNDA.n1598 585
R870 GNDA.n1596 GNDA.n1550 585
R871 GNDA.n1550 GNDA.n1549 585
R872 GNDA.n1595 GNDA.n1594 585
R873 GNDA.n1594 GNDA.n1593 585
R874 GNDA.n1592 GNDA.n1551 585
R875 GNDA.n1592 GNDA.n66 585
R876 GNDA.n1591 GNDA.n1590 585
R877 GNDA.n1591 GNDA.n67 585
R878 GNDA.n1589 GNDA.n1552 585
R879 GNDA.n1555 GNDA.n1552 585
R880 GNDA.n1588 GNDA.n1587 585
R881 GNDA.n1587 GNDA.n1586 585
R882 GNDA.n1554 GNDA.n1553 585
R883 GNDA.n1585 GNDA.n1554 585
R884 GNDA.n1583 GNDA.n1582 585
R885 GNDA.n1584 GNDA.n1583 585
R886 GNDA.n1581 GNDA.n1556 585
R887 GNDA.n1556 GNDA.n53 585
R888 GNDA.n161 GNDA.n21 585
R889 GNDA.n21 GNDA.n20 585
R890 GNDA.n1875 GNDA.n1874 585
R891 GNDA.n1874 GNDA.n1873 585
R892 GNDA.n164 GNDA.n163 585
R893 GNDA.n1872 GNDA.n164 585
R894 GNDA.n1870 GNDA.n1869 585
R895 GNDA.n1871 GNDA.n1870 585
R896 GNDA.n1864 GNDA.n165 585
R897 GNDA.n1856 GNDA.n165 585
R898 GNDA.n1859 GNDA.n1858 585
R899 GNDA.n1858 GNDA.n1857 585
R900 GNDA.n167 GNDA.n166 585
R901 GNDA.n181 GNDA.n167 585
R902 GNDA.n179 GNDA.n178 585
R903 GNDA.n180 GNDA.n179 585
R904 GNDA.n173 GNDA.n171 585
R905 GNDA.n171 GNDA.n168 585
R906 GNDA.n170 GNDA.n140 585
R907 GNDA.n170 GNDA.n169 585
R908 GNDA.n1931 GNDA.n138 585
R909 GNDA.n138 GNDA.n137 585
R910 GNDA.n1934 GNDA.n1933 585
R911 GNDA.n1935 GNDA.n1934 585
R912 GNDA.n2052 GNDA.n2051 585
R913 GNDA.n1621 GNDA.n1619 585
R914 GNDA.n1625 GNDA.n1618 585
R915 GNDA.n1633 GNDA.n1618 585
R916 GNDA.n1624 GNDA.n1623 585
R917 GNDA.n186 GNDA.n184 585
R918 GNDA.n1851 GNDA.n183 585
R919 GNDA.n1855 GNDA.n183 585
R920 GNDA.n1849 GNDA.n1848 585
R921 GNDA.n197 GNDA.n196 585
R922 GNDA.n1819 GNDA.n1818 585
R923 GNDA.n1818 GNDA.n1817 585
R924 GNDA.n1830 GNDA.n1825 585
R925 GNDA.n1829 GNDA.n1828 585
R926 GNDA.n1828 GNDA.n1827 585
R927 GNDA.n663 GNDA.n662 585
R928 GNDA.n660 GNDA.n659 585
R929 GNDA.n658 GNDA.n657 585
R930 GNDA.n632 GNDA.n482 585
R931 GNDA.n638 GNDA.n637 585
R932 GNDA.n640 GNDA.n631 585
R933 GNDA.n642 GNDA.n641 585
R934 GNDA.n628 GNDA.n627 585
R935 GNDA.n648 GNDA.n647 585
R936 GNDA.n651 GNDA.n650 585
R937 GNDA.n626 GNDA.n505 585
R938 GNDA.n624 GNDA.n623 585
R939 GNDA.n787 GNDA.n786 585
R940 GNDA.n784 GNDA.n783 585
R941 GNDA.n669 GNDA.n668 585
R942 GNDA.n777 GNDA.n776 585
R943 GNDA.n774 GNDA.n773 585
R944 GNDA.n763 GNDA.n762 585
R945 GNDA.n765 GNDA.n764 585
R946 GNDA.n760 GNDA.n676 585
R947 GNDA.n759 GNDA.n758 585
R948 GNDA.n749 GNDA.n678 585
R949 GNDA.n751 GNDA.n750 585
R950 GNDA.n747 GNDA.n746 585
R951 GNDA.n976 GNDA.n857 585
R952 GNDA.n974 GNDA.n973 585
R953 GNDA.n893 GNDA.n858 585
R954 GNDA.n891 GNDA.n890 585
R955 GNDA.n903 GNDA.n902 585
R956 GNDA.n905 GNDA.n888 585
R957 GNDA.n907 GNDA.n906 585
R958 GNDA.n884 GNDA.n883 585
R959 GNDA.n914 GNDA.n913 585
R960 GNDA.n917 GNDA.n916 585
R961 GNDA.n882 GNDA.n878 585
R962 GNDA.n880 GNDA.n788 585
R963 GNDA.n1558 GNDA.n1557 585
R964 GNDA.n1560 GNDA.n1559 585
R965 GNDA.n1562 GNDA.n1561 585
R966 GNDA.n1564 GNDA.n1563 585
R967 GNDA.n1566 GNDA.n1565 585
R968 GNDA.n1568 GNDA.n1567 585
R969 GNDA.n1570 GNDA.n1569 585
R970 GNDA.n1572 GNDA.n1571 585
R971 GNDA.n1574 GNDA.n1573 585
R972 GNDA.n1576 GNDA.n1575 585
R973 GNDA.n1578 GNDA.n1577 585
R974 GNDA.n1580 GNDA.n1579 585
R975 GNDA.n1979 GNDA.n1978 585
R976 GNDA.n1981 GNDA.n1980 585
R977 GNDA.n1983 GNDA.n1982 585
R978 GNDA.n1985 GNDA.n1984 585
R979 GNDA.n1987 GNDA.n1986 585
R980 GNDA.n1989 GNDA.n1988 585
R981 GNDA.n1991 GNDA.n1990 585
R982 GNDA.n1993 GNDA.n1992 585
R983 GNDA.n1995 GNDA.n1994 585
R984 GNDA.n1997 GNDA.n1996 585
R985 GNDA.n1999 GNDA.n1998 585
R986 GNDA.n2001 GNDA.n2000 585
R987 GNDA.n2029 GNDA.n31 585
R988 GNDA.n102 GNDA.n33 585
R989 GNDA.n104 GNDA.n103 585
R990 GNDA.n106 GNDA.n105 585
R991 GNDA.n108 GNDA.n107 585
R992 GNDA.n110 GNDA.n109 585
R993 GNDA.n112 GNDA.n111 585
R994 GNDA.n114 GNDA.n113 585
R995 GNDA.n116 GNDA.n115 585
R996 GNDA.n118 GNDA.n117 585
R997 GNDA.n120 GNDA.n119 585
R998 GNDA.n122 GNDA.n121 585
R999 GNDA.n1318 GNDA.n1091 585
R1000 GNDA.n1321 GNDA.n1320 585
R1001 GNDA.n1317 GNDA.n1287 585
R1002 GNDA.n1315 GNDA.n1314 585
R1003 GNDA.n1309 GNDA.n1288 585
R1004 GNDA.n1304 GNDA.n1303 585
R1005 GNDA.n1301 GNDA.n1289 585
R1006 GNDA.n1299 GNDA.n1298 585
R1007 GNDA.n1293 GNDA.n1291 585
R1008 GNDA.n1264 GNDA.n1262 585
R1009 GNDA.n1378 GNDA.n1377 585
R1010 GNDA.n1380 GNDA.n1261 585
R1011 GNDA.n527 GNDA.n463 585
R1012 GNDA.n529 GNDA.n525 585
R1013 GNDA.n531 GNDA.n530 585
R1014 GNDA.n532 GNDA.n524 585
R1015 GNDA.n534 GNDA.n533 585
R1016 GNDA.n536 GNDA.n522 585
R1017 GNDA.n538 GNDA.n537 585
R1018 GNDA.n539 GNDA.n521 585
R1019 GNDA.n541 GNDA.n540 585
R1020 GNDA.n543 GNDA.n520 585
R1021 GNDA.n544 GNDA.n519 585
R1022 GNDA.n547 GNDA.n546 585
R1023 GNDA.n840 GNDA.n839 585
R1024 GNDA.n837 GNDA.n813 585
R1025 GNDA.n836 GNDA.n835 585
R1026 GNDA.n834 GNDA.n833 585
R1027 GNDA.n832 GNDA.n815 585
R1028 GNDA.n830 GNDA.n829 585
R1029 GNDA.n828 GNDA.n816 585
R1030 GNDA.n827 GNDA.n826 585
R1031 GNDA.n824 GNDA.n817 585
R1032 GNDA.n822 GNDA.n821 585
R1033 GNDA.n820 GNDA.n819 585
R1034 GNDA.n466 GNDA.n462 585
R1035 GNDA.n1003 GNDA.n1002 585
R1036 GNDA.n1004 GNDA.n849 585
R1037 GNDA.n1006 GNDA.n1005 585
R1038 GNDA.n1008 GNDA.n847 585
R1039 GNDA.n1010 GNDA.n1009 585
R1040 GNDA.n1011 GNDA.n846 585
R1041 GNDA.n1013 GNDA.n1012 585
R1042 GNDA.n1015 GNDA.n844 585
R1043 GNDA.n1017 GNDA.n1016 585
R1044 GNDA.n1018 GNDA.n843 585
R1045 GNDA.n1020 GNDA.n1019 585
R1046 GNDA.n1022 GNDA.n842 585
R1047 GNDA.n1431 GNDA.n1430 585
R1048 GNDA.n1430 GNDA.n1429 585
R1049 GNDA.n1228 GNDA.n1227 585
R1050 GNDA.n1428 GNDA.n1228 585
R1051 GNDA.n1426 GNDA.n1425 585
R1052 GNDA.n1427 GNDA.n1426 585
R1053 GNDA.n1424 GNDA.n1230 585
R1054 GNDA.n1230 GNDA.n1229 585
R1055 GNDA.n1423 GNDA.n1422 585
R1056 GNDA.n1422 GNDA.n1421 585
R1057 GNDA.n1232 GNDA.n1231 585
R1058 GNDA.n1420 GNDA.n1232 585
R1059 GNDA.n1418 GNDA.n1417 585
R1060 GNDA.n1419 GNDA.n1418 585
R1061 GNDA.n1416 GNDA.n1246 585
R1062 GNDA.n1246 GNDA.n1245 585
R1063 GNDA.n1415 GNDA.n1414 585
R1064 GNDA.n1414 GNDA.n1413 585
R1065 GNDA.n1248 GNDA.n1247 585
R1066 GNDA.n1412 GNDA.n1248 585
R1067 GNDA.n1410 GNDA.n1409 585
R1068 GNDA.n1411 GNDA.n1410 585
R1069 GNDA.n1408 GNDA.n1250 585
R1070 GNDA.n1250 GNDA.n1249 585
R1071 GNDA.n438 GNDA.n437 585
R1072 GNDA.n437 GNDA.n55 585
R1073 GNDA.n439 GNDA.n284 585
R1074 GNDA.n284 GNDA.n283 585
R1075 GNDA.n441 GNDA.n440 585
R1076 GNDA.n442 GNDA.n441 585
R1077 GNDA.n282 GNDA.n281 585
R1078 GNDA.n443 GNDA.n282 585
R1079 GNDA.n446 GNDA.n445 585
R1080 GNDA.n445 GNDA.n444 585
R1081 GNDA.n447 GNDA.n280 585
R1082 GNDA.n280 GNDA.n58 585
R1083 GNDA.n449 GNDA.n448 585
R1084 GNDA.n449 GNDA.n57 585
R1085 GNDA.n450 GNDA.n279 585
R1086 GNDA.n451 GNDA.n450 585
R1087 GNDA.n454 GNDA.n453 585
R1088 GNDA.n453 GNDA.n452 585
R1089 GNDA.n455 GNDA.n278 585
R1090 GNDA.n278 GNDA.n277 585
R1091 GNDA.n457 GNDA.n456 585
R1092 GNDA.n458 GNDA.n457 585
R1093 GNDA.n262 GNDA.n259 585
R1094 GNDA.n459 GNDA.n262 585
R1095 GNDA.n436 GNDA.n285 585
R1096 GNDA.n436 GNDA.n23 585
R1097 GNDA.n435 GNDA.n286 585
R1098 GNDA.n433 GNDA.n432 585
R1099 GNDA.n431 GNDA.n287 585
R1100 GNDA.n430 GNDA.n429 585
R1101 GNDA.n427 GNDA.n288 585
R1102 GNDA.n425 GNDA.n424 585
R1103 GNDA.n423 GNDA.n289 585
R1104 GNDA.n422 GNDA.n421 585
R1105 GNDA.n419 GNDA.n290 585
R1106 GNDA.n417 GNDA.n416 585
R1107 GNDA.n412 GNDA.n292 585
R1108 GNDA.n410 GNDA.n409 585
R1109 GNDA.n329 GNDA.n293 585
R1110 GNDA.n327 GNDA.n326 585
R1111 GNDA.n339 GNDA.n338 585
R1112 GNDA.n341 GNDA.n324 585
R1113 GNDA.n343 GNDA.n342 585
R1114 GNDA.n320 GNDA.n319 585
R1115 GNDA.n350 GNDA.n349 585
R1116 GNDA.n353 GNDA.n352 585
R1117 GNDA.n318 GNDA.n313 585
R1118 GNDA.n316 GNDA.n315 585
R1119 GNDA.n415 GNDA.n414 585
R1120 GNDA.n415 GNDA.n291 585
R1121 GNDA.n1116 GNDA.n274 585
R1122 GNDA.n1151 GNDA.n1150 585
R1123 GNDA.n1148 GNDA.n1118 585
R1124 GNDA.n1146 GNDA.n1145 585
R1125 GNDA.n1140 GNDA.n1119 585
R1126 GNDA.n1135 GNDA.n1134 585
R1127 GNDA.n1132 GNDA.n1120 585
R1128 GNDA.n1130 GNDA.n1129 585
R1129 GNDA.n1124 GNDA.n1122 585
R1130 GNDA.n1094 GNDA.n1093 585
R1131 GNDA.n1208 GNDA.n1207 585
R1132 GNDA.n1211 GNDA.n1210 585
R1133 GNDA.n1477 GNDA.n275 585
R1134 GNDA.n1477 GNDA.n1476 585
R1135 GNDA.n1514 GNDA.n261 585
R1136 GNDA.n1503 GNDA.n260 585
R1137 GNDA.n1504 GNDA.n263 585
R1138 GNDA.n1507 GNDA.n1506 585
R1139 GNDA.n1501 GNDA.n265 585
R1140 GNDA.n1499 GNDA.n1498 585
R1141 GNDA.n267 GNDA.n266 585
R1142 GNDA.n1492 GNDA.n1491 585
R1143 GNDA.n1489 GNDA.n269 585
R1144 GNDA.n1487 GNDA.n1486 585
R1145 GNDA.n271 GNDA.n270 585
R1146 GNDA.n1480 GNDA.n1479 585
R1147 GNDA.n460 GNDA.n275 585
R1148 GNDA.n1476 GNDA.n460 585
R1149 GNDA.n1481 GNDA.n1480 585
R1150 GNDA.n1483 GNDA.n271 585
R1151 GNDA.n1486 GNDA.n1485 585
R1152 GNDA.n269 GNDA.n268 585
R1153 GNDA.n1493 GNDA.n1492 585
R1154 GNDA.n1495 GNDA.n267 585
R1155 GNDA.n1498 GNDA.n1497 585
R1156 GNDA.n265 GNDA.n264 585
R1157 GNDA.n1508 GNDA.n1507 585
R1158 GNDA.n1510 GNDA.n263 585
R1159 GNDA.n1511 GNDA.n260 585
R1160 GNDA.n1514 GNDA.n1513 585
R1161 GNDA.n1048 GNDA.n665 585
R1162 GNDA.n1051 GNDA.n665 585
R1163 GNDA.n1025 GNDA.n812 585
R1164 GNDA.n1026 GNDA.n810 585
R1165 GNDA.n1027 GNDA.n809 585
R1166 GNDA.n807 GNDA.n805 585
R1167 GNDA.n1033 GNDA.n804 585
R1168 GNDA.n1034 GNDA.n802 585
R1169 GNDA.n1035 GNDA.n801 585
R1170 GNDA.n799 GNDA.n797 585
R1171 GNDA.n1040 GNDA.n796 585
R1172 GNDA.n1041 GNDA.n794 585
R1173 GNDA.n793 GNDA.n790 585
R1174 GNDA.n1046 GNDA.n789 585
R1175 GNDA.n1049 GNDA.n1048 585
R1176 GNDA.n1051 GNDA.n1049 585
R1177 GNDA.n1046 GNDA.n1045 585
R1178 GNDA.n1043 GNDA.n790 585
R1179 GNDA.n1042 GNDA.n1041 585
R1180 GNDA.n1040 GNDA.n1039 585
R1181 GNDA.n1038 GNDA.n797 585
R1182 GNDA.n1036 GNDA.n1035 585
R1183 GNDA.n1034 GNDA.n798 585
R1184 GNDA.n1033 GNDA.n1032 585
R1185 GNDA.n1030 GNDA.n805 585
R1186 GNDA.n1028 GNDA.n1027 585
R1187 GNDA.n1026 GNDA.n806 585
R1188 GNDA.n1025 GNDA.n1024 585
R1189 GNDA.n1940 GNDA.n135 585
R1190 GNDA.n1940 GNDA.n1939 585
R1191 GNDA.n1977 GNDA.n1976 585
R1192 GNDA.n1965 GNDA.n101 585
R1193 GNDA.n1966 GNDA.n123 585
R1194 GNDA.n1969 GNDA.n1968 585
R1195 GNDA.n1964 GNDA.n125 585
R1196 GNDA.n1962 GNDA.n1961 585
R1197 GNDA.n127 GNDA.n126 585
R1198 GNDA.n1955 GNDA.n1954 585
R1199 GNDA.n1952 GNDA.n129 585
R1200 GNDA.n1950 GNDA.n1949 585
R1201 GNDA.n131 GNDA.n130 585
R1202 GNDA.n1943 GNDA.n1942 585
R1203 GNDA.n1936 GNDA.n135 585
R1204 GNDA.n1937 GNDA.n1936 585
R1205 GNDA.n1944 GNDA.n1943 585
R1206 GNDA.n1946 GNDA.n131 585
R1207 GNDA.n1949 GNDA.n1948 585
R1208 GNDA.n129 GNDA.n128 585
R1209 GNDA.n1956 GNDA.n1955 585
R1210 GNDA.n1958 GNDA.n127 585
R1211 GNDA.n1961 GNDA.n1960 585
R1212 GNDA.n125 GNDA.n124 585
R1213 GNDA.n1970 GNDA.n1969 585
R1214 GNDA.n1972 GNDA.n123 585
R1215 GNDA.n1973 GNDA.n101 585
R1216 GNDA.n1976 GNDA.n1975 585
R1217 GNDA.n1748 GNDA.n134 585
R1218 GNDA.n136 GNDA.n134 585
R1219 GNDA.n11 GNDA.n8 585
R1220 GNDA.n8 GNDA.n7 585
R1221 GNDA.n2070 GNDA.n2069 585
R1222 GNDA.n2071 GNDA.n2070 585
R1223 GNDA.n9 GNDA.n5 585
R1224 GNDA.n2072 GNDA.n5 585
R1225 GNDA.n2075 GNDA.n2074 585
R1226 GNDA.n2074 GNDA.n2073 585
R1227 GNDA.n13 GNDA.n4 585
R1228 GNDA.n6 GNDA.n4 585
R1229 GNDA.n2057 GNDA.n2056 585
R1230 GNDA.n2056 GNDA.n2055 585
R1231 GNDA.n17 GNDA.n16 585
R1232 GNDA.n18 GNDA.n17 585
R1233 GNDA.n1807 GNDA.n1806 585
R1234 GNDA.n1806 GNDA.n1805 585
R1235 GNDA.n1734 GNDA.n1731 585
R1236 GNDA.n1731 GNDA.n1729 585
R1237 GNDA.n1813 GNDA.n1812 585
R1238 GNDA.n1814 GNDA.n1813 585
R1239 GNDA.n1732 GNDA.n1730 585
R1240 GNDA.n1730 GNDA.n1728 585
R1241 GNDA.n1717 GNDA.n198 585
R1242 GNDA.n1722 GNDA.n198 585
R1243 GNDA.n1720 GNDA.n1719 585
R1244 GNDA.n1721 GNDA.n1720 585
R1245 GNDA.n1638 GNDA.n199 585
R1246 GNDA.n1634 GNDA.n199 585
R1247 GNDA.n1645 GNDA.n1644 585
R1248 GNDA.n1646 GNDA.n1645 585
R1249 GNDA.n1636 GNDA.n1615 585
R1250 GNDA.n1647 GNDA.n1615 585
R1251 GNDA.n1650 GNDA.n1649 585
R1252 GNDA.n1649 GNDA.n1648 585
R1253 GNDA.n1611 GNDA.n1608 585
R1254 GNDA.n1616 GNDA.n1608 585
R1255 GNDA.n1657 GNDA.n1656 585
R1256 GNDA.n1658 GNDA.n1657 585
R1257 GNDA.n1609 GNDA.n222 585
R1258 GNDA.n1659 GNDA.n222 585
R1259 GNDA.n1662 GNDA.n1661 585
R1260 GNDA.n1661 GNDA.n1660 585
R1261 GNDA.n221 GNDA.n219 585
R1262 GNDA.n1607 GNDA.n221 585
R1263 GNDA.n1605 GNDA.n1604 585
R1264 GNDA.n1606 GNDA.n1605 585
R1265 GNDA.n1603 GNDA.n1547 585
R1266 GNDA.n1547 GNDA.n1544 585
R1267 GNDA.n1603 GNDA.n1602 585
R1268 GNDA.n1602 GNDA.n1601 585
R1269 GNDA.n1725 GNDA.n1724 585
R1270 GNDA.n1724 GNDA.n1723 585
R1271 GNDA.n2003 GNDA.n97 585
R1272 GNDA.n2004 GNDA.n95 585
R1273 GNDA.n2007 GNDA.n94 585
R1274 GNDA.n2008 GNDA.n92 585
R1275 GNDA.n2011 GNDA.n91 585
R1276 GNDA.n2012 GNDA.n89 585
R1277 GNDA.n2015 GNDA.n88 585
R1278 GNDA.n2016 GNDA.n86 585
R1279 GNDA.n2019 GNDA.n85 585
R1280 GNDA.n2021 GNDA.n83 585
R1281 GNDA.n2022 GNDA.n82 585
R1282 GNDA.n2023 GNDA.n80 585
R1283 GNDA.n1726 GNDA.n1725 585
R1284 GNDA.n1727 GNDA.n1726 585
R1285 GNDA.n2024 GNDA.n2023 585
R1286 GNDA.n2022 GNDA.n77 585
R1287 GNDA.n2021 GNDA.n2020 585
R1288 GNDA.n2019 GNDA.n2018 585
R1289 GNDA.n2017 GNDA.n2016 585
R1290 GNDA.n2015 GNDA.n2014 585
R1291 GNDA.n2013 GNDA.n2012 585
R1292 GNDA.n2011 GNDA.n2010 585
R1293 GNDA.n2009 GNDA.n2008 585
R1294 GNDA.n2007 GNDA.n2006 585
R1295 GNDA.n2005 GNDA.n2004 585
R1296 GNDA.n2003 GNDA.n2002 585
R1297 GNDA.n1052 GNDA.n664 585
R1298 GNDA.n1052 GNDA.n1051 585
R1299 GNDA.n1089 GNDA.n465 585
R1300 GNDA.n1078 GNDA.n464 585
R1301 GNDA.n1079 GNDA.n467 585
R1302 GNDA.n1082 GNDA.n1081 585
R1303 GNDA.n1076 GNDA.n469 585
R1304 GNDA.n1074 GNDA.n1073 585
R1305 GNDA.n471 GNDA.n470 585
R1306 GNDA.n1067 GNDA.n1066 585
R1307 GNDA.n1064 GNDA.n473 585
R1308 GNDA.n1062 GNDA.n1061 585
R1309 GNDA.n475 GNDA.n474 585
R1310 GNDA.n1055 GNDA.n1054 585
R1311 GNDA.n1050 GNDA.n664 585
R1312 GNDA.n1051 GNDA.n1050 585
R1313 GNDA.n1056 GNDA.n1055 585
R1314 GNDA.n1058 GNDA.n475 585
R1315 GNDA.n1061 GNDA.n1060 585
R1316 GNDA.n473 GNDA.n472 585
R1317 GNDA.n1068 GNDA.n1067 585
R1318 GNDA.n1070 GNDA.n471 585
R1319 GNDA.n1073 GNDA.n1072 585
R1320 GNDA.n469 GNDA.n468 585
R1321 GNDA.n1083 GNDA.n1082 585
R1322 GNDA.n1085 GNDA.n467 585
R1323 GNDA.n1086 GNDA.n464 585
R1324 GNDA.n1089 GNDA.n1088 585
R1325 GNDA.n1474 GNDA.n276 585
R1326 GNDA.n1476 GNDA.n276 585
R1327 GNDA.n1451 GNDA.n1226 585
R1328 GNDA.n1452 GNDA.n1225 585
R1329 GNDA.n1453 GNDA.n1224 585
R1330 GNDA.n1239 GNDA.n1222 585
R1331 GNDA.n1459 GNDA.n1221 585
R1332 GNDA.n1460 GNDA.n1220 585
R1333 GNDA.n1461 GNDA.n1219 585
R1334 GNDA.n1236 GNDA.n1217 585
R1335 GNDA.n1466 GNDA.n1216 585
R1336 GNDA.n1467 GNDA.n1215 585
R1337 GNDA.n1233 GNDA.n1213 585
R1338 GNDA.n1472 GNDA.n1212 585
R1339 GNDA.n1475 GNDA.n1474 585
R1340 GNDA.n1476 GNDA.n1475 585
R1341 GNDA.n1472 GNDA.n1471 585
R1342 GNDA.n1469 GNDA.n1213 585
R1343 GNDA.n1468 GNDA.n1467 585
R1344 GNDA.n1466 GNDA.n1465 585
R1345 GNDA.n1464 GNDA.n1217 585
R1346 GNDA.n1462 GNDA.n1461 585
R1347 GNDA.n1460 GNDA.n1218 585
R1348 GNDA.n1459 GNDA.n1458 585
R1349 GNDA.n1456 GNDA.n1222 585
R1350 GNDA.n1454 GNDA.n1453 585
R1351 GNDA.n1452 GNDA.n1223 585
R1352 GNDA.n1451 GNDA.n1450 585
R1353 GNDA.n1516 GNDA.n258 585
R1354 GNDA.n258 GNDA.n257 585
R1355 GNDA.n1518 GNDA.n1517 585
R1356 GNDA.n1519 GNDA.n1518 585
R1357 GNDA.n256 GNDA.n255 585
R1358 GNDA.n1520 GNDA.n256 585
R1359 GNDA.n1523 GNDA.n1522 585
R1360 GNDA.n1522 GNDA.n1521 585
R1361 GNDA.n1524 GNDA.n252 585
R1362 GNDA.n252 GNDA.n250 585
R1363 GNDA.n1526 GNDA.n1525 585
R1364 GNDA.n1527 GNDA.n1526 585
R1365 GNDA.n1438 GNDA.n251 585
R1366 GNDA.n251 GNDA.n248 585
R1367 GNDA.n1441 GNDA.n1440 585
R1368 GNDA.n1440 GNDA.n1439 585
R1369 GNDA.n1442 GNDA.n1436 585
R1370 GNDA.n1436 GNDA.n1435 585
R1371 GNDA.n1444 GNDA.n1443 585
R1372 GNDA.n1445 GNDA.n1444 585
R1373 GNDA.n1437 GNDA.n1433 585
R1374 GNDA.n1446 GNDA.n1433 585
R1375 GNDA.n1448 GNDA.n1434 585
R1376 GNDA.n1448 GNDA.n1447 585
R1377 GNDA.n245 GNDA.n244 585
R1378 GNDA.n1529 GNDA.n1528 585
R1379 GNDA.n1528 GNDA.t16 585
R1380 GNDA.n1938 GNDA.n68 370.214
R1381 GNDA.n71 GNDA.n70 370.214
R1382 GNDA.n1938 GNDA.n69 365.957
R1383 GNDA.n2026 GNDA.n71 365.957
R1384 GNDA.t16 GNDA.n53 337.541
R1385 GNDA.t16 GNDA.n246 172.876
R1386 GNDA.t16 GNDA.n69 327.661
R1387 GNDA.t16 GNDA.n2026 327.661
R1388 GNDA.t16 GNDA.n62 172.876
R1389 GNDA.t16 GNDA.n64 172.876
R1390 GNDA.t16 GNDA.n56 172.876
R1391 GNDA.t16 GNDA.n1242 172.615
R1392 GNDA.t16 GNDA.n68 323.404
R1393 GNDA.t16 GNDA.n70 323.404
R1394 GNDA.t16 GNDA.n61 172.615
R1395 GNDA.t16 GNDA.n63 172.615
R1396 GNDA.t16 GNDA.n247 172.615
R1397 GNDA.n517 GNDA.t11 305.584
R1398 GNDA.t3 GNDA.t0 297.408
R1399 GNDA.t33 GNDA.n1543 271.354
R1400 GNDA.n413 GNDA.n23 263.904
R1401 GNDA.n980 GNDA.n979 263.904
R1402 GNDA.n2050 GNDA.n22 263.904
R1403 GNDA.n1541 GNDA.t26 260
R1404 GNDA.t26 GNDA.n223 260
R1405 GNDA.t16 GNDA.n249 257.779
R1406 GNDA.n1450 GNDA.n1448 257.466
R1407 GNDA.n2002 GNDA.n2001 257.466
R1408 GNDA.n1088 GNDA.n466 257.466
R1409 GNDA.n1975 GNDA.n122 257.466
R1410 GNDA.n1024 GNDA.n1022 257.466
R1411 GNDA.n1579 GNDA.n1556 257.466
R1412 GNDA.n546 GNDA.n518 257.466
R1413 GNDA.n1406 GNDA.n1250 257.466
R1414 GNDA.n1513 GNDA.n262 257.466
R1415 GNDA.n1000 GNDA.n23 254.34
R1416 GNDA.n994 GNDA.n23 254.34
R1417 GNDA.n992 GNDA.n23 254.34
R1418 GNDA.n986 GNDA.n23 254.34
R1419 GNDA.n984 GNDA.n23 254.34
R1420 GNDA.n978 GNDA.n23 254.34
R1421 GNDA.n32 GNDA.n23 254.34
R1422 GNDA.n2035 GNDA.n23 254.34
R1423 GNDA.n29 GNDA.n23 254.34
R1424 GNDA.n2042 GNDA.n23 254.34
R1425 GNDA.n26 GNDA.n23 254.34
R1426 GNDA.n2049 GNDA.n23 254.34
R1427 GNDA.n478 GNDA.n51 254.34
R1428 GNDA.n481 GNDA.n51 254.34
R1429 GNDA.n639 GNDA.n51 254.34
R1430 GNDA.n630 GNDA.n51 254.34
R1431 GNDA.n649 GNDA.n51 254.34
R1432 GNDA.n625 GNDA.n51 254.34
R1433 GNDA.n785 GNDA.n51 254.34
R1434 GNDA.n775 GNDA.n51 254.34
R1435 GNDA.n673 GNDA.n51 254.34
R1436 GNDA.n761 GNDA.n51 254.34
R1437 GNDA.n677 GNDA.n51 254.34
R1438 GNDA.n748 GNDA.n51 254.34
R1439 GNDA.n975 GNDA.n51 254.34
R1440 GNDA.n889 GNDA.n51 254.34
R1441 GNDA.n904 GNDA.n51 254.34
R1442 GNDA.n887 GNDA.n51 254.34
R1443 GNDA.n915 GNDA.n51 254.34
R1444 GNDA.n881 GNDA.n51 254.34
R1445 GNDA.n2027 GNDA.n50 254.34
R1446 GNDA.n2027 GNDA.n49 254.34
R1447 GNDA.n2027 GNDA.n48 254.34
R1448 GNDA.n2027 GNDA.n47 254.34
R1449 GNDA.n2027 GNDA.n46 254.34
R1450 GNDA.n2027 GNDA.n45 254.34
R1451 GNDA.n2027 GNDA.n44 254.34
R1452 GNDA.n2027 GNDA.n43 254.34
R1453 GNDA.n2027 GNDA.n42 254.34
R1454 GNDA.n2027 GNDA.n41 254.34
R1455 GNDA.n2027 GNDA.n40 254.34
R1456 GNDA.n2027 GNDA.n39 254.34
R1457 GNDA.n2028 GNDA.n2027 254.34
R1458 GNDA.n2027 GNDA.n38 254.34
R1459 GNDA.n2027 GNDA.n37 254.34
R1460 GNDA.n2027 GNDA.n36 254.34
R1461 GNDA.n2027 GNDA.n35 254.34
R1462 GNDA.n2027 GNDA.n34 254.34
R1463 GNDA.n1319 GNDA.n54 254.34
R1464 GNDA.n1316 GNDA.n54 254.34
R1465 GNDA.n1302 GNDA.n54 254.34
R1466 GNDA.n1300 GNDA.n54 254.34
R1467 GNDA.n1290 GNDA.n54 254.34
R1468 GNDA.n1379 GNDA.n54 254.34
R1469 GNDA.n528 GNDA.n65 254.34
R1470 GNDA.n526 GNDA.n65 254.34
R1471 GNDA.n535 GNDA.n65 254.34
R1472 GNDA.n523 GNDA.n65 254.34
R1473 GNDA.n542 GNDA.n65 254.34
R1474 GNDA.n545 GNDA.n65 254.34
R1475 GNDA.n838 GNDA.n65 254.34
R1476 GNDA.n814 GNDA.n65 254.34
R1477 GNDA.n831 GNDA.n65 254.34
R1478 GNDA.n825 GNDA.n65 254.34
R1479 GNDA.n823 GNDA.n65 254.34
R1480 GNDA.n818 GNDA.n65 254.34
R1481 GNDA.n851 GNDA.n65 254.34
R1482 GNDA.n1007 GNDA.n65 254.34
R1483 GNDA.n848 GNDA.n65 254.34
R1484 GNDA.n1014 GNDA.n65 254.34
R1485 GNDA.n845 GNDA.n65 254.34
R1486 GNDA.n1021 GNDA.n65 254.34
R1487 GNDA.n434 GNDA.n23 254.34
R1488 GNDA.n428 GNDA.n23 254.34
R1489 GNDA.n426 GNDA.n23 254.34
R1490 GNDA.n420 GNDA.n23 254.34
R1491 GNDA.n418 GNDA.n23 254.34
R1492 GNDA.n411 GNDA.n54 254.34
R1493 GNDA.n325 GNDA.n54 254.34
R1494 GNDA.n340 GNDA.n54 254.34
R1495 GNDA.n323 GNDA.n54 254.34
R1496 GNDA.n351 GNDA.n54 254.34
R1497 GNDA.n317 GNDA.n54 254.34
R1498 GNDA.n1149 GNDA.n54 254.34
R1499 GNDA.n1147 GNDA.n54 254.34
R1500 GNDA.n1133 GNDA.n54 254.34
R1501 GNDA.n1131 GNDA.n54 254.34
R1502 GNDA.n1121 GNDA.n54 254.34
R1503 GNDA.n1209 GNDA.n54 254.34
R1504 GNDA.n1502 GNDA.n247 254.34
R1505 GNDA.n1505 GNDA.n247 254.34
R1506 GNDA.n1500 GNDA.n247 254.34
R1507 GNDA.n1490 GNDA.n247 254.34
R1508 GNDA.n1488 GNDA.n247 254.34
R1509 GNDA.n1478 GNDA.n247 254.34
R1510 GNDA.n1482 GNDA.n56 254.34
R1511 GNDA.n1484 GNDA.n56 254.34
R1512 GNDA.n1494 GNDA.n56 254.34
R1513 GNDA.n1496 GNDA.n56 254.34
R1514 GNDA.n1509 GNDA.n56 254.34
R1515 GNDA.n1512 GNDA.n56 254.34
R1516 GNDA.n811 GNDA.n61 254.34
R1517 GNDA.n808 GNDA.n61 254.34
R1518 GNDA.n803 GNDA.n61 254.34
R1519 GNDA.n800 GNDA.n61 254.34
R1520 GNDA.n795 GNDA.n61 254.34
R1521 GNDA.n792 GNDA.n61 254.34
R1522 GNDA.n1044 GNDA.n62 254.34
R1523 GNDA.n791 GNDA.n62 254.34
R1524 GNDA.n1037 GNDA.n62 254.34
R1525 GNDA.n1031 GNDA.n62 254.34
R1526 GNDA.n1029 GNDA.n62 254.34
R1527 GNDA.n1023 GNDA.n62 254.34
R1528 GNDA.n100 GNDA.n68 254.34
R1529 GNDA.n1967 GNDA.n68 254.34
R1530 GNDA.n1963 GNDA.n68 254.34
R1531 GNDA.n1953 GNDA.n68 254.34
R1532 GNDA.n1951 GNDA.n68 254.34
R1533 GNDA.n1941 GNDA.n68 254.34
R1534 GNDA.n1945 GNDA.n69 254.34
R1535 GNDA.n1947 GNDA.n69 254.34
R1536 GNDA.n1957 GNDA.n69 254.34
R1537 GNDA.n1959 GNDA.n69 254.34
R1538 GNDA.n1971 GNDA.n69 254.34
R1539 GNDA.n1974 GNDA.n69 254.34
R1540 GNDA.n96 GNDA.n70 254.34
R1541 GNDA.n93 GNDA.n70 254.34
R1542 GNDA.n90 GNDA.n70 254.34
R1543 GNDA.n87 GNDA.n70 254.34
R1544 GNDA.n84 GNDA.n70 254.34
R1545 GNDA.n81 GNDA.n70 254.34
R1546 GNDA.n2026 GNDA.n2025 254.34
R1547 GNDA.n2026 GNDA.n76 254.34
R1548 GNDA.n2026 GNDA.n75 254.34
R1549 GNDA.n2026 GNDA.n74 254.34
R1550 GNDA.n2026 GNDA.n73 254.34
R1551 GNDA.n2026 GNDA.n72 254.34
R1552 GNDA.n1077 GNDA.n63 254.34
R1553 GNDA.n1080 GNDA.n63 254.34
R1554 GNDA.n1075 GNDA.n63 254.34
R1555 GNDA.n1065 GNDA.n63 254.34
R1556 GNDA.n1063 GNDA.n63 254.34
R1557 GNDA.n1053 GNDA.n63 254.34
R1558 GNDA.n1057 GNDA.n64 254.34
R1559 GNDA.n1059 GNDA.n64 254.34
R1560 GNDA.n1069 GNDA.n64 254.34
R1561 GNDA.n1071 GNDA.n64 254.34
R1562 GNDA.n1084 GNDA.n64 254.34
R1563 GNDA.n1087 GNDA.n64 254.34
R1564 GNDA.n1242 GNDA.n1241 254.34
R1565 GNDA.n1242 GNDA.n1240 254.34
R1566 GNDA.n1242 GNDA.n1238 254.34
R1567 GNDA.n1242 GNDA.n1237 254.34
R1568 GNDA.n1242 GNDA.n1235 254.34
R1569 GNDA.n1242 GNDA.n1234 254.34
R1570 GNDA.n1470 GNDA.n246 254.34
R1571 GNDA.n1214 GNDA.n246 254.34
R1572 GNDA.n1463 GNDA.n246 254.34
R1573 GNDA.n1457 GNDA.n246 254.34
R1574 GNDA.n1455 GNDA.n246 254.34
R1575 GNDA.n1449 GNDA.n246 254.34
R1576 GNDA.n261 GNDA.n258 251.614
R1577 GNDA.n1978 GNDA.n1977 251.614
R1578 GNDA.n839 GNDA.n812 251.614
R1579 GNDA.n2030 GNDA.n2029 251.614
R1580 GNDA.n1002 GNDA.n1001 251.614
R1581 GNDA.n1557 GNDA.n97 251.614
R1582 GNDA.n527 GNDA.n465 251.614
R1583 GNDA.n1430 GNDA.n1226 251.614
R1584 GNDA.n437 GNDA.n436 251.614
R1585 GNDA.n1817 GNDA.n1816 250.349
R1586 GNDA.n1827 GNDA.n1826 250.349
R1587 GNDA.n184 GNDA.n183 246.25
R1588 GNDA.n1848 GNDA.n183 246.25
R1589 GNDA.n1619 GNDA.n1618 246.25
R1590 GNDA.n1623 GNDA.n1618 246.25
R1591 GNDA.n1543 GNDA.n1542 241.643
R1592 GNDA.n1633 GNDA.n1632 241.643
R1593 GNDA.n1633 GNDA.n1617 241.643
R1594 GNDA.n1855 GNDA.n1854 241.643
R1595 GNDA.n1855 GNDA.n182 241.643
R1596 GNDA.t16 GNDA.n52 221.698
R1597 GNDA.n1715 GNDA.n202 221.667
R1598 GNDA.n1154 GNDA.n1153 221.667
R1599 GNDA.n781 GNDA.n670 221.667
R1600 GNDA.n1878 GNDA.n1877 221.667
R1601 GNDA.n970 GNDA.n861 221.667
R1602 GNDA.n493 GNDA.n484 221.667
R1603 GNDA.n1324 GNDA.n1323 221.667
R1604 GNDA.n406 GNDA.n296 221.667
R1605 GNDA.n2067 GNDA.n12 221.667
R1606 GNDA.n23 GNDA.t6 217.377
R1607 GNDA.n1828 GNDA.n1825 197
R1608 GNDA.n1818 GNDA.n197 197
R1609 GNDA.n1210 GNDA.n461 195.049
R1610 GNDA.n1730 GNDA.n78 195.049
R1611 GNDA.n747 GNDA.n476 195.049
R1612 GNDA.n1934 GNDA.n132 195.049
R1613 GNDA.n880 GNDA.n666 195.049
R1614 GNDA.n1605 GNDA.n1545 195.049
R1615 GNDA.n624 GNDA.n507 195.049
R1616 GNDA.n1381 GNDA.n1380 195.049
R1617 GNDA.n316 GNDA.n272 195.049
R1618 GNDA.n1447 GNDA.t16 187.726
R1619 GNDA.t16 GNDA.n459 187.726
R1620 GNDA.n1477 GNDA.n274 187.249
R1621 GNDA.n1940 GNDA.n134 187.249
R1622 GNDA.n786 GNDA.n665 187.249
R1623 GNDA.n2051 GNDA.n21 187.249
R1624 GNDA.n977 GNDA.n976 187.249
R1625 GNDA.n1724 GNDA.n198 187.249
R1626 GNDA.n1052 GNDA.n663 187.249
R1627 GNDA.n1318 GNDA.n276 187.249
R1628 GNDA.n414 GNDA.n412 187.249
R1629 GNDA.n1701 GNDA.n207 185
R1630 GNDA.n1703 GNDA.n1702 185
R1631 GNDA.n1705 GNDA.n205 185
R1632 GNDA.n1707 GNDA.n1706 185
R1633 GNDA.n1708 GNDA.n204 185
R1634 GNDA.n1710 GNDA.n1709 185
R1635 GNDA.n1712 GNDA.n203 185
R1636 GNDA.n1713 GNDA.n201 185
R1637 GNDA.n1716 GNDA.n1715 185
R1638 GNDA.n1700 GNDA.n1699 185
R1639 GNDA.n1697 GNDA.n208 185
R1640 GNDA.n1697 GNDA.t20 185
R1641 GNDA.n1696 GNDA.n209 185
R1642 GNDA.n1694 GNDA.n1693 185
R1643 GNDA.n1692 GNDA.n210 185
R1644 GNDA.n1691 GNDA.n1690 185
R1645 GNDA.n1688 GNDA.n211 185
R1646 GNDA.n1686 GNDA.n1685 185
R1647 GNDA.n1684 GNDA.n212 185
R1648 GNDA.n1667 GNDA.n1666 185
R1649 GNDA.n1668 GNDA.n216 185
R1650 GNDA.n1670 GNDA.n1669 185
R1651 GNDA.n1672 GNDA.n215 185
R1652 GNDA.n1675 GNDA.n1674 185
R1653 GNDA.n1676 GNDA.n214 185
R1654 GNDA.n1678 GNDA.n1677 185
R1655 GNDA.n1680 GNDA.n213 185
R1656 GNDA.n1683 GNDA.n1682 185
R1657 GNDA.n1171 GNDA.n1170 185
R1658 GNDA.n1169 GNDA.n1168 185
R1659 GNDA.n1167 GNDA.n1166 185
R1660 GNDA.n1165 GNDA.n1164 185
R1661 GNDA.n1163 GNDA.n1162 185
R1662 GNDA.n1161 GNDA.n1160 185
R1663 GNDA.n1159 GNDA.n1158 185
R1664 GNDA.n1157 GNDA.n1156 185
R1665 GNDA.n1155 GNDA.n1154 185
R1666 GNDA.n1173 GNDA.n1172 185
R1667 GNDA.n1174 GNDA.n1104 185
R1668 GNDA.t23 GNDA.n1104 185
R1669 GNDA.n1176 GNDA.n1175 185
R1670 GNDA.n1178 GNDA.n1177 185
R1671 GNDA.n1180 GNDA.n1179 185
R1672 GNDA.n1182 GNDA.n1181 185
R1673 GNDA.n1184 GNDA.n1183 185
R1674 GNDA.n1186 GNDA.n1185 185
R1675 GNDA.n1188 GNDA.n1187 185
R1676 GNDA.n1115 GNDA.n1095 185
R1677 GNDA.n1203 GNDA.n1202 185
R1678 GNDA.n1201 GNDA.n1114 185
R1679 GNDA.n1200 GNDA.n1199 185
R1680 GNDA.n1198 GNDA.n1197 185
R1681 GNDA.n1196 GNDA.n1195 185
R1682 GNDA.n1194 GNDA.n1193 185
R1683 GNDA.n1192 GNDA.n1191 185
R1684 GNDA.n1190 GNDA.n1189 185
R1685 GNDA.n708 GNDA.n688 185
R1686 GNDA.n707 GNDA.n706 185
R1687 GNDA.n705 GNDA.n704 185
R1688 GNDA.n703 GNDA.n690 185
R1689 GNDA.n701 GNDA.n700 185
R1690 GNDA.n699 GNDA.n691 185
R1691 GNDA.n698 GNDA.n697 185
R1692 GNDA.n695 GNDA.n693 185
R1693 GNDA.n692 GNDA.n670 185
R1694 GNDA.n711 GNDA.n710 185
R1695 GNDA.n712 GNDA.n687 185
R1696 GNDA.n687 GNDA.t17 185
R1697 GNDA.n714 GNDA.n713 185
R1698 GNDA.n716 GNDA.n686 185
R1699 GNDA.n719 GNDA.n718 185
R1700 GNDA.n720 GNDA.n685 185
R1701 GNDA.n722 GNDA.n721 185
R1702 GNDA.n724 GNDA.n684 185
R1703 GNDA.n727 GNDA.n726 185
R1704 GNDA.n744 GNDA.n679 185
R1705 GNDA.n743 GNDA.n742 185
R1706 GNDA.n740 GNDA.n680 185
R1707 GNDA.n738 GNDA.n737 185
R1708 GNDA.n736 GNDA.n681 185
R1709 GNDA.n735 GNDA.n734 185
R1710 GNDA.n732 GNDA.n682 185
R1711 GNDA.n730 GNDA.n729 185
R1712 GNDA.n728 GNDA.n683 185
R1713 GNDA.n782 GNDA.n781 185
R1714 GNDA.n779 GNDA.n778 185
R1715 GNDA.n672 GNDA.n671 185
R1716 GNDA.n772 GNDA.n771 185
R1717 GNDA.n769 GNDA.n674 185
R1718 GNDA.n767 GNDA.n766 185
R1719 GNDA.n757 GNDA.n675 185
R1720 GNDA.n756 GNDA.n755 185
R1721 GNDA.n753 GNDA.n752 185
R1722 GNDA.n753 GNDA.t17 185
R1723 GNDA.n1853 GNDA.n1852 185
R1724 GNDA.n1852 GNDA.n1851 185
R1725 GNDA.n1846 GNDA.n185 185
R1726 GNDA.n1853 GNDA.n185 185
R1727 GNDA.n1631 GNDA.n1630 185
R1728 GNDA.n1628 GNDA.n1627 185
R1729 GNDA.n1895 GNDA.n1894 185
R1730 GNDA.n1893 GNDA.n1892 185
R1731 GNDA.n1891 GNDA.n1890 185
R1732 GNDA.n1889 GNDA.n1888 185
R1733 GNDA.n1887 GNDA.n1886 185
R1734 GNDA.n1885 GNDA.n1884 185
R1735 GNDA.n1883 GNDA.n1882 185
R1736 GNDA.n1881 GNDA.n1880 185
R1737 GNDA.n1879 GNDA.n1878 185
R1738 GNDA.n1897 GNDA.n1896 185
R1739 GNDA.n1898 GNDA.n150 185
R1740 GNDA.t24 GNDA.n150 185
R1741 GNDA.n1900 GNDA.n1899 185
R1742 GNDA.n1902 GNDA.n1901 185
R1743 GNDA.n1904 GNDA.n1903 185
R1744 GNDA.n1906 GNDA.n1905 185
R1745 GNDA.n1908 GNDA.n1907 185
R1746 GNDA.n1910 GNDA.n1909 185
R1747 GNDA.n1912 GNDA.n1911 185
R1748 GNDA.n141 GNDA.n139 185
R1749 GNDA.n1927 GNDA.n1926 185
R1750 GNDA.n1925 GNDA.n160 185
R1751 GNDA.n1924 GNDA.n1923 185
R1752 GNDA.n1922 GNDA.n1921 185
R1753 GNDA.n1920 GNDA.n1919 185
R1754 GNDA.n1918 GNDA.n1917 185
R1755 GNDA.n1916 GNDA.n1915 185
R1756 GNDA.n1914 GNDA.n1913 185
R1757 GNDA.n1877 GNDA.n1876 185
R1758 GNDA.n1868 GNDA.n1867 185
R1759 GNDA.n1866 GNDA.n1865 185
R1760 GNDA.n1863 GNDA.n1862 185
R1761 GNDA.n1861 GNDA.n1860 185
R1762 GNDA.n177 GNDA.n176 185
R1763 GNDA.n175 GNDA.n174 185
R1764 GNDA.n172 GNDA.n142 185
R1765 GNDA.n1930 GNDA.n1929 185
R1766 GNDA.n1929 GNDA.t24 185
R1767 GNDA.n956 GNDA.n866 185
R1768 GNDA.n958 GNDA.n957 185
R1769 GNDA.n960 GNDA.n864 185
R1770 GNDA.n962 GNDA.n961 185
R1771 GNDA.n963 GNDA.n863 185
R1772 GNDA.n965 GNDA.n964 185
R1773 GNDA.n967 GNDA.n862 185
R1774 GNDA.n968 GNDA.n860 185
R1775 GNDA.n971 GNDA.n970 185
R1776 GNDA.n955 GNDA.n954 185
R1777 GNDA.n952 GNDA.n867 185
R1778 GNDA.n952 GNDA.t19 185
R1779 GNDA.n951 GNDA.n868 185
R1780 GNDA.n949 GNDA.n948 185
R1781 GNDA.n947 GNDA.n869 185
R1782 GNDA.n946 GNDA.n945 185
R1783 GNDA.n943 GNDA.n870 185
R1784 GNDA.n941 GNDA.n940 185
R1785 GNDA.n939 GNDA.n871 185
R1786 GNDA.n922 GNDA.n921 185
R1787 GNDA.n923 GNDA.n875 185
R1788 GNDA.n925 GNDA.n924 185
R1789 GNDA.n927 GNDA.n874 185
R1790 GNDA.n930 GNDA.n929 185
R1791 GNDA.n931 GNDA.n873 185
R1792 GNDA.n933 GNDA.n932 185
R1793 GNDA.n935 GNDA.n872 185
R1794 GNDA.n938 GNDA.n937 185
R1795 GNDA.n861 GNDA.n859 185
R1796 GNDA.n895 GNDA.n894 185
R1797 GNDA.n901 GNDA.n900 185
R1798 GNDA.n898 GNDA.n897 185
R1799 GNDA.n896 GNDA.n886 185
R1800 GNDA.n909 GNDA.n908 185
R1801 GNDA.n912 GNDA.n911 185
R1802 GNDA.n879 GNDA.n877 185
R1803 GNDA.n919 GNDA.n918 185
R1804 GNDA.n919 GNDA.t19 185
R1805 GNDA.n587 GNDA.n586 185
R1806 GNDA.n585 GNDA.n584 185
R1807 GNDA.n583 GNDA.n582 185
R1808 GNDA.n581 GNDA.n580 185
R1809 GNDA.n579 GNDA.n578 185
R1810 GNDA.n577 GNDA.n576 185
R1811 GNDA.n575 GNDA.n574 185
R1812 GNDA.n573 GNDA.n572 185
R1813 GNDA.n493 GNDA.n479 185
R1814 GNDA.n589 GNDA.n588 185
R1815 GNDA.n590 GNDA.n491 185
R1816 GNDA.t15 GNDA.n491 185
R1817 GNDA.n592 GNDA.n591 185
R1818 GNDA.n594 GNDA.n593 185
R1819 GNDA.n596 GNDA.n595 185
R1820 GNDA.n598 GNDA.n597 185
R1821 GNDA.n600 GNDA.n599 185
R1822 GNDA.n602 GNDA.n601 185
R1823 GNDA.n604 GNDA.n603 185
R1824 GNDA.n621 GNDA.n503 185
R1825 GNDA.n620 GNDA.n619 185
R1826 GNDA.n618 GNDA.n617 185
R1827 GNDA.n616 GNDA.n615 185
R1828 GNDA.n614 GNDA.n613 185
R1829 GNDA.n612 GNDA.n611 185
R1830 GNDA.n610 GNDA.n609 185
R1831 GNDA.n608 GNDA.n607 185
R1832 GNDA.n606 GNDA.n605 185
R1833 GNDA.n484 GNDA.n480 185
R1834 GNDA.n656 GNDA.n655 185
R1835 GNDA.n636 GNDA.n483 185
R1836 GNDA.n635 GNDA.n634 185
R1837 GNDA.n633 GNDA.n629 185
R1838 GNDA.n644 GNDA.n643 185
R1839 GNDA.n646 GNDA.n645 185
R1840 GNDA.n506 GNDA.n504 185
R1841 GNDA.n653 GNDA.n652 185
R1842 GNDA.t15 GNDA.n653 185
R1843 GNDA.n1341 GNDA.n1340 185
R1844 GNDA.n1339 GNDA.n1338 185
R1845 GNDA.n1337 GNDA.n1336 185
R1846 GNDA.n1335 GNDA.n1334 185
R1847 GNDA.n1333 GNDA.n1332 185
R1848 GNDA.n1331 GNDA.n1330 185
R1849 GNDA.n1329 GNDA.n1328 185
R1850 GNDA.n1327 GNDA.n1326 185
R1851 GNDA.n1325 GNDA.n1324 185
R1852 GNDA.n1343 GNDA.n1342 185
R1853 GNDA.n1344 GNDA.n1274 185
R1854 GNDA.t21 GNDA.n1274 185
R1855 GNDA.n1346 GNDA.n1345 185
R1856 GNDA.n1348 GNDA.n1347 185
R1857 GNDA.n1350 GNDA.n1349 185
R1858 GNDA.n1352 GNDA.n1351 185
R1859 GNDA.n1354 GNDA.n1353 185
R1860 GNDA.n1356 GNDA.n1355 185
R1861 GNDA.n1358 GNDA.n1357 185
R1862 GNDA.n1285 GNDA.n1265 185
R1863 GNDA.n1373 GNDA.n1372 185
R1864 GNDA.n1371 GNDA.n1284 185
R1865 GNDA.n1370 GNDA.n1369 185
R1866 GNDA.n1368 GNDA.n1367 185
R1867 GNDA.n1366 GNDA.n1365 185
R1868 GNDA.n1364 GNDA.n1363 185
R1869 GNDA.n1362 GNDA.n1361 185
R1870 GNDA.n1360 GNDA.n1359 185
R1871 GNDA.n1323 GNDA.n1322 185
R1872 GNDA.n1313 GNDA.n1312 185
R1873 GNDA.n1311 GNDA.n1310 185
R1874 GNDA.n1308 GNDA.n1307 185
R1875 GNDA.n1306 GNDA.n1305 185
R1876 GNDA.n1297 GNDA.n1296 185
R1877 GNDA.n1295 GNDA.n1294 185
R1878 GNDA.n1292 GNDA.n1266 185
R1879 GNDA.n1376 GNDA.n1375 185
R1880 GNDA.n1375 GNDA.t21 185
R1881 GNDA.n392 GNDA.n301 185
R1882 GNDA.n394 GNDA.n393 185
R1883 GNDA.n396 GNDA.n299 185
R1884 GNDA.n398 GNDA.n397 185
R1885 GNDA.n399 GNDA.n298 185
R1886 GNDA.n401 GNDA.n400 185
R1887 GNDA.n403 GNDA.n297 185
R1888 GNDA.n404 GNDA.n295 185
R1889 GNDA.n407 GNDA.n406 185
R1890 GNDA.n391 GNDA.n390 185
R1891 GNDA.n388 GNDA.n302 185
R1892 GNDA.n388 GNDA.t18 185
R1893 GNDA.n387 GNDA.n303 185
R1894 GNDA.n385 GNDA.n384 185
R1895 GNDA.n383 GNDA.n304 185
R1896 GNDA.n382 GNDA.n381 185
R1897 GNDA.n379 GNDA.n305 185
R1898 GNDA.n377 GNDA.n376 185
R1899 GNDA.n375 GNDA.n306 185
R1900 GNDA.n358 GNDA.n357 185
R1901 GNDA.n359 GNDA.n310 185
R1902 GNDA.n361 GNDA.n360 185
R1903 GNDA.n363 GNDA.n309 185
R1904 GNDA.n366 GNDA.n365 185
R1905 GNDA.n367 GNDA.n308 185
R1906 GNDA.n369 GNDA.n368 185
R1907 GNDA.n371 GNDA.n307 185
R1908 GNDA.n374 GNDA.n373 185
R1909 GNDA.n296 GNDA.n294 185
R1910 GNDA.n331 GNDA.n330 185
R1911 GNDA.n337 GNDA.n336 185
R1912 GNDA.n334 GNDA.n333 185
R1913 GNDA.n332 GNDA.n322 185
R1914 GNDA.n345 GNDA.n344 185
R1915 GNDA.n348 GNDA.n347 185
R1916 GNDA.n314 GNDA.n312 185
R1917 GNDA.n355 GNDA.n354 185
R1918 GNDA.n355 GNDA.t18 185
R1919 GNDA.n1153 GNDA.n1152 185
R1920 GNDA.n1144 GNDA.n1143 185
R1921 GNDA.n1142 GNDA.n1141 185
R1922 GNDA.n1139 GNDA.n1138 185
R1923 GNDA.n1137 GNDA.n1136 185
R1924 GNDA.n1128 GNDA.n1127 185
R1925 GNDA.n1126 GNDA.n1125 185
R1926 GNDA.n1123 GNDA.n1096 185
R1927 GNDA.n1206 GNDA.n1205 185
R1928 GNDA.n1205 GNDA.t23 185
R1929 GNDA.n1766 GNDA.n1744 185
R1930 GNDA.n1765 GNDA.n1764 185
R1931 GNDA.n1763 GNDA.n1762 185
R1932 GNDA.n1761 GNDA.n1746 185
R1933 GNDA.n1759 GNDA.n1758 185
R1934 GNDA.n1757 GNDA.n1747 185
R1935 GNDA.n1756 GNDA.n1755 185
R1936 GNDA.n1753 GNDA.n1751 185
R1937 GNDA.n1750 GNDA.n12 185
R1938 GNDA.n1769 GNDA.n1768 185
R1939 GNDA.n1770 GNDA.n1743 185
R1940 GNDA.n1743 GNDA.t22 185
R1941 GNDA.n1772 GNDA.n1771 185
R1942 GNDA.n1774 GNDA.n1742 185
R1943 GNDA.n1777 GNDA.n1776 185
R1944 GNDA.n1778 GNDA.n1741 185
R1945 GNDA.n1780 GNDA.n1779 185
R1946 GNDA.n1782 GNDA.n1740 185
R1947 GNDA.n1785 GNDA.n1784 185
R1948 GNDA.n1802 GNDA.n1801 185
R1949 GNDA.n1800 GNDA.n1799 185
R1950 GNDA.n1798 GNDA.n1736 185
R1951 GNDA.n1796 GNDA.n1795 185
R1952 GNDA.n1794 GNDA.n1737 185
R1953 GNDA.n1793 GNDA.n1792 185
R1954 GNDA.n1790 GNDA.n1738 185
R1955 GNDA.n1788 GNDA.n1787 185
R1956 GNDA.n1786 GNDA.n1739 185
R1957 GNDA.n2068 GNDA.n2067 185
R1958 GNDA.n2065 GNDA.n10 185
R1959 GNDA.n2064 GNDA.n3 185
R1960 GNDA.n2062 GNDA.n2 185
R1961 GNDA.n2061 GNDA.n14 185
R1962 GNDA.n2059 GNDA.n2058 185
R1963 GNDA.n1804 GNDA.n15 185
R1964 GNDA.n1809 GNDA.n1808 185
R1965 GNDA.n1811 GNDA.n1810 185
R1966 GNDA.n1810 GNDA.t22 185
R1967 GNDA.n202 GNDA.n200 185
R1968 GNDA.n1643 GNDA.n1642 185
R1969 GNDA.n1640 GNDA.n1637 185
R1970 GNDA.n1635 GNDA.n1614 185
R1971 GNDA.n1652 GNDA.n1651 185
R1972 GNDA.n1655 GNDA.n1654 185
R1973 GNDA.n1613 GNDA.n1610 185
R1974 GNDA.n220 GNDA.n218 185
R1975 GNDA.n1664 GNDA.n1663 185
R1976 GNDA.n1664 GNDA.t20 185
R1977 GNDA.n1429 GNDA.t16 183.71
R1978 GNDA.t16 GNDA.n257 183.71
R1979 GNDA.n1601 GNDA.n1600 179.756
R1980 GNDA.n1600 GNDA.n1599 179.756
R1981 GNDA.n1599 GNDA.n1549 179.756
R1982 GNDA.n1593 GNDA.n1549 179.756
R1983 GNDA.n1593 GNDA.n66 179.756
R1984 GNDA.n1555 GNDA.n67 179.756
R1985 GNDA.n1586 GNDA.n1555 179.756
R1986 GNDA.n1586 GNDA.n1585 179.756
R1987 GNDA.n1585 GNDA.n1584 179.756
R1988 GNDA.n1584 GNDA.n53 179.756
R1989 GNDA.n568 GNDA.n52 179.756
R1990 GNDA.n568 GNDA.n567 179.756
R1991 GNDA.n567 GNDA.n566 179.756
R1992 GNDA.n566 GNDA.n510 179.756
R1993 GNDA.n560 GNDA.n510 179.756
R1994 GNDA.n560 GNDA.n59 179.756
R1995 GNDA.n516 GNDA.n60 179.756
R1996 GNDA.n553 GNDA.n516 179.756
R1997 GNDA.n553 GNDA.n552 179.756
R1998 GNDA.n552 GNDA.n551 179.756
R1999 GNDA.n551 GNDA.n517 179.756
R2000 GNDA.n1382 GNDA.n1259 179.756
R2001 GNDA.n1387 GNDA.n1259 179.756
R2002 GNDA.n1388 GNDA.n1387 179.756
R2003 GNDA.n1390 GNDA.n1388 179.756
R2004 GNDA.n1390 GNDA.n1389 179.756
R2005 GNDA.n1389 GNDA.n1243 179.756
R2006 GNDA.n1397 GNDA.n1244 179.756
R2007 GNDA.n1397 GNDA.n1253 179.756
R2008 GNDA.n1403 GNDA.n1253 179.756
R2009 GNDA.n1404 GNDA.n1403 179.756
R2010 GNDA.n1405 GNDA.n1404 179.756
R2011 GNDA.n1487 GNDA.n270 175.546
R2012 GNDA.n1491 GNDA.n1489 175.546
R2013 GNDA.n1499 GNDA.n266 175.546
R2014 GNDA.n1506 GNDA.n1501 175.546
R2015 GNDA.n1504 GNDA.n1503 175.546
R2016 GNDA.n1448 GNDA.n1433 175.546
R2017 GNDA.n1444 GNDA.n1433 175.546
R2018 GNDA.n1444 GNDA.n1436 175.546
R2019 GNDA.n1440 GNDA.n1436 175.546
R2020 GNDA.n1440 GNDA.n251 175.546
R2021 GNDA.n1526 GNDA.n251 175.546
R2022 GNDA.n1526 GNDA.n252 175.546
R2023 GNDA.n1522 GNDA.n252 175.546
R2024 GNDA.n1522 GNDA.n256 175.546
R2025 GNDA.n1518 GNDA.n256 175.546
R2026 GNDA.n1518 GNDA.n258 175.546
R2027 GNDA.n1469 GNDA.n1468 175.546
R2028 GNDA.n1465 GNDA.n1464 175.546
R2029 GNDA.n1462 GNDA.n1218 175.546
R2030 GNDA.n1458 GNDA.n1456 175.546
R2031 GNDA.n1454 GNDA.n1223 175.546
R2032 GNDA.n1208 GNDA.n1093 175.546
R2033 GNDA.n1130 GNDA.n1122 175.546
R2034 GNDA.n1134 GNDA.n1132 175.546
R2035 GNDA.n1146 GNDA.n1119 175.546
R2036 GNDA.n1150 GNDA.n1148 175.546
R2037 GNDA.n2020 GNDA.n77 175.546
R2038 GNDA.n2018 GNDA.n2017 175.546
R2039 GNDA.n2014 GNDA.n2013 175.546
R2040 GNDA.n2010 GNDA.n2009 175.546
R2041 GNDA.n2006 GNDA.n2005 175.546
R2042 GNDA.n1813 GNDA.n1730 175.546
R2043 GNDA.n1813 GNDA.n1731 175.546
R2044 GNDA.n1806 GNDA.n1731 175.546
R2045 GNDA.n1806 GNDA.n17 175.546
R2046 GNDA.n2056 GNDA.n17 175.546
R2047 GNDA.n2056 GNDA.n4 175.546
R2048 GNDA.n2074 GNDA.n4 175.546
R2049 GNDA.n2074 GNDA.n5 175.546
R2050 GNDA.n2070 GNDA.n5 175.546
R2051 GNDA.n2070 GNDA.n8 175.546
R2052 GNDA.n134 GNDA.n8 175.546
R2053 GNDA.n1950 GNDA.n130 175.546
R2054 GNDA.n1954 GNDA.n1952 175.546
R2055 GNDA.n1962 GNDA.n126 175.546
R2056 GNDA.n1968 GNDA.n1964 175.546
R2057 GNDA.n1966 GNDA.n1965 175.546
R2058 GNDA.n1998 GNDA.n1997 175.546
R2059 GNDA.n1994 GNDA.n1993 175.546
R2060 GNDA.n1990 GNDA.n1989 175.546
R2061 GNDA.n1986 GNDA.n1985 175.546
R2062 GNDA.n1982 GNDA.n1981 175.546
R2063 GNDA.n794 GNDA.n793 175.546
R2064 GNDA.n799 GNDA.n796 175.546
R2065 GNDA.n802 GNDA.n801 175.546
R2066 GNDA.n807 GNDA.n804 175.546
R2067 GNDA.n810 GNDA.n809 175.546
R2068 GNDA.n822 GNDA.n819 175.546
R2069 GNDA.n826 GNDA.n824 175.546
R2070 GNDA.n830 GNDA.n816 175.546
R2071 GNDA.n833 GNDA.n832 175.546
R2072 GNDA.n837 GNDA.n836 175.546
R2073 GNDA.n1060 GNDA.n1058 175.546
R2074 GNDA.n1068 GNDA.n472 175.546
R2075 GNDA.n1072 GNDA.n1070 175.546
R2076 GNDA.n1083 GNDA.n468 175.546
R2077 GNDA.n1086 GNDA.n1085 175.546
R2078 GNDA.n750 GNDA.n749 175.546
R2079 GNDA.n760 GNDA.n759 175.546
R2080 GNDA.n764 GNDA.n763 175.546
R2081 GNDA.n776 GNDA.n774 175.546
R2082 GNDA.n784 GNDA.n668 175.546
R2083 GNDA.n1934 GNDA.n138 175.546
R2084 GNDA.n170 GNDA.n138 175.546
R2085 GNDA.n171 GNDA.n170 175.546
R2086 GNDA.n179 GNDA.n171 175.546
R2087 GNDA.n179 GNDA.n167 175.546
R2088 GNDA.n1858 GNDA.n167 175.546
R2089 GNDA.n1858 GNDA.n165 175.546
R2090 GNDA.n1870 GNDA.n165 175.546
R2091 GNDA.n1870 GNDA.n164 175.546
R2092 GNDA.n1874 GNDA.n164 175.546
R2093 GNDA.n1874 GNDA.n21 175.546
R2094 GNDA.n1948 GNDA.n1946 175.546
R2095 GNDA.n1956 GNDA.n128 175.546
R2096 GNDA.n1960 GNDA.n1958 175.546
R2097 GNDA.n1970 GNDA.n124 175.546
R2098 GNDA.n1973 GNDA.n1972 175.546
R2099 GNDA.n119 GNDA.n118 175.546
R2100 GNDA.n115 GNDA.n114 175.546
R2101 GNDA.n111 GNDA.n110 175.546
R2102 GNDA.n107 GNDA.n106 175.546
R2103 GNDA.n103 GNDA.n33 175.546
R2104 GNDA.n2048 GNDA.n24 175.546
R2105 GNDA.n2044 GNDA.n2043 175.546
R2106 GNDA.n2041 GNDA.n27 175.546
R2107 GNDA.n2037 GNDA.n2036 175.546
R2108 GNDA.n2034 GNDA.n30 175.546
R2109 GNDA.n983 GNDA.n856 175.546
R2110 GNDA.n987 GNDA.n985 175.546
R2111 GNDA.n991 GNDA.n854 175.546
R2112 GNDA.n995 GNDA.n993 175.546
R2113 GNDA.n999 GNDA.n852 175.546
R2114 GNDA.n1020 GNDA.n843 175.546
R2115 GNDA.n1016 GNDA.n1015 175.546
R2116 GNDA.n1013 GNDA.n846 175.546
R2117 GNDA.n1009 GNDA.n1008 175.546
R2118 GNDA.n1006 GNDA.n849 175.546
R2119 GNDA.n1043 GNDA.n1042 175.546
R2120 GNDA.n1039 GNDA.n1038 175.546
R2121 GNDA.n1036 GNDA.n798 175.546
R2122 GNDA.n1032 GNDA.n1030 175.546
R2123 GNDA.n1028 GNDA.n806 175.546
R2124 GNDA.n916 GNDA.n882 175.546
R2125 GNDA.n914 GNDA.n883 175.546
R2126 GNDA.n906 GNDA.n905 175.546
R2127 GNDA.n903 GNDA.n890 175.546
R2128 GNDA.n974 GNDA.n858 175.546
R2129 GNDA.n1605 GNDA.n221 175.546
R2130 GNDA.n1661 GNDA.n221 175.546
R2131 GNDA.n1661 GNDA.n222 175.546
R2132 GNDA.n1657 GNDA.n222 175.546
R2133 GNDA.n1657 GNDA.n1608 175.546
R2134 GNDA.n1649 GNDA.n1608 175.546
R2135 GNDA.n1649 GNDA.n1615 175.546
R2136 GNDA.n1645 GNDA.n1615 175.546
R2137 GNDA.n1645 GNDA.n199 175.546
R2138 GNDA.n1720 GNDA.n199 175.546
R2139 GNDA.n1720 GNDA.n198 175.546
R2140 GNDA.n83 GNDA.n82 175.546
R2141 GNDA.n86 GNDA.n85 175.546
R2142 GNDA.n89 GNDA.n88 175.546
R2143 GNDA.n92 GNDA.n91 175.546
R2144 GNDA.n95 GNDA.n94 175.546
R2145 GNDA.n1577 GNDA.n1576 175.546
R2146 GNDA.n1573 GNDA.n1572 175.546
R2147 GNDA.n1569 GNDA.n1568 175.546
R2148 GNDA.n1565 GNDA.n1564 175.546
R2149 GNDA.n1561 GNDA.n1560 175.546
R2150 GNDA.n1602 GNDA.n1548 175.546
R2151 GNDA.n1598 GNDA.n1548 175.546
R2152 GNDA.n1598 GNDA.n1550 175.546
R2153 GNDA.n1594 GNDA.n1550 175.546
R2154 GNDA.n1594 GNDA.n1592 175.546
R2155 GNDA.n1592 GNDA.n1591 175.546
R2156 GNDA.n1591 GNDA.n1552 175.546
R2157 GNDA.n1587 GNDA.n1552 175.546
R2158 GNDA.n1587 GNDA.n1554 175.546
R2159 GNDA.n1583 GNDA.n1554 175.546
R2160 GNDA.n1583 GNDA.n1556 175.546
R2161 GNDA.n1062 GNDA.n474 175.546
R2162 GNDA.n1066 GNDA.n1064 175.546
R2163 GNDA.n1074 GNDA.n470 175.546
R2164 GNDA.n1081 GNDA.n1076 175.546
R2165 GNDA.n1079 GNDA.n1078 175.546
R2166 GNDA.n544 GNDA.n543 175.546
R2167 GNDA.n541 GNDA.n521 175.546
R2168 GNDA.n537 GNDA.n536 175.546
R2169 GNDA.n534 GNDA.n524 175.546
R2170 GNDA.n530 GNDA.n529 175.546
R2171 GNDA.n569 GNDA.n509 175.546
R2172 GNDA.n565 GNDA.n509 175.546
R2173 GNDA.n565 GNDA.n511 175.546
R2174 GNDA.n561 GNDA.n511 175.546
R2175 GNDA.n561 GNDA.n559 175.546
R2176 GNDA.n559 GNDA.n558 175.546
R2177 GNDA.n558 GNDA.n513 175.546
R2178 GNDA.n554 GNDA.n513 175.546
R2179 GNDA.n554 GNDA.n515 175.546
R2180 GNDA.n550 GNDA.n515 175.546
R2181 GNDA.n550 GNDA.n518 175.546
R2182 GNDA.n650 GNDA.n626 175.546
R2183 GNDA.n648 GNDA.n627 175.546
R2184 GNDA.n641 GNDA.n640 175.546
R2185 GNDA.n638 GNDA.n632 175.546
R2186 GNDA.n659 GNDA.n658 175.546
R2187 GNDA.n1233 GNDA.n1215 175.546
R2188 GNDA.n1236 GNDA.n1216 175.546
R2189 GNDA.n1220 GNDA.n1219 175.546
R2190 GNDA.n1239 GNDA.n1221 175.546
R2191 GNDA.n1225 GNDA.n1224 175.546
R2192 GNDA.n1410 GNDA.n1250 175.546
R2193 GNDA.n1410 GNDA.n1248 175.546
R2194 GNDA.n1414 GNDA.n1248 175.546
R2195 GNDA.n1414 GNDA.n1246 175.546
R2196 GNDA.n1418 GNDA.n1246 175.546
R2197 GNDA.n1418 GNDA.n1232 175.546
R2198 GNDA.n1422 GNDA.n1232 175.546
R2199 GNDA.n1422 GNDA.n1230 175.546
R2200 GNDA.n1426 GNDA.n1230 175.546
R2201 GNDA.n1426 GNDA.n1228 175.546
R2202 GNDA.n1430 GNDA.n1228 175.546
R2203 GNDA.n1386 GNDA.n1260 175.546
R2204 GNDA.n1386 GNDA.n1258 175.546
R2205 GNDA.n1391 GNDA.n1258 175.546
R2206 GNDA.n1391 GNDA.n1256 175.546
R2207 GNDA.n1395 GNDA.n1256 175.546
R2208 GNDA.n1396 GNDA.n1395 175.546
R2209 GNDA.n1398 GNDA.n1396 175.546
R2210 GNDA.n1398 GNDA.n1254 175.546
R2211 GNDA.n1402 GNDA.n1254 175.546
R2212 GNDA.n1402 GNDA.n1252 175.546
R2213 GNDA.n1406 GNDA.n1252 175.546
R2214 GNDA.n1378 GNDA.n1262 175.546
R2215 GNDA.n1299 GNDA.n1291 175.546
R2216 GNDA.n1303 GNDA.n1301 175.546
R2217 GNDA.n1315 GNDA.n1288 175.546
R2218 GNDA.n1320 GNDA.n1317 175.546
R2219 GNDA.n1485 GNDA.n1483 175.546
R2220 GNDA.n1493 GNDA.n268 175.546
R2221 GNDA.n1497 GNDA.n1495 175.546
R2222 GNDA.n1508 GNDA.n264 175.546
R2223 GNDA.n1511 GNDA.n1510 175.546
R2224 GNDA.n352 GNDA.n318 175.546
R2225 GNDA.n350 GNDA.n319 175.546
R2226 GNDA.n342 GNDA.n341 175.546
R2227 GNDA.n339 GNDA.n326 175.546
R2228 GNDA.n410 GNDA.n293 175.546
R2229 GNDA.n417 GNDA.n291 175.546
R2230 GNDA.n421 GNDA.n419 175.546
R2231 GNDA.n425 GNDA.n289 175.546
R2232 GNDA.n429 GNDA.n427 175.546
R2233 GNDA.n433 GNDA.n287 175.546
R2234 GNDA.n436 GNDA.n435 175.546
R2235 GNDA.n457 GNDA.n262 175.546
R2236 GNDA.n457 GNDA.n278 175.546
R2237 GNDA.n453 GNDA.n278 175.546
R2238 GNDA.n453 GNDA.n450 175.546
R2239 GNDA.n450 GNDA.n449 175.546
R2240 GNDA.n449 GNDA.n280 175.546
R2241 GNDA.n445 GNDA.n280 175.546
R2242 GNDA.n445 GNDA.n282 175.546
R2243 GNDA.n441 GNDA.n282 175.546
R2244 GNDA.n441 GNDA.n284 175.546
R2245 GNDA.n437 GNDA.n284 175.546
R2246 GNDA.n1666 GNDA.n1664 163.333
R2247 GNDA.n1205 GNDA.n1095 163.333
R2248 GNDA.n753 GNDA.n679 163.333
R2249 GNDA.n1929 GNDA.n141 163.333
R2250 GNDA.n921 GNDA.n919 163.333
R2251 GNDA.n653 GNDA.n503 163.333
R2252 GNDA.n1375 GNDA.n1265 163.333
R2253 GNDA.n357 GNDA.n355 163.333
R2254 GNDA.n1810 GNDA.n1802 163.333
R2255 GNDA.n1528 GNDA.n245 157.601
R2256 GNDA.t2 GNDA.t5 155.788
R2257 GNDA.n1664 GNDA.n218 150
R2258 GNDA.n1654 GNDA.n1613 150
R2259 GNDA.n1652 GNDA.n1614 150
R2260 GNDA.n1642 GNDA.n1640 150
R2261 GNDA.n1670 GNDA.n216 150
R2262 GNDA.n1674 GNDA.n1672 150
R2263 GNDA.n1678 GNDA.n214 150
R2264 GNDA.n1682 GNDA.n1680 150
R2265 GNDA.n1686 GNDA.n212 150
R2266 GNDA.n1690 GNDA.n1688 150
R2267 GNDA.n1694 GNDA.n210 150
R2268 GNDA.n1697 GNDA.n1696 150
R2269 GNDA.n1699 GNDA.n1697 150
R2270 GNDA.n1713 GNDA.n1712 150
R2271 GNDA.n1710 GNDA.n204 150
R2272 GNDA.n1706 GNDA.n1705 150
R2273 GNDA.n1703 GNDA.n207 150
R2274 GNDA.n1205 GNDA.n1096 150
R2275 GNDA.n1127 GNDA.n1126 150
R2276 GNDA.n1138 GNDA.n1137 150
R2277 GNDA.n1143 GNDA.n1142 150
R2278 GNDA.n1203 GNDA.n1114 150
R2279 GNDA.n1199 GNDA.n1198 150
R2280 GNDA.n1195 GNDA.n1194 150
R2281 GNDA.n1191 GNDA.n1190 150
R2282 GNDA.n1187 GNDA.n1186 150
R2283 GNDA.n1183 GNDA.n1182 150
R2284 GNDA.n1179 GNDA.n1178 150
R2285 GNDA.n1175 GNDA.n1104 150
R2286 GNDA.n1172 GNDA.n1104 150
R2287 GNDA.n1158 GNDA.n1157 150
R2288 GNDA.n1162 GNDA.n1161 150
R2289 GNDA.n1166 GNDA.n1165 150
R2290 GNDA.n1170 GNDA.n1169 150
R2291 GNDA.n755 GNDA.n753 150
R2292 GNDA.n767 GNDA.n675 150
R2293 GNDA.n771 GNDA.n769 150
R2294 GNDA.n779 GNDA.n671 150
R2295 GNDA.n742 GNDA.n740 150
R2296 GNDA.n738 GNDA.n681 150
R2297 GNDA.n734 GNDA.n732 150
R2298 GNDA.n730 GNDA.n683 150
R2299 GNDA.n726 GNDA.n724 150
R2300 GNDA.n722 GNDA.n685 150
R2301 GNDA.n718 GNDA.n716 150
R2302 GNDA.n714 GNDA.n687 150
R2303 GNDA.n710 GNDA.n687 150
R2304 GNDA.n697 GNDA.n695 150
R2305 GNDA.n701 GNDA.n691 150
R2306 GNDA.n704 GNDA.n703 150
R2307 GNDA.n708 GNDA.n707 150
R2308 GNDA.n1929 GNDA.n142 150
R2309 GNDA.n176 GNDA.n175 150
R2310 GNDA.n1862 GNDA.n1861 150
R2311 GNDA.n1867 GNDA.n1866 150
R2312 GNDA.n1927 GNDA.n160 150
R2313 GNDA.n1923 GNDA.n1922 150
R2314 GNDA.n1919 GNDA.n1918 150
R2315 GNDA.n1915 GNDA.n1914 150
R2316 GNDA.n1911 GNDA.n1910 150
R2317 GNDA.n1907 GNDA.n1906 150
R2318 GNDA.n1903 GNDA.n1902 150
R2319 GNDA.n1899 GNDA.n150 150
R2320 GNDA.n1896 GNDA.n150 150
R2321 GNDA.n1882 GNDA.n1881 150
R2322 GNDA.n1886 GNDA.n1885 150
R2323 GNDA.n1890 GNDA.n1889 150
R2324 GNDA.n1894 GNDA.n1893 150
R2325 GNDA.n919 GNDA.n877 150
R2326 GNDA.n911 GNDA.n909 150
R2327 GNDA.n898 GNDA.n896 150
R2328 GNDA.n900 GNDA.n895 150
R2329 GNDA.n925 GNDA.n875 150
R2330 GNDA.n929 GNDA.n927 150
R2331 GNDA.n933 GNDA.n873 150
R2332 GNDA.n937 GNDA.n935 150
R2333 GNDA.n941 GNDA.n871 150
R2334 GNDA.n945 GNDA.n943 150
R2335 GNDA.n949 GNDA.n869 150
R2336 GNDA.n952 GNDA.n951 150
R2337 GNDA.n954 GNDA.n952 150
R2338 GNDA.n968 GNDA.n967 150
R2339 GNDA.n965 GNDA.n863 150
R2340 GNDA.n961 GNDA.n960 150
R2341 GNDA.n958 GNDA.n866 150
R2342 GNDA.n653 GNDA.n504 150
R2343 GNDA.n645 GNDA.n644 150
R2344 GNDA.n634 GNDA.n633 150
R2345 GNDA.n655 GNDA.n483 150
R2346 GNDA.n619 GNDA.n618 150
R2347 GNDA.n615 GNDA.n614 150
R2348 GNDA.n611 GNDA.n610 150
R2349 GNDA.n607 GNDA.n606 150
R2350 GNDA.n603 GNDA.n602 150
R2351 GNDA.n599 GNDA.n598 150
R2352 GNDA.n595 GNDA.n594 150
R2353 GNDA.n591 GNDA.n491 150
R2354 GNDA.n588 GNDA.n491 150
R2355 GNDA.n574 GNDA.n573 150
R2356 GNDA.n578 GNDA.n577 150
R2357 GNDA.n582 GNDA.n581 150
R2358 GNDA.n586 GNDA.n585 150
R2359 GNDA.n1375 GNDA.n1266 150
R2360 GNDA.n1296 GNDA.n1295 150
R2361 GNDA.n1307 GNDA.n1306 150
R2362 GNDA.n1312 GNDA.n1311 150
R2363 GNDA.n1373 GNDA.n1284 150
R2364 GNDA.n1369 GNDA.n1368 150
R2365 GNDA.n1365 GNDA.n1364 150
R2366 GNDA.n1361 GNDA.n1360 150
R2367 GNDA.n1357 GNDA.n1356 150
R2368 GNDA.n1353 GNDA.n1352 150
R2369 GNDA.n1349 GNDA.n1348 150
R2370 GNDA.n1345 GNDA.n1274 150
R2371 GNDA.n1342 GNDA.n1274 150
R2372 GNDA.n1328 GNDA.n1327 150
R2373 GNDA.n1332 GNDA.n1331 150
R2374 GNDA.n1336 GNDA.n1335 150
R2375 GNDA.n1340 GNDA.n1339 150
R2376 GNDA.n355 GNDA.n312 150
R2377 GNDA.n347 GNDA.n345 150
R2378 GNDA.n334 GNDA.n332 150
R2379 GNDA.n336 GNDA.n331 150
R2380 GNDA.n361 GNDA.n310 150
R2381 GNDA.n365 GNDA.n363 150
R2382 GNDA.n369 GNDA.n308 150
R2383 GNDA.n373 GNDA.n371 150
R2384 GNDA.n377 GNDA.n306 150
R2385 GNDA.n381 GNDA.n379 150
R2386 GNDA.n385 GNDA.n304 150
R2387 GNDA.n388 GNDA.n387 150
R2388 GNDA.n390 GNDA.n388 150
R2389 GNDA.n404 GNDA.n403 150
R2390 GNDA.n401 GNDA.n298 150
R2391 GNDA.n397 GNDA.n396 150
R2392 GNDA.n394 GNDA.n301 150
R2393 GNDA.n1810 GNDA.n1809 150
R2394 GNDA.n2059 GNDA.n15 150
R2395 GNDA.n2062 GNDA.n2061 150
R2396 GNDA.n2065 GNDA.n2064 150
R2397 GNDA.n1799 GNDA.n1798 150
R2398 GNDA.n1796 GNDA.n1737 150
R2399 GNDA.n1792 GNDA.n1790 150
R2400 GNDA.n1788 GNDA.n1739 150
R2401 GNDA.n1784 GNDA.n1782 150
R2402 GNDA.n1780 GNDA.n1741 150
R2403 GNDA.n1776 GNDA.n1774 150
R2404 GNDA.n1772 GNDA.n1743 150
R2405 GNDA.n1768 GNDA.n1743 150
R2406 GNDA.n1755 GNDA.n1753 150
R2407 GNDA.n1759 GNDA.n1747 150
R2408 GNDA.n1762 GNDA.n1761 150
R2409 GNDA.n1766 GNDA.n1765 150
R2410 GNDA.n1606 GNDA.n1544 137.035
R2411 GNDA.n1728 GNDA.n1727 137.035
R2412 GNDA.n1937 GNDA.n1935 137.035
R2413 GNDA.n1852 GNDA.n187 134.268
R2414 GNDA.n187 GNDA.n185 134.268
R2415 GNDA.n2050 GNDA.n2049 133.517
R2416 GNDA.n979 GNDA.n978 133.517
R2417 GNDA.n1723 GNDA.n1722 130.25
R2418 GNDA.n1939 GNDA.n136 130.25
R2419 GNDA.n2052 GNDA.n20 130.25
R2420 GNDA.n1479 GNDA.n1477 126.782
R2421 GNDA.n1942 GNDA.n1940 126.782
R2422 GNDA.n789 GNDA.n665 126.782
R2423 GNDA.n1724 GNDA.n80 126.782
R2424 GNDA.n1054 GNDA.n1052 126.782
R2425 GNDA.n1212 GNDA.n276 126.782
R2426 GNDA.n1471 GNDA.n461 124.832
R2427 GNDA.n2024 GNDA.n78 124.832
R2428 GNDA.n1056 GNDA.n476 124.832
R2429 GNDA.n1944 GNDA.n132 124.832
R2430 GNDA.n1045 GNDA.n666 124.832
R2431 GNDA.n1602 GNDA.n1545 124.832
R2432 GNDA.n569 GNDA.n507 124.832
R2433 GNDA.n1381 GNDA.n1260 124.832
R2434 GNDA.n1481 GNDA.n272 124.832
R2435 GNDA.n1607 GNDA.n1606 122.109
R2436 GNDA.n1660 GNDA.n1607 122.109
R2437 GNDA.n1660 GNDA.n1659 122.109
R2438 GNDA.n1648 GNDA.n1647 122.109
R2439 GNDA.n1647 GNDA.n1646 122.109
R2440 GNDA.n1646 GNDA.n1634 122.109
R2441 GNDA.n1722 GNDA.n1721 122.109
R2442 GNDA.n1814 GNDA.n1729 122.109
R2443 GNDA.n1805 GNDA.n1729 122.109
R2444 GNDA.n1805 GNDA.n18 122.109
R2445 GNDA.n2055 GNDA.n18 122.109
R2446 GNDA.n2073 GNDA.n6 122.109
R2447 GNDA.n2073 GNDA.n2072 122.109
R2448 GNDA.n2072 GNDA.n2071 122.109
R2449 GNDA.n2071 GNDA.n7 122.109
R2450 GNDA.n1935 GNDA.n137 122.109
R2451 GNDA.n169 GNDA.n168 122.109
R2452 GNDA.n180 GNDA.n168 122.109
R2453 GNDA.n181 GNDA.n180 122.109
R2454 GNDA.n1872 GNDA.n1871 122.109
R2455 GNDA.n1873 GNDA.n1872 122.109
R2456 GNDA.n1873 GNDA.n20 122.109
R2457 GNDA.t16 GNDA.n67 121.835
R2458 GNDA.t16 GNDA.n60 121.835
R2459 GNDA.t16 GNDA.n1244 121.835
R2460 GNDA.t8 GNDA.n1658 118.04
R2461 GNDA.n1721 GNDA.t25 118.04
R2462 GNDA.n1939 GNDA.n1938 118.04
R2463 GNDA.n1727 GNDA.n71 116.683
R2464 GNDA.t37 GNDA.n137 112.612
R2465 GNDA.n1856 GNDA.t4 112.612
R2466 GNDA.n241 GNDA.t1 111.338
R2467 GNDA.n1533 GNDA.t9 110.826
R2468 GNDA.n241 GNDA.t7 110.659
R2469 GNDA.n1532 GNDA.t12 110.591
R2470 GNDA.n1 GNDA.n51 14.555
R2471 GNDA.n0 GNDA.n54 14.555
R2472 GNDA.n1848 GNDA.n182 101.718
R2473 GNDA.n1623 GNDA.n1617 101.718
R2474 GNDA.n1632 GNDA.n1619 101.718
R2475 GNDA.n1854 GNDA.n184 101.718
R2476 GNDA.n1852 GNDA.n1847 91.069
R2477 GNDA.n1850 GNDA.n185 91.069
R2478 GNDA.n1630 GNDA.n1622 91.069
R2479 GNDA.n1630 GNDA.n1629 91.069
R2480 GNDA.n1627 GNDA.n1620 91.069
R2481 GNDA.n1627 GNDA.n1626 91.069
R2482 GNDA.n1411 GNDA.n1249 90.3496
R2483 GNDA.n1412 GNDA.n1411 90.3496
R2484 GNDA.n1413 GNDA.n1412 90.3496
R2485 GNDA.n1413 GNDA.n1245 90.3496
R2486 GNDA.n1419 GNDA.n1245 90.3496
R2487 GNDA.n1421 GNDA.n1420 90.3496
R2488 GNDA.n1421 GNDA.n1229 90.3496
R2489 GNDA.n1427 GNDA.n1229 90.3496
R2490 GNDA.n1428 GNDA.n1427 90.3496
R2491 GNDA.n1429 GNDA.n1428 90.3496
R2492 GNDA.n1447 GNDA.n1446 90.3496
R2493 GNDA.n1446 GNDA.n1445 90.3496
R2494 GNDA.n1445 GNDA.n1435 90.3496
R2495 GNDA.n1439 GNDA.n1435 90.3496
R2496 GNDA.n1439 GNDA.n248 90.3496
R2497 GNDA.n1527 GNDA.n250 90.3496
R2498 GNDA.n1521 GNDA.n250 90.3496
R2499 GNDA.n1521 GNDA.n1520 90.3496
R2500 GNDA.n1520 GNDA.n1519 90.3496
R2501 GNDA.n1519 GNDA.n257 90.3496
R2502 GNDA.n459 GNDA.n458 90.3496
R2503 GNDA.n458 GNDA.n277 90.3496
R2504 GNDA.n452 GNDA.n277 90.3496
R2505 GNDA.n452 GNDA.n451 90.3496
R2506 GNDA.n451 GNDA.n57 90.3496
R2507 GNDA.n444 GNDA.n58 90.3496
R2508 GNDA.n444 GNDA.n443 90.3496
R2509 GNDA.n443 GNDA.n442 90.3496
R2510 GNDA.n442 GNDA.n283 90.3496
R2511 GNDA.n283 GNDA.n55 90.3496
R2512 GNDA.n1826 GNDA.n1825 84.306
R2513 GNDA.n1816 GNDA.n197 84.306
R2514 GNDA.n1616 GNDA.t35 77.3363
R2515 GNDA.n1827 GNDA.n136 77.3363
R2516 GNDA.n1478 GNDA.n270 76.3222
R2517 GNDA.n1489 GNDA.n1488 76.3222
R2518 GNDA.n1490 GNDA.n266 76.3222
R2519 GNDA.n1501 GNDA.n1500 76.3222
R2520 GNDA.n1505 GNDA.n1504 76.3222
R2521 GNDA.n1502 GNDA.n261 76.3222
R2522 GNDA.n1471 GNDA.n1470 76.3222
R2523 GNDA.n1468 GNDA.n1214 76.3222
R2524 GNDA.n1464 GNDA.n1463 76.3222
R2525 GNDA.n1457 GNDA.n1218 76.3222
R2526 GNDA.n1456 GNDA.n1455 76.3222
R2527 GNDA.n1449 GNDA.n1223 76.3222
R2528 GNDA.n1209 GNDA.n1208 76.3222
R2529 GNDA.n1122 GNDA.n1121 76.3222
R2530 GNDA.n1132 GNDA.n1131 76.3222
R2531 GNDA.n1133 GNDA.n1119 76.3222
R2532 GNDA.n1148 GNDA.n1147 76.3222
R2533 GNDA.n1149 GNDA.n274 76.3222
R2534 GNDA.n2025 GNDA.n2024 76.3222
R2535 GNDA.n2020 GNDA.n76 76.3222
R2536 GNDA.n2017 GNDA.n75 76.3222
R2537 GNDA.n2013 GNDA.n74 76.3222
R2538 GNDA.n2009 GNDA.n73 76.3222
R2539 GNDA.n2005 GNDA.n72 76.3222
R2540 GNDA.n1941 GNDA.n130 76.3222
R2541 GNDA.n1952 GNDA.n1951 76.3222
R2542 GNDA.n1953 GNDA.n126 76.3222
R2543 GNDA.n1964 GNDA.n1963 76.3222
R2544 GNDA.n1967 GNDA.n1966 76.3222
R2545 GNDA.n1977 GNDA.n100 76.3222
R2546 GNDA.n1998 GNDA.n39 76.3222
R2547 GNDA.n1994 GNDA.n40 76.3222
R2548 GNDA.n1990 GNDA.n41 76.3222
R2549 GNDA.n1986 GNDA.n42 76.3222
R2550 GNDA.n1982 GNDA.n43 76.3222
R2551 GNDA.n1978 GNDA.n44 76.3222
R2552 GNDA.n793 GNDA.n792 76.3222
R2553 GNDA.n796 GNDA.n795 76.3222
R2554 GNDA.n801 GNDA.n800 76.3222
R2555 GNDA.n804 GNDA.n803 76.3222
R2556 GNDA.n809 GNDA.n808 76.3222
R2557 GNDA.n812 GNDA.n811 76.3222
R2558 GNDA.n819 GNDA.n818 76.3222
R2559 GNDA.n824 GNDA.n823 76.3222
R2560 GNDA.n825 GNDA.n816 76.3222
R2561 GNDA.n832 GNDA.n831 76.3222
R2562 GNDA.n836 GNDA.n814 76.3222
R2563 GNDA.n839 GNDA.n838 76.3222
R2564 GNDA.n1057 GNDA.n1056 76.3222
R2565 GNDA.n1060 GNDA.n1059 76.3222
R2566 GNDA.n1069 GNDA.n1068 76.3222
R2567 GNDA.n1072 GNDA.n1071 76.3222
R2568 GNDA.n1084 GNDA.n1083 76.3222
R2569 GNDA.n1087 GNDA.n1086 76.3222
R2570 GNDA.n750 GNDA.n748 76.3222
R2571 GNDA.n759 GNDA.n677 76.3222
R2572 GNDA.n764 GNDA.n761 76.3222
R2573 GNDA.n774 GNDA.n673 76.3222
R2574 GNDA.n775 GNDA.n668 76.3222
R2575 GNDA.n786 GNDA.n785 76.3222
R2576 GNDA.n1945 GNDA.n1944 76.3222
R2577 GNDA.n1948 GNDA.n1947 76.3222
R2578 GNDA.n1957 GNDA.n1956 76.3222
R2579 GNDA.n1960 GNDA.n1959 76.3222
R2580 GNDA.n1971 GNDA.n1970 76.3222
R2581 GNDA.n1974 GNDA.n1973 76.3222
R2582 GNDA.n119 GNDA.n34 76.3222
R2583 GNDA.n115 GNDA.n35 76.3222
R2584 GNDA.n111 GNDA.n36 76.3222
R2585 GNDA.n107 GNDA.n37 76.3222
R2586 GNDA.n103 GNDA.n38 76.3222
R2587 GNDA.n2029 GNDA.n2028 76.3222
R2588 GNDA.n2049 GNDA.n2048 76.3222
R2589 GNDA.n2044 GNDA.n26 76.3222
R2590 GNDA.n2042 GNDA.n2041 76.3222
R2591 GNDA.n2037 GNDA.n29 76.3222
R2592 GNDA.n2035 GNDA.n2034 76.3222
R2593 GNDA.n2030 GNDA.n32 76.3222
R2594 GNDA.n978 GNDA.n856 76.3222
R2595 GNDA.n985 GNDA.n984 76.3222
R2596 GNDA.n986 GNDA.n854 76.3222
R2597 GNDA.n993 GNDA.n992 76.3222
R2598 GNDA.n994 GNDA.n852 76.3222
R2599 GNDA.n1001 GNDA.n1000 76.3222
R2600 GNDA.n1021 GNDA.n1020 76.3222
R2601 GNDA.n1016 GNDA.n845 76.3222
R2602 GNDA.n1014 GNDA.n1013 76.3222
R2603 GNDA.n1009 GNDA.n848 76.3222
R2604 GNDA.n1007 GNDA.n1006 76.3222
R2605 GNDA.n1002 GNDA.n851 76.3222
R2606 GNDA.n1045 GNDA.n1044 76.3222
R2607 GNDA.n1042 GNDA.n791 76.3222
R2608 GNDA.n1038 GNDA.n1037 76.3222
R2609 GNDA.n1031 GNDA.n798 76.3222
R2610 GNDA.n1030 GNDA.n1029 76.3222
R2611 GNDA.n1023 GNDA.n806 76.3222
R2612 GNDA.n882 GNDA.n881 76.3222
R2613 GNDA.n915 GNDA.n914 76.3222
R2614 GNDA.n906 GNDA.n887 76.3222
R2615 GNDA.n904 GNDA.n903 76.3222
R2616 GNDA.n889 GNDA.n858 76.3222
R2617 GNDA.n976 GNDA.n975 76.3222
R2618 GNDA.n1000 GNDA.n999 76.3222
R2619 GNDA.n995 GNDA.n994 76.3222
R2620 GNDA.n992 GNDA.n991 76.3222
R2621 GNDA.n987 GNDA.n986 76.3222
R2622 GNDA.n984 GNDA.n983 76.3222
R2623 GNDA.n32 GNDA.n30 76.3222
R2624 GNDA.n2036 GNDA.n2035 76.3222
R2625 GNDA.n29 GNDA.n27 76.3222
R2626 GNDA.n2043 GNDA.n2042 76.3222
R2627 GNDA.n26 GNDA.n24 76.3222
R2628 GNDA.n82 GNDA.n81 76.3222
R2629 GNDA.n85 GNDA.n84 76.3222
R2630 GNDA.n88 GNDA.n87 76.3222
R2631 GNDA.n91 GNDA.n90 76.3222
R2632 GNDA.n94 GNDA.n93 76.3222
R2633 GNDA.n97 GNDA.n96 76.3222
R2634 GNDA.n1577 GNDA.n45 76.3222
R2635 GNDA.n1573 GNDA.n46 76.3222
R2636 GNDA.n1569 GNDA.n47 76.3222
R2637 GNDA.n1565 GNDA.n48 76.3222
R2638 GNDA.n1561 GNDA.n49 76.3222
R2639 GNDA.n1557 GNDA.n50 76.3222
R2640 GNDA.n1053 GNDA.n474 76.3222
R2641 GNDA.n1064 GNDA.n1063 76.3222
R2642 GNDA.n1065 GNDA.n470 76.3222
R2643 GNDA.n1076 GNDA.n1075 76.3222
R2644 GNDA.n1080 GNDA.n1079 76.3222
R2645 GNDA.n1077 GNDA.n465 76.3222
R2646 GNDA.n545 GNDA.n544 76.3222
R2647 GNDA.n542 GNDA.n541 76.3222
R2648 GNDA.n537 GNDA.n523 76.3222
R2649 GNDA.n535 GNDA.n534 76.3222
R2650 GNDA.n530 GNDA.n526 76.3222
R2651 GNDA.n528 GNDA.n527 76.3222
R2652 GNDA.n626 GNDA.n625 76.3222
R2653 GNDA.n649 GNDA.n648 76.3222
R2654 GNDA.n641 GNDA.n630 76.3222
R2655 GNDA.n639 GNDA.n638 76.3222
R2656 GNDA.n658 GNDA.n481 76.3222
R2657 GNDA.n663 GNDA.n478 76.3222
R2658 GNDA.n1234 GNDA.n1233 76.3222
R2659 GNDA.n1235 GNDA.n1216 76.3222
R2660 GNDA.n1237 GNDA.n1219 76.3222
R2661 GNDA.n1238 GNDA.n1221 76.3222
R2662 GNDA.n1240 GNDA.n1224 76.3222
R2663 GNDA.n1241 GNDA.n1226 76.3222
R2664 GNDA.n1379 GNDA.n1378 76.3222
R2665 GNDA.n1291 GNDA.n1290 76.3222
R2666 GNDA.n1301 GNDA.n1300 76.3222
R2667 GNDA.n1302 GNDA.n1288 76.3222
R2668 GNDA.n1317 GNDA.n1316 76.3222
R2669 GNDA.n1319 GNDA.n1318 76.3222
R2670 GNDA.n659 GNDA.n478 76.3222
R2671 GNDA.n632 GNDA.n481 76.3222
R2672 GNDA.n640 GNDA.n639 76.3222
R2673 GNDA.n630 GNDA.n627 76.3222
R2674 GNDA.n650 GNDA.n649 76.3222
R2675 GNDA.n625 GNDA.n624 76.3222
R2676 GNDA.n785 GNDA.n784 76.3222
R2677 GNDA.n776 GNDA.n775 76.3222
R2678 GNDA.n763 GNDA.n673 76.3222
R2679 GNDA.n761 GNDA.n760 76.3222
R2680 GNDA.n749 GNDA.n677 76.3222
R2681 GNDA.n748 GNDA.n747 76.3222
R2682 GNDA.n975 GNDA.n974 76.3222
R2683 GNDA.n890 GNDA.n889 76.3222
R2684 GNDA.n905 GNDA.n904 76.3222
R2685 GNDA.n887 GNDA.n883 76.3222
R2686 GNDA.n916 GNDA.n915 76.3222
R2687 GNDA.n881 GNDA.n880 76.3222
R2688 GNDA.n1560 GNDA.n50 76.3222
R2689 GNDA.n1564 GNDA.n49 76.3222
R2690 GNDA.n1568 GNDA.n48 76.3222
R2691 GNDA.n1572 GNDA.n47 76.3222
R2692 GNDA.n1576 GNDA.n46 76.3222
R2693 GNDA.n1579 GNDA.n45 76.3222
R2694 GNDA.n1981 GNDA.n44 76.3222
R2695 GNDA.n1985 GNDA.n43 76.3222
R2696 GNDA.n1989 GNDA.n42 76.3222
R2697 GNDA.n1993 GNDA.n41 76.3222
R2698 GNDA.n1997 GNDA.n40 76.3222
R2699 GNDA.n2001 GNDA.n39 76.3222
R2700 GNDA.n2028 GNDA.n33 76.3222
R2701 GNDA.n106 GNDA.n38 76.3222
R2702 GNDA.n110 GNDA.n37 76.3222
R2703 GNDA.n114 GNDA.n36 76.3222
R2704 GNDA.n118 GNDA.n35 76.3222
R2705 GNDA.n122 GNDA.n34 76.3222
R2706 GNDA.n1320 GNDA.n1319 76.3222
R2707 GNDA.n1316 GNDA.n1315 76.3222
R2708 GNDA.n1303 GNDA.n1302 76.3222
R2709 GNDA.n1300 GNDA.n1299 76.3222
R2710 GNDA.n1290 GNDA.n1262 76.3222
R2711 GNDA.n1380 GNDA.n1379 76.3222
R2712 GNDA.n529 GNDA.n528 76.3222
R2713 GNDA.n526 GNDA.n524 76.3222
R2714 GNDA.n536 GNDA.n535 76.3222
R2715 GNDA.n523 GNDA.n521 76.3222
R2716 GNDA.n543 GNDA.n542 76.3222
R2717 GNDA.n546 GNDA.n545 76.3222
R2718 GNDA.n838 GNDA.n837 76.3222
R2719 GNDA.n833 GNDA.n814 76.3222
R2720 GNDA.n831 GNDA.n830 76.3222
R2721 GNDA.n826 GNDA.n825 76.3222
R2722 GNDA.n823 GNDA.n822 76.3222
R2723 GNDA.n818 GNDA.n466 76.3222
R2724 GNDA.n851 GNDA.n849 76.3222
R2725 GNDA.n1008 GNDA.n1007 76.3222
R2726 GNDA.n848 GNDA.n846 76.3222
R2727 GNDA.n1015 GNDA.n1014 76.3222
R2728 GNDA.n845 GNDA.n843 76.3222
R2729 GNDA.n1022 GNDA.n1021 76.3222
R2730 GNDA.n1482 GNDA.n1481 76.3222
R2731 GNDA.n1485 GNDA.n1484 76.3222
R2732 GNDA.n1494 GNDA.n1493 76.3222
R2733 GNDA.n1497 GNDA.n1496 76.3222
R2734 GNDA.n1509 GNDA.n1508 76.3222
R2735 GNDA.n1512 GNDA.n1511 76.3222
R2736 GNDA.n318 GNDA.n317 76.3222
R2737 GNDA.n351 GNDA.n350 76.3222
R2738 GNDA.n342 GNDA.n323 76.3222
R2739 GNDA.n340 GNDA.n339 76.3222
R2740 GNDA.n325 GNDA.n293 76.3222
R2741 GNDA.n412 GNDA.n411 76.3222
R2742 GNDA.n418 GNDA.n417 76.3222
R2743 GNDA.n421 GNDA.n420 76.3222
R2744 GNDA.n426 GNDA.n425 76.3222
R2745 GNDA.n429 GNDA.n428 76.3222
R2746 GNDA.n434 GNDA.n433 76.3222
R2747 GNDA.n435 GNDA.n434 76.3222
R2748 GNDA.n428 GNDA.n287 76.3222
R2749 GNDA.n427 GNDA.n426 76.3222
R2750 GNDA.n420 GNDA.n289 76.3222
R2751 GNDA.n419 GNDA.n418 76.3222
R2752 GNDA.n411 GNDA.n410 76.3222
R2753 GNDA.n326 GNDA.n325 76.3222
R2754 GNDA.n341 GNDA.n340 76.3222
R2755 GNDA.n323 GNDA.n319 76.3222
R2756 GNDA.n352 GNDA.n351 76.3222
R2757 GNDA.n317 GNDA.n316 76.3222
R2758 GNDA.n1150 GNDA.n1149 76.3222
R2759 GNDA.n1147 GNDA.n1146 76.3222
R2760 GNDA.n1134 GNDA.n1133 76.3222
R2761 GNDA.n1131 GNDA.n1130 76.3222
R2762 GNDA.n1121 GNDA.n1093 76.3222
R2763 GNDA.n1210 GNDA.n1209 76.3222
R2764 GNDA.n1503 GNDA.n1502 76.3222
R2765 GNDA.n1506 GNDA.n1505 76.3222
R2766 GNDA.n1500 GNDA.n1499 76.3222
R2767 GNDA.n1491 GNDA.n1490 76.3222
R2768 GNDA.n1488 GNDA.n1487 76.3222
R2769 GNDA.n1479 GNDA.n1478 76.3222
R2770 GNDA.n1483 GNDA.n1482 76.3222
R2771 GNDA.n1484 GNDA.n268 76.3222
R2772 GNDA.n1495 GNDA.n1494 76.3222
R2773 GNDA.n1496 GNDA.n264 76.3222
R2774 GNDA.n1510 GNDA.n1509 76.3222
R2775 GNDA.n1513 GNDA.n1512 76.3222
R2776 GNDA.n811 GNDA.n810 76.3222
R2777 GNDA.n808 GNDA.n807 76.3222
R2778 GNDA.n803 GNDA.n802 76.3222
R2779 GNDA.n800 GNDA.n799 76.3222
R2780 GNDA.n795 GNDA.n794 76.3222
R2781 GNDA.n792 GNDA.n789 76.3222
R2782 GNDA.n1044 GNDA.n1043 76.3222
R2783 GNDA.n1039 GNDA.n791 76.3222
R2784 GNDA.n1037 GNDA.n1036 76.3222
R2785 GNDA.n1032 GNDA.n1031 76.3222
R2786 GNDA.n1029 GNDA.n1028 76.3222
R2787 GNDA.n1024 GNDA.n1023 76.3222
R2788 GNDA.n1965 GNDA.n100 76.3222
R2789 GNDA.n1968 GNDA.n1967 76.3222
R2790 GNDA.n1963 GNDA.n1962 76.3222
R2791 GNDA.n1954 GNDA.n1953 76.3222
R2792 GNDA.n1951 GNDA.n1950 76.3222
R2793 GNDA.n1942 GNDA.n1941 76.3222
R2794 GNDA.n1946 GNDA.n1945 76.3222
R2795 GNDA.n1947 GNDA.n128 76.3222
R2796 GNDA.n1958 GNDA.n1957 76.3222
R2797 GNDA.n1959 GNDA.n124 76.3222
R2798 GNDA.n1972 GNDA.n1971 76.3222
R2799 GNDA.n1975 GNDA.n1974 76.3222
R2800 GNDA.n96 GNDA.n95 76.3222
R2801 GNDA.n93 GNDA.n92 76.3222
R2802 GNDA.n90 GNDA.n89 76.3222
R2803 GNDA.n87 GNDA.n86 76.3222
R2804 GNDA.n84 GNDA.n83 76.3222
R2805 GNDA.n81 GNDA.n80 76.3222
R2806 GNDA.n2025 GNDA.n77 76.3222
R2807 GNDA.n2018 GNDA.n76 76.3222
R2808 GNDA.n2014 GNDA.n75 76.3222
R2809 GNDA.n2010 GNDA.n74 76.3222
R2810 GNDA.n2006 GNDA.n73 76.3222
R2811 GNDA.n2002 GNDA.n72 76.3222
R2812 GNDA.n1078 GNDA.n1077 76.3222
R2813 GNDA.n1081 GNDA.n1080 76.3222
R2814 GNDA.n1075 GNDA.n1074 76.3222
R2815 GNDA.n1066 GNDA.n1065 76.3222
R2816 GNDA.n1063 GNDA.n1062 76.3222
R2817 GNDA.n1054 GNDA.n1053 76.3222
R2818 GNDA.n1058 GNDA.n1057 76.3222
R2819 GNDA.n1059 GNDA.n472 76.3222
R2820 GNDA.n1070 GNDA.n1069 76.3222
R2821 GNDA.n1071 GNDA.n468 76.3222
R2822 GNDA.n1085 GNDA.n1084 76.3222
R2823 GNDA.n1088 GNDA.n1087 76.3222
R2824 GNDA.n1241 GNDA.n1225 76.3222
R2825 GNDA.n1240 GNDA.n1239 76.3222
R2826 GNDA.n1238 GNDA.n1220 76.3222
R2827 GNDA.n1237 GNDA.n1236 76.3222
R2828 GNDA.n1235 GNDA.n1215 76.3222
R2829 GNDA.n1234 GNDA.n1212 76.3222
R2830 GNDA.n1470 GNDA.n1469 76.3222
R2831 GNDA.n1465 GNDA.n1214 76.3222
R2832 GNDA.n1463 GNDA.n1462 76.3222
R2833 GNDA.n1458 GNDA.n1457 76.3222
R2834 GNDA.n1455 GNDA.n1454 76.3222
R2835 GNDA.n1450 GNDA.n1449 76.3222
R2836 GNDA.n1699 GNDA.n1698 76.062
R2837 GNDA.n1698 GNDA.n207 76.062
R2838 GNDA.n1172 GNDA.n1105 76.062
R2839 GNDA.n1170 GNDA.n1105 76.062
R2840 GNDA.n710 GNDA.n709 76.062
R2841 GNDA.n709 GNDA.n708 76.062
R2842 GNDA.n1896 GNDA.n151 76.062
R2843 GNDA.n1894 GNDA.n151 76.062
R2844 GNDA.n954 GNDA.n953 76.062
R2845 GNDA.n953 GNDA.n866 76.062
R2846 GNDA.n588 GNDA.n492 76.062
R2847 GNDA.n586 GNDA.n492 76.062
R2848 GNDA.n1342 GNDA.n1275 76.062
R2849 GNDA.n1340 GNDA.n1275 76.062
R2850 GNDA.n390 GNDA.n389 76.062
R2851 GNDA.n389 GNDA.n301 76.062
R2852 GNDA.n1768 GNDA.n1767 76.062
R2853 GNDA.n1767 GNDA.n1766 76.062
R2854 GNDA.n1601 GNDA.n19 75.897
R2855 GNDA.n1682 GNDA.n1681 74.5978
R2856 GNDA.n1681 GNDA.n212 74.5978
R2857 GNDA.n1190 GNDA.n1110 74.5978
R2858 GNDA.n1187 GNDA.n1110 74.5978
R2859 GNDA.n725 GNDA.n683 74.5978
R2860 GNDA.n726 GNDA.n725 74.5978
R2861 GNDA.n1914 GNDA.n156 74.5978
R2862 GNDA.n1911 GNDA.n156 74.5978
R2863 GNDA.n937 GNDA.n936 74.5978
R2864 GNDA.n936 GNDA.n871 74.5978
R2865 GNDA.n606 GNDA.n498 74.5978
R2866 GNDA.n603 GNDA.n498 74.5978
R2867 GNDA.n1360 GNDA.n1280 74.5978
R2868 GNDA.n1357 GNDA.n1280 74.5978
R2869 GNDA.n373 GNDA.n372 74.5978
R2870 GNDA.n372 GNDA.n306 74.5978
R2871 GNDA.n1783 GNDA.n1739 74.5978
R2872 GNDA.n1784 GNDA.n1783 74.5978
R2873 GNDA.n2053 GNDA.t13 73.5411
R2874 GNDA.n1817 GNDA.n1728 71.9092
R2875 GNDA.n1857 GNDA.t36 71.9092
R2876 GNDA.n249 GNDA.n245 69.4466
R2877 GNDA.n1704 GNDA.t20 65.8183
R2878 GNDA.n206 GNDA.t20 65.8183
R2879 GNDA.n1711 GNDA.t20 65.8183
R2880 GNDA.n1714 GNDA.t20 65.8183
R2881 GNDA.n1695 GNDA.t20 65.8183
R2882 GNDA.n1689 GNDA.t20 65.8183
R2883 GNDA.n1687 GNDA.t20 65.8183
R2884 GNDA.n1665 GNDA.t20 65.8183
R2885 GNDA.n1671 GNDA.t20 65.8183
R2886 GNDA.n1673 GNDA.t20 65.8183
R2887 GNDA.n1679 GNDA.t20 65.8183
R2888 GNDA.t23 GNDA.n1109 65.8183
R2889 GNDA.t23 GNDA.n1108 65.8183
R2890 GNDA.t23 GNDA.n1107 65.8183
R2891 GNDA.t23 GNDA.n1106 65.8183
R2892 GNDA.t23 GNDA.n1102 65.8183
R2893 GNDA.t23 GNDA.n1100 65.8183
R2894 GNDA.t23 GNDA.n1098 65.8183
R2895 GNDA.t23 GNDA.n1204 65.8183
R2896 GNDA.t23 GNDA.n1113 65.8183
R2897 GNDA.t23 GNDA.n1112 65.8183
R2898 GNDA.t23 GNDA.n1111 65.8183
R2899 GNDA.n689 GNDA.t17 65.8183
R2900 GNDA.n702 GNDA.t17 65.8183
R2901 GNDA.n696 GNDA.t17 65.8183
R2902 GNDA.n694 GNDA.t17 65.8183
R2903 GNDA.n715 GNDA.t17 65.8183
R2904 GNDA.n717 GNDA.t17 65.8183
R2905 GNDA.n723 GNDA.t17 65.8183
R2906 GNDA.n741 GNDA.t17 65.8183
R2907 GNDA.n739 GNDA.t17 65.8183
R2908 GNDA.n733 GNDA.t17 65.8183
R2909 GNDA.n731 GNDA.t17 65.8183
R2910 GNDA.n780 GNDA.t17 65.8183
R2911 GNDA.n770 GNDA.t17 65.8183
R2912 GNDA.n768 GNDA.t17 65.8183
R2913 GNDA.n754 GNDA.t17 65.8183
R2914 GNDA.t24 GNDA.n155 65.8183
R2915 GNDA.t24 GNDA.n154 65.8183
R2916 GNDA.t24 GNDA.n153 65.8183
R2917 GNDA.t24 GNDA.n152 65.8183
R2918 GNDA.t24 GNDA.n148 65.8183
R2919 GNDA.t24 GNDA.n146 65.8183
R2920 GNDA.t24 GNDA.n144 65.8183
R2921 GNDA.t24 GNDA.n1928 65.8183
R2922 GNDA.t24 GNDA.n159 65.8183
R2923 GNDA.t24 GNDA.n158 65.8183
R2924 GNDA.t24 GNDA.n157 65.8183
R2925 GNDA.t24 GNDA.n149 65.8183
R2926 GNDA.t24 GNDA.n147 65.8183
R2927 GNDA.t24 GNDA.n145 65.8183
R2928 GNDA.t24 GNDA.n143 65.8183
R2929 GNDA.n959 GNDA.t19 65.8183
R2930 GNDA.n865 GNDA.t19 65.8183
R2931 GNDA.n966 GNDA.t19 65.8183
R2932 GNDA.n969 GNDA.t19 65.8183
R2933 GNDA.n950 GNDA.t19 65.8183
R2934 GNDA.n944 GNDA.t19 65.8183
R2935 GNDA.n942 GNDA.t19 65.8183
R2936 GNDA.n920 GNDA.t19 65.8183
R2937 GNDA.n926 GNDA.t19 65.8183
R2938 GNDA.n928 GNDA.t19 65.8183
R2939 GNDA.n934 GNDA.t19 65.8183
R2940 GNDA.n892 GNDA.t19 65.8183
R2941 GNDA.n899 GNDA.t19 65.8183
R2942 GNDA.n885 GNDA.t19 65.8183
R2943 GNDA.n910 GNDA.t19 65.8183
R2944 GNDA.t15 GNDA.n497 65.8183
R2945 GNDA.t15 GNDA.n496 65.8183
R2946 GNDA.t15 GNDA.n495 65.8183
R2947 GNDA.t15 GNDA.n494 65.8183
R2948 GNDA.t15 GNDA.n490 65.8183
R2949 GNDA.t15 GNDA.n488 65.8183
R2950 GNDA.t15 GNDA.n486 65.8183
R2951 GNDA.t15 GNDA.n502 65.8183
R2952 GNDA.t15 GNDA.n501 65.8183
R2953 GNDA.t15 GNDA.n500 65.8183
R2954 GNDA.t15 GNDA.n499 65.8183
R2955 GNDA.n654 GNDA.t15 65.8183
R2956 GNDA.t15 GNDA.n489 65.8183
R2957 GNDA.t15 GNDA.n487 65.8183
R2958 GNDA.t15 GNDA.n485 65.8183
R2959 GNDA.t21 GNDA.n1279 65.8183
R2960 GNDA.t21 GNDA.n1278 65.8183
R2961 GNDA.t21 GNDA.n1277 65.8183
R2962 GNDA.t21 GNDA.n1276 65.8183
R2963 GNDA.t21 GNDA.n1272 65.8183
R2964 GNDA.t21 GNDA.n1270 65.8183
R2965 GNDA.t21 GNDA.n1268 65.8183
R2966 GNDA.t21 GNDA.n1374 65.8183
R2967 GNDA.t21 GNDA.n1283 65.8183
R2968 GNDA.t21 GNDA.n1282 65.8183
R2969 GNDA.t21 GNDA.n1281 65.8183
R2970 GNDA.t21 GNDA.n1273 65.8183
R2971 GNDA.t21 GNDA.n1271 65.8183
R2972 GNDA.t21 GNDA.n1269 65.8183
R2973 GNDA.t21 GNDA.n1267 65.8183
R2974 GNDA.n395 GNDA.t18 65.8183
R2975 GNDA.n300 GNDA.t18 65.8183
R2976 GNDA.n402 GNDA.t18 65.8183
R2977 GNDA.n405 GNDA.t18 65.8183
R2978 GNDA.n386 GNDA.t18 65.8183
R2979 GNDA.n380 GNDA.t18 65.8183
R2980 GNDA.n378 GNDA.t18 65.8183
R2981 GNDA.n356 GNDA.t18 65.8183
R2982 GNDA.n362 GNDA.t18 65.8183
R2983 GNDA.n364 GNDA.t18 65.8183
R2984 GNDA.n370 GNDA.t18 65.8183
R2985 GNDA.n328 GNDA.t18 65.8183
R2986 GNDA.n335 GNDA.t18 65.8183
R2987 GNDA.n321 GNDA.t18 65.8183
R2988 GNDA.n346 GNDA.t18 65.8183
R2989 GNDA.t23 GNDA.n1103 65.8183
R2990 GNDA.t23 GNDA.n1101 65.8183
R2991 GNDA.t23 GNDA.n1099 65.8183
R2992 GNDA.t23 GNDA.n1097 65.8183
R2993 GNDA.n1745 GNDA.t22 65.8183
R2994 GNDA.n1760 GNDA.t22 65.8183
R2995 GNDA.n1754 GNDA.t22 65.8183
R2996 GNDA.n1752 GNDA.t22 65.8183
R2997 GNDA.n1773 GNDA.t22 65.8183
R2998 GNDA.n1775 GNDA.t22 65.8183
R2999 GNDA.n1781 GNDA.t22 65.8183
R3000 GNDA.n1735 GNDA.t22 65.8183
R3001 GNDA.n1797 GNDA.t22 65.8183
R3002 GNDA.n1791 GNDA.t22 65.8183
R3003 GNDA.n1789 GNDA.t22 65.8183
R3004 GNDA.n2066 GNDA.t22 65.8183
R3005 GNDA.n2063 GNDA.t22 65.8183
R3006 GNDA.n2060 GNDA.t22 65.8183
R3007 GNDA.n1803 GNDA.t22 65.8183
R3008 GNDA.n1641 GNDA.t20 65.8183
R3009 GNDA.n1639 GNDA.t20 65.8183
R3010 GNDA.n1653 GNDA.t20 65.8183
R3011 GNDA.n1612 GNDA.t20 65.8183
R3012 GNDA.t6 GNDA.t14 64.8893
R3013 GNDA.t14 GNDA.t3 64.8893
R3014 GNDA.n1723 GNDA.t31 63.7686
R3015 GNDA.n1857 GNDA.t16 63.7686
R3016 GNDA.t29 GNDA.n1937 62.4118
R3017 GNDA.n1 GNDA.t16 32.9056
R3018 GNDA.n0 GNDA.t16 32.9056
R3019 GNDA.t16 GNDA.n1616 58.3415
R3020 GNDA.n2055 GNDA.t16 58.3415
R3021 GNDA.t16 GNDA.n66 57.9215
R3022 GNDA.t16 GNDA.n59 57.9215
R3023 GNDA.t16 GNDA.n1243 57.9215
R3024 GNDA.n414 GNDA.n413 57.1945
R3025 GNDA.n413 GNDA.n291 57.1945
R3026 GNDA.n979 GNDA.n977 57.1945
R3027 GNDA.n2051 GNDA.n2050 57.1945
R3028 GNDA.t10 GNDA.n6 55.628
R3029 GNDA.n1681 GNDA.t20 55.2026
R3030 GNDA.t23 GNDA.n1110 55.2026
R3031 GNDA.n725 GNDA.t17 55.2026
R3032 GNDA.t24 GNDA.n156 55.2026
R3033 GNDA.n936 GNDA.t19 55.2026
R3034 GNDA.t15 GNDA.n498 55.2026
R3035 GNDA.t21 GNDA.n1280 55.2026
R3036 GNDA.n372 GNDA.t18 55.2026
R3037 GNDA.n1783 GNDA.t22 55.2026
R3038 GNDA.n1698 GNDA.t20 54.4705
R3039 GNDA.t23 GNDA.n1105 54.4705
R3040 GNDA.n709 GNDA.t17 54.4705
R3041 GNDA.t24 GNDA.n151 54.4705
R3042 GNDA.n953 GNDA.t19 54.4705
R3043 GNDA.t15 GNDA.n492 54.4705
R3044 GNDA.t21 GNDA.n1275 54.4705
R3045 GNDA.n389 GNDA.t18 54.4705
R3046 GNDA.n1767 GNDA.t22 54.4705
R3047 GNDA.t31 GNDA.n71 54.2712
R3048 GNDA.n1938 GNDA.t29 54.2712
R3049 GNDA.n1612 GNDA.n218 53.3664
R3050 GNDA.n1654 GNDA.n1653 53.3664
R3051 GNDA.n1639 GNDA.n1614 53.3664
R3052 GNDA.n1642 GNDA.n1641 53.3664
R3053 GNDA.n1666 GNDA.n1665 53.3664
R3054 GNDA.n1671 GNDA.n1670 53.3664
R3055 GNDA.n1674 GNDA.n1673 53.3664
R3056 GNDA.n1679 GNDA.n1678 53.3664
R3057 GNDA.n1687 GNDA.n1686 53.3664
R3058 GNDA.n1690 GNDA.n1689 53.3664
R3059 GNDA.n1695 GNDA.n1694 53.3664
R3060 GNDA.n1714 GNDA.n1713 53.3664
R3061 GNDA.n1711 GNDA.n1710 53.3664
R3062 GNDA.n1706 GNDA.n206 53.3664
R3063 GNDA.n1704 GNDA.n1703 53.3664
R3064 GNDA.n1705 GNDA.n1704 53.3664
R3065 GNDA.n206 GNDA.n204 53.3664
R3066 GNDA.n1712 GNDA.n1711 53.3664
R3067 GNDA.n1715 GNDA.n1714 53.3664
R3068 GNDA.n1696 GNDA.n1695 53.3664
R3069 GNDA.n1689 GNDA.n210 53.3664
R3070 GNDA.n1688 GNDA.n1687 53.3664
R3071 GNDA.n1665 GNDA.n216 53.3664
R3072 GNDA.n1672 GNDA.n1671 53.3664
R3073 GNDA.n1673 GNDA.n214 53.3664
R3074 GNDA.n1680 GNDA.n1679 53.3664
R3075 GNDA.n1097 GNDA.n1096 53.3664
R3076 GNDA.n1127 GNDA.n1099 53.3664
R3077 GNDA.n1138 GNDA.n1101 53.3664
R3078 GNDA.n1143 GNDA.n1103 53.3664
R3079 GNDA.n1204 GNDA.n1095 53.3664
R3080 GNDA.n1114 GNDA.n1113 53.3664
R3081 GNDA.n1198 GNDA.n1112 53.3664
R3082 GNDA.n1194 GNDA.n1111 53.3664
R3083 GNDA.n1186 GNDA.n1098 53.3664
R3084 GNDA.n1182 GNDA.n1100 53.3664
R3085 GNDA.n1178 GNDA.n1102 53.3664
R3086 GNDA.n1157 GNDA.n1106 53.3664
R3087 GNDA.n1161 GNDA.n1107 53.3664
R3088 GNDA.n1165 GNDA.n1108 53.3664
R3089 GNDA.n1169 GNDA.n1109 53.3664
R3090 GNDA.n1166 GNDA.n1109 53.3664
R3091 GNDA.n1162 GNDA.n1108 53.3664
R3092 GNDA.n1158 GNDA.n1107 53.3664
R3093 GNDA.n1154 GNDA.n1106 53.3664
R3094 GNDA.n1175 GNDA.n1102 53.3664
R3095 GNDA.n1179 GNDA.n1100 53.3664
R3096 GNDA.n1183 GNDA.n1098 53.3664
R3097 GNDA.n1204 GNDA.n1203 53.3664
R3098 GNDA.n1199 GNDA.n1113 53.3664
R3099 GNDA.n1195 GNDA.n1112 53.3664
R3100 GNDA.n1191 GNDA.n1111 53.3664
R3101 GNDA.n755 GNDA.n754 53.3664
R3102 GNDA.n768 GNDA.n767 53.3664
R3103 GNDA.n771 GNDA.n770 53.3664
R3104 GNDA.n780 GNDA.n779 53.3664
R3105 GNDA.n741 GNDA.n679 53.3664
R3106 GNDA.n740 GNDA.n739 53.3664
R3107 GNDA.n733 GNDA.n681 53.3664
R3108 GNDA.n732 GNDA.n731 53.3664
R3109 GNDA.n724 GNDA.n723 53.3664
R3110 GNDA.n717 GNDA.n685 53.3664
R3111 GNDA.n716 GNDA.n715 53.3664
R3112 GNDA.n695 GNDA.n694 53.3664
R3113 GNDA.n696 GNDA.n691 53.3664
R3114 GNDA.n703 GNDA.n702 53.3664
R3115 GNDA.n707 GNDA.n689 53.3664
R3116 GNDA.n704 GNDA.n689 53.3664
R3117 GNDA.n702 GNDA.n701 53.3664
R3118 GNDA.n697 GNDA.n696 53.3664
R3119 GNDA.n694 GNDA.n670 53.3664
R3120 GNDA.n715 GNDA.n714 53.3664
R3121 GNDA.n718 GNDA.n717 53.3664
R3122 GNDA.n723 GNDA.n722 53.3664
R3123 GNDA.n742 GNDA.n741 53.3664
R3124 GNDA.n739 GNDA.n738 53.3664
R3125 GNDA.n734 GNDA.n733 53.3664
R3126 GNDA.n731 GNDA.n730 53.3664
R3127 GNDA.n781 GNDA.n780 53.3664
R3128 GNDA.n770 GNDA.n671 53.3664
R3129 GNDA.n769 GNDA.n768 53.3664
R3130 GNDA.n754 GNDA.n675 53.3664
R3131 GNDA.n143 GNDA.n142 53.3664
R3132 GNDA.n176 GNDA.n145 53.3664
R3133 GNDA.n1862 GNDA.n147 53.3664
R3134 GNDA.n1867 GNDA.n149 53.3664
R3135 GNDA.n1928 GNDA.n141 53.3664
R3136 GNDA.n160 GNDA.n159 53.3664
R3137 GNDA.n1922 GNDA.n158 53.3664
R3138 GNDA.n1918 GNDA.n157 53.3664
R3139 GNDA.n1910 GNDA.n144 53.3664
R3140 GNDA.n1906 GNDA.n146 53.3664
R3141 GNDA.n1902 GNDA.n148 53.3664
R3142 GNDA.n1881 GNDA.n152 53.3664
R3143 GNDA.n1885 GNDA.n153 53.3664
R3144 GNDA.n1889 GNDA.n154 53.3664
R3145 GNDA.n1893 GNDA.n155 53.3664
R3146 GNDA.n1890 GNDA.n155 53.3664
R3147 GNDA.n1886 GNDA.n154 53.3664
R3148 GNDA.n1882 GNDA.n153 53.3664
R3149 GNDA.n1878 GNDA.n152 53.3664
R3150 GNDA.n1899 GNDA.n148 53.3664
R3151 GNDA.n1903 GNDA.n146 53.3664
R3152 GNDA.n1907 GNDA.n144 53.3664
R3153 GNDA.n1928 GNDA.n1927 53.3664
R3154 GNDA.n1923 GNDA.n159 53.3664
R3155 GNDA.n1919 GNDA.n158 53.3664
R3156 GNDA.n1915 GNDA.n157 53.3664
R3157 GNDA.n1877 GNDA.n149 53.3664
R3158 GNDA.n1866 GNDA.n147 53.3664
R3159 GNDA.n1861 GNDA.n145 53.3664
R3160 GNDA.n175 GNDA.n143 53.3664
R3161 GNDA.n910 GNDA.n877 53.3664
R3162 GNDA.n909 GNDA.n885 53.3664
R3163 GNDA.n899 GNDA.n898 53.3664
R3164 GNDA.n895 GNDA.n892 53.3664
R3165 GNDA.n921 GNDA.n920 53.3664
R3166 GNDA.n926 GNDA.n925 53.3664
R3167 GNDA.n929 GNDA.n928 53.3664
R3168 GNDA.n934 GNDA.n933 53.3664
R3169 GNDA.n942 GNDA.n941 53.3664
R3170 GNDA.n945 GNDA.n944 53.3664
R3171 GNDA.n950 GNDA.n949 53.3664
R3172 GNDA.n969 GNDA.n968 53.3664
R3173 GNDA.n966 GNDA.n965 53.3664
R3174 GNDA.n961 GNDA.n865 53.3664
R3175 GNDA.n959 GNDA.n958 53.3664
R3176 GNDA.n960 GNDA.n959 53.3664
R3177 GNDA.n865 GNDA.n863 53.3664
R3178 GNDA.n967 GNDA.n966 53.3664
R3179 GNDA.n970 GNDA.n969 53.3664
R3180 GNDA.n951 GNDA.n950 53.3664
R3181 GNDA.n944 GNDA.n869 53.3664
R3182 GNDA.n943 GNDA.n942 53.3664
R3183 GNDA.n920 GNDA.n875 53.3664
R3184 GNDA.n927 GNDA.n926 53.3664
R3185 GNDA.n928 GNDA.n873 53.3664
R3186 GNDA.n935 GNDA.n934 53.3664
R3187 GNDA.n892 GNDA.n861 53.3664
R3188 GNDA.n900 GNDA.n899 53.3664
R3189 GNDA.n896 GNDA.n885 53.3664
R3190 GNDA.n911 GNDA.n910 53.3664
R3191 GNDA.n504 GNDA.n485 53.3664
R3192 GNDA.n644 GNDA.n487 53.3664
R3193 GNDA.n634 GNDA.n489 53.3664
R3194 GNDA.n655 GNDA.n654 53.3664
R3195 GNDA.n503 GNDA.n502 53.3664
R3196 GNDA.n618 GNDA.n501 53.3664
R3197 GNDA.n614 GNDA.n500 53.3664
R3198 GNDA.n610 GNDA.n499 53.3664
R3199 GNDA.n602 GNDA.n486 53.3664
R3200 GNDA.n598 GNDA.n488 53.3664
R3201 GNDA.n594 GNDA.n490 53.3664
R3202 GNDA.n573 GNDA.n494 53.3664
R3203 GNDA.n577 GNDA.n495 53.3664
R3204 GNDA.n581 GNDA.n496 53.3664
R3205 GNDA.n585 GNDA.n497 53.3664
R3206 GNDA.n582 GNDA.n497 53.3664
R3207 GNDA.n578 GNDA.n496 53.3664
R3208 GNDA.n574 GNDA.n495 53.3664
R3209 GNDA.n494 GNDA.n493 53.3664
R3210 GNDA.n591 GNDA.n490 53.3664
R3211 GNDA.n595 GNDA.n488 53.3664
R3212 GNDA.n599 GNDA.n486 53.3664
R3213 GNDA.n619 GNDA.n502 53.3664
R3214 GNDA.n615 GNDA.n501 53.3664
R3215 GNDA.n611 GNDA.n500 53.3664
R3216 GNDA.n607 GNDA.n499 53.3664
R3217 GNDA.n654 GNDA.n484 53.3664
R3218 GNDA.n489 GNDA.n483 53.3664
R3219 GNDA.n633 GNDA.n487 53.3664
R3220 GNDA.n645 GNDA.n485 53.3664
R3221 GNDA.n1267 GNDA.n1266 53.3664
R3222 GNDA.n1296 GNDA.n1269 53.3664
R3223 GNDA.n1307 GNDA.n1271 53.3664
R3224 GNDA.n1312 GNDA.n1273 53.3664
R3225 GNDA.n1374 GNDA.n1265 53.3664
R3226 GNDA.n1284 GNDA.n1283 53.3664
R3227 GNDA.n1368 GNDA.n1282 53.3664
R3228 GNDA.n1364 GNDA.n1281 53.3664
R3229 GNDA.n1356 GNDA.n1268 53.3664
R3230 GNDA.n1352 GNDA.n1270 53.3664
R3231 GNDA.n1348 GNDA.n1272 53.3664
R3232 GNDA.n1327 GNDA.n1276 53.3664
R3233 GNDA.n1331 GNDA.n1277 53.3664
R3234 GNDA.n1335 GNDA.n1278 53.3664
R3235 GNDA.n1339 GNDA.n1279 53.3664
R3236 GNDA.n1336 GNDA.n1279 53.3664
R3237 GNDA.n1332 GNDA.n1278 53.3664
R3238 GNDA.n1328 GNDA.n1277 53.3664
R3239 GNDA.n1324 GNDA.n1276 53.3664
R3240 GNDA.n1345 GNDA.n1272 53.3664
R3241 GNDA.n1349 GNDA.n1270 53.3664
R3242 GNDA.n1353 GNDA.n1268 53.3664
R3243 GNDA.n1374 GNDA.n1373 53.3664
R3244 GNDA.n1369 GNDA.n1283 53.3664
R3245 GNDA.n1365 GNDA.n1282 53.3664
R3246 GNDA.n1361 GNDA.n1281 53.3664
R3247 GNDA.n1323 GNDA.n1273 53.3664
R3248 GNDA.n1311 GNDA.n1271 53.3664
R3249 GNDA.n1306 GNDA.n1269 53.3664
R3250 GNDA.n1295 GNDA.n1267 53.3664
R3251 GNDA.n346 GNDA.n312 53.3664
R3252 GNDA.n345 GNDA.n321 53.3664
R3253 GNDA.n335 GNDA.n334 53.3664
R3254 GNDA.n331 GNDA.n328 53.3664
R3255 GNDA.n357 GNDA.n356 53.3664
R3256 GNDA.n362 GNDA.n361 53.3664
R3257 GNDA.n365 GNDA.n364 53.3664
R3258 GNDA.n370 GNDA.n369 53.3664
R3259 GNDA.n378 GNDA.n377 53.3664
R3260 GNDA.n381 GNDA.n380 53.3664
R3261 GNDA.n386 GNDA.n385 53.3664
R3262 GNDA.n405 GNDA.n404 53.3664
R3263 GNDA.n402 GNDA.n401 53.3664
R3264 GNDA.n397 GNDA.n300 53.3664
R3265 GNDA.n395 GNDA.n394 53.3664
R3266 GNDA.n396 GNDA.n395 53.3664
R3267 GNDA.n300 GNDA.n298 53.3664
R3268 GNDA.n403 GNDA.n402 53.3664
R3269 GNDA.n406 GNDA.n405 53.3664
R3270 GNDA.n387 GNDA.n386 53.3664
R3271 GNDA.n380 GNDA.n304 53.3664
R3272 GNDA.n379 GNDA.n378 53.3664
R3273 GNDA.n356 GNDA.n310 53.3664
R3274 GNDA.n363 GNDA.n362 53.3664
R3275 GNDA.n364 GNDA.n308 53.3664
R3276 GNDA.n371 GNDA.n370 53.3664
R3277 GNDA.n328 GNDA.n296 53.3664
R3278 GNDA.n336 GNDA.n335 53.3664
R3279 GNDA.n332 GNDA.n321 53.3664
R3280 GNDA.n347 GNDA.n346 53.3664
R3281 GNDA.n1153 GNDA.n1103 53.3664
R3282 GNDA.n1142 GNDA.n1101 53.3664
R3283 GNDA.n1137 GNDA.n1099 53.3664
R3284 GNDA.n1126 GNDA.n1097 53.3664
R3285 GNDA.n1809 GNDA.n1803 53.3664
R3286 GNDA.n2060 GNDA.n2059 53.3664
R3287 GNDA.n2063 GNDA.n2062 53.3664
R3288 GNDA.n2066 GNDA.n2065 53.3664
R3289 GNDA.n1802 GNDA.n1735 53.3664
R3290 GNDA.n1798 GNDA.n1797 53.3664
R3291 GNDA.n1791 GNDA.n1737 53.3664
R3292 GNDA.n1790 GNDA.n1789 53.3664
R3293 GNDA.n1782 GNDA.n1781 53.3664
R3294 GNDA.n1775 GNDA.n1741 53.3664
R3295 GNDA.n1774 GNDA.n1773 53.3664
R3296 GNDA.n1753 GNDA.n1752 53.3664
R3297 GNDA.n1754 GNDA.n1747 53.3664
R3298 GNDA.n1761 GNDA.n1760 53.3664
R3299 GNDA.n1765 GNDA.n1745 53.3664
R3300 GNDA.n1762 GNDA.n1745 53.3664
R3301 GNDA.n1760 GNDA.n1759 53.3664
R3302 GNDA.n1755 GNDA.n1754 53.3664
R3303 GNDA.n1752 GNDA.n12 53.3664
R3304 GNDA.n1773 GNDA.n1772 53.3664
R3305 GNDA.n1776 GNDA.n1775 53.3664
R3306 GNDA.n1781 GNDA.n1780 53.3664
R3307 GNDA.n1799 GNDA.n1735 53.3664
R3308 GNDA.n1797 GNDA.n1796 53.3664
R3309 GNDA.n1792 GNDA.n1791 53.3664
R3310 GNDA.n1789 GNDA.n1788 53.3664
R3311 GNDA.n2067 GNDA.n2066 53.3664
R3312 GNDA.n2064 GNDA.n2063 53.3664
R3313 GNDA.n2061 GNDA.n2060 53.3664
R3314 GNDA.n1803 GNDA.n15 53.3664
R3315 GNDA.n1641 GNDA.n202 53.3664
R3316 GNDA.n1640 GNDA.n1639 53.3664
R3317 GNDA.n1653 GNDA.n1652 53.3664
R3318 GNDA.n1613 GNDA.n1612 53.3664
R3319 GNDA.n1817 GNDA.n1814 50.2009
R3320 GNDA.t36 GNDA.n1856 50.2009
R3321 GNDA.n2027 GNDA.t16 47.6748
R3322 GNDA.t16 GNDA.n65 47.6748
R3323 GNDA.n1420 GNDA.t16 47.1828
R3324 GNDA.t16 GNDA.n1527 47.1828
R3325 GNDA.t16 GNDA.n58 47.1828
R3326 GNDA.n2053 GNDA.t0 45.4226
R3327 GNDA.n1658 GNDA.t35 44.7739
R3328 GNDA.n1827 GNDA.n7 44.7739
R3329 GNDA.t16 GNDA.n1419 43.1673
R3330 GNDA.t16 GNDA.n248 43.1673
R3331 GNDA.t16 GNDA.n57 43.1673
R3332 GNDA.t16 GNDA.t5 41.9433
R3333 GNDA.t16 GNDA.n23 41.0967
R3334 GNDA.n1648 GNDA.n1633 36.6332
R3335 GNDA.n1846 GNDA.n1845 33.0535
R3336 GNDA.n1628 GNDA.n191 32.3962
R3337 GNDA.t16 GNDA.t11 31.9569
R3338 GNDA.n1855 GNDA.n181 31.2062
R3339 GNDA.n1701 GNDA.n1700 27.5561
R3340 GNDA.n1173 GNDA.n1171 27.5561
R3341 GNDA.n711 GNDA.n688 27.5561
R3342 GNDA.n1897 GNDA.n1895 27.5561
R3343 GNDA.n956 GNDA.n955 27.5561
R3344 GNDA.n589 GNDA.n587 27.5561
R3345 GNDA.n1343 GNDA.n1341 27.5561
R3346 GNDA.n392 GNDA.n391 27.5561
R3347 GNDA.n1769 GNDA.n1744 27.5561
R3348 GNDA.n1633 GNDA.t16 27.1359
R3349 GNDA.t16 GNDA.n1855 27.1359
R3350 GNDA.n1051 GNDA.n1 8.60107
R3351 GNDA.n1476 GNDA.n0 8.60107
R3352 GNDA.n1684 GNDA.n1683 26.6672
R3353 GNDA.n1189 GNDA.n1188 26.6672
R3354 GNDA.n728 GNDA.n727 26.6672
R3355 GNDA.n1913 GNDA.n1912 26.6672
R3356 GNDA.n939 GNDA.n938 26.6672
R3357 GNDA.n605 GNDA.n604 26.6672
R3358 GNDA.n1359 GNDA.n1358 26.6672
R3359 GNDA.n375 GNDA.n374 26.6672
R3360 GNDA.n1786 GNDA.n1785 26.6672
R3361 GNDA.n187 GNDA.n186 25.3679
R3362 GNDA.n1382 GNDA.t2 23.9678
R3363 GNDA.t16 GNDA.n55 20.0781
R3364 GNDA.n1581 GNDA.n1580 17.455
R3365 GNDA.n548 GNDA.n547 17.455
R3366 GNDA.n1408 GNDA.n1407 17.455
R3367 GNDA.n2031 GNDA.n31 17.0672
R3368 GNDA.n1003 GNDA.n850 17.0672
R3369 GNDA.n438 GNDA.n285 17.0672
R3370 GNDA.n254 GNDA.n253 16.9605
R3371 GNDA.n841 GNDA.n275 16.7235
R3372 GNDA.n1048 GNDA.n99 16.7235
R3373 GNDA.n664 GNDA.n98 16.7235
R3374 GNDA.n1474 GNDA.n1090 16.7235
R3375 GNDA.n1716 GNDA.n201 16.0005
R3376 GNDA.n203 GNDA.n201 16.0005
R3377 GNDA.n1709 GNDA.n203 16.0005
R3378 GNDA.n1709 GNDA.n1708 16.0005
R3379 GNDA.n1708 GNDA.n1707 16.0005
R3380 GNDA.n1707 GNDA.n205 16.0005
R3381 GNDA.n1702 GNDA.n205 16.0005
R3382 GNDA.n1702 GNDA.n1701 16.0005
R3383 GNDA.n1685 GNDA.n1684 16.0005
R3384 GNDA.n1685 GNDA.n211 16.0005
R3385 GNDA.n1691 GNDA.n211 16.0005
R3386 GNDA.n1692 GNDA.n1691 16.0005
R3387 GNDA.n1693 GNDA.n1692 16.0005
R3388 GNDA.n1693 GNDA.n209 16.0005
R3389 GNDA.n209 GNDA.n208 16.0005
R3390 GNDA.n1700 GNDA.n208 16.0005
R3391 GNDA.n1668 GNDA.n1667 16.0005
R3392 GNDA.n1669 GNDA.n1668 16.0005
R3393 GNDA.n1669 GNDA.n215 16.0005
R3394 GNDA.n1675 GNDA.n215 16.0005
R3395 GNDA.n1676 GNDA.n1675 16.0005
R3396 GNDA.n1677 GNDA.n1676 16.0005
R3397 GNDA.n1677 GNDA.n213 16.0005
R3398 GNDA.n1683 GNDA.n213 16.0005
R3399 GNDA.n1156 GNDA.n1155 16.0005
R3400 GNDA.n1159 GNDA.n1156 16.0005
R3401 GNDA.n1160 GNDA.n1159 16.0005
R3402 GNDA.n1163 GNDA.n1160 16.0005
R3403 GNDA.n1164 GNDA.n1163 16.0005
R3404 GNDA.n1167 GNDA.n1164 16.0005
R3405 GNDA.n1168 GNDA.n1167 16.0005
R3406 GNDA.n1171 GNDA.n1168 16.0005
R3407 GNDA.n1188 GNDA.n1185 16.0005
R3408 GNDA.n1185 GNDA.n1184 16.0005
R3409 GNDA.n1184 GNDA.n1181 16.0005
R3410 GNDA.n1181 GNDA.n1180 16.0005
R3411 GNDA.n1180 GNDA.n1177 16.0005
R3412 GNDA.n1177 GNDA.n1176 16.0005
R3413 GNDA.n1176 GNDA.n1174 16.0005
R3414 GNDA.n1174 GNDA.n1173 16.0005
R3415 GNDA.n1202 GNDA.n1115 16.0005
R3416 GNDA.n1202 GNDA.n1201 16.0005
R3417 GNDA.n1201 GNDA.n1200 16.0005
R3418 GNDA.n1200 GNDA.n1197 16.0005
R3419 GNDA.n1197 GNDA.n1196 16.0005
R3420 GNDA.n1196 GNDA.n1193 16.0005
R3421 GNDA.n1193 GNDA.n1192 16.0005
R3422 GNDA.n1192 GNDA.n1189 16.0005
R3423 GNDA.n693 GNDA.n692 16.0005
R3424 GNDA.n698 GNDA.n693 16.0005
R3425 GNDA.n699 GNDA.n698 16.0005
R3426 GNDA.n700 GNDA.n699 16.0005
R3427 GNDA.n700 GNDA.n690 16.0005
R3428 GNDA.n705 GNDA.n690 16.0005
R3429 GNDA.n706 GNDA.n705 16.0005
R3430 GNDA.n706 GNDA.n688 16.0005
R3431 GNDA.n727 GNDA.n684 16.0005
R3432 GNDA.n721 GNDA.n684 16.0005
R3433 GNDA.n721 GNDA.n720 16.0005
R3434 GNDA.n720 GNDA.n719 16.0005
R3435 GNDA.n719 GNDA.n686 16.0005
R3436 GNDA.n713 GNDA.n686 16.0005
R3437 GNDA.n713 GNDA.n712 16.0005
R3438 GNDA.n712 GNDA.n711 16.0005
R3439 GNDA.n744 GNDA.n743 16.0005
R3440 GNDA.n743 GNDA.n680 16.0005
R3441 GNDA.n737 GNDA.n680 16.0005
R3442 GNDA.n737 GNDA.n736 16.0005
R3443 GNDA.n736 GNDA.n735 16.0005
R3444 GNDA.n735 GNDA.n682 16.0005
R3445 GNDA.n729 GNDA.n682 16.0005
R3446 GNDA.n729 GNDA.n728 16.0005
R3447 GNDA.n1880 GNDA.n1879 16.0005
R3448 GNDA.n1883 GNDA.n1880 16.0005
R3449 GNDA.n1884 GNDA.n1883 16.0005
R3450 GNDA.n1887 GNDA.n1884 16.0005
R3451 GNDA.n1888 GNDA.n1887 16.0005
R3452 GNDA.n1891 GNDA.n1888 16.0005
R3453 GNDA.n1892 GNDA.n1891 16.0005
R3454 GNDA.n1895 GNDA.n1892 16.0005
R3455 GNDA.n1912 GNDA.n1909 16.0005
R3456 GNDA.n1909 GNDA.n1908 16.0005
R3457 GNDA.n1908 GNDA.n1905 16.0005
R3458 GNDA.n1905 GNDA.n1904 16.0005
R3459 GNDA.n1904 GNDA.n1901 16.0005
R3460 GNDA.n1901 GNDA.n1900 16.0005
R3461 GNDA.n1900 GNDA.n1898 16.0005
R3462 GNDA.n1898 GNDA.n1897 16.0005
R3463 GNDA.n1926 GNDA.n139 16.0005
R3464 GNDA.n1926 GNDA.n1925 16.0005
R3465 GNDA.n1925 GNDA.n1924 16.0005
R3466 GNDA.n1924 GNDA.n1921 16.0005
R3467 GNDA.n1921 GNDA.n1920 16.0005
R3468 GNDA.n1920 GNDA.n1917 16.0005
R3469 GNDA.n1917 GNDA.n1916 16.0005
R3470 GNDA.n1916 GNDA.n1913 16.0005
R3471 GNDA.n971 GNDA.n860 16.0005
R3472 GNDA.n862 GNDA.n860 16.0005
R3473 GNDA.n964 GNDA.n862 16.0005
R3474 GNDA.n964 GNDA.n963 16.0005
R3475 GNDA.n963 GNDA.n962 16.0005
R3476 GNDA.n962 GNDA.n864 16.0005
R3477 GNDA.n957 GNDA.n864 16.0005
R3478 GNDA.n957 GNDA.n956 16.0005
R3479 GNDA.n940 GNDA.n939 16.0005
R3480 GNDA.n940 GNDA.n870 16.0005
R3481 GNDA.n946 GNDA.n870 16.0005
R3482 GNDA.n947 GNDA.n946 16.0005
R3483 GNDA.n948 GNDA.n947 16.0005
R3484 GNDA.n948 GNDA.n868 16.0005
R3485 GNDA.n868 GNDA.n867 16.0005
R3486 GNDA.n955 GNDA.n867 16.0005
R3487 GNDA.n923 GNDA.n922 16.0005
R3488 GNDA.n924 GNDA.n923 16.0005
R3489 GNDA.n924 GNDA.n874 16.0005
R3490 GNDA.n930 GNDA.n874 16.0005
R3491 GNDA.n931 GNDA.n930 16.0005
R3492 GNDA.n932 GNDA.n931 16.0005
R3493 GNDA.n932 GNDA.n872 16.0005
R3494 GNDA.n938 GNDA.n872 16.0005
R3495 GNDA.n572 GNDA.n479 16.0005
R3496 GNDA.n575 GNDA.n572 16.0005
R3497 GNDA.n576 GNDA.n575 16.0005
R3498 GNDA.n579 GNDA.n576 16.0005
R3499 GNDA.n580 GNDA.n579 16.0005
R3500 GNDA.n583 GNDA.n580 16.0005
R3501 GNDA.n584 GNDA.n583 16.0005
R3502 GNDA.n587 GNDA.n584 16.0005
R3503 GNDA.n604 GNDA.n601 16.0005
R3504 GNDA.n601 GNDA.n600 16.0005
R3505 GNDA.n600 GNDA.n597 16.0005
R3506 GNDA.n597 GNDA.n596 16.0005
R3507 GNDA.n596 GNDA.n593 16.0005
R3508 GNDA.n593 GNDA.n592 16.0005
R3509 GNDA.n592 GNDA.n590 16.0005
R3510 GNDA.n590 GNDA.n589 16.0005
R3511 GNDA.n621 GNDA.n620 16.0005
R3512 GNDA.n620 GNDA.n617 16.0005
R3513 GNDA.n617 GNDA.n616 16.0005
R3514 GNDA.n616 GNDA.n613 16.0005
R3515 GNDA.n613 GNDA.n612 16.0005
R3516 GNDA.n612 GNDA.n609 16.0005
R3517 GNDA.n609 GNDA.n608 16.0005
R3518 GNDA.n608 GNDA.n605 16.0005
R3519 GNDA.n1326 GNDA.n1325 16.0005
R3520 GNDA.n1329 GNDA.n1326 16.0005
R3521 GNDA.n1330 GNDA.n1329 16.0005
R3522 GNDA.n1333 GNDA.n1330 16.0005
R3523 GNDA.n1334 GNDA.n1333 16.0005
R3524 GNDA.n1337 GNDA.n1334 16.0005
R3525 GNDA.n1338 GNDA.n1337 16.0005
R3526 GNDA.n1341 GNDA.n1338 16.0005
R3527 GNDA.n1358 GNDA.n1355 16.0005
R3528 GNDA.n1355 GNDA.n1354 16.0005
R3529 GNDA.n1354 GNDA.n1351 16.0005
R3530 GNDA.n1351 GNDA.n1350 16.0005
R3531 GNDA.n1350 GNDA.n1347 16.0005
R3532 GNDA.n1347 GNDA.n1346 16.0005
R3533 GNDA.n1346 GNDA.n1344 16.0005
R3534 GNDA.n1344 GNDA.n1343 16.0005
R3535 GNDA.n1372 GNDA.n1285 16.0005
R3536 GNDA.n1372 GNDA.n1371 16.0005
R3537 GNDA.n1371 GNDA.n1370 16.0005
R3538 GNDA.n1370 GNDA.n1367 16.0005
R3539 GNDA.n1367 GNDA.n1366 16.0005
R3540 GNDA.n1366 GNDA.n1363 16.0005
R3541 GNDA.n1363 GNDA.n1362 16.0005
R3542 GNDA.n1362 GNDA.n1359 16.0005
R3543 GNDA.n407 GNDA.n295 16.0005
R3544 GNDA.n297 GNDA.n295 16.0005
R3545 GNDA.n400 GNDA.n297 16.0005
R3546 GNDA.n400 GNDA.n399 16.0005
R3547 GNDA.n399 GNDA.n398 16.0005
R3548 GNDA.n398 GNDA.n299 16.0005
R3549 GNDA.n393 GNDA.n299 16.0005
R3550 GNDA.n393 GNDA.n392 16.0005
R3551 GNDA.n376 GNDA.n375 16.0005
R3552 GNDA.n376 GNDA.n305 16.0005
R3553 GNDA.n382 GNDA.n305 16.0005
R3554 GNDA.n383 GNDA.n382 16.0005
R3555 GNDA.n384 GNDA.n383 16.0005
R3556 GNDA.n384 GNDA.n303 16.0005
R3557 GNDA.n303 GNDA.n302 16.0005
R3558 GNDA.n391 GNDA.n302 16.0005
R3559 GNDA.n359 GNDA.n358 16.0005
R3560 GNDA.n360 GNDA.n359 16.0005
R3561 GNDA.n360 GNDA.n309 16.0005
R3562 GNDA.n366 GNDA.n309 16.0005
R3563 GNDA.n367 GNDA.n366 16.0005
R3564 GNDA.n368 GNDA.n367 16.0005
R3565 GNDA.n368 GNDA.n307 16.0005
R3566 GNDA.n374 GNDA.n307 16.0005
R3567 GNDA.n1751 GNDA.n1750 16.0005
R3568 GNDA.n1756 GNDA.n1751 16.0005
R3569 GNDA.n1757 GNDA.n1756 16.0005
R3570 GNDA.n1758 GNDA.n1757 16.0005
R3571 GNDA.n1758 GNDA.n1746 16.0005
R3572 GNDA.n1763 GNDA.n1746 16.0005
R3573 GNDA.n1764 GNDA.n1763 16.0005
R3574 GNDA.n1764 GNDA.n1744 16.0005
R3575 GNDA.n1785 GNDA.n1740 16.0005
R3576 GNDA.n1779 GNDA.n1740 16.0005
R3577 GNDA.n1779 GNDA.n1778 16.0005
R3578 GNDA.n1778 GNDA.n1777 16.0005
R3579 GNDA.n1777 GNDA.n1742 16.0005
R3580 GNDA.n1771 GNDA.n1742 16.0005
R3581 GNDA.n1771 GNDA.n1770 16.0005
R3582 GNDA.n1770 GNDA.n1769 16.0005
R3583 GNDA.n1801 GNDA.n1800 16.0005
R3584 GNDA.n1800 GNDA.n1736 16.0005
R3585 GNDA.n1795 GNDA.n1736 16.0005
R3586 GNDA.n1795 GNDA.n1794 16.0005
R3587 GNDA.n1794 GNDA.n1793 16.0005
R3588 GNDA.n1793 GNDA.n1738 16.0005
R3589 GNDA.n1787 GNDA.n1738 16.0005
R3590 GNDA.n1787 GNDA.n1786 16.0005
R3591 GNDA.n1830 GNDA.n1824 12.8005
R3592 GNDA.n1830 GNDA.n1829 12.8005
R3593 GNDA.n1815 GNDA.n196 12.8005
R3594 GNDA.n1819 GNDA.n196 12.8005
R3595 GNDA.n253 GNDA.n244 12.8005
R3596 GNDA.n1529 GNDA.n244 12.8005
R3597 GNDA.n820 GNDA.n462 11.6369
R3598 GNDA.n821 GNDA.n820 11.6369
R3599 GNDA.n821 GNDA.n817 11.6369
R3600 GNDA.n827 GNDA.n817 11.6369
R3601 GNDA.n828 GNDA.n827 11.6369
R3602 GNDA.n829 GNDA.n828 11.6369
R3603 GNDA.n829 GNDA.n815 11.6369
R3604 GNDA.n834 GNDA.n815 11.6369
R3605 GNDA.n835 GNDA.n834 11.6369
R3606 GNDA.n835 GNDA.n813 11.6369
R3607 GNDA.n840 GNDA.n813 11.6369
R3608 GNDA.n2000 GNDA.n1999 11.6369
R3609 GNDA.n1999 GNDA.n1996 11.6369
R3610 GNDA.n1996 GNDA.n1995 11.6369
R3611 GNDA.n1995 GNDA.n1992 11.6369
R3612 GNDA.n1992 GNDA.n1991 11.6369
R3613 GNDA.n1991 GNDA.n1988 11.6369
R3614 GNDA.n1988 GNDA.n1987 11.6369
R3615 GNDA.n1987 GNDA.n1984 11.6369
R3616 GNDA.n1984 GNDA.n1983 11.6369
R3617 GNDA.n1983 GNDA.n1980 11.6369
R3618 GNDA.n1980 GNDA.n1979 11.6369
R3619 GNDA.n121 GNDA.n120 11.6369
R3620 GNDA.n120 GNDA.n117 11.6369
R3621 GNDA.n117 GNDA.n116 11.6369
R3622 GNDA.n116 GNDA.n113 11.6369
R3623 GNDA.n113 GNDA.n112 11.6369
R3624 GNDA.n112 GNDA.n109 11.6369
R3625 GNDA.n109 GNDA.n108 11.6369
R3626 GNDA.n108 GNDA.n105 11.6369
R3627 GNDA.n105 GNDA.n104 11.6369
R3628 GNDA.n104 GNDA.n102 11.6369
R3629 GNDA.n102 GNDA.n31 11.6369
R3630 GNDA.n2047 GNDA.n2046 11.6369
R3631 GNDA.n2046 GNDA.n2045 11.6369
R3632 GNDA.n2045 GNDA.n25 11.6369
R3633 GNDA.n2040 GNDA.n25 11.6369
R3634 GNDA.n2040 GNDA.n2039 11.6369
R3635 GNDA.n2039 GNDA.n2038 11.6369
R3636 GNDA.n2038 GNDA.n28 11.6369
R3637 GNDA.n2033 GNDA.n28 11.6369
R3638 GNDA.n2033 GNDA.n2032 11.6369
R3639 GNDA.n2032 GNDA.n2031 11.6369
R3640 GNDA.n1019 GNDA.n842 11.6369
R3641 GNDA.n1019 GNDA.n1018 11.6369
R3642 GNDA.n1018 GNDA.n1017 11.6369
R3643 GNDA.n1017 GNDA.n844 11.6369
R3644 GNDA.n1012 GNDA.n844 11.6369
R3645 GNDA.n1012 GNDA.n1011 11.6369
R3646 GNDA.n1011 GNDA.n1010 11.6369
R3647 GNDA.n1010 GNDA.n847 11.6369
R3648 GNDA.n1005 GNDA.n847 11.6369
R3649 GNDA.n1005 GNDA.n1004 11.6369
R3650 GNDA.n1004 GNDA.n1003 11.6369
R3651 GNDA.n982 GNDA.n981 11.6369
R3652 GNDA.n982 GNDA.n855 11.6369
R3653 GNDA.n988 GNDA.n855 11.6369
R3654 GNDA.n989 GNDA.n988 11.6369
R3655 GNDA.n990 GNDA.n989 11.6369
R3656 GNDA.n990 GNDA.n853 11.6369
R3657 GNDA.n996 GNDA.n853 11.6369
R3658 GNDA.n997 GNDA.n996 11.6369
R3659 GNDA.n998 GNDA.n997 11.6369
R3660 GNDA.n998 GNDA.n850 11.6369
R3661 GNDA.n1580 GNDA.n1578 11.6369
R3662 GNDA.n1578 GNDA.n1575 11.6369
R3663 GNDA.n1575 GNDA.n1574 11.6369
R3664 GNDA.n1574 GNDA.n1571 11.6369
R3665 GNDA.n1571 GNDA.n1570 11.6369
R3666 GNDA.n1570 GNDA.n1567 11.6369
R3667 GNDA.n1567 GNDA.n1566 11.6369
R3668 GNDA.n1566 GNDA.n1563 11.6369
R3669 GNDA.n1563 GNDA.n1562 11.6369
R3670 GNDA.n1562 GNDA.n1559 11.6369
R3671 GNDA.n1559 GNDA.n1558 11.6369
R3672 GNDA.n1597 GNDA.n1546 11.6369
R3673 GNDA.n1597 GNDA.n1596 11.6369
R3674 GNDA.n1596 GNDA.n1595 11.6369
R3675 GNDA.n1595 GNDA.n1551 11.6369
R3676 GNDA.n1590 GNDA.n1551 11.6369
R3677 GNDA.n1590 GNDA.n1589 11.6369
R3678 GNDA.n1589 GNDA.n1588 11.6369
R3679 GNDA.n1588 GNDA.n1553 11.6369
R3680 GNDA.n1582 GNDA.n1553 11.6369
R3681 GNDA.n1582 GNDA.n1581 11.6369
R3682 GNDA.n547 GNDA.n519 11.6369
R3683 GNDA.n520 GNDA.n519 11.6369
R3684 GNDA.n540 GNDA.n520 11.6369
R3685 GNDA.n540 GNDA.n539 11.6369
R3686 GNDA.n539 GNDA.n538 11.6369
R3687 GNDA.n538 GNDA.n522 11.6369
R3688 GNDA.n533 GNDA.n522 11.6369
R3689 GNDA.n533 GNDA.n532 11.6369
R3690 GNDA.n532 GNDA.n531 11.6369
R3691 GNDA.n531 GNDA.n525 11.6369
R3692 GNDA.n525 GNDA.n463 11.6369
R3693 GNDA.n564 GNDA.n508 11.6369
R3694 GNDA.n564 GNDA.n563 11.6369
R3695 GNDA.n563 GNDA.n562 11.6369
R3696 GNDA.n562 GNDA.n512 11.6369
R3697 GNDA.n557 GNDA.n512 11.6369
R3698 GNDA.n557 GNDA.n556 11.6369
R3699 GNDA.n556 GNDA.n555 11.6369
R3700 GNDA.n555 GNDA.n514 11.6369
R3701 GNDA.n549 GNDA.n514 11.6369
R3702 GNDA.n549 GNDA.n548 11.6369
R3703 GNDA.n1409 GNDA.n1408 11.6369
R3704 GNDA.n1409 GNDA.n1247 11.6369
R3705 GNDA.n1415 GNDA.n1247 11.6369
R3706 GNDA.n1416 GNDA.n1415 11.6369
R3707 GNDA.n1417 GNDA.n1416 11.6369
R3708 GNDA.n1417 GNDA.n1231 11.6369
R3709 GNDA.n1423 GNDA.n1231 11.6369
R3710 GNDA.n1424 GNDA.n1423 11.6369
R3711 GNDA.n1425 GNDA.n1424 11.6369
R3712 GNDA.n1425 GNDA.n1227 11.6369
R3713 GNDA.n1431 GNDA.n1227 11.6369
R3714 GNDA.n1385 GNDA.n1257 11.6369
R3715 GNDA.n1392 GNDA.n1257 11.6369
R3716 GNDA.n1393 GNDA.n1392 11.6369
R3717 GNDA.n1394 GNDA.n1393 11.6369
R3718 GNDA.n1394 GNDA.n1255 11.6369
R3719 GNDA.n1399 GNDA.n1255 11.6369
R3720 GNDA.n1400 GNDA.n1399 11.6369
R3721 GNDA.n1401 GNDA.n1400 11.6369
R3722 GNDA.n1401 GNDA.n1251 11.6369
R3723 GNDA.n1407 GNDA.n1251 11.6369
R3724 GNDA.n456 GNDA.n259 11.6369
R3725 GNDA.n456 GNDA.n455 11.6369
R3726 GNDA.n455 GNDA.n454 11.6369
R3727 GNDA.n454 GNDA.n279 11.6369
R3728 GNDA.n448 GNDA.n279 11.6369
R3729 GNDA.n448 GNDA.n447 11.6369
R3730 GNDA.n447 GNDA.n446 11.6369
R3731 GNDA.n446 GNDA.n281 11.6369
R3732 GNDA.n440 GNDA.n281 11.6369
R3733 GNDA.n440 GNDA.n439 11.6369
R3734 GNDA.n439 GNDA.n438 11.6369
R3735 GNDA.n416 GNDA.n290 11.6369
R3736 GNDA.n422 GNDA.n290 11.6369
R3737 GNDA.n423 GNDA.n422 11.6369
R3738 GNDA.n424 GNDA.n423 11.6369
R3739 GNDA.n424 GNDA.n288 11.6369
R3740 GNDA.n430 GNDA.n288 11.6369
R3741 GNDA.n431 GNDA.n430 11.6369
R3742 GNDA.n432 GNDA.n431 11.6369
R3743 GNDA.n432 GNDA.n286 11.6369
R3744 GNDA.n286 GNDA.n285 11.6369
R3745 GNDA.n1437 GNDA.n1434 11.6369
R3746 GNDA.n1443 GNDA.n1437 11.6369
R3747 GNDA.n1443 GNDA.n1442 11.6369
R3748 GNDA.n1442 GNDA.n1441 11.6369
R3749 GNDA.n1441 GNDA.n1438 11.6369
R3750 GNDA.n1525 GNDA.n1524 11.6369
R3751 GNDA.n1524 GNDA.n1523 11.6369
R3752 GNDA.n1523 GNDA.n255 11.6369
R3753 GNDA.n1517 GNDA.n255 11.6369
R3754 GNDA.n1517 GNDA.n1516 11.6369
R3755 GNDA.n1627 GNDA.t32 9.6005
R3756 GNDA.n1630 GNDA.t34 9.6005
R3757 GNDA.n185 GNDA.t30 9.6005
R3758 GNDA.n1852 GNDA.t28 9.6005
R3759 GNDA.n169 GNDA.t37 9.49788
R3760 GNDA.n1871 GNDA.t4 9.49788
R3761 GNDA.t27 GNDA.n2052 9.49788
R3762 GNDA.n1832 GNDA.n1824 9.36264
R3763 GNDA.n1815 GNDA.n194 9.36264
R3764 GNDA.n253 GNDA.n242 9.36264
R3765 GNDA.n1831 GNDA.n1830 9.3005
R3766 GNDA.n1829 GNDA.n1823 9.3005
R3767 GNDA.n196 GNDA.n195 9.3005
R3768 GNDA.n1820 GNDA.n1819 9.3005
R3769 GNDA.n244 GNDA.n243 9.3005
R3770 GNDA.n1530 GNDA.n1529 9.3005
R3771 GNDA.n1544 GNDA.t33 8.14111
R3772 GNDA.t16 GNDA.t10 8.14111
R3773 GNDA.n1540 GNDA.n1539 6.98357
R3774 GNDA.n1090 GNDA.n462 6.72373
R3775 GNDA.n2000 GNDA.n98 6.72373
R3776 GNDA.n121 GNDA.n99 6.72373
R3777 GNDA.n842 GNDA.n841 6.72373
R3778 GNDA.n1515 GNDA.n259 6.72373
R3779 GNDA.n1434 GNDA.n1432 6.72373
R3780 GNDA.n841 GNDA.n840 6.20656
R3781 GNDA.n1979 GNDA.n99 6.20656
R3782 GNDA.n1558 GNDA.n98 6.20656
R3783 GNDA.n1090 GNDA.n463 6.20656
R3784 GNDA.n1432 GNDA.n1431 6.20656
R3785 GNDA.n1516 GNDA.n1515 6.20656
R3786 GNDA.n1525 GNDA.n254 6.07727
R3787 GNDA.n1853 GNDA.n186 5.81868
R3788 GNDA.n1851 GNDA.n186 5.81868
R3789 GNDA.n1438 GNDA.n254 5.5601
R3790 GNDA.n1667 GNDA.n217 5.51161
R3791 GNDA.n1115 GNDA.n1092 5.51161
R3792 GNDA.n745 GNDA.n744 5.51161
R3793 GNDA.n1932 GNDA.n139 5.51161
R3794 GNDA.n922 GNDA.n876 5.51161
R3795 GNDA.n622 GNDA.n621 5.51161
R3796 GNDA.n1285 GNDA.n1263 5.51161
R3797 GNDA.n358 GNDA.n311 5.51161
R3798 GNDA.n1801 GNDA.n1733 5.51161
R3799 GNDA.n623 GNDA.n571 5.1717
R3800 GNDA.n1384 GNDA.n1261 5.1717
R3801 GNDA.n1604 GNDA.n1603 5.1717
R3802 GNDA.n161 GNDA.n22 4.9157
R3803 GNDA.n980 GNDA.n857 4.9157
R3804 GNDA.n415 GNDA.n292 4.9157
R3805 GNDA.n1821 GNDA.n1820 4.5005
R3806 GNDA.n1833 GNDA.n1823 4.5005
R3807 GNDA.n1838 GNDA.n1837 4.5005
R3808 GNDA.n1843 GNDA.n192 4.5005
R3809 GNDA.n1845 GNDA.n1844 4.5005
R3810 GNDA.n1844 GNDA.n1843 4.5005
R3811 GNDA.n1531 GNDA.n1530 4.5005
R3812 GNDA.n1480 GNDA.n271 4.26717
R3813 GNDA.n1486 GNDA.n271 4.26717
R3814 GNDA.n1486 GNDA.n269 4.26717
R3815 GNDA.n1492 GNDA.n269 4.26717
R3816 GNDA.n1492 GNDA.n267 4.26717
R3817 GNDA.n1498 GNDA.n267 4.26717
R3818 GNDA.n1498 GNDA.n265 4.26717
R3819 GNDA.n1507 GNDA.n265 4.26717
R3820 GNDA.n1507 GNDA.n263 4.26717
R3821 GNDA.n263 GNDA.n260 4.26717
R3822 GNDA.n1514 GNDA.n260 4.26717
R3823 GNDA.n1046 GNDA.n790 4.26717
R3824 GNDA.n1041 GNDA.n790 4.26717
R3825 GNDA.n1041 GNDA.n1040 4.26717
R3826 GNDA.n1040 GNDA.n797 4.26717
R3827 GNDA.n1035 GNDA.n797 4.26717
R3828 GNDA.n1035 GNDA.n1034 4.26717
R3829 GNDA.n1034 GNDA.n1033 4.26717
R3830 GNDA.n1033 GNDA.n805 4.26717
R3831 GNDA.n1027 GNDA.n805 4.26717
R3832 GNDA.n1027 GNDA.n1026 4.26717
R3833 GNDA.n1026 GNDA.n1025 4.26717
R3834 GNDA.n1943 GNDA.n131 4.26717
R3835 GNDA.n1949 GNDA.n131 4.26717
R3836 GNDA.n1949 GNDA.n129 4.26717
R3837 GNDA.n1955 GNDA.n129 4.26717
R3838 GNDA.n1955 GNDA.n127 4.26717
R3839 GNDA.n1961 GNDA.n127 4.26717
R3840 GNDA.n1961 GNDA.n125 4.26717
R3841 GNDA.n1969 GNDA.n125 4.26717
R3842 GNDA.n1969 GNDA.n123 4.26717
R3843 GNDA.n123 GNDA.n101 4.26717
R3844 GNDA.n1976 GNDA.n101 4.26717
R3845 GNDA.n2023 GNDA.n2022 4.26717
R3846 GNDA.n2022 GNDA.n2021 4.26717
R3847 GNDA.n2021 GNDA.n2019 4.26717
R3848 GNDA.n2019 GNDA.n2016 4.26717
R3849 GNDA.n2016 GNDA.n2015 4.26717
R3850 GNDA.n2015 GNDA.n2012 4.26717
R3851 GNDA.n2012 GNDA.n2011 4.26717
R3852 GNDA.n2011 GNDA.n2008 4.26717
R3853 GNDA.n2008 GNDA.n2007 4.26717
R3854 GNDA.n2007 GNDA.n2004 4.26717
R3855 GNDA.n2004 GNDA.n2003 4.26717
R3856 GNDA.n1055 GNDA.n475 4.26717
R3857 GNDA.n1061 GNDA.n475 4.26717
R3858 GNDA.n1061 GNDA.n473 4.26717
R3859 GNDA.n1067 GNDA.n473 4.26717
R3860 GNDA.n1067 GNDA.n471 4.26717
R3861 GNDA.n1073 GNDA.n471 4.26717
R3862 GNDA.n1073 GNDA.n469 4.26717
R3863 GNDA.n1082 GNDA.n469 4.26717
R3864 GNDA.n1082 GNDA.n467 4.26717
R3865 GNDA.n467 GNDA.n464 4.26717
R3866 GNDA.n1089 GNDA.n464 4.26717
R3867 GNDA.n1472 GNDA.n1213 4.26717
R3868 GNDA.n1467 GNDA.n1213 4.26717
R3869 GNDA.n1467 GNDA.n1466 4.26717
R3870 GNDA.n1466 GNDA.n1217 4.26717
R3871 GNDA.n1461 GNDA.n1217 4.26717
R3872 GNDA.n1461 GNDA.n1460 4.26717
R3873 GNDA.n1460 GNDA.n1459 4.26717
R3874 GNDA.n1459 GNDA.n1222 4.26717
R3875 GNDA.n1453 GNDA.n1222 4.26717
R3876 GNDA.n1453 GNDA.n1452 4.26717
R3877 GNDA.n1452 GNDA.n1451 4.26717
R3878 GNDA.n1659 GNDA.t8 4.07081
R3879 GNDA.n1634 GNDA.t25 4.07081
R3880 GNDA.n1515 GNDA.n1514 3.98272
R3881 GNDA.n1025 GNDA.n841 3.98272
R3882 GNDA.n1976 GNDA.n99 3.98272
R3883 GNDA.n2003 GNDA.n98 3.98272
R3884 GNDA.n1090 GNDA.n1089 3.98272
R3885 GNDA.n1451 GNDA.n1432 3.98272
R3886 GNDA.n752 GNDA.n678 3.7893
R3887 GNDA.n758 GNDA.n756 3.7893
R3888 GNDA.n757 GNDA.n676 3.7893
R3889 GNDA.n766 GNDA.n765 3.7893
R3890 GNDA.n762 GNDA.n674 3.7893
R3891 GNDA.n777 GNDA.n672 3.7893
R3892 GNDA.n778 GNDA.n669 3.7893
R3893 GNDA.n783 GNDA.n782 3.7893
R3894 GNDA.n1930 GNDA.n140 3.7893
R3895 GNDA.n173 GNDA.n172 3.7893
R3896 GNDA.n178 GNDA.n174 3.7893
R3897 GNDA.n177 GNDA.n166 3.7893
R3898 GNDA.n1860 GNDA.n1859 3.7893
R3899 GNDA.n1869 GNDA.n1865 3.7893
R3900 GNDA.n1868 GNDA.n163 3.7893
R3901 GNDA.n1876 GNDA.n1875 3.7893
R3902 GNDA.n918 GNDA.n917 3.7893
R3903 GNDA.n913 GNDA.n879 3.7893
R3904 GNDA.n912 GNDA.n884 3.7893
R3905 GNDA.n908 GNDA.n907 3.7893
R3906 GNDA.n888 GNDA.n886 3.7893
R3907 GNDA.n901 GNDA.n891 3.7893
R3908 GNDA.n894 GNDA.n893 3.7893
R3909 GNDA.n973 GNDA.n859 3.7893
R3910 GNDA.n652 GNDA.n651 3.7893
R3911 GNDA.n647 GNDA.n506 3.7893
R3912 GNDA.n646 GNDA.n628 3.7893
R3913 GNDA.n643 GNDA.n642 3.7893
R3914 GNDA.n631 GNDA.n629 3.7893
R3915 GNDA.n636 GNDA.n482 3.7893
R3916 GNDA.n657 GNDA.n656 3.7893
R3917 GNDA.n660 GNDA.n480 3.7893
R3918 GNDA.n1376 GNDA.n1264 3.7893
R3919 GNDA.n1293 GNDA.n1292 3.7893
R3920 GNDA.n1298 GNDA.n1294 3.7893
R3921 GNDA.n1297 GNDA.n1289 3.7893
R3922 GNDA.n1305 GNDA.n1304 3.7893
R3923 GNDA.n1314 GNDA.n1310 3.7893
R3924 GNDA.n1313 GNDA.n1287 3.7893
R3925 GNDA.n1322 GNDA.n1321 3.7893
R3926 GNDA.n354 GNDA.n353 3.7893
R3927 GNDA.n349 GNDA.n314 3.7893
R3928 GNDA.n348 GNDA.n320 3.7893
R3929 GNDA.n344 GNDA.n343 3.7893
R3930 GNDA.n324 GNDA.n322 3.7893
R3931 GNDA.n337 GNDA.n327 3.7893
R3932 GNDA.n330 GNDA.n329 3.7893
R3933 GNDA.n409 GNDA.n294 3.7893
R3934 GNDA.n1206 GNDA.n1094 3.7893
R3935 GNDA.n1124 GNDA.n1123 3.7893
R3936 GNDA.n1129 GNDA.n1125 3.7893
R3937 GNDA.n1128 GNDA.n1120 3.7893
R3938 GNDA.n1136 GNDA.n1135 3.7893
R3939 GNDA.n1145 GNDA.n1141 3.7893
R3940 GNDA.n1144 GNDA.n1118 3.7893
R3941 GNDA.n1152 GNDA.n1151 3.7893
R3942 GNDA.n1811 GNDA.n1734 3.7893
R3943 GNDA.n1808 GNDA.n1807 3.7893
R3944 GNDA.n1804 GNDA.n16 3.7893
R3945 GNDA.n2058 GNDA.n2057 3.7893
R3946 GNDA.n14 GNDA.n13 3.7893
R3947 GNDA.n9 GNDA.n3 3.7893
R3948 GNDA.n2069 GNDA.n10 3.7893
R3949 GNDA.n2068 GNDA.n11 3.7893
R3950 GNDA.n1663 GNDA.n1662 3.7893
R3951 GNDA.n1609 GNDA.n220 3.7893
R3952 GNDA.n1656 GNDA.n1610 3.7893
R3953 GNDA.n1655 GNDA.n1611 3.7893
R3954 GNDA.n1651 GNDA.n1650 3.7893
R3955 GNDA.n1644 GNDA.n1637 3.7893
R3956 GNDA.n1643 GNDA.n1638 3.7893
R3957 GNDA.n1719 GNDA.n200 3.7893
R3958 GNDA.n238 GNDA.n237 3.4105
R3959 GNDA.n1539 GNDA.n234 3.4105
R3960 GNDA.n1537 GNDA.n234 3.4105
R3961 GNDA.n1539 GNDA.n1538 3.4105
R3962 GNDA.n1538 GNDA.n1537 3.4105
R3963 GNDA.n229 GNDA.n226 3.4105
R3964 GNDA.n230 GNDA.n229 3.4105
R3965 GNDA.n231 GNDA.n230 3.4105
R3966 GNDA.n773 GNDA 2.9189
R3967 GNDA.n1864 GNDA 2.9189
R3968 GNDA.n902 GNDA 2.9189
R3969 GNDA.n637 GNDA 2.9189
R3970 GNDA.n1309 GNDA 2.9189
R3971 GNDA.n338 GNDA 2.9189
R3972 GNDA.n1140 GNDA 2.9189
R3973 GNDA GNDA.n2075 2.9189
R3974 GNDA.n1636 GNDA 2.9189
R3975 GNDA.n1850 GNDA.n1849 2.86505
R3976 GNDA.n1849 GNDA.n1847 2.86505
R3977 GNDA.n1847 GNDA.n1846 2.86505
R3978 GNDA.n1851 GNDA.n1850 2.86505
R3979 GNDA.n1621 GNDA.n1620 2.86505
R3980 GNDA.n1622 GNDA.n1621 2.86505
R3981 GNDA.n1626 GNDA.n1624 2.86505
R3982 GNDA.n1629 GNDA.n1624 2.86505
R3983 GNDA.n1625 GNDA.n1622 2.86505
R3984 GNDA.n1629 GNDA.n1628 2.86505
R3985 GNDA.n1631 GNDA.n1620 2.86505
R3986 GNDA.n1626 GNDA.n1625 2.86505
R3987 GNDA.n746 GNDA.n477 2.6629
R3988 GNDA.n787 GNDA.n667 2.6629
R3989 GNDA.n1933 GNDA.n133 2.6629
R3990 GNDA.n162 GNDA.n161 2.6629
R3991 GNDA.n1047 GNDA.n788 2.6629
R3992 GNDA.n972 GNDA.n857 2.6629
R3993 GNDA.n662 GNDA.n661 2.6629
R3994 GNDA.n1286 GNDA.n1091 2.6629
R3995 GNDA.n315 GNDA.n273 2.6629
R3996 GNDA.n408 GNDA.n292 2.6629
R3997 GNDA.n1473 GNDA.n1211 2.6629
R3998 GNDA.n1117 GNDA.n1116 2.6629
R3999 GNDA.n1732 GNDA.n79 2.6629
R4000 GNDA.n1749 GNDA.n1748 2.6629
R4001 GNDA.n1718 GNDA.n1717 2.6629
R4002 GNDA.n746 GNDA.n745 2.4581
R4003 GNDA.n1047 GNDA.n787 2.4581
R4004 GNDA.n1933 GNDA.n1932 2.4581
R4005 GNDA.n876 GNDA.n788 2.4581
R4006 GNDA.n623 GNDA.n622 2.4581
R4007 GNDA.n662 GNDA.n477 2.4581
R4008 GNDA.n1263 GNDA.n1261 2.4581
R4009 GNDA.n1473 GNDA.n1091 2.4581
R4010 GNDA.n315 GNDA.n311 2.4581
R4011 GNDA.n1211 GNDA.n1092 2.4581
R4012 GNDA.n1116 GNDA.n273 2.4581
R4013 GNDA.n1733 GNDA.n1732 2.4581
R4014 GNDA.n1748 GNDA.n133 2.4581
R4015 GNDA.n1604 GNDA.n217 2.4581
R4016 GNDA.n1717 GNDA.n79 2.4581
R4017 GNDA.n1541 GNDA.n1540 2.44675
R4018 GNDA.n1540 GNDA.n223 2.44675
R4019 GNDA.n1836 GNDA.n1835 2.26187
R4020 GNDA.n1839 GNDA.n1822 2.24063
R4021 GNDA.n1840 GNDA.n193 2.24063
R4022 GNDA.n1845 GNDA.n189 2.24063
R4023 GNDA.n190 GNDA.n188 2.24063
R4024 GNDA.n1835 GNDA.n1834 2.24063
R4025 GNDA.n1842 GNDA.n1841 2.24063
R4026 GNDA.n1821 GNDA.n194 2.22018
R4027 GNDA.n1833 GNDA.n1832 2.22018
R4028 GNDA.n1531 GNDA.n242 2.22018
R4029 GNDA.n1480 GNDA.n273 2.18124
R4030 GNDA.n1047 GNDA.n1046 2.18124
R4031 GNDA.n1943 GNDA.n133 2.18124
R4032 GNDA.n2023 GNDA.n79 2.18124
R4033 GNDA.n1055 GNDA.n477 2.18124
R4034 GNDA.n1473 GNDA.n1472 2.18124
R4035 GNDA.n751 GNDA.n745 2.1509
R4036 GNDA.n1932 GNDA.n1931 2.1509
R4037 GNDA.n878 GNDA.n876 2.1509
R4038 GNDA.n622 GNDA.n505 2.1509
R4039 GNDA.n1377 GNDA.n1263 2.1509
R4040 GNDA.n313 GNDA.n311 2.1509
R4041 GNDA.n1207 GNDA.n1092 2.1509
R4042 GNDA.n1812 GNDA.n1733 2.1509
R4043 GNDA.n219 GNDA.n217 2.1509
R4044 GNDA.n1718 GNDA.n1716 2.13383
R4045 GNDA.n1155 GNDA.n1117 2.13383
R4046 GNDA.n692 GNDA.n667 2.13383
R4047 GNDA.n1879 GNDA.n162 2.13383
R4048 GNDA.n972 GNDA.n971 2.13383
R4049 GNDA.n661 GNDA.n479 2.13383
R4050 GNDA.n1325 GNDA.n1286 2.13383
R4051 GNDA.n408 GNDA.n407 2.13383
R4052 GNDA.n1750 GNDA.n1749 2.13383
R4053 GNDA.n275 GNDA.n273 2.08643
R4054 GNDA.n1048 GNDA.n1047 2.08643
R4055 GNDA.n135 GNDA.n133 2.08643
R4056 GNDA.n1725 GNDA.n79 2.08643
R4057 GNDA.n664 GNDA.n477 2.08643
R4058 GNDA.n1474 GNDA.n1473 2.08643
R4059 GNDA.n1475 GNDA.n461 1.951
R4060 GNDA.n1726 GNDA.n78 1.951
R4061 GNDA.n1050 GNDA.n476 1.951
R4062 GNDA.n1936 GNDA.n132 1.951
R4063 GNDA.n1049 GNDA.n666 1.951
R4064 GNDA.n1547 GNDA.n1545 1.951
R4065 GNDA.n570 GNDA.n507 1.951
R4066 GNDA.n1383 GNDA.n1381 1.951
R4067 GNDA.n460 GNDA.n272 1.951
R4068 GNDA.n783 GNDA.n667 1.9461
R4069 GNDA.n1875 GNDA.n162 1.9461
R4070 GNDA.n973 GNDA.n972 1.9461
R4071 GNDA.n661 GNDA.n660 1.9461
R4072 GNDA.n1321 GNDA.n1286 1.9461
R4073 GNDA.n409 GNDA.n408 1.9461
R4074 GNDA.n1151 GNDA.n1117 1.9461
R4075 GNDA.n1749 GNDA.n11 1.9461
R4076 GNDA.n1719 GNDA.n1718 1.9461
R4077 GNDA.n239 GNDA.n236 1.72394
R4078 GNDA.n240 GNDA.n239 1.70387
R4079 GNDA.n1535 GNDA.n1534 1.70194
R4080 GNDA.n235 GNDA.n224 1.70194
R4081 GNDA.n232 GNDA.n226 1.70194
R4082 GNDA.n228 GNDA.n227 1.70194
R4083 GNDA.n1536 GNDA.n236 1.69525
R4084 GNDA.n233 GNDA.n225 1.69525
R4085 GNDA.n2047 GNDA.n22 1.52512
R4086 GNDA.n981 GNDA.n980 1.52512
R4087 GNDA.n416 GNDA.n415 1.52512
R4088 GNDA.n1603 GNDA.n1546 1.42272
R4089 GNDA.n571 GNDA.n508 1.42272
R4090 GNDA.n1385 GNDA.n1384 1.42272
R4091 GNDA.n1532 GNDA.n1531 1.22446
R4092 GNDA.n1531 GNDA.n241 1.22446
R4093 GNDA.n226 GNDA.n191 1.13952
R4094 GNDA GNDA.n772 0.8709
R4095 GNDA GNDA.n1863 0.8709
R4096 GNDA.n897 GNDA 0.8709
R4097 GNDA GNDA.n635 0.8709
R4098 GNDA GNDA.n1308 0.8709
R4099 GNDA.n333 GNDA 0.8709
R4100 GNDA GNDA.n1139 0.8709
R4101 GNDA GNDA.n2 0.8709
R4102 GNDA GNDA.n1635 0.8709
R4103 GNDA.n752 GNDA.n751 0.8197
R4104 GNDA.n756 GNDA.n678 0.8197
R4105 GNDA.n758 GNDA.n757 0.8197
R4106 GNDA.n766 GNDA.n676 0.8197
R4107 GNDA.n765 GNDA.n674 0.8197
R4108 GNDA.n773 GNDA.n672 0.8197
R4109 GNDA.n778 GNDA.n777 0.8197
R4110 GNDA.n782 GNDA.n669 0.8197
R4111 GNDA.n1931 GNDA.n1930 0.8197
R4112 GNDA.n172 GNDA.n140 0.8197
R4113 GNDA.n174 GNDA.n173 0.8197
R4114 GNDA.n178 GNDA.n177 0.8197
R4115 GNDA.n1860 GNDA.n166 0.8197
R4116 GNDA.n1865 GNDA.n1864 0.8197
R4117 GNDA.n1869 GNDA.n1868 0.8197
R4118 GNDA.n1876 GNDA.n163 0.8197
R4119 GNDA.n918 GNDA.n878 0.8197
R4120 GNDA.n917 GNDA.n879 0.8197
R4121 GNDA.n913 GNDA.n912 0.8197
R4122 GNDA.n908 GNDA.n884 0.8197
R4123 GNDA.n907 GNDA.n886 0.8197
R4124 GNDA.n902 GNDA.n901 0.8197
R4125 GNDA.n894 GNDA.n891 0.8197
R4126 GNDA.n893 GNDA.n859 0.8197
R4127 GNDA.n652 GNDA.n505 0.8197
R4128 GNDA.n651 GNDA.n506 0.8197
R4129 GNDA.n647 GNDA.n646 0.8197
R4130 GNDA.n643 GNDA.n628 0.8197
R4131 GNDA.n642 GNDA.n629 0.8197
R4132 GNDA.n637 GNDA.n636 0.8197
R4133 GNDA.n656 GNDA.n482 0.8197
R4134 GNDA.n657 GNDA.n480 0.8197
R4135 GNDA.n1377 GNDA.n1376 0.8197
R4136 GNDA.n1292 GNDA.n1264 0.8197
R4137 GNDA.n1294 GNDA.n1293 0.8197
R4138 GNDA.n1298 GNDA.n1297 0.8197
R4139 GNDA.n1305 GNDA.n1289 0.8197
R4140 GNDA.n1310 GNDA.n1309 0.8197
R4141 GNDA.n1314 GNDA.n1313 0.8197
R4142 GNDA.n1322 GNDA.n1287 0.8197
R4143 GNDA.n354 GNDA.n313 0.8197
R4144 GNDA.n353 GNDA.n314 0.8197
R4145 GNDA.n349 GNDA.n348 0.8197
R4146 GNDA.n344 GNDA.n320 0.8197
R4147 GNDA.n343 GNDA.n322 0.8197
R4148 GNDA.n338 GNDA.n337 0.8197
R4149 GNDA.n330 GNDA.n327 0.8197
R4150 GNDA.n329 GNDA.n294 0.8197
R4151 GNDA.n1207 GNDA.n1206 0.8197
R4152 GNDA.n1123 GNDA.n1094 0.8197
R4153 GNDA.n1125 GNDA.n1124 0.8197
R4154 GNDA.n1129 GNDA.n1128 0.8197
R4155 GNDA.n1136 GNDA.n1120 0.8197
R4156 GNDA.n1141 GNDA.n1140 0.8197
R4157 GNDA.n1145 GNDA.n1144 0.8197
R4158 GNDA.n1152 GNDA.n1118 0.8197
R4159 GNDA.n1812 GNDA.n1811 0.8197
R4160 GNDA.n1808 GNDA.n1734 0.8197
R4161 GNDA.n1807 GNDA.n1804 0.8197
R4162 GNDA.n2058 GNDA.n16 0.8197
R4163 GNDA.n2057 GNDA.n14 0.8197
R4164 GNDA.n2075 GNDA.n3 0.8197
R4165 GNDA.n10 GNDA.n9 0.8197
R4166 GNDA.n2069 GNDA.n2068 0.8197
R4167 GNDA.n1663 GNDA.n219 0.8197
R4168 GNDA.n1662 GNDA.n220 0.8197
R4169 GNDA.n1610 GNDA.n1609 0.8197
R4170 GNDA.n1656 GNDA.n1655 0.8197
R4171 GNDA.n1651 GNDA.n1611 0.8197
R4172 GNDA.n1637 GNDA.n1636 0.8197
R4173 GNDA.n1644 GNDA.n1643 0.8197
R4174 GNDA.n1638 GNDA.n200 0.8197
R4175 GNDA.n1841 GNDA.n1840 0.71925
R4176 GNDA.n1843 GNDA.n191 0.65675
R4177 GNDA GNDA.n1536 0.580769
R4178 GNDA.n762 GNDA 0.5125
R4179 GNDA.n1859 GNDA 0.5125
R4180 GNDA GNDA.n888 0.5125
R4181 GNDA GNDA.n631 0.5125
R4182 GNDA.n1304 GNDA 0.5125
R4183 GNDA GNDA.n324 0.5125
R4184 GNDA.n1135 GNDA 0.5125
R4185 GNDA.n13 GNDA 0.5125
R4186 GNDA.n1650 GNDA 0.5125
R4187 GNDA.n1534 GNDA.n1533 0.379106
R4188 GNDA.n772 GNDA 0.3077
R4189 GNDA.n1863 GNDA 0.3077
R4190 GNDA.n897 GNDA 0.3077
R4191 GNDA.n635 GNDA 0.3077
R4192 GNDA.n1308 GNDA 0.3077
R4193 GNDA.n333 GNDA 0.3077
R4194 GNDA.n1139 GNDA 0.3077
R4195 GNDA GNDA.n2 0.3077
R4196 GNDA.n1635 GNDA 0.3077
R4197 GNDA.n1538 GNDA 0.259
R4198 GNDA.n1533 GNDA.n1532 0.234875
R4199 GNDA.n1822 GNDA.n1821 0.188
R4200 GNDA.n1834 GNDA.n1833 0.188
R4201 GNDA.n1831 GNDA.n1823 0.1255
R4202 GNDA.n1820 GNDA.n195 0.1255
R4203 GNDA.n1530 GNDA.n243 0.1255
R4204 GNDA.n1537 GNDA.n224 0.0666765
R4205 GNDA.n1539 GNDA.n224 0.0666765
R4206 GNDA.n1832 GNDA.n1831 0.0626438
R4207 GNDA.n195 GNDA.n194 0.0626438
R4208 GNDA.n243 GNDA.n242 0.0626438
R4209 GNDA.n227 GNDA.n226 0.0437692
R4210 GNDA.n1845 GNDA.n188 0.0421667
R4211 GNDA.n234 GNDA.n233 0.0402692
R4212 GNDA.n238 GNDA.n236 0.0224982
R4213 GNDA.n227 GNDA.n225 0.0224982
R4214 GNDA.n1534 GNDA.n240 0.0224982
R4215 GNDA.n240 GNDA.n238 0.0224982
R4216 GNDA.n230 GNDA.n225 0.0224982
R4217 GNDA.n1834 GNDA.n193 0.0217373
R4218 GNDA.n1839 GNDA.n1838 0.0217373
R4219 GNDA.n1841 GNDA.n189 0.0217373
R4220 GNDA.n1844 GNDA.n190 0.0217373
R4221 GNDA.n1837 GNDA.n193 0.0217373
R4222 GNDA.n1840 GNDA.n1839 0.0217373
R4223 GNDA.n192 GNDA.n189 0.0217373
R4224 GNDA.n192 GNDA.n190 0.0217373
R4225 GNDA.n1837 GNDA.n1836 0.0217373
R4226 GNDA.n1838 GNDA.n1835 0.0217373
R4227 GNDA.n1836 GNDA.n1822 0.0217373
R4228 GNDA.n1843 GNDA.n1842 0.0217373
R4229 GNDA.n1842 GNDA.n188 0.0217373
R4230 GNDA.n1535 GNDA.n237 0.00911526
R4231 GNDA.n1536 GNDA.n1535 0.00911526
R4232 GNDA.n231 GNDA.n228 0.00911526
R4233 GNDA.n232 GNDA.n231 0.00911526
R4234 GNDA.n1538 GNDA.n235 0.00911526
R4235 GNDA.n239 GNDA.n237 0.00911526
R4236 GNDA.n235 GNDA.n234 0.00911526
R4237 GNDA.n229 GNDA.n228 0.00911526
R4238 GNDA.n233 GNDA.n232 0.00911526
R4239 a_36200_n1130.n11 a_36200_n1130.t13 310.488
R4240 a_36200_n1130.n6 a_36200_n1130.t14 310.488
R4241 a_36200_n1130.n1 a_36200_n1130.t18 310.488
R4242 a_36200_n1130.n9 a_36200_n1130.n5 297.433
R4243 a_36200_n1130.n4 a_36200_n1130.n0 297.433
R4244 a_36200_n1130.n15 a_36200_n1130.n14 297.433
R4245 a_36200_n1130.n13 a_36200_n1130.t11 184.097
R4246 a_36200_n1130.n8 a_36200_n1130.t7 184.097
R4247 a_36200_n1130.n3 a_36200_n1130.t9 184.097
R4248 a_36200_n1130.n12 a_36200_n1130.n11 167.094
R4249 a_36200_n1130.n7 a_36200_n1130.n6 167.094
R4250 a_36200_n1130.n2 a_36200_n1130.n1 167.094
R4251 a_36200_n1130.n14 a_36200_n1130.n13 161.3
R4252 a_36200_n1130.n9 a_36200_n1130.n8 161.3
R4253 a_36200_n1130.n4 a_36200_n1130.n3 161.3
R4254 a_36200_n1130.n11 a_36200_n1130.t16 120.501
R4255 a_36200_n1130.n12 a_36200_n1130.t3 120.501
R4256 a_36200_n1130.n6 a_36200_n1130.t17 120.501
R4257 a_36200_n1130.n7 a_36200_n1130.t1 120.501
R4258 a_36200_n1130.n1 a_36200_n1130.t15 120.501
R4259 a_36200_n1130.n2 a_36200_n1130.t5 120.501
R4260 a_36200_n1130.n14 a_36200_n1130.t0 50.2014
R4261 a_36200_n1130.n13 a_36200_n1130.n12 40.7027
R4262 a_36200_n1130.n8 a_36200_n1130.n7 40.7027
R4263 a_36200_n1130.n3 a_36200_n1130.n2 40.7027
R4264 a_36200_n1130.n5 a_36200_n1130.t8 39.4005
R4265 a_36200_n1130.n5 a_36200_n1130.t2 39.4005
R4266 a_36200_n1130.n0 a_36200_n1130.t10 39.4005
R4267 a_36200_n1130.n0 a_36200_n1130.t6 39.4005
R4268 a_36200_n1130.t12 a_36200_n1130.n15 39.4005
R4269 a_36200_n1130.n15 a_36200_n1130.t4 39.4005
R4270 a_36200_n1130.n10 a_36200_n1130.n9 6.6255
R4271 a_36200_n1130.n10 a_36200_n1130.n4 6.6255
R4272 a_36200_n1130.n14 a_36200_n1130.n10 4.5005
R4273 1st_Vout_2.n5 1st_Vout_2.t27 362.341
R4274 1st_Vout_2 1st_Vout_2.t21 354.812
R4275 1st_Vout_2.n7 1st_Vout_2.n6 302.183
R4276 1st_Vout_2 1st_Vout_2.n15 302.183
R4277 1st_Vout_2.n11 1st_Vout_2.n10 297.683
R4278 1st_Vout_2.n13 1st_Vout_2.t28 194.809
R4279 1st_Vout_2.n13 1st_Vout_2.t24 194.809
R4280 1st_Vout_2.n8 1st_Vout_2.t32 194.809
R4281 1st_Vout_2.n8 1st_Vout_2.t19 194.809
R4282 1st_Vout_2.n14 1st_Vout_2.n13 166.03
R4283 1st_Vout_2.n9 1st_Vout_2.n8 166.03
R4284 1st_Vout_2.n11 1st_Vout_2.t0 49.5035
R4285 1st_Vout_2.n15 1st_Vout_2.t2 39.4005
R4286 1st_Vout_2.n15 1st_Vout_2.t5 39.4005
R4287 1st_Vout_2.n6 1st_Vout_2.t4 39.4005
R4288 1st_Vout_2.n6 1st_Vout_2.t1 39.4005
R4289 1st_Vout_2.n10 1st_Vout_2.t3 39.4005
R4290 1st_Vout_2.n10 1st_Vout_2.t6 39.4005
R4291 1st_Vout_2.n5 1st_Vout_2.n4 33.8685
R4292 1st_Vout_2.n0 1st_Vout_2.t22 4.8295
R4293 1st_Vout_2.n0 1st_Vout_2.t31 4.8295
R4294 1st_Vout_2.n2 1st_Vout_2.t13 4.8295
R4295 1st_Vout_2.n1 1st_Vout_2.t26 4.8295
R4296 1st_Vout_2.n2 1st_Vout_2.t18 4.8295
R4297 1st_Vout_2.n2 1st_Vout_2.t29 4.8295
R4298 1st_Vout_2.n3 1st_Vout_2.t11 4.8295
R4299 1st_Vout_2.n3 1st_Vout_2.t25 4.8295
R4300 1st_Vout_2.n3 1st_Vout_2.t23 4.8295
R4301 1st_Vout_2.n0 1st_Vout_2.t20 4.5005
R4302 1st_Vout_2.n0 1st_Vout_2.t17 4.5005
R4303 1st_Vout_2.n2 1st_Vout_2.t12 4.5005
R4304 1st_Vout_2.n1 1st_Vout_2.t10 4.5005
R4305 1st_Vout_2.n2 1st_Vout_2.t16 4.5005
R4306 1st_Vout_2.n2 1st_Vout_2.t15 4.5005
R4307 1st_Vout_2.n3 1st_Vout_2.t8 4.5005
R4308 1st_Vout_2.n3 1st_Vout_2.t7 4.5005
R4309 1st_Vout_2.n3 1st_Vout_2.t14 4.5005
R4310 1st_Vout_2.n4 1st_Vout_2.t30 4.5005
R4311 1st_Vout_2.n4 1st_Vout_2.t9 4.5005
R4312 1st_Vout_2.n12 1st_Vout_2.n11 4.5005
R4313 1st_Vout_2.n7 1st_Vout_2.n5 2.90725
R4314 1st_Vout_2 1st_Vout_2.n14 1.03175
R4315 1st_Vout_2.n3 1st_Vout_2.n2 0.8935
R4316 1st_Vout_2.n2 1st_Vout_2.n0 0.8935
R4317 1st_Vout_2.n12 1st_Vout_2.n9 0.7505
R4318 1st_Vout_2.n4 1st_Vout_2.n3 0.6585
R4319 1st_Vout_2.n2 1st_Vout_2.n1 0.6585
R4320 1st_Vout_2.n9 1st_Vout_2.n7 0.3755
R4321 1st_Vout_2.n14 1st_Vout_2.n12 0.3755
R4322 V_mir1.n11 V_mir1.t14 310.488
R4323 V_mir1.n6 V_mir1.t15 310.488
R4324 V_mir1.n1 V_mir1.t16 310.488
R4325 V_mir1.n9 V_mir1.n5 297.433
R4326 V_mir1.n4 V_mir1.n0 297.433
R4327 V_mir1.n15 V_mir1.n14 297.433
R4328 V_mir1.n13 V_mir1.t3 184.097
R4329 V_mir1.n8 V_mir1.t5 184.097
R4330 V_mir1.n3 V_mir1.t1 184.097
R4331 V_mir1.n12 V_mir1.n11 167.094
R4332 V_mir1.n7 V_mir1.n6 167.094
R4333 V_mir1.n2 V_mir1.n1 167.094
R4334 V_mir1.n14 V_mir1.n13 161.3
R4335 V_mir1.n9 V_mir1.n8 161.3
R4336 V_mir1.n4 V_mir1.n3 161.3
R4337 V_mir1.n11 V_mir1.t17 120.501
R4338 V_mir1.n12 V_mir1.t11 120.501
R4339 V_mir1.n6 V_mir1.t18 120.501
R4340 V_mir1.n7 V_mir1.t7 120.501
R4341 V_mir1.n1 V_mir1.t13 120.501
R4342 V_mir1.n2 V_mir1.t9 120.501
R4343 V_mir1.n9 V_mir1.t0 50.2014
R4344 V_mir1.n13 V_mir1.n12 40.7027
R4345 V_mir1.n8 V_mir1.n7 40.7027
R4346 V_mir1.n3 V_mir1.n2 40.7027
R4347 V_mir1.n5 V_mir1.t8 39.4005
R4348 V_mir1.n5 V_mir1.t6 39.4005
R4349 V_mir1.n0 V_mir1.t10 39.4005
R4350 V_mir1.n0 V_mir1.t2 39.4005
R4351 V_mir1.t12 V_mir1.n15 39.4005
R4352 V_mir1.n15 V_mir1.t4 39.4005
R4353 V_mir1.n10 V_mir1.n4 6.6255
R4354 V_mir1.n14 V_mir1.n10 6.6255
R4355 V_mir1.n10 V_mir1.n9 4.5005
R4356 cap_res2 cap_res2.t0 118.561
R4357 cap_res2 cap_res2.t13 0.206125
R4358 cap_res2.t2 cap_res2.t18 0.1603
R4359 cap_res2.t20 cap_res2.t5 0.1603
R4360 cap_res2.t12 cap_res2.t3 0.1603
R4361 cap_res2.t17 cap_res2.t4 0.1603
R4362 cap_res2.t10 cap_res2.t1 0.1603
R4363 cap_res2.n1 cap_res2.t8 0.159278
R4364 cap_res2.n2 cap_res2.t15 0.159278
R4365 cap_res2.n3 cap_res2.t11 0.159278
R4366 cap_res2.n4 cap_res2.t19 0.159278
R4367 cap_res2.n4 cap_res2.t2 0.1368
R4368 cap_res2.n4 cap_res2.t6 0.1368
R4369 cap_res2.n3 cap_res2.t20 0.1368
R4370 cap_res2.n3 cap_res2.t16 0.1368
R4371 cap_res2.n2 cap_res2.t12 0.1368
R4372 cap_res2.n2 cap_res2.t9 0.1368
R4373 cap_res2.n1 cap_res2.t17 0.1368
R4374 cap_res2.n1 cap_res2.t14 0.1368
R4375 cap_res2.n0 cap_res2.t10 0.1368
R4376 cap_res2.n0 cap_res2.t7 0.1368
R4377 cap_res2.t8 cap_res2.n0 0.00152174
R4378 cap_res2.t15 cap_res2.n1 0.00152174
R4379 cap_res2.t11 cap_res2.n2 0.00152174
R4380 cap_res2.t19 cap_res2.n3 0.00152174
R4381 cap_res2.t13 cap_res2.n4 0.00152174
R4382 Vin-.n7 Vin-.t8 539.797
R4383 Vin-.n6 Vin-.n5 314.526
R4384 Vin-.n8 Vin-.t0 117.817
R4385 Vin-.n4 Vin-.n2 107.079
R4386 Vin-.n4 Vin-.n3 104.829
R4387 Vin-.n1 Vin-.n0 83.5719
R4388 Vin-.n13 Vin-.n1 73.682
R4389 Vin-.n5 Vin-.t1 39.4005
R4390 Vin-.n5 Vin-.t2 39.4005
R4391 Vin-.n10 Vin-.t3 36.6632
R4392 Vin-.t3 Vin-.n1 25.7843
R4393 Vin-.n9 Vin-.n8 24.3755
R4394 Vin-.n8 Vin-.n7 14.0317
R4395 Vin-.n3 Vin-.t7 13.1338
R4396 Vin-.n3 Vin-.t4 13.1338
R4397 Vin-.n2 Vin-.t5 13.1338
R4398 Vin-.n2 Vin-.t6 13.1338
R4399 Vin-.n7 Vin-.n6 10.1567
R4400 Vin-.n6 Vin-.n4 2.0005
R4401 Vin-.n11 Vin-.n10 1.80777
R4402 Vin-.n12 Vin-.n11 1.5505
R4403 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter Vin-.n13 1.07742
R4404 Vin-.n10 Vin-.n9 1.04793
R4405 Vin-.n13 Vin-.n12 0.763532
R4406 Vin-.n11 Vin-.n0 0.590702
R4407 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter Vin-.n0 0.498483
R4408 Vin-.n12 Vin-.n9 0.0106786
R4409 START_UP.n2 START_UP.t6 238.322
R4410 START_UP.n2 START_UP.t7 238.322
R4411 START_UP.n3 START_UP.n2 167.332
R4412 START_UP.n1 START_UP.t1 130.001
R4413 START_UP.n4 START_UP.n0 108.546
R4414 START_UP.n5 START_UP.n4 105.171
R4415 START_UP.n1 START_UP.t0 81.7084
R4416 START_UP.n3 START_UP.n1 50.9489
R4417 START_UP.n0 START_UP.t2 13.1338
R4418 START_UP.n0 START_UP.t3 13.1338
R4419 START_UP.n5 START_UP.t4 13.1338
R4420 START_UP.t5 START_UP.n5 13.1338
R4421 START_UP.n4 START_UP.n3 2.17238
R4422 V1.n5 V1.t7 537.609
R4423 V1.t0 V1.n5 115.737
R4424 V1.n2 V1.n0 107.266
R4425 V1.n2 V1.n1 105.016
R4426 V1.n4 V1.n3 105.016
R4427 V1.n0 V1.t5 13.1338
R4428 V1.n0 V1.t2 13.1338
R4429 V1.n1 V1.t3 13.1338
R4430 V1.n1 V1.t4 13.1338
R4431 V1.n3 V1.t1 13.1338
R4432 V1.n3 V1.t6 13.1338
R4433 V1.n5 V1.n4 8.7505
R4434 V1.n4 V1.n2 2.2505
R4435 a_38370_n6700.t0 a_38370_n6700.t1 178.133
R4436 a_38490_n7778.t0 a_38490_n7778.t1 178.133
R4437 V_p_2.n0 V_p_2.t1 142.327
R4438 V_p_2.t0 V_p_2.n0 9.6005
R4439 V_p_2.n0 V_p_2.t2 9.6005
R4440 a_38040_n7928.t0 a_38040_n7928.t1 178.133
R4441 V_p_1.n0 V_p_1.t1 99.603
R4442 V_p_1.n0 V_p_1.t2 9.6005
R4443 V_p_1.t0 V_p_1.n0 9.6005
R4444 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 172.969
R4445 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 83.5719
R4446 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 83.5719
R4447 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 83.5719
R4448 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 83.5719
R4449 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R4450 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 83.5719
R4451 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 83.5719
R4452 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R4453 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 83.5719
R4454 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R4455 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 83.5719
R4456 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 83.5719
R4457 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R4458 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 83.5719
R4459 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 83.5719
R4460 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 83.5719
R4461 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 83.5719
R4462 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R4463 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R4464 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R4465 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.682
R4466 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.682
R4467 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 73.3165
R4468 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 73.3165
R4469 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 73.3165
R4470 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 73.3165
R4471 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 73.3165
R4472 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.3165
R4473 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 73.19
R4474 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 73.19
R4475 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 73.19
R4476 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 73.19
R4477 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 73.19
R4478 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.19
R4479 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 36.6632
R4480 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 36.6632
R4481 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 26.074
R4482 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 26.074
R4483 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 26.074
R4484 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 26.074
R4485 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 26.074
R4486 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 26.074
R4487 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 25.7843
R4488 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R4489 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 25.7843
R4490 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 25.7843
R4491 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 25.7843
R4492 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R4493 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R4494 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 25.7843
R4495 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4496 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4497 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4498 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 9.3005
R4499 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4500 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4501 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4502 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 9.3005
R4503 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4504 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4505 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4506 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 9.3005
R4507 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4508 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4509 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4510 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R4511 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4512 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4513 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4514 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R4515 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 9.3005
R4516 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4517 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4518 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4519 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R4520 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R4521 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4522 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4523 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4524 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 9.3005
R4525 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R4526 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4527 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4528 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4529 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R4530 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 9.3005
R4531 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4532 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4533 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4534 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 9.3005
R4535 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4536 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4537 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4538 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R4539 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4540 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4541 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4542 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R4543 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 9.3005
R4544 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4545 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4546 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4547 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R4548 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 9.3005
R4549 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 4.64654
R4550 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 4.64654
R4551 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 4.64654
R4552 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 4.64654
R4553 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R4554 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 4.64654
R4555 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 4.64654
R4556 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 4.64654
R4557 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 4.64654
R4558 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 2.36206
R4559 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 2.36206
R4560 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 2.36206
R4561 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.36206
R4562 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 2.19742
R4563 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 2.19742
R4564 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 2.19742
R4565 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 2.19742
R4566 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.80777
R4567 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.80777
R4568 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.5505
R4569 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R4570 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R4571 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.5505
R4572 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 1.5505
R4573 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R4574 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 1.5505
R4575 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 1.5505
R4576 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.5505
R4577 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 1.5505
R4578 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 1.5505
R4579 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.5505
R4580 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 1.5505
R4581 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 1.5505
R4582 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 1.5505
R4583 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.5505
R4584 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 1.5505
R4585 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 1.5505
R4586 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 1.19225
R4587 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 1.19225
R4588 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.19225
R4589 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 1.19225
R4590 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 1.19225
R4591 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 1.19225
R4592 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 1.07742
R4593 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 1.07742
R4594 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R4595 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 1.07024
R4596 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 1.07024
R4597 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 1.07024
R4598 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R4599 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R4600 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.04793
R4601 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.04793
R4602 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.0237
R4603 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 1.0237
R4604 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 1.0237
R4605 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 1.0237
R4606 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.0237
R4607 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.0237
R4608 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 0.959578
R4609 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 0.959578
R4610 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.959578
R4611 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.959578
R4612 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.959578
R4613 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 0.959578
R4614 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.885803
R4615 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.885803
R4616 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.885803
R4617 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.885803
R4618 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 0.885803
R4619 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R4620 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 0.812055
R4621 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 0.812055
R4622 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.77514
R4623 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 0.77514
R4624 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.77514
R4625 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.77514
R4626 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.77514
R4627 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R4628 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.763532
R4629 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.763532
R4630 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.756696
R4631 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4632 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4633 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.756696
R4634 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4635 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 0.756696
R4636 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.647417
R4637 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.647417
R4638 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.590702
R4639 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.590702
R4640 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.590702
R4641 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 0.590702
R4642 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.590702
R4643 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R4644 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 0.590702
R4645 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.590702
R4646 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4647 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4648 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 0.498483
R4649 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.498483
R4650 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4651 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4652 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4653 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.498483
R4654 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.290206
R4655 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 0.290206
R4656 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R4657 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.290206
R4658 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.290206
R4659 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.290206
R4660 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.154071
R4661 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 0.154071
R4662 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.154071
R4663 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 0.154071
R4664 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.137464
R4665 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 0.137464
R4666 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.134964
R4667 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 0.134964
R4668 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R4669 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.0183571
R4670 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R4671 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R4672 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 0.0183571
R4673 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R4674 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R4675 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.0183571
R4676 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.0183571
R4677 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.0183571
R4678 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.0183571
R4679 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.0183571
R4680 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.0183571
R4681 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 0.0183571
R4682 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.0183571
R4683 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.0183571
R4684 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 0.0183571
R4685 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.0183571
R4686 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0106786
R4687 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 0.0106786
R4688 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 0.0106786
R4689 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 0.0106786
R4690 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.0106786
R4691 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R4692 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.00992001
R4693 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00992001
R4694 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 0.00992001
R4695 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.00992001
R4696 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R4697 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 0.00992001
R4698 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 0.00992001
R4699 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00992001
R4700 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 0.00992001
R4701 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R4702 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R4703 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.00992001
R4704 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.00992001
R4705 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.00992001
R4706 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.00992001
R4707 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.00992001
R4708 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.00992001
R4709 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R4710 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00817857
R4711 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.00817857
R4712 a_32970_n7928.t0 a_32970_n7928.t1 178.133
R4713 a_33090_n6320.t0 a_33090_n6320.t1 178.133
R4714 a_37920_n6320.t0 a_37920_n6320.t1 178.133
C0 1st_Vout_2 V_CUR_REF_REG 1.06368f
C1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter Vin+ 1.06291f
C2 V_TOP cap_res1 0.607363f
C3 CURRENT_OUTPUT V_CUR_REF_REG 0.01137f
C4 V_CUR_REF_REG sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.793278f
C5 cap_res2 1st_Vout_2 7.29943f
C6 1st_Vout_2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.4193f
C7 VDDA Vin+ 1.80314f
C8 VDDA V_CUR_REF_REG 3.96867f
C9 V_TOP Vin+ 2.13673f
C10 VDDA 1st_Vout_2 1.34874f
C11 VDDA CURRENT_OUTPUT 3.5212f
C12 V_CUR_REF_REG V_TOP 0.756389f
C13 VDDA cap_res2 0.531875f
C14 VDDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.036669f
C15 1st_Vout_2 V_TOP 0.074293f
C16 CURRENT_OUTPUT V_TOP 0.019757f
C17 cap_res2 V_TOP 0.01893f
C18 V_TOP sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.025706f
C19 V_CUR_REF_REG Vin+ 1.57773f
C20 VDDA V_TOP 16.5127f
C21 1st_Vout_2 Vin+ 0.317284f
C22 VDDA cap_res1 1.26357f
C23 CURRENT_OUTPUT GNDA 1.25602f
C24 VDDA GNDA 46.483517f
C25 cap_res2 GNDA 6.728005f
C26 cap_res1 GNDA 6.013068f
C27 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 16.8331f
C28 1st_Vout_2 GNDA 7.427619f
C29 Vin+ GNDA 4.339304f
C30 V_TOP GNDA 10.622867f
C31 V_CUR_REF_REG GNDA 5.067328f
C32 V1.t5 GNDA 0.035662f
C33 V1.t2 GNDA 0.035662f
C34 V1.n0 GNDA 0.099479f
C35 V1.t3 GNDA 0.035662f
C36 V1.t4 GNDA 0.035662f
C37 V1.n1 GNDA 0.089537f
C38 V1.n2 GNDA 1.09957f
C39 V1.t1 GNDA 0.035662f
C40 V1.t6 GNDA 0.035662f
C41 V1.n3 GNDA 0.089537f
C42 V1.n4 GNDA 0.826974f
C43 V1.t7 GNDA 0.058965f
C44 V1.n5 GNDA 1.8495f
C45 V1.t0 GNDA 0.172471f
C46 START_UP.t4 GNDA 0.058627f
C47 START_UP.t2 GNDA 0.058627f
C48 START_UP.t3 GNDA 0.058627f
C49 START_UP.n0 GNDA 0.170978f
C50 START_UP.t0 GNDA 2.33703f
C51 START_UP.t1 GNDA 0.061434f
C52 START_UP.n1 GNDA 1.7713f
C53 START_UP.t7 GNDA 0.022031f
C54 START_UP.t6 GNDA 0.022031f
C55 START_UP.n2 GNDA 0.063205f
C56 START_UP.n3 GNDA 1.43522f
C57 START_UP.n4 GNDA 1.93784f
C58 START_UP.n5 GNDA 0.14442f
C59 START_UP.t5 GNDA 0.058627f
C60 Vin-.n0 GNDA 0.056136f
C61 Vin-.n1 GNDA 0.383665f
C62 Vin-.t5 GNDA 0.032904f
C63 Vin-.t6 GNDA 0.032904f
C64 Vin-.n2 GNDA 0.088024f
C65 Vin-.t7 GNDA 0.032904f
C66 Vin-.t4 GNDA 0.032904f
C67 Vin-.n3 GNDA 0.079838f
C68 Vin-.n4 GNDA 0.9026f
C69 Vin-.t1 GNDA 0.010968f
C70 Vin-.t2 GNDA 0.010968f
C71 Vin-.n5 GNDA 0.030918f
C72 Vin-.n6 GNDA 0.636189f
C73 Vin-.t8 GNDA 0.053296f
C74 Vin-.n7 GNDA 0.598388f
C75 Vin-.t0 GNDA 0.138906f
C76 Vin-.n8 GNDA 0.734816f
C77 Vin-.n9 GNDA 1.7887f
C78 Vin-.t3 GNDA 0.399528f
C79 Vin-.n10 GNDA 0.357045f
C80 Vin-.n11 GNDA 0.148745f
C81 Vin-.n12 GNDA 0.702909f
C82 Vin-.n13 GNDA 0.44709f
C83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.09965f
C84 cap_res2.t6 GNDA 0.315239f
C85 cap_res2.t18 GNDA 0.331845f
C86 cap_res2.t2 GNDA 0.333048f
C87 cap_res2.t16 GNDA 0.315239f
C88 cap_res2.t5 GNDA 0.331845f
C89 cap_res2.t20 GNDA 0.333048f
C90 cap_res2.t9 GNDA 0.315239f
C91 cap_res2.t3 GNDA 0.331845f
C92 cap_res2.t12 GNDA 0.333048f
C93 cap_res2.t14 GNDA 0.315239f
C94 cap_res2.t4 GNDA 0.331845f
C95 cap_res2.t17 GNDA 0.333048f
C96 cap_res2.t7 GNDA 0.315239f
C97 cap_res2.t1 GNDA 0.331845f
C98 cap_res2.t10 GNDA 0.333048f
C99 cap_res2.n0 GNDA 0.222436f
C100 cap_res2.t8 GNDA 0.177138f
C101 cap_res2.n1 GNDA 0.241348f
C102 cap_res2.t15 GNDA 0.177138f
C103 cap_res2.n2 GNDA 0.241348f
C104 cap_res2.t11 GNDA 0.177138f
C105 cap_res2.n3 GNDA 0.241348f
C106 cap_res2.t19 GNDA 0.177138f
C107 cap_res2.n4 GNDA 0.241348f
C108 cap_res2.t13 GNDA 0.167759f
C109 cap_res2.t0 GNDA 0.083968f
C110 1st_Vout_2.n0 GNDA 0.302322f
C111 1st_Vout_2.n1 GNDA 0.132617f
C112 1st_Vout_2.n2 GNDA 0.546201f
C113 1st_Vout_2.n3 GNDA 0.509114f
C114 1st_Vout_2.n4 GNDA 0.544617f
C115 1st_Vout_2.t22 GNDA 0.201167f
C116 1st_Vout_2.t20 GNDA 0.197798f
C117 1st_Vout_2.t31 GNDA 0.201167f
C118 1st_Vout_2.t17 GNDA 0.197798f
C119 1st_Vout_2.t13 GNDA 0.201167f
C120 1st_Vout_2.t12 GNDA 0.197798f
C121 1st_Vout_2.t26 GNDA 0.201167f
C122 1st_Vout_2.t10 GNDA 0.197798f
C123 1st_Vout_2.t18 GNDA 0.201167f
C124 1st_Vout_2.t16 GNDA 0.197798f
C125 1st_Vout_2.t29 GNDA 0.201167f
C126 1st_Vout_2.t15 GNDA 0.197798f
C127 1st_Vout_2.t11 GNDA 0.201167f
C128 1st_Vout_2.t8 GNDA 0.197798f
C129 1st_Vout_2.t25 GNDA 0.201167f
C130 1st_Vout_2.t7 GNDA 0.197798f
C131 1st_Vout_2.t23 GNDA 0.201167f
C132 1st_Vout_2.t14 GNDA 0.197798f
C133 1st_Vout_2.t30 GNDA 0.197798f
C134 1st_Vout_2.t9 GNDA 0.197798f
C135 1st_Vout_2.t27 GNDA 0.01171f
C136 1st_Vout_2.n5 GNDA 0.57223f
C137 1st_Vout_2.n6 GNDA 0.010843f
C138 1st_Vout_2.n7 GNDA 0.103269f
C139 1st_Vout_2.n8 GNDA 0.014831f
C140 1st_Vout_2.n9 GNDA 0.057383f
C141 1st_Vout_2.n10 GNDA 0.010155f
C142 1st_Vout_2.t0 GNDA 0.045272f
C143 1st_Vout_2.n11 GNDA 0.144597f
C144 1st_Vout_2.n12 GNDA 0.035604f
C145 1st_Vout_2.n13 GNDA 0.014831f
C146 1st_Vout_2.n14 GNDA 0.057383f
C147 1st_Vout_2.n15 GNDA 0.010843f
C148 1st_Vout_2.t21 GNDA 0.011835f
C149 Vin+.t6 GNDA 0.080172f
C150 Vin+.t4 GNDA 0.050158f
C151 Vin+.t5 GNDA 0.050158f
C152 Vin+.n0 GNDA 0.124769f
C153 Vin+.t2 GNDA 0.050158f
C154 Vin+.t3 GNDA 0.050158f
C155 Vin+.n1 GNDA 0.119903f
C156 Vin+.n2 GNDA 1.73187f
C157 Vin+.t1 GNDA 0.336693f
C158 Vin+.t0 GNDA 0.14593f
C159 Vin+.n3 GNDA 2.14622f
C160 Vin+.n4 GNDA 0.876731f
C161 V_TOP.t16 GNDA 0.172467f
C162 V_TOP.n0 GNDA 0.022579f
C163 V_TOP.t39 GNDA 0.171428f
C164 V_TOP.t28 GNDA 0.173018f
C165 V_TOP.t36 GNDA 0.173764f
C166 V_TOP.n1 GNDA 0.218626f
C167 V_TOP.t41 GNDA 0.173764f
C168 V_TOP.n2 GNDA 0.119759f
C169 V_TOP.t48 GNDA 0.173764f
C170 V_TOP.n3 GNDA 0.119759f
C171 V_TOP.t15 GNDA 0.173764f
C172 V_TOP.n4 GNDA 0.119759f
C173 V_TOP.t26 GNDA 0.173764f
C174 V_TOP.n5 GNDA 0.119759f
C175 V_TOP.n6 GNDA 0.033868f
C176 V_TOP.t34 GNDA 0.172666f
C177 V_TOP.n7 GNDA 0.076954f
C178 V_TOP.t7 GNDA 0.173299f
C179 V_TOP.t47 GNDA 0.510295f
C180 V_TOP.t46 GNDA 0.501749f
C181 V_TOP.t25 GNDA 0.510295f
C182 V_TOP.t27 GNDA 0.501749f
C183 V_TOP.n8 GNDA 0.336406f
C184 V_TOP.n9 GNDA 0.430484f
C185 V_TOP.t35 GNDA 0.510295f
C186 V_TOP.t33 GNDA 0.501749f
C187 V_TOP.t19 GNDA 0.510295f
C188 V_TOP.t20 GNDA 0.501749f
C189 V_TOP.n10 GNDA 0.336406f
C190 V_TOP.n11 GNDA 0.524562f
C191 V_TOP.t44 GNDA 0.510295f
C192 V_TOP.t43 GNDA 0.501749f
C193 V_TOP.t23 GNDA 0.510295f
C194 V_TOP.t24 GNDA 0.501749f
C195 V_TOP.n12 GNDA 0.336406f
C196 V_TOP.n13 GNDA 0.524562f
C197 V_TOP.t32 GNDA 0.510295f
C198 V_TOP.t30 GNDA 0.501749f
C199 V_TOP.t17 GNDA 0.510295f
C200 V_TOP.t18 GNDA 0.501749f
C201 V_TOP.n14 GNDA 0.336406f
C202 V_TOP.n15 GNDA 0.524562f
C203 V_TOP.t40 GNDA 0.510295f
C204 V_TOP.t29 GNDA 0.501749f
C205 V_TOP.n16 GNDA 0.430484f
C206 V_TOP.t37 GNDA 0.501749f
C207 V_TOP.n17 GNDA 0.219515f
C208 V_TOP.t21 GNDA 0.501749f
C209 V_TOP.n18 GNDA 1.05142f
C210 V_TOP.t2 GNDA 0.141186f
C211 V_TOP.n19 GNDA 1.66799f
C212 V_TOP.t1 GNDA 0.012544f
C213 V_TOP.t4 GNDA 0.012544f
C214 V_TOP.n20 GNDA 0.025684f
C215 V_TOP.t3 GNDA 0.012544f
C216 V_TOP.t0 GNDA 0.012544f
C217 V_TOP.n21 GNDA 0.029192f
C218 V_TOP.n22 GNDA 0.344015f
C219 V_TOP.t10 GNDA 0.012544f
C220 V_TOP.t6 GNDA 0.012544f
C221 V_TOP.n23 GNDA 0.025684f
C222 V_TOP.n24 GNDA 0.212647f
C223 V_TOP.n25 GNDA 0.723899f
C224 V_TOP.t12 GNDA 0.012544f
C225 V_TOP.t8 GNDA 0.012544f
C226 V_TOP.n26 GNDA 0.027096f
C227 V_TOP.n27 GNDA 0.266427f
C228 V_TOP.t13 GNDA 0.012544f
C229 V_TOP.t9 GNDA 0.012544f
C230 V_TOP.n28 GNDA 0.027096f
C231 V_TOP.n29 GNDA 0.273954f
C232 V_TOP.t5 GNDA 0.012544f
C233 V_TOP.t11 GNDA 0.012544f
C234 V_TOP.n30 GNDA 0.027096f
C235 V_TOP.n31 GNDA 0.25537f
C236 V_TOP.n32 GNDA 0.505711f
C237 V_TOP.n33 GNDA 0.12042f
C238 V_TOP.n34 GNDA 0.070666f
C239 V_TOP.n35 GNDA 0.033868f
C240 V_TOP.t45 GNDA 0.172427f
C241 V_TOP.n36 GNDA 0.113569f
C242 V_TOP.t14 GNDA 0.173764f
C243 V_TOP.n37 GNDA 0.119759f
C244 V_TOP.t22 GNDA 0.173764f
C245 V_TOP.n38 GNDA 0.119759f
C246 V_TOP.t31 GNDA 0.173764f
C247 V_TOP.n39 GNDA 0.119759f
C248 V_TOP.t38 GNDA 0.173764f
C249 V_TOP.n40 GNDA 0.119759f
C250 V_TOP.t42 GNDA 0.173764f
C251 V_TOP.n41 GNDA 0.119759f
C252 V_TOP.t49 GNDA 0.173764f
C253 V_TOP.n42 GNDA 0.10847f
C254 CURRENT_OUTPUT.t9 GNDA 0.02211f
C255 CURRENT_OUTPUT.t2 GNDA 0.02211f
C256 CURRENT_OUTPUT.n0 GNDA 0.045394f
C257 CURRENT_OUTPUT.t0 GNDA 0.02211f
C258 CURRENT_OUTPUT.t3 GNDA 0.02211f
C259 CURRENT_OUTPUT.n1 GNDA 0.051982f
C260 CURRENT_OUTPUT.t8 GNDA 0.02211f
C261 CURRENT_OUTPUT.t5 GNDA 0.02211f
C262 CURRENT_OUTPUT.n2 GNDA 0.051451f
C263 CURRENT_OUTPUT.n3 GNDA 0.964476f
C264 CURRENT_OUTPUT.t4 GNDA 0.02211f
C265 CURRENT_OUTPUT.t1 GNDA 0.02211f
C266 CURRENT_OUTPUT.n4 GNDA 0.045357f
C267 CURRENT_OUTPUT.n5 GNDA -0.865603f
C268 CURRENT_OUTPUT.n6 GNDA 1.2771f
C269 CURRENT_OUTPUT.t6 GNDA 0.02211f
C270 CURRENT_OUTPUT.t10 GNDA 0.02211f
C271 CURRENT_OUTPUT.n7 GNDA 0.051451f
C272 CURRENT_OUTPUT.n8 GNDA 0.559603f
C273 CURRENT_OUTPUT.t7 GNDA 0.02211f
C274 CURRENT_OUTPUT.t11 GNDA 0.02211f
C275 CURRENT_OUTPUT.n9 GNDA 0.051451f
C276 CURRENT_OUTPUT.n10 GNDA 0.49798f
C277 CURRENT_OUTPUT.n11 GNDA 0.097284f
C278 CURRENT_OUTPUT.n12 GNDA 0.296205f
C279 cap_res1.t16 GNDA 0.355848f
C280 cap_res1.t5 GNDA 0.357137f
C281 cap_res1.t6 GNDA 0.33804f
C282 cap_res1.t18 GNDA 0.355848f
C283 cap_res1.t19 GNDA 0.357137f
C284 cap_res1.t10 GNDA 0.33804f
C285 cap_res1.t13 GNDA 0.355848f
C286 cap_res1.t14 GNDA 0.357137f
C287 cap_res1.t4 GNDA 0.33804f
C288 cap_res1.t15 GNDA 0.355848f
C289 cap_res1.t17 GNDA 0.357137f
C290 cap_res1.t8 GNDA 0.33804f
C291 cap_res1.t11 GNDA 0.355848f
C292 cap_res1.t12 GNDA 0.357137f
C293 cap_res1.t2 GNDA 0.33804f
C294 cap_res1.n0 GNDA 0.238525f
C295 cap_res1.t1 GNDA 0.18995f
C296 cap_res1.n1 GNDA 0.258805f
C297 cap_res1.t7 GNDA 0.18995f
C298 cap_res1.n2 GNDA 0.258805f
C299 cap_res1.t3 GNDA 0.18995f
C300 cap_res1.n3 GNDA 0.258805f
C301 cap_res1.t9 GNDA 0.18995f
C302 cap_res1.n4 GNDA 0.258805f
C303 cap_res1.t20 GNDA 0.201666f
C304 cap_res1.t0 GNDA 0.081828f
C305 1st_Vout_1.n0 GNDA 2.83353f
C306 1st_Vout_1.n1 GNDA 0.431786f
C307 1st_Vout_1.n2 GNDA 0.969511f
C308 1st_Vout_1.n3 GNDA 3.5912f
C309 1st_Vout_1.n4 GNDA 0.703222f
C310 1st_Vout_1.t17 GNDA 0.01671f
C311 1st_Vout_1.n5 GNDA 0.014961f
C312 1st_Vout_1.t8 GNDA 0.010934f
C313 1st_Vout_1.t21 GNDA 0.010934f
C314 1st_Vout_1.n6 GNDA 0.020826f
C315 1st_Vout_1.t12 GNDA 0.282502f
C316 1st_Vout_1.t20 GNDA 0.287314f
C317 1st_Vout_1.t18 GNDA 0.282502f
C318 1st_Vout_1.t32 GNDA 0.282502f
C319 1st_Vout_1.t31 GNDA 0.287314f
C320 1st_Vout_1.t13 GNDA 0.287314f
C321 1st_Vout_1.t11 GNDA 0.282502f
C322 1st_Vout_1.t25 GNDA 0.282502f
C323 1st_Vout_1.t24 GNDA 0.287314f
C324 1st_Vout_1.t16 GNDA 0.287314f
C325 1st_Vout_1.t15 GNDA 0.282502f
C326 1st_Vout_1.t30 GNDA 0.282502f
C327 1st_Vout_1.t29 GNDA 0.287314f
C328 1st_Vout_1.t10 GNDA 0.287314f
C329 1st_Vout_1.t9 GNDA 0.282502f
C330 1st_Vout_1.t23 GNDA 0.282502f
C331 1st_Vout_1.t22 GNDA 0.287314f
C332 1st_Vout_1.t26 GNDA 0.287314f
C333 1st_Vout_1.t7 GNDA 0.282502f
C334 1st_Vout_1.t27 GNDA 0.282502f
C335 1st_Vout_1.t19 GNDA 0.016978f
C336 1st_Vout_1.n7 GNDA 0.014961f
C337 1st_Vout_1.t14 GNDA 0.010934f
C338 1st_Vout_1.t28 GNDA 0.010934f
C339 1st_Vout_1.n8 GNDA 0.020826f
C340 1st_Vout_1.n9 GNDA 0.014533f
C341 1st_Vout_1.n10 GNDA 0.207089f
C342 1st_Vout_1.t6 GNDA 0.064412f
C343 V_CUR_REF_REG.n0 GNDA 0.018468f
C344 V_CUR_REF_REG.n1 GNDA 0.018353f
C345 V_CUR_REF_REG.n2 GNDA 0.213743f
C346 V_CUR_REF_REG.n3 GNDA 0.018353f
C347 V_CUR_REF_REG.n4 GNDA 0.112795f
C348 V_CUR_REF_REG.n5 GNDA 0.018353f
C349 V_CUR_REF_REG.n6 GNDA 0.112795f
C350 V_CUR_REF_REG.n7 GNDA 0.018353f
C351 V_CUR_REF_REG.n8 GNDA 0.112795f
C352 V_CUR_REF_REG.n9 GNDA 0.018353f
C353 V_CUR_REF_REG.n10 GNDA 0.455835f
C354 V_CUR_REF_REG.t0 GNDA 0.278272f
C355 V_CUR_REF_REG.n11 GNDA 2.15625f
C356 V_CUR_REF_REG.t13 GNDA 0.042841f
C357 VDDA.n1 GNDA 0.038807f
C358 VDDA.n2 GNDA 0.038807f
C359 VDDA.n4 GNDA 0.038807f
C360 VDDA.n5 GNDA 0.038807f
C361 VDDA.n7 GNDA 0.038807f
C362 VDDA.n8 GNDA 0.038807f
C363 VDDA.n9 GNDA 0.014329f
C364 VDDA.n10 GNDA 0.078542f
C365 VDDA.t117 GNDA 0.0135f
C366 VDDA.n11 GNDA 0.02599f
C367 VDDA.t119 GNDA 0.023074f
C368 VDDA.n13 GNDA 0.02599f
C369 VDDA.t116 GNDA 0.023074f
C370 VDDA.t114 GNDA 0.0135f
C371 VDDA.n14 GNDA 0.014329f
C372 VDDA.n15 GNDA 0.078542f
C373 VDDA.t99 GNDA 0.0135f
C374 VDDA.n16 GNDA 0.02599f
C375 VDDA.t101 GNDA 0.023074f
C376 VDDA.n18 GNDA 0.02599f
C377 VDDA.t110 GNDA 0.023074f
C378 VDDA.t108 GNDA 0.0135f
C379 VDDA.n19 GNDA 0.014329f
C380 VDDA.n20 GNDA 0.078542f
C381 VDDA.n21 GNDA 0.014329f
C382 VDDA.n22 GNDA 0.078542f
C383 VDDA.n23 GNDA 0.014329f
C384 VDDA.n24 GNDA 0.078542f
C385 VDDA.n25 GNDA 0.014329f
C386 VDDA.n26 GNDA 0.097031f
C387 VDDA.n27 GNDA 0.032894f
C388 VDDA.n28 GNDA 0.043682f
C389 VDDA.n29 GNDA 0.025597f
C390 VDDA.n30 GNDA 0.065794f
C391 VDDA.t109 GNDA 0.080177f
C392 VDDA.t162 GNDA 0.051079f
C393 VDDA.t190 GNDA 0.051079f
C394 VDDA.t168 GNDA 0.051079f
C395 VDDA.t184 GNDA 0.051079f
C396 VDDA.t198 GNDA 0.051079f
C397 VDDA.t178 GNDA 0.051079f
C398 VDDA.t194 GNDA 0.051079f
C399 VDDA.t172 GNDA 0.051079f
C400 VDDA.t186 GNDA 0.051079f
C401 VDDA.t166 GNDA 0.051079f
C402 VDDA.t100 GNDA 0.065489f
C403 VDDA.n31 GNDA 0.080481f
C404 VDDA.n32 GNDA 0.025597f
C405 VDDA.n33 GNDA 0.043682f
C406 VDDA.n34 GNDA 0.031481f
C407 VDDA.n35 GNDA 0.053069f
C408 VDDA.n36 GNDA 0.014329f
C409 VDDA.n37 GNDA 0.078542f
C410 VDDA.n38 GNDA 0.014329f
C411 VDDA.n39 GNDA 0.078542f
C412 VDDA.n40 GNDA 0.014329f
C413 VDDA.n41 GNDA 0.078542f
C414 VDDA.n42 GNDA 0.014329f
C415 VDDA.n43 GNDA 0.078542f
C416 VDDA.n44 GNDA 0.053069f
C417 VDDA.n45 GNDA 0.031481f
C418 VDDA.n46 GNDA 0.043682f
C419 VDDA.n47 GNDA 0.025597f
C420 VDDA.n48 GNDA 0.065794f
C421 VDDA.t115 GNDA 0.080177f
C422 VDDA.t164 GNDA 0.051079f
C423 VDDA.t182 GNDA 0.051079f
C424 VDDA.t174 GNDA 0.051079f
C425 VDDA.t188 GNDA 0.051079f
C426 VDDA.t160 GNDA 0.051079f
C427 VDDA.t180 GNDA 0.051079f
C428 VDDA.t196 GNDA 0.051079f
C429 VDDA.t176 GNDA 0.051079f
C430 VDDA.t192 GNDA 0.051079f
C431 VDDA.t170 GNDA 0.051079f
C432 VDDA.t118 GNDA 0.065489f
C433 VDDA.n49 GNDA 0.080481f
C434 VDDA.n50 GNDA 0.025597f
C435 VDDA.n51 GNDA 0.043682f
C436 VDDA.n52 GNDA 0.031481f
C437 VDDA.n53 GNDA 0.247053f
C438 VDDA.t42 GNDA 0.019901f
C439 VDDA.t152 GNDA 0.019901f
C440 VDDA.n54 GNDA 0.077433f
C441 VDDA.n55 GNDA 0.266192f
C442 VDDA.n56 GNDA 0.01871f
C443 VDDA.n58 GNDA 0.013267f
C444 VDDA.n61 GNDA 0.013267f
C445 VDDA.n62 GNDA 0.013267f
C446 VDDA.t105 GNDA 0.094896f
C447 VDDA.t78 GNDA 0.019901f
C448 VDDA.t86 GNDA 0.019901f
C449 VDDA.n63 GNDA 0.077433f
C450 VDDA.n64 GNDA 0.266192f
C451 VDDA.t142 GNDA 0.019901f
C452 VDDA.t69 GNDA 0.019901f
C453 VDDA.n65 GNDA 0.077433f
C454 VDDA.n66 GNDA 0.266192f
C455 VDDA.t76 GNDA 0.019901f
C456 VDDA.t136 GNDA 0.019901f
C457 VDDA.n67 GNDA 0.077433f
C458 VDDA.n68 GNDA 0.266192f
C459 VDDA.t25 GNDA 0.019901f
C460 VDDA.t9 GNDA 0.019901f
C461 VDDA.n69 GNDA 0.077433f
C462 VDDA.n70 GNDA 0.266192f
C463 VDDA.t6 GNDA 0.019901f
C464 VDDA.t74 GNDA 0.019901f
C465 VDDA.n71 GNDA 0.077433f
C466 VDDA.n72 GNDA 0.266192f
C467 VDDA.t64 GNDA 0.019901f
C468 VDDA.t93 GNDA 0.019901f
C469 VDDA.n73 GNDA 0.077433f
C470 VDDA.n74 GNDA 0.266192f
C471 VDDA.t21 GNDA 0.019901f
C472 VDDA.t80 GNDA 0.019901f
C473 VDDA.n75 GNDA 0.077433f
C474 VDDA.n76 GNDA 0.37925f
C475 VDDA.n77 GNDA 0.038327f
C476 VDDA.n80 GNDA 0.023079f
C477 VDDA.n81 GNDA 0.023079f
C478 VDDA.n82 GNDA 0.013267f
C479 VDDA.n83 GNDA 0.023218f
C480 VDDA.n85 GNDA 0.025023f
C481 VDDA.n86 GNDA 0.01871f
C482 VDDA.n88 GNDA 0.023218f
C483 VDDA.n89 GNDA 0.013267f
C484 VDDA.n90 GNDA 0.013267f
C485 VDDA.n91 GNDA 0.023218f
C486 VDDA.n92 GNDA 0.023218f
C487 VDDA.n93 GNDA 0.01871f
C488 VDDA.n94 GNDA 0.026509f
C489 VDDA.n95 GNDA 0.013267f
C490 VDDA.n96 GNDA 0.186075f
C491 VDDA.t106 GNDA 0.197352f
C492 VDDA.t20 GNDA 0.202991f
C493 VDDA.t79 GNDA 0.202991f
C494 VDDA.t63 GNDA 0.202991f
C495 VDDA.t92 GNDA 0.202991f
C496 VDDA.t5 GNDA 0.202991f
C497 VDDA.t73 GNDA 0.202991f
C498 VDDA.t24 GNDA 0.202991f
C499 VDDA.t8 GNDA 0.202991f
C500 VDDA.t75 GNDA 0.202991f
C501 VDDA.t135 GNDA 0.202991f
C502 VDDA.t141 GNDA 0.202991f
C503 VDDA.t68 GNDA 0.202991f
C504 VDDA.t77 GNDA 0.202991f
C505 VDDA.t85 GNDA 0.202991f
C506 VDDA.t41 GNDA 0.202991f
C507 VDDA.t151 GNDA 0.202991f
C508 VDDA.t112 GNDA 0.197352f
C509 VDDA.n98 GNDA 0.013267f
C510 VDDA.n99 GNDA 0.013267f
C511 VDDA.n100 GNDA 0.023218f
C512 VDDA.n102 GNDA 0.023218f
C513 VDDA.n103 GNDA 0.025023f
C514 VDDA.n105 GNDA 0.01871f
C515 VDDA.n106 GNDA 0.013267f
C516 VDDA.n107 GNDA 0.023218f
C517 VDDA.n109 GNDA 0.023079f
C518 VDDA.n110 GNDA 0.023079f
C519 VDDA.n111 GNDA 0.023218f
C520 VDDA.n112 GNDA 0.013267f
C521 VDDA.n113 GNDA 0.186075f
C522 VDDA.n114 GNDA 0.010297f
C523 VDDA.n115 GNDA 0.029479f
C524 VDDA.t111 GNDA 0.094896f
C525 VDDA.n116 GNDA 0.036375f
C526 VDDA.n117 GNDA 0.224466f
C527 VDDA.n118 GNDA 0.22135f
C528 VDDA.n119 GNDA 0.025793f
C529 VDDA.t104 GNDA 0.023074f
C530 VDDA.n120 GNDA 0.027319f
C531 VDDA.t98 GNDA 0.026323f
C532 VDDA.t96 GNDA 0.012982f
C533 VDDA.n121 GNDA 0.066189f
C534 VDDA.n122 GNDA 0.019524f
C535 VDDA.n123 GNDA 0.027123f
C536 VDDA.n124 GNDA 0.068643f
C537 VDDA.t97 GNDA 0.081971f
C538 VDDA.t33 GNDA 0.051079f
C539 VDDA.t87 GNDA 0.051079f
C540 VDDA.t103 GNDA 0.065489f
C541 VDDA.n125 GNDA 0.080481f
C542 VDDA.n126 GNDA 0.025597f
C543 VDDA.t102 GNDA 0.012923f
C544 VDDA.n128 GNDA 0.0818f
C545 VDDA.n129 GNDA 0.427736f
C546 VDDA.n130 GNDA 0.353662f
C547 VDDA.n132 GNDA 0.387956f
C548 VDDA.n134 GNDA 0.036183f
C549 VDDA.n135 GNDA 0.293209f
C550 VDDA.n136 GNDA 0.014043f
C551 VDDA.n137 GNDA 0.177339f
C552 VDDA.n138 GNDA 0.025793f
C553 VDDA.t128 GNDA 0.023074f
C554 VDDA.n139 GNDA 0.025793f
C555 VDDA.t122 GNDA 0.023074f
C556 VDDA.n140 GNDA 0.014043f
C557 VDDA.n141 GNDA 0.177339f
C558 VDDA.n142 GNDA 0.025793f
C559 VDDA.t131 GNDA 0.023074f
C560 VDDA.n143 GNDA 0.025793f
C561 VDDA.t125 GNDA 0.023074f
C562 VDDA.n144 GNDA 0.014043f
C563 VDDA.n145 GNDA 0.177339f
C564 VDDA.n146 GNDA 0.014043f
C565 VDDA.n147 GNDA 0.177339f
C566 VDDA.n148 GNDA 0.014043f
C567 VDDA.n149 GNDA 0.177339f
C568 VDDA.n150 GNDA 0.014043f
C569 VDDA.n151 GNDA 0.177339f
C570 VDDA.n152 GNDA 0.014043f
C571 VDDA.n153 GNDA 0.177339f
C572 VDDA.n154 GNDA 0.014043f
C573 VDDA.n155 GNDA 0.177339f
C574 VDDA.n156 GNDA 0.014043f
C575 VDDA.n157 GNDA 0.177339f
C576 VDDA.n158 GNDA 0.014043f
C577 VDDA.n159 GNDA 0.241638f
C578 VDDA.t123 GNDA 0.016536f
C579 VDDA.n160 GNDA 0.059302f
C580 VDDA.n161 GNDA 0.019705f
C581 VDDA.n162 GNDA 0.025597f
C582 VDDA.n163 GNDA 0.067233f
C583 VDDA.t124 GNDA 0.083381f
C584 VDDA.t145 GNDA 0.055723f
C585 VDDA.t45 GNDA 0.055723f
C586 VDDA.t156 GNDA 0.055723f
C587 VDDA.t137 GNDA 0.055723f
C588 VDDA.t18 GNDA 0.055723f
C589 VDDA.t81 GNDA 0.055723f
C590 VDDA.t3 GNDA 0.055723f
C591 VDDA.t35 GNDA 0.055723f
C592 VDDA.t158 GNDA 0.055723f
C593 VDDA.t10 GNDA 0.055723f
C594 VDDA.t147 GNDA 0.055723f
C595 VDDA.t51 GNDA 0.055723f
C596 VDDA.t154 GNDA 0.055723f
C597 VDDA.t59 GNDA 0.055723f
C598 VDDA.t83 GNDA 0.055723f
C599 VDDA.t47 GNDA 0.055723f
C600 VDDA.t53 GNDA 0.055723f
C601 VDDA.t43 GNDA 0.055723f
C602 VDDA.t130 GNDA 0.069408f
C603 VDDA.n164 GNDA 0.085849f
C604 VDDA.n165 GNDA 0.025597f
C605 VDDA.t129 GNDA 0.016536f
C606 VDDA.n167 GNDA 0.073038f
C607 VDDA.n168 GNDA 0.180271f
C608 VDDA.n169 GNDA 0.014043f
C609 VDDA.n170 GNDA 0.177339f
C610 VDDA.n171 GNDA 0.014043f
C611 VDDA.n172 GNDA 0.177339f
C612 VDDA.n173 GNDA 0.014043f
C613 VDDA.n174 GNDA 0.177339f
C614 VDDA.n175 GNDA 0.014043f
C615 VDDA.n176 GNDA 0.177339f
C616 VDDA.n177 GNDA 0.014043f
C617 VDDA.n178 GNDA 0.177339f
C618 VDDA.n179 GNDA 0.014043f
C619 VDDA.n180 GNDA 0.177339f
C620 VDDA.n181 GNDA 0.014043f
C621 VDDA.n182 GNDA 0.177339f
C622 VDDA.n183 GNDA 0.014043f
C623 VDDA.n184 GNDA 0.177339f
C624 VDDA.n185 GNDA 0.180271f
C625 VDDA.t120 GNDA 0.016536f
C626 VDDA.n186 GNDA 0.054776f
C627 VDDA.n187 GNDA 0.019705f
C628 VDDA.n188 GNDA 0.025597f
C629 VDDA.n189 GNDA 0.070586f
C630 VDDA.t121 GNDA 0.084671f
C631 VDDA.t1 GNDA 0.055723f
C632 VDDA.t39 GNDA 0.055723f
C633 VDDA.t12 GNDA 0.055723f
C634 VDDA.t14 GNDA 0.055723f
C635 VDDA.t139 GNDA 0.055723f
C636 VDDA.t200 GNDA 0.055723f
C637 VDDA.t88 GNDA 0.055723f
C638 VDDA.t22 GNDA 0.055723f
C639 VDDA.t71 GNDA 0.055723f
C640 VDDA.t16 GNDA 0.055723f
C641 VDDA.t29 GNDA 0.055723f
C642 VDDA.t65 GNDA 0.055723f
C643 VDDA.t55 GNDA 0.055723f
C644 VDDA.t37 GNDA 0.055723f
C645 VDDA.t94 GNDA 0.055723f
C646 VDDA.t149 GNDA 0.055723f
C647 VDDA.t31 GNDA 0.055723f
C648 VDDA.t132 GNDA 0.055723f
C649 VDDA.t127 GNDA 0.068843f
C650 VDDA.n190 GNDA 0.081771f
C651 VDDA.n191 GNDA 0.025597f
C652 VDDA.t126 GNDA 0.016536f
C653 VDDA.n193 GNDA 0.073038f
C654 VDDA.n194 GNDA 0.378698f
C655 VDDA.n195 GNDA 0.347691f
C656 VDDA.n197 GNDA 0.293209f
C657 VDDA.n199 GNDA 0.036183f
C658 VDDA.n200 GNDA 0.381603f
C659 VDDA.t205 GNDA 0.735431f
C660 VDDA.t204 GNDA 0.783652f
C661 VDDA.t203 GNDA 0.783652f
C662 VDDA.t202 GNDA 0.744502f
C663 VDDA.n201 GNDA 1.44119f
C664 VDDA.n202 GNDA 0.760732f
C665 VDDA.n203 GNDA 0.982356f
C666 VDDA.n204 GNDA 0.523732f
C667 VDDA.n206 GNDA 0.381603f
C668 VDDA.n208 GNDA 0.036183f
C669 VDDA.n209 GNDA 0.551922f
C670 VDDA.t50 GNDA 0.352266f
C671 VDDA.t91 GNDA 0.370823f
C672 VDDA.t34 GNDA 0.372167f
C673 VDDA.t153 GNDA 0.352266f
C674 VDDA.t26 GNDA 0.370823f
C675 VDDA.t70 GNDA 0.372167f
C676 VDDA.t28 GNDA 0.352266f
C677 VDDA.t90 GNDA 0.370823f
C678 VDDA.t7 GNDA 0.372167f
C679 VDDA.t27 GNDA 0.352266f
C680 VDDA.t67 GNDA 0.370823f
C681 VDDA.t0 GNDA 0.372167f
C682 VDDA.t144 GNDA 0.352266f
C683 VDDA.t61 GNDA 0.370823f
C684 VDDA.t143 GNDA 0.372167f
C685 VDDA.n210 GNDA 0.248563f
C686 VDDA.t62 GNDA 0.197944f
C687 VDDA.n211 GNDA 0.269697f
C688 VDDA.t58 GNDA 0.197944f
C689 VDDA.n212 GNDA 0.269697f
C690 VDDA.t49 GNDA 0.197944f
C691 VDDA.n213 GNDA 0.269697f
C692 VDDA.t134 GNDA 0.197944f
C693 VDDA.n214 GNDA 0.269697f
C694 VDDA.t57 GNDA 0.523916f
C695 V2.t24 GNDA 0.029604f
C696 V2.t13 GNDA 0.029569f
C697 V2.n0 GNDA 0.15465f
C698 V2.t21 GNDA 0.029569f
C699 V2.n1 GNDA 0.081084f
C700 V2.t11 GNDA 0.029569f
C701 V2.n2 GNDA 0.081084f
C702 V2.t19 GNDA 0.029569f
C703 V2.n3 GNDA 0.081084f
C704 V2.t29 GNDA 0.029569f
C705 V2.n4 GNDA 0.081084f
C706 V2.t15 GNDA 0.029569f
C707 V2.n5 GNDA 0.081084f
C708 V2.t22 GNDA 0.029569f
C709 V2.n6 GNDA 0.081084f
C710 V2.t18 GNDA 0.029569f
C711 V2.n7 GNDA 0.081084f
C712 V2.t27 GNDA 0.029569f
C713 V2.n8 GNDA 0.200801f
C714 V2.t26 GNDA 0.029569f
C715 V2.n9 GNDA 0.200801f
C716 V2.t16 GNDA 0.029569f
C717 V2.n10 GNDA 0.081084f
C718 V2.t23 GNDA 0.029569f
C719 V2.n11 GNDA 0.081084f
C720 V2.t12 GNDA 0.029569f
C721 V2.n12 GNDA 0.081084f
C722 V2.t20 GNDA 0.029569f
C723 V2.n13 GNDA 0.081084f
C724 V2.t10 GNDA 0.029569f
C725 V2.n14 GNDA 0.081084f
C726 V2.t17 GNDA 0.029569f
C727 V2.n15 GNDA 0.081084f
C728 V2.t25 GNDA 0.029569f
C729 V2.n16 GNDA 0.081084f
C730 V2.t14 GNDA 0.029569f
C731 V2.n17 GNDA 0.081084f
C732 V2.t28 GNDA 0.029569f
C733 V2.n18 GNDA 0.642575f
C734 V2.t5 GNDA 0.263098f
C735 V2.t2 GNDA 0.017102f
C736 V2.t6 GNDA 0.017102f
C737 V2.n19 GNDA 0.036943f
C738 V2.n20 GNDA 0.891145f
C739 V2.t3 GNDA 0.017102f
C740 V2.t9 GNDA 0.017102f
C741 V2.n21 GNDA 0.036943f
C742 V2.n22 GNDA 0.373516f
C743 V2.t4 GNDA 0.017102f
C744 V2.t0 GNDA 0.017102f
C745 V2.n23 GNDA 0.036943f
C746 V2.n24 GNDA 0.36582f
C747 V2.t7 GNDA 0.017102f
C748 V2.t8 GNDA 0.017102f
C749 V2.n25 GNDA 0.036943f
C750 V2.n26 GNDA 0.496771f
C751 V2.n27 GNDA 2.55195f
C752 V2.t1 GNDA 0.266609f
.ends

