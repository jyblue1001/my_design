* PEX produced on Thu Feb 20 09:58:47 AM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from vco2_3.ext - technology: sky130A

.subckt current_starved_VCO_magic VDDA V_OSC V_CONT GNDA
X0 a_4510_n870.t1 VDDA.t14 GNDA.t7 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X1 a_3310_n50.t2 a_2390_720.t3 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X2 a_4510_n870.t0 V_OSC.t2 a_3880_n330.t1 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.2 as=0.28 ps=2.2 w=0.7 l=0.15
X3 a_3910_n870.t0 VDDA.t15 GNDA.t6 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X4 a_3310_n50.t1 a_3280_n330.t2 V_OSC.t1 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.56 pd=3.6 as=0.56 ps=3.6 w=1.4 l=0.15
X5 a_4510_n870.t2 V_CONT.t0 GNDA.t8 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X6 a_4510_n50.t2 a_2390_720.t4 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X7 a_3910_n870.t2 a_3880_n330.t2 a_3280_n330.t1 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.2 as=0.28 ps=2.2 w=0.7 l=0.15
X8 a_3910_n50.t1 a_2390_720.t5 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X9 a_3910_n870.t1 V_CONT.t1 GNDA.t9 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X10 a_4510_n50.t1 V_OSC.t3 a_3880_n330.t0 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.56 pd=3.6 as=0.56 ps=3.6 w=1.4 l=0.15
X11 GNDA.t3 V_CONT.t2 a_2390_720.t0 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X12 a_3310_n50.t0 GNDA.t11 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X13 a_3910_n50.t2 a_3880_n330.t3 a_3280_n330.t0 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.56 pd=3.6 as=0.56 ps=3.6 w=1.4 l=0.15
X14 a_4510_n50.t0 GNDA.t12 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X15 VDDA.t3 a_2390_720.t1 a_2390_720.t2 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X16 a_3910_n50.t0 GNDA.t13 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X17 a_3310_n870.t0 VDDA.t16 GNDA.t5 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X18 a_3310_n870.t1 a_3280_n330.t3 V_OSC.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.2 as=0.28 ps=2.2 w=0.7 l=0.15
X19 a_3310_n870.t2 V_CONT.t3 GNDA.t10 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
R0 VDDA.n23 VDDA.n22 831.25
R1 VDDA.n21 VDDA.n18 831.25
R2 VDDA.n22 VDDA.n20 585
R3 VDDA.n26 VDDA.n21 585
R4 VDDA.n7 VDDA.t14 537.866
R5 VDDA.n16 VDDA.t16 537.866
R6 VDDA.n14 VDDA.t15 537.866
R7 VDDA.t5 VDDA.n24 465.079
R8 VDDA.n25 VDDA.t5 465.079
R9 VDDA.t7 VDDA.n5 464.281
R10 VDDA.n10 VDDA.t7 464.281
R11 VDDA.t1 VDDA.n31 464.281
R12 VDDA.n33 VDDA.t1 464.281
R13 VDDA.n16 VDDA.t13 359.752
R14 VDDA.n14 VDDA.t9 359.752
R15 VDDA.n7 VDDA.t11 359.752
R16 VDDA.n41 VDDA.n40 238.367
R17 VDDA.n13 VDDA.n8 238.367
R18 VDDA.n37 VDDA.n4 238.367
R19 VDDA.n32 VDDA.n15 238.367
R20 VDDA.n28 VDDA.n18 238.367
R21 VDDA.n23 VDDA.n17 238.367
R22 VDDA.n39 VDDA.t6 205.201
R23 VDDA.t0 VDDA.n38 205.201
R24 VDDA.t4 VDDA.n29 205.201
R25 VDDA.n29 VDDA.t2 205.201
R26 VDDA.t4 VDDA.n16 185.002
R27 VDDA.t0 VDDA.n14 185.002
R28 VDDA.n7 VDDA.t6 185.002
R29 VDDA.n36 VDDA.n35 185
R30 VDDA.n34 VDDA.n30 185
R31 VDDA.n20 VDDA.n19 185
R32 VDDA.n27 VDDA.n26 185
R33 VDDA.n9 VDDA.n6 185
R34 VDDA.n12 VDDA.n11 185
R35 VDDA.n12 VDDA.n6 150
R36 VDDA.n27 VDDA.n19 150
R37 VDDA.n36 VDDA.n30 150
R38 VDDA.n39 VDDA.t8 148.201
R39 VDDA.n38 VDDA.t12 148.201
R40 VDDA.n22 VDDA.t3 123.126
R41 VDDA.t3 VDDA.n21 123.126
R42 VDDA.t6 VDDA.t10 102.6
R43 VDDA.t8 VDDA.t0 102.6
R44 VDDA.t12 VDDA.t4 102.6
R45 VDDA.n18 VDDA.n16 90.5056
R46 VDDA.n8 VDDA.n7 74.7688
R47 VDDA.n32 VDDA.n14 74.7687
R48 VDDA.n38 VDDA.n37 65.8183
R49 VDDA.n38 VDDA.n15 65.8183
R50 VDDA.n29 VDDA.n17 65.8183
R51 VDDA.n29 VDDA.n28 65.8183
R52 VDDA.n40 VDDA.n39 65.8183
R53 VDDA.n39 VDDA.n13 65.8183
R54 VDDA.n19 VDDA.n17 53.3664
R55 VDDA.n28 VDDA.n27 53.3664
R56 VDDA.n37 VDDA.n36 53.3664
R57 VDDA.n30 VDDA.n15 53.3664
R58 VDDA.n40 VDDA.n6 53.3664
R59 VDDA.n13 VDDA.n12 53.3664
R60 VDDA.n45 VDDA.n44 32.0005
R61 VDDA.n45 VDDA.n2 32.0005
R62 VDDA.n49 VDDA.n2 32.0005
R63 VDDA.n50 VDDA.n49 32.0005
R64 VDDA.n51 VDDA.n50 32.0005
R65 VDDA.n42 VDDA.n41 31.5568
R66 VDDA.n43 VDDA.n4 24.991
R67 VDDA.n23 VDDA.n0 23.6611
R68 VDDA.n44 VDDA.n43 22.4005
R69 VDDA.n51 VDDA.n0 16.0005
R70 VDDA.n44 VDDA.n3 9.3005
R71 VDDA.n46 VDDA.n45 9.3005
R72 VDDA.n47 VDDA.n2 9.3005
R73 VDDA.n49 VDDA.n48 9.3005
R74 VDDA.n50 VDDA.n1 9.3005
R75 VDDA.n52 VDDA.n51 9.3005
R76 VDDA.n35 VDDA.n34 9.14336
R77 VDDA.n11 VDDA.n9 9.14336
R78 VDDA.n53 VDDA.n0 7.37301
R79 VDDA.n43 VDDA.n42 7.05917
R80 VDDA.n26 VDDA.n20 5.81868
R81 VDDA.n31 VDDA.n4 5.33286
R82 VDDA.n33 VDDA.n32 5.33286
R83 VDDA.n41 VDDA.n5 5.33286
R84 VDDA.n10 VDDA.n8 5.33286
R85 VDDA.n35 VDDA.n31 3.75335
R86 VDDA.n34 VDDA.n33 3.75335
R87 VDDA.n9 VDDA.n5 3.75335
R88 VDDA.n11 VDDA.n10 3.75335
R89 VDDA.n24 VDDA.n23 3.40194
R90 VDDA.n25 VDDA.n18 3.40194
R91 VDDA.n24 VDDA.n20 2.39444
R92 VDDA.n26 VDDA.n25 2.39444
R93 VDDA VDDA.n53 0.712019
R94 VDDA.n42 VDDA.n3 0.203454
R95 VDDA.n53 VDDA.n52 0.196483
R96 VDDA.n46 VDDA.n3 0.15675
R97 VDDA.n47 VDDA.n46 0.15675
R98 VDDA.n48 VDDA.n47 0.15675
R99 VDDA.n48 VDDA.n1 0.15675
R100 VDDA.n52 VDDA.n1 0.15675
R101 GNDA.n7 GNDA.t4 2131.25
R102 GNDA.t0 GNDA.n29 2131.25
R103 GNDA.n29 GNDA.n28 1173.78
R104 GNDA.n8 GNDA.n7 1173.78
R105 GNDA.n31 GNDA.n30 1173.78
R106 GNDA.n28 GNDA.t13 728.899
R107 GNDA.n8 GNDA.t12 728.899
R108 GNDA.n31 GNDA.t11 728.899
R109 GNDA.n33 GNDA.n2 686.717
R110 GNDA.n26 GNDA.n4 686.717
R111 GNDA.n11 GNDA.n10 686.717
R112 GNDA.n12 GNDA.n11 686.717
R113 GNDA.n24 GNDA.n4 686.717
R114 GNDA.n34 GNDA.n2 686.717
R115 GNDA.n7 GNDA.t1 618.75
R116 GNDA.n29 GNDA.t4 618.75
R117 GNDA.n30 GNDA.t0 618.75
R118 GNDA.n30 GNDA.t2 618.75
R119 GNDA.t3 GNDA.n33 260
R120 GNDA.n34 GNDA.t3 260
R121 GNDA.n11 GNDA.n7 241.643
R122 GNDA.n29 GNDA.n4 241.643
R123 GNDA.n30 GNDA.n2 241.643
R124 GNDA.n27 GNDA.t6 233
R125 GNDA.n9 GNDA.t7 233
R126 GNDA.n32 GNDA.t5 233
R127 GNDA.n3 GNDA.t10 128.562
R128 GNDA.n25 GNDA.t9 127.754
R129 GNDA.n6 GNDA.t8 127.754
R130 GNDA.n22 GNDA.n12 41.9648
R131 GNDA.n27 GNDA.n26 35.6576
R132 GNDA.n24 GNDA.n23 35.6576
R133 GNDA.n10 GNDA.n9 35.6576
R134 GNDA.n33 GNDA.n32 34.3278
R135 GNDA.n35 GNDA.n34 34.3278
R136 GNDA.n19 GNDA.n5 32.0005
R137 GNDA.n19 GNDA.n18 32.0005
R138 GNDA.n18 GNDA.n17 32.0005
R139 GNDA.n17 GNDA.n14 32.0005
R140 GNDA.n14 GNDA.n1 32.0005
R141 GNDA.n35 GNDA.n1 25.6005
R142 GNDA.n23 GNDA.n5 12.8005
R143 GNDA.n21 GNDA.n5 9.3005
R144 GNDA.n20 GNDA.n19 9.3005
R145 GNDA.n18 GNDA.n13 9.3005
R146 GNDA.n17 GNDA.n16 9.3005
R147 GNDA.n15 GNDA.n14 9.3005
R148 GNDA.n1 GNDA.n0 9.3005
R149 GNDA.n23 GNDA.n22 7.49828
R150 GNDA.n36 GNDA.n35 6.86152
R151 GNDA.n25 GNDA.n24 4.49344
R152 GNDA.n26 GNDA.n25 4.49344
R153 GNDA.n12 GNDA.n6 4.49344
R154 GNDA.n10 GNDA.n6 4.49344
R155 GNDA.n28 GNDA.n27 3.8278
R156 GNDA.n9 GNDA.n8 3.8278
R157 GNDA.n32 GNDA.n31 3.8278
R158 GNDA.n34 GNDA.n3 2.8779
R159 GNDA.n33 GNDA.n3 2.8779
R160 GNDA GNDA.n36 1.17078
R161 GNDA.n36 GNDA.n0 0.206966
R162 GNDA.n22 GNDA.n21 0.194576
R163 GNDA.n21 GNDA.n20 0.15675
R164 GNDA.n20 GNDA.n13 0.15675
R165 GNDA.n16 GNDA.n13 0.15675
R166 GNDA.n16 GNDA.n15 0.15675
R167 GNDA.n15 GNDA.n0 0.15675
R168 a_4510_n870.n0 a_4510_n870.t0 274.752
R169 a_4510_n870.n0 a_4510_n870.t1 233
R170 a_4510_n870.t2 a_4510_n870.n0 184.191
R171 a_2390_720.n0 a_2390_720.t4 600.206
R172 a_2390_720.n1 a_2390_720.n0 568.072
R173 a_2390_720.t0 a_2390_720.n5 458.399
R174 a_2390_720.n2 a_2390_720.n1 392.486
R175 a_2390_720.n4 a_2390_720.t2 289.791
R176 a_2390_720.n5 a_2390_720.n2 168.067
R177 a_2390_720.n4 a_2390_720.n3 97.9242
R178 a_2390_720.n3 a_2390_720.n2 37.7572
R179 a_2390_720.n0 a_2390_720.t5 32.1338
R180 a_2390_720.n1 a_2390_720.t3 32.1338
R181 a_2390_720.n3 a_2390_720.t1 32.1338
R182 a_2390_720.n5 a_2390_720.n4 28.3357
R183 a_3310_n50.n0 a_3310_n50.t0 348.81
R184 a_3310_n50.n0 a_3310_n50.t2 316.159
R185 a_3310_n50.t1 a_3310_n50.n0 295.204
R186 V_OSC.n2 V_OSC.n1 386.233
R187 V_OSC.n1 V_OSC.t3 289.2
R188 V_OSC.n0 V_OSC.t1 246.294
R189 V_OSC.n0 V_OSC.t0 238.487
R190 V_OSC.n1 V_OSC.t2 176.733
R191 V_OSC.n2 V_OSC.n0 75.6755
R192 V_OSC V_OSC.n2 0.063
R193 a_3880_n330.n1 a_3880_n330.n0 437.733
R194 a_3880_n330.n0 a_3880_n330.t3 289.2
R195 a_3880_n330.t0 a_3880_n330.n1 246.294
R196 a_3880_n330.n1 a_3880_n330.t1 238.487
R197 a_3880_n330.n0 a_3880_n330.t2 176.733
R198 a_3910_n870.n0 a_3910_n870.t2 274.752
R199 a_3910_n870.n0 a_3910_n870.t0 233
R200 a_3910_n870.t1 a_3910_n870.n0 184.191
R201 a_3280_n330.n1 a_3280_n330.n0 437.733
R202 a_3280_n330.n0 a_3280_n330.t2 289.2
R203 a_3280_n330.t0 a_3280_n330.n1 246.294
R204 a_3280_n330.n1 a_3280_n330.t1 238.487
R205 a_3280_n330.n0 a_3280_n330.t3 176.733
R206 V_CONT.n0 V_CONT.t0 1156.8
R207 V_CONT.n1 V_CONT.n0 964
R208 V_CONT V_CONT.n2 565.011
R209 V_CONT.n2 V_CONT.n1 417.733
R210 V_CONT.n1 V_CONT.t3 192.8
R211 V_CONT.n0 V_CONT.t1 192.8
R212 V_CONT.n2 V_CONT.t2 192.8
R213 a_4510_n50.n0 a_4510_n50.t0 348.81
R214 a_4510_n50.n0 a_4510_n50.t2 316.159
R215 a_4510_n50.t1 a_4510_n50.n0 295.204
R216 a_3910_n50.n0 a_3910_n50.t0 348.81
R217 a_3910_n50.n0 a_3910_n50.t1 316.159
R218 a_3910_n50.t2 a_3910_n50.n0 295.204
R219 a_3310_n870.n0 a_3310_n870.t1 274.752
R220 a_3310_n870.n0 a_3310_n870.t0 233
R221 a_3310_n870.t2 a_3310_n870.n0 184.191
C0 V_OSC V_CONT 0.073017f
C1 VDDA V_CONT 0.090222f
C2 V_OSC VDDA 0.430141f
C3 V_CONT GNDA 1.58413f
C4 V_OSC GNDA 2.62496f
C5 VDDA GNDA 12.370811f
C6 a_2390_720.t3 GNDA 0.284469f
C7 a_2390_720.t5 GNDA 0.284469f
C8 a_2390_720.t4 GNDA 0.473934f
C9 a_2390_720.n0 GNDA 0.231971f
C10 a_2390_720.n1 GNDA 0.207751f
C11 a_2390_720.n2 GNDA 0.043218f
C12 a_2390_720.t2 GNDA 0.099803f
C13 a_2390_720.t1 GNDA 0.284469f
C14 a_2390_720.n3 GNDA 0.16127f
C15 a_2390_720.n4 GNDA 0.175764f
C16 a_2390_720.n5 GNDA 0.260394f
C17 a_2390_720.t0 GNDA 0.192487f
C18 VDDA.n4 GNDA 0.012737f
C19 VDDA.t10 GNDA 0.17048f
C20 VDDA.t6 GNDA 0.175868f
C21 VDDA.n7 GNDA 0.073352f
C22 VDDA.n8 GNDA 0.018249f
C23 VDDA.t7 GNDA 0.014205f
C24 VDDA.n14 GNDA 0.073352f
C25 VDDA.n16 GNDA 0.074722f
C26 VDDA.t2 GNDA 0.34096f
C27 VDDA.n18 GNDA 0.026557f
C28 VDDA.n20 GNDA 0.014817f
C29 VDDA.n23 GNDA 0.019264f
C30 VDDA.t5 GNDA 0.014212f
C31 VDDA.n26 GNDA 0.014817f
C32 VDDA.n29 GNDA 0.227307f
C33 VDDA.t4 GNDA 0.175868f
C34 VDDA.t12 GNDA 0.13891f
C35 VDDA.n32 GNDA 0.018249f
C36 VDDA.t1 GNDA 0.014205f
C37 VDDA.n38 GNDA 0.195736f
C38 VDDA.t0 GNDA 0.175868f
C39 VDDA.t8 GNDA 0.13891f
C40 VDDA.n39 GNDA 0.195736f
C41 VDDA.n41 GNDA 0.015859f
C42 VDDA.n42 GNDA 0.088482f
C43 VDDA.n53 GNDA 0.019789f
.ends

