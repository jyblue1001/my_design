magic
tech sky130A
timestamp 1753019775
<< nwell >>
rect 56025 4340 56365 4730
rect 56495 4340 56835 4560
rect 56965 4340 57305 4730
rect 57435 4340 57775 4730
rect 54865 3670 55745 4060
rect 55945 3670 56825 4060
rect 56975 3670 57855 4060
rect 58060 3670 58940 4060
rect 54890 2730 55710 3370
rect 56215 3285 57585 3375
rect 55970 2925 56790 3015
rect 57010 2925 57830 3015
rect 58090 2730 58910 3370
rect 54890 2200 55710 2440
rect 58090 2200 58910 2440
<< nmos >>
rect 56590 2535 56605 2585
rect 56645 2535 56660 2585
rect 56700 2535 56715 2585
rect 56755 2535 56770 2585
rect 56810 2535 56825 2585
rect 56865 2535 56880 2585
rect 56920 2535 56935 2585
rect 56975 2535 56990 2585
rect 57030 2535 57045 2585
rect 57085 2535 57100 2585
rect 57140 2535 57155 2585
rect 57195 2535 57210 2585
rect 56070 2030 56085 2180
rect 56125 2030 56140 2180
rect 56180 2030 56195 2180
rect 56235 2030 56250 2180
rect 56290 2030 56305 2180
rect 56345 2030 56360 2180
rect 56400 2030 56415 2180
rect 56455 2030 56470 2180
rect 56510 2030 56525 2180
rect 56565 2030 56580 2180
rect 56620 2030 56635 2180
rect 56675 2030 56690 2180
rect 57110 2030 57125 2180
rect 57165 2030 57180 2180
rect 57220 2030 57235 2180
rect 57275 2030 57290 2180
rect 57330 2030 57345 2180
rect 57385 2030 57400 2180
rect 57440 2030 57455 2180
rect 57495 2030 57510 2180
rect 57550 2030 57565 2180
rect 57605 2030 57620 2180
rect 57660 2030 57675 2180
rect 57715 2030 57730 2180
rect 54990 1560 55005 1860
rect 55045 1560 55060 1860
rect 55100 1560 55115 1860
rect 55155 1560 55170 1860
rect 55210 1560 55225 1860
rect 55265 1560 55280 1860
rect 55320 1560 55335 1860
rect 55375 1560 55390 1860
rect 55430 1560 55445 1860
rect 55485 1560 55500 1860
rect 55540 1560 55555 1860
rect 55595 1560 55610 1860
rect 56070 1560 56085 1710
rect 56125 1560 56140 1710
rect 56180 1560 56195 1710
rect 56235 1560 56250 1710
rect 56290 1560 56305 1710
rect 56345 1560 56360 1710
rect 56400 1560 56415 1710
rect 56455 1560 56470 1710
rect 56510 1560 56525 1710
rect 56565 1560 56580 1710
rect 56620 1560 56635 1710
rect 56675 1560 56690 1710
rect 56810 1560 56825 1710
rect 56865 1560 56880 1710
rect 56920 1560 56935 1710
rect 56975 1560 56990 1710
rect 57110 1560 57125 1710
rect 57165 1560 57180 1710
rect 57220 1560 57235 1710
rect 57275 1560 57290 1710
rect 57330 1560 57345 1710
rect 57385 1560 57400 1710
rect 57440 1560 57455 1710
rect 57495 1560 57510 1710
rect 57550 1560 57565 1710
rect 57605 1560 57620 1710
rect 57660 1560 57675 1710
rect 57715 1560 57730 1710
rect 58190 1560 58205 1860
rect 58245 1560 58260 1860
rect 58300 1560 58315 1860
rect 58355 1560 58370 1860
rect 58410 1560 58425 1860
rect 58465 1560 58480 1860
rect 58520 1560 58535 1860
rect 58575 1560 58590 1860
rect 58630 1560 58645 1860
rect 58685 1560 58700 1860
rect 58740 1560 58755 1860
rect 58795 1560 58810 1860
rect 55025 470 55085 1170
rect 55125 470 55185 1170
rect 55225 470 55285 1170
rect 55325 470 55385 1170
rect 55425 470 55485 1170
rect 55525 470 55585 1170
rect 56260 910 56275 1160
rect 56315 910 56330 1160
rect 56370 910 56385 1160
rect 56425 910 56440 1160
rect 56480 910 56495 1160
rect 56535 910 56550 1160
rect 56590 910 56605 1160
rect 56645 910 56660 1160
rect 56700 910 56715 1160
rect 56755 910 56770 1160
rect 56810 910 56825 1160
rect 56865 910 56880 1160
rect 56920 910 56935 1160
rect 56975 910 56990 1160
rect 57030 910 57045 1160
rect 57085 910 57100 1160
rect 57140 910 57155 1160
rect 57195 910 57210 1160
rect 57250 910 57265 1160
rect 57305 910 57320 1160
rect 57360 910 57375 1160
rect 57415 910 57430 1160
rect 57470 910 57485 1160
rect 56470 545 56485 695
rect 56525 545 56540 695
rect 56580 545 56595 695
rect 56635 545 56650 695
rect 56690 545 56705 695
rect 56745 545 56760 695
rect 56910 545 57210 695
rect 58220 470 58280 1170
rect 58320 470 58380 1170
rect 58420 470 58480 1170
rect 58520 470 58580 1170
rect 58620 470 58680 1170
rect 58720 470 58780 1170
<< pmos >>
rect 56125 4360 56145 4710
rect 56185 4360 56205 4710
rect 56245 4360 56265 4710
rect 56595 4360 56615 4540
rect 56655 4360 56675 4540
rect 56715 4360 56735 4540
rect 57065 4360 57085 4710
rect 57125 4360 57145 4710
rect 57185 4360 57205 4710
rect 57535 4360 57555 4710
rect 57595 4360 57615 4710
rect 57655 4360 57675 4710
rect 54965 3690 54985 4040
rect 55025 3690 55045 4040
rect 55085 3690 55105 4040
rect 55145 3690 55165 4040
rect 55205 3690 55225 4040
rect 55265 3690 55285 4040
rect 55325 3690 55345 4040
rect 55385 3690 55405 4040
rect 55445 3690 55465 4040
rect 55505 3690 55525 4040
rect 55565 3690 55585 4040
rect 55625 3690 55645 4040
rect 56045 3690 56065 4040
rect 56105 3690 56125 4040
rect 56165 3690 56185 4040
rect 56225 3690 56245 4040
rect 56285 3690 56305 4040
rect 56345 3690 56365 4040
rect 56405 3690 56425 4040
rect 56465 3690 56485 4040
rect 56525 3690 56545 4040
rect 56585 3690 56605 4040
rect 56645 3690 56665 4040
rect 56705 3690 56725 4040
rect 57075 3690 57095 4040
rect 57135 3690 57155 4040
rect 57195 3690 57215 4040
rect 57255 3690 57275 4040
rect 57315 3690 57335 4040
rect 57375 3690 57395 4040
rect 57435 3690 57455 4040
rect 57495 3690 57515 4040
rect 57555 3690 57575 4040
rect 57615 3690 57635 4040
rect 57675 3690 57695 4040
rect 57735 3690 57755 4040
rect 58160 3690 58180 4040
rect 58220 3690 58240 4040
rect 58280 3690 58300 4040
rect 58340 3690 58360 4040
rect 58400 3690 58420 4040
rect 58460 3690 58480 4040
rect 58520 3690 58540 4040
rect 58580 3690 58600 4040
rect 58640 3690 58660 4040
rect 58700 3690 58720 4040
rect 58760 3690 58780 4040
rect 58820 3690 58840 4040
rect 54990 2750 55005 3350
rect 55045 2750 55060 3350
rect 55100 2750 55115 3350
rect 55155 2750 55170 3350
rect 55210 2750 55225 3350
rect 55265 2750 55280 3350
rect 55320 2750 55335 3350
rect 55375 2750 55390 3350
rect 55430 2750 55445 3350
rect 55485 2750 55500 3350
rect 55540 2750 55555 3350
rect 55595 2750 55610 3350
rect 56315 3305 56330 3355
rect 56370 3305 56385 3355
rect 56425 3305 56440 3355
rect 56480 3305 56495 3355
rect 56535 3305 56550 3355
rect 56590 3305 56605 3355
rect 56645 3305 56660 3355
rect 56700 3305 56715 3355
rect 56755 3305 56770 3355
rect 56810 3305 56825 3355
rect 56865 3305 56880 3355
rect 56920 3305 56935 3355
rect 56975 3305 56990 3355
rect 57030 3305 57045 3355
rect 57085 3305 57100 3355
rect 57140 3305 57155 3355
rect 57195 3305 57210 3355
rect 57250 3305 57265 3355
rect 57305 3305 57320 3355
rect 57360 3305 57375 3355
rect 57415 3305 57430 3355
rect 57470 3305 57485 3355
rect 56070 2945 56085 2995
rect 56125 2945 56140 2995
rect 56180 2945 56195 2995
rect 56235 2945 56250 2995
rect 56290 2945 56305 2995
rect 56345 2945 56360 2995
rect 56400 2945 56415 2995
rect 56455 2945 56470 2995
rect 56510 2945 56525 2995
rect 56565 2945 56580 2995
rect 56620 2945 56635 2995
rect 56675 2945 56690 2995
rect 57110 2945 57125 2995
rect 57165 2945 57180 2995
rect 57220 2945 57235 2995
rect 57275 2945 57290 2995
rect 57330 2945 57345 2995
rect 57385 2945 57400 2995
rect 57440 2945 57455 2995
rect 57495 2945 57510 2995
rect 57550 2945 57565 2995
rect 57605 2945 57620 2995
rect 57660 2945 57675 2995
rect 57715 2945 57730 2995
rect 58190 2750 58205 3350
rect 58245 2750 58260 3350
rect 58300 2750 58315 3350
rect 58355 2750 58370 3350
rect 58410 2750 58425 3350
rect 58465 2750 58480 3350
rect 58520 2750 58535 3350
rect 58575 2750 58590 3350
rect 58630 2750 58645 3350
rect 58685 2750 58700 3350
rect 58740 2750 58755 3350
rect 58795 2750 58810 3350
rect 54990 2220 55005 2420
rect 55045 2220 55060 2420
rect 55100 2220 55115 2420
rect 55155 2220 55170 2420
rect 55210 2220 55225 2420
rect 55265 2220 55280 2420
rect 55320 2220 55335 2420
rect 55375 2220 55390 2420
rect 55430 2220 55445 2420
rect 55485 2220 55500 2420
rect 55540 2220 55555 2420
rect 55595 2220 55610 2420
rect 58190 2220 58205 2420
rect 58245 2220 58260 2420
rect 58300 2220 58315 2420
rect 58355 2220 58370 2420
rect 58410 2220 58425 2420
rect 58465 2220 58480 2420
rect 58520 2220 58535 2420
rect 58575 2220 58590 2420
rect 58630 2220 58645 2420
rect 58685 2220 58700 2420
rect 58740 2220 58755 2420
rect 58795 2220 58810 2420
<< ndiff >>
rect 56550 2570 56590 2585
rect 56550 2550 56560 2570
rect 56580 2550 56590 2570
rect 56550 2535 56590 2550
rect 56605 2570 56645 2585
rect 56605 2550 56615 2570
rect 56635 2550 56645 2570
rect 56605 2535 56645 2550
rect 56660 2570 56700 2585
rect 56660 2550 56670 2570
rect 56690 2550 56700 2570
rect 56660 2535 56700 2550
rect 56715 2570 56755 2585
rect 56715 2550 56725 2570
rect 56745 2550 56755 2570
rect 56715 2535 56755 2550
rect 56770 2570 56810 2585
rect 56770 2550 56780 2570
rect 56800 2550 56810 2570
rect 56770 2535 56810 2550
rect 56825 2570 56865 2585
rect 56825 2550 56835 2570
rect 56855 2550 56865 2570
rect 56825 2535 56865 2550
rect 56880 2570 56920 2585
rect 56880 2550 56890 2570
rect 56910 2550 56920 2570
rect 56880 2535 56920 2550
rect 56935 2570 56975 2585
rect 56935 2550 56945 2570
rect 56965 2550 56975 2570
rect 56935 2535 56975 2550
rect 56990 2570 57030 2585
rect 56990 2550 57000 2570
rect 57020 2550 57030 2570
rect 56990 2535 57030 2550
rect 57045 2570 57085 2585
rect 57045 2550 57055 2570
rect 57075 2550 57085 2570
rect 57045 2535 57085 2550
rect 57100 2570 57140 2585
rect 57100 2550 57110 2570
rect 57130 2550 57140 2570
rect 57100 2535 57140 2550
rect 57155 2570 57195 2585
rect 57155 2550 57165 2570
rect 57185 2550 57195 2570
rect 57155 2535 57195 2550
rect 57210 2570 57250 2585
rect 57210 2550 57220 2570
rect 57240 2550 57250 2570
rect 57210 2535 57250 2550
rect 56030 2165 56070 2180
rect 56030 2045 56040 2165
rect 56060 2045 56070 2165
rect 56030 2030 56070 2045
rect 56085 2165 56125 2180
rect 56085 2045 56095 2165
rect 56115 2045 56125 2165
rect 56085 2030 56125 2045
rect 56140 2165 56180 2180
rect 56140 2045 56150 2165
rect 56170 2045 56180 2165
rect 56140 2030 56180 2045
rect 56195 2165 56235 2180
rect 56195 2045 56205 2165
rect 56225 2045 56235 2165
rect 56195 2030 56235 2045
rect 56250 2165 56290 2180
rect 56250 2045 56260 2165
rect 56280 2045 56290 2165
rect 56250 2030 56290 2045
rect 56305 2165 56345 2180
rect 56305 2045 56315 2165
rect 56335 2045 56345 2165
rect 56305 2030 56345 2045
rect 56360 2165 56400 2180
rect 56360 2045 56370 2165
rect 56390 2045 56400 2165
rect 56360 2030 56400 2045
rect 56415 2165 56455 2180
rect 56415 2045 56425 2165
rect 56445 2045 56455 2165
rect 56415 2030 56455 2045
rect 56470 2165 56510 2180
rect 56470 2045 56480 2165
rect 56500 2045 56510 2165
rect 56470 2030 56510 2045
rect 56525 2165 56565 2180
rect 56525 2045 56535 2165
rect 56555 2045 56565 2165
rect 56525 2030 56565 2045
rect 56580 2165 56620 2180
rect 56580 2045 56590 2165
rect 56610 2045 56620 2165
rect 56580 2030 56620 2045
rect 56635 2165 56675 2180
rect 56635 2045 56645 2165
rect 56665 2045 56675 2165
rect 56635 2030 56675 2045
rect 56690 2165 56730 2180
rect 56690 2045 56700 2165
rect 56720 2045 56730 2165
rect 56690 2030 56730 2045
rect 57070 2165 57110 2180
rect 57070 2045 57080 2165
rect 57100 2045 57110 2165
rect 57070 2030 57110 2045
rect 57125 2165 57165 2180
rect 57125 2045 57135 2165
rect 57155 2045 57165 2165
rect 57125 2030 57165 2045
rect 57180 2165 57220 2180
rect 57180 2045 57190 2165
rect 57210 2045 57220 2165
rect 57180 2030 57220 2045
rect 57235 2165 57275 2180
rect 57235 2045 57245 2165
rect 57265 2045 57275 2165
rect 57235 2030 57275 2045
rect 57290 2165 57330 2180
rect 57290 2045 57300 2165
rect 57320 2045 57330 2165
rect 57290 2030 57330 2045
rect 57345 2165 57385 2180
rect 57345 2045 57355 2165
rect 57375 2045 57385 2165
rect 57345 2030 57385 2045
rect 57400 2165 57440 2180
rect 57400 2045 57410 2165
rect 57430 2045 57440 2165
rect 57400 2030 57440 2045
rect 57455 2165 57495 2180
rect 57455 2045 57465 2165
rect 57485 2045 57495 2165
rect 57455 2030 57495 2045
rect 57510 2165 57550 2180
rect 57510 2045 57520 2165
rect 57540 2045 57550 2165
rect 57510 2030 57550 2045
rect 57565 2165 57605 2180
rect 57565 2045 57575 2165
rect 57595 2045 57605 2165
rect 57565 2030 57605 2045
rect 57620 2165 57660 2180
rect 57620 2045 57630 2165
rect 57650 2045 57660 2165
rect 57620 2030 57660 2045
rect 57675 2165 57715 2180
rect 57675 2045 57685 2165
rect 57705 2045 57715 2165
rect 57675 2030 57715 2045
rect 57730 2165 57770 2180
rect 57730 2045 57740 2165
rect 57760 2045 57770 2165
rect 57730 2030 57770 2045
rect 54950 1845 54990 1860
rect 54950 1575 54960 1845
rect 54980 1575 54990 1845
rect 54950 1560 54990 1575
rect 55005 1845 55045 1860
rect 55005 1575 55015 1845
rect 55035 1575 55045 1845
rect 55005 1560 55045 1575
rect 55060 1845 55100 1860
rect 55060 1575 55070 1845
rect 55090 1575 55100 1845
rect 55060 1560 55100 1575
rect 55115 1845 55155 1860
rect 55115 1575 55125 1845
rect 55145 1575 55155 1845
rect 55115 1560 55155 1575
rect 55170 1845 55210 1860
rect 55170 1575 55180 1845
rect 55200 1575 55210 1845
rect 55170 1560 55210 1575
rect 55225 1845 55265 1860
rect 55225 1575 55235 1845
rect 55255 1575 55265 1845
rect 55225 1560 55265 1575
rect 55280 1845 55320 1860
rect 55280 1575 55290 1845
rect 55310 1575 55320 1845
rect 55280 1560 55320 1575
rect 55335 1845 55375 1860
rect 55335 1575 55345 1845
rect 55365 1575 55375 1845
rect 55335 1560 55375 1575
rect 55390 1845 55430 1860
rect 55390 1575 55400 1845
rect 55420 1575 55430 1845
rect 55390 1560 55430 1575
rect 55445 1845 55485 1860
rect 55445 1575 55455 1845
rect 55475 1575 55485 1845
rect 55445 1560 55485 1575
rect 55500 1845 55540 1860
rect 55500 1575 55510 1845
rect 55530 1575 55540 1845
rect 55500 1560 55540 1575
rect 55555 1845 55595 1860
rect 55555 1575 55565 1845
rect 55585 1575 55595 1845
rect 55555 1560 55595 1575
rect 55610 1845 55650 1860
rect 55610 1575 55620 1845
rect 55640 1575 55650 1845
rect 58150 1845 58190 1860
rect 55610 1560 55650 1575
rect 56030 1695 56070 1710
rect 56030 1575 56040 1695
rect 56060 1575 56070 1695
rect 56030 1560 56070 1575
rect 56085 1695 56125 1710
rect 56085 1575 56095 1695
rect 56115 1575 56125 1695
rect 56085 1560 56125 1575
rect 56140 1695 56180 1710
rect 56140 1575 56150 1695
rect 56170 1575 56180 1695
rect 56140 1560 56180 1575
rect 56195 1695 56235 1710
rect 56195 1575 56205 1695
rect 56225 1575 56235 1695
rect 56195 1560 56235 1575
rect 56250 1695 56290 1710
rect 56250 1575 56260 1695
rect 56280 1575 56290 1695
rect 56250 1560 56290 1575
rect 56305 1695 56345 1710
rect 56305 1575 56315 1695
rect 56335 1575 56345 1695
rect 56305 1560 56345 1575
rect 56360 1695 56400 1710
rect 56360 1575 56370 1695
rect 56390 1575 56400 1695
rect 56360 1560 56400 1575
rect 56415 1695 56455 1710
rect 56415 1575 56425 1695
rect 56445 1575 56455 1695
rect 56415 1560 56455 1575
rect 56470 1695 56510 1710
rect 56470 1575 56480 1695
rect 56500 1575 56510 1695
rect 56470 1560 56510 1575
rect 56525 1695 56565 1710
rect 56525 1575 56535 1695
rect 56555 1575 56565 1695
rect 56525 1560 56565 1575
rect 56580 1695 56620 1710
rect 56580 1575 56590 1695
rect 56610 1575 56620 1695
rect 56580 1560 56620 1575
rect 56635 1695 56675 1710
rect 56635 1575 56645 1695
rect 56665 1575 56675 1695
rect 56635 1560 56675 1575
rect 56690 1695 56730 1710
rect 56770 1695 56810 1710
rect 56690 1575 56700 1695
rect 56720 1575 56730 1695
rect 56770 1575 56780 1695
rect 56800 1575 56810 1695
rect 56690 1560 56730 1575
rect 56770 1560 56810 1575
rect 56825 1695 56865 1710
rect 56825 1575 56835 1695
rect 56855 1575 56865 1695
rect 56825 1560 56865 1575
rect 56880 1695 56920 1710
rect 56880 1575 56890 1695
rect 56910 1575 56920 1695
rect 56880 1560 56920 1575
rect 56935 1695 56975 1710
rect 56935 1575 56945 1695
rect 56965 1575 56975 1695
rect 56935 1560 56975 1575
rect 56990 1695 57030 1710
rect 57070 1695 57110 1710
rect 56990 1575 57000 1695
rect 57020 1575 57030 1695
rect 57070 1575 57080 1695
rect 57100 1575 57110 1695
rect 56990 1560 57030 1575
rect 57070 1560 57110 1575
rect 57125 1695 57165 1710
rect 57125 1575 57135 1695
rect 57155 1575 57165 1695
rect 57125 1560 57165 1575
rect 57180 1695 57220 1710
rect 57180 1575 57190 1695
rect 57210 1575 57220 1695
rect 57180 1560 57220 1575
rect 57235 1695 57275 1710
rect 57235 1575 57245 1695
rect 57265 1575 57275 1695
rect 57235 1560 57275 1575
rect 57290 1695 57330 1710
rect 57290 1575 57300 1695
rect 57320 1575 57330 1695
rect 57290 1560 57330 1575
rect 57345 1695 57385 1710
rect 57345 1575 57355 1695
rect 57375 1575 57385 1695
rect 57345 1560 57385 1575
rect 57400 1695 57440 1710
rect 57400 1575 57410 1695
rect 57430 1575 57440 1695
rect 57400 1560 57440 1575
rect 57455 1695 57495 1710
rect 57455 1575 57465 1695
rect 57485 1575 57495 1695
rect 57455 1560 57495 1575
rect 57510 1695 57550 1710
rect 57510 1575 57520 1695
rect 57540 1575 57550 1695
rect 57510 1560 57550 1575
rect 57565 1695 57605 1710
rect 57565 1575 57575 1695
rect 57595 1575 57605 1695
rect 57565 1560 57605 1575
rect 57620 1695 57660 1710
rect 57620 1575 57630 1695
rect 57650 1575 57660 1695
rect 57620 1560 57660 1575
rect 57675 1695 57715 1710
rect 57675 1575 57685 1695
rect 57705 1575 57715 1695
rect 57675 1560 57715 1575
rect 57730 1695 57770 1710
rect 57730 1575 57740 1695
rect 57760 1575 57770 1695
rect 57730 1560 57770 1575
rect 58150 1575 58160 1845
rect 58180 1575 58190 1845
rect 58150 1560 58190 1575
rect 58205 1845 58245 1860
rect 58205 1575 58215 1845
rect 58235 1575 58245 1845
rect 58205 1560 58245 1575
rect 58260 1845 58300 1860
rect 58260 1575 58270 1845
rect 58290 1575 58300 1845
rect 58260 1560 58300 1575
rect 58315 1845 58355 1860
rect 58315 1575 58325 1845
rect 58345 1575 58355 1845
rect 58315 1560 58355 1575
rect 58370 1845 58410 1860
rect 58370 1575 58380 1845
rect 58400 1575 58410 1845
rect 58370 1560 58410 1575
rect 58425 1845 58465 1860
rect 58425 1575 58435 1845
rect 58455 1575 58465 1845
rect 58425 1560 58465 1575
rect 58480 1845 58520 1860
rect 58480 1575 58490 1845
rect 58510 1575 58520 1845
rect 58480 1560 58520 1575
rect 58535 1845 58575 1860
rect 58535 1575 58545 1845
rect 58565 1575 58575 1845
rect 58535 1560 58575 1575
rect 58590 1845 58630 1860
rect 58590 1575 58600 1845
rect 58620 1575 58630 1845
rect 58590 1560 58630 1575
rect 58645 1845 58685 1860
rect 58645 1575 58655 1845
rect 58675 1575 58685 1845
rect 58645 1560 58685 1575
rect 58700 1845 58740 1860
rect 58700 1575 58710 1845
rect 58730 1575 58740 1845
rect 58700 1560 58740 1575
rect 58755 1845 58795 1860
rect 58755 1575 58765 1845
rect 58785 1575 58795 1845
rect 58755 1560 58795 1575
rect 58810 1845 58850 1860
rect 58810 1575 58820 1845
rect 58840 1575 58850 1845
rect 58810 1560 58850 1575
rect 54985 1155 55025 1170
rect 54985 485 54995 1155
rect 55015 485 55025 1155
rect 54985 470 55025 485
rect 55085 1155 55125 1170
rect 55085 485 55095 1155
rect 55115 485 55125 1155
rect 55085 470 55125 485
rect 55185 1155 55225 1170
rect 55185 485 55195 1155
rect 55215 485 55225 1155
rect 55185 470 55225 485
rect 55285 1155 55325 1170
rect 55285 485 55295 1155
rect 55315 485 55325 1155
rect 55285 470 55325 485
rect 55385 1155 55425 1170
rect 55385 485 55395 1155
rect 55415 485 55425 1155
rect 55385 470 55425 485
rect 55485 1155 55525 1170
rect 55485 485 55495 1155
rect 55515 485 55525 1155
rect 55485 470 55525 485
rect 55585 1155 55625 1170
rect 55585 485 55595 1155
rect 55615 485 55625 1155
rect 56220 1145 56260 1160
rect 56220 925 56230 1145
rect 56250 925 56260 1145
rect 56220 910 56260 925
rect 56275 1145 56315 1160
rect 56275 925 56285 1145
rect 56305 925 56315 1145
rect 56275 910 56315 925
rect 56330 1145 56370 1160
rect 56330 925 56340 1145
rect 56360 925 56370 1145
rect 56330 910 56370 925
rect 56385 1145 56425 1160
rect 56385 925 56395 1145
rect 56415 925 56425 1145
rect 56385 910 56425 925
rect 56440 1145 56480 1160
rect 56440 925 56450 1145
rect 56470 925 56480 1145
rect 56440 910 56480 925
rect 56495 1145 56535 1160
rect 56495 925 56505 1145
rect 56525 925 56535 1145
rect 56495 910 56535 925
rect 56550 1145 56590 1160
rect 56550 925 56560 1145
rect 56580 925 56590 1145
rect 56550 910 56590 925
rect 56605 1145 56645 1160
rect 56605 925 56615 1145
rect 56635 925 56645 1145
rect 56605 910 56645 925
rect 56660 1145 56700 1160
rect 56660 925 56670 1145
rect 56690 925 56700 1145
rect 56660 910 56700 925
rect 56715 1145 56755 1160
rect 56715 925 56725 1145
rect 56745 925 56755 1145
rect 56715 910 56755 925
rect 56770 1145 56810 1160
rect 56770 925 56780 1145
rect 56800 925 56810 1145
rect 56770 910 56810 925
rect 56825 1145 56865 1160
rect 56825 925 56835 1145
rect 56855 925 56865 1145
rect 56825 910 56865 925
rect 56880 1145 56920 1160
rect 56880 925 56890 1145
rect 56910 925 56920 1145
rect 56880 910 56920 925
rect 56935 1145 56975 1160
rect 56935 925 56945 1145
rect 56965 925 56975 1145
rect 56935 910 56975 925
rect 56990 1145 57030 1160
rect 56990 925 57000 1145
rect 57020 925 57030 1145
rect 56990 910 57030 925
rect 57045 1145 57085 1160
rect 57045 925 57055 1145
rect 57075 925 57085 1145
rect 57045 910 57085 925
rect 57100 1145 57140 1160
rect 57100 925 57110 1145
rect 57130 925 57140 1145
rect 57100 910 57140 925
rect 57155 1145 57195 1160
rect 57155 925 57165 1145
rect 57185 925 57195 1145
rect 57155 910 57195 925
rect 57210 1145 57250 1160
rect 57210 925 57220 1145
rect 57240 925 57250 1145
rect 57210 910 57250 925
rect 57265 1145 57305 1160
rect 57265 925 57275 1145
rect 57295 925 57305 1145
rect 57265 910 57305 925
rect 57320 1145 57360 1160
rect 57320 925 57330 1145
rect 57350 925 57360 1145
rect 57320 910 57360 925
rect 57375 1145 57415 1160
rect 57375 925 57385 1145
rect 57405 925 57415 1145
rect 57375 910 57415 925
rect 57430 1145 57470 1160
rect 57430 925 57440 1145
rect 57460 925 57470 1145
rect 57430 910 57470 925
rect 57485 1145 57525 1160
rect 57485 925 57495 1145
rect 57515 925 57525 1145
rect 57485 910 57525 925
rect 58180 1155 58220 1170
rect 56430 680 56470 695
rect 56430 560 56440 680
rect 56460 560 56470 680
rect 56430 545 56470 560
rect 56485 680 56525 695
rect 56485 560 56495 680
rect 56515 560 56525 680
rect 56485 545 56525 560
rect 56540 680 56580 695
rect 56540 560 56550 680
rect 56570 560 56580 680
rect 56540 545 56580 560
rect 56595 680 56635 695
rect 56595 560 56605 680
rect 56625 560 56635 680
rect 56595 545 56635 560
rect 56650 680 56690 695
rect 56650 560 56660 680
rect 56680 560 56690 680
rect 56650 545 56690 560
rect 56705 680 56745 695
rect 56705 560 56715 680
rect 56735 560 56745 680
rect 56705 545 56745 560
rect 56760 680 56800 695
rect 56760 560 56770 680
rect 56790 560 56800 680
rect 56760 545 56800 560
rect 56870 680 56910 695
rect 56870 560 56880 680
rect 56900 560 56910 680
rect 56870 545 56910 560
rect 57210 680 57250 695
rect 57210 560 57220 680
rect 57240 560 57250 680
rect 57210 545 57250 560
rect 55585 470 55625 485
rect 58180 485 58190 1155
rect 58210 485 58220 1155
rect 58180 470 58220 485
rect 58280 1155 58320 1170
rect 58280 485 58290 1155
rect 58310 485 58320 1155
rect 58280 470 58320 485
rect 58380 1155 58420 1170
rect 58380 485 58390 1155
rect 58410 485 58420 1155
rect 58380 470 58420 485
rect 58480 1155 58520 1170
rect 58480 485 58490 1155
rect 58510 485 58520 1155
rect 58480 470 58520 485
rect 58580 1155 58620 1170
rect 58580 485 58590 1155
rect 58610 485 58620 1155
rect 58580 470 58620 485
rect 58680 1155 58720 1170
rect 58680 485 58690 1155
rect 58710 485 58720 1155
rect 58680 470 58720 485
rect 58780 1155 58820 1170
rect 58780 485 58790 1155
rect 58810 485 58820 1155
rect 58780 470 58820 485
<< pdiff >>
rect 56085 4695 56125 4710
rect 56085 4375 56095 4695
rect 56115 4375 56125 4695
rect 56085 4360 56125 4375
rect 56145 4695 56185 4710
rect 56145 4375 56155 4695
rect 56175 4375 56185 4695
rect 56145 4360 56185 4375
rect 56205 4695 56245 4710
rect 56205 4375 56215 4695
rect 56235 4375 56245 4695
rect 56205 4360 56245 4375
rect 56265 4695 56305 4710
rect 56265 4375 56275 4695
rect 56295 4375 56305 4695
rect 57025 4695 57065 4710
rect 56265 4360 56305 4375
rect 56555 4525 56595 4540
rect 56555 4375 56565 4525
rect 56585 4375 56595 4525
rect 56555 4360 56595 4375
rect 56615 4525 56655 4540
rect 56615 4375 56625 4525
rect 56645 4375 56655 4525
rect 56615 4360 56655 4375
rect 56675 4525 56715 4540
rect 56675 4375 56685 4525
rect 56705 4375 56715 4525
rect 56675 4360 56715 4375
rect 56735 4525 56775 4540
rect 56735 4375 56745 4525
rect 56765 4375 56775 4525
rect 56735 4360 56775 4375
rect 57025 4375 57035 4695
rect 57055 4375 57065 4695
rect 57025 4360 57065 4375
rect 57085 4695 57125 4710
rect 57085 4375 57095 4695
rect 57115 4375 57125 4695
rect 57085 4360 57125 4375
rect 57145 4695 57185 4710
rect 57145 4375 57155 4695
rect 57175 4375 57185 4695
rect 57145 4360 57185 4375
rect 57205 4695 57245 4710
rect 57205 4375 57215 4695
rect 57235 4375 57245 4695
rect 57205 4360 57245 4375
rect 57495 4695 57535 4710
rect 57495 4375 57505 4695
rect 57525 4375 57535 4695
rect 57495 4360 57535 4375
rect 57555 4695 57595 4710
rect 57555 4375 57565 4695
rect 57585 4375 57595 4695
rect 57555 4360 57595 4375
rect 57615 4695 57655 4710
rect 57615 4375 57625 4695
rect 57645 4375 57655 4695
rect 57615 4360 57655 4375
rect 57675 4695 57715 4710
rect 57675 4375 57685 4695
rect 57705 4375 57715 4695
rect 57675 4360 57715 4375
rect 54925 4025 54965 4040
rect 54925 3705 54935 4025
rect 54955 3705 54965 4025
rect 54925 3690 54965 3705
rect 54985 4025 55025 4040
rect 54985 3705 54995 4025
rect 55015 3705 55025 4025
rect 54985 3690 55025 3705
rect 55045 4025 55085 4040
rect 55045 3705 55055 4025
rect 55075 3705 55085 4025
rect 55045 3690 55085 3705
rect 55105 4025 55145 4040
rect 55105 3705 55115 4025
rect 55135 3705 55145 4025
rect 55105 3690 55145 3705
rect 55165 4025 55205 4040
rect 55165 3705 55175 4025
rect 55195 3705 55205 4025
rect 55165 3690 55205 3705
rect 55225 4025 55265 4040
rect 55225 3705 55235 4025
rect 55255 3705 55265 4025
rect 55225 3690 55265 3705
rect 55285 4025 55325 4040
rect 55285 3705 55295 4025
rect 55315 3705 55325 4025
rect 55285 3690 55325 3705
rect 55345 4025 55385 4040
rect 55345 3705 55355 4025
rect 55375 3705 55385 4025
rect 55345 3690 55385 3705
rect 55405 4025 55445 4040
rect 55405 3705 55415 4025
rect 55435 3705 55445 4025
rect 55405 3690 55445 3705
rect 55465 4025 55505 4040
rect 55465 3705 55475 4025
rect 55495 3705 55505 4025
rect 55465 3690 55505 3705
rect 55525 4025 55565 4040
rect 55525 3705 55535 4025
rect 55555 3705 55565 4025
rect 55525 3690 55565 3705
rect 55585 4025 55625 4040
rect 55585 3705 55595 4025
rect 55615 3705 55625 4025
rect 55585 3690 55625 3705
rect 55645 4025 55685 4040
rect 55645 3705 55655 4025
rect 55675 3705 55685 4025
rect 55645 3690 55685 3705
rect 56005 4025 56045 4040
rect 56005 3705 56015 4025
rect 56035 3705 56045 4025
rect 56005 3690 56045 3705
rect 56065 4025 56105 4040
rect 56065 3705 56075 4025
rect 56095 3705 56105 4025
rect 56065 3690 56105 3705
rect 56125 4025 56165 4040
rect 56125 3705 56135 4025
rect 56155 3705 56165 4025
rect 56125 3690 56165 3705
rect 56185 4025 56225 4040
rect 56185 3705 56195 4025
rect 56215 3705 56225 4025
rect 56185 3690 56225 3705
rect 56245 4025 56285 4040
rect 56245 3705 56255 4025
rect 56275 3705 56285 4025
rect 56245 3690 56285 3705
rect 56305 4025 56345 4040
rect 56305 3705 56315 4025
rect 56335 3705 56345 4025
rect 56305 3690 56345 3705
rect 56365 4025 56405 4040
rect 56365 3705 56375 4025
rect 56395 3705 56405 4025
rect 56365 3690 56405 3705
rect 56425 4025 56465 4040
rect 56425 3705 56435 4025
rect 56455 3705 56465 4025
rect 56425 3690 56465 3705
rect 56485 4025 56525 4040
rect 56485 3705 56495 4025
rect 56515 3705 56525 4025
rect 56485 3690 56525 3705
rect 56545 4025 56585 4040
rect 56545 3705 56555 4025
rect 56575 3705 56585 4025
rect 56545 3690 56585 3705
rect 56605 4025 56645 4040
rect 56605 3705 56615 4025
rect 56635 3705 56645 4025
rect 56605 3690 56645 3705
rect 56665 4025 56705 4040
rect 56665 3705 56675 4025
rect 56695 3705 56705 4025
rect 56665 3690 56705 3705
rect 56725 4025 56765 4040
rect 56725 3705 56735 4025
rect 56755 3705 56765 4025
rect 56725 3690 56765 3705
rect 57035 4025 57075 4040
rect 57035 3705 57045 4025
rect 57065 3705 57075 4025
rect 57035 3690 57075 3705
rect 57095 4025 57135 4040
rect 57095 3705 57105 4025
rect 57125 3705 57135 4025
rect 57095 3690 57135 3705
rect 57155 4025 57195 4040
rect 57155 3705 57165 4025
rect 57185 3705 57195 4025
rect 57155 3690 57195 3705
rect 57215 4025 57255 4040
rect 57215 3705 57225 4025
rect 57245 3705 57255 4025
rect 57215 3690 57255 3705
rect 57275 4025 57315 4040
rect 57275 3705 57285 4025
rect 57305 3705 57315 4025
rect 57275 3690 57315 3705
rect 57335 4025 57375 4040
rect 57335 3705 57345 4025
rect 57365 3705 57375 4025
rect 57335 3690 57375 3705
rect 57395 4025 57435 4040
rect 57395 3705 57405 4025
rect 57425 3705 57435 4025
rect 57395 3690 57435 3705
rect 57455 4025 57495 4040
rect 57455 3705 57465 4025
rect 57485 3705 57495 4025
rect 57455 3690 57495 3705
rect 57515 4025 57555 4040
rect 57515 3705 57525 4025
rect 57545 3705 57555 4025
rect 57515 3690 57555 3705
rect 57575 4025 57615 4040
rect 57575 3705 57585 4025
rect 57605 3705 57615 4025
rect 57575 3690 57615 3705
rect 57635 4025 57675 4040
rect 57635 3705 57645 4025
rect 57665 3705 57675 4025
rect 57635 3690 57675 3705
rect 57695 4025 57735 4040
rect 57695 3705 57705 4025
rect 57725 3705 57735 4025
rect 57695 3690 57735 3705
rect 57755 4025 57795 4040
rect 57755 3705 57765 4025
rect 57785 3705 57795 4025
rect 57755 3690 57795 3705
rect 58120 4025 58160 4040
rect 58120 3705 58130 4025
rect 58150 3705 58160 4025
rect 58120 3690 58160 3705
rect 58180 4025 58220 4040
rect 58180 3705 58190 4025
rect 58210 3705 58220 4025
rect 58180 3690 58220 3705
rect 58240 4025 58280 4040
rect 58240 3705 58250 4025
rect 58270 3705 58280 4025
rect 58240 3690 58280 3705
rect 58300 4025 58340 4040
rect 58300 3705 58310 4025
rect 58330 3705 58340 4025
rect 58300 3690 58340 3705
rect 58360 4025 58400 4040
rect 58360 3705 58370 4025
rect 58390 3705 58400 4025
rect 58360 3690 58400 3705
rect 58420 4025 58460 4040
rect 58420 3705 58430 4025
rect 58450 3705 58460 4025
rect 58420 3690 58460 3705
rect 58480 4025 58520 4040
rect 58480 3705 58490 4025
rect 58510 3705 58520 4025
rect 58480 3690 58520 3705
rect 58540 4025 58580 4040
rect 58540 3705 58550 4025
rect 58570 3705 58580 4025
rect 58540 3690 58580 3705
rect 58600 4025 58640 4040
rect 58600 3705 58610 4025
rect 58630 3705 58640 4025
rect 58600 3690 58640 3705
rect 58660 4025 58700 4040
rect 58660 3705 58670 4025
rect 58690 3705 58700 4025
rect 58660 3690 58700 3705
rect 58720 4025 58760 4040
rect 58720 3705 58730 4025
rect 58750 3705 58760 4025
rect 58720 3690 58760 3705
rect 58780 4025 58820 4040
rect 58780 3705 58790 4025
rect 58810 3705 58820 4025
rect 58780 3690 58820 3705
rect 58840 4025 58880 4040
rect 58840 3705 58850 4025
rect 58870 3705 58880 4025
rect 58840 3690 58880 3705
rect 54950 3335 54990 3350
rect 54950 2765 54960 3335
rect 54980 2765 54990 3335
rect 54950 2750 54990 2765
rect 55005 3335 55045 3350
rect 55005 2765 55015 3335
rect 55035 2765 55045 3335
rect 55005 2750 55045 2765
rect 55060 3335 55100 3350
rect 55060 2765 55070 3335
rect 55090 2765 55100 3335
rect 55060 2750 55100 2765
rect 55115 3335 55155 3350
rect 55115 2765 55125 3335
rect 55145 2765 55155 3335
rect 55115 2750 55155 2765
rect 55170 3335 55210 3350
rect 55170 2765 55180 3335
rect 55200 2765 55210 3335
rect 55170 2750 55210 2765
rect 55225 3335 55265 3350
rect 55225 2765 55235 3335
rect 55255 2765 55265 3335
rect 55225 2750 55265 2765
rect 55280 3335 55320 3350
rect 55280 2765 55290 3335
rect 55310 2765 55320 3335
rect 55280 2750 55320 2765
rect 55335 3335 55375 3350
rect 55335 2765 55345 3335
rect 55365 2765 55375 3335
rect 55335 2750 55375 2765
rect 55390 3335 55430 3350
rect 55390 2765 55400 3335
rect 55420 2765 55430 3335
rect 55390 2750 55430 2765
rect 55445 3335 55485 3350
rect 55445 2765 55455 3335
rect 55475 2765 55485 3335
rect 55445 2750 55485 2765
rect 55500 3335 55540 3350
rect 55500 2765 55510 3335
rect 55530 2765 55540 3335
rect 55500 2750 55540 2765
rect 55555 3335 55595 3350
rect 55555 2765 55565 3335
rect 55585 2765 55595 3335
rect 55555 2750 55595 2765
rect 55610 3335 55650 3350
rect 55610 2765 55620 3335
rect 55640 2765 55650 3335
rect 56275 3340 56315 3355
rect 56275 3320 56285 3340
rect 56305 3320 56315 3340
rect 56275 3305 56315 3320
rect 56330 3340 56370 3355
rect 56330 3320 56340 3340
rect 56360 3320 56370 3340
rect 56330 3305 56370 3320
rect 56385 3340 56425 3355
rect 56385 3320 56395 3340
rect 56415 3320 56425 3340
rect 56385 3305 56425 3320
rect 56440 3340 56480 3355
rect 56440 3320 56450 3340
rect 56470 3320 56480 3340
rect 56440 3305 56480 3320
rect 56495 3340 56535 3355
rect 56495 3320 56505 3340
rect 56525 3320 56535 3340
rect 56495 3305 56535 3320
rect 56550 3340 56590 3355
rect 56550 3320 56560 3340
rect 56580 3320 56590 3340
rect 56550 3305 56590 3320
rect 56605 3340 56645 3355
rect 56605 3320 56615 3340
rect 56635 3320 56645 3340
rect 56605 3305 56645 3320
rect 56660 3340 56700 3355
rect 56660 3320 56670 3340
rect 56690 3320 56700 3340
rect 56660 3305 56700 3320
rect 56715 3340 56755 3355
rect 56715 3320 56725 3340
rect 56745 3320 56755 3340
rect 56715 3305 56755 3320
rect 56770 3340 56810 3355
rect 56770 3320 56780 3340
rect 56800 3320 56810 3340
rect 56770 3305 56810 3320
rect 56825 3340 56865 3355
rect 56825 3320 56835 3340
rect 56855 3320 56865 3340
rect 56825 3305 56865 3320
rect 56880 3340 56920 3355
rect 56880 3320 56890 3340
rect 56910 3320 56920 3340
rect 56880 3305 56920 3320
rect 56935 3340 56975 3355
rect 56935 3320 56945 3340
rect 56965 3320 56975 3340
rect 56935 3305 56975 3320
rect 56990 3340 57030 3355
rect 56990 3320 57000 3340
rect 57020 3320 57030 3340
rect 56990 3305 57030 3320
rect 57045 3340 57085 3355
rect 57045 3320 57055 3340
rect 57075 3320 57085 3340
rect 57045 3305 57085 3320
rect 57100 3340 57140 3355
rect 57100 3320 57110 3340
rect 57130 3320 57140 3340
rect 57100 3305 57140 3320
rect 57155 3340 57195 3355
rect 57155 3320 57165 3340
rect 57185 3320 57195 3340
rect 57155 3305 57195 3320
rect 57210 3340 57250 3355
rect 57210 3320 57220 3340
rect 57240 3320 57250 3340
rect 57210 3305 57250 3320
rect 57265 3340 57305 3355
rect 57265 3320 57275 3340
rect 57295 3320 57305 3340
rect 57265 3305 57305 3320
rect 57320 3340 57360 3355
rect 57320 3320 57330 3340
rect 57350 3320 57360 3340
rect 57320 3305 57360 3320
rect 57375 3340 57415 3355
rect 57375 3320 57385 3340
rect 57405 3320 57415 3340
rect 57375 3305 57415 3320
rect 57430 3340 57470 3355
rect 57430 3320 57440 3340
rect 57460 3320 57470 3340
rect 57430 3305 57470 3320
rect 57485 3340 57525 3355
rect 57485 3320 57495 3340
rect 57515 3320 57525 3340
rect 57485 3305 57525 3320
rect 58150 3335 58190 3350
rect 56030 2980 56070 2995
rect 56030 2960 56040 2980
rect 56060 2960 56070 2980
rect 56030 2945 56070 2960
rect 56085 2980 56125 2995
rect 56085 2960 56095 2980
rect 56115 2960 56125 2980
rect 56085 2945 56125 2960
rect 56140 2980 56180 2995
rect 56140 2960 56150 2980
rect 56170 2960 56180 2980
rect 56140 2945 56180 2960
rect 56195 2980 56235 2995
rect 56195 2960 56205 2980
rect 56225 2960 56235 2980
rect 56195 2945 56235 2960
rect 56250 2980 56290 2995
rect 56250 2960 56260 2980
rect 56280 2960 56290 2980
rect 56250 2945 56290 2960
rect 56305 2980 56345 2995
rect 56305 2960 56315 2980
rect 56335 2960 56345 2980
rect 56305 2945 56345 2960
rect 56360 2980 56400 2995
rect 56360 2960 56370 2980
rect 56390 2960 56400 2980
rect 56360 2945 56400 2960
rect 56415 2980 56455 2995
rect 56415 2960 56425 2980
rect 56445 2960 56455 2980
rect 56415 2945 56455 2960
rect 56470 2980 56510 2995
rect 56470 2960 56480 2980
rect 56500 2960 56510 2980
rect 56470 2945 56510 2960
rect 56525 2980 56565 2995
rect 56525 2960 56535 2980
rect 56555 2960 56565 2980
rect 56525 2945 56565 2960
rect 56580 2980 56620 2995
rect 56580 2960 56590 2980
rect 56610 2960 56620 2980
rect 56580 2945 56620 2960
rect 56635 2980 56675 2995
rect 56635 2960 56645 2980
rect 56665 2960 56675 2980
rect 56635 2945 56675 2960
rect 56690 2980 56730 2995
rect 56690 2960 56700 2980
rect 56720 2960 56730 2980
rect 56690 2945 56730 2960
rect 57070 2980 57110 2995
rect 57070 2960 57080 2980
rect 57100 2960 57110 2980
rect 57070 2945 57110 2960
rect 57125 2980 57165 2995
rect 57125 2960 57135 2980
rect 57155 2960 57165 2980
rect 57125 2945 57165 2960
rect 57180 2980 57220 2995
rect 57180 2960 57190 2980
rect 57210 2960 57220 2980
rect 57180 2945 57220 2960
rect 57235 2980 57275 2995
rect 57235 2960 57245 2980
rect 57265 2960 57275 2980
rect 57235 2945 57275 2960
rect 57290 2980 57330 2995
rect 57290 2960 57300 2980
rect 57320 2960 57330 2980
rect 57290 2945 57330 2960
rect 57345 2980 57385 2995
rect 57345 2960 57355 2980
rect 57375 2960 57385 2980
rect 57345 2945 57385 2960
rect 57400 2980 57440 2995
rect 57400 2960 57410 2980
rect 57430 2960 57440 2980
rect 57400 2945 57440 2960
rect 57455 2980 57495 2995
rect 57455 2960 57465 2980
rect 57485 2960 57495 2980
rect 57455 2945 57495 2960
rect 57510 2980 57550 2995
rect 57510 2960 57520 2980
rect 57540 2960 57550 2980
rect 57510 2945 57550 2960
rect 57565 2980 57605 2995
rect 57565 2960 57575 2980
rect 57595 2960 57605 2980
rect 57565 2945 57605 2960
rect 57620 2980 57660 2995
rect 57620 2960 57630 2980
rect 57650 2960 57660 2980
rect 57620 2945 57660 2960
rect 57675 2980 57715 2995
rect 57675 2960 57685 2980
rect 57705 2960 57715 2980
rect 57675 2945 57715 2960
rect 57730 2980 57770 2995
rect 57730 2960 57740 2980
rect 57760 2960 57770 2980
rect 57730 2945 57770 2960
rect 55610 2750 55650 2765
rect 58150 2765 58160 3335
rect 58180 2765 58190 3335
rect 58150 2750 58190 2765
rect 58205 3335 58245 3350
rect 58205 2765 58215 3335
rect 58235 2765 58245 3335
rect 58205 2750 58245 2765
rect 58260 3335 58300 3350
rect 58260 2765 58270 3335
rect 58290 2765 58300 3335
rect 58260 2750 58300 2765
rect 58315 3335 58355 3350
rect 58315 2765 58325 3335
rect 58345 2765 58355 3335
rect 58315 2750 58355 2765
rect 58370 3335 58410 3350
rect 58370 2765 58380 3335
rect 58400 2765 58410 3335
rect 58370 2750 58410 2765
rect 58425 3335 58465 3350
rect 58425 2765 58435 3335
rect 58455 2765 58465 3335
rect 58425 2750 58465 2765
rect 58480 3335 58520 3350
rect 58480 2765 58490 3335
rect 58510 2765 58520 3335
rect 58480 2750 58520 2765
rect 58535 3335 58575 3350
rect 58535 2765 58545 3335
rect 58565 2765 58575 3335
rect 58535 2750 58575 2765
rect 58590 3335 58630 3350
rect 58590 2765 58600 3335
rect 58620 2765 58630 3335
rect 58590 2750 58630 2765
rect 58645 3335 58685 3350
rect 58645 2765 58655 3335
rect 58675 2765 58685 3335
rect 58645 2750 58685 2765
rect 58700 3335 58740 3350
rect 58700 2765 58710 3335
rect 58730 2765 58740 3335
rect 58700 2750 58740 2765
rect 58755 3335 58795 3350
rect 58755 2765 58765 3335
rect 58785 2765 58795 3335
rect 58755 2750 58795 2765
rect 58810 3335 58850 3350
rect 58810 2765 58820 3335
rect 58840 2765 58850 3335
rect 58810 2750 58850 2765
rect 54950 2405 54990 2420
rect 54950 2235 54960 2405
rect 54980 2235 54990 2405
rect 54950 2220 54990 2235
rect 55005 2405 55045 2420
rect 55005 2235 55015 2405
rect 55035 2235 55045 2405
rect 55005 2220 55045 2235
rect 55060 2405 55100 2420
rect 55060 2235 55070 2405
rect 55090 2235 55100 2405
rect 55060 2220 55100 2235
rect 55115 2405 55155 2420
rect 55115 2235 55125 2405
rect 55145 2235 55155 2405
rect 55115 2220 55155 2235
rect 55170 2405 55210 2420
rect 55170 2235 55180 2405
rect 55200 2235 55210 2405
rect 55170 2220 55210 2235
rect 55225 2405 55265 2420
rect 55225 2235 55235 2405
rect 55255 2235 55265 2405
rect 55225 2220 55265 2235
rect 55280 2405 55320 2420
rect 55280 2235 55290 2405
rect 55310 2235 55320 2405
rect 55280 2220 55320 2235
rect 55335 2405 55375 2420
rect 55335 2235 55345 2405
rect 55365 2235 55375 2405
rect 55335 2220 55375 2235
rect 55390 2405 55430 2420
rect 55390 2235 55400 2405
rect 55420 2235 55430 2405
rect 55390 2220 55430 2235
rect 55445 2405 55485 2420
rect 55445 2235 55455 2405
rect 55475 2235 55485 2405
rect 55445 2220 55485 2235
rect 55500 2405 55540 2420
rect 55500 2235 55510 2405
rect 55530 2235 55540 2405
rect 55500 2220 55540 2235
rect 55555 2405 55595 2420
rect 55555 2235 55565 2405
rect 55585 2235 55595 2405
rect 55555 2220 55595 2235
rect 55610 2405 55650 2420
rect 55610 2235 55620 2405
rect 55640 2235 55650 2405
rect 58150 2405 58190 2420
rect 55610 2220 55650 2235
rect 58150 2235 58160 2405
rect 58180 2235 58190 2405
rect 58150 2220 58190 2235
rect 58205 2405 58245 2420
rect 58205 2235 58215 2405
rect 58235 2235 58245 2405
rect 58205 2220 58245 2235
rect 58260 2405 58300 2420
rect 58260 2235 58270 2405
rect 58290 2235 58300 2405
rect 58260 2220 58300 2235
rect 58315 2405 58355 2420
rect 58315 2235 58325 2405
rect 58345 2235 58355 2405
rect 58315 2220 58355 2235
rect 58370 2405 58410 2420
rect 58370 2235 58380 2405
rect 58400 2235 58410 2405
rect 58370 2220 58410 2235
rect 58425 2405 58465 2420
rect 58425 2235 58435 2405
rect 58455 2235 58465 2405
rect 58425 2220 58465 2235
rect 58480 2405 58520 2420
rect 58480 2235 58490 2405
rect 58510 2235 58520 2405
rect 58480 2220 58520 2235
rect 58535 2405 58575 2420
rect 58535 2235 58545 2405
rect 58565 2235 58575 2405
rect 58535 2220 58575 2235
rect 58590 2405 58630 2420
rect 58590 2235 58600 2405
rect 58620 2235 58630 2405
rect 58590 2220 58630 2235
rect 58645 2405 58685 2420
rect 58645 2235 58655 2405
rect 58675 2235 58685 2405
rect 58645 2220 58685 2235
rect 58700 2405 58740 2420
rect 58700 2235 58710 2405
rect 58730 2235 58740 2405
rect 58700 2220 58740 2235
rect 58755 2405 58795 2420
rect 58755 2235 58765 2405
rect 58785 2235 58795 2405
rect 58755 2220 58795 2235
rect 58810 2405 58850 2420
rect 58810 2235 58820 2405
rect 58840 2235 58850 2405
rect 58810 2220 58850 2235
<< ndiffc >>
rect 56560 2550 56580 2570
rect 56615 2550 56635 2570
rect 56670 2550 56690 2570
rect 56725 2550 56745 2570
rect 56780 2550 56800 2570
rect 56835 2550 56855 2570
rect 56890 2550 56910 2570
rect 56945 2550 56965 2570
rect 57000 2550 57020 2570
rect 57055 2550 57075 2570
rect 57110 2550 57130 2570
rect 57165 2550 57185 2570
rect 57220 2550 57240 2570
rect 56040 2045 56060 2165
rect 56095 2045 56115 2165
rect 56150 2045 56170 2165
rect 56205 2045 56225 2165
rect 56260 2045 56280 2165
rect 56315 2045 56335 2165
rect 56370 2045 56390 2165
rect 56425 2045 56445 2165
rect 56480 2045 56500 2165
rect 56535 2045 56555 2165
rect 56590 2045 56610 2165
rect 56645 2045 56665 2165
rect 56700 2045 56720 2165
rect 57080 2045 57100 2165
rect 57135 2045 57155 2165
rect 57190 2045 57210 2165
rect 57245 2045 57265 2165
rect 57300 2045 57320 2165
rect 57355 2045 57375 2165
rect 57410 2045 57430 2165
rect 57465 2045 57485 2165
rect 57520 2045 57540 2165
rect 57575 2045 57595 2165
rect 57630 2045 57650 2165
rect 57685 2045 57705 2165
rect 57740 2045 57760 2165
rect 54960 1575 54980 1845
rect 55015 1575 55035 1845
rect 55070 1575 55090 1845
rect 55125 1575 55145 1845
rect 55180 1575 55200 1845
rect 55235 1575 55255 1845
rect 55290 1575 55310 1845
rect 55345 1575 55365 1845
rect 55400 1575 55420 1845
rect 55455 1575 55475 1845
rect 55510 1575 55530 1845
rect 55565 1575 55585 1845
rect 55620 1575 55640 1845
rect 56040 1575 56060 1695
rect 56095 1575 56115 1695
rect 56150 1575 56170 1695
rect 56205 1575 56225 1695
rect 56260 1575 56280 1695
rect 56315 1575 56335 1695
rect 56370 1575 56390 1695
rect 56425 1575 56445 1695
rect 56480 1575 56500 1695
rect 56535 1575 56555 1695
rect 56590 1575 56610 1695
rect 56645 1575 56665 1695
rect 56700 1575 56720 1695
rect 56780 1575 56800 1695
rect 56835 1575 56855 1695
rect 56890 1575 56910 1695
rect 56945 1575 56965 1695
rect 57000 1575 57020 1695
rect 57080 1575 57100 1695
rect 57135 1575 57155 1695
rect 57190 1575 57210 1695
rect 57245 1575 57265 1695
rect 57300 1575 57320 1695
rect 57355 1575 57375 1695
rect 57410 1575 57430 1695
rect 57465 1575 57485 1695
rect 57520 1575 57540 1695
rect 57575 1575 57595 1695
rect 57630 1575 57650 1695
rect 57685 1575 57705 1695
rect 57740 1575 57760 1695
rect 58160 1575 58180 1845
rect 58215 1575 58235 1845
rect 58270 1575 58290 1845
rect 58325 1575 58345 1845
rect 58380 1575 58400 1845
rect 58435 1575 58455 1845
rect 58490 1575 58510 1845
rect 58545 1575 58565 1845
rect 58600 1575 58620 1845
rect 58655 1575 58675 1845
rect 58710 1575 58730 1845
rect 58765 1575 58785 1845
rect 58820 1575 58840 1845
rect 54995 485 55015 1155
rect 55095 485 55115 1155
rect 55195 485 55215 1155
rect 55295 485 55315 1155
rect 55395 485 55415 1155
rect 55495 485 55515 1155
rect 55595 485 55615 1155
rect 56230 925 56250 1145
rect 56285 925 56305 1145
rect 56340 925 56360 1145
rect 56395 925 56415 1145
rect 56450 925 56470 1145
rect 56505 925 56525 1145
rect 56560 925 56580 1145
rect 56615 925 56635 1145
rect 56670 925 56690 1145
rect 56725 925 56745 1145
rect 56780 925 56800 1145
rect 56835 925 56855 1145
rect 56890 925 56910 1145
rect 56945 925 56965 1145
rect 57000 925 57020 1145
rect 57055 925 57075 1145
rect 57110 925 57130 1145
rect 57165 925 57185 1145
rect 57220 925 57240 1145
rect 57275 925 57295 1145
rect 57330 925 57350 1145
rect 57385 925 57405 1145
rect 57440 925 57460 1145
rect 57495 925 57515 1145
rect 56440 560 56460 680
rect 56495 560 56515 680
rect 56550 560 56570 680
rect 56605 560 56625 680
rect 56660 560 56680 680
rect 56715 560 56735 680
rect 56770 560 56790 680
rect 56880 560 56900 680
rect 57220 560 57240 680
rect 58190 485 58210 1155
rect 58290 485 58310 1155
rect 58390 485 58410 1155
rect 58490 485 58510 1155
rect 58590 485 58610 1155
rect 58690 485 58710 1155
rect 58790 485 58810 1155
<< pdiffc >>
rect 56095 4375 56115 4695
rect 56155 4375 56175 4695
rect 56215 4375 56235 4695
rect 56275 4375 56295 4695
rect 56565 4375 56585 4525
rect 56625 4375 56645 4525
rect 56685 4375 56705 4525
rect 56745 4375 56765 4525
rect 57035 4375 57055 4695
rect 57095 4375 57115 4695
rect 57155 4375 57175 4695
rect 57215 4375 57235 4695
rect 57505 4375 57525 4695
rect 57565 4375 57585 4695
rect 57625 4375 57645 4695
rect 57685 4375 57705 4695
rect 54935 3705 54955 4025
rect 54995 3705 55015 4025
rect 55055 3705 55075 4025
rect 55115 3705 55135 4025
rect 55175 3705 55195 4025
rect 55235 3705 55255 4025
rect 55295 3705 55315 4025
rect 55355 3705 55375 4025
rect 55415 3705 55435 4025
rect 55475 3705 55495 4025
rect 55535 3705 55555 4025
rect 55595 3705 55615 4025
rect 55655 3705 55675 4025
rect 56015 3705 56035 4025
rect 56075 3705 56095 4025
rect 56135 3705 56155 4025
rect 56195 3705 56215 4025
rect 56255 3705 56275 4025
rect 56315 3705 56335 4025
rect 56375 3705 56395 4025
rect 56435 3705 56455 4025
rect 56495 3705 56515 4025
rect 56555 3705 56575 4025
rect 56615 3705 56635 4025
rect 56675 3705 56695 4025
rect 56735 3705 56755 4025
rect 57045 3705 57065 4025
rect 57105 3705 57125 4025
rect 57165 3705 57185 4025
rect 57225 3705 57245 4025
rect 57285 3705 57305 4025
rect 57345 3705 57365 4025
rect 57405 3705 57425 4025
rect 57465 3705 57485 4025
rect 57525 3705 57545 4025
rect 57585 3705 57605 4025
rect 57645 3705 57665 4025
rect 57705 3705 57725 4025
rect 57765 3705 57785 4025
rect 58130 3705 58150 4025
rect 58190 3705 58210 4025
rect 58250 3705 58270 4025
rect 58310 3705 58330 4025
rect 58370 3705 58390 4025
rect 58430 3705 58450 4025
rect 58490 3705 58510 4025
rect 58550 3705 58570 4025
rect 58610 3705 58630 4025
rect 58670 3705 58690 4025
rect 58730 3705 58750 4025
rect 58790 3705 58810 4025
rect 58850 3705 58870 4025
rect 54960 2765 54980 3335
rect 55015 2765 55035 3335
rect 55070 2765 55090 3335
rect 55125 2765 55145 3335
rect 55180 2765 55200 3335
rect 55235 2765 55255 3335
rect 55290 2765 55310 3335
rect 55345 2765 55365 3335
rect 55400 2765 55420 3335
rect 55455 2765 55475 3335
rect 55510 2765 55530 3335
rect 55565 2765 55585 3335
rect 55620 2765 55640 3335
rect 56285 3320 56305 3340
rect 56340 3320 56360 3340
rect 56395 3320 56415 3340
rect 56450 3320 56470 3340
rect 56505 3320 56525 3340
rect 56560 3320 56580 3340
rect 56615 3320 56635 3340
rect 56670 3320 56690 3340
rect 56725 3320 56745 3340
rect 56780 3320 56800 3340
rect 56835 3320 56855 3340
rect 56890 3320 56910 3340
rect 56945 3320 56965 3340
rect 57000 3320 57020 3340
rect 57055 3320 57075 3340
rect 57110 3320 57130 3340
rect 57165 3320 57185 3340
rect 57220 3320 57240 3340
rect 57275 3320 57295 3340
rect 57330 3320 57350 3340
rect 57385 3320 57405 3340
rect 57440 3320 57460 3340
rect 57495 3320 57515 3340
rect 56040 2960 56060 2980
rect 56095 2960 56115 2980
rect 56150 2960 56170 2980
rect 56205 2960 56225 2980
rect 56260 2960 56280 2980
rect 56315 2960 56335 2980
rect 56370 2960 56390 2980
rect 56425 2960 56445 2980
rect 56480 2960 56500 2980
rect 56535 2960 56555 2980
rect 56590 2960 56610 2980
rect 56645 2960 56665 2980
rect 56700 2960 56720 2980
rect 57080 2960 57100 2980
rect 57135 2960 57155 2980
rect 57190 2960 57210 2980
rect 57245 2960 57265 2980
rect 57300 2960 57320 2980
rect 57355 2960 57375 2980
rect 57410 2960 57430 2980
rect 57465 2960 57485 2980
rect 57520 2960 57540 2980
rect 57575 2960 57595 2980
rect 57630 2960 57650 2980
rect 57685 2960 57705 2980
rect 57740 2960 57760 2980
rect 58160 2765 58180 3335
rect 58215 2765 58235 3335
rect 58270 2765 58290 3335
rect 58325 2765 58345 3335
rect 58380 2765 58400 3335
rect 58435 2765 58455 3335
rect 58490 2765 58510 3335
rect 58545 2765 58565 3335
rect 58600 2765 58620 3335
rect 58655 2765 58675 3335
rect 58710 2765 58730 3335
rect 58765 2765 58785 3335
rect 58820 2765 58840 3335
rect 54960 2235 54980 2405
rect 55015 2235 55035 2405
rect 55070 2235 55090 2405
rect 55125 2235 55145 2405
rect 55180 2235 55200 2405
rect 55235 2235 55255 2405
rect 55290 2235 55310 2405
rect 55345 2235 55365 2405
rect 55400 2235 55420 2405
rect 55455 2235 55475 2405
rect 55510 2235 55530 2405
rect 55565 2235 55585 2405
rect 55620 2235 55640 2405
rect 58160 2235 58180 2405
rect 58215 2235 58235 2405
rect 58270 2235 58290 2405
rect 58325 2235 58345 2405
rect 58380 2235 58400 2405
rect 58435 2235 58455 2405
rect 58490 2235 58510 2405
rect 58545 2235 58565 2405
rect 58600 2235 58620 2405
rect 58655 2235 58675 2405
rect 58710 2235 58730 2405
rect 58765 2235 58785 2405
rect 58820 2235 58840 2405
<< psubdiff >>
rect 56510 2570 56550 2585
rect 56510 2550 56520 2570
rect 56540 2550 56550 2570
rect 56510 2535 56550 2550
rect 57250 2570 57290 2585
rect 57250 2550 57260 2570
rect 57280 2550 57290 2570
rect 57250 2535 57290 2550
rect 55990 2165 56030 2180
rect 55990 2045 56000 2165
rect 56020 2045 56030 2165
rect 55990 2030 56030 2045
rect 56730 2165 56770 2180
rect 56730 2045 56740 2165
rect 56760 2045 56770 2165
rect 56730 2030 56770 2045
rect 57030 2165 57070 2180
rect 57030 2045 57040 2165
rect 57060 2045 57070 2165
rect 57030 2030 57070 2045
rect 57770 2165 57810 2180
rect 57770 2045 57780 2165
rect 57800 2045 57810 2165
rect 57770 2030 57810 2045
rect 54910 1845 54950 1860
rect 54910 1575 54920 1845
rect 54940 1575 54950 1845
rect 54910 1560 54950 1575
rect 55650 1845 55690 1860
rect 55650 1575 55660 1845
rect 55680 1575 55690 1845
rect 58110 1845 58150 1860
rect 55650 1560 55690 1575
rect 55990 1695 56030 1710
rect 55990 1575 56000 1695
rect 56020 1575 56030 1695
rect 55990 1560 56030 1575
rect 56730 1695 56770 1710
rect 56730 1575 56740 1695
rect 56760 1575 56770 1695
rect 56730 1560 56770 1575
rect 57030 1695 57070 1710
rect 57030 1575 57040 1695
rect 57060 1575 57070 1695
rect 57030 1560 57070 1575
rect 57770 1695 57810 1710
rect 57770 1575 57780 1695
rect 57800 1575 57810 1695
rect 57770 1560 57810 1575
rect 58110 1575 58120 1845
rect 58140 1575 58150 1845
rect 58110 1560 58150 1575
rect 58850 1845 58890 1860
rect 58850 1575 58860 1845
rect 58880 1575 58890 1845
rect 58850 1560 58890 1575
rect 54945 1155 54985 1170
rect 54945 485 54955 1155
rect 54975 485 54985 1155
rect 54945 470 54985 485
rect 55625 1155 55665 1170
rect 55625 485 55635 1155
rect 55655 485 55665 1155
rect 56180 1145 56220 1160
rect 56180 925 56190 1145
rect 56210 925 56220 1145
rect 56180 910 56220 925
rect 57525 1145 57565 1160
rect 57525 925 57535 1145
rect 57555 925 57565 1145
rect 57525 910 57565 925
rect 58140 1155 58180 1170
rect 56390 680 56430 695
rect 56390 560 56400 680
rect 56420 560 56430 680
rect 56390 545 56430 560
rect 56800 680 56840 695
rect 56800 560 56810 680
rect 56830 560 56840 680
rect 56800 545 56840 560
rect 55625 470 55665 485
rect 58140 485 58150 1155
rect 58170 485 58180 1155
rect 58140 470 58180 485
rect 58820 1155 58860 1170
rect 58820 485 58830 1155
rect 58850 485 58860 1155
rect 58820 470 58860 485
<< nsubdiff >>
rect 56045 4695 56085 4710
rect 56045 4375 56055 4695
rect 56075 4375 56085 4695
rect 56045 4360 56085 4375
rect 56305 4695 56345 4710
rect 56305 4375 56315 4695
rect 56335 4375 56345 4695
rect 56985 4695 57025 4710
rect 56305 4360 56345 4375
rect 56515 4525 56555 4540
rect 56515 4375 56525 4525
rect 56545 4375 56555 4525
rect 56515 4360 56555 4375
rect 56775 4525 56815 4540
rect 56775 4375 56785 4525
rect 56805 4375 56815 4525
rect 56775 4360 56815 4375
rect 56985 4375 56995 4695
rect 57015 4375 57025 4695
rect 56985 4360 57025 4375
rect 57245 4695 57285 4710
rect 57245 4375 57255 4695
rect 57275 4375 57285 4695
rect 57245 4360 57285 4375
rect 57455 4695 57495 4710
rect 57455 4375 57465 4695
rect 57485 4375 57495 4695
rect 57455 4360 57495 4375
rect 57715 4695 57755 4710
rect 57715 4375 57725 4695
rect 57745 4375 57755 4695
rect 57715 4360 57755 4375
rect 54885 4025 54925 4040
rect 54885 3705 54895 4025
rect 54915 3705 54925 4025
rect 54885 3690 54925 3705
rect 55685 4025 55725 4040
rect 55685 3705 55695 4025
rect 55715 3705 55725 4025
rect 55685 3690 55725 3705
rect 55965 4025 56005 4040
rect 55965 3705 55975 4025
rect 55995 3705 56005 4025
rect 55965 3690 56005 3705
rect 56765 4025 56805 4040
rect 56765 3705 56775 4025
rect 56795 3705 56805 4025
rect 56765 3690 56805 3705
rect 56995 4025 57035 4040
rect 56995 3705 57005 4025
rect 57025 3705 57035 4025
rect 56995 3690 57035 3705
rect 57795 4025 57835 4040
rect 57795 3705 57805 4025
rect 57825 3705 57835 4025
rect 57795 3690 57835 3705
rect 58080 4025 58120 4040
rect 58080 3705 58090 4025
rect 58110 3705 58120 4025
rect 58080 3690 58120 3705
rect 58880 4025 58920 4040
rect 58880 3705 58890 4025
rect 58910 3705 58920 4025
rect 58880 3690 58920 3705
rect 54910 3335 54950 3350
rect 54910 2765 54920 3335
rect 54940 2765 54950 3335
rect 54910 2750 54950 2765
rect 55650 3335 55690 3350
rect 55650 2765 55660 3335
rect 55680 2765 55690 3335
rect 56235 3340 56275 3355
rect 56235 3320 56245 3340
rect 56265 3320 56275 3340
rect 56235 3305 56275 3320
rect 57525 3340 57565 3355
rect 57525 3320 57535 3340
rect 57555 3320 57565 3340
rect 57525 3305 57565 3320
rect 58110 3335 58150 3350
rect 55990 2980 56030 2995
rect 55990 2960 56000 2980
rect 56020 2960 56030 2980
rect 55990 2945 56030 2960
rect 56730 2980 56770 2995
rect 56730 2960 56740 2980
rect 56760 2960 56770 2980
rect 56730 2945 56770 2960
rect 57030 2980 57070 2995
rect 57030 2960 57040 2980
rect 57060 2960 57070 2980
rect 57030 2945 57070 2960
rect 57770 2980 57810 2995
rect 57770 2960 57780 2980
rect 57800 2960 57810 2980
rect 57770 2945 57810 2960
rect 55650 2750 55690 2765
rect 58110 2765 58120 3335
rect 58140 2765 58150 3335
rect 58110 2750 58150 2765
rect 58850 3335 58890 3350
rect 58850 2765 58860 3335
rect 58880 2765 58890 3335
rect 58850 2750 58890 2765
rect 54910 2405 54950 2420
rect 54910 2235 54920 2405
rect 54940 2235 54950 2405
rect 54910 2220 54950 2235
rect 55650 2405 55690 2420
rect 55650 2235 55660 2405
rect 55680 2235 55690 2405
rect 58110 2405 58150 2420
rect 55650 2220 55690 2235
rect 58110 2235 58120 2405
rect 58140 2235 58150 2405
rect 58110 2220 58150 2235
rect 58850 2405 58890 2420
rect 58850 2235 58860 2405
rect 58880 2235 58890 2405
rect 58850 2220 58890 2235
<< psubdiffcont >>
rect 56520 2550 56540 2570
rect 57260 2550 57280 2570
rect 56000 2045 56020 2165
rect 56740 2045 56760 2165
rect 57040 2045 57060 2165
rect 57780 2045 57800 2165
rect 54920 1575 54940 1845
rect 55660 1575 55680 1845
rect 56000 1575 56020 1695
rect 56740 1575 56760 1695
rect 57040 1575 57060 1695
rect 57780 1575 57800 1695
rect 58120 1575 58140 1845
rect 58860 1575 58880 1845
rect 54955 485 54975 1155
rect 55635 485 55655 1155
rect 56190 925 56210 1145
rect 57535 925 57555 1145
rect 56400 560 56420 680
rect 56810 560 56830 680
rect 58150 485 58170 1155
rect 58830 485 58850 1155
<< nsubdiffcont >>
rect 56055 4375 56075 4695
rect 56315 4375 56335 4695
rect 56525 4375 56545 4525
rect 56785 4375 56805 4525
rect 56995 4375 57015 4695
rect 57255 4375 57275 4695
rect 57465 4375 57485 4695
rect 57725 4375 57745 4695
rect 54895 3705 54915 4025
rect 55695 3705 55715 4025
rect 55975 3705 55995 4025
rect 56775 3705 56795 4025
rect 57005 3705 57025 4025
rect 57805 3705 57825 4025
rect 58090 3705 58110 4025
rect 58890 3705 58910 4025
rect 54920 2765 54940 3335
rect 55660 2765 55680 3335
rect 56245 3320 56265 3340
rect 57535 3320 57555 3340
rect 56000 2960 56020 2980
rect 56740 2960 56760 2980
rect 57040 2960 57060 2980
rect 57780 2960 57800 2980
rect 58120 2765 58140 3335
rect 58860 2765 58880 3335
rect 54920 2235 54940 2405
rect 55660 2235 55680 2405
rect 58120 2235 58140 2405
rect 58860 2235 58880 2405
<< poly >>
rect 56085 4755 56125 4765
rect 56085 4735 56095 4755
rect 56115 4740 56125 4755
rect 56265 4755 56305 4765
rect 56265 4740 56275 4755
rect 56115 4735 56145 4740
rect 56085 4725 56145 4735
rect 56245 4735 56275 4740
rect 56295 4735 56305 4755
rect 56245 4725 56305 4735
rect 57025 4755 57065 4765
rect 57025 4735 57035 4755
rect 57055 4740 57065 4755
rect 57205 4755 57245 4765
rect 57205 4740 57215 4755
rect 57055 4735 57085 4740
rect 57025 4725 57085 4735
rect 57185 4735 57215 4740
rect 57235 4735 57245 4755
rect 57185 4725 57245 4735
rect 57495 4755 57535 4765
rect 57495 4735 57505 4755
rect 57525 4740 57535 4755
rect 57675 4755 57715 4765
rect 57675 4740 57685 4755
rect 57525 4735 57555 4740
rect 57495 4725 57555 4735
rect 57655 4735 57685 4740
rect 57705 4735 57715 4755
rect 57655 4725 57715 4735
rect 56125 4710 56145 4725
rect 56185 4710 56205 4725
rect 56245 4710 56265 4725
rect 57065 4710 57085 4725
rect 57125 4710 57145 4725
rect 57185 4710 57205 4725
rect 57535 4710 57555 4725
rect 57595 4710 57615 4725
rect 57655 4710 57675 4725
rect 56555 4585 56595 4595
rect 56555 4565 56565 4585
rect 56585 4570 56595 4585
rect 56735 4585 56775 4595
rect 56735 4570 56745 4585
rect 56585 4565 56615 4570
rect 56555 4555 56615 4565
rect 56715 4565 56745 4570
rect 56765 4565 56775 4585
rect 56715 4555 56775 4565
rect 56595 4540 56615 4555
rect 56655 4540 56675 4555
rect 56715 4540 56735 4555
rect 56125 4345 56145 4360
rect 56185 4315 56205 4360
rect 56245 4345 56265 4360
rect 56595 4345 56615 4360
rect 56655 4315 56675 4360
rect 56715 4345 56735 4360
rect 57065 4345 57085 4360
rect 56150 4305 56205 4315
rect 56150 4285 56160 4305
rect 56180 4285 56205 4305
rect 56150 4275 56205 4285
rect 56630 4305 56675 4315
rect 56630 4285 56635 4305
rect 56655 4300 56675 4305
rect 57125 4315 57145 4360
rect 57185 4345 57205 4360
rect 57535 4345 57555 4360
rect 57125 4305 57170 4315
rect 57595 4305 57615 4360
rect 57655 4345 57675 4360
rect 57125 4300 57145 4305
rect 56655 4285 56660 4300
rect 56630 4275 56660 4285
rect 57140 4285 57145 4300
rect 57165 4285 57170 4305
rect 57140 4275 57170 4285
rect 57576 4295 57615 4305
rect 57576 4275 57581 4295
rect 57601 4290 57615 4295
rect 57601 4275 57606 4290
rect 57576 4265 57606 4275
rect 54930 4085 54960 4095
rect 54930 4065 54935 4085
rect 54955 4070 54960 4085
rect 55650 4085 55680 4095
rect 55650 4070 55655 4085
rect 54955 4065 54985 4070
rect 54930 4055 54985 4065
rect 55625 4065 55655 4070
rect 55675 4065 55680 4085
rect 55625 4055 55680 4065
rect 56010 4085 56040 4095
rect 56010 4065 56015 4085
rect 56035 4070 56040 4085
rect 56730 4085 56760 4095
rect 56730 4070 56735 4085
rect 56035 4065 56065 4070
rect 56010 4055 56065 4065
rect 56705 4065 56735 4070
rect 56755 4065 56760 4085
rect 56705 4055 56760 4065
rect 57040 4085 57070 4095
rect 57040 4065 57045 4085
rect 57065 4070 57070 4085
rect 57760 4085 57790 4095
rect 57760 4070 57765 4085
rect 57065 4065 57095 4070
rect 57040 4055 57095 4065
rect 57735 4065 57765 4070
rect 57785 4065 57790 4085
rect 57735 4055 57790 4065
rect 58125 4085 58155 4095
rect 58125 4065 58130 4085
rect 58150 4070 58155 4085
rect 58845 4085 58875 4095
rect 58845 4070 58850 4085
rect 58150 4065 58180 4070
rect 58125 4055 58180 4065
rect 58820 4065 58850 4070
rect 58870 4065 58875 4085
rect 58820 4055 58875 4065
rect 54965 4040 54985 4055
rect 55025 4040 55045 4055
rect 55085 4040 55105 4055
rect 55145 4040 55165 4055
rect 55205 4040 55225 4055
rect 55265 4040 55285 4055
rect 55325 4040 55345 4055
rect 55385 4040 55405 4055
rect 55445 4040 55465 4055
rect 55505 4040 55525 4055
rect 55565 4040 55585 4055
rect 55625 4040 55645 4055
rect 56045 4040 56065 4055
rect 56105 4040 56125 4055
rect 56165 4040 56185 4055
rect 56225 4040 56245 4055
rect 56285 4040 56305 4055
rect 56345 4040 56365 4055
rect 56405 4040 56425 4055
rect 56465 4040 56485 4055
rect 56525 4040 56545 4055
rect 56585 4040 56605 4055
rect 56645 4040 56665 4055
rect 56705 4040 56725 4055
rect 57075 4040 57095 4055
rect 57135 4040 57155 4055
rect 57195 4040 57215 4055
rect 57255 4040 57275 4055
rect 57315 4040 57335 4055
rect 57375 4040 57395 4055
rect 57435 4040 57455 4055
rect 57495 4040 57515 4055
rect 57555 4040 57575 4055
rect 57615 4040 57635 4055
rect 57675 4040 57695 4055
rect 57735 4040 57755 4055
rect 58160 4040 58180 4055
rect 58220 4040 58240 4055
rect 58280 4040 58300 4055
rect 58340 4040 58360 4055
rect 58400 4040 58420 4055
rect 58460 4040 58480 4055
rect 58520 4040 58540 4055
rect 58580 4040 58600 4055
rect 58640 4040 58660 4055
rect 58700 4040 58720 4055
rect 58760 4040 58780 4055
rect 58820 4040 58840 4055
rect 54965 3675 54985 3690
rect 55025 3680 55045 3690
rect 55085 3680 55105 3690
rect 55145 3680 55165 3690
rect 55205 3680 55225 3690
rect 55265 3680 55285 3690
rect 55325 3680 55345 3690
rect 55385 3680 55405 3690
rect 55445 3680 55465 3690
rect 55505 3680 55525 3690
rect 55565 3680 55585 3690
rect 55025 3665 55585 3680
rect 55325 3545 55345 3665
rect 55625 3660 55645 3690
rect 56045 3675 56065 3690
rect 56105 3680 56125 3690
rect 56165 3680 56185 3690
rect 56225 3680 56245 3690
rect 56285 3680 56305 3690
rect 56345 3680 56365 3690
rect 56405 3680 56425 3690
rect 56465 3680 56485 3690
rect 56525 3680 56545 3690
rect 56585 3680 56605 3690
rect 56645 3680 56665 3690
rect 56105 3665 56665 3680
rect 56705 3675 56725 3690
rect 57075 3675 57095 3690
rect 57135 3680 57155 3690
rect 57195 3680 57215 3690
rect 57255 3680 57275 3690
rect 57315 3680 57335 3690
rect 57375 3680 57395 3690
rect 57435 3680 57455 3690
rect 57495 3680 57515 3690
rect 57555 3680 57575 3690
rect 57615 3680 57635 3690
rect 57675 3680 57695 3690
rect 57135 3665 57695 3680
rect 57735 3675 57755 3690
rect 56405 3590 56425 3665
rect 57375 3590 57395 3665
rect 58160 3660 58180 3690
rect 58220 3680 58240 3690
rect 58280 3680 58300 3690
rect 58340 3680 58360 3690
rect 58400 3680 58420 3690
rect 58460 3680 58480 3690
rect 58520 3680 58540 3690
rect 58580 3680 58600 3690
rect 58640 3680 58660 3690
rect 58700 3680 58720 3690
rect 58760 3680 58780 3690
rect 58220 3665 58780 3680
rect 58820 3675 58840 3690
rect 56395 3580 56435 3590
rect 56395 3560 56405 3580
rect 56425 3560 56435 3580
rect 56395 3550 56435 3560
rect 57365 3580 57405 3590
rect 57365 3560 57375 3580
rect 57395 3560 57405 3580
rect 57365 3550 57405 3560
rect 58460 3545 58480 3665
rect 55315 3535 55355 3545
rect 55315 3515 55325 3535
rect 55345 3515 55355 3535
rect 55315 3505 55355 3515
rect 58450 3535 58490 3545
rect 58450 3515 58460 3535
rect 58480 3515 58490 3535
rect 58450 3505 58490 3515
rect 54955 3395 54985 3405
rect 54955 3375 54960 3395
rect 54980 3380 54985 3395
rect 55615 3395 55645 3405
rect 55615 3380 55620 3395
rect 54980 3375 55005 3380
rect 54955 3365 55005 3375
rect 55595 3375 55620 3380
rect 55640 3375 55645 3395
rect 55595 3365 55645 3375
rect 58155 3395 58185 3405
rect 58155 3375 58160 3395
rect 58180 3380 58185 3395
rect 58815 3395 58845 3405
rect 58815 3380 58820 3395
rect 58180 3375 58205 3380
rect 54990 3350 55005 3365
rect 55045 3350 55060 3365
rect 55100 3350 55115 3365
rect 55155 3350 55170 3365
rect 55210 3350 55225 3365
rect 55265 3350 55280 3365
rect 55320 3350 55335 3365
rect 55375 3350 55390 3365
rect 55430 3350 55445 3365
rect 55485 3350 55500 3365
rect 55540 3350 55555 3365
rect 55595 3350 55610 3365
rect 56315 3355 56330 3370
rect 56370 3355 56385 3370
rect 56425 3355 56440 3370
rect 56480 3355 56495 3370
rect 56535 3355 56550 3370
rect 56590 3355 56605 3370
rect 56645 3355 56660 3370
rect 56700 3355 56715 3370
rect 56755 3355 56770 3370
rect 56810 3355 56825 3370
rect 56865 3355 56880 3370
rect 56920 3355 56935 3370
rect 56975 3355 56990 3370
rect 57030 3355 57045 3370
rect 57085 3355 57100 3370
rect 57140 3355 57155 3370
rect 57195 3355 57210 3370
rect 57250 3355 57265 3370
rect 57305 3355 57320 3370
rect 57360 3355 57375 3370
rect 57415 3355 57430 3370
rect 57470 3355 57485 3370
rect 58155 3365 58205 3375
rect 58795 3375 58820 3380
rect 58840 3375 58845 3395
rect 58795 3365 58845 3375
rect 58190 3350 58205 3365
rect 58245 3350 58260 3365
rect 58300 3350 58315 3365
rect 58355 3350 58370 3365
rect 58410 3350 58425 3365
rect 58465 3350 58480 3365
rect 58520 3350 58535 3365
rect 58575 3350 58590 3365
rect 58630 3350 58645 3365
rect 58685 3350 58700 3365
rect 58740 3350 58755 3365
rect 58795 3350 58810 3365
rect 56315 3290 56330 3305
rect 56280 3280 56330 3290
rect 56370 3295 56385 3305
rect 56425 3295 56440 3305
rect 56480 3295 56495 3305
rect 56535 3295 56550 3305
rect 56590 3295 56605 3305
rect 56645 3295 56660 3305
rect 56700 3295 56715 3305
rect 56755 3295 56770 3305
rect 56810 3295 56825 3305
rect 56865 3295 56880 3305
rect 56920 3295 56935 3305
rect 56975 3295 56990 3305
rect 57030 3295 57045 3305
rect 57085 3295 57100 3305
rect 57140 3295 57155 3305
rect 57195 3295 57210 3305
rect 57250 3295 57265 3305
rect 57305 3295 57320 3305
rect 57360 3295 57375 3305
rect 57415 3295 57430 3305
rect 56370 3280 57430 3295
rect 57470 3290 57485 3305
rect 57470 3280 57520 3290
rect 56280 3260 56285 3280
rect 56305 3275 56330 3280
rect 56305 3260 56310 3275
rect 56280 3250 56310 3260
rect 56810 3160 56825 3280
rect 57470 3275 57495 3280
rect 57490 3260 57495 3275
rect 57515 3260 57520 3280
rect 57490 3250 57520 3260
rect 56795 3150 56835 3160
rect 56795 3130 56805 3150
rect 56825 3130 56835 3150
rect 56795 3120 56835 3130
rect 55990 3065 56020 3075
rect 55990 3045 55995 3065
rect 56015 3050 56020 3065
rect 56740 3065 56770 3075
rect 56740 3050 56745 3065
rect 56015 3045 56745 3050
rect 56765 3045 56770 3065
rect 55990 3035 56770 3045
rect 57030 3065 57060 3075
rect 57030 3045 57035 3065
rect 57055 3050 57060 3065
rect 57780 3065 57810 3075
rect 57780 3050 57785 3065
rect 57055 3045 57785 3050
rect 57805 3045 57810 3065
rect 57030 3035 57810 3045
rect 56070 2995 56085 3010
rect 56125 2995 56140 3010
rect 56180 2995 56195 3035
rect 56235 2995 56250 3035
rect 56290 2995 56305 3010
rect 56345 2995 56360 3010
rect 56400 2995 56415 3035
rect 56455 2995 56470 3035
rect 56510 2995 56525 3010
rect 56565 2995 56580 3010
rect 56620 2995 56635 3035
rect 56675 2995 56690 3010
rect 57110 2995 57125 3010
rect 57165 2995 57180 3035
rect 57220 2995 57235 3010
rect 57275 2995 57290 3010
rect 57330 2995 57345 3035
rect 57385 2995 57400 3035
rect 57440 2995 57455 3010
rect 57495 2995 57510 3010
rect 57550 2995 57565 3035
rect 57605 2995 57620 3035
rect 57660 2995 57675 3010
rect 57715 2995 57730 3010
rect 56070 2930 56085 2945
rect 56035 2920 56085 2930
rect 56035 2900 56040 2920
rect 56060 2915 56085 2920
rect 56060 2900 56065 2915
rect 56035 2890 56065 2900
rect 56125 2905 56140 2945
rect 56180 2930 56195 2945
rect 56235 2930 56250 2945
rect 56290 2905 56305 2945
rect 56345 2905 56360 2945
rect 56400 2930 56415 2945
rect 56455 2930 56470 2945
rect 56510 2905 56525 2945
rect 56565 2905 56580 2945
rect 56620 2930 56635 2945
rect 56675 2930 56690 2945
rect 57110 2930 57125 2945
rect 57165 2930 57180 2945
rect 56675 2920 56725 2930
rect 56675 2915 56700 2920
rect 56125 2890 56580 2905
rect 56695 2900 56700 2915
rect 56720 2900 56725 2920
rect 56695 2890 56725 2900
rect 57075 2920 57125 2930
rect 57075 2900 57080 2920
rect 57100 2915 57125 2920
rect 57100 2900 57105 2915
rect 57075 2890 57105 2900
rect 57220 2905 57235 2945
rect 57275 2905 57290 2945
rect 57330 2930 57345 2945
rect 57385 2930 57400 2945
rect 57440 2905 57455 2945
rect 57495 2905 57510 2945
rect 57550 2930 57565 2945
rect 57605 2930 57620 2945
rect 57660 2905 57675 2945
rect 57715 2930 57730 2945
rect 57715 2920 57765 2930
rect 57715 2915 57740 2920
rect 57220 2890 57675 2905
rect 57735 2900 57740 2915
rect 57760 2900 57765 2920
rect 57735 2890 57765 2900
rect 56125 2845 56140 2890
rect 56095 2835 56140 2845
rect 56095 2815 56100 2835
rect 56120 2825 56140 2835
rect 56565 2845 56580 2890
rect 57220 2845 57235 2890
rect 56565 2835 56610 2845
rect 56565 2825 56585 2835
rect 56120 2815 56125 2825
rect 56095 2805 56125 2815
rect 56580 2815 56585 2825
rect 56605 2815 56610 2835
rect 56580 2805 56610 2815
rect 57190 2835 57235 2845
rect 57190 2815 57195 2835
rect 57215 2825 57235 2835
rect 57215 2815 57220 2825
rect 57190 2805 57220 2815
rect 54990 2735 55005 2750
rect 55045 2740 55060 2750
rect 55100 2740 55115 2750
rect 55155 2740 55170 2750
rect 55210 2740 55225 2750
rect 55265 2740 55280 2750
rect 55320 2740 55335 2750
rect 55375 2740 55390 2750
rect 55430 2740 55445 2750
rect 55485 2740 55500 2750
rect 55540 2740 55555 2750
rect 55045 2725 55555 2740
rect 55595 2735 55610 2750
rect 58190 2735 58205 2750
rect 58245 2740 58260 2750
rect 58300 2740 58315 2750
rect 58355 2740 58370 2750
rect 58410 2740 58425 2750
rect 58465 2740 58480 2750
rect 58520 2740 58535 2750
rect 58575 2740 58590 2750
rect 58630 2740 58645 2750
rect 58685 2740 58700 2750
rect 58740 2740 58755 2750
rect 58245 2725 58755 2740
rect 58795 2735 58810 2750
rect 55320 2645 55335 2725
rect 58465 2645 58480 2725
rect 55310 2635 55350 2645
rect 55310 2615 55320 2635
rect 55340 2615 55350 2635
rect 55310 2605 55350 2615
rect 56715 2630 56755 2640
rect 56715 2610 56725 2630
rect 56745 2610 56755 2630
rect 56935 2630 56975 2640
rect 56935 2610 56945 2630
rect 56965 2610 56975 2630
rect 58450 2635 58490 2645
rect 58450 2615 58460 2635
rect 58480 2615 58490 2635
rect 56590 2585 56605 2600
rect 56645 2595 57155 2610
rect 58450 2605 58490 2615
rect 56645 2585 56660 2595
rect 56700 2585 56715 2595
rect 56755 2585 56770 2595
rect 56810 2585 56825 2595
rect 56865 2585 56880 2595
rect 56920 2585 56935 2595
rect 56975 2585 56990 2595
rect 57030 2585 57045 2595
rect 57085 2585 57100 2595
rect 57140 2585 57155 2595
rect 57195 2585 57210 2600
rect 56590 2520 56605 2535
rect 56645 2520 56660 2535
rect 56700 2520 56715 2535
rect 56755 2520 56770 2535
rect 56810 2520 56825 2535
rect 56865 2520 56880 2535
rect 56920 2520 56935 2535
rect 56975 2520 56990 2535
rect 57030 2520 57045 2535
rect 57085 2520 57100 2535
rect 57140 2520 57155 2535
rect 57195 2520 57210 2535
rect 56550 2510 56605 2520
rect 56550 2490 56560 2510
rect 56580 2505 56605 2510
rect 57195 2510 57250 2520
rect 57195 2505 57220 2510
rect 56580 2490 56590 2505
rect 56550 2480 56590 2490
rect 57210 2490 57220 2505
rect 57240 2490 57250 2510
rect 57210 2480 57250 2490
rect 54955 2465 54985 2475
rect 54955 2445 54960 2465
rect 54980 2450 54985 2465
rect 55615 2465 55645 2475
rect 55615 2450 55620 2465
rect 54980 2445 55005 2450
rect 54955 2435 55005 2445
rect 55595 2445 55620 2450
rect 55640 2445 55645 2465
rect 55595 2435 55645 2445
rect 58155 2465 58185 2475
rect 58155 2445 58160 2465
rect 58180 2450 58185 2465
rect 58815 2465 58845 2475
rect 58815 2450 58820 2465
rect 58180 2445 58205 2450
rect 58155 2435 58205 2445
rect 58795 2445 58820 2450
rect 58840 2445 58845 2465
rect 58795 2435 58845 2445
rect 54990 2420 55005 2435
rect 55045 2420 55060 2435
rect 55100 2420 55115 2435
rect 55155 2420 55170 2435
rect 55210 2420 55225 2435
rect 55265 2420 55280 2435
rect 55320 2420 55335 2435
rect 55375 2420 55390 2435
rect 55430 2420 55445 2435
rect 55485 2420 55500 2435
rect 55540 2420 55555 2435
rect 55595 2420 55610 2435
rect 58190 2420 58205 2435
rect 58245 2420 58260 2435
rect 58300 2420 58315 2435
rect 58355 2420 58370 2435
rect 58410 2420 58425 2435
rect 58465 2420 58480 2435
rect 58520 2420 58535 2435
rect 58575 2420 58590 2435
rect 58630 2420 58645 2435
rect 58685 2420 58700 2435
rect 58740 2420 58755 2435
rect 58795 2420 58810 2435
rect 56635 2265 56665 2275
rect 56635 2250 56640 2265
rect 56620 2245 56640 2250
rect 56660 2245 56665 2265
rect 56620 2235 56665 2245
rect 57135 2265 57165 2275
rect 57135 2245 57140 2265
rect 57160 2250 57165 2265
rect 57160 2245 57180 2250
rect 57135 2235 57180 2245
rect 57785 2240 57815 2250
rect 57785 2235 57790 2240
rect 54990 2205 55005 2220
rect 55045 2210 55060 2220
rect 55100 2210 55115 2220
rect 55155 2210 55170 2220
rect 55210 2210 55225 2220
rect 55265 2210 55280 2220
rect 55320 2210 55335 2220
rect 55375 2210 55390 2220
rect 55430 2210 55445 2220
rect 55485 2210 55500 2220
rect 55540 2210 55555 2220
rect 55045 2195 55555 2210
rect 55595 2205 55610 2220
rect 56620 2205 56635 2235
rect 55320 2055 55335 2195
rect 56070 2180 56085 2195
rect 56125 2190 56635 2205
rect 57165 2205 57180 2235
rect 57660 2220 57790 2235
rect 57810 2220 57815 2240
rect 57660 2205 57675 2220
rect 57785 2210 57815 2220
rect 58190 2205 58205 2220
rect 58245 2210 58260 2220
rect 58300 2210 58315 2220
rect 58355 2210 58370 2220
rect 58410 2210 58425 2220
rect 58465 2210 58480 2220
rect 58520 2210 58535 2220
rect 58575 2210 58590 2220
rect 58630 2210 58645 2220
rect 58685 2210 58700 2220
rect 58740 2210 58755 2220
rect 56125 2180 56140 2190
rect 56180 2180 56195 2190
rect 56235 2180 56250 2190
rect 56290 2180 56305 2190
rect 56345 2180 56360 2190
rect 56400 2180 56415 2190
rect 56455 2180 56470 2190
rect 56510 2180 56525 2190
rect 56565 2180 56580 2190
rect 56620 2180 56635 2190
rect 56675 2180 56690 2195
rect 57110 2180 57125 2195
rect 57165 2190 57675 2205
rect 58245 2195 58755 2210
rect 58795 2205 58810 2220
rect 57165 2180 57180 2190
rect 57220 2180 57235 2190
rect 57275 2180 57290 2190
rect 57330 2180 57345 2190
rect 57385 2180 57400 2190
rect 57440 2180 57455 2190
rect 57495 2180 57510 2190
rect 57550 2180 57565 2190
rect 57605 2180 57620 2190
rect 57660 2180 57675 2190
rect 57715 2180 57730 2195
rect 55310 2045 55350 2055
rect 55310 2025 55320 2045
rect 55340 2025 55350 2045
rect 58465 2055 58480 2195
rect 58450 2045 58490 2055
rect 55310 2015 55350 2025
rect 56070 2015 56085 2030
rect 56125 2015 56140 2030
rect 56180 2015 56195 2030
rect 56235 2015 56250 2030
rect 56290 2015 56305 2030
rect 56345 2015 56360 2030
rect 56400 2015 56415 2030
rect 56455 2015 56470 2030
rect 56510 2015 56525 2030
rect 56565 2015 56580 2030
rect 56620 2015 56635 2030
rect 56675 2015 56690 2030
rect 57110 2015 57125 2030
rect 57165 2015 57180 2030
rect 57220 2015 57235 2030
rect 57275 2015 57290 2030
rect 57330 2015 57345 2030
rect 57385 2015 57400 2030
rect 57440 2015 57455 2030
rect 57495 2015 57510 2030
rect 57550 2015 57565 2030
rect 57605 2015 57620 2030
rect 57660 2015 57675 2030
rect 57715 2015 57730 2030
rect 58450 2025 58460 2045
rect 58480 2025 58490 2045
rect 58450 2015 58490 2025
rect 55320 1885 55335 2015
rect 56035 2005 56085 2015
rect 56035 1985 56040 2005
rect 56060 2000 56085 2005
rect 56675 2005 56725 2015
rect 56675 2000 56700 2005
rect 56060 1985 56065 2000
rect 56035 1975 56065 1985
rect 56695 1985 56700 2000
rect 56720 1985 56725 2005
rect 56695 1975 56725 1985
rect 57075 2005 57125 2015
rect 57075 1985 57080 2005
rect 57100 2000 57125 2005
rect 57715 2005 57765 2015
rect 57715 2000 57740 2005
rect 57100 1985 57105 2000
rect 57075 1975 57105 1985
rect 57735 1985 57740 2000
rect 57760 1985 57765 2005
rect 57735 1975 57765 1985
rect 58465 1885 58480 2015
rect 54990 1860 55005 1875
rect 55045 1870 55555 1885
rect 55045 1860 55060 1870
rect 55100 1860 55115 1870
rect 55155 1860 55170 1870
rect 55210 1860 55225 1870
rect 55265 1860 55280 1870
rect 55320 1860 55335 1870
rect 55375 1860 55390 1870
rect 55430 1860 55445 1870
rect 55485 1860 55500 1870
rect 55540 1860 55555 1870
rect 55595 1860 55610 1875
rect 58190 1860 58205 1875
rect 58245 1870 58755 1885
rect 58245 1860 58260 1870
rect 58300 1860 58315 1870
rect 58355 1860 58370 1870
rect 58410 1860 58425 1870
rect 58465 1860 58480 1870
rect 58520 1860 58535 1870
rect 58575 1860 58590 1870
rect 58630 1860 58645 1870
rect 58685 1860 58700 1870
rect 58740 1860 58755 1870
rect 58795 1860 58810 1875
rect 55990 1780 56020 1790
rect 55990 1760 55995 1780
rect 56015 1765 56020 1780
rect 56690 1780 56720 1790
rect 56690 1765 56695 1780
rect 56015 1760 56140 1765
rect 55990 1750 56140 1760
rect 56125 1735 56140 1750
rect 56620 1760 56695 1765
rect 56715 1760 56720 1780
rect 56620 1750 56720 1760
rect 56859 1780 56889 1790
rect 56859 1760 56864 1780
rect 56884 1760 56889 1780
rect 56859 1750 56889 1760
rect 56911 1780 56941 1790
rect 56911 1760 56916 1780
rect 56936 1760 56941 1780
rect 56911 1750 56941 1760
rect 57080 1780 57110 1790
rect 57080 1760 57085 1780
rect 57105 1765 57110 1780
rect 57780 1780 57810 1790
rect 57780 1765 57785 1780
rect 57105 1760 57180 1765
rect 57080 1750 57180 1760
rect 56620 1735 56635 1750
rect 56070 1710 56085 1725
rect 56125 1720 56635 1735
rect 56125 1710 56140 1720
rect 56180 1710 56195 1720
rect 56235 1710 56250 1720
rect 56290 1710 56305 1720
rect 56345 1710 56360 1720
rect 56400 1710 56415 1720
rect 56455 1710 56470 1720
rect 56510 1710 56525 1720
rect 56565 1710 56580 1720
rect 56620 1710 56635 1720
rect 56675 1710 56690 1725
rect 56810 1710 56825 1725
rect 56865 1710 56880 1750
rect 56920 1710 56935 1750
rect 57165 1735 57180 1750
rect 57660 1760 57785 1765
rect 57805 1760 57810 1780
rect 57660 1750 57810 1760
rect 57660 1735 57675 1750
rect 56975 1710 56990 1725
rect 57110 1710 57125 1725
rect 57165 1720 57675 1735
rect 57165 1710 57180 1720
rect 57220 1710 57235 1720
rect 57275 1710 57290 1720
rect 57330 1710 57345 1720
rect 57385 1710 57400 1720
rect 57440 1710 57455 1720
rect 57495 1710 57510 1720
rect 57550 1710 57565 1720
rect 57605 1710 57620 1720
rect 57660 1710 57675 1720
rect 57715 1710 57730 1725
rect 54990 1545 55005 1560
rect 55045 1545 55060 1560
rect 55100 1545 55115 1560
rect 55155 1545 55170 1560
rect 55210 1545 55225 1560
rect 55265 1545 55280 1560
rect 55320 1545 55335 1560
rect 55375 1545 55390 1560
rect 55430 1545 55445 1560
rect 55485 1545 55500 1560
rect 55540 1545 55555 1560
rect 55595 1545 55610 1560
rect 56070 1545 56085 1560
rect 56125 1545 56140 1560
rect 56180 1545 56195 1560
rect 56235 1545 56250 1560
rect 56290 1545 56305 1560
rect 56345 1545 56360 1560
rect 56400 1545 56415 1560
rect 56455 1545 56470 1560
rect 56510 1545 56525 1560
rect 56565 1545 56580 1560
rect 56620 1545 56635 1560
rect 56675 1545 56690 1560
rect 56810 1545 56825 1560
rect 56865 1545 56880 1560
rect 56920 1545 56935 1560
rect 56975 1545 56990 1560
rect 57110 1545 57125 1560
rect 57165 1545 57180 1560
rect 57220 1545 57235 1560
rect 57275 1545 57290 1560
rect 57330 1545 57345 1560
rect 57385 1545 57400 1560
rect 57440 1545 57455 1560
rect 57495 1545 57510 1560
rect 57550 1545 57565 1560
rect 57605 1545 57620 1560
rect 57660 1545 57675 1560
rect 57715 1545 57730 1560
rect 58190 1545 58205 1560
rect 58245 1545 58260 1560
rect 58300 1545 58315 1560
rect 58355 1545 58370 1560
rect 58410 1545 58425 1560
rect 58465 1545 58480 1560
rect 58520 1545 58535 1560
rect 58575 1545 58590 1560
rect 58630 1545 58645 1560
rect 58685 1545 58700 1560
rect 58740 1545 58755 1560
rect 58795 1545 58810 1560
rect 54955 1535 55005 1545
rect 54955 1515 54960 1535
rect 54980 1530 55005 1535
rect 55595 1535 55645 1545
rect 55595 1530 55620 1535
rect 54980 1515 54985 1530
rect 54955 1505 54985 1515
rect 55615 1515 55620 1530
rect 55640 1515 55645 1535
rect 55615 1505 55645 1515
rect 56035 1535 56085 1545
rect 56035 1515 56040 1535
rect 56060 1530 56085 1535
rect 56675 1535 56825 1545
rect 56675 1530 56740 1535
rect 56060 1515 56065 1530
rect 56035 1505 56065 1515
rect 56735 1515 56740 1530
rect 56760 1530 56825 1535
rect 56975 1535 57125 1545
rect 56975 1530 57040 1535
rect 56760 1515 56765 1530
rect 56735 1505 56765 1515
rect 57035 1515 57040 1530
rect 57060 1530 57125 1535
rect 57715 1535 57765 1545
rect 57715 1530 57740 1535
rect 57060 1515 57065 1530
rect 57035 1505 57065 1515
rect 57735 1515 57740 1530
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 58155 1535 58205 1545
rect 58155 1515 58160 1535
rect 58180 1530 58205 1535
rect 58795 1535 58845 1545
rect 58795 1530 58820 1535
rect 58180 1515 58185 1530
rect 58155 1505 58185 1515
rect 58815 1515 58820 1530
rect 58840 1515 58845 1535
rect 58815 1505 58845 1515
rect 57405 1260 57445 1270
rect 57405 1240 57415 1260
rect 57435 1240 57445 1260
rect 57405 1230 57445 1240
rect 55340 1215 55370 1225
rect 55340 1195 55345 1215
rect 55365 1195 55370 1215
rect 56830 1205 56860 1215
rect 55025 1170 55085 1185
rect 55125 1180 55485 1195
rect 56830 1185 56835 1205
rect 56855 1185 56860 1205
rect 55125 1170 55185 1180
rect 55225 1170 55285 1180
rect 55325 1170 55385 1180
rect 55425 1170 55485 1180
rect 55525 1170 55585 1185
rect 56260 1160 56275 1175
rect 56315 1170 57375 1185
rect 56315 1160 56330 1170
rect 56370 1160 56385 1170
rect 56425 1160 56440 1170
rect 56480 1160 56495 1170
rect 56535 1160 56550 1170
rect 56590 1160 56605 1170
rect 56645 1160 56660 1170
rect 56700 1160 56715 1170
rect 56755 1160 56770 1170
rect 56810 1160 56825 1170
rect 56865 1160 56880 1170
rect 56920 1160 56935 1170
rect 56975 1160 56990 1170
rect 57030 1160 57045 1170
rect 57085 1160 57100 1170
rect 57140 1160 57155 1170
rect 57195 1160 57210 1170
rect 57250 1160 57265 1170
rect 57305 1160 57320 1170
rect 57360 1160 57375 1170
rect 57415 1160 57430 1230
rect 58435 1215 58465 1225
rect 58435 1195 58440 1215
rect 58460 1195 58465 1215
rect 57470 1160 57485 1175
rect 58220 1170 58280 1185
rect 58320 1180 58680 1195
rect 58320 1170 58380 1180
rect 58420 1170 58480 1180
rect 58520 1170 58580 1180
rect 58620 1170 58680 1180
rect 58720 1170 58780 1185
rect 56260 895 56275 910
rect 56315 895 56330 910
rect 56370 895 56385 910
rect 56425 895 56440 910
rect 56480 895 56495 910
rect 56535 895 56550 910
rect 56590 895 56605 910
rect 56645 895 56660 910
rect 56700 895 56715 910
rect 56755 895 56770 910
rect 56810 895 56825 910
rect 56865 895 56880 910
rect 56920 895 56935 910
rect 56975 895 56990 910
rect 57030 895 57045 910
rect 57085 895 57100 910
rect 57140 895 57155 910
rect 57195 895 57210 910
rect 57250 895 57265 910
rect 57305 895 57320 910
rect 57360 895 57375 910
rect 57415 895 57430 910
rect 57470 895 57485 910
rect 56220 885 56275 895
rect 56220 865 56230 885
rect 56250 880 56275 885
rect 57470 885 57525 895
rect 57470 880 57495 885
rect 56250 865 56260 880
rect 56220 855 56260 865
rect 57485 865 57495 880
rect 57515 865 57525 885
rect 57485 855 57525 865
rect 56595 740 56635 750
rect 56595 720 56605 740
rect 56625 720 56635 740
rect 57040 740 57080 750
rect 57040 720 57050 740
rect 57070 720 57080 740
rect 56470 695 56485 710
rect 56525 705 56705 720
rect 57040 710 57080 720
rect 56525 695 56540 705
rect 56580 695 56595 705
rect 56635 695 56650 705
rect 56690 695 56705 705
rect 56745 695 56760 710
rect 56910 695 57210 710
rect 56470 530 56485 545
rect 56525 530 56540 545
rect 56580 530 56595 545
rect 56635 530 56650 545
rect 56690 530 56705 545
rect 56745 530 56760 545
rect 56910 530 57210 545
rect 56435 520 56485 530
rect 56435 500 56440 520
rect 56460 515 56485 520
rect 56745 520 56795 530
rect 56745 515 56770 520
rect 56460 500 56465 515
rect 56435 490 56465 500
rect 56765 500 56770 515
rect 56790 500 56795 520
rect 56765 490 56795 500
rect 55025 455 55085 470
rect 55125 455 55185 470
rect 55225 455 55285 470
rect 55325 455 55385 470
rect 55425 455 55485 470
rect 55525 455 55585 470
rect 58220 455 58280 470
rect 58320 455 58380 470
rect 58420 455 58480 470
rect 58520 455 58580 470
rect 58620 455 58680 470
rect 58720 455 58780 470
rect 54990 445 55085 455
rect 54990 425 54995 445
rect 55015 440 55085 445
rect 55525 445 55620 455
rect 55525 440 55595 445
rect 55015 425 55020 440
rect 54990 415 55020 425
rect 55590 425 55595 440
rect 55615 425 55620 445
rect 55590 415 55620 425
rect 58185 445 58280 455
rect 58185 425 58190 445
rect 58210 440 58280 445
rect 58720 445 58815 455
rect 58720 440 58790 445
rect 58210 425 58215 440
rect 58185 415 58215 425
rect 58785 425 58790 440
rect 58810 425 58815 445
rect 58785 415 58815 425
<< polycont >>
rect 56095 4735 56115 4755
rect 56275 4735 56295 4755
rect 57035 4735 57055 4755
rect 57215 4735 57235 4755
rect 57505 4735 57525 4755
rect 57685 4735 57705 4755
rect 56565 4565 56585 4585
rect 56745 4565 56765 4585
rect 56160 4285 56180 4305
rect 56635 4285 56655 4305
rect 57145 4285 57165 4305
rect 57581 4275 57601 4295
rect 54935 4065 54955 4085
rect 55655 4065 55675 4085
rect 56015 4065 56035 4085
rect 56735 4065 56755 4085
rect 57045 4065 57065 4085
rect 57765 4065 57785 4085
rect 58130 4065 58150 4085
rect 58850 4065 58870 4085
rect 56405 3560 56425 3580
rect 57375 3560 57395 3580
rect 55325 3515 55345 3535
rect 58460 3515 58480 3535
rect 54960 3375 54980 3395
rect 55620 3375 55640 3395
rect 58160 3375 58180 3395
rect 58820 3375 58840 3395
rect 56285 3260 56305 3280
rect 57495 3260 57515 3280
rect 56805 3130 56825 3150
rect 55995 3045 56015 3065
rect 56745 3045 56765 3065
rect 57035 3045 57055 3065
rect 57785 3045 57805 3065
rect 56040 2900 56060 2920
rect 56700 2900 56720 2920
rect 57080 2900 57100 2920
rect 57740 2900 57760 2920
rect 56100 2815 56120 2835
rect 56585 2815 56605 2835
rect 57195 2815 57215 2835
rect 55320 2615 55340 2635
rect 56725 2610 56745 2630
rect 56945 2610 56965 2630
rect 58460 2615 58480 2635
rect 56560 2490 56580 2510
rect 57220 2490 57240 2510
rect 54960 2445 54980 2465
rect 55620 2445 55640 2465
rect 58160 2445 58180 2465
rect 58820 2445 58840 2465
rect 56640 2245 56660 2265
rect 57140 2245 57160 2265
rect 57790 2220 57810 2240
rect 55320 2025 55340 2045
rect 58460 2025 58480 2045
rect 56040 1985 56060 2005
rect 56700 1985 56720 2005
rect 57080 1985 57100 2005
rect 57740 1985 57760 2005
rect 55995 1760 56015 1780
rect 56695 1760 56715 1780
rect 56864 1760 56884 1780
rect 56916 1760 56936 1780
rect 57085 1760 57105 1780
rect 57785 1760 57805 1780
rect 54960 1515 54980 1535
rect 55620 1515 55640 1535
rect 56040 1515 56060 1535
rect 56740 1515 56760 1535
rect 57040 1515 57060 1535
rect 57740 1515 57760 1535
rect 58160 1515 58180 1535
rect 58820 1515 58840 1535
rect 57415 1240 57435 1260
rect 55345 1195 55365 1215
rect 56835 1185 56855 1205
rect 58440 1195 58460 1215
rect 56230 865 56250 885
rect 57495 865 57515 885
rect 56605 720 56625 740
rect 57050 720 57070 740
rect 56440 500 56460 520
rect 56770 500 56790 520
rect 54995 425 55015 445
rect 55595 425 55615 445
rect 58190 425 58210 445
rect 58790 425 58810 445
<< xpolycontact >>
rect 54554 3065 54695 3285
rect 54554 2720 54695 2940
rect 59105 3065 59246 3285
rect 59105 2720 59246 2940
rect 54450 1929 54485 2149
rect 54450 1550 54485 1770
rect 54510 1929 54545 2149
rect 54510 1550 54545 1770
rect 54570 1929 54605 2149
rect 54570 1550 54605 1770
rect 54630 1929 54665 2149
rect 59135 1929 59170 2149
rect 54630 1550 54665 1770
rect 59135 1550 59170 1770
rect 59195 1929 59230 2149
rect 59195 1550 59230 1770
rect 59255 1929 59290 2149
rect 59255 1550 59290 1770
rect 59315 1929 59350 2149
rect 59315 1550 59350 1770
rect 54735 890 54770 1110
rect 54735 423 54770 643
rect 54795 890 54830 1110
rect 54795 423 54830 643
rect 58975 890 59010 1110
rect 58975 423 59010 643
rect 59035 890 59070 1110
rect 59035 423 59070 643
<< ppolyres >>
rect 54554 2940 54695 3065
rect 59105 2940 59246 3065
<< xpolyres >>
rect 54450 1770 54485 1929
rect 54510 1770 54545 1929
rect 54570 1770 54605 1929
rect 54630 1770 54665 1929
rect 59135 1770 59170 1929
rect 59195 1770 59230 1929
rect 59255 1770 59290 1929
rect 59315 1770 59350 1929
rect 54735 643 54770 890
rect 54795 643 54830 890
rect 58975 643 59010 890
rect 59035 643 59070 890
<< locali >>
rect 56085 4755 56125 4765
rect 56085 4735 56095 4755
rect 56115 4735 56125 4755
rect 56085 4725 56125 4735
rect 56265 4755 56305 4765
rect 56265 4735 56275 4755
rect 56295 4735 56305 4755
rect 56265 4725 56305 4735
rect 57025 4755 57065 4765
rect 57025 4735 57035 4755
rect 57055 4735 57065 4755
rect 57025 4725 57065 4735
rect 57205 4755 57245 4765
rect 57205 4735 57215 4755
rect 57235 4735 57245 4755
rect 57205 4725 57245 4735
rect 57495 4755 57535 4765
rect 57495 4735 57505 4755
rect 57525 4735 57535 4755
rect 57495 4725 57535 4735
rect 57675 4755 57715 4765
rect 57675 4735 57685 4755
rect 57705 4735 57715 4755
rect 57675 4725 57715 4735
rect 56050 4695 56120 4705
rect 56050 4375 56055 4695
rect 56075 4375 56095 4695
rect 56115 4375 56120 4695
rect 56050 4365 56120 4375
rect 56150 4695 56180 4705
rect 56150 4375 56155 4695
rect 56175 4375 56180 4695
rect 56150 4365 56180 4375
rect 56210 4695 56240 4705
rect 56210 4375 56215 4695
rect 56235 4375 56240 4695
rect 56210 4365 56240 4375
rect 56270 4695 56340 4705
rect 56270 4375 56275 4695
rect 56295 4375 56315 4695
rect 56335 4375 56340 4695
rect 56990 4695 57060 4705
rect 56555 4585 56595 4595
rect 56555 4565 56565 4585
rect 56585 4565 56595 4585
rect 56555 4555 56595 4565
rect 56735 4585 56775 4595
rect 56735 4565 56745 4585
rect 56765 4565 56775 4585
rect 56735 4555 56775 4565
rect 56270 4365 56340 4375
rect 56520 4525 56590 4535
rect 56520 4375 56525 4525
rect 56545 4375 56565 4525
rect 56585 4375 56590 4525
rect 56520 4365 56590 4375
rect 56620 4525 56650 4535
rect 56620 4375 56625 4525
rect 56645 4375 56650 4525
rect 56620 4365 56650 4375
rect 56680 4525 56710 4535
rect 56680 4375 56685 4525
rect 56705 4375 56710 4525
rect 56680 4365 56710 4375
rect 56740 4525 56810 4535
rect 56740 4375 56745 4525
rect 56765 4375 56785 4525
rect 56805 4375 56810 4525
rect 56740 4365 56810 4375
rect 56990 4375 56995 4695
rect 57015 4375 57035 4695
rect 57055 4375 57060 4695
rect 56990 4365 57060 4375
rect 57090 4695 57120 4705
rect 57090 4375 57095 4695
rect 57115 4375 57120 4695
rect 57090 4365 57120 4375
rect 57150 4695 57180 4705
rect 57150 4375 57155 4695
rect 57175 4375 57180 4695
rect 57150 4365 57180 4375
rect 57210 4695 57280 4705
rect 57210 4375 57215 4695
rect 57235 4375 57255 4695
rect 57275 4375 57280 4695
rect 57210 4365 57280 4375
rect 57460 4695 57530 4705
rect 57460 4375 57465 4695
rect 57485 4375 57505 4695
rect 57525 4375 57530 4695
rect 57460 4365 57530 4375
rect 57560 4695 57590 4705
rect 57560 4375 57565 4695
rect 57585 4375 57590 4695
rect 57560 4365 57590 4375
rect 57620 4695 57650 4705
rect 57620 4375 57625 4695
rect 57645 4375 57650 4695
rect 57620 4365 57650 4375
rect 57680 4695 57750 4705
rect 57680 4375 57685 4695
rect 57705 4375 57725 4695
rect 57745 4375 57750 4695
rect 57680 4365 57750 4375
rect 56150 4305 56190 4315
rect 56150 4285 56160 4305
rect 56180 4285 56190 4305
rect 56150 4275 56190 4285
rect 56630 4305 56660 4315
rect 56630 4285 56635 4305
rect 56655 4285 56660 4305
rect 56630 4275 56660 4285
rect 57140 4305 57170 4315
rect 57140 4285 57145 4305
rect 57165 4285 57170 4305
rect 57140 4275 57170 4285
rect 57576 4295 57606 4305
rect 57576 4275 57581 4295
rect 57601 4275 57606 4295
rect 57576 4265 57606 4275
rect 54930 4085 54960 4095
rect 54930 4065 54935 4085
rect 54955 4065 54960 4085
rect 54930 4055 54960 4065
rect 55650 4085 55680 4095
rect 55650 4065 55655 4085
rect 55675 4065 55680 4085
rect 55650 4055 55680 4065
rect 56010 4085 56040 4095
rect 56010 4065 56015 4085
rect 56035 4065 56040 4085
rect 56010 4055 56040 4065
rect 56730 4085 56760 4095
rect 56730 4065 56735 4085
rect 56755 4065 56760 4085
rect 56730 4055 56760 4065
rect 57040 4085 57070 4095
rect 57040 4065 57045 4085
rect 57065 4065 57070 4085
rect 57040 4055 57070 4065
rect 57760 4085 57790 4095
rect 57760 4065 57765 4085
rect 57785 4065 57790 4085
rect 57760 4055 57790 4065
rect 58125 4085 58155 4095
rect 58125 4065 58130 4085
rect 58150 4065 58155 4085
rect 58125 4055 58155 4065
rect 58845 4085 58875 4095
rect 58845 4065 58850 4085
rect 58870 4065 58875 4085
rect 58845 4055 58875 4065
rect 54890 4025 54960 4035
rect 54890 3705 54895 4025
rect 54915 3705 54935 4025
rect 54955 3705 54960 4025
rect 54890 3695 54960 3705
rect 54990 4025 55020 4035
rect 54990 3705 54995 4025
rect 55015 3705 55020 4025
rect 54990 3695 55020 3705
rect 55050 4025 55080 4035
rect 55050 3705 55055 4025
rect 55075 3705 55080 4025
rect 55050 3695 55080 3705
rect 55110 4025 55140 4035
rect 55110 3705 55115 4025
rect 55135 3705 55140 4025
rect 55110 3695 55140 3705
rect 55170 4025 55200 4035
rect 55170 3705 55175 4025
rect 55195 3705 55200 4025
rect 55170 3695 55200 3705
rect 55230 4025 55260 4035
rect 55230 3705 55235 4025
rect 55255 3705 55260 4025
rect 55230 3695 55260 3705
rect 55290 4025 55320 4035
rect 55290 3705 55295 4025
rect 55315 3705 55320 4025
rect 55290 3695 55320 3705
rect 55350 4025 55380 4035
rect 55350 3705 55355 4025
rect 55375 3705 55380 4025
rect 55350 3695 55380 3705
rect 55410 4025 55440 4035
rect 55410 3705 55415 4025
rect 55435 3705 55440 4025
rect 55410 3695 55440 3705
rect 55470 4025 55500 4035
rect 55470 3705 55475 4025
rect 55495 3705 55500 4025
rect 55470 3695 55500 3705
rect 55530 4025 55560 4035
rect 55530 3705 55535 4025
rect 55555 3705 55560 4025
rect 55530 3695 55560 3705
rect 55590 4025 55620 4035
rect 55590 3705 55595 4025
rect 55615 3705 55620 4025
rect 55590 3695 55620 3705
rect 55650 4025 55720 4035
rect 55650 3705 55655 4025
rect 55675 3705 55695 4025
rect 55715 3705 55720 4025
rect 55650 3695 55720 3705
rect 55970 4025 56040 4035
rect 55970 3705 55975 4025
rect 55995 3705 56015 4025
rect 56035 3705 56040 4025
rect 55970 3695 56040 3705
rect 56070 4025 56100 4035
rect 56070 3705 56075 4025
rect 56095 3705 56100 4025
rect 56070 3695 56100 3705
rect 56130 4025 56160 4035
rect 56130 3705 56135 4025
rect 56155 3705 56160 4025
rect 56130 3695 56160 3705
rect 56190 4025 56220 4035
rect 56190 3705 56195 4025
rect 56215 3705 56220 4025
rect 56190 3695 56220 3705
rect 56250 4025 56280 4035
rect 56250 3705 56255 4025
rect 56275 3705 56280 4025
rect 56250 3695 56280 3705
rect 56310 4025 56340 4035
rect 56310 3705 56315 4025
rect 56335 3705 56340 4025
rect 56310 3695 56340 3705
rect 56370 4025 56400 4035
rect 56370 3705 56375 4025
rect 56395 3705 56400 4025
rect 56370 3695 56400 3705
rect 56430 4025 56460 4035
rect 56430 3705 56435 4025
rect 56455 3705 56460 4025
rect 56430 3695 56460 3705
rect 56490 4025 56520 4035
rect 56490 3705 56495 4025
rect 56515 3705 56520 4025
rect 56490 3695 56520 3705
rect 56550 4025 56580 4035
rect 56550 3705 56555 4025
rect 56575 3705 56580 4025
rect 56550 3695 56580 3705
rect 56610 4025 56640 4035
rect 56610 3705 56615 4025
rect 56635 3705 56640 4025
rect 56610 3695 56640 3705
rect 56670 4025 56700 4035
rect 56670 3705 56675 4025
rect 56695 3705 56700 4025
rect 56670 3695 56700 3705
rect 56730 4025 56800 4035
rect 56730 3705 56735 4025
rect 56755 3705 56775 4025
rect 56795 3705 56800 4025
rect 56730 3695 56800 3705
rect 57000 4025 57070 4035
rect 57000 3705 57005 4025
rect 57025 3705 57045 4025
rect 57065 3705 57070 4025
rect 57000 3695 57070 3705
rect 57100 4025 57130 4035
rect 57100 3705 57105 4025
rect 57125 3705 57130 4025
rect 57100 3695 57130 3705
rect 57160 4025 57190 4035
rect 57160 3705 57165 4025
rect 57185 3705 57190 4025
rect 57160 3695 57190 3705
rect 57220 4025 57250 4035
rect 57220 3705 57225 4025
rect 57245 3705 57250 4025
rect 57220 3695 57250 3705
rect 57280 4025 57310 4035
rect 57280 3705 57285 4025
rect 57305 3705 57310 4025
rect 57280 3695 57310 3705
rect 57340 4025 57370 4035
rect 57340 3705 57345 4025
rect 57365 3705 57370 4025
rect 57340 3695 57370 3705
rect 57400 4025 57430 4035
rect 57400 3705 57405 4025
rect 57425 3705 57430 4025
rect 57400 3695 57430 3705
rect 57460 4025 57490 4035
rect 57460 3705 57465 4025
rect 57485 3705 57490 4025
rect 57460 3695 57490 3705
rect 57520 4025 57550 4035
rect 57520 3705 57525 4025
rect 57545 3705 57550 4025
rect 57520 3695 57550 3705
rect 57580 4025 57610 4035
rect 57580 3705 57585 4025
rect 57605 3705 57610 4025
rect 57580 3695 57610 3705
rect 57640 4025 57670 4035
rect 57640 3705 57645 4025
rect 57665 3705 57670 4025
rect 57640 3695 57670 3705
rect 57700 4025 57730 4035
rect 57700 3705 57705 4025
rect 57725 3705 57730 4025
rect 57700 3695 57730 3705
rect 57760 4025 57830 4035
rect 57760 3705 57765 4025
rect 57785 3705 57805 4025
rect 57825 3705 57830 4025
rect 57760 3695 57830 3705
rect 58085 4025 58155 4035
rect 58085 3705 58090 4025
rect 58110 3705 58130 4025
rect 58150 3705 58155 4025
rect 58085 3695 58155 3705
rect 58185 4025 58215 4035
rect 58185 3705 58190 4025
rect 58210 3705 58215 4025
rect 58185 3695 58215 3705
rect 58245 4025 58275 4035
rect 58245 3705 58250 4025
rect 58270 3705 58275 4025
rect 58245 3695 58275 3705
rect 58305 4025 58335 4035
rect 58305 3705 58310 4025
rect 58330 3705 58335 4025
rect 58305 3695 58335 3705
rect 58365 4025 58395 4035
rect 58365 3705 58370 4025
rect 58390 3705 58395 4025
rect 58365 3695 58395 3705
rect 58425 4025 58455 4035
rect 58425 3705 58430 4025
rect 58450 3705 58455 4025
rect 58425 3695 58455 3705
rect 58485 4025 58515 4035
rect 58485 3705 58490 4025
rect 58510 3705 58515 4025
rect 58485 3695 58515 3705
rect 58545 4025 58575 4035
rect 58545 3705 58550 4025
rect 58570 3705 58575 4025
rect 58545 3695 58575 3705
rect 58605 4025 58635 4035
rect 58605 3705 58610 4025
rect 58630 3705 58635 4025
rect 58605 3695 58635 3705
rect 58665 4025 58695 4035
rect 58665 3705 58670 4025
rect 58690 3705 58695 4025
rect 58665 3695 58695 3705
rect 58725 4025 58755 4035
rect 58725 3705 58730 4025
rect 58750 3705 58755 4025
rect 58725 3695 58755 3705
rect 58785 4025 58815 4035
rect 58785 3705 58790 4025
rect 58810 3705 58815 4025
rect 58785 3695 58815 3705
rect 58845 4025 58915 4035
rect 58845 3705 58850 4025
rect 58870 3705 58890 4025
rect 58910 3705 58915 4025
rect 58845 3695 58915 3705
rect 56395 3580 56435 3590
rect 56395 3560 56405 3580
rect 56425 3560 56435 3580
rect 56395 3550 56435 3560
rect 57365 3580 57405 3590
rect 57365 3560 57375 3580
rect 57395 3560 57405 3580
rect 57365 3550 57405 3560
rect 55315 3535 55355 3545
rect 55315 3515 55325 3535
rect 55345 3515 55355 3535
rect 55315 3505 55355 3515
rect 58450 3535 58490 3545
rect 58450 3515 58460 3535
rect 58480 3515 58490 3535
rect 58450 3505 58490 3515
rect 54955 3395 54985 3405
rect 54955 3375 54960 3395
rect 54980 3375 54985 3395
rect 54955 3365 54985 3375
rect 55615 3395 55645 3405
rect 55615 3375 55620 3395
rect 55640 3375 55645 3395
rect 55615 3365 55645 3375
rect 58155 3395 58185 3405
rect 58155 3375 58160 3395
rect 58180 3375 58185 3395
rect 58155 3365 58185 3375
rect 58815 3395 58845 3405
rect 58815 3375 58820 3395
rect 58840 3375 58845 3395
rect 58815 3365 58845 3375
rect 54915 3335 54985 3345
rect 54554 3315 54695 3325
rect 54554 3295 54560 3315
rect 54580 3295 54615 3315
rect 54635 3295 54670 3315
rect 54690 3295 54695 3315
rect 54554 3285 54695 3295
rect 54915 2765 54920 3335
rect 54940 2765 54960 3335
rect 54980 2765 54985 3335
rect 54915 2755 54985 2765
rect 55010 3335 55040 3345
rect 55010 2765 55015 3335
rect 55035 2765 55040 3335
rect 55010 2755 55040 2765
rect 55065 3335 55095 3345
rect 55065 2765 55070 3335
rect 55090 2765 55095 3335
rect 55065 2755 55095 2765
rect 55120 3335 55150 3345
rect 55120 2765 55125 3335
rect 55145 2765 55150 3335
rect 55120 2755 55150 2765
rect 55175 3335 55205 3345
rect 55175 2765 55180 3335
rect 55200 2765 55205 3335
rect 55175 2755 55205 2765
rect 55230 3335 55260 3345
rect 55230 2765 55235 3335
rect 55255 2765 55260 3335
rect 55230 2755 55260 2765
rect 55285 3335 55315 3345
rect 55285 2765 55290 3335
rect 55310 2765 55315 3335
rect 55285 2755 55315 2765
rect 55340 3335 55370 3345
rect 55340 2765 55345 3335
rect 55365 2765 55370 3335
rect 55340 2755 55370 2765
rect 55395 3335 55425 3345
rect 55395 2765 55400 3335
rect 55420 2765 55425 3335
rect 55395 2755 55425 2765
rect 55450 3335 55480 3345
rect 55450 2765 55455 3335
rect 55475 2765 55480 3335
rect 55450 2755 55480 2765
rect 55505 3335 55535 3345
rect 55505 2765 55510 3335
rect 55530 2765 55535 3335
rect 55505 2755 55535 2765
rect 55560 3335 55590 3345
rect 55560 2765 55565 3335
rect 55585 2765 55590 3335
rect 55560 2755 55590 2765
rect 55615 3335 55685 3345
rect 55615 2765 55620 3335
rect 55640 2765 55660 3335
rect 55680 2765 55685 3335
rect 56240 3340 56310 3350
rect 56240 3320 56245 3340
rect 56265 3320 56285 3340
rect 56305 3320 56310 3340
rect 56240 3310 56310 3320
rect 56335 3340 56365 3350
rect 56335 3320 56340 3340
rect 56360 3320 56365 3340
rect 56335 3310 56365 3320
rect 56390 3340 56420 3350
rect 56390 3320 56395 3340
rect 56415 3320 56420 3340
rect 56390 3310 56420 3320
rect 56445 3340 56475 3350
rect 56445 3320 56450 3340
rect 56470 3320 56475 3340
rect 56445 3310 56475 3320
rect 56500 3340 56530 3350
rect 56500 3320 56505 3340
rect 56525 3320 56530 3340
rect 56500 3310 56530 3320
rect 56555 3340 56585 3350
rect 56555 3320 56560 3340
rect 56580 3320 56585 3340
rect 56555 3310 56585 3320
rect 56610 3340 56640 3350
rect 56610 3320 56615 3340
rect 56635 3320 56640 3340
rect 56610 3310 56640 3320
rect 56665 3340 56695 3350
rect 56665 3320 56670 3340
rect 56690 3320 56695 3340
rect 56665 3310 56695 3320
rect 56720 3340 56750 3350
rect 56720 3320 56725 3340
rect 56745 3320 56750 3340
rect 56720 3310 56750 3320
rect 56775 3340 56805 3350
rect 56775 3320 56780 3340
rect 56800 3320 56805 3340
rect 56775 3310 56805 3320
rect 56830 3340 56860 3350
rect 56830 3320 56835 3340
rect 56855 3320 56860 3340
rect 56830 3310 56860 3320
rect 56885 3340 56915 3350
rect 56885 3320 56890 3340
rect 56910 3320 56915 3340
rect 56885 3310 56915 3320
rect 56940 3340 56970 3350
rect 56940 3320 56945 3340
rect 56965 3320 56970 3340
rect 56940 3310 56970 3320
rect 56995 3340 57025 3350
rect 56995 3320 57000 3340
rect 57020 3320 57025 3340
rect 56995 3310 57025 3320
rect 57050 3340 57080 3350
rect 57050 3320 57055 3340
rect 57075 3320 57080 3340
rect 57050 3310 57080 3320
rect 57105 3340 57135 3350
rect 57105 3320 57110 3340
rect 57130 3320 57135 3340
rect 57105 3310 57135 3320
rect 57160 3340 57190 3350
rect 57160 3320 57165 3340
rect 57185 3320 57190 3340
rect 57160 3310 57190 3320
rect 57215 3340 57245 3350
rect 57215 3320 57220 3340
rect 57240 3320 57245 3340
rect 57215 3310 57245 3320
rect 57270 3340 57300 3350
rect 57270 3320 57275 3340
rect 57295 3320 57300 3340
rect 57270 3310 57300 3320
rect 57325 3340 57355 3350
rect 57325 3320 57330 3340
rect 57350 3320 57355 3340
rect 57325 3310 57355 3320
rect 57380 3340 57410 3350
rect 57380 3320 57385 3340
rect 57405 3320 57410 3340
rect 57380 3310 57410 3320
rect 57435 3340 57465 3350
rect 57435 3320 57440 3340
rect 57460 3320 57465 3340
rect 57435 3310 57465 3320
rect 57490 3340 57560 3350
rect 57490 3320 57495 3340
rect 57515 3320 57535 3340
rect 57555 3320 57560 3340
rect 57490 3310 57560 3320
rect 58115 3335 58185 3345
rect 56280 3280 56310 3290
rect 56280 3260 56285 3280
rect 56305 3260 56310 3280
rect 56280 3250 56310 3260
rect 57490 3280 57520 3290
rect 57490 3260 57495 3280
rect 57515 3260 57520 3280
rect 57490 3250 57520 3260
rect 56795 3150 56835 3160
rect 56795 3130 56805 3150
rect 56825 3130 56835 3150
rect 56795 3120 56835 3130
rect 55990 3065 56020 3075
rect 55990 3045 55995 3065
rect 56015 3045 56020 3065
rect 55990 3035 56020 3045
rect 56740 3065 56770 3075
rect 56740 3045 56745 3065
rect 56765 3045 56770 3065
rect 56740 3035 56770 3045
rect 57030 3065 57060 3075
rect 57030 3045 57035 3065
rect 57055 3045 57060 3065
rect 57030 3035 57060 3045
rect 57780 3065 57810 3075
rect 57780 3045 57785 3065
rect 57805 3045 57810 3065
rect 57780 3035 57810 3045
rect 55995 2980 56065 2990
rect 55995 2960 56000 2980
rect 56020 2960 56040 2980
rect 56060 2960 56065 2980
rect 55995 2950 56065 2960
rect 56090 2980 56120 2990
rect 56090 2960 56095 2980
rect 56115 2960 56120 2980
rect 56090 2950 56120 2960
rect 56145 2980 56175 2990
rect 56145 2960 56150 2980
rect 56170 2960 56175 2980
rect 56145 2950 56175 2960
rect 56200 2980 56230 2990
rect 56200 2960 56205 2980
rect 56225 2960 56230 2980
rect 56200 2950 56230 2960
rect 56255 2980 56285 2990
rect 56255 2960 56260 2980
rect 56280 2960 56285 2980
rect 56255 2950 56285 2960
rect 56310 2980 56340 2990
rect 56310 2960 56315 2980
rect 56335 2960 56340 2980
rect 56310 2950 56340 2960
rect 56365 2980 56395 2990
rect 56365 2960 56370 2980
rect 56390 2960 56395 2980
rect 56365 2950 56395 2960
rect 56420 2980 56450 2990
rect 56420 2960 56425 2980
rect 56445 2960 56450 2980
rect 56420 2950 56450 2960
rect 56475 2980 56505 2990
rect 56475 2960 56480 2980
rect 56500 2960 56505 2980
rect 56475 2950 56505 2960
rect 56530 2980 56560 2990
rect 56530 2960 56535 2980
rect 56555 2960 56560 2980
rect 56530 2950 56560 2960
rect 56585 2980 56615 2990
rect 56585 2960 56590 2980
rect 56610 2960 56615 2980
rect 56585 2950 56615 2960
rect 56640 2980 56670 2990
rect 56640 2960 56645 2980
rect 56665 2960 56670 2980
rect 56640 2950 56670 2960
rect 56695 2980 56765 2990
rect 56695 2960 56700 2980
rect 56720 2960 56740 2980
rect 56760 2960 56765 2980
rect 56695 2950 56765 2960
rect 57035 2980 57105 2990
rect 57035 2960 57040 2980
rect 57060 2960 57080 2980
rect 57100 2960 57105 2980
rect 57035 2950 57105 2960
rect 57130 2980 57160 2990
rect 57130 2960 57135 2980
rect 57155 2960 57160 2980
rect 57130 2950 57160 2960
rect 57185 2980 57215 2990
rect 57185 2960 57190 2980
rect 57210 2960 57215 2980
rect 57185 2950 57215 2960
rect 57240 2980 57270 2990
rect 57240 2960 57245 2980
rect 57265 2960 57270 2980
rect 57240 2950 57270 2960
rect 57295 2980 57325 2990
rect 57295 2960 57300 2980
rect 57320 2960 57325 2980
rect 57295 2950 57325 2960
rect 57350 2980 57380 2990
rect 57350 2960 57355 2980
rect 57375 2960 57380 2980
rect 57350 2950 57380 2960
rect 57405 2980 57435 2990
rect 57405 2960 57410 2980
rect 57430 2960 57435 2980
rect 57405 2950 57435 2960
rect 57460 2980 57490 2990
rect 57460 2960 57465 2980
rect 57485 2960 57490 2980
rect 57460 2950 57490 2960
rect 57515 2980 57545 2990
rect 57515 2960 57520 2980
rect 57540 2960 57545 2980
rect 57515 2950 57545 2960
rect 57570 2980 57600 2990
rect 57570 2960 57575 2980
rect 57595 2960 57600 2980
rect 57570 2950 57600 2960
rect 57625 2980 57655 2990
rect 57625 2960 57630 2980
rect 57650 2960 57655 2980
rect 57625 2950 57655 2960
rect 57680 2980 57710 2990
rect 57680 2960 57685 2980
rect 57705 2960 57710 2980
rect 57680 2950 57710 2960
rect 57735 2980 57805 2990
rect 57735 2960 57740 2980
rect 57760 2960 57780 2980
rect 57800 2960 57805 2980
rect 57735 2950 57805 2960
rect 56035 2920 56065 2930
rect 56035 2900 56040 2920
rect 56060 2900 56065 2920
rect 56035 2890 56065 2900
rect 56695 2920 56725 2930
rect 56695 2900 56700 2920
rect 56720 2900 56725 2920
rect 56695 2890 56725 2900
rect 57075 2920 57105 2930
rect 57075 2900 57080 2920
rect 57100 2900 57105 2920
rect 57075 2890 57105 2900
rect 57735 2920 57765 2930
rect 57735 2900 57740 2920
rect 57760 2900 57765 2920
rect 57735 2890 57765 2900
rect 56095 2835 56125 2845
rect 56095 2815 56100 2835
rect 56120 2815 56125 2835
rect 56095 2805 56125 2815
rect 56580 2835 56610 2845
rect 56580 2815 56585 2835
rect 56605 2815 56610 2835
rect 56580 2805 56610 2815
rect 57190 2835 57220 2845
rect 57190 2815 57195 2835
rect 57215 2815 57220 2835
rect 57190 2805 57220 2815
rect 55615 2755 55685 2765
rect 58115 2765 58120 3335
rect 58140 2765 58160 3335
rect 58180 2765 58185 3335
rect 58115 2755 58185 2765
rect 58210 3335 58240 3345
rect 58210 2765 58215 3335
rect 58235 2765 58240 3335
rect 58210 2755 58240 2765
rect 58265 3335 58295 3345
rect 58265 2765 58270 3335
rect 58290 2765 58295 3335
rect 58265 2755 58295 2765
rect 58320 3335 58350 3345
rect 58320 2765 58325 3335
rect 58345 2765 58350 3335
rect 58320 2755 58350 2765
rect 58375 3335 58405 3345
rect 58375 2765 58380 3335
rect 58400 2765 58405 3335
rect 58375 2755 58405 2765
rect 58430 3335 58460 3345
rect 58430 2765 58435 3335
rect 58455 2765 58460 3335
rect 58430 2755 58460 2765
rect 58485 3335 58515 3345
rect 58485 2765 58490 3335
rect 58510 2765 58515 3335
rect 58485 2755 58515 2765
rect 58540 3335 58570 3345
rect 58540 2765 58545 3335
rect 58565 2765 58570 3335
rect 58540 2755 58570 2765
rect 58595 3335 58625 3345
rect 58595 2765 58600 3335
rect 58620 2765 58625 3335
rect 58595 2755 58625 2765
rect 58650 3335 58680 3345
rect 58650 2765 58655 3335
rect 58675 2765 58680 3335
rect 58650 2755 58680 2765
rect 58705 3335 58735 3345
rect 58705 2765 58710 3335
rect 58730 2765 58735 3335
rect 58705 2755 58735 2765
rect 58760 3335 58790 3345
rect 58760 2765 58765 3335
rect 58785 2765 58790 3335
rect 58760 2755 58790 2765
rect 58815 3335 58885 3345
rect 58815 2765 58820 3335
rect 58840 2765 58860 3335
rect 58880 2765 58885 3335
rect 59105 3315 59246 3325
rect 59105 3295 59110 3315
rect 59130 3295 59165 3315
rect 59185 3295 59220 3315
rect 59240 3295 59246 3315
rect 59105 3285 59246 3295
rect 58815 2755 58885 2765
rect 54554 2710 54695 2720
rect 54554 2690 54560 2710
rect 54580 2690 54615 2710
rect 54635 2690 54670 2710
rect 54690 2690 54695 2710
rect 54554 2680 54695 2690
rect 59105 2710 59246 2720
rect 59105 2690 59110 2710
rect 59130 2690 59165 2710
rect 59185 2690 59220 2710
rect 59240 2690 59246 2710
rect 59105 2680 59246 2690
rect 55310 2635 55350 2645
rect 55310 2615 55320 2635
rect 55340 2615 55350 2635
rect 55310 2605 55350 2615
rect 56715 2630 56755 2640
rect 56715 2610 56725 2630
rect 56745 2610 56755 2630
rect 56715 2600 56755 2610
rect 56935 2630 56975 2640
rect 56935 2610 56945 2630
rect 56965 2610 56975 2630
rect 56935 2600 56975 2610
rect 58450 2635 58490 2645
rect 58450 2615 58460 2635
rect 58480 2615 58490 2635
rect 58450 2605 58490 2615
rect 56515 2570 56585 2580
rect 56515 2550 56520 2570
rect 56540 2550 56560 2570
rect 56580 2550 56585 2570
rect 56515 2540 56585 2550
rect 56610 2570 56640 2580
rect 56610 2550 56615 2570
rect 56635 2550 56640 2570
rect 56610 2540 56640 2550
rect 56665 2570 56695 2580
rect 56665 2550 56670 2570
rect 56690 2550 56695 2570
rect 56665 2540 56695 2550
rect 56720 2570 56750 2580
rect 56720 2550 56725 2570
rect 56745 2550 56750 2570
rect 56720 2540 56750 2550
rect 56775 2570 56805 2580
rect 56775 2550 56780 2570
rect 56800 2550 56805 2570
rect 56775 2540 56805 2550
rect 56830 2570 56860 2580
rect 56830 2550 56835 2570
rect 56855 2550 56860 2570
rect 56830 2540 56860 2550
rect 56885 2570 56915 2580
rect 56885 2550 56890 2570
rect 56910 2550 56915 2570
rect 56885 2540 56915 2550
rect 56940 2570 56970 2580
rect 56940 2550 56945 2570
rect 56965 2550 56970 2570
rect 56940 2540 56970 2550
rect 56995 2570 57025 2580
rect 56995 2550 57000 2570
rect 57020 2550 57025 2570
rect 56995 2540 57025 2550
rect 57050 2570 57080 2580
rect 57050 2550 57055 2570
rect 57075 2550 57080 2570
rect 57050 2540 57080 2550
rect 57105 2570 57135 2580
rect 57105 2550 57110 2570
rect 57130 2550 57135 2570
rect 57105 2540 57135 2550
rect 57160 2570 57190 2580
rect 57160 2550 57165 2570
rect 57185 2550 57190 2570
rect 57160 2540 57190 2550
rect 57215 2570 57285 2580
rect 57215 2550 57220 2570
rect 57240 2550 57260 2570
rect 57280 2550 57285 2570
rect 57215 2540 57285 2550
rect 56550 2510 56590 2520
rect 56550 2490 56560 2510
rect 56580 2490 56590 2510
rect 56550 2480 56590 2490
rect 57210 2510 57250 2520
rect 57210 2490 57220 2510
rect 57240 2490 57250 2510
rect 57210 2480 57250 2490
rect 54955 2465 54985 2475
rect 54955 2445 54960 2465
rect 54980 2445 54985 2465
rect 54955 2435 54985 2445
rect 55615 2465 55645 2475
rect 55615 2445 55620 2465
rect 55640 2445 55645 2465
rect 55615 2435 55645 2445
rect 58155 2465 58185 2475
rect 58155 2445 58160 2465
rect 58180 2445 58185 2465
rect 58155 2435 58185 2445
rect 58815 2465 58845 2475
rect 58815 2445 58820 2465
rect 58840 2445 58845 2465
rect 58815 2435 58845 2445
rect 54915 2405 54985 2415
rect 54915 2235 54920 2405
rect 54940 2235 54960 2405
rect 54980 2235 54985 2405
rect 54915 2225 54985 2235
rect 55010 2405 55040 2415
rect 55010 2235 55015 2405
rect 55035 2235 55040 2405
rect 55010 2225 55040 2235
rect 55065 2405 55095 2415
rect 55065 2235 55070 2405
rect 55090 2235 55095 2405
rect 55065 2225 55095 2235
rect 55120 2405 55150 2415
rect 55120 2235 55125 2405
rect 55145 2235 55150 2405
rect 55120 2225 55150 2235
rect 55175 2405 55205 2415
rect 55175 2235 55180 2405
rect 55200 2235 55205 2405
rect 55175 2225 55205 2235
rect 55230 2405 55260 2415
rect 55230 2235 55235 2405
rect 55255 2235 55260 2405
rect 55230 2225 55260 2235
rect 55285 2405 55315 2415
rect 55285 2235 55290 2405
rect 55310 2235 55315 2405
rect 55285 2225 55315 2235
rect 55340 2405 55370 2415
rect 55340 2235 55345 2405
rect 55365 2235 55370 2405
rect 55340 2225 55370 2235
rect 55395 2405 55425 2415
rect 55395 2235 55400 2405
rect 55420 2235 55425 2405
rect 55395 2225 55425 2235
rect 55450 2405 55480 2415
rect 55450 2235 55455 2405
rect 55475 2235 55480 2405
rect 55450 2225 55480 2235
rect 55505 2405 55535 2415
rect 55505 2235 55510 2405
rect 55530 2235 55535 2405
rect 55505 2225 55535 2235
rect 55560 2405 55590 2415
rect 55560 2235 55565 2405
rect 55585 2235 55590 2405
rect 55560 2225 55590 2235
rect 55615 2405 55685 2415
rect 55615 2235 55620 2405
rect 55640 2235 55660 2405
rect 55680 2235 55685 2405
rect 58115 2405 58185 2415
rect 56635 2265 56665 2275
rect 56635 2245 56640 2265
rect 56660 2245 56665 2265
rect 56635 2235 56665 2245
rect 57135 2265 57165 2275
rect 57135 2245 57140 2265
rect 57160 2245 57165 2265
rect 57135 2235 57165 2245
rect 57785 2240 57815 2250
rect 55615 2225 55685 2235
rect 57785 2220 57790 2240
rect 57810 2220 57815 2240
rect 58115 2235 58120 2405
rect 58140 2235 58160 2405
rect 58180 2235 58185 2405
rect 58115 2225 58185 2235
rect 58210 2405 58240 2415
rect 58210 2235 58215 2405
rect 58235 2235 58240 2405
rect 58210 2225 58240 2235
rect 58265 2405 58295 2415
rect 58265 2235 58270 2405
rect 58290 2235 58295 2405
rect 58265 2225 58295 2235
rect 58320 2405 58350 2415
rect 58320 2235 58325 2405
rect 58345 2235 58350 2405
rect 58320 2225 58350 2235
rect 58375 2405 58405 2415
rect 58375 2235 58380 2405
rect 58400 2235 58405 2405
rect 58375 2225 58405 2235
rect 58430 2405 58460 2415
rect 58430 2235 58435 2405
rect 58455 2235 58460 2405
rect 58430 2225 58460 2235
rect 58485 2405 58515 2415
rect 58485 2235 58490 2405
rect 58510 2235 58515 2405
rect 58485 2225 58515 2235
rect 58540 2405 58570 2415
rect 58540 2235 58545 2405
rect 58565 2235 58570 2405
rect 58540 2225 58570 2235
rect 58595 2405 58625 2415
rect 58595 2235 58600 2405
rect 58620 2235 58625 2405
rect 58595 2225 58625 2235
rect 58650 2405 58680 2415
rect 58650 2235 58655 2405
rect 58675 2235 58680 2405
rect 58650 2225 58680 2235
rect 58705 2405 58735 2415
rect 58705 2235 58710 2405
rect 58730 2235 58735 2405
rect 58705 2225 58735 2235
rect 58760 2405 58790 2415
rect 58760 2235 58765 2405
rect 58785 2235 58790 2405
rect 58760 2225 58790 2235
rect 58815 2405 58885 2415
rect 58815 2235 58820 2405
rect 58840 2235 58860 2405
rect 58880 2235 58885 2405
rect 58815 2225 58885 2235
rect 57785 2210 57815 2220
rect 55060 2195 55100 2205
rect 54450 2166 54665 2186
rect 54450 2149 54485 2166
rect 54630 2149 54665 2166
rect 55060 2175 55070 2195
rect 55090 2175 55100 2195
rect 55060 2165 55100 2175
rect 55170 2195 55210 2205
rect 55170 2175 55180 2195
rect 55200 2175 55210 2195
rect 55170 2165 55210 2175
rect 55280 2195 55320 2205
rect 55280 2175 55290 2195
rect 55310 2175 55320 2195
rect 55280 2165 55320 2175
rect 55390 2195 55430 2205
rect 55390 2175 55400 2195
rect 55420 2175 55430 2195
rect 55390 2165 55430 2175
rect 55500 2195 55540 2205
rect 55500 2175 55510 2195
rect 55530 2175 55540 2195
rect 58260 2195 58300 2205
rect 58260 2175 58270 2195
rect 58290 2175 58300 2195
rect 55500 2165 55540 2175
rect 55995 2165 56065 2175
rect 54545 2099 54570 2149
rect 55310 2045 55350 2055
rect 55310 2025 55320 2045
rect 55340 2025 55350 2045
rect 55995 2045 56000 2165
rect 56020 2045 56040 2165
rect 56060 2045 56065 2165
rect 55995 2035 56065 2045
rect 56090 2165 56120 2175
rect 56090 2045 56095 2165
rect 56115 2045 56120 2165
rect 56090 2035 56120 2045
rect 56145 2165 56175 2175
rect 56145 2045 56150 2165
rect 56170 2045 56175 2165
rect 56145 2035 56175 2045
rect 56200 2165 56230 2175
rect 56200 2045 56205 2165
rect 56225 2045 56230 2165
rect 56200 2035 56230 2045
rect 56255 2165 56285 2175
rect 56255 2045 56260 2165
rect 56280 2045 56285 2165
rect 56255 2035 56285 2045
rect 56310 2165 56340 2175
rect 56310 2045 56315 2165
rect 56335 2045 56340 2165
rect 56310 2035 56340 2045
rect 56365 2165 56395 2175
rect 56365 2045 56370 2165
rect 56390 2045 56395 2165
rect 56365 2035 56395 2045
rect 56420 2165 56450 2175
rect 56420 2045 56425 2165
rect 56445 2045 56450 2165
rect 56420 2035 56450 2045
rect 56475 2165 56505 2175
rect 56475 2045 56480 2165
rect 56500 2045 56505 2165
rect 56475 2035 56505 2045
rect 56530 2165 56560 2175
rect 56530 2045 56535 2165
rect 56555 2045 56560 2165
rect 56530 2035 56560 2045
rect 56585 2165 56615 2175
rect 56585 2045 56590 2165
rect 56610 2045 56615 2165
rect 56585 2035 56615 2045
rect 56640 2165 56670 2175
rect 56640 2045 56645 2165
rect 56665 2045 56670 2165
rect 56640 2035 56670 2045
rect 56695 2165 56765 2175
rect 56695 2045 56700 2165
rect 56720 2045 56740 2165
rect 56760 2045 56765 2165
rect 56695 2035 56765 2045
rect 57035 2165 57105 2175
rect 57035 2045 57040 2165
rect 57060 2045 57080 2165
rect 57100 2045 57105 2165
rect 57035 2035 57105 2045
rect 57130 2165 57160 2175
rect 57130 2045 57135 2165
rect 57155 2045 57160 2165
rect 57130 2035 57160 2045
rect 57185 2165 57215 2175
rect 57185 2045 57190 2165
rect 57210 2045 57215 2165
rect 57185 2035 57215 2045
rect 57240 2165 57270 2175
rect 57240 2045 57245 2165
rect 57265 2045 57270 2165
rect 57240 2035 57270 2045
rect 57295 2165 57325 2175
rect 57295 2045 57300 2165
rect 57320 2045 57325 2165
rect 57295 2035 57325 2045
rect 57350 2165 57380 2175
rect 57350 2045 57355 2165
rect 57375 2045 57380 2165
rect 57350 2035 57380 2045
rect 57405 2165 57435 2175
rect 57405 2045 57410 2165
rect 57430 2045 57435 2165
rect 57405 2035 57435 2045
rect 57460 2165 57490 2175
rect 57460 2045 57465 2165
rect 57485 2045 57490 2165
rect 57460 2035 57490 2045
rect 57515 2165 57545 2175
rect 57515 2045 57520 2165
rect 57540 2045 57545 2165
rect 57515 2035 57545 2045
rect 57570 2165 57600 2175
rect 57570 2045 57575 2165
rect 57595 2045 57600 2165
rect 57570 2035 57600 2045
rect 57625 2165 57655 2175
rect 57625 2045 57630 2165
rect 57650 2045 57655 2165
rect 57625 2035 57655 2045
rect 57680 2165 57710 2175
rect 57680 2045 57685 2165
rect 57705 2045 57710 2165
rect 57680 2035 57710 2045
rect 57735 2165 57805 2175
rect 58260 2165 58300 2175
rect 58370 2195 58410 2205
rect 58370 2175 58380 2195
rect 58400 2175 58410 2195
rect 58370 2165 58410 2175
rect 58480 2195 58520 2205
rect 58480 2175 58490 2195
rect 58510 2175 58520 2195
rect 58480 2165 58520 2175
rect 58590 2195 58630 2205
rect 58590 2175 58600 2195
rect 58620 2175 58630 2195
rect 58590 2165 58630 2175
rect 58700 2195 58740 2205
rect 58700 2175 58710 2195
rect 58730 2175 58740 2195
rect 58700 2165 58740 2175
rect 59135 2166 59350 2186
rect 57735 2045 57740 2165
rect 57760 2045 57780 2165
rect 57800 2045 57805 2165
rect 59135 2149 59170 2166
rect 59315 2149 59350 2166
rect 57735 2035 57805 2045
rect 58450 2045 58490 2055
rect 55310 2015 55350 2025
rect 56035 2005 56065 2035
rect 56035 1985 56040 2005
rect 56060 1985 56065 2005
rect 56035 1975 56065 1985
rect 56695 2005 56725 2015
rect 56695 1985 56700 2005
rect 56720 1985 56725 2005
rect 56695 1975 56725 1985
rect 57075 2005 57105 2015
rect 57075 1985 57080 2005
rect 57100 1985 57105 2005
rect 57075 1975 57105 1985
rect 57735 2005 57765 2035
rect 58450 2025 58460 2045
rect 58480 2025 58490 2045
rect 58450 2015 58490 2025
rect 57735 1985 57740 2005
rect 57760 1985 57765 2005
rect 57735 1975 57765 1985
rect 59230 2099 59255 2149
rect 54915 1845 54985 1855
rect 54450 1540 54485 1550
rect 54450 1515 54455 1540
rect 54480 1515 54485 1540
rect 54450 1505 54485 1515
rect 54510 1540 54545 1550
rect 54510 1515 54515 1540
rect 54540 1515 54545 1540
rect 54510 1505 54545 1515
rect 54570 1540 54605 1550
rect 54570 1515 54575 1540
rect 54600 1515 54605 1540
rect 54570 1505 54605 1515
rect 54915 1575 54920 1845
rect 54940 1575 54960 1845
rect 54980 1575 54985 1845
rect 54915 1565 54985 1575
rect 55010 1845 55040 1855
rect 55010 1575 55015 1845
rect 55035 1575 55040 1845
rect 55010 1565 55040 1575
rect 55065 1845 55095 1855
rect 55065 1575 55070 1845
rect 55090 1575 55095 1845
rect 55065 1565 55095 1575
rect 55120 1845 55150 1855
rect 55120 1575 55125 1845
rect 55145 1575 55150 1845
rect 55120 1565 55150 1575
rect 55175 1845 55205 1855
rect 55175 1575 55180 1845
rect 55200 1575 55205 1845
rect 55175 1565 55205 1575
rect 55230 1845 55260 1855
rect 55230 1575 55235 1845
rect 55255 1575 55260 1845
rect 55230 1565 55260 1575
rect 55285 1845 55315 1855
rect 55285 1575 55290 1845
rect 55310 1575 55315 1845
rect 55285 1565 55315 1575
rect 55340 1845 55370 1855
rect 55340 1575 55345 1845
rect 55365 1575 55370 1845
rect 55340 1565 55370 1575
rect 55395 1845 55425 1855
rect 55395 1575 55400 1845
rect 55420 1575 55425 1845
rect 55395 1565 55425 1575
rect 55450 1845 55480 1855
rect 55450 1575 55455 1845
rect 55475 1575 55480 1845
rect 55450 1565 55480 1575
rect 55505 1845 55535 1855
rect 55505 1575 55510 1845
rect 55530 1575 55535 1845
rect 55505 1565 55535 1575
rect 55560 1845 55590 1855
rect 55560 1575 55565 1845
rect 55585 1575 55590 1845
rect 55560 1565 55590 1575
rect 55615 1845 55685 1855
rect 55615 1575 55620 1845
rect 55640 1575 55660 1845
rect 55680 1575 55685 1845
rect 58115 1845 58185 1855
rect 55990 1780 56020 1790
rect 55990 1760 55995 1780
rect 56015 1760 56020 1780
rect 55990 1750 56020 1760
rect 56690 1780 56720 1790
rect 56690 1760 56695 1780
rect 56715 1760 56720 1780
rect 56690 1750 56720 1760
rect 56859 1780 56889 1790
rect 56859 1760 56864 1780
rect 56884 1760 56889 1780
rect 56859 1750 56889 1760
rect 56911 1780 56941 1790
rect 56911 1760 56916 1780
rect 56936 1760 56941 1780
rect 56911 1750 56941 1760
rect 57080 1780 57110 1790
rect 57080 1760 57085 1780
rect 57105 1760 57110 1780
rect 57080 1750 57110 1760
rect 57780 1780 57810 1790
rect 57780 1760 57785 1780
rect 57805 1760 57810 1780
rect 57780 1750 57810 1760
rect 55615 1565 55685 1575
rect 55995 1695 56065 1705
rect 55995 1575 56000 1695
rect 56020 1575 56040 1695
rect 56060 1575 56065 1695
rect 55995 1565 56065 1575
rect 56090 1695 56120 1705
rect 56090 1575 56095 1695
rect 56115 1575 56120 1695
rect 56090 1565 56120 1575
rect 56145 1695 56175 1705
rect 56145 1575 56150 1695
rect 56170 1575 56175 1695
rect 56145 1565 56175 1575
rect 56200 1695 56230 1705
rect 56200 1575 56205 1695
rect 56225 1575 56230 1695
rect 56200 1565 56230 1575
rect 56255 1695 56285 1705
rect 56255 1575 56260 1695
rect 56280 1575 56285 1695
rect 56255 1565 56285 1575
rect 56310 1695 56340 1705
rect 56310 1575 56315 1695
rect 56335 1575 56340 1695
rect 56310 1565 56340 1575
rect 56365 1695 56395 1705
rect 56365 1575 56370 1695
rect 56390 1575 56395 1695
rect 56365 1565 56395 1575
rect 56420 1695 56450 1705
rect 56420 1575 56425 1695
rect 56445 1575 56450 1695
rect 56420 1565 56450 1575
rect 56475 1695 56505 1705
rect 56475 1575 56480 1695
rect 56500 1575 56505 1695
rect 56475 1565 56505 1575
rect 56530 1695 56560 1705
rect 56530 1575 56535 1695
rect 56555 1575 56560 1695
rect 56530 1565 56560 1575
rect 56585 1695 56615 1705
rect 56585 1575 56590 1695
rect 56610 1575 56615 1695
rect 56585 1565 56615 1575
rect 56640 1695 56670 1705
rect 56640 1575 56645 1695
rect 56665 1575 56670 1695
rect 56640 1565 56670 1575
rect 56695 1695 56805 1705
rect 56695 1575 56700 1695
rect 56720 1575 56740 1695
rect 56760 1575 56780 1695
rect 56800 1575 56805 1695
rect 56695 1565 56805 1575
rect 56830 1695 56860 1705
rect 56830 1575 56835 1695
rect 56855 1575 56860 1695
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1575 56890 1695
rect 56910 1575 56915 1695
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1575 56945 1695
rect 56965 1575 56970 1695
rect 56940 1565 56970 1575
rect 56995 1695 57105 1705
rect 56995 1575 57000 1695
rect 57020 1575 57040 1695
rect 57060 1575 57080 1695
rect 57100 1575 57105 1695
rect 56995 1565 57105 1575
rect 57130 1695 57160 1705
rect 57130 1575 57135 1695
rect 57155 1575 57160 1695
rect 57130 1565 57160 1575
rect 57185 1695 57215 1705
rect 57185 1575 57190 1695
rect 57210 1575 57215 1695
rect 57185 1565 57215 1575
rect 57240 1695 57270 1705
rect 57240 1575 57245 1695
rect 57265 1575 57270 1695
rect 57240 1565 57270 1575
rect 57295 1695 57325 1705
rect 57295 1575 57300 1695
rect 57320 1575 57325 1695
rect 57295 1565 57325 1575
rect 57350 1695 57380 1705
rect 57350 1575 57355 1695
rect 57375 1575 57380 1695
rect 57350 1565 57380 1575
rect 57405 1695 57435 1705
rect 57405 1575 57410 1695
rect 57430 1575 57435 1695
rect 57405 1565 57435 1575
rect 57460 1695 57490 1705
rect 57460 1575 57465 1695
rect 57485 1575 57490 1695
rect 57460 1565 57490 1575
rect 57515 1695 57545 1705
rect 57515 1575 57520 1695
rect 57540 1575 57545 1695
rect 57515 1565 57545 1575
rect 57570 1695 57600 1705
rect 57570 1575 57575 1695
rect 57595 1575 57600 1695
rect 57570 1565 57600 1575
rect 57625 1695 57655 1705
rect 57625 1575 57630 1695
rect 57650 1575 57655 1695
rect 57625 1565 57655 1575
rect 57680 1695 57710 1705
rect 57680 1575 57685 1695
rect 57705 1575 57710 1695
rect 57680 1565 57710 1575
rect 57735 1695 57805 1705
rect 57735 1575 57740 1695
rect 57760 1575 57780 1695
rect 57800 1575 57805 1695
rect 57735 1565 57805 1575
rect 58115 1575 58120 1845
rect 58140 1575 58160 1845
rect 58180 1575 58185 1845
rect 58115 1565 58185 1575
rect 58210 1845 58240 1855
rect 58210 1575 58215 1845
rect 58235 1575 58240 1845
rect 58210 1565 58240 1575
rect 58265 1845 58295 1855
rect 58265 1575 58270 1845
rect 58290 1575 58295 1845
rect 58265 1565 58295 1575
rect 58320 1845 58350 1855
rect 58320 1575 58325 1845
rect 58345 1575 58350 1845
rect 58320 1565 58350 1575
rect 58375 1845 58405 1855
rect 58375 1575 58380 1845
rect 58400 1575 58405 1845
rect 58375 1565 58405 1575
rect 58430 1845 58460 1855
rect 58430 1575 58435 1845
rect 58455 1575 58460 1845
rect 58430 1565 58460 1575
rect 58485 1845 58515 1855
rect 58485 1575 58490 1845
rect 58510 1575 58515 1845
rect 58485 1565 58515 1575
rect 58540 1845 58570 1855
rect 58540 1575 58545 1845
rect 58565 1575 58570 1845
rect 58540 1565 58570 1575
rect 58595 1845 58625 1855
rect 58595 1575 58600 1845
rect 58620 1575 58625 1845
rect 58595 1565 58625 1575
rect 58650 1845 58680 1855
rect 58650 1575 58655 1845
rect 58675 1575 58680 1845
rect 58650 1565 58680 1575
rect 58705 1845 58735 1855
rect 58705 1575 58710 1845
rect 58730 1575 58735 1845
rect 58705 1565 58735 1575
rect 58760 1845 58790 1855
rect 58760 1575 58765 1845
rect 58785 1575 58790 1845
rect 58760 1565 58790 1575
rect 58815 1845 58885 1855
rect 58815 1575 58820 1845
rect 58840 1575 58860 1845
rect 58880 1575 58885 1845
rect 58815 1565 58885 1575
rect 54630 1540 54665 1550
rect 54630 1515 54635 1540
rect 54660 1515 54665 1540
rect 54630 1505 54665 1515
rect 54955 1535 54985 1545
rect 54955 1515 54960 1535
rect 54980 1515 54985 1535
rect 54955 1505 54985 1515
rect 55615 1535 55645 1545
rect 55615 1515 55620 1535
rect 55640 1515 55645 1535
rect 55615 1505 55645 1515
rect 56035 1535 56065 1545
rect 56035 1515 56040 1535
rect 56060 1515 56065 1535
rect 56035 1505 56065 1515
rect 56735 1535 56765 1545
rect 56735 1515 56740 1535
rect 56760 1515 56765 1535
rect 56735 1505 56765 1515
rect 57035 1535 57065 1545
rect 57035 1515 57040 1535
rect 57060 1515 57065 1535
rect 57035 1505 57065 1515
rect 57735 1535 57765 1565
rect 57735 1515 57740 1535
rect 57760 1515 57765 1535
rect 57735 1505 57765 1515
rect 58155 1535 58185 1545
rect 58155 1515 58160 1535
rect 58180 1515 58185 1535
rect 58155 1505 58185 1515
rect 58815 1535 58845 1545
rect 58815 1515 58820 1535
rect 58840 1515 58845 1535
rect 58815 1505 58845 1515
rect 59135 1540 59170 1550
rect 59135 1515 59140 1540
rect 59165 1515 59170 1540
rect 59135 1505 59170 1515
rect 59195 1540 59230 1550
rect 59195 1515 59200 1540
rect 59225 1515 59230 1540
rect 59195 1505 59230 1515
rect 59255 1540 59290 1550
rect 59255 1515 59260 1540
rect 59285 1515 59290 1540
rect 59255 1505 59290 1515
rect 59315 1540 59350 1550
rect 59315 1515 59320 1540
rect 59345 1515 59350 1540
rect 59315 1505 59350 1515
rect 57405 1260 57445 1270
rect 57405 1240 57415 1260
rect 57435 1240 57445 1260
rect 57405 1230 57445 1240
rect 55340 1215 55370 1225
rect 58435 1215 58465 1225
rect 55340 1195 55345 1215
rect 55365 1195 55370 1215
rect 55340 1185 55370 1195
rect 56830 1205 56860 1215
rect 56830 1185 56835 1205
rect 56855 1185 56860 1205
rect 58435 1195 58440 1215
rect 58460 1195 58465 1215
rect 58435 1185 58465 1195
rect 56830 1175 56860 1185
rect 54950 1155 55020 1165
rect 54735 1145 54770 1155
rect 54735 1120 54740 1145
rect 54765 1120 54770 1145
rect 54735 1110 54770 1120
rect 54795 1145 54830 1155
rect 54795 1120 54800 1145
rect 54825 1120 54830 1145
rect 54795 1110 54830 1120
rect 54770 423 54795 473
rect 54950 485 54955 1155
rect 54975 485 54995 1155
rect 55015 485 55020 1155
rect 54950 475 55020 485
rect 55090 1155 55120 1165
rect 55090 485 55095 1155
rect 55115 485 55120 1155
rect 55090 475 55120 485
rect 55190 1155 55220 1165
rect 55190 485 55195 1155
rect 55215 485 55220 1155
rect 55190 475 55220 485
rect 55290 1155 55320 1165
rect 55290 485 55295 1155
rect 55315 485 55320 1155
rect 55290 475 55320 485
rect 55390 1155 55420 1165
rect 55390 485 55395 1155
rect 55415 485 55420 1155
rect 55390 475 55420 485
rect 55490 1155 55520 1165
rect 55490 485 55495 1155
rect 55515 485 55520 1155
rect 55490 475 55520 485
rect 55590 1155 55660 1165
rect 58145 1155 58215 1165
rect 55590 485 55595 1155
rect 55615 485 55635 1155
rect 55655 485 55660 1155
rect 56185 1145 56255 1155
rect 56185 925 56190 1145
rect 56210 925 56230 1145
rect 56250 925 56255 1145
rect 56185 915 56255 925
rect 56280 1145 56310 1155
rect 56280 925 56285 1145
rect 56305 925 56310 1145
rect 56280 915 56310 925
rect 56335 1145 56365 1155
rect 56335 925 56340 1145
rect 56360 925 56365 1145
rect 56335 915 56365 925
rect 56390 1145 56420 1155
rect 56390 925 56395 1145
rect 56415 925 56420 1145
rect 56390 915 56420 925
rect 56445 1145 56475 1155
rect 56445 925 56450 1145
rect 56470 925 56475 1145
rect 56445 915 56475 925
rect 56500 1145 56530 1155
rect 56500 925 56505 1145
rect 56525 925 56530 1145
rect 56500 915 56530 925
rect 56555 1145 56585 1155
rect 56555 925 56560 1145
rect 56580 925 56585 1145
rect 56555 915 56585 925
rect 56610 1145 56640 1155
rect 56610 925 56615 1145
rect 56635 925 56640 1145
rect 56610 915 56640 925
rect 56665 1145 56695 1155
rect 56665 925 56670 1145
rect 56690 925 56695 1145
rect 56665 915 56695 925
rect 56720 1145 56750 1155
rect 56720 925 56725 1145
rect 56745 925 56750 1145
rect 56720 915 56750 925
rect 56775 1145 56805 1155
rect 56775 925 56780 1145
rect 56800 925 56805 1145
rect 56775 915 56805 925
rect 56830 1145 56860 1155
rect 56830 925 56835 1145
rect 56855 925 56860 1145
rect 56830 915 56860 925
rect 56885 1145 56915 1155
rect 56885 925 56890 1145
rect 56910 925 56915 1145
rect 56885 915 56915 925
rect 56940 1145 56970 1155
rect 56940 925 56945 1145
rect 56965 925 56970 1145
rect 56940 915 56970 925
rect 56995 1145 57025 1155
rect 56995 925 57000 1145
rect 57020 925 57025 1145
rect 56995 915 57025 925
rect 57050 1145 57080 1155
rect 57050 925 57055 1145
rect 57075 925 57080 1145
rect 57050 915 57080 925
rect 57105 1145 57135 1155
rect 57105 925 57110 1145
rect 57130 925 57135 1145
rect 57105 915 57135 925
rect 57160 1145 57190 1155
rect 57160 925 57165 1145
rect 57185 925 57190 1145
rect 57160 915 57190 925
rect 57215 1145 57245 1155
rect 57215 925 57220 1145
rect 57240 925 57245 1145
rect 57215 915 57245 925
rect 57270 1145 57300 1155
rect 57270 925 57275 1145
rect 57295 925 57300 1145
rect 57270 915 57300 925
rect 57325 1145 57355 1155
rect 57325 925 57330 1145
rect 57350 925 57355 1145
rect 57325 915 57355 925
rect 57380 1145 57410 1155
rect 57380 925 57385 1145
rect 57405 925 57410 1145
rect 57380 915 57410 925
rect 57435 1145 57465 1155
rect 57435 925 57440 1145
rect 57460 925 57465 1145
rect 57435 915 57465 925
rect 57490 1145 57560 1155
rect 57490 925 57495 1145
rect 57515 925 57535 1145
rect 57555 925 57560 1145
rect 57490 915 57560 925
rect 56220 885 56260 895
rect 56220 865 56230 885
rect 56250 865 56260 885
rect 56220 855 56260 865
rect 57485 885 57525 895
rect 57485 865 57495 885
rect 57515 865 57525 885
rect 57485 855 57525 865
rect 56595 740 56635 750
rect 56595 720 56605 740
rect 56625 720 56635 740
rect 56595 710 56635 720
rect 57040 740 57080 750
rect 57040 720 57050 740
rect 57070 720 57080 740
rect 57040 710 57080 720
rect 56395 680 56465 690
rect 56395 560 56400 680
rect 56420 560 56440 680
rect 56460 560 56465 680
rect 56395 550 56465 560
rect 56490 680 56520 690
rect 56490 560 56495 680
rect 56515 560 56520 680
rect 56490 550 56520 560
rect 56545 680 56575 690
rect 56545 560 56550 680
rect 56570 560 56575 680
rect 56545 550 56575 560
rect 56600 680 56630 690
rect 56600 560 56605 680
rect 56625 560 56630 680
rect 56600 550 56630 560
rect 56655 680 56685 690
rect 56655 560 56660 680
rect 56680 560 56685 680
rect 56655 550 56685 560
rect 56710 680 56740 690
rect 56710 560 56715 680
rect 56735 560 56740 680
rect 56710 550 56740 560
rect 56765 680 56835 690
rect 56765 560 56770 680
rect 56790 560 56810 680
rect 56830 560 56835 680
rect 56765 550 56835 560
rect 56875 680 56905 690
rect 56875 560 56880 680
rect 56900 560 56905 680
rect 56875 550 56905 560
rect 57215 680 57245 690
rect 57215 560 57220 680
rect 57240 560 57245 680
rect 57215 550 57245 560
rect 56435 520 56465 530
rect 56435 500 56440 520
rect 56460 500 56465 520
rect 56435 490 56465 500
rect 56765 520 56795 530
rect 56765 500 56770 520
rect 56790 500 56795 520
rect 56765 490 56795 500
rect 55590 475 55660 485
rect 58145 485 58150 1155
rect 58170 485 58190 1155
rect 58210 485 58215 1155
rect 58145 475 58215 485
rect 58285 1155 58315 1165
rect 58285 485 58290 1155
rect 58310 485 58315 1155
rect 58285 475 58315 485
rect 58385 1155 58415 1165
rect 58385 485 58390 1155
rect 58410 485 58415 1155
rect 58385 475 58415 485
rect 58485 1155 58515 1165
rect 58485 485 58490 1155
rect 58510 485 58515 1155
rect 58485 475 58515 485
rect 58585 1155 58615 1165
rect 58585 485 58590 1155
rect 58610 485 58615 1155
rect 58585 475 58615 485
rect 58685 1155 58715 1165
rect 58685 485 58690 1155
rect 58710 485 58715 1155
rect 58685 475 58715 485
rect 58785 1155 58855 1165
rect 58785 485 58790 1155
rect 58810 485 58830 1155
rect 58850 485 58855 1155
rect 58975 1145 59010 1155
rect 58975 1120 58980 1145
rect 59005 1120 59010 1145
rect 58975 1110 59010 1120
rect 59035 1145 59070 1155
rect 59035 1120 59040 1145
rect 59065 1120 59070 1145
rect 59035 1110 59070 1120
rect 58785 475 58855 485
rect 54990 445 55020 455
rect 54990 425 54995 445
rect 55015 425 55020 445
rect 54990 415 55020 425
rect 55590 445 55620 455
rect 55590 425 55595 445
rect 55615 425 55620 445
rect 55590 415 55620 425
rect 58185 445 58215 455
rect 58185 425 58190 445
rect 58210 425 58215 445
rect 58185 415 58215 425
rect 58785 445 58815 455
rect 58785 425 58790 445
rect 58810 425 58815 445
rect 58785 415 58815 425
rect 59010 423 59035 473
<< viali >>
rect 56095 4735 56115 4755
rect 56275 4735 56295 4755
rect 57035 4735 57055 4755
rect 57215 4735 57235 4755
rect 57505 4735 57525 4755
rect 57685 4735 57705 4755
rect 56095 4375 56115 4695
rect 56155 4375 56175 4695
rect 56215 4375 56235 4695
rect 56275 4375 56295 4695
rect 56565 4565 56585 4585
rect 56745 4565 56765 4585
rect 56565 4375 56585 4525
rect 56625 4375 56645 4525
rect 56685 4375 56705 4525
rect 56745 4375 56765 4525
rect 57035 4375 57055 4695
rect 57095 4375 57115 4695
rect 57155 4375 57175 4695
rect 57215 4375 57235 4695
rect 57505 4375 57525 4695
rect 57565 4375 57585 4695
rect 57625 4375 57645 4695
rect 57685 4375 57705 4695
rect 56160 4285 56180 4305
rect 56635 4285 56655 4305
rect 57145 4285 57165 4305
rect 57581 4275 57601 4295
rect 54935 4065 54955 4085
rect 55655 4065 55675 4085
rect 56015 4065 56035 4085
rect 56735 4065 56755 4085
rect 57045 4065 57065 4085
rect 57765 4065 57785 4085
rect 58130 4065 58150 4085
rect 58850 4065 58870 4085
rect 54935 3705 54955 4025
rect 54995 3705 55015 4025
rect 55055 3705 55075 4025
rect 55115 3705 55135 4025
rect 55175 3705 55195 4025
rect 55235 3705 55255 4025
rect 55295 3705 55315 4025
rect 55355 3705 55375 4025
rect 55415 3705 55435 4025
rect 55475 3705 55495 4025
rect 55535 3705 55555 4025
rect 55595 3705 55615 4025
rect 55655 3705 55675 4025
rect 56015 3705 56035 4025
rect 56075 3705 56095 4025
rect 56135 3705 56155 4025
rect 56195 3705 56215 4025
rect 56255 3705 56275 4025
rect 56315 3705 56335 4025
rect 56375 3705 56395 4025
rect 56435 3705 56455 4025
rect 56495 3705 56515 4025
rect 56555 3705 56575 4025
rect 56615 3705 56635 4025
rect 56675 3705 56695 4025
rect 56735 3705 56755 4025
rect 57045 3705 57065 4025
rect 57105 3705 57125 4025
rect 57165 3705 57185 4025
rect 57225 3705 57245 4025
rect 57285 3705 57305 4025
rect 57345 3705 57365 4025
rect 57405 3705 57425 4025
rect 57465 3705 57485 4025
rect 57525 3705 57545 4025
rect 57585 3705 57605 4025
rect 57645 3705 57665 4025
rect 57705 3705 57725 4025
rect 57765 3705 57785 4025
rect 58130 3705 58150 4025
rect 58190 3705 58210 4025
rect 58250 3705 58270 4025
rect 58310 3705 58330 4025
rect 58370 3705 58390 4025
rect 58430 3705 58450 4025
rect 58490 3705 58510 4025
rect 58550 3705 58570 4025
rect 58610 3705 58630 4025
rect 58670 3705 58690 4025
rect 58730 3705 58750 4025
rect 58790 3705 58810 4025
rect 58850 3705 58870 4025
rect 56405 3560 56425 3580
rect 57375 3560 57395 3580
rect 55325 3515 55345 3535
rect 58460 3515 58480 3535
rect 54960 3375 54980 3395
rect 55620 3375 55640 3395
rect 58160 3375 58180 3395
rect 58820 3375 58840 3395
rect 54560 3295 54580 3315
rect 54615 3295 54635 3315
rect 54670 3295 54690 3315
rect 54960 2765 54980 3335
rect 55015 2765 55035 3335
rect 55070 2765 55090 3335
rect 55125 2765 55145 3335
rect 55180 2765 55200 3335
rect 55235 2765 55255 3335
rect 55290 2765 55310 3335
rect 55345 2765 55365 3335
rect 55400 2765 55420 3335
rect 55455 2765 55475 3335
rect 55510 2765 55530 3335
rect 55565 2765 55585 3335
rect 55620 2765 55640 3335
rect 56285 3320 56305 3340
rect 56340 3320 56360 3340
rect 56395 3320 56415 3340
rect 56450 3320 56470 3340
rect 56505 3320 56525 3340
rect 56560 3320 56580 3340
rect 56615 3320 56635 3340
rect 56670 3320 56690 3340
rect 56725 3320 56745 3340
rect 56780 3320 56800 3340
rect 56835 3320 56855 3340
rect 56890 3320 56910 3340
rect 56945 3320 56965 3340
rect 57000 3320 57020 3340
rect 57055 3320 57075 3340
rect 57110 3320 57130 3340
rect 57165 3320 57185 3340
rect 57220 3320 57240 3340
rect 57275 3320 57295 3340
rect 57330 3320 57350 3340
rect 57385 3320 57405 3340
rect 57440 3320 57460 3340
rect 57495 3320 57515 3340
rect 56285 3260 56305 3280
rect 57495 3260 57515 3280
rect 56805 3130 56825 3150
rect 55995 3045 56015 3065
rect 56745 3045 56765 3065
rect 57035 3045 57055 3065
rect 57785 3045 57805 3065
rect 56040 2960 56060 2980
rect 56095 2960 56115 2980
rect 56150 2960 56170 2980
rect 56205 2960 56225 2980
rect 56260 2960 56280 2980
rect 56315 2960 56335 2980
rect 56370 2960 56390 2980
rect 56425 2960 56445 2980
rect 56480 2960 56500 2980
rect 56535 2960 56555 2980
rect 56590 2960 56610 2980
rect 56645 2960 56665 2980
rect 56700 2960 56720 2980
rect 57080 2960 57100 2980
rect 57135 2960 57155 2980
rect 57190 2960 57210 2980
rect 57245 2960 57265 2980
rect 57300 2960 57320 2980
rect 57355 2960 57375 2980
rect 57410 2960 57430 2980
rect 57465 2960 57485 2980
rect 57520 2960 57540 2980
rect 57575 2960 57595 2980
rect 57630 2960 57650 2980
rect 57685 2960 57705 2980
rect 57740 2960 57760 2980
rect 56040 2900 56060 2920
rect 56700 2900 56720 2920
rect 57080 2900 57100 2920
rect 57740 2900 57760 2920
rect 56100 2815 56120 2835
rect 56585 2815 56605 2835
rect 57195 2815 57215 2835
rect 58160 2765 58180 3335
rect 58215 2765 58235 3335
rect 58270 2765 58290 3335
rect 58325 2765 58345 3335
rect 58380 2765 58400 3335
rect 58435 2765 58455 3335
rect 58490 2765 58510 3335
rect 58545 2765 58565 3335
rect 58600 2765 58620 3335
rect 58655 2765 58675 3335
rect 58710 2765 58730 3335
rect 58765 2765 58785 3335
rect 58820 2765 58840 3335
rect 59110 3295 59130 3315
rect 59165 3295 59185 3315
rect 59220 3295 59240 3315
rect 54560 2690 54580 2710
rect 54615 2690 54635 2710
rect 54670 2690 54690 2710
rect 59110 2690 59130 2710
rect 59165 2690 59185 2710
rect 59220 2690 59240 2710
rect 55320 2615 55340 2635
rect 56725 2610 56745 2630
rect 56945 2610 56965 2630
rect 58460 2615 58480 2635
rect 56560 2550 56580 2570
rect 56615 2550 56635 2570
rect 56670 2550 56690 2570
rect 56725 2550 56745 2570
rect 56780 2550 56800 2570
rect 56835 2550 56855 2570
rect 56890 2550 56910 2570
rect 56945 2550 56965 2570
rect 57000 2550 57020 2570
rect 57055 2550 57075 2570
rect 57110 2550 57130 2570
rect 57165 2550 57185 2570
rect 57220 2550 57240 2570
rect 56560 2490 56580 2510
rect 57220 2490 57240 2510
rect 54960 2445 54980 2465
rect 55620 2445 55640 2465
rect 58160 2445 58180 2465
rect 58820 2445 58840 2465
rect 54960 2235 54980 2405
rect 55015 2235 55035 2405
rect 55070 2235 55090 2405
rect 55125 2235 55145 2405
rect 55180 2235 55200 2405
rect 55235 2235 55255 2405
rect 55290 2235 55310 2405
rect 55345 2235 55365 2405
rect 55400 2235 55420 2405
rect 55455 2235 55475 2405
rect 55510 2235 55530 2405
rect 55565 2235 55585 2405
rect 55620 2235 55640 2405
rect 56640 2245 56660 2265
rect 57140 2245 57160 2265
rect 57790 2220 57810 2240
rect 58160 2235 58180 2405
rect 58215 2235 58235 2405
rect 58270 2235 58290 2405
rect 58325 2235 58345 2405
rect 58380 2235 58400 2405
rect 58435 2235 58455 2405
rect 58490 2235 58510 2405
rect 58545 2235 58565 2405
rect 58600 2235 58620 2405
rect 58655 2235 58675 2405
rect 58710 2235 58730 2405
rect 58765 2235 58785 2405
rect 58820 2235 58840 2405
rect 55070 2175 55090 2195
rect 55180 2175 55200 2195
rect 55290 2175 55310 2195
rect 55400 2175 55420 2195
rect 55510 2175 55530 2195
rect 58270 2175 58290 2195
rect 55320 2025 55340 2045
rect 56040 2045 56060 2165
rect 56095 2045 56115 2165
rect 56150 2045 56170 2165
rect 56205 2045 56225 2165
rect 56260 2045 56280 2165
rect 56315 2045 56335 2165
rect 56370 2045 56390 2165
rect 56425 2045 56445 2165
rect 56480 2045 56500 2165
rect 56535 2045 56555 2165
rect 56590 2045 56610 2165
rect 56645 2045 56665 2165
rect 56700 2045 56720 2165
rect 57080 2045 57100 2165
rect 57135 2045 57155 2165
rect 57190 2045 57210 2165
rect 57245 2045 57265 2165
rect 57300 2045 57320 2165
rect 57355 2045 57375 2165
rect 57410 2045 57430 2165
rect 57465 2045 57485 2165
rect 57520 2045 57540 2165
rect 57575 2045 57595 2165
rect 57630 2045 57650 2165
rect 57685 2045 57705 2165
rect 58380 2175 58400 2195
rect 58490 2175 58510 2195
rect 58600 2175 58620 2195
rect 58710 2175 58730 2195
rect 57740 2045 57760 2165
rect 56040 1985 56060 2005
rect 56700 1985 56720 2005
rect 57080 1985 57100 2005
rect 58460 2025 58480 2045
rect 57740 1985 57760 2005
rect 54455 1515 54480 1540
rect 54515 1515 54540 1540
rect 54575 1515 54600 1540
rect 54960 1575 54980 1845
rect 55015 1575 55035 1845
rect 55070 1575 55090 1845
rect 55125 1575 55145 1845
rect 55180 1575 55200 1845
rect 55235 1575 55255 1845
rect 55290 1575 55310 1845
rect 55345 1575 55365 1845
rect 55400 1575 55420 1845
rect 55455 1575 55475 1845
rect 55510 1575 55530 1845
rect 55565 1575 55585 1845
rect 55620 1575 55640 1845
rect 55995 1760 56015 1780
rect 56695 1760 56715 1780
rect 56864 1760 56884 1780
rect 56916 1760 56936 1780
rect 57085 1760 57105 1780
rect 57785 1760 57805 1780
rect 56040 1575 56060 1695
rect 56095 1575 56115 1695
rect 56150 1575 56170 1695
rect 56205 1575 56225 1695
rect 56260 1575 56280 1695
rect 56315 1575 56335 1695
rect 56370 1575 56390 1695
rect 56425 1575 56445 1695
rect 56480 1575 56500 1695
rect 56535 1575 56555 1695
rect 56590 1575 56610 1695
rect 56645 1575 56665 1695
rect 56700 1575 56720 1695
rect 56780 1575 56800 1695
rect 56835 1575 56855 1695
rect 56890 1575 56910 1695
rect 56945 1575 56965 1695
rect 57000 1575 57020 1695
rect 57080 1575 57100 1695
rect 57135 1575 57155 1695
rect 57190 1575 57210 1695
rect 57245 1575 57265 1695
rect 57300 1575 57320 1695
rect 57355 1575 57375 1695
rect 57410 1575 57430 1695
rect 57465 1575 57485 1695
rect 57520 1575 57540 1695
rect 57575 1575 57595 1695
rect 57630 1575 57650 1695
rect 57685 1575 57705 1695
rect 57740 1575 57760 1695
rect 58160 1575 58180 1845
rect 58215 1575 58235 1845
rect 58270 1575 58290 1845
rect 58325 1575 58345 1845
rect 58380 1575 58400 1845
rect 58435 1575 58455 1845
rect 58490 1575 58510 1845
rect 58545 1575 58565 1845
rect 58600 1575 58620 1845
rect 58655 1575 58675 1845
rect 58710 1575 58730 1845
rect 58765 1575 58785 1845
rect 58820 1575 58840 1845
rect 54635 1515 54660 1540
rect 54960 1515 54980 1535
rect 55620 1515 55640 1535
rect 56040 1515 56060 1535
rect 56740 1515 56760 1535
rect 57040 1515 57060 1535
rect 57740 1515 57760 1535
rect 58160 1515 58180 1535
rect 58820 1515 58840 1535
rect 59140 1515 59165 1540
rect 59200 1515 59225 1540
rect 59260 1515 59285 1540
rect 59320 1515 59345 1540
rect 57415 1240 57435 1260
rect 55345 1195 55365 1215
rect 56835 1185 56855 1205
rect 58440 1195 58460 1215
rect 54740 1120 54765 1145
rect 54800 1120 54825 1145
rect 54995 485 55015 1155
rect 55095 485 55115 1155
rect 55195 485 55215 1155
rect 55295 485 55315 1155
rect 55395 485 55415 1155
rect 55495 485 55515 1155
rect 55595 485 55615 1155
rect 56230 925 56250 1145
rect 56285 925 56305 1145
rect 56340 925 56360 1145
rect 56395 925 56415 1145
rect 56450 925 56470 1145
rect 56505 925 56525 1145
rect 56560 925 56580 1145
rect 56615 925 56635 1145
rect 56670 925 56690 1145
rect 56725 925 56745 1145
rect 56780 925 56800 1145
rect 56835 925 56855 1145
rect 56890 925 56910 1145
rect 56945 925 56965 1145
rect 57000 925 57020 1145
rect 57055 925 57075 1145
rect 57110 925 57130 1145
rect 57165 925 57185 1145
rect 57220 925 57240 1145
rect 57275 925 57295 1145
rect 57330 925 57350 1145
rect 57385 925 57405 1145
rect 57440 925 57460 1145
rect 57495 925 57515 1145
rect 56230 865 56250 885
rect 57495 865 57515 885
rect 56605 720 56625 740
rect 57050 720 57070 740
rect 56440 560 56460 680
rect 56495 560 56515 680
rect 56550 560 56570 680
rect 56605 560 56625 680
rect 56660 560 56680 680
rect 56715 560 56735 680
rect 56770 560 56790 680
rect 56880 560 56900 680
rect 57220 560 57240 680
rect 56440 500 56460 520
rect 56770 500 56790 520
rect 58190 485 58210 1155
rect 58290 485 58310 1155
rect 58390 485 58410 1155
rect 58490 485 58510 1155
rect 58590 485 58610 1155
rect 58690 485 58710 1155
rect 58790 485 58810 1155
rect 58980 1120 59005 1145
rect 59040 1120 59065 1145
rect 54995 425 55015 445
rect 55595 425 55615 445
rect 58190 425 58210 445
rect 58790 425 58810 445
<< metal1 >>
rect 56880 6185 56920 6190
rect 56880 6155 56885 6185
rect 56915 6155 56920 6185
rect 56880 6150 56920 6155
rect 56205 4815 56245 4820
rect 56205 4785 56210 4815
rect 56240 4785 56245 4815
rect 56085 4760 56125 4765
rect 56085 4730 56090 4760
rect 56120 4730 56125 4760
rect 56085 4725 56125 4730
rect 56205 4760 56245 4785
rect 56675 4815 56715 4820
rect 56675 4785 56680 4815
rect 56710 4785 56715 4815
rect 56675 4780 56715 4785
rect 56205 4730 56210 4760
rect 56240 4730 56245 4760
rect 56205 4725 56245 4730
rect 56265 4760 56305 4765
rect 56265 4730 56270 4760
rect 56300 4730 56305 4760
rect 56265 4725 56305 4730
rect 56090 4695 56120 4725
rect 56090 4375 56095 4695
rect 56115 4375 56120 4695
rect 56090 4365 56120 4375
rect 56150 4695 56180 4705
rect 56150 4375 56155 4695
rect 56175 4375 56180 4695
rect 56150 4315 56180 4375
rect 56210 4695 56240 4725
rect 56210 4375 56215 4695
rect 56235 4375 56240 4695
rect 56210 4360 56240 4375
rect 56270 4695 56300 4725
rect 56270 4375 56275 4695
rect 56295 4375 56300 4695
rect 56555 4590 56595 4595
rect 56555 4560 56560 4590
rect 56590 4560 56595 4590
rect 56555 4555 56595 4560
rect 56615 4590 56655 4595
rect 56615 4560 56620 4590
rect 56650 4560 56655 4590
rect 56615 4555 56655 4560
rect 56270 4365 56300 4375
rect 56560 4525 56590 4555
rect 56560 4375 56565 4525
rect 56585 4375 56590 4525
rect 56560 4365 56590 4375
rect 56620 4525 56650 4555
rect 56620 4375 56625 4525
rect 56645 4375 56650 4525
rect 56620 4365 56650 4375
rect 56680 4525 56710 4780
rect 56890 4765 56910 6150
rect 57085 4815 57125 4820
rect 57085 4785 57090 4815
rect 57120 4785 57125 4815
rect 57085 4780 57125 4785
rect 57555 4815 57595 4820
rect 57555 4785 57560 4815
rect 57590 4785 57595 4815
rect 56880 4760 56920 4765
rect 56880 4730 56885 4760
rect 56915 4730 56920 4760
rect 56880 4725 56920 4730
rect 57025 4760 57065 4765
rect 57025 4730 57030 4760
rect 57060 4730 57065 4760
rect 57025 4725 57065 4730
rect 56890 4595 56910 4725
rect 57030 4695 57060 4725
rect 56735 4590 56775 4595
rect 56735 4560 56740 4590
rect 56770 4560 56775 4590
rect 56735 4555 56775 4560
rect 56880 4590 56920 4595
rect 56880 4560 56885 4590
rect 56915 4560 56920 4590
rect 56880 4555 56920 4560
rect 56680 4375 56685 4525
rect 56705 4375 56710 4525
rect 56680 4360 56710 4375
rect 56740 4525 56770 4555
rect 56740 4375 56745 4525
rect 56765 4375 56770 4525
rect 56740 4365 56770 4375
rect 56205 4355 56245 4360
rect 56205 4325 56210 4355
rect 56240 4325 56245 4355
rect 56205 4320 56245 4325
rect 56675 4355 56715 4360
rect 56675 4325 56680 4355
rect 56710 4325 56715 4355
rect 56675 4320 56715 4325
rect 56150 4310 56190 4315
rect 56150 4280 56155 4310
rect 56185 4280 56190 4310
rect 56150 4275 56190 4280
rect 56630 4310 56660 4315
rect 56630 4275 56660 4280
rect 56825 4310 56865 4315
rect 56825 4280 56830 4310
rect 56860 4280 56865 4310
rect 56825 4275 56865 4280
rect 54925 4200 54965 4205
rect 54925 4170 54930 4200
rect 54960 4170 54965 4200
rect 54925 4165 54965 4170
rect 55045 4200 55085 4205
rect 55045 4170 55050 4200
rect 55080 4170 55085 4200
rect 55045 4165 55085 4170
rect 55165 4200 55205 4205
rect 55165 4170 55170 4200
rect 55200 4170 55205 4200
rect 55165 4165 55205 4170
rect 55285 4200 55325 4205
rect 55285 4170 55290 4200
rect 55320 4170 55325 4200
rect 55285 4165 55325 4170
rect 55405 4200 55445 4205
rect 55405 4170 55410 4200
rect 55440 4170 55445 4200
rect 55405 4165 55445 4170
rect 55525 4200 55565 4205
rect 55525 4170 55530 4200
rect 55560 4170 55565 4200
rect 55525 4165 55565 4170
rect 55645 4200 55685 4205
rect 55645 4170 55650 4200
rect 55680 4170 55685 4200
rect 55645 4165 55685 4170
rect 55755 4200 55795 4205
rect 55755 4170 55760 4200
rect 55790 4170 55795 4200
rect 55755 4165 55795 4170
rect 54930 4085 54960 4165
rect 54930 4065 54935 4085
rect 54955 4065 54960 4085
rect 54930 4025 54960 4065
rect 54985 4075 55025 4080
rect 54985 4045 54990 4075
rect 55020 4045 55025 4075
rect 54985 4040 55025 4045
rect 54930 3705 54935 4025
rect 54955 3705 54960 4025
rect 54930 3645 54960 3705
rect 54990 4025 55020 4040
rect 54990 3705 54995 4025
rect 55015 3705 55020 4025
rect 54990 3690 55020 3705
rect 55050 4025 55080 4165
rect 55105 4075 55145 4080
rect 55105 4045 55110 4075
rect 55140 4045 55145 4075
rect 55105 4040 55145 4045
rect 55050 3705 55055 4025
rect 55075 3705 55080 4025
rect 54985 3685 55025 3690
rect 54985 3655 54990 3685
rect 55020 3655 55025 3685
rect 54985 3650 55025 3655
rect 55050 3645 55080 3705
rect 55110 4025 55140 4040
rect 55110 3705 55115 4025
rect 55135 3705 55140 4025
rect 55110 3690 55140 3705
rect 55170 4025 55200 4165
rect 55225 4075 55265 4080
rect 55225 4045 55230 4075
rect 55260 4045 55265 4075
rect 55225 4040 55265 4045
rect 55170 3705 55175 4025
rect 55195 3705 55200 4025
rect 55105 3685 55145 3690
rect 55105 3655 55110 3685
rect 55140 3655 55145 3685
rect 55105 3650 55145 3655
rect 55170 3645 55200 3705
rect 55230 4025 55260 4040
rect 55230 3705 55235 4025
rect 55255 3705 55260 4025
rect 55230 3690 55260 3705
rect 55290 4025 55320 4165
rect 55345 4075 55385 4080
rect 55345 4045 55350 4075
rect 55380 4045 55385 4075
rect 55345 4040 55385 4045
rect 55290 3705 55295 4025
rect 55315 3705 55320 4025
rect 55225 3685 55265 3690
rect 55225 3655 55230 3685
rect 55260 3655 55265 3685
rect 55225 3650 55265 3655
rect 55290 3645 55320 3705
rect 55350 4025 55380 4040
rect 55350 3705 55355 4025
rect 55375 3705 55380 4025
rect 55350 3690 55380 3705
rect 55410 4025 55440 4165
rect 55465 4075 55505 4080
rect 55465 4045 55470 4075
rect 55500 4045 55505 4075
rect 55465 4040 55505 4045
rect 55410 3705 55415 4025
rect 55435 3705 55440 4025
rect 55345 3685 55385 3690
rect 55345 3655 55350 3685
rect 55380 3655 55385 3685
rect 55345 3650 55385 3655
rect 55410 3645 55440 3705
rect 55470 4025 55500 4040
rect 55470 3705 55475 4025
rect 55495 3705 55500 4025
rect 55470 3690 55500 3705
rect 55530 4025 55560 4165
rect 55650 4085 55680 4165
rect 55585 4075 55625 4080
rect 55585 4045 55590 4075
rect 55620 4045 55625 4075
rect 55585 4040 55625 4045
rect 55650 4065 55655 4085
rect 55675 4065 55680 4085
rect 55530 3705 55535 4025
rect 55555 3705 55560 4025
rect 55465 3685 55505 3690
rect 55465 3655 55470 3685
rect 55500 3655 55505 3685
rect 55465 3650 55505 3655
rect 55530 3645 55560 3705
rect 55590 4025 55620 4040
rect 55590 3705 55595 4025
rect 55615 3705 55620 4025
rect 55590 3690 55620 3705
rect 55650 4025 55680 4065
rect 55650 3705 55655 4025
rect 55675 3705 55680 4025
rect 55585 3685 55625 3690
rect 55585 3655 55590 3685
rect 55620 3655 55625 3685
rect 55585 3650 55625 3655
rect 55650 3645 55680 3705
rect 54925 3640 54965 3645
rect 54925 3610 54930 3640
rect 54960 3610 54965 3640
rect 54925 3605 54965 3610
rect 55045 3640 55085 3645
rect 55045 3610 55050 3640
rect 55080 3610 55085 3640
rect 55045 3605 55085 3610
rect 55165 3640 55205 3645
rect 55165 3610 55170 3640
rect 55200 3610 55205 3640
rect 55165 3605 55205 3610
rect 55285 3640 55325 3645
rect 55285 3610 55290 3640
rect 55320 3610 55325 3640
rect 55285 3605 55325 3610
rect 55405 3640 55445 3645
rect 55405 3610 55410 3640
rect 55440 3610 55445 3640
rect 55405 3605 55445 3610
rect 55525 3640 55565 3645
rect 55525 3610 55530 3640
rect 55560 3610 55565 3640
rect 55525 3605 55565 3610
rect 55645 3640 55685 3645
rect 55645 3610 55650 3640
rect 55680 3610 55685 3640
rect 55645 3605 55685 3610
rect 55710 3640 55750 3645
rect 55710 3610 55715 3640
rect 55745 3610 55750 3640
rect 55710 3605 55750 3610
rect 55315 3540 55355 3545
rect 55315 3510 55320 3540
rect 55350 3510 55355 3540
rect 55315 3505 55355 3510
rect 54950 3480 54990 3485
rect 54950 3450 54955 3480
rect 54985 3450 54990 3480
rect 54950 3445 54990 3450
rect 55060 3480 55100 3485
rect 55060 3450 55065 3480
rect 55095 3450 55100 3480
rect 55060 3445 55100 3450
rect 55170 3480 55210 3485
rect 55170 3450 55175 3480
rect 55205 3450 55210 3480
rect 55170 3445 55210 3450
rect 55280 3480 55320 3485
rect 55280 3450 55285 3480
rect 55315 3450 55320 3480
rect 55280 3445 55320 3450
rect 55390 3480 55430 3485
rect 55390 3450 55395 3480
rect 55425 3450 55430 3480
rect 55390 3445 55430 3450
rect 55500 3480 55540 3485
rect 55500 3450 55505 3480
rect 55535 3450 55540 3480
rect 55500 3445 55540 3450
rect 55610 3480 55650 3485
rect 55610 3450 55615 3480
rect 55645 3450 55650 3480
rect 55610 3445 55650 3450
rect 54605 3400 54645 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 54955 3395 54985 3445
rect 54955 3375 54960 3395
rect 54980 3375 54985 3395
rect 54615 3325 54635 3365
rect 54955 3335 54985 3375
rect 55005 3385 55045 3390
rect 55005 3355 55010 3385
rect 55040 3355 55045 3385
rect 55005 3350 55045 3355
rect 54554 3315 54695 3325
rect 54554 3295 54560 3315
rect 54580 3295 54615 3315
rect 54635 3295 54670 3315
rect 54690 3295 54695 3315
rect 54554 3285 54695 3295
rect 54955 2765 54960 3335
rect 54980 2765 54985 3335
rect 54554 2710 54695 2720
rect 54554 2690 54560 2710
rect 54580 2690 54615 2710
rect 54635 2690 54670 2710
rect 54690 2690 54695 2710
rect 54955 2705 54985 2765
rect 55010 3335 55040 3350
rect 55010 2765 55015 3335
rect 55035 2765 55040 3335
rect 55010 2750 55040 2765
rect 55065 3335 55095 3445
rect 55115 3385 55155 3390
rect 55115 3355 55120 3385
rect 55150 3355 55155 3385
rect 55115 3350 55155 3355
rect 55065 2765 55070 3335
rect 55090 2765 55095 3335
rect 55005 2745 55045 2750
rect 55005 2715 55010 2745
rect 55040 2715 55045 2745
rect 55005 2710 55045 2715
rect 55065 2705 55095 2765
rect 55120 3335 55150 3350
rect 55120 2765 55125 3335
rect 55145 2765 55150 3335
rect 55120 2750 55150 2765
rect 55175 3335 55205 3445
rect 55225 3385 55265 3390
rect 55225 3355 55230 3385
rect 55260 3355 55265 3385
rect 55225 3350 55265 3355
rect 55175 2765 55180 3335
rect 55200 2765 55205 3335
rect 55115 2745 55155 2750
rect 55115 2715 55120 2745
rect 55150 2715 55155 2745
rect 55115 2710 55155 2715
rect 55175 2705 55205 2765
rect 55230 3335 55260 3350
rect 55230 2765 55235 3335
rect 55255 2765 55260 3335
rect 55230 2750 55260 2765
rect 55285 3335 55315 3445
rect 55335 3385 55375 3390
rect 55335 3355 55340 3385
rect 55370 3355 55375 3385
rect 55335 3350 55375 3355
rect 55285 2765 55290 3335
rect 55310 2765 55315 3335
rect 55225 2745 55265 2750
rect 55225 2715 55230 2745
rect 55260 2715 55265 2745
rect 55225 2710 55265 2715
rect 55285 2705 55315 2765
rect 55340 3335 55370 3350
rect 55340 2765 55345 3335
rect 55365 2765 55370 3335
rect 55340 2750 55370 2765
rect 55395 3335 55425 3445
rect 55445 3385 55485 3390
rect 55445 3355 55450 3385
rect 55480 3355 55485 3385
rect 55445 3350 55485 3355
rect 55395 2765 55400 3335
rect 55420 2765 55425 3335
rect 55335 2745 55375 2750
rect 55335 2715 55340 2745
rect 55370 2715 55375 2745
rect 55335 2710 55375 2715
rect 55395 2705 55425 2765
rect 55450 3335 55480 3350
rect 55450 2765 55455 3335
rect 55475 2765 55480 3335
rect 55450 2750 55480 2765
rect 55505 3335 55535 3445
rect 55615 3395 55645 3445
rect 55555 3385 55595 3390
rect 55555 3355 55560 3385
rect 55590 3355 55595 3385
rect 55555 3350 55595 3355
rect 55615 3375 55620 3395
rect 55640 3375 55645 3395
rect 55505 2765 55510 3335
rect 55530 2765 55535 3335
rect 55445 2745 55485 2750
rect 55445 2715 55450 2745
rect 55480 2715 55485 2745
rect 55445 2710 55485 2715
rect 54554 2680 54695 2690
rect 54950 2700 54990 2705
rect 54615 2645 54635 2680
rect 54950 2670 54955 2700
rect 54985 2670 54990 2700
rect 54950 2665 54990 2670
rect 55060 2700 55100 2705
rect 55060 2670 55065 2700
rect 55095 2670 55100 2700
rect 55060 2665 55100 2670
rect 55170 2700 55210 2705
rect 55170 2670 55175 2700
rect 55205 2670 55210 2700
rect 55170 2665 55210 2670
rect 55280 2700 55320 2705
rect 55280 2670 55285 2700
rect 55315 2670 55320 2700
rect 55280 2665 55320 2670
rect 55390 2700 55430 2705
rect 55390 2670 55395 2700
rect 55425 2670 55430 2700
rect 55390 2665 55430 2670
rect 54605 2640 54645 2645
rect 54605 2610 54610 2640
rect 54640 2610 54645 2640
rect 54605 2605 54645 2610
rect 55310 2640 55350 2645
rect 55310 2610 55315 2640
rect 55345 2610 55350 2640
rect 55310 2605 55350 2610
rect 55455 2600 55475 2710
rect 55505 2705 55535 2765
rect 55560 3335 55590 3350
rect 55560 2765 55565 3335
rect 55585 2765 55590 3335
rect 55560 2750 55590 2765
rect 55615 3335 55645 3375
rect 55615 2765 55620 3335
rect 55640 2765 55645 3335
rect 55555 2745 55595 2750
rect 55555 2715 55560 2745
rect 55590 2715 55595 2745
rect 55555 2710 55595 2715
rect 55615 2705 55645 2765
rect 55500 2700 55540 2705
rect 55500 2670 55505 2700
rect 55535 2670 55540 2700
rect 55500 2665 55540 2670
rect 55610 2700 55650 2705
rect 55610 2670 55615 2700
rect 55645 2670 55650 2700
rect 55610 2665 55650 2670
rect 55720 2645 55740 3605
rect 55765 3485 55785 4165
rect 56005 4140 56045 4145
rect 56005 4110 56010 4140
rect 56040 4110 56045 4140
rect 56005 4105 56045 4110
rect 56125 4140 56165 4145
rect 56125 4110 56130 4140
rect 56160 4110 56165 4140
rect 56125 4105 56165 4110
rect 56245 4140 56285 4145
rect 56245 4110 56250 4140
rect 56280 4110 56285 4140
rect 56245 4105 56285 4110
rect 56365 4140 56405 4145
rect 56365 4110 56370 4140
rect 56400 4110 56405 4140
rect 56365 4105 56405 4110
rect 56485 4140 56525 4145
rect 56485 4110 56490 4140
rect 56520 4110 56525 4140
rect 56485 4105 56525 4110
rect 56605 4140 56645 4145
rect 56605 4110 56610 4140
rect 56640 4110 56645 4140
rect 56605 4105 56645 4110
rect 56725 4140 56765 4145
rect 56725 4110 56730 4140
rect 56760 4110 56765 4140
rect 56725 4105 56765 4110
rect 56010 4085 56040 4105
rect 56010 4065 56015 4085
rect 56035 4065 56040 4085
rect 56010 4025 56040 4065
rect 56065 4075 56105 4080
rect 56065 4045 56070 4075
rect 56100 4045 56105 4075
rect 56065 4040 56105 4045
rect 56010 3705 56015 4025
rect 56035 3705 56040 4025
rect 56010 3690 56040 3705
rect 56070 4025 56100 4040
rect 56070 3705 56075 4025
rect 56095 3705 56100 4025
rect 56005 3685 56045 3690
rect 56005 3655 56010 3685
rect 56040 3655 56045 3685
rect 56005 3650 56045 3655
rect 56070 3645 56100 3705
rect 56130 4025 56160 4105
rect 56185 4075 56225 4080
rect 56185 4045 56190 4075
rect 56220 4045 56225 4075
rect 56185 4040 56225 4045
rect 56130 3705 56135 4025
rect 56155 3705 56160 4025
rect 56130 3690 56160 3705
rect 56190 4025 56220 4040
rect 56190 3705 56195 4025
rect 56215 3705 56220 4025
rect 56125 3685 56165 3690
rect 56125 3655 56130 3685
rect 56160 3655 56165 3685
rect 56125 3650 56165 3655
rect 56190 3645 56220 3705
rect 56250 4025 56280 4105
rect 56305 4075 56345 4080
rect 56305 4045 56310 4075
rect 56340 4045 56345 4075
rect 56305 4040 56345 4045
rect 56250 3705 56255 4025
rect 56275 3705 56280 4025
rect 56250 3690 56280 3705
rect 56310 4025 56340 4040
rect 56310 3705 56315 4025
rect 56335 3705 56340 4025
rect 56245 3685 56285 3690
rect 56245 3655 56250 3685
rect 56280 3655 56285 3685
rect 56245 3650 56285 3655
rect 56310 3645 56340 3705
rect 56370 4025 56400 4105
rect 56425 4075 56465 4080
rect 56425 4045 56430 4075
rect 56460 4045 56465 4075
rect 56425 4040 56465 4045
rect 56370 3705 56375 4025
rect 56395 3705 56400 4025
rect 56370 3690 56400 3705
rect 56430 4025 56460 4040
rect 56430 3705 56435 4025
rect 56455 3705 56460 4025
rect 56365 3685 56405 3690
rect 56365 3655 56370 3685
rect 56400 3655 56405 3685
rect 56365 3650 56405 3655
rect 56430 3645 56460 3705
rect 56490 4025 56520 4105
rect 56545 4075 56585 4080
rect 56545 4045 56550 4075
rect 56580 4045 56585 4075
rect 56545 4040 56585 4045
rect 56490 3705 56495 4025
rect 56515 3705 56520 4025
rect 56490 3690 56520 3705
rect 56550 4025 56580 4040
rect 56550 3705 56555 4025
rect 56575 3705 56580 4025
rect 56485 3685 56525 3690
rect 56485 3655 56490 3685
rect 56520 3655 56525 3685
rect 56485 3650 56525 3655
rect 56550 3645 56580 3705
rect 56610 4025 56640 4105
rect 56730 4085 56760 4105
rect 56665 4075 56705 4080
rect 56665 4045 56670 4075
rect 56700 4045 56705 4075
rect 56665 4040 56705 4045
rect 56730 4065 56735 4085
rect 56755 4065 56760 4085
rect 56610 3705 56615 4025
rect 56635 3705 56640 4025
rect 56610 3690 56640 3705
rect 56670 4025 56700 4040
rect 56670 3705 56675 4025
rect 56695 3705 56700 4025
rect 56605 3685 56645 3690
rect 56605 3655 56610 3685
rect 56640 3655 56645 3685
rect 56605 3650 56645 3655
rect 56670 3645 56700 3705
rect 56730 4025 56760 4065
rect 56730 3705 56735 4025
rect 56755 3705 56760 4025
rect 56730 3690 56760 3705
rect 56725 3685 56765 3690
rect 56725 3655 56730 3685
rect 56760 3655 56765 3685
rect 56725 3650 56765 3655
rect 56065 3640 56105 3645
rect 56065 3610 56070 3640
rect 56100 3610 56105 3640
rect 56065 3605 56105 3610
rect 56185 3640 56225 3645
rect 56185 3610 56190 3640
rect 56220 3610 56225 3640
rect 56185 3605 56225 3610
rect 56305 3640 56345 3645
rect 56305 3610 56310 3640
rect 56340 3610 56345 3640
rect 56305 3605 56345 3610
rect 56425 3640 56465 3645
rect 56425 3610 56430 3640
rect 56460 3610 56465 3640
rect 56425 3605 56465 3610
rect 56545 3640 56585 3645
rect 56545 3610 56550 3640
rect 56580 3610 56585 3640
rect 56545 3605 56585 3610
rect 56665 3640 56705 3645
rect 56665 3610 56670 3640
rect 56700 3610 56705 3640
rect 56665 3605 56705 3610
rect 56845 3590 56865 4275
rect 56890 4205 56910 4555
rect 57030 4375 57035 4695
rect 57055 4375 57060 4695
rect 57030 4365 57060 4375
rect 57090 4695 57120 4780
rect 57145 4760 57185 4765
rect 57145 4730 57150 4760
rect 57180 4730 57185 4760
rect 57145 4725 57185 4730
rect 57205 4760 57245 4765
rect 57205 4730 57210 4760
rect 57240 4730 57245 4760
rect 57205 4725 57245 4730
rect 57495 4760 57535 4765
rect 57495 4730 57500 4760
rect 57530 4730 57535 4760
rect 57495 4725 57535 4730
rect 57555 4760 57595 4785
rect 57555 4730 57560 4760
rect 57590 4730 57595 4760
rect 57555 4725 57595 4730
rect 57675 4760 57715 4765
rect 57675 4730 57680 4760
rect 57710 4730 57715 4760
rect 57675 4725 57715 4730
rect 57090 4375 57095 4695
rect 57115 4375 57120 4695
rect 57090 4360 57120 4375
rect 57150 4695 57180 4725
rect 57150 4375 57155 4695
rect 57175 4375 57180 4695
rect 57150 4365 57180 4375
rect 57210 4695 57240 4725
rect 57210 4375 57215 4695
rect 57235 4375 57240 4695
rect 57210 4365 57240 4375
rect 57500 4695 57530 4725
rect 57500 4375 57505 4695
rect 57525 4375 57530 4695
rect 57500 4365 57530 4375
rect 57560 4695 57590 4725
rect 57560 4375 57565 4695
rect 57585 4375 57590 4695
rect 57560 4360 57590 4375
rect 57620 4695 57650 4705
rect 57620 4375 57625 4695
rect 57645 4375 57650 4695
rect 57085 4355 57125 4360
rect 57085 4325 57090 4355
rect 57120 4325 57125 4355
rect 57085 4320 57125 4325
rect 57555 4355 57595 4360
rect 57555 4325 57560 4355
rect 57590 4325 57595 4355
rect 57555 4320 57595 4325
rect 57140 4305 57170 4315
rect 57140 4285 57145 4305
rect 57165 4285 57170 4305
rect 56935 4255 56975 4260
rect 56935 4225 56940 4255
rect 56970 4225 56975 4255
rect 57140 4250 57170 4285
rect 57576 4300 57606 4305
rect 57576 4265 57606 4270
rect 57620 4250 57650 4375
rect 57680 4695 57710 4725
rect 57680 4375 57685 4695
rect 57705 4375 57710 4695
rect 57680 4365 57710 4375
rect 56935 4220 56975 4225
rect 57135 4245 57175 4250
rect 56880 4200 56920 4205
rect 56880 4170 56885 4200
rect 56915 4170 56920 4200
rect 56880 4165 56920 4170
rect 56395 3585 56435 3590
rect 56395 3555 56400 3585
rect 56430 3555 56435 3585
rect 56395 3550 56435 3555
rect 56835 3585 56875 3590
rect 56835 3555 56840 3585
rect 56870 3555 56875 3585
rect 56835 3550 56875 3555
rect 56935 3545 56955 4220
rect 57135 4215 57140 4245
rect 57170 4215 57175 4245
rect 57135 4210 57175 4215
rect 57615 4245 57655 4250
rect 57615 4215 57620 4245
rect 57650 4215 57655 4245
rect 57615 4210 57655 4215
rect 58005 4200 58045 4205
rect 58005 4170 58010 4200
rect 58040 4170 58045 4200
rect 58005 4165 58045 4170
rect 58120 4200 58160 4205
rect 58120 4170 58125 4200
rect 58155 4170 58160 4200
rect 58120 4165 58160 4170
rect 58240 4200 58280 4205
rect 58240 4170 58245 4200
rect 58275 4170 58280 4200
rect 58240 4165 58280 4170
rect 58360 4200 58400 4205
rect 58360 4170 58365 4200
rect 58395 4170 58400 4200
rect 58360 4165 58400 4170
rect 58480 4200 58520 4205
rect 58480 4170 58485 4200
rect 58515 4170 58520 4200
rect 58480 4165 58520 4170
rect 58600 4200 58640 4205
rect 58600 4170 58605 4200
rect 58635 4170 58640 4200
rect 58600 4165 58640 4170
rect 58720 4200 58760 4205
rect 58720 4170 58725 4200
rect 58755 4170 58760 4200
rect 58720 4165 58760 4170
rect 58840 4200 58880 4205
rect 58840 4170 58845 4200
rect 58875 4170 58880 4200
rect 58840 4165 58880 4170
rect 57035 4140 57075 4145
rect 57035 4110 57040 4140
rect 57070 4110 57075 4140
rect 57035 4105 57075 4110
rect 57155 4140 57195 4145
rect 57155 4110 57160 4140
rect 57190 4110 57195 4140
rect 57155 4105 57195 4110
rect 57275 4140 57315 4145
rect 57275 4110 57280 4140
rect 57310 4110 57315 4140
rect 57275 4105 57315 4110
rect 57395 4140 57435 4145
rect 57395 4110 57400 4140
rect 57430 4110 57435 4140
rect 57395 4105 57435 4110
rect 57515 4140 57555 4145
rect 57515 4110 57520 4140
rect 57550 4110 57555 4140
rect 57515 4105 57555 4110
rect 57635 4140 57675 4145
rect 57635 4110 57640 4140
rect 57670 4110 57675 4140
rect 57635 4105 57675 4110
rect 57755 4140 57795 4145
rect 57755 4110 57760 4140
rect 57790 4110 57795 4140
rect 57755 4105 57795 4110
rect 57040 4085 57070 4105
rect 57040 4065 57045 4085
rect 57065 4065 57070 4085
rect 57040 4025 57070 4065
rect 57095 4075 57135 4080
rect 57095 4045 57100 4075
rect 57130 4045 57135 4075
rect 57095 4040 57135 4045
rect 57040 3705 57045 4025
rect 57065 3705 57070 4025
rect 57040 3690 57070 3705
rect 57100 4025 57130 4040
rect 57100 3705 57105 4025
rect 57125 3705 57130 4025
rect 57035 3685 57075 3690
rect 57035 3655 57040 3685
rect 57070 3655 57075 3685
rect 57035 3650 57075 3655
rect 57100 3645 57130 3705
rect 57160 4025 57190 4105
rect 57215 4075 57255 4080
rect 57215 4045 57220 4075
rect 57250 4045 57255 4075
rect 57215 4040 57255 4045
rect 57160 3705 57165 4025
rect 57185 3705 57190 4025
rect 57160 3690 57190 3705
rect 57220 4025 57250 4040
rect 57220 3705 57225 4025
rect 57245 3705 57250 4025
rect 57155 3685 57195 3690
rect 57155 3655 57160 3685
rect 57190 3655 57195 3685
rect 57155 3650 57195 3655
rect 57220 3645 57250 3705
rect 57280 4025 57310 4105
rect 57335 4075 57375 4080
rect 57335 4045 57340 4075
rect 57370 4045 57375 4075
rect 57335 4040 57375 4045
rect 57280 3705 57285 4025
rect 57305 3705 57310 4025
rect 57280 3690 57310 3705
rect 57340 4025 57370 4040
rect 57340 3705 57345 4025
rect 57365 3705 57370 4025
rect 57275 3685 57315 3690
rect 57275 3655 57280 3685
rect 57310 3655 57315 3685
rect 57275 3650 57315 3655
rect 57340 3645 57370 3705
rect 57400 4025 57430 4105
rect 57455 4075 57495 4080
rect 57455 4045 57460 4075
rect 57490 4045 57495 4075
rect 57455 4040 57495 4045
rect 57400 3705 57405 4025
rect 57425 3705 57430 4025
rect 57400 3690 57430 3705
rect 57460 4025 57490 4040
rect 57460 3705 57465 4025
rect 57485 3705 57490 4025
rect 57395 3685 57435 3690
rect 57395 3655 57400 3685
rect 57430 3655 57435 3685
rect 57395 3650 57435 3655
rect 57460 3645 57490 3705
rect 57520 4025 57550 4105
rect 57575 4075 57615 4080
rect 57575 4045 57580 4075
rect 57610 4045 57615 4075
rect 57575 4040 57615 4045
rect 57520 3705 57525 4025
rect 57545 3705 57550 4025
rect 57520 3690 57550 3705
rect 57580 4025 57610 4040
rect 57580 3705 57585 4025
rect 57605 3705 57610 4025
rect 57515 3685 57555 3690
rect 57515 3655 57520 3685
rect 57550 3655 57555 3685
rect 57515 3650 57555 3655
rect 57580 3645 57610 3705
rect 57640 4025 57670 4105
rect 57760 4085 57790 4105
rect 57695 4075 57735 4080
rect 57695 4045 57700 4075
rect 57730 4045 57735 4075
rect 57695 4040 57735 4045
rect 57760 4065 57765 4085
rect 57785 4065 57790 4085
rect 57640 3705 57645 4025
rect 57665 3705 57670 4025
rect 57640 3690 57670 3705
rect 57700 4025 57730 4040
rect 57700 3705 57705 4025
rect 57725 3705 57730 4025
rect 57635 3685 57675 3690
rect 57635 3655 57640 3685
rect 57670 3655 57675 3685
rect 57635 3650 57675 3655
rect 57700 3645 57730 3705
rect 57760 4025 57790 4065
rect 57760 3705 57765 4025
rect 57785 3705 57790 4025
rect 57760 3690 57790 3705
rect 57755 3685 57795 3690
rect 57755 3655 57760 3685
rect 57790 3655 57795 3685
rect 57755 3650 57795 3655
rect 57095 3640 57135 3645
rect 57095 3610 57100 3640
rect 57130 3610 57135 3640
rect 57095 3605 57135 3610
rect 57215 3640 57255 3645
rect 57215 3610 57220 3640
rect 57250 3610 57255 3640
rect 57215 3605 57255 3610
rect 57335 3640 57375 3645
rect 57335 3610 57340 3640
rect 57370 3610 57375 3640
rect 57335 3605 57375 3610
rect 57455 3640 57495 3645
rect 57455 3610 57460 3640
rect 57490 3610 57495 3640
rect 57455 3605 57495 3610
rect 57575 3640 57615 3645
rect 57575 3610 57580 3640
rect 57610 3610 57615 3640
rect 57575 3605 57615 3610
rect 57695 3640 57735 3645
rect 57695 3610 57700 3640
rect 57730 3610 57735 3640
rect 57695 3605 57735 3610
rect 57365 3585 57405 3590
rect 57365 3555 57370 3585
rect 57400 3555 57405 3585
rect 57365 3550 57405 3555
rect 56925 3540 56965 3545
rect 56925 3510 56930 3540
rect 56960 3510 56965 3540
rect 56925 3505 56965 3510
rect 58015 3485 58035 4165
rect 58125 4085 58155 4165
rect 58125 4065 58130 4085
rect 58150 4065 58155 4085
rect 58125 4025 58155 4065
rect 58180 4075 58220 4080
rect 58180 4045 58185 4075
rect 58215 4045 58220 4075
rect 58180 4040 58220 4045
rect 58125 3705 58130 4025
rect 58150 3705 58155 4025
rect 58125 3645 58155 3705
rect 58185 4025 58215 4040
rect 58185 3705 58190 4025
rect 58210 3705 58215 4025
rect 58185 3690 58215 3705
rect 58245 4025 58275 4165
rect 58300 4075 58340 4080
rect 58300 4045 58305 4075
rect 58335 4045 58340 4075
rect 58300 4040 58340 4045
rect 58245 3705 58250 4025
rect 58270 3705 58275 4025
rect 58180 3685 58220 3690
rect 58180 3655 58185 3685
rect 58215 3655 58220 3685
rect 58180 3650 58220 3655
rect 58245 3645 58275 3705
rect 58305 4025 58335 4040
rect 58305 3705 58310 4025
rect 58330 3705 58335 4025
rect 58305 3690 58335 3705
rect 58365 4025 58395 4165
rect 58420 4075 58460 4080
rect 58420 4045 58425 4075
rect 58455 4045 58460 4075
rect 58420 4040 58460 4045
rect 58365 3705 58370 4025
rect 58390 3705 58395 4025
rect 58300 3685 58340 3690
rect 58300 3655 58305 3685
rect 58335 3655 58340 3685
rect 58300 3650 58340 3655
rect 58365 3645 58395 3705
rect 58425 4025 58455 4040
rect 58425 3705 58430 4025
rect 58450 3705 58455 4025
rect 58425 3690 58455 3705
rect 58485 4025 58515 4165
rect 58540 4075 58580 4080
rect 58540 4045 58545 4075
rect 58575 4045 58580 4075
rect 58540 4040 58580 4045
rect 58485 3705 58490 4025
rect 58510 3705 58515 4025
rect 58420 3685 58460 3690
rect 58420 3655 58425 3685
rect 58455 3655 58460 3685
rect 58420 3650 58460 3655
rect 58485 3645 58515 3705
rect 58545 4025 58575 4040
rect 58545 3705 58550 4025
rect 58570 3705 58575 4025
rect 58545 3690 58575 3705
rect 58605 4025 58635 4165
rect 58660 4075 58700 4080
rect 58660 4045 58665 4075
rect 58695 4045 58700 4075
rect 58660 4040 58700 4045
rect 58605 3705 58610 4025
rect 58630 3705 58635 4025
rect 58540 3685 58580 3690
rect 58540 3655 58545 3685
rect 58575 3655 58580 3685
rect 58540 3650 58580 3655
rect 58605 3645 58635 3705
rect 58665 4025 58695 4040
rect 58665 3705 58670 4025
rect 58690 3705 58695 4025
rect 58665 3690 58695 3705
rect 58725 4025 58755 4165
rect 58845 4085 58875 4165
rect 58780 4075 58820 4080
rect 58780 4045 58785 4075
rect 58815 4045 58820 4075
rect 58780 4040 58820 4045
rect 58845 4065 58850 4085
rect 58870 4065 58875 4085
rect 58725 3705 58730 4025
rect 58750 3705 58755 4025
rect 58660 3685 58700 3690
rect 58660 3655 58665 3685
rect 58695 3655 58700 3685
rect 58660 3650 58700 3655
rect 58725 3645 58755 3705
rect 58785 4025 58815 4040
rect 58785 3705 58790 4025
rect 58810 3705 58815 4025
rect 58785 3690 58815 3705
rect 58845 4025 58875 4065
rect 58845 3705 58850 4025
rect 58870 3705 58875 4025
rect 58780 3685 58820 3690
rect 58780 3655 58785 3685
rect 58815 3655 58820 3685
rect 58780 3650 58820 3655
rect 58845 3645 58875 3705
rect 58050 3640 58090 3645
rect 58050 3610 58055 3640
rect 58085 3610 58090 3640
rect 58050 3605 58090 3610
rect 58120 3640 58160 3645
rect 58120 3610 58125 3640
rect 58155 3610 58160 3640
rect 58120 3605 58160 3610
rect 58240 3640 58280 3645
rect 58240 3610 58245 3640
rect 58275 3610 58280 3640
rect 58240 3605 58280 3610
rect 58360 3640 58400 3645
rect 58360 3610 58365 3640
rect 58395 3610 58400 3640
rect 58360 3605 58400 3610
rect 58480 3640 58520 3645
rect 58480 3610 58485 3640
rect 58515 3610 58520 3640
rect 58480 3605 58520 3610
rect 58600 3640 58640 3645
rect 58600 3610 58605 3640
rect 58635 3610 58640 3640
rect 58600 3605 58640 3610
rect 58720 3640 58760 3645
rect 58720 3610 58725 3640
rect 58755 3610 58760 3640
rect 58720 3605 58760 3610
rect 58840 3640 58880 3645
rect 58840 3610 58845 3640
rect 58875 3610 58880 3640
rect 58840 3605 58880 3610
rect 55755 3480 55795 3485
rect 55755 3450 55760 3480
rect 55790 3450 55795 3480
rect 55755 3445 55795 3450
rect 56275 3480 56315 3485
rect 56275 3450 56280 3480
rect 56310 3450 56315 3480
rect 56275 3445 56315 3450
rect 56385 3480 56425 3485
rect 56385 3450 56390 3480
rect 56420 3450 56425 3480
rect 56385 3445 56425 3450
rect 56495 3480 56535 3485
rect 56495 3450 56500 3480
rect 56530 3450 56535 3480
rect 56495 3445 56535 3450
rect 56605 3480 56645 3485
rect 56605 3450 56610 3480
rect 56640 3450 56645 3480
rect 56605 3445 56645 3450
rect 56715 3480 56755 3485
rect 56715 3450 56720 3480
rect 56750 3450 56755 3480
rect 56715 3445 56755 3450
rect 56825 3480 56865 3485
rect 56825 3450 56830 3480
rect 56860 3450 56865 3480
rect 56825 3445 56865 3450
rect 56935 3480 56975 3485
rect 56935 3450 56940 3480
rect 56970 3450 56975 3480
rect 56935 3445 56975 3450
rect 57045 3480 57085 3485
rect 57045 3450 57050 3480
rect 57080 3450 57085 3480
rect 57045 3445 57085 3450
rect 57155 3480 57195 3485
rect 57155 3450 57160 3480
rect 57190 3450 57195 3480
rect 57155 3445 57195 3450
rect 57265 3480 57305 3485
rect 57265 3450 57270 3480
rect 57300 3450 57305 3480
rect 57265 3445 57305 3450
rect 57375 3480 57415 3485
rect 57375 3450 57380 3480
rect 57410 3450 57415 3480
rect 57375 3445 57415 3450
rect 57485 3480 57525 3485
rect 57485 3450 57490 3480
rect 57520 3450 57525 3480
rect 57485 3445 57525 3450
rect 58005 3480 58045 3485
rect 58005 3450 58010 3480
rect 58040 3450 58045 3480
rect 58005 3445 58045 3450
rect 55765 2800 55785 3445
rect 56280 3340 56310 3445
rect 56330 3435 56370 3440
rect 56330 3405 56335 3435
rect 56365 3405 56370 3435
rect 56330 3400 56370 3405
rect 56280 3320 56285 3340
rect 56305 3320 56310 3340
rect 56280 3280 56310 3320
rect 56335 3340 56365 3400
rect 56335 3320 56340 3340
rect 56360 3320 56365 3340
rect 56335 3305 56365 3320
rect 56390 3340 56420 3445
rect 56440 3390 56480 3395
rect 56440 3360 56445 3390
rect 56475 3360 56480 3390
rect 56440 3355 56480 3360
rect 56390 3320 56395 3340
rect 56415 3320 56420 3340
rect 56280 3260 56285 3280
rect 56305 3260 56310 3280
rect 56330 3300 56370 3305
rect 56330 3270 56335 3300
rect 56365 3270 56370 3300
rect 56330 3265 56370 3270
rect 56140 3255 56180 3260
rect 56140 3225 56145 3255
rect 56175 3225 56180 3255
rect 56140 3220 56180 3225
rect 56030 3120 56070 3125
rect 56030 3090 56035 3120
rect 56065 3090 56070 3120
rect 56030 3085 56070 3090
rect 55935 3070 55975 3075
rect 55935 3040 55940 3070
rect 55970 3040 55975 3070
rect 55935 3035 55975 3040
rect 55990 3070 56020 3075
rect 55990 3035 56020 3040
rect 55755 2795 55795 2800
rect 55755 2765 55760 2795
rect 55790 2765 55795 2795
rect 55755 2760 55795 2765
rect 55710 2640 55750 2645
rect 55710 2610 55715 2640
rect 55745 2610 55750 2640
rect 55710 2605 55750 2610
rect 54295 2595 54335 2600
rect 54295 2565 54300 2595
rect 54330 2565 54335 2595
rect 54295 2560 54335 2565
rect 55445 2595 55485 2600
rect 55445 2565 55450 2595
rect 55480 2565 55485 2595
rect 55445 2560 55485 2565
rect 54245 2500 54285 2505
rect 54245 2470 54250 2500
rect 54280 2470 54285 2500
rect 54245 2465 54285 2470
rect 54255 400 54275 2465
rect 54305 1920 54325 2560
rect 54950 2545 54990 2550
rect 54950 2515 54955 2545
rect 54985 2515 54990 2545
rect 54950 2510 54990 2515
rect 55610 2545 55650 2550
rect 55610 2515 55615 2545
rect 55645 2515 55650 2545
rect 55610 2510 55650 2515
rect 54955 2465 54985 2510
rect 55005 2500 55045 2505
rect 55005 2470 55010 2500
rect 55040 2470 55045 2500
rect 55005 2465 55045 2470
rect 55115 2500 55155 2505
rect 55115 2470 55120 2500
rect 55150 2470 55155 2500
rect 55115 2465 55155 2470
rect 55225 2500 55265 2505
rect 55225 2470 55230 2500
rect 55260 2470 55265 2500
rect 55225 2465 55265 2470
rect 55335 2500 55375 2505
rect 55335 2470 55340 2500
rect 55370 2470 55375 2500
rect 55335 2465 55375 2470
rect 55445 2500 55485 2505
rect 55445 2470 55450 2500
rect 55480 2470 55485 2500
rect 55445 2465 55485 2470
rect 55555 2500 55595 2505
rect 55555 2470 55560 2500
rect 55590 2470 55595 2500
rect 55555 2465 55595 2470
rect 55615 2465 55645 2510
rect 54955 2445 54960 2465
rect 54980 2445 54985 2465
rect 54955 2405 54985 2445
rect 54955 2235 54960 2405
rect 54980 2235 54985 2405
rect 54760 2200 54800 2205
rect 54760 2170 54765 2200
rect 54795 2170 54800 2200
rect 54760 2165 54800 2170
rect 54290 1910 54340 1920
rect 54290 1880 54300 1910
rect 54330 1880 54340 1910
rect 54290 1870 54340 1880
rect 54305 1210 54325 1870
rect 54450 1545 54485 1550
rect 54450 1505 54485 1510
rect 54510 1545 54545 1550
rect 54510 1505 54545 1510
rect 54570 1545 54605 1550
rect 54570 1505 54605 1510
rect 54630 1545 54665 1550
rect 54630 1505 54665 1510
rect 54460 1425 54480 1505
rect 54580 1490 54600 1505
rect 54770 1490 54790 2165
rect 54955 2115 54985 2235
rect 55010 2405 55040 2465
rect 55060 2455 55100 2460
rect 55060 2425 55065 2455
rect 55095 2425 55100 2455
rect 55060 2420 55100 2425
rect 55010 2235 55015 2405
rect 55035 2235 55040 2405
rect 55010 2160 55040 2235
rect 55065 2405 55095 2420
rect 55065 2235 55070 2405
rect 55090 2235 55095 2405
rect 55065 2205 55095 2235
rect 55120 2405 55150 2465
rect 55170 2455 55210 2460
rect 55170 2425 55175 2455
rect 55205 2425 55210 2455
rect 55170 2420 55210 2425
rect 55120 2235 55125 2405
rect 55145 2235 55150 2405
rect 55060 2200 55100 2205
rect 55060 2170 55065 2200
rect 55095 2170 55100 2200
rect 55060 2165 55100 2170
rect 55120 2160 55150 2235
rect 55175 2405 55205 2420
rect 55175 2235 55180 2405
rect 55200 2235 55205 2405
rect 55175 2205 55205 2235
rect 55230 2405 55260 2465
rect 55280 2455 55320 2460
rect 55280 2425 55285 2455
rect 55315 2425 55320 2455
rect 55280 2420 55320 2425
rect 55230 2235 55235 2405
rect 55255 2235 55260 2405
rect 55170 2200 55210 2205
rect 55170 2170 55175 2200
rect 55205 2170 55210 2200
rect 55170 2165 55210 2170
rect 55230 2160 55260 2235
rect 55285 2405 55315 2420
rect 55285 2235 55290 2405
rect 55310 2235 55315 2405
rect 55285 2205 55315 2235
rect 55340 2405 55370 2465
rect 55390 2455 55430 2460
rect 55390 2425 55395 2455
rect 55425 2425 55430 2455
rect 55390 2420 55430 2425
rect 55340 2235 55345 2405
rect 55365 2235 55370 2405
rect 55280 2200 55320 2205
rect 55280 2170 55285 2200
rect 55315 2170 55320 2200
rect 55280 2165 55320 2170
rect 55340 2160 55370 2235
rect 55395 2405 55425 2420
rect 55395 2235 55400 2405
rect 55420 2235 55425 2405
rect 55395 2205 55425 2235
rect 55450 2405 55480 2465
rect 55500 2455 55540 2460
rect 55500 2425 55505 2455
rect 55535 2425 55540 2455
rect 55500 2420 55540 2425
rect 55450 2235 55455 2405
rect 55475 2235 55480 2405
rect 55390 2200 55430 2205
rect 55390 2170 55395 2200
rect 55425 2170 55430 2200
rect 55390 2165 55430 2170
rect 55450 2160 55480 2235
rect 55505 2405 55535 2420
rect 55505 2235 55510 2405
rect 55530 2235 55535 2405
rect 55505 2205 55535 2235
rect 55560 2405 55590 2465
rect 55560 2235 55565 2405
rect 55585 2235 55590 2405
rect 55500 2200 55540 2205
rect 55500 2170 55505 2200
rect 55535 2170 55540 2200
rect 55500 2165 55540 2170
rect 55560 2160 55590 2235
rect 55615 2445 55620 2465
rect 55640 2445 55645 2465
rect 55615 2405 55645 2445
rect 55615 2235 55620 2405
rect 55640 2235 55645 2405
rect 55005 2155 55045 2160
rect 55005 2125 55010 2155
rect 55040 2125 55045 2155
rect 55005 2120 55045 2125
rect 55115 2155 55155 2160
rect 55115 2125 55120 2155
rect 55150 2125 55155 2155
rect 55115 2120 55155 2125
rect 55225 2155 55265 2160
rect 55225 2125 55230 2155
rect 55260 2125 55265 2155
rect 55225 2120 55265 2125
rect 55335 2155 55375 2160
rect 55335 2125 55340 2155
rect 55370 2125 55375 2155
rect 55335 2120 55375 2125
rect 55445 2155 55485 2160
rect 55445 2125 55450 2155
rect 55480 2125 55485 2155
rect 55445 2120 55485 2125
rect 55555 2155 55595 2160
rect 55555 2125 55560 2155
rect 55590 2125 55595 2155
rect 55555 2120 55595 2125
rect 55615 2115 55645 2235
rect 54950 2110 54990 2115
rect 54950 2080 54955 2110
rect 54985 2080 54990 2110
rect 54950 2075 54990 2080
rect 55610 2110 55650 2115
rect 55610 2080 55615 2110
rect 55645 2080 55650 2110
rect 55610 2075 55650 2080
rect 55720 2055 55740 2605
rect 55765 2550 55785 2760
rect 55755 2545 55795 2550
rect 55755 2515 55760 2545
rect 55790 2515 55795 2545
rect 55755 2510 55795 2515
rect 55310 2050 55350 2055
rect 55310 2020 55315 2050
rect 55345 2020 55350 2050
rect 55310 2015 55350 2020
rect 55710 2050 55750 2055
rect 55710 2020 55715 2050
rect 55745 2020 55750 2050
rect 55710 2015 55750 2020
rect 54950 1985 54990 1990
rect 54950 1955 54955 1985
rect 54985 1955 54990 1985
rect 54950 1950 54990 1955
rect 55610 1985 55650 1990
rect 55610 1955 55615 1985
rect 55645 1955 55650 1985
rect 55610 1950 55650 1955
rect 54805 1895 54845 1900
rect 54805 1865 54810 1895
rect 54840 1865 54845 1895
rect 54805 1860 54845 1865
rect 54815 1545 54835 1860
rect 54955 1845 54985 1950
rect 55005 1940 55045 1945
rect 55005 1910 55010 1940
rect 55040 1910 55045 1940
rect 55005 1905 55045 1910
rect 55115 1940 55155 1945
rect 55115 1910 55120 1940
rect 55150 1910 55155 1940
rect 55115 1905 55155 1910
rect 55225 1940 55265 1945
rect 55225 1910 55230 1940
rect 55260 1910 55265 1940
rect 55225 1905 55265 1910
rect 55335 1940 55375 1945
rect 55335 1910 55340 1940
rect 55370 1910 55375 1940
rect 55335 1905 55375 1910
rect 55445 1940 55485 1945
rect 55445 1910 55450 1940
rect 55480 1910 55485 1940
rect 55445 1905 55485 1910
rect 55555 1940 55595 1945
rect 55555 1910 55560 1940
rect 55590 1910 55595 1940
rect 55555 1905 55595 1910
rect 54955 1575 54960 1845
rect 54980 1575 54985 1845
rect 54805 1540 54845 1545
rect 54805 1510 54810 1540
rect 54840 1510 54845 1540
rect 54805 1505 54845 1510
rect 54955 1535 54985 1575
rect 54955 1515 54960 1535
rect 54980 1515 54985 1535
rect 55010 1845 55040 1905
rect 55060 1895 55100 1900
rect 55060 1865 55065 1895
rect 55095 1865 55100 1895
rect 55060 1860 55100 1865
rect 55010 1575 55015 1845
rect 55035 1575 55040 1845
rect 55010 1515 55040 1575
rect 55065 1845 55095 1860
rect 55065 1575 55070 1845
rect 55090 1575 55095 1845
rect 55065 1560 55095 1575
rect 55120 1845 55150 1905
rect 55170 1895 55210 1900
rect 55170 1865 55175 1895
rect 55205 1865 55210 1895
rect 55170 1860 55210 1865
rect 55120 1575 55125 1845
rect 55145 1575 55150 1845
rect 55060 1555 55100 1560
rect 55060 1525 55065 1555
rect 55095 1525 55100 1555
rect 55060 1520 55100 1525
rect 55120 1515 55150 1575
rect 55175 1845 55205 1860
rect 55175 1575 55180 1845
rect 55200 1575 55205 1845
rect 55175 1560 55205 1575
rect 55230 1845 55260 1905
rect 55280 1895 55320 1900
rect 55280 1865 55285 1895
rect 55315 1865 55320 1895
rect 55280 1860 55320 1865
rect 55230 1575 55235 1845
rect 55255 1575 55260 1845
rect 55170 1555 55210 1560
rect 55170 1525 55175 1555
rect 55205 1525 55210 1555
rect 55170 1520 55210 1525
rect 55230 1515 55260 1575
rect 55285 1845 55315 1860
rect 55285 1575 55290 1845
rect 55310 1575 55315 1845
rect 55285 1560 55315 1575
rect 55340 1845 55370 1905
rect 55390 1895 55430 1900
rect 55390 1865 55395 1895
rect 55425 1865 55430 1895
rect 55390 1860 55430 1865
rect 55340 1575 55345 1845
rect 55365 1575 55370 1845
rect 55280 1555 55320 1560
rect 55280 1525 55285 1555
rect 55315 1525 55320 1555
rect 55280 1520 55320 1525
rect 55340 1515 55370 1575
rect 55395 1845 55425 1860
rect 55395 1575 55400 1845
rect 55420 1575 55425 1845
rect 55395 1560 55425 1575
rect 55450 1845 55480 1905
rect 55500 1895 55540 1900
rect 55500 1865 55505 1895
rect 55535 1865 55540 1895
rect 55500 1860 55540 1865
rect 55450 1575 55455 1845
rect 55475 1575 55480 1845
rect 55390 1555 55430 1560
rect 55390 1525 55395 1555
rect 55425 1525 55430 1555
rect 55390 1520 55430 1525
rect 55450 1515 55480 1575
rect 55505 1845 55535 1860
rect 55505 1575 55510 1845
rect 55530 1575 55535 1845
rect 55505 1560 55535 1575
rect 55560 1845 55590 1905
rect 55560 1575 55565 1845
rect 55585 1575 55590 1845
rect 55500 1555 55540 1560
rect 55500 1525 55505 1555
rect 55535 1525 55540 1555
rect 55500 1520 55540 1525
rect 55560 1515 55590 1575
rect 55615 1845 55645 1950
rect 55615 1575 55620 1845
rect 55640 1575 55645 1845
rect 55615 1535 55645 1575
rect 55615 1515 55620 1535
rect 55640 1515 55645 1535
rect 55765 1515 55785 2510
rect 55845 1935 55885 1940
rect 55845 1905 55850 1935
rect 55880 1905 55885 1935
rect 55845 1900 55885 1905
rect 54570 1485 54610 1490
rect 54570 1455 54575 1485
rect 54605 1455 54610 1485
rect 54570 1450 54610 1455
rect 54760 1485 54800 1490
rect 54760 1455 54765 1485
rect 54795 1455 54800 1485
rect 54955 1470 54985 1515
rect 55005 1510 55045 1515
rect 55005 1480 55010 1510
rect 55040 1480 55045 1510
rect 55005 1475 55045 1480
rect 55115 1510 55155 1515
rect 55115 1480 55120 1510
rect 55150 1480 55155 1510
rect 55115 1475 55155 1480
rect 55225 1510 55265 1515
rect 55225 1480 55230 1510
rect 55260 1480 55265 1510
rect 55225 1475 55265 1480
rect 55335 1510 55375 1515
rect 55335 1480 55340 1510
rect 55370 1480 55375 1510
rect 55335 1475 55375 1480
rect 55445 1510 55485 1515
rect 55445 1480 55450 1510
rect 55480 1480 55485 1510
rect 55445 1475 55485 1480
rect 55555 1510 55595 1515
rect 55555 1480 55560 1510
rect 55590 1480 55595 1510
rect 55555 1475 55595 1480
rect 55615 1470 55645 1515
rect 55755 1510 55795 1515
rect 55755 1480 55760 1510
rect 55790 1480 55795 1510
rect 55755 1475 55795 1480
rect 55855 1470 55875 1900
rect 54760 1450 54800 1455
rect 54950 1465 54990 1470
rect 54950 1435 54955 1465
rect 54985 1435 54990 1465
rect 54950 1430 54990 1435
rect 55610 1465 55650 1470
rect 55610 1435 55615 1465
rect 55645 1435 55650 1465
rect 55610 1430 55650 1435
rect 55845 1465 55885 1470
rect 55845 1435 55850 1465
rect 55880 1435 55885 1465
rect 55845 1430 55885 1435
rect 54450 1420 54490 1425
rect 54450 1390 54455 1420
rect 54485 1390 54490 1420
rect 54450 1385 54490 1390
rect 54730 1325 54770 1330
rect 54730 1295 54735 1325
rect 54765 1295 54770 1325
rect 54730 1290 54770 1295
rect 55335 1325 55375 1330
rect 55335 1295 55340 1325
rect 55370 1295 55375 1325
rect 55335 1290 55375 1295
rect 54295 1205 54335 1210
rect 54295 1175 54300 1205
rect 54330 1175 54335 1205
rect 54295 1170 54335 1175
rect 54740 1155 54760 1290
rect 54985 1250 55025 1255
rect 54985 1220 54990 1250
rect 55020 1220 55025 1250
rect 54985 1215 55025 1220
rect 55185 1250 55225 1255
rect 55185 1220 55190 1250
rect 55220 1220 55225 1250
rect 55345 1225 55365 1290
rect 55385 1250 55425 1255
rect 55185 1215 55225 1220
rect 55340 1215 55370 1225
rect 55385 1220 55390 1250
rect 55420 1220 55425 1250
rect 55385 1215 55425 1220
rect 55585 1250 55625 1255
rect 55585 1220 55590 1250
rect 55620 1220 55625 1250
rect 55585 1215 55625 1220
rect 54795 1205 54835 1210
rect 54795 1175 54800 1205
rect 54830 1175 54835 1205
rect 54795 1170 54835 1175
rect 54805 1155 54825 1170
rect 54990 1155 55020 1215
rect 55085 1205 55125 1210
rect 55085 1175 55090 1205
rect 55120 1175 55125 1205
rect 55085 1170 55125 1175
rect 54735 1150 54770 1155
rect 54735 1110 54770 1115
rect 54795 1150 54830 1155
rect 54795 1110 54830 1115
rect 54990 485 54995 1155
rect 55015 485 55020 1155
rect 54990 445 55020 485
rect 55090 1155 55120 1170
rect 55090 485 55095 1155
rect 55115 485 55120 1155
rect 55090 470 55120 485
rect 55190 1155 55220 1215
rect 55285 1205 55325 1210
rect 55285 1175 55290 1205
rect 55320 1175 55325 1205
rect 55340 1195 55345 1215
rect 55365 1195 55370 1215
rect 55340 1185 55370 1195
rect 55285 1170 55325 1175
rect 55190 485 55195 1155
rect 55215 485 55220 1155
rect 54990 425 54995 445
rect 55015 425 55020 445
rect 55085 465 55125 470
rect 55085 435 55090 465
rect 55120 435 55125 465
rect 55085 430 55125 435
rect 54990 400 55020 425
rect 55190 400 55220 485
rect 55290 1155 55320 1170
rect 55290 485 55295 1155
rect 55315 485 55320 1155
rect 55290 470 55320 485
rect 55390 1155 55420 1215
rect 55485 1205 55525 1210
rect 55485 1175 55490 1205
rect 55520 1175 55525 1205
rect 55485 1170 55525 1175
rect 55390 485 55395 1155
rect 55415 485 55420 1155
rect 55285 465 55325 470
rect 55285 435 55290 465
rect 55320 435 55325 465
rect 55285 430 55325 435
rect 55390 400 55420 485
rect 55490 1155 55520 1170
rect 55490 485 55495 1155
rect 55515 485 55520 1155
rect 55490 470 55520 485
rect 55590 1155 55620 1215
rect 55590 485 55595 1155
rect 55615 485 55620 1155
rect 55855 895 55875 1430
rect 55945 1425 55965 3035
rect 56035 2980 56065 3085
rect 56150 3080 56170 3220
rect 56280 3215 56310 3260
rect 56390 3215 56420 3320
rect 56445 3340 56475 3355
rect 56445 3320 56450 3340
rect 56470 3320 56475 3340
rect 56445 3260 56475 3320
rect 56500 3340 56530 3445
rect 56550 3435 56590 3440
rect 56550 3405 56555 3435
rect 56585 3405 56590 3435
rect 56550 3400 56590 3405
rect 56500 3320 56505 3340
rect 56525 3320 56530 3340
rect 56440 3255 56480 3260
rect 56440 3225 56445 3255
rect 56475 3225 56480 3255
rect 56440 3220 56480 3225
rect 56500 3215 56530 3320
rect 56555 3340 56585 3400
rect 56555 3320 56560 3340
rect 56580 3320 56585 3340
rect 56555 3305 56585 3320
rect 56610 3340 56640 3445
rect 56660 3390 56700 3395
rect 56660 3360 56665 3390
rect 56695 3360 56700 3390
rect 56660 3355 56700 3360
rect 56610 3320 56615 3340
rect 56635 3320 56640 3340
rect 56550 3300 56590 3305
rect 56550 3270 56555 3300
rect 56585 3270 56590 3300
rect 56550 3265 56590 3270
rect 56610 3215 56640 3320
rect 56665 3340 56695 3355
rect 56665 3320 56670 3340
rect 56690 3320 56695 3340
rect 56665 3260 56695 3320
rect 56720 3340 56750 3445
rect 56770 3435 56810 3440
rect 56770 3405 56775 3435
rect 56805 3405 56810 3435
rect 56770 3400 56810 3405
rect 56720 3320 56725 3340
rect 56745 3320 56750 3340
rect 56660 3255 56700 3260
rect 56660 3225 56665 3255
rect 56695 3225 56700 3255
rect 56660 3220 56700 3225
rect 56720 3215 56750 3320
rect 56775 3340 56805 3400
rect 56775 3320 56780 3340
rect 56800 3320 56805 3340
rect 56775 3305 56805 3320
rect 56830 3340 56860 3445
rect 56880 3390 56920 3395
rect 56880 3360 56885 3390
rect 56915 3360 56920 3390
rect 56880 3355 56920 3360
rect 56830 3320 56835 3340
rect 56855 3320 56860 3340
rect 56770 3300 56810 3305
rect 56770 3270 56775 3300
rect 56805 3270 56810 3300
rect 56770 3265 56810 3270
rect 56830 3215 56860 3320
rect 56885 3340 56915 3355
rect 56885 3320 56890 3340
rect 56910 3320 56915 3340
rect 56885 3260 56915 3320
rect 56940 3340 56970 3445
rect 56990 3435 57030 3440
rect 56990 3405 56995 3435
rect 57025 3405 57030 3435
rect 56990 3400 57030 3405
rect 56940 3320 56945 3340
rect 56965 3320 56970 3340
rect 56880 3255 56920 3260
rect 56880 3225 56885 3255
rect 56915 3225 56920 3255
rect 56880 3220 56920 3225
rect 56940 3215 56970 3320
rect 56995 3340 57025 3400
rect 56995 3320 57000 3340
rect 57020 3320 57025 3340
rect 56995 3305 57025 3320
rect 57050 3340 57080 3445
rect 57100 3390 57140 3395
rect 57100 3360 57105 3390
rect 57135 3360 57140 3390
rect 57100 3355 57140 3360
rect 57050 3320 57055 3340
rect 57075 3320 57080 3340
rect 56990 3300 57030 3305
rect 56990 3270 56995 3300
rect 57025 3270 57030 3300
rect 56990 3265 57030 3270
rect 57050 3215 57080 3320
rect 57105 3340 57135 3355
rect 57105 3320 57110 3340
rect 57130 3320 57135 3340
rect 57105 3260 57135 3320
rect 57160 3340 57190 3445
rect 57210 3435 57250 3440
rect 57210 3405 57215 3435
rect 57245 3405 57250 3435
rect 57210 3400 57250 3405
rect 57160 3320 57165 3340
rect 57185 3320 57190 3340
rect 57100 3255 57140 3260
rect 57100 3225 57105 3255
rect 57135 3225 57140 3255
rect 57100 3220 57140 3225
rect 57160 3215 57190 3320
rect 57215 3340 57245 3400
rect 57215 3320 57220 3340
rect 57240 3320 57245 3340
rect 57215 3305 57245 3320
rect 57270 3340 57300 3445
rect 57320 3390 57360 3395
rect 57320 3360 57325 3390
rect 57355 3360 57360 3390
rect 57320 3355 57360 3360
rect 57270 3320 57275 3340
rect 57295 3320 57300 3340
rect 57210 3300 57250 3305
rect 57210 3270 57215 3300
rect 57245 3270 57250 3300
rect 57210 3265 57250 3270
rect 57270 3215 57300 3320
rect 57325 3340 57355 3355
rect 57325 3320 57330 3340
rect 57350 3320 57355 3340
rect 57325 3260 57355 3320
rect 57380 3340 57410 3445
rect 57430 3435 57470 3440
rect 57430 3405 57435 3435
rect 57465 3405 57470 3435
rect 57430 3400 57470 3405
rect 57380 3320 57385 3340
rect 57405 3320 57410 3340
rect 57320 3255 57360 3260
rect 57320 3225 57325 3255
rect 57355 3225 57360 3255
rect 57320 3220 57360 3225
rect 57380 3215 57410 3320
rect 57435 3340 57465 3400
rect 57435 3320 57440 3340
rect 57460 3320 57465 3340
rect 57435 3305 57465 3320
rect 57490 3340 57520 3445
rect 57490 3320 57495 3340
rect 57515 3320 57520 3340
rect 57430 3300 57470 3305
rect 57430 3270 57435 3300
rect 57465 3270 57470 3300
rect 57430 3265 57470 3270
rect 57490 3280 57520 3320
rect 57490 3260 57495 3280
rect 57515 3260 57520 3280
rect 57620 3305 57660 3310
rect 57620 3275 57625 3305
rect 57655 3275 57660 3305
rect 57620 3270 57660 3275
rect 57490 3215 57520 3260
rect 56275 3210 56315 3215
rect 56275 3180 56280 3210
rect 56310 3180 56315 3210
rect 56275 3175 56315 3180
rect 56385 3210 56425 3215
rect 56385 3180 56390 3210
rect 56420 3180 56425 3210
rect 56385 3175 56425 3180
rect 56495 3210 56535 3215
rect 56495 3180 56500 3210
rect 56530 3180 56535 3210
rect 56495 3175 56535 3180
rect 56605 3210 56645 3215
rect 56605 3180 56610 3210
rect 56640 3180 56645 3210
rect 56605 3175 56645 3180
rect 56715 3210 56755 3215
rect 56715 3180 56720 3210
rect 56750 3180 56755 3210
rect 56715 3175 56755 3180
rect 56825 3210 56865 3215
rect 56825 3180 56830 3210
rect 56860 3180 56865 3210
rect 56825 3175 56865 3180
rect 56935 3210 56975 3215
rect 56935 3180 56940 3210
rect 56970 3180 56975 3210
rect 56935 3175 56975 3180
rect 57045 3210 57085 3215
rect 57045 3180 57050 3210
rect 57080 3180 57085 3210
rect 57045 3175 57085 3180
rect 57155 3210 57195 3215
rect 57155 3180 57160 3210
rect 57190 3180 57195 3210
rect 57155 3175 57195 3180
rect 57265 3210 57305 3215
rect 57265 3180 57270 3210
rect 57300 3180 57305 3210
rect 57265 3175 57305 3180
rect 57375 3210 57415 3215
rect 57375 3180 57380 3210
rect 57410 3180 57415 3210
rect 57375 3175 57415 3180
rect 57485 3210 57525 3215
rect 57485 3180 57490 3210
rect 57520 3180 57525 3210
rect 57485 3175 57525 3180
rect 56795 3150 56835 3160
rect 56795 3130 56805 3150
rect 56825 3130 56835 3150
rect 56690 3120 56730 3125
rect 56795 3120 56835 3130
rect 57070 3120 57110 3125
rect 56690 3090 56695 3120
rect 56725 3090 56730 3120
rect 56690 3085 56730 3090
rect 56140 3075 56180 3080
rect 56140 3045 56145 3075
rect 56175 3045 56180 3075
rect 56140 3040 56180 3045
rect 56250 3075 56290 3080
rect 56250 3045 56255 3075
rect 56285 3045 56290 3075
rect 56250 3040 56290 3045
rect 56360 3075 56400 3080
rect 56360 3045 56365 3075
rect 56395 3045 56400 3075
rect 56360 3040 56400 3045
rect 56470 3075 56510 3080
rect 56470 3045 56475 3075
rect 56505 3045 56510 3075
rect 56470 3040 56510 3045
rect 56580 3075 56620 3080
rect 56580 3045 56585 3075
rect 56615 3045 56620 3075
rect 56580 3040 56620 3045
rect 56085 3030 56125 3035
rect 56085 3000 56090 3030
rect 56120 3000 56125 3030
rect 56085 2995 56125 3000
rect 56035 2960 56040 2980
rect 56060 2960 56065 2980
rect 56035 2920 56065 2960
rect 56035 2900 56040 2920
rect 56060 2900 56065 2920
rect 56090 2980 56120 2995
rect 56090 2960 56095 2980
rect 56115 2960 56120 2980
rect 56090 2900 56120 2960
rect 56145 2980 56175 3040
rect 56195 3030 56235 3035
rect 56195 3000 56200 3030
rect 56230 3000 56235 3030
rect 56195 2995 56235 3000
rect 56145 2960 56150 2980
rect 56170 2960 56175 2980
rect 56145 2945 56175 2960
rect 56200 2980 56230 2995
rect 56200 2960 56205 2980
rect 56225 2960 56230 2980
rect 56140 2940 56180 2945
rect 56140 2910 56145 2940
rect 56175 2910 56180 2940
rect 56140 2905 56180 2910
rect 56200 2900 56230 2960
rect 56255 2980 56285 3040
rect 56305 3030 56345 3035
rect 56305 3000 56310 3030
rect 56340 3000 56345 3030
rect 56305 2995 56345 3000
rect 56255 2960 56260 2980
rect 56280 2960 56285 2980
rect 56255 2945 56285 2960
rect 56310 2980 56340 2995
rect 56310 2960 56315 2980
rect 56335 2960 56340 2980
rect 56250 2940 56290 2945
rect 56250 2910 56255 2940
rect 56285 2910 56290 2940
rect 56250 2905 56290 2910
rect 56310 2900 56340 2960
rect 56365 2980 56395 3040
rect 56415 3030 56455 3035
rect 56415 3000 56420 3030
rect 56450 3000 56455 3030
rect 56415 2995 56455 3000
rect 56365 2960 56370 2980
rect 56390 2960 56395 2980
rect 56365 2945 56395 2960
rect 56420 2980 56450 2995
rect 56420 2960 56425 2980
rect 56445 2960 56450 2980
rect 56360 2940 56400 2945
rect 56360 2910 56365 2940
rect 56395 2910 56400 2940
rect 56360 2905 56400 2910
rect 56420 2900 56450 2960
rect 56475 2980 56505 3040
rect 56525 3030 56565 3035
rect 56525 3000 56530 3030
rect 56560 3000 56565 3030
rect 56525 2995 56565 3000
rect 56475 2960 56480 2980
rect 56500 2960 56505 2980
rect 56475 2945 56505 2960
rect 56530 2980 56560 2995
rect 56530 2960 56535 2980
rect 56555 2960 56560 2980
rect 56470 2940 56510 2945
rect 56470 2910 56475 2940
rect 56505 2910 56510 2940
rect 56470 2905 56510 2910
rect 56530 2900 56560 2960
rect 56585 2980 56615 3040
rect 56635 3030 56675 3035
rect 56635 3000 56640 3030
rect 56670 3000 56675 3030
rect 56635 2995 56675 3000
rect 56585 2960 56590 2980
rect 56610 2960 56615 2980
rect 56585 2945 56615 2960
rect 56640 2980 56670 2995
rect 56640 2960 56645 2980
rect 56665 2960 56670 2980
rect 56580 2940 56620 2945
rect 56580 2910 56585 2940
rect 56615 2910 56620 2940
rect 56580 2905 56620 2910
rect 56640 2900 56670 2960
rect 56695 2980 56725 3085
rect 56740 3070 56770 3075
rect 56740 3035 56770 3040
rect 56695 2960 56700 2980
rect 56720 2960 56725 2980
rect 56695 2920 56725 2960
rect 56695 2900 56700 2920
rect 56720 2900 56725 2920
rect 56805 2900 56825 3120
rect 57070 3090 57075 3120
rect 57105 3090 57110 3120
rect 57070 3085 57110 3090
rect 57030 3070 57060 3075
rect 57030 3035 57060 3040
rect 57075 2980 57105 3085
rect 57630 3080 57650 3270
rect 57730 3120 57770 3125
rect 57730 3090 57735 3120
rect 57765 3090 57770 3120
rect 57730 3085 57770 3090
rect 57180 3075 57220 3080
rect 57180 3045 57185 3075
rect 57215 3045 57220 3075
rect 57180 3040 57220 3045
rect 57290 3075 57330 3080
rect 57290 3045 57295 3075
rect 57325 3045 57330 3075
rect 57290 3040 57330 3045
rect 57400 3075 57440 3080
rect 57400 3045 57405 3075
rect 57435 3045 57440 3075
rect 57400 3040 57440 3045
rect 57510 3075 57550 3080
rect 57510 3045 57515 3075
rect 57545 3045 57550 3075
rect 57510 3040 57550 3045
rect 57620 3075 57660 3080
rect 57620 3045 57625 3075
rect 57655 3045 57660 3075
rect 57620 3040 57660 3045
rect 57125 3030 57165 3035
rect 57125 3000 57130 3030
rect 57160 3000 57165 3030
rect 57125 2995 57165 3000
rect 57075 2960 57080 2980
rect 57100 2960 57105 2980
rect 57075 2920 57105 2960
rect 57075 2900 57080 2920
rect 57100 2900 57105 2920
rect 57130 2980 57160 2995
rect 57130 2960 57135 2980
rect 57155 2960 57160 2980
rect 57130 2900 57160 2960
rect 57185 2980 57215 3040
rect 57185 2960 57190 2980
rect 57210 2960 57215 2980
rect 57185 2945 57215 2960
rect 57240 2980 57270 2990
rect 57240 2960 57245 2980
rect 57265 2960 57270 2980
rect 57180 2940 57220 2945
rect 57180 2910 57185 2940
rect 57215 2910 57220 2940
rect 57180 2905 57220 2910
rect 56035 2800 56065 2900
rect 56085 2895 56125 2900
rect 56085 2865 56090 2895
rect 56120 2865 56125 2895
rect 56085 2860 56125 2865
rect 56195 2895 56235 2900
rect 56195 2865 56200 2895
rect 56230 2865 56235 2895
rect 56195 2860 56235 2865
rect 56305 2895 56345 2900
rect 56305 2865 56310 2895
rect 56340 2865 56345 2895
rect 56305 2860 56345 2865
rect 56415 2895 56455 2900
rect 56415 2865 56420 2895
rect 56450 2865 56455 2895
rect 56415 2860 56455 2865
rect 56525 2895 56565 2900
rect 56525 2865 56530 2895
rect 56560 2865 56565 2895
rect 56525 2860 56565 2865
rect 56635 2895 56675 2900
rect 56635 2865 56640 2895
rect 56670 2865 56675 2895
rect 56635 2860 56675 2865
rect 56095 2840 56125 2845
rect 56095 2805 56125 2810
rect 56580 2840 56610 2845
rect 56580 2805 56610 2810
rect 56695 2800 56725 2900
rect 56795 2895 56835 2900
rect 56795 2865 56800 2895
rect 56830 2865 56835 2895
rect 56795 2860 56835 2865
rect 57075 2800 57105 2900
rect 57125 2895 57165 2900
rect 57125 2865 57130 2895
rect 57160 2865 57165 2895
rect 57125 2860 57165 2865
rect 57190 2840 57220 2845
rect 57190 2805 57220 2810
rect 56030 2795 56070 2800
rect 56030 2765 56035 2795
rect 56065 2765 56070 2795
rect 56030 2760 56070 2765
rect 56690 2795 56730 2800
rect 56690 2765 56695 2795
rect 56725 2765 56730 2795
rect 56690 2760 56730 2765
rect 57070 2795 57110 2800
rect 57070 2765 57075 2795
rect 57105 2765 57110 2795
rect 57070 2760 57110 2765
rect 57240 2740 57270 2960
rect 57295 2980 57325 3040
rect 57345 3030 57385 3035
rect 57345 3000 57350 3030
rect 57380 3000 57385 3030
rect 57345 2995 57385 3000
rect 57295 2960 57300 2980
rect 57320 2960 57325 2980
rect 57295 2945 57325 2960
rect 57350 2980 57380 2995
rect 57350 2960 57355 2980
rect 57375 2960 57380 2980
rect 57290 2940 57330 2945
rect 57290 2910 57295 2940
rect 57325 2910 57330 2940
rect 57290 2905 57330 2910
rect 57350 2900 57380 2960
rect 57405 2980 57435 3040
rect 57405 2960 57410 2980
rect 57430 2960 57435 2980
rect 57405 2945 57435 2960
rect 57460 2980 57490 2990
rect 57460 2960 57465 2980
rect 57485 2960 57490 2980
rect 57400 2940 57440 2945
rect 57400 2910 57405 2940
rect 57435 2910 57440 2940
rect 57400 2905 57440 2910
rect 57345 2895 57385 2900
rect 57345 2865 57350 2895
rect 57380 2865 57385 2895
rect 57345 2860 57385 2865
rect 56605 2735 56645 2740
rect 56605 2705 56610 2735
rect 56640 2705 56645 2735
rect 56605 2700 56645 2705
rect 56825 2735 56865 2740
rect 56825 2705 56830 2735
rect 56860 2705 56865 2735
rect 56825 2700 56865 2705
rect 57045 2735 57085 2740
rect 57045 2705 57050 2735
rect 57080 2705 57085 2735
rect 57045 2700 57085 2705
rect 57235 2735 57275 2740
rect 57235 2705 57240 2735
rect 57270 2705 57275 2735
rect 57235 2700 57275 2705
rect 56550 2680 56590 2685
rect 56550 2650 56555 2680
rect 56585 2650 56590 2680
rect 56550 2645 56590 2650
rect 56305 2640 56345 2645
rect 56305 2610 56310 2640
rect 56340 2610 56345 2640
rect 56305 2605 56345 2610
rect 56030 2315 56070 2320
rect 56030 2285 56035 2315
rect 56065 2285 56070 2315
rect 56030 2280 56070 2285
rect 56035 2175 56065 2280
rect 56140 2260 56180 2265
rect 56140 2230 56145 2260
rect 56175 2230 56180 2260
rect 56140 2225 56180 2230
rect 56250 2260 56290 2265
rect 56250 2230 56255 2260
rect 56285 2230 56290 2260
rect 56250 2225 56290 2230
rect 56085 2215 56125 2220
rect 56085 2185 56090 2215
rect 56120 2185 56125 2215
rect 56085 2180 56125 2185
rect 56030 2165 56065 2175
rect 56030 2045 56040 2165
rect 56060 2045 56065 2165
rect 56030 2035 56065 2045
rect 56035 2030 56065 2035
rect 56090 2165 56120 2180
rect 56090 2045 56095 2165
rect 56115 2045 56120 2165
rect 56035 2005 56065 2015
rect 56035 1985 56040 2005
rect 56060 1985 56065 2005
rect 56090 1985 56120 2045
rect 56145 2165 56175 2225
rect 56195 2215 56235 2220
rect 56195 2185 56200 2215
rect 56230 2185 56235 2215
rect 56195 2180 56235 2185
rect 56145 2045 56150 2165
rect 56170 2045 56175 2165
rect 56145 2030 56175 2045
rect 56200 2165 56230 2180
rect 56200 2045 56205 2165
rect 56225 2045 56230 2165
rect 56140 2025 56180 2030
rect 56140 1995 56145 2025
rect 56175 1995 56180 2025
rect 56140 1990 56180 1995
rect 56200 1985 56230 2045
rect 56255 2165 56285 2225
rect 56315 2220 56335 2605
rect 56555 2570 56585 2645
rect 56555 2550 56560 2570
rect 56580 2550 56585 2570
rect 56555 2520 56585 2550
rect 56610 2570 56640 2700
rect 56660 2680 56700 2685
rect 56660 2650 56665 2680
rect 56695 2650 56700 2680
rect 56660 2645 56700 2650
rect 56770 2680 56810 2685
rect 56770 2650 56775 2680
rect 56805 2650 56810 2680
rect 56770 2645 56810 2650
rect 56610 2550 56615 2570
rect 56635 2550 56640 2570
rect 56550 2515 56590 2520
rect 56550 2485 56555 2515
rect 56585 2485 56590 2515
rect 56550 2480 56590 2485
rect 56610 2465 56640 2550
rect 56665 2570 56695 2645
rect 56715 2635 56755 2640
rect 56715 2605 56720 2635
rect 56750 2605 56755 2635
rect 56715 2600 56755 2605
rect 56665 2550 56670 2570
rect 56690 2550 56695 2570
rect 56665 2520 56695 2550
rect 56720 2570 56750 2600
rect 56720 2550 56725 2570
rect 56745 2550 56750 2570
rect 56660 2515 56700 2520
rect 56660 2485 56665 2515
rect 56695 2485 56700 2515
rect 56660 2480 56700 2485
rect 56605 2460 56645 2465
rect 56605 2430 56610 2460
rect 56640 2430 56645 2460
rect 56605 2425 56645 2430
rect 56720 2420 56750 2550
rect 56775 2570 56805 2645
rect 56775 2550 56780 2570
rect 56800 2550 56805 2570
rect 56775 2520 56805 2550
rect 56830 2570 56860 2700
rect 56880 2680 56920 2685
rect 56880 2650 56885 2680
rect 56915 2650 56920 2680
rect 56880 2645 56920 2650
rect 56990 2680 57030 2685
rect 56990 2650 56995 2680
rect 57025 2650 57030 2680
rect 56990 2645 57030 2650
rect 56830 2550 56835 2570
rect 56855 2550 56860 2570
rect 56770 2515 56810 2520
rect 56770 2485 56775 2515
rect 56805 2485 56810 2515
rect 56770 2480 56810 2485
rect 56830 2465 56860 2550
rect 56885 2570 56915 2645
rect 56935 2635 56975 2640
rect 56935 2605 56940 2635
rect 56970 2605 56975 2635
rect 56935 2600 56975 2605
rect 56885 2550 56890 2570
rect 56910 2550 56915 2570
rect 56885 2520 56915 2550
rect 56940 2570 56970 2600
rect 56940 2550 56945 2570
rect 56965 2550 56970 2570
rect 56880 2515 56920 2520
rect 56880 2485 56885 2515
rect 56915 2485 56920 2515
rect 56880 2480 56920 2485
rect 56825 2460 56865 2465
rect 56825 2430 56830 2460
rect 56860 2430 56865 2460
rect 56825 2425 56865 2430
rect 56940 2420 56970 2550
rect 56995 2570 57025 2645
rect 56995 2550 57000 2570
rect 57020 2550 57025 2570
rect 56995 2520 57025 2550
rect 57050 2570 57080 2700
rect 57100 2680 57140 2685
rect 57100 2650 57105 2680
rect 57135 2650 57140 2680
rect 57100 2645 57140 2650
rect 57210 2680 57250 2685
rect 57210 2650 57215 2680
rect 57245 2650 57250 2680
rect 57210 2645 57250 2650
rect 57050 2550 57055 2570
rect 57075 2550 57080 2570
rect 56990 2515 57030 2520
rect 56990 2485 56995 2515
rect 57025 2485 57030 2515
rect 56990 2480 57030 2485
rect 57050 2465 57080 2550
rect 57105 2570 57135 2645
rect 57155 2635 57195 2640
rect 57155 2605 57160 2635
rect 57190 2605 57195 2635
rect 57155 2600 57195 2605
rect 57105 2550 57110 2570
rect 57130 2550 57135 2570
rect 57105 2520 57135 2550
rect 57160 2570 57190 2600
rect 57160 2550 57165 2570
rect 57185 2550 57190 2570
rect 57100 2515 57140 2520
rect 57100 2485 57105 2515
rect 57135 2485 57140 2515
rect 57100 2480 57140 2485
rect 57045 2460 57085 2465
rect 57045 2430 57050 2460
rect 57080 2430 57085 2460
rect 57045 2425 57085 2430
rect 57160 2420 57190 2550
rect 57215 2570 57245 2645
rect 57350 2640 57380 2860
rect 57460 2740 57490 2960
rect 57515 2980 57545 3040
rect 57565 3030 57605 3035
rect 57565 3000 57570 3030
rect 57600 3000 57605 3030
rect 57565 2995 57605 3000
rect 57515 2960 57520 2980
rect 57540 2960 57545 2980
rect 57515 2945 57545 2960
rect 57570 2980 57600 2995
rect 57570 2960 57575 2980
rect 57595 2960 57600 2980
rect 57510 2940 57550 2945
rect 57510 2910 57515 2940
rect 57545 2910 57550 2940
rect 57510 2905 57550 2910
rect 57570 2900 57600 2960
rect 57625 2980 57655 3040
rect 57625 2960 57630 2980
rect 57650 2960 57655 2980
rect 57625 2945 57655 2960
rect 57680 2980 57710 2990
rect 57680 2960 57685 2980
rect 57705 2960 57710 2980
rect 57620 2940 57660 2945
rect 57620 2910 57625 2940
rect 57655 2910 57660 2940
rect 57620 2905 57660 2910
rect 57565 2895 57605 2900
rect 57565 2865 57570 2895
rect 57600 2865 57605 2895
rect 57565 2860 57605 2865
rect 57680 2740 57710 2960
rect 57735 2980 57765 3085
rect 57780 3070 57810 3075
rect 57780 3035 57810 3040
rect 57825 3070 57865 3075
rect 57825 3040 57830 3070
rect 57860 3040 57865 3070
rect 57825 3035 57865 3040
rect 57735 2960 57740 2980
rect 57760 2960 57765 2980
rect 57735 2920 57765 2960
rect 57735 2900 57740 2920
rect 57760 2900 57765 2920
rect 57735 2800 57765 2900
rect 57730 2795 57770 2800
rect 57730 2765 57735 2795
rect 57765 2765 57770 2795
rect 57730 2760 57770 2765
rect 57455 2735 57495 2740
rect 57455 2705 57460 2735
rect 57490 2705 57495 2735
rect 57455 2700 57495 2705
rect 57675 2735 57715 2740
rect 57675 2705 57680 2735
rect 57710 2705 57715 2735
rect 57675 2700 57715 2705
rect 57455 2640 57495 2645
rect 57345 2635 57385 2640
rect 57345 2605 57350 2635
rect 57380 2605 57385 2635
rect 57455 2610 57460 2640
rect 57490 2610 57495 2640
rect 57455 2605 57495 2610
rect 57345 2600 57385 2605
rect 57215 2550 57220 2570
rect 57240 2550 57245 2570
rect 57215 2520 57245 2550
rect 57210 2515 57250 2520
rect 57210 2485 57215 2515
rect 57245 2485 57250 2515
rect 57210 2480 57250 2485
rect 56715 2415 56755 2420
rect 56715 2385 56720 2415
rect 56750 2385 56755 2415
rect 56715 2380 56755 2385
rect 56935 2415 56975 2420
rect 56935 2385 56940 2415
rect 56970 2385 56975 2415
rect 56935 2380 56975 2385
rect 57155 2415 57195 2420
rect 57155 2385 57160 2415
rect 57190 2385 57195 2415
rect 57155 2380 57195 2385
rect 56690 2315 56730 2320
rect 56690 2285 56695 2315
rect 56725 2285 56730 2315
rect 56690 2280 56730 2285
rect 57070 2315 57110 2320
rect 57070 2285 57075 2315
rect 57105 2285 57110 2315
rect 57070 2280 57110 2285
rect 56635 2270 56665 2275
rect 56360 2260 56400 2265
rect 56360 2230 56365 2260
rect 56395 2230 56400 2260
rect 56360 2225 56400 2230
rect 56470 2260 56510 2265
rect 56470 2230 56475 2260
rect 56505 2230 56510 2260
rect 56470 2225 56510 2230
rect 56580 2260 56620 2265
rect 56580 2230 56585 2260
rect 56615 2230 56620 2260
rect 56635 2235 56665 2240
rect 56580 2225 56620 2230
rect 56305 2215 56345 2220
rect 56305 2185 56310 2215
rect 56340 2185 56345 2215
rect 56305 2180 56345 2185
rect 56255 2045 56260 2165
rect 56280 2045 56285 2165
rect 56255 2030 56285 2045
rect 56310 2165 56340 2180
rect 56310 2045 56315 2165
rect 56335 2045 56340 2165
rect 56250 2025 56290 2030
rect 56250 1995 56255 2025
rect 56285 1995 56290 2025
rect 56250 1990 56290 1995
rect 56310 1985 56340 2045
rect 56365 2165 56395 2225
rect 56415 2215 56455 2220
rect 56415 2185 56420 2215
rect 56450 2185 56455 2215
rect 56415 2180 56455 2185
rect 56365 2045 56370 2165
rect 56390 2045 56395 2165
rect 56365 2030 56395 2045
rect 56420 2165 56450 2180
rect 56420 2045 56425 2165
rect 56445 2045 56450 2165
rect 56360 2025 56400 2030
rect 56360 1995 56365 2025
rect 56395 1995 56400 2025
rect 56360 1990 56400 1995
rect 56035 1940 56065 1985
rect 56085 1980 56125 1985
rect 56085 1950 56090 1980
rect 56120 1950 56125 1980
rect 56085 1945 56125 1950
rect 56195 1980 56235 1985
rect 56195 1950 56200 1980
rect 56230 1950 56235 1980
rect 56195 1945 56235 1950
rect 56305 1980 56345 1985
rect 56305 1950 56310 1980
rect 56340 1950 56345 1980
rect 56305 1945 56345 1950
rect 56030 1935 56070 1940
rect 56030 1905 56035 1935
rect 56065 1905 56070 1935
rect 56030 1900 56070 1905
rect 56030 1850 56070 1855
rect 56030 1820 56035 1850
rect 56065 1820 56070 1850
rect 56030 1815 56070 1820
rect 55990 1785 56020 1790
rect 55990 1750 56020 1755
rect 56035 1695 56065 1815
rect 56370 1810 56390 1990
rect 56420 1985 56450 2045
rect 56475 2165 56505 2225
rect 56525 2215 56565 2220
rect 56525 2185 56530 2215
rect 56560 2185 56565 2215
rect 56525 2180 56565 2185
rect 56475 2045 56480 2165
rect 56500 2045 56505 2165
rect 56475 2030 56505 2045
rect 56530 2165 56560 2180
rect 56530 2045 56535 2165
rect 56555 2045 56560 2165
rect 56470 2025 56510 2030
rect 56470 1995 56475 2025
rect 56505 1995 56510 2025
rect 56470 1990 56510 1995
rect 56530 1985 56560 2045
rect 56585 2165 56615 2225
rect 56635 2215 56675 2220
rect 56635 2185 56640 2215
rect 56670 2185 56675 2215
rect 56635 2180 56675 2185
rect 56585 2045 56590 2165
rect 56610 2045 56615 2165
rect 56585 2030 56615 2045
rect 56640 2165 56670 2180
rect 56640 2045 56645 2165
rect 56665 2045 56670 2165
rect 56580 2025 56620 2030
rect 56580 1995 56585 2025
rect 56615 1995 56620 2025
rect 56580 1990 56620 1995
rect 56640 1985 56670 2045
rect 56695 2175 56725 2280
rect 57075 2175 57105 2280
rect 57135 2270 57165 2275
rect 57135 2235 57165 2240
rect 57180 2260 57220 2265
rect 57180 2230 57185 2260
rect 57215 2230 57220 2260
rect 57180 2225 57220 2230
rect 57290 2260 57330 2265
rect 57290 2230 57295 2260
rect 57325 2230 57330 2260
rect 57290 2225 57330 2230
rect 57400 2260 57440 2265
rect 57400 2230 57405 2260
rect 57435 2230 57440 2260
rect 57400 2225 57440 2230
rect 57125 2215 57165 2220
rect 57125 2185 57130 2215
rect 57160 2185 57165 2215
rect 57125 2180 57165 2185
rect 56695 2165 56765 2175
rect 56695 2045 56700 2165
rect 56720 2045 56765 2165
rect 56695 2035 56765 2045
rect 57035 2165 57105 2175
rect 57035 2045 57080 2165
rect 57100 2045 57105 2165
rect 57035 2035 57105 2045
rect 56695 2005 56725 2035
rect 56695 1985 56700 2005
rect 56720 1985 56725 2005
rect 56415 1980 56455 1985
rect 56415 1950 56420 1980
rect 56450 1950 56455 1980
rect 56415 1945 56455 1950
rect 56525 1980 56565 1985
rect 56525 1950 56530 1980
rect 56560 1950 56565 1980
rect 56525 1945 56565 1950
rect 56635 1980 56675 1985
rect 56635 1950 56640 1980
rect 56670 1950 56675 1980
rect 56635 1945 56675 1950
rect 56695 1940 56725 1985
rect 57075 2005 57105 2035
rect 57075 1985 57080 2005
rect 57100 1985 57105 2005
rect 57130 2165 57160 2180
rect 57130 2045 57135 2165
rect 57155 2045 57160 2165
rect 57130 1985 57160 2045
rect 57185 2165 57215 2225
rect 57235 2215 57275 2220
rect 57235 2185 57240 2215
rect 57270 2185 57275 2215
rect 57235 2180 57275 2185
rect 57185 2045 57190 2165
rect 57210 2045 57215 2165
rect 57185 2030 57215 2045
rect 57240 2165 57270 2180
rect 57240 2045 57245 2165
rect 57265 2045 57270 2165
rect 57180 2025 57220 2030
rect 57180 1995 57185 2025
rect 57215 1995 57220 2025
rect 57180 1990 57220 1995
rect 57240 1985 57270 2045
rect 57295 2165 57325 2225
rect 57345 2215 57385 2220
rect 57345 2185 57350 2215
rect 57380 2185 57385 2215
rect 57345 2180 57385 2185
rect 57295 2045 57300 2165
rect 57320 2045 57325 2165
rect 57295 2030 57325 2045
rect 57350 2165 57380 2180
rect 57350 2045 57355 2165
rect 57375 2045 57380 2165
rect 57290 2025 57330 2030
rect 57290 1995 57295 2025
rect 57325 1995 57330 2025
rect 57290 1990 57330 1995
rect 57350 1985 57380 2045
rect 57405 2165 57435 2225
rect 57465 2220 57485 2605
rect 57730 2315 57770 2320
rect 57730 2285 57735 2315
rect 57765 2285 57770 2315
rect 57730 2280 57770 2285
rect 57510 2260 57550 2265
rect 57510 2230 57515 2260
rect 57545 2230 57550 2260
rect 57510 2225 57550 2230
rect 57620 2260 57660 2265
rect 57620 2230 57625 2260
rect 57655 2230 57660 2260
rect 57620 2225 57660 2230
rect 57455 2215 57495 2220
rect 57455 2185 57460 2215
rect 57490 2185 57495 2215
rect 57455 2180 57495 2185
rect 57405 2045 57410 2165
rect 57430 2045 57435 2165
rect 57405 2030 57435 2045
rect 57460 2165 57490 2180
rect 57460 2045 57465 2165
rect 57485 2045 57490 2165
rect 57400 2025 57440 2030
rect 57400 1995 57405 2025
rect 57435 1995 57440 2025
rect 57400 1990 57440 1995
rect 57075 1940 57105 1985
rect 57125 1980 57165 1985
rect 57125 1950 57130 1980
rect 57160 1950 57165 1980
rect 57125 1945 57165 1950
rect 57235 1980 57275 1985
rect 57235 1950 57240 1980
rect 57270 1950 57275 1980
rect 57235 1945 57275 1950
rect 57345 1980 57385 1985
rect 57345 1950 57350 1980
rect 57380 1950 57385 1980
rect 57345 1945 57385 1950
rect 56690 1935 56730 1940
rect 56690 1905 56695 1935
rect 56725 1905 56730 1935
rect 56690 1900 56730 1905
rect 57070 1935 57110 1940
rect 57070 1905 57075 1935
rect 57105 1905 57110 1935
rect 57070 1900 57110 1905
rect 56730 1850 56770 1855
rect 56730 1820 56735 1850
rect 56765 1820 56770 1850
rect 57030 1850 57070 1855
rect 56730 1815 56770 1820
rect 56815 1840 56855 1845
rect 56365 1805 56395 1810
rect 56085 1795 56125 1800
rect 56085 1765 56090 1795
rect 56120 1765 56125 1795
rect 56085 1760 56125 1765
rect 56195 1795 56235 1800
rect 56195 1765 56200 1795
rect 56230 1765 56235 1795
rect 56195 1760 56235 1765
rect 56305 1795 56345 1800
rect 56305 1765 56310 1795
rect 56340 1765 56345 1795
rect 56365 1770 56395 1775
rect 56415 1795 56455 1800
rect 56305 1760 56345 1765
rect 56415 1765 56420 1795
rect 56450 1765 56455 1795
rect 56415 1760 56455 1765
rect 56525 1795 56565 1800
rect 56525 1765 56530 1795
rect 56560 1765 56565 1795
rect 56525 1760 56565 1765
rect 56635 1795 56675 1800
rect 56635 1765 56640 1795
rect 56670 1765 56675 1795
rect 56635 1760 56675 1765
rect 56690 1785 56720 1790
rect 56035 1575 56040 1695
rect 56060 1575 56065 1695
rect 56035 1535 56065 1575
rect 56090 1695 56120 1760
rect 56140 1750 56180 1755
rect 56140 1720 56145 1750
rect 56175 1720 56180 1750
rect 56140 1715 56180 1720
rect 56090 1575 56095 1695
rect 56115 1575 56120 1695
rect 56090 1560 56120 1575
rect 56145 1695 56175 1715
rect 56145 1575 56150 1695
rect 56170 1575 56175 1695
rect 56035 1515 56040 1535
rect 56060 1515 56065 1535
rect 56085 1555 56125 1560
rect 56085 1525 56090 1555
rect 56120 1525 56125 1555
rect 56085 1520 56125 1525
rect 56145 1515 56175 1575
rect 56200 1695 56230 1760
rect 56250 1750 56290 1755
rect 56250 1720 56255 1750
rect 56285 1720 56290 1750
rect 56250 1715 56290 1720
rect 56200 1575 56205 1695
rect 56225 1575 56230 1695
rect 56200 1560 56230 1575
rect 56255 1695 56285 1715
rect 56255 1575 56260 1695
rect 56280 1575 56285 1695
rect 56195 1555 56235 1560
rect 56195 1525 56200 1555
rect 56230 1525 56235 1555
rect 56195 1520 56235 1525
rect 56255 1515 56285 1575
rect 56310 1695 56340 1760
rect 56360 1750 56400 1755
rect 56360 1720 56365 1750
rect 56395 1720 56400 1750
rect 56360 1715 56400 1720
rect 56310 1575 56315 1695
rect 56335 1575 56340 1695
rect 56310 1560 56340 1575
rect 56365 1695 56395 1715
rect 56365 1575 56370 1695
rect 56390 1575 56395 1695
rect 56305 1555 56345 1560
rect 56305 1525 56310 1555
rect 56340 1525 56345 1555
rect 56305 1520 56345 1525
rect 56365 1515 56395 1575
rect 56420 1695 56450 1760
rect 56470 1750 56510 1755
rect 56470 1720 56475 1750
rect 56505 1720 56510 1750
rect 56470 1715 56510 1720
rect 56420 1575 56425 1695
rect 56445 1575 56450 1695
rect 56420 1560 56450 1575
rect 56475 1695 56505 1715
rect 56475 1575 56480 1695
rect 56500 1575 56505 1695
rect 56415 1555 56455 1560
rect 56415 1525 56420 1555
rect 56450 1525 56455 1555
rect 56415 1520 56455 1525
rect 56475 1515 56505 1575
rect 56530 1695 56560 1760
rect 56580 1750 56620 1755
rect 56580 1720 56585 1750
rect 56615 1720 56620 1750
rect 56580 1715 56620 1720
rect 56530 1575 56535 1695
rect 56555 1575 56560 1695
rect 56530 1560 56560 1575
rect 56585 1695 56615 1715
rect 56585 1575 56590 1695
rect 56610 1575 56615 1695
rect 56525 1555 56565 1560
rect 56525 1525 56530 1555
rect 56560 1525 56565 1555
rect 56525 1520 56565 1525
rect 56585 1515 56615 1575
rect 56640 1695 56670 1760
rect 56690 1750 56720 1755
rect 56735 1705 56765 1815
rect 56815 1810 56820 1840
rect 56850 1810 56855 1840
rect 56815 1805 56855 1810
rect 56945 1840 56985 1845
rect 56945 1810 56950 1840
rect 56980 1810 56985 1840
rect 57030 1820 57035 1850
rect 57065 1820 57070 1850
rect 57030 1815 57070 1820
rect 56945 1805 56985 1810
rect 56830 1705 56845 1805
rect 56859 1785 56889 1790
rect 56859 1750 56889 1755
rect 56911 1785 56941 1790
rect 56911 1755 56914 1785
rect 56911 1750 56941 1755
rect 56955 1705 56970 1805
rect 57035 1705 57065 1815
rect 57410 1810 57430 1990
rect 57460 1985 57490 2045
rect 57515 2165 57545 2225
rect 57565 2215 57605 2220
rect 57565 2185 57570 2215
rect 57600 2185 57605 2215
rect 57565 2180 57605 2185
rect 57515 2045 57520 2165
rect 57540 2045 57545 2165
rect 57515 2030 57545 2045
rect 57570 2165 57600 2180
rect 57570 2045 57575 2165
rect 57595 2045 57600 2165
rect 57510 2025 57550 2030
rect 57510 1995 57515 2025
rect 57545 1995 57550 2025
rect 57510 1990 57550 1995
rect 57570 1985 57600 2045
rect 57625 2165 57655 2225
rect 57675 2215 57715 2220
rect 57675 2185 57680 2215
rect 57710 2185 57715 2215
rect 57675 2180 57715 2185
rect 57625 2045 57630 2165
rect 57650 2045 57655 2165
rect 57625 2030 57655 2045
rect 57680 2165 57710 2180
rect 57680 2045 57685 2165
rect 57705 2045 57710 2165
rect 57620 2025 57660 2030
rect 57620 1995 57625 2025
rect 57655 1995 57660 2025
rect 57620 1990 57660 1995
rect 57680 1985 57710 2045
rect 57735 2165 57765 2280
rect 57785 2245 57815 2250
rect 57785 2210 57815 2215
rect 57735 2045 57740 2165
rect 57760 2045 57765 2165
rect 57735 2035 57765 2045
rect 57735 2005 57765 2015
rect 57735 1985 57740 2005
rect 57760 1985 57765 2005
rect 57455 1980 57495 1985
rect 57455 1950 57460 1980
rect 57490 1950 57495 1980
rect 57455 1945 57495 1950
rect 57565 1980 57605 1985
rect 57565 1950 57570 1980
rect 57600 1950 57605 1980
rect 57565 1945 57605 1950
rect 57675 1980 57715 1985
rect 57675 1950 57680 1980
rect 57710 1950 57715 1980
rect 57675 1945 57715 1950
rect 57735 1940 57765 1985
rect 57730 1935 57770 1940
rect 57730 1905 57735 1935
rect 57765 1905 57770 1935
rect 57730 1900 57770 1905
rect 57730 1850 57770 1855
rect 57730 1820 57735 1850
rect 57765 1820 57770 1850
rect 57730 1815 57770 1820
rect 57405 1805 57435 1810
rect 57125 1795 57165 1800
rect 57080 1785 57110 1790
rect 57125 1765 57130 1795
rect 57160 1765 57165 1795
rect 57125 1760 57165 1765
rect 57235 1795 57275 1800
rect 57235 1765 57240 1795
rect 57270 1765 57275 1795
rect 57235 1760 57275 1765
rect 57345 1795 57385 1800
rect 57345 1765 57350 1795
rect 57380 1765 57385 1795
rect 57405 1770 57435 1775
rect 57455 1795 57495 1800
rect 57345 1760 57385 1765
rect 57455 1765 57460 1795
rect 57490 1765 57495 1795
rect 57455 1760 57495 1765
rect 57565 1795 57605 1800
rect 57565 1765 57570 1795
rect 57600 1765 57605 1795
rect 57565 1760 57605 1765
rect 57675 1795 57715 1800
rect 57675 1765 57680 1795
rect 57710 1765 57715 1795
rect 57675 1760 57715 1765
rect 57080 1750 57110 1755
rect 56640 1575 56645 1695
rect 56665 1575 56670 1695
rect 56640 1560 56670 1575
rect 56695 1695 56805 1705
rect 56695 1575 56700 1695
rect 56720 1575 56780 1695
rect 56800 1575 56805 1695
rect 56695 1565 56805 1575
rect 56830 1695 56860 1705
rect 56830 1575 56835 1695
rect 56855 1575 56860 1695
rect 56830 1565 56860 1575
rect 56885 1695 56915 1705
rect 56885 1575 56890 1695
rect 56910 1575 56915 1695
rect 56885 1565 56915 1575
rect 56940 1695 56970 1705
rect 56940 1575 56945 1695
rect 56965 1575 56970 1695
rect 56940 1565 56970 1575
rect 56995 1695 57105 1705
rect 56995 1575 57000 1695
rect 57020 1575 57080 1695
rect 57100 1575 57105 1695
rect 56995 1565 57105 1575
rect 57130 1695 57160 1760
rect 57180 1750 57220 1755
rect 57180 1720 57185 1750
rect 57215 1720 57220 1750
rect 57180 1715 57220 1720
rect 57130 1575 57135 1695
rect 57155 1575 57160 1695
rect 56635 1555 56675 1560
rect 56635 1525 56640 1555
rect 56670 1525 56675 1555
rect 56635 1520 56675 1525
rect 56735 1535 56765 1565
rect 56735 1515 56740 1535
rect 56760 1515 56765 1535
rect 56035 1470 56065 1515
rect 56140 1510 56180 1515
rect 56140 1480 56145 1510
rect 56175 1480 56180 1510
rect 56140 1475 56180 1480
rect 56250 1510 56290 1515
rect 56250 1480 56255 1510
rect 56285 1480 56290 1510
rect 56250 1475 56290 1480
rect 56360 1510 56400 1515
rect 56360 1480 56365 1510
rect 56395 1480 56400 1510
rect 56360 1475 56400 1480
rect 56470 1510 56510 1515
rect 56470 1480 56475 1510
rect 56505 1480 56510 1510
rect 56470 1475 56510 1480
rect 56580 1510 56620 1515
rect 56580 1480 56585 1510
rect 56615 1480 56620 1510
rect 56580 1475 56620 1480
rect 56735 1470 56765 1515
rect 56030 1465 56070 1470
rect 56030 1435 56035 1465
rect 56065 1435 56070 1465
rect 56030 1430 56070 1435
rect 56730 1465 56770 1470
rect 56730 1435 56735 1465
rect 56765 1435 56770 1465
rect 56730 1430 56770 1435
rect 56835 1425 56855 1565
rect 55935 1420 55975 1425
rect 55935 1390 55940 1420
rect 55970 1390 55975 1420
rect 55935 1385 55975 1390
rect 56825 1420 56865 1425
rect 56825 1390 56830 1420
rect 56860 1390 56865 1420
rect 56825 1385 56865 1390
rect 56330 1265 56370 1270
rect 56330 1235 56335 1265
rect 56365 1235 56370 1265
rect 56330 1230 56370 1235
rect 56185 1145 56255 1155
rect 56185 925 56230 1145
rect 56250 925 56255 1145
rect 56185 915 56255 925
rect 56225 895 56255 915
rect 56280 1145 56310 1155
rect 56280 925 56285 1145
rect 56305 925 56310 1145
rect 56280 895 56310 925
rect 56335 1145 56365 1230
rect 56835 1215 56855 1385
rect 56890 1270 56910 1565
rect 56945 1425 56965 1565
rect 57035 1535 57065 1565
rect 57130 1560 57160 1575
rect 57185 1695 57215 1715
rect 57185 1575 57190 1695
rect 57210 1575 57215 1695
rect 57035 1515 57040 1535
rect 57060 1515 57065 1535
rect 57125 1555 57165 1560
rect 57125 1525 57130 1555
rect 57160 1525 57165 1555
rect 57125 1520 57165 1525
rect 57185 1515 57215 1575
rect 57240 1695 57270 1760
rect 57290 1750 57330 1755
rect 57290 1720 57295 1750
rect 57325 1720 57330 1750
rect 57290 1715 57330 1720
rect 57240 1575 57245 1695
rect 57265 1575 57270 1695
rect 57240 1560 57270 1575
rect 57295 1695 57325 1715
rect 57295 1575 57300 1695
rect 57320 1575 57325 1695
rect 57235 1555 57275 1560
rect 57235 1525 57240 1555
rect 57270 1525 57275 1555
rect 57235 1520 57275 1525
rect 57295 1515 57325 1575
rect 57350 1695 57380 1760
rect 57400 1750 57440 1755
rect 57400 1720 57405 1750
rect 57435 1720 57440 1750
rect 57400 1715 57440 1720
rect 57350 1575 57355 1695
rect 57375 1575 57380 1695
rect 57350 1560 57380 1575
rect 57405 1695 57435 1715
rect 57405 1575 57410 1695
rect 57430 1575 57435 1695
rect 57345 1555 57385 1560
rect 57345 1525 57350 1555
rect 57380 1525 57385 1555
rect 57345 1520 57385 1525
rect 57405 1515 57435 1575
rect 57460 1695 57490 1760
rect 57510 1750 57550 1755
rect 57510 1720 57515 1750
rect 57545 1720 57550 1750
rect 57510 1715 57550 1720
rect 57460 1575 57465 1695
rect 57485 1575 57490 1695
rect 57460 1560 57490 1575
rect 57515 1695 57545 1715
rect 57515 1575 57520 1695
rect 57540 1575 57545 1695
rect 57455 1555 57495 1560
rect 57455 1525 57460 1555
rect 57490 1525 57495 1555
rect 57455 1520 57495 1525
rect 57515 1515 57545 1575
rect 57570 1695 57600 1760
rect 57620 1750 57660 1755
rect 57620 1720 57625 1750
rect 57655 1720 57660 1750
rect 57620 1715 57660 1720
rect 57570 1575 57575 1695
rect 57595 1575 57600 1695
rect 57570 1560 57600 1575
rect 57625 1695 57655 1715
rect 57625 1575 57630 1695
rect 57650 1575 57655 1695
rect 57565 1555 57605 1560
rect 57565 1525 57570 1555
rect 57600 1525 57605 1555
rect 57565 1520 57605 1525
rect 57625 1515 57655 1575
rect 57680 1695 57710 1760
rect 57680 1575 57685 1695
rect 57705 1575 57710 1695
rect 57680 1560 57710 1575
rect 57735 1695 57765 1815
rect 57780 1785 57810 1790
rect 57780 1750 57810 1755
rect 57735 1575 57740 1695
rect 57760 1575 57765 1695
rect 57675 1555 57715 1560
rect 57675 1525 57680 1555
rect 57710 1525 57715 1555
rect 57675 1520 57715 1525
rect 57735 1535 57765 1575
rect 57735 1515 57740 1535
rect 57760 1515 57765 1535
rect 57035 1470 57065 1515
rect 57180 1510 57220 1515
rect 57180 1480 57185 1510
rect 57215 1480 57220 1510
rect 57180 1475 57220 1480
rect 57290 1510 57330 1515
rect 57290 1480 57295 1510
rect 57325 1480 57330 1510
rect 57290 1475 57330 1480
rect 57400 1510 57440 1515
rect 57400 1480 57405 1510
rect 57435 1480 57440 1510
rect 57400 1475 57440 1480
rect 57510 1510 57550 1515
rect 57510 1480 57515 1510
rect 57545 1480 57550 1510
rect 57510 1475 57550 1480
rect 57620 1510 57660 1515
rect 57620 1480 57625 1510
rect 57655 1480 57660 1510
rect 57620 1475 57660 1480
rect 57030 1465 57070 1470
rect 57030 1435 57035 1465
rect 57065 1435 57070 1465
rect 57030 1430 57070 1435
rect 56935 1420 56975 1425
rect 56935 1390 56940 1420
rect 56970 1390 56975 1420
rect 56935 1385 56975 1390
rect 56880 1265 56920 1270
rect 56880 1235 56885 1265
rect 56915 1235 56920 1265
rect 56880 1230 56920 1235
rect 57200 1215 57220 1475
rect 57735 1470 57765 1515
rect 57730 1465 57770 1470
rect 57730 1435 57735 1465
rect 57765 1435 57770 1465
rect 57730 1430 57770 1435
rect 57835 1425 57855 3035
rect 58015 2800 58035 3445
rect 58005 2795 58045 2800
rect 58005 2765 58010 2795
rect 58040 2765 58045 2795
rect 58005 2760 58045 2765
rect 58015 2550 58035 2760
rect 58060 2645 58080 3605
rect 58450 3540 58490 3545
rect 58450 3510 58455 3540
rect 58485 3510 58490 3540
rect 58450 3505 58490 3510
rect 58150 3480 58190 3485
rect 58150 3450 58155 3480
rect 58185 3450 58190 3480
rect 58150 3445 58190 3450
rect 58260 3480 58300 3485
rect 58260 3450 58265 3480
rect 58295 3450 58300 3480
rect 58260 3445 58300 3450
rect 58370 3480 58410 3485
rect 58370 3450 58375 3480
rect 58405 3450 58410 3480
rect 58370 3445 58410 3450
rect 58480 3480 58520 3485
rect 58480 3450 58485 3480
rect 58515 3450 58520 3480
rect 58480 3445 58520 3450
rect 58590 3480 58630 3485
rect 58590 3450 58595 3480
rect 58625 3450 58630 3480
rect 58590 3445 58630 3450
rect 58700 3480 58740 3485
rect 58700 3450 58705 3480
rect 58735 3450 58740 3480
rect 58700 3445 58740 3450
rect 58810 3480 58850 3485
rect 58810 3450 58815 3480
rect 58845 3450 58850 3480
rect 58810 3445 58850 3450
rect 58155 3395 58185 3445
rect 58155 3375 58160 3395
rect 58180 3375 58185 3395
rect 58155 3335 58185 3375
rect 58205 3385 58245 3390
rect 58205 3355 58210 3385
rect 58240 3355 58245 3385
rect 58205 3350 58245 3355
rect 58155 2765 58160 3335
rect 58180 2765 58185 3335
rect 58155 2705 58185 2765
rect 58210 3335 58240 3350
rect 58210 2765 58215 3335
rect 58235 2765 58240 3335
rect 58210 2750 58240 2765
rect 58265 3335 58295 3445
rect 58315 3385 58355 3390
rect 58315 3355 58320 3385
rect 58350 3355 58355 3385
rect 58315 3350 58355 3355
rect 58265 2765 58270 3335
rect 58290 2765 58295 3335
rect 58205 2745 58245 2750
rect 58205 2715 58210 2745
rect 58240 2715 58245 2745
rect 58205 2710 58245 2715
rect 58265 2705 58295 2765
rect 58320 3335 58350 3350
rect 58320 2765 58325 3335
rect 58345 2765 58350 3335
rect 58320 2750 58350 2765
rect 58375 3335 58405 3445
rect 58425 3385 58465 3390
rect 58425 3355 58430 3385
rect 58460 3355 58465 3385
rect 58425 3350 58465 3355
rect 58375 2765 58380 3335
rect 58400 2765 58405 3335
rect 58315 2745 58355 2750
rect 58315 2715 58320 2745
rect 58350 2715 58355 2745
rect 58315 2710 58355 2715
rect 58150 2700 58190 2705
rect 58150 2670 58155 2700
rect 58185 2670 58190 2700
rect 58150 2665 58190 2670
rect 58260 2700 58300 2705
rect 58260 2670 58265 2700
rect 58295 2670 58300 2700
rect 58260 2665 58300 2670
rect 58050 2640 58090 2645
rect 58050 2610 58055 2640
rect 58085 2610 58090 2640
rect 58050 2605 58090 2610
rect 58005 2545 58045 2550
rect 57915 2515 57955 2520
rect 57915 2485 57920 2515
rect 57950 2485 57955 2515
rect 58005 2515 58010 2545
rect 58040 2515 58045 2545
rect 58005 2510 58045 2515
rect 57915 2480 57955 2485
rect 57870 2460 57910 2465
rect 57870 2430 57875 2460
rect 57905 2430 57910 2460
rect 57870 2425 57910 2430
rect 57825 1420 57865 1425
rect 57825 1390 57830 1420
rect 57860 1390 57865 1420
rect 57825 1385 57865 1390
rect 57880 1270 57900 2425
rect 57925 1940 57945 2480
rect 57960 2245 58000 2250
rect 57960 2215 57965 2245
rect 57995 2215 58000 2245
rect 57960 2210 58000 2215
rect 57915 1935 57955 1940
rect 57915 1905 57920 1935
rect 57950 1905 57955 1935
rect 57915 1900 57955 1905
rect 57925 1470 57945 1900
rect 57915 1465 57955 1470
rect 57915 1435 57920 1465
rect 57950 1435 57955 1465
rect 57915 1430 57955 1435
rect 57405 1265 57445 1270
rect 57405 1235 57410 1265
rect 57440 1235 57445 1265
rect 57405 1230 57445 1235
rect 57870 1265 57910 1270
rect 57870 1235 57875 1265
rect 57905 1235 57910 1265
rect 57870 1230 57910 1235
rect 56440 1210 56480 1215
rect 56440 1180 56445 1210
rect 56475 1180 56480 1210
rect 56440 1175 56480 1180
rect 56550 1210 56590 1215
rect 56550 1180 56555 1210
rect 56585 1180 56590 1210
rect 56550 1175 56590 1180
rect 56660 1210 56700 1215
rect 56660 1180 56665 1210
rect 56695 1180 56700 1210
rect 56660 1175 56700 1180
rect 56770 1210 56810 1215
rect 56770 1180 56775 1210
rect 56805 1180 56810 1210
rect 56770 1175 56810 1180
rect 56830 1205 56860 1215
rect 56830 1185 56835 1205
rect 56855 1185 56860 1205
rect 56830 1175 56860 1185
rect 56880 1210 56920 1215
rect 56880 1180 56885 1210
rect 56915 1180 56920 1210
rect 56880 1175 56920 1180
rect 56990 1210 57030 1215
rect 56990 1180 56995 1210
rect 57025 1180 57030 1210
rect 56990 1175 57030 1180
rect 57100 1210 57140 1215
rect 57100 1180 57105 1210
rect 57135 1180 57140 1210
rect 57100 1175 57140 1180
rect 57200 1210 57250 1215
rect 57200 1180 57215 1210
rect 57245 1180 57250 1210
rect 57200 1175 57250 1180
rect 57320 1210 57360 1215
rect 57320 1180 57325 1210
rect 57355 1180 57360 1210
rect 57320 1175 57360 1180
rect 57430 1210 57470 1215
rect 57430 1180 57435 1210
rect 57465 1180 57470 1210
rect 57430 1175 57470 1180
rect 56335 925 56340 1145
rect 56360 925 56365 1145
rect 56335 915 56365 925
rect 56390 1145 56420 1155
rect 56390 925 56395 1145
rect 56415 925 56420 1145
rect 56390 895 56420 925
rect 56445 1145 56475 1175
rect 56445 925 56450 1145
rect 56470 925 56475 1145
rect 55845 890 55885 895
rect 55845 860 55850 890
rect 55880 860 55885 890
rect 55845 855 55885 860
rect 56220 890 56260 895
rect 56220 860 56225 890
rect 56255 860 56260 890
rect 56220 855 56260 860
rect 56275 890 56315 895
rect 56275 860 56280 890
rect 56310 860 56315 890
rect 56275 855 56315 860
rect 56385 890 56425 895
rect 56385 860 56390 890
rect 56420 860 56425 890
rect 56385 855 56425 860
rect 55485 465 55525 470
rect 55485 435 55490 465
rect 55520 435 55525 465
rect 55485 430 55525 435
rect 55590 445 55620 485
rect 55590 425 55595 445
rect 55615 425 55620 445
rect 55590 400 55620 425
rect 55855 400 55875 855
rect 56445 850 56475 925
rect 56500 1145 56530 1155
rect 56500 925 56505 1145
rect 56525 925 56530 1145
rect 56500 895 56530 925
rect 56555 1145 56585 1175
rect 56555 925 56560 1145
rect 56580 925 56585 1145
rect 56495 890 56535 895
rect 56495 860 56500 890
rect 56530 860 56535 890
rect 56495 855 56535 860
rect 56555 850 56585 925
rect 56610 1145 56640 1155
rect 56610 925 56615 1145
rect 56635 925 56640 1145
rect 56610 895 56640 925
rect 56665 1145 56695 1175
rect 56665 925 56670 1145
rect 56690 925 56695 1145
rect 56605 890 56645 895
rect 56605 860 56610 890
rect 56640 860 56645 890
rect 56605 855 56645 860
rect 56665 850 56695 925
rect 56720 1145 56750 1155
rect 56720 925 56725 1145
rect 56745 925 56750 1145
rect 56720 895 56750 925
rect 56775 1145 56805 1175
rect 56775 925 56780 1145
rect 56800 925 56805 1145
rect 56715 890 56755 895
rect 56715 860 56720 890
rect 56750 860 56755 890
rect 56715 855 56755 860
rect 56775 850 56805 925
rect 56830 1145 56860 1155
rect 56830 925 56835 1145
rect 56855 925 56860 1145
rect 56830 895 56860 925
rect 56885 1145 56915 1175
rect 56885 925 56890 1145
rect 56910 925 56915 1145
rect 56825 890 56865 895
rect 56825 860 56830 890
rect 56860 860 56865 890
rect 56825 855 56865 860
rect 56885 850 56915 925
rect 56940 1145 56970 1155
rect 56940 925 56945 1145
rect 56965 925 56970 1145
rect 56940 895 56970 925
rect 56995 1145 57025 1175
rect 56995 925 57000 1145
rect 57020 925 57025 1145
rect 56935 890 56975 895
rect 56935 860 56940 890
rect 56970 860 56975 890
rect 56935 855 56975 860
rect 56995 850 57025 925
rect 57050 1145 57080 1155
rect 57050 925 57055 1145
rect 57075 925 57080 1145
rect 57050 895 57080 925
rect 57105 1145 57135 1175
rect 57105 925 57110 1145
rect 57130 925 57135 1145
rect 57045 890 57085 895
rect 57045 860 57050 890
rect 57080 860 57085 890
rect 57045 855 57085 860
rect 57105 850 57135 925
rect 57160 1145 57190 1155
rect 57160 925 57165 1145
rect 57185 925 57190 1145
rect 57160 895 57190 925
rect 57215 1145 57245 1175
rect 57215 925 57220 1145
rect 57240 925 57245 1145
rect 57155 890 57195 895
rect 57155 860 57160 890
rect 57190 860 57195 890
rect 57155 855 57195 860
rect 57215 850 57245 925
rect 57270 1145 57300 1155
rect 57270 925 57275 1145
rect 57295 925 57300 1145
rect 57270 895 57300 925
rect 57325 1145 57355 1175
rect 57325 925 57330 1145
rect 57350 925 57355 1145
rect 57265 890 57305 895
rect 57265 860 57270 890
rect 57300 860 57305 890
rect 57265 855 57305 860
rect 57325 850 57355 925
rect 57380 1145 57410 1155
rect 57380 925 57385 1145
rect 57405 925 57410 1145
rect 57380 895 57410 925
rect 57435 1145 57465 1175
rect 57435 925 57440 1145
rect 57460 925 57465 1145
rect 57375 890 57415 895
rect 57375 860 57380 890
rect 57410 860 57415 890
rect 57375 855 57415 860
rect 57435 850 57465 925
rect 57490 1145 57520 1155
rect 57490 925 57495 1145
rect 57515 925 57520 1145
rect 57490 895 57520 925
rect 57485 890 57525 895
rect 57485 860 57490 890
rect 57520 860 57525 890
rect 57925 885 57945 1430
rect 57485 855 57525 860
rect 57915 880 57955 885
rect 57915 850 57920 880
rect 57950 850 57955 880
rect 56440 845 56480 850
rect 56440 815 56445 845
rect 56475 815 56480 845
rect 56440 810 56480 815
rect 56550 845 56590 850
rect 56550 815 56555 845
rect 56585 815 56590 845
rect 56550 810 56590 815
rect 56660 845 56700 850
rect 56660 815 56665 845
rect 56695 815 56700 845
rect 56660 810 56700 815
rect 56770 845 56810 850
rect 56770 815 56775 845
rect 56805 815 56810 845
rect 56770 810 56810 815
rect 56880 845 56920 850
rect 56880 815 56885 845
rect 56915 815 56920 845
rect 56880 810 56920 815
rect 56990 845 57030 850
rect 56990 815 56995 845
rect 57025 815 57030 845
rect 56990 810 57030 815
rect 57100 845 57140 850
rect 57100 815 57105 845
rect 57135 815 57140 845
rect 57100 810 57140 815
rect 57210 845 57250 850
rect 57210 815 57215 845
rect 57245 815 57250 845
rect 57210 810 57250 815
rect 57320 845 57360 850
rect 57320 815 57325 845
rect 57355 815 57360 845
rect 57320 810 57360 815
rect 57430 845 57470 850
rect 57915 845 57955 850
rect 57430 815 57435 845
rect 57465 815 57470 845
rect 57430 810 57470 815
rect 56540 790 56580 795
rect 56540 760 56545 790
rect 56575 760 56580 790
rect 56540 755 56580 760
rect 56650 790 56690 795
rect 56650 760 56655 790
rect 56685 760 56690 790
rect 56650 755 56690 760
rect 56870 790 56910 795
rect 56870 760 56875 790
rect 56905 760 56910 790
rect 56870 755 56910 760
rect 56485 745 56525 750
rect 56485 715 56490 745
rect 56520 715 56525 745
rect 56485 710 56525 715
rect 56395 680 56465 690
rect 56395 560 56440 680
rect 56460 560 56465 680
rect 56395 550 56465 560
rect 56435 520 56465 550
rect 56435 500 56440 520
rect 56460 500 56465 520
rect 56490 680 56520 710
rect 56490 560 56495 680
rect 56515 560 56520 680
rect 56490 500 56520 560
rect 56545 680 56575 755
rect 56595 745 56635 750
rect 56595 715 56600 745
rect 56630 715 56635 745
rect 56595 710 56635 715
rect 56545 560 56550 680
rect 56570 560 56575 680
rect 56545 545 56575 560
rect 56600 680 56630 710
rect 56600 560 56605 680
rect 56625 560 56630 680
rect 56540 540 56580 545
rect 56540 510 56545 540
rect 56575 510 56580 540
rect 56540 505 56580 510
rect 56600 500 56630 560
rect 56655 680 56685 755
rect 56705 745 56745 750
rect 56705 715 56710 745
rect 56740 715 56745 745
rect 56705 710 56745 715
rect 56655 560 56660 680
rect 56680 560 56685 680
rect 56655 545 56685 560
rect 56710 680 56740 710
rect 56710 560 56715 680
rect 56735 560 56740 680
rect 56650 540 56690 545
rect 56650 510 56655 540
rect 56685 510 56690 540
rect 56650 505 56690 510
rect 56710 500 56740 560
rect 56765 680 56835 690
rect 56765 560 56770 680
rect 56790 560 56835 680
rect 56765 550 56835 560
rect 56875 680 56905 755
rect 57040 745 57080 750
rect 57040 715 57045 745
rect 57075 715 57080 745
rect 57040 710 57080 715
rect 56875 560 56880 680
rect 56900 560 56905 680
rect 56765 520 56795 550
rect 56875 545 56905 560
rect 57215 680 57245 810
rect 57215 560 57220 680
rect 57240 560 57245 680
rect 57215 550 57245 560
rect 56765 500 56770 520
rect 56790 500 56795 520
rect 56870 540 56910 545
rect 56870 510 56875 540
rect 56905 510 56910 540
rect 56870 505 56910 510
rect 56435 400 56465 500
rect 56485 495 56525 500
rect 56485 465 56490 495
rect 56520 465 56525 495
rect 56485 460 56525 465
rect 56595 495 56635 500
rect 56595 465 56600 495
rect 56630 465 56635 495
rect 56595 460 56635 465
rect 56705 495 56745 500
rect 56705 465 56710 495
rect 56740 465 56745 495
rect 56705 460 56745 465
rect 56765 400 56795 500
rect 57925 400 57945 845
rect 57970 750 57990 2210
rect 58015 1515 58035 2510
rect 58060 2055 58080 2605
rect 58325 2600 58345 2710
rect 58375 2705 58405 2765
rect 58430 3335 58460 3350
rect 58430 2765 58435 3335
rect 58455 2765 58460 3335
rect 58430 2750 58460 2765
rect 58485 3335 58515 3445
rect 58535 3385 58575 3390
rect 58535 3355 58540 3385
rect 58570 3355 58575 3385
rect 58535 3350 58575 3355
rect 58485 2765 58490 3335
rect 58510 2765 58515 3335
rect 58425 2745 58465 2750
rect 58425 2715 58430 2745
rect 58460 2715 58465 2745
rect 58425 2710 58465 2715
rect 58485 2705 58515 2765
rect 58540 3335 58570 3350
rect 58540 2765 58545 3335
rect 58565 2765 58570 3335
rect 58540 2750 58570 2765
rect 58595 3335 58625 3445
rect 58645 3385 58685 3390
rect 58645 3355 58650 3385
rect 58680 3355 58685 3385
rect 58645 3350 58685 3355
rect 58595 2765 58600 3335
rect 58620 2765 58625 3335
rect 58535 2745 58575 2750
rect 58535 2715 58540 2745
rect 58570 2715 58575 2745
rect 58535 2710 58575 2715
rect 58595 2705 58625 2765
rect 58650 3335 58680 3350
rect 58650 2765 58655 3335
rect 58675 2765 58680 3335
rect 58650 2750 58680 2765
rect 58705 3335 58735 3445
rect 58815 3395 58845 3445
rect 58755 3385 58795 3390
rect 58755 3355 58760 3385
rect 58790 3355 58795 3385
rect 58755 3350 58795 3355
rect 58815 3375 58820 3395
rect 58840 3375 58845 3395
rect 58705 2765 58710 3335
rect 58730 2765 58735 3335
rect 58645 2745 58685 2750
rect 58645 2715 58650 2745
rect 58680 2715 58685 2745
rect 58645 2710 58685 2715
rect 58705 2705 58735 2765
rect 58760 3335 58790 3350
rect 58760 2765 58765 3335
rect 58785 2765 58790 3335
rect 58760 2750 58790 2765
rect 58815 3335 58845 3375
rect 59155 3400 59195 3405
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58815 2765 58820 3335
rect 58840 2765 58845 3335
rect 59165 3325 59185 3365
rect 59105 3315 59246 3325
rect 59105 3295 59110 3315
rect 59130 3295 59165 3315
rect 59185 3295 59220 3315
rect 59240 3295 59246 3315
rect 59105 3285 59246 3295
rect 58755 2745 58795 2750
rect 58755 2715 58760 2745
rect 58790 2715 58795 2745
rect 58755 2710 58795 2715
rect 58815 2705 58845 2765
rect 59105 2710 59246 2720
rect 58370 2700 58410 2705
rect 58370 2670 58375 2700
rect 58405 2670 58410 2700
rect 58370 2665 58410 2670
rect 58480 2700 58520 2705
rect 58480 2670 58485 2700
rect 58515 2670 58520 2700
rect 58480 2665 58520 2670
rect 58590 2700 58630 2705
rect 58590 2670 58595 2700
rect 58625 2670 58630 2700
rect 58590 2665 58630 2670
rect 58700 2700 58740 2705
rect 58700 2670 58705 2700
rect 58735 2670 58740 2700
rect 58700 2665 58740 2670
rect 58810 2700 58850 2705
rect 58810 2670 58815 2700
rect 58845 2670 58850 2700
rect 59105 2690 59110 2710
rect 59130 2690 59165 2710
rect 59185 2690 59220 2710
rect 59240 2690 59246 2710
rect 59105 2680 59246 2690
rect 58810 2665 58850 2670
rect 59165 2645 59185 2680
rect 58450 2640 58490 2645
rect 58450 2610 58455 2640
rect 58485 2610 58490 2640
rect 58450 2605 58490 2610
rect 59155 2640 59195 2645
rect 59155 2610 59160 2640
rect 59190 2610 59195 2640
rect 59155 2605 59195 2610
rect 58315 2595 58355 2600
rect 58315 2565 58320 2595
rect 58350 2565 58355 2595
rect 58315 2560 58355 2565
rect 59465 2595 59505 2600
rect 59465 2565 59470 2595
rect 59500 2565 59505 2595
rect 59465 2560 59505 2565
rect 58150 2545 58190 2550
rect 58150 2515 58155 2545
rect 58185 2515 58190 2545
rect 58150 2510 58190 2515
rect 58810 2545 58850 2550
rect 58810 2515 58815 2545
rect 58845 2515 58850 2545
rect 58810 2510 58850 2515
rect 58155 2465 58185 2510
rect 58205 2500 58245 2505
rect 58205 2470 58210 2500
rect 58240 2470 58245 2500
rect 58205 2465 58245 2470
rect 58315 2500 58355 2505
rect 58315 2470 58320 2500
rect 58350 2470 58355 2500
rect 58315 2465 58355 2470
rect 58425 2500 58465 2505
rect 58425 2470 58430 2500
rect 58460 2470 58465 2500
rect 58425 2465 58465 2470
rect 58535 2500 58575 2505
rect 58535 2470 58540 2500
rect 58570 2470 58575 2500
rect 58535 2465 58575 2470
rect 58645 2500 58685 2505
rect 58645 2470 58650 2500
rect 58680 2470 58685 2500
rect 58645 2465 58685 2470
rect 58755 2500 58795 2505
rect 58755 2470 58760 2500
rect 58790 2470 58795 2500
rect 58755 2465 58795 2470
rect 58815 2465 58845 2510
rect 58155 2445 58160 2465
rect 58180 2445 58185 2465
rect 58155 2405 58185 2445
rect 58155 2235 58160 2405
rect 58180 2235 58185 2405
rect 58155 2115 58185 2235
rect 58210 2405 58240 2465
rect 58260 2455 58300 2460
rect 58260 2425 58265 2455
rect 58295 2425 58300 2455
rect 58260 2420 58300 2425
rect 58210 2235 58215 2405
rect 58235 2235 58240 2405
rect 58210 2160 58240 2235
rect 58265 2405 58295 2420
rect 58265 2235 58270 2405
rect 58290 2235 58295 2405
rect 58265 2205 58295 2235
rect 58320 2405 58350 2465
rect 58370 2455 58410 2460
rect 58370 2425 58375 2455
rect 58405 2425 58410 2455
rect 58370 2420 58410 2425
rect 58320 2235 58325 2405
rect 58345 2235 58350 2405
rect 58260 2200 58300 2205
rect 58260 2170 58265 2200
rect 58295 2170 58300 2200
rect 58260 2165 58300 2170
rect 58320 2160 58350 2235
rect 58375 2405 58405 2420
rect 58375 2235 58380 2405
rect 58400 2235 58405 2405
rect 58375 2205 58405 2235
rect 58430 2405 58460 2465
rect 58480 2455 58520 2460
rect 58480 2425 58485 2455
rect 58515 2425 58520 2455
rect 58480 2420 58520 2425
rect 58430 2235 58435 2405
rect 58455 2235 58460 2405
rect 58370 2200 58410 2205
rect 58370 2170 58375 2200
rect 58405 2170 58410 2200
rect 58370 2165 58410 2170
rect 58430 2160 58460 2235
rect 58485 2405 58515 2420
rect 58485 2235 58490 2405
rect 58510 2235 58515 2405
rect 58485 2205 58515 2235
rect 58540 2405 58570 2465
rect 58590 2455 58630 2460
rect 58590 2425 58595 2455
rect 58625 2425 58630 2455
rect 58590 2420 58630 2425
rect 58540 2235 58545 2405
rect 58565 2235 58570 2405
rect 58480 2200 58520 2205
rect 58480 2170 58485 2200
rect 58515 2170 58520 2200
rect 58480 2165 58520 2170
rect 58540 2160 58570 2235
rect 58595 2405 58625 2420
rect 58595 2235 58600 2405
rect 58620 2235 58625 2405
rect 58595 2205 58625 2235
rect 58650 2405 58680 2465
rect 58700 2455 58740 2460
rect 58700 2425 58705 2455
rect 58735 2425 58740 2455
rect 58700 2420 58740 2425
rect 58650 2235 58655 2405
rect 58675 2235 58680 2405
rect 58590 2200 58630 2205
rect 58590 2170 58595 2200
rect 58625 2170 58630 2200
rect 58590 2165 58630 2170
rect 58650 2160 58680 2235
rect 58705 2405 58735 2420
rect 58705 2235 58710 2405
rect 58730 2235 58735 2405
rect 58705 2205 58735 2235
rect 58760 2405 58790 2465
rect 58760 2235 58765 2405
rect 58785 2235 58790 2405
rect 58700 2200 58740 2205
rect 58700 2170 58705 2200
rect 58735 2170 58740 2200
rect 58700 2165 58740 2170
rect 58760 2160 58790 2235
rect 58815 2445 58820 2465
rect 58840 2445 58845 2465
rect 58815 2405 58845 2445
rect 58815 2235 58820 2405
rect 58840 2235 58845 2405
rect 58205 2155 58245 2160
rect 58205 2125 58210 2155
rect 58240 2125 58245 2155
rect 58205 2120 58245 2125
rect 58315 2155 58355 2160
rect 58315 2125 58320 2155
rect 58350 2125 58355 2155
rect 58315 2120 58355 2125
rect 58425 2155 58465 2160
rect 58425 2125 58430 2155
rect 58460 2125 58465 2155
rect 58425 2120 58465 2125
rect 58535 2155 58575 2160
rect 58535 2125 58540 2155
rect 58570 2125 58575 2155
rect 58535 2120 58575 2125
rect 58645 2155 58685 2160
rect 58645 2125 58650 2155
rect 58680 2125 58685 2155
rect 58645 2120 58685 2125
rect 58755 2155 58795 2160
rect 58755 2125 58760 2155
rect 58790 2125 58795 2155
rect 58755 2120 58795 2125
rect 58815 2115 58845 2235
rect 59000 2200 59040 2205
rect 59000 2170 59005 2200
rect 59035 2170 59040 2200
rect 59000 2165 59040 2170
rect 58150 2110 58190 2115
rect 58150 2080 58155 2110
rect 58185 2080 58190 2110
rect 58150 2075 58190 2080
rect 58810 2110 58850 2115
rect 58810 2080 58815 2110
rect 58845 2080 58850 2110
rect 58810 2075 58850 2080
rect 58050 2050 58090 2055
rect 58050 2020 58055 2050
rect 58085 2020 58090 2050
rect 58050 2015 58090 2020
rect 58450 2050 58490 2055
rect 58450 2020 58455 2050
rect 58485 2020 58490 2050
rect 58450 2015 58490 2020
rect 58150 1985 58190 1990
rect 58150 1955 58155 1985
rect 58185 1955 58190 1985
rect 58150 1950 58190 1955
rect 58810 1985 58850 1990
rect 58810 1955 58815 1985
rect 58845 1955 58850 1985
rect 58810 1950 58850 1955
rect 58155 1845 58185 1950
rect 58205 1940 58245 1945
rect 58205 1910 58210 1940
rect 58240 1910 58245 1940
rect 58205 1905 58245 1910
rect 58315 1940 58355 1945
rect 58315 1910 58320 1940
rect 58350 1910 58355 1940
rect 58315 1905 58355 1910
rect 58425 1940 58465 1945
rect 58425 1910 58430 1940
rect 58460 1910 58465 1940
rect 58425 1905 58465 1910
rect 58535 1940 58575 1945
rect 58535 1910 58540 1940
rect 58570 1910 58575 1940
rect 58535 1905 58575 1910
rect 58645 1940 58685 1945
rect 58645 1910 58650 1940
rect 58680 1910 58685 1940
rect 58645 1905 58685 1910
rect 58755 1940 58795 1945
rect 58755 1910 58760 1940
rect 58790 1910 58795 1940
rect 58755 1905 58795 1910
rect 58155 1575 58160 1845
rect 58180 1575 58185 1845
rect 58155 1535 58185 1575
rect 58155 1515 58160 1535
rect 58180 1515 58185 1535
rect 58210 1845 58240 1905
rect 58260 1895 58300 1900
rect 58260 1865 58265 1895
rect 58295 1865 58300 1895
rect 58260 1860 58300 1865
rect 58210 1575 58215 1845
rect 58235 1575 58240 1845
rect 58210 1515 58240 1575
rect 58265 1845 58295 1860
rect 58265 1575 58270 1845
rect 58290 1575 58295 1845
rect 58265 1560 58295 1575
rect 58320 1845 58350 1905
rect 58370 1895 58410 1900
rect 58370 1865 58375 1895
rect 58405 1865 58410 1895
rect 58370 1860 58410 1865
rect 58320 1575 58325 1845
rect 58345 1575 58350 1845
rect 58260 1555 58300 1560
rect 58260 1525 58265 1555
rect 58295 1525 58300 1555
rect 58260 1520 58300 1525
rect 58320 1515 58350 1575
rect 58375 1845 58405 1860
rect 58375 1575 58380 1845
rect 58400 1575 58405 1845
rect 58375 1560 58405 1575
rect 58430 1845 58460 1905
rect 58480 1895 58520 1900
rect 58480 1865 58485 1895
rect 58515 1865 58520 1895
rect 58480 1860 58520 1865
rect 58430 1575 58435 1845
rect 58455 1575 58460 1845
rect 58370 1555 58410 1560
rect 58370 1525 58375 1555
rect 58405 1525 58410 1555
rect 58370 1520 58410 1525
rect 58430 1515 58460 1575
rect 58485 1845 58515 1860
rect 58485 1575 58490 1845
rect 58510 1575 58515 1845
rect 58485 1560 58515 1575
rect 58540 1845 58570 1905
rect 58590 1895 58630 1900
rect 58590 1865 58595 1895
rect 58625 1865 58630 1895
rect 58590 1860 58630 1865
rect 58540 1575 58545 1845
rect 58565 1575 58570 1845
rect 58480 1555 58520 1560
rect 58480 1525 58485 1555
rect 58515 1525 58520 1555
rect 58480 1520 58520 1525
rect 58540 1515 58570 1575
rect 58595 1845 58625 1860
rect 58595 1575 58600 1845
rect 58620 1575 58625 1845
rect 58595 1560 58625 1575
rect 58650 1845 58680 1905
rect 58700 1895 58740 1900
rect 58700 1865 58705 1895
rect 58735 1865 58740 1895
rect 58700 1860 58740 1865
rect 58650 1575 58655 1845
rect 58675 1575 58680 1845
rect 58590 1555 58630 1560
rect 58590 1525 58595 1555
rect 58625 1525 58630 1555
rect 58590 1520 58630 1525
rect 58650 1515 58680 1575
rect 58705 1845 58735 1860
rect 58705 1575 58710 1845
rect 58730 1575 58735 1845
rect 58705 1560 58735 1575
rect 58760 1845 58790 1905
rect 58760 1575 58765 1845
rect 58785 1575 58790 1845
rect 58700 1555 58740 1560
rect 58700 1525 58705 1555
rect 58735 1525 58740 1555
rect 58700 1520 58740 1525
rect 58760 1515 58790 1575
rect 58815 1845 58845 1950
rect 58955 1895 58995 1900
rect 58955 1865 58960 1895
rect 58990 1865 58995 1895
rect 58955 1860 58995 1865
rect 58815 1575 58820 1845
rect 58840 1575 58845 1845
rect 58815 1535 58845 1575
rect 58965 1545 58985 1860
rect 58815 1515 58820 1535
rect 58840 1515 58845 1535
rect 58005 1510 58045 1515
rect 58005 1480 58010 1510
rect 58040 1480 58045 1510
rect 58005 1475 58045 1480
rect 58155 1470 58185 1515
rect 58205 1510 58245 1515
rect 58205 1480 58210 1510
rect 58240 1480 58245 1510
rect 58205 1475 58245 1480
rect 58315 1510 58355 1515
rect 58315 1480 58320 1510
rect 58350 1480 58355 1510
rect 58315 1475 58355 1480
rect 58425 1510 58465 1515
rect 58425 1480 58430 1510
rect 58460 1480 58465 1510
rect 58425 1475 58465 1480
rect 58535 1510 58575 1515
rect 58535 1480 58540 1510
rect 58570 1480 58575 1510
rect 58535 1475 58575 1480
rect 58645 1510 58685 1515
rect 58645 1480 58650 1510
rect 58680 1480 58685 1510
rect 58645 1475 58685 1480
rect 58755 1510 58795 1515
rect 58755 1480 58760 1510
rect 58790 1480 58795 1510
rect 58755 1475 58795 1480
rect 58815 1470 58845 1515
rect 58955 1540 58995 1545
rect 58955 1510 58960 1540
rect 58990 1510 58995 1540
rect 58955 1505 58995 1510
rect 59010 1490 59030 2165
rect 59475 1920 59495 2560
rect 59515 2500 59555 2505
rect 59515 2470 59520 2500
rect 59550 2470 59555 2500
rect 59515 2465 59555 2470
rect 59460 1910 59510 1920
rect 59460 1880 59470 1910
rect 59500 1880 59510 1910
rect 59460 1870 59510 1880
rect 59135 1545 59170 1550
rect 59135 1505 59170 1510
rect 59195 1545 59230 1550
rect 59195 1505 59230 1510
rect 59255 1545 59290 1550
rect 59255 1505 59290 1510
rect 59315 1545 59350 1551
rect 59315 1505 59350 1510
rect 59200 1490 59220 1505
rect 59000 1485 59040 1490
rect 58150 1465 58190 1470
rect 58150 1435 58155 1465
rect 58185 1435 58190 1465
rect 58150 1430 58190 1435
rect 58810 1465 58850 1470
rect 58810 1435 58815 1465
rect 58845 1435 58850 1465
rect 59000 1455 59005 1485
rect 59035 1455 59040 1485
rect 59000 1450 59040 1455
rect 59190 1485 59230 1490
rect 59190 1455 59195 1485
rect 59225 1455 59230 1485
rect 59190 1450 59230 1455
rect 58810 1430 58850 1435
rect 59320 1425 59340 1505
rect 59310 1420 59350 1425
rect 59310 1390 59315 1420
rect 59345 1390 59350 1420
rect 59310 1385 59350 1390
rect 58430 1325 58470 1330
rect 58430 1295 58435 1325
rect 58465 1295 58470 1325
rect 58430 1290 58470 1295
rect 59035 1325 59075 1330
rect 59035 1295 59040 1325
rect 59070 1295 59075 1325
rect 59035 1290 59075 1295
rect 58180 1250 58220 1255
rect 58180 1220 58185 1250
rect 58215 1220 58220 1250
rect 58180 1215 58220 1220
rect 58380 1250 58420 1255
rect 58380 1220 58385 1250
rect 58415 1220 58420 1250
rect 58440 1225 58460 1290
rect 58580 1250 58620 1255
rect 58380 1215 58420 1220
rect 58435 1215 58465 1225
rect 58580 1220 58585 1250
rect 58615 1220 58620 1250
rect 58580 1215 58620 1220
rect 58780 1250 58820 1255
rect 58780 1220 58785 1250
rect 58815 1220 58820 1250
rect 58780 1215 58820 1220
rect 58185 1155 58215 1215
rect 58280 1205 58320 1210
rect 58280 1175 58285 1205
rect 58315 1175 58320 1205
rect 58280 1170 58320 1175
rect 57960 745 58000 750
rect 57960 715 57965 745
rect 57995 715 58000 745
rect 57960 710 58000 715
rect 58185 485 58190 1155
rect 58210 485 58215 1155
rect 58185 445 58215 485
rect 58285 1155 58315 1170
rect 58285 485 58290 1155
rect 58310 485 58315 1155
rect 58285 470 58315 485
rect 58385 1155 58415 1215
rect 58435 1195 58440 1215
rect 58460 1195 58465 1215
rect 58435 1185 58465 1195
rect 58480 1205 58520 1210
rect 58480 1175 58485 1205
rect 58515 1175 58520 1205
rect 58480 1170 58520 1175
rect 58385 485 58390 1155
rect 58410 485 58415 1155
rect 58185 425 58190 445
rect 58210 425 58215 445
rect 58280 465 58320 470
rect 58280 435 58285 465
rect 58315 435 58320 465
rect 58280 430 58320 435
rect 58185 400 58215 425
rect 58385 400 58415 485
rect 58485 1155 58515 1170
rect 58485 485 58490 1155
rect 58510 485 58515 1155
rect 58485 470 58515 485
rect 58585 1155 58615 1215
rect 58680 1205 58720 1210
rect 58680 1175 58685 1205
rect 58715 1175 58720 1205
rect 58680 1170 58720 1175
rect 58585 485 58590 1155
rect 58610 485 58615 1155
rect 58480 465 58520 470
rect 58480 435 58485 465
rect 58515 435 58520 465
rect 58480 430 58520 435
rect 58585 400 58615 485
rect 58685 1155 58715 1170
rect 58685 485 58690 1155
rect 58710 485 58715 1155
rect 58685 470 58715 485
rect 58785 1155 58815 1215
rect 58970 1205 59010 1210
rect 58970 1175 58975 1205
rect 59005 1175 59010 1205
rect 58970 1170 59010 1175
rect 58980 1155 59000 1170
rect 59045 1155 59065 1290
rect 59475 1210 59495 1870
rect 59465 1205 59505 1210
rect 59465 1175 59470 1205
rect 59500 1175 59505 1205
rect 59465 1170 59505 1175
rect 58785 485 58790 1155
rect 58810 485 58815 1155
rect 58975 1150 59010 1155
rect 58975 1110 59010 1115
rect 59035 1150 59070 1155
rect 59035 1110 59070 1115
rect 58680 465 58720 470
rect 58680 435 58685 465
rect 58715 435 58720 465
rect 58680 430 58720 435
rect 58785 445 58815 485
rect 58785 425 58790 445
rect 58810 425 58815 445
rect 58785 400 58815 425
rect 59525 400 59545 2465
rect 54245 395 54285 400
rect 54245 365 54250 395
rect 54280 365 54285 395
rect 54245 360 54285 365
rect 54985 395 55025 400
rect 54985 365 54990 395
rect 55020 365 55025 395
rect 54985 360 55025 365
rect 55185 395 55225 400
rect 55185 365 55190 395
rect 55220 365 55225 395
rect 55185 360 55225 365
rect 55385 395 55425 400
rect 55385 365 55390 395
rect 55420 365 55425 395
rect 55385 360 55425 365
rect 55585 395 55625 400
rect 55585 365 55590 395
rect 55620 365 55625 395
rect 55585 360 55625 365
rect 55845 395 55885 400
rect 55845 365 55850 395
rect 55880 365 55885 395
rect 55845 360 55885 365
rect 56430 395 56470 400
rect 56430 365 56435 395
rect 56465 365 56470 395
rect 56430 360 56470 365
rect 56760 395 56800 400
rect 56760 365 56765 395
rect 56795 365 56800 395
rect 56760 360 56800 365
rect 56880 395 56920 400
rect 56880 365 56885 395
rect 56915 365 56920 395
rect 56880 360 56920 365
rect 57915 395 57955 400
rect 57915 365 57920 395
rect 57950 365 57955 395
rect 57915 360 57955 365
rect 58180 395 58220 400
rect 58180 365 58185 395
rect 58215 365 58220 395
rect 58180 360 58220 365
rect 58380 395 58420 400
rect 58380 365 58385 395
rect 58415 365 58420 395
rect 58380 360 58420 365
rect 58580 395 58620 400
rect 58580 365 58585 395
rect 58615 365 58620 395
rect 58580 360 58620 365
rect 58780 395 58820 400
rect 58780 365 58785 395
rect 58815 365 58820 395
rect 58780 360 58820 365
rect 59515 395 59555 400
rect 59515 365 59520 395
rect 59550 365 59555 395
rect 59515 360 59555 365
rect 56890 -510 56910 360
rect 56880 -515 56920 -510
rect 56880 -545 56885 -515
rect 56915 -545 56920 -515
rect 56880 -550 56920 -545
<< via1 >>
rect 56885 6155 56915 6185
rect 56210 4785 56240 4815
rect 56090 4755 56120 4760
rect 56090 4735 56095 4755
rect 56095 4735 56115 4755
rect 56115 4735 56120 4755
rect 56090 4730 56120 4735
rect 56680 4785 56710 4815
rect 56210 4730 56240 4760
rect 56270 4755 56300 4760
rect 56270 4735 56275 4755
rect 56275 4735 56295 4755
rect 56295 4735 56300 4755
rect 56270 4730 56300 4735
rect 56560 4585 56590 4590
rect 56560 4565 56565 4585
rect 56565 4565 56585 4585
rect 56585 4565 56590 4585
rect 56560 4560 56590 4565
rect 56620 4560 56650 4590
rect 57090 4785 57120 4815
rect 57560 4785 57590 4815
rect 56885 4730 56915 4760
rect 57030 4755 57060 4760
rect 57030 4735 57035 4755
rect 57035 4735 57055 4755
rect 57055 4735 57060 4755
rect 57030 4730 57060 4735
rect 56740 4585 56770 4590
rect 56740 4565 56745 4585
rect 56745 4565 56765 4585
rect 56765 4565 56770 4585
rect 56740 4560 56770 4565
rect 56885 4560 56915 4590
rect 56210 4325 56240 4355
rect 56680 4325 56710 4355
rect 56155 4305 56185 4310
rect 56155 4285 56160 4305
rect 56160 4285 56180 4305
rect 56180 4285 56185 4305
rect 56155 4280 56185 4285
rect 56630 4305 56660 4310
rect 56630 4285 56635 4305
rect 56635 4285 56655 4305
rect 56655 4285 56660 4305
rect 56630 4280 56660 4285
rect 56830 4280 56860 4310
rect 54930 4170 54960 4200
rect 55050 4170 55080 4200
rect 55170 4170 55200 4200
rect 55290 4170 55320 4200
rect 55410 4170 55440 4200
rect 55530 4170 55560 4200
rect 55650 4170 55680 4200
rect 55760 4170 55790 4200
rect 54990 4045 55020 4075
rect 55110 4045 55140 4075
rect 54990 3655 55020 3685
rect 55230 4045 55260 4075
rect 55110 3655 55140 3685
rect 55350 4045 55380 4075
rect 55230 3655 55260 3685
rect 55470 4045 55500 4075
rect 55350 3655 55380 3685
rect 55590 4045 55620 4075
rect 55470 3655 55500 3685
rect 55590 3655 55620 3685
rect 54930 3610 54960 3640
rect 55050 3610 55080 3640
rect 55170 3610 55200 3640
rect 55290 3610 55320 3640
rect 55410 3610 55440 3640
rect 55530 3610 55560 3640
rect 55650 3610 55680 3640
rect 55715 3610 55745 3640
rect 55320 3535 55350 3540
rect 55320 3515 55325 3535
rect 55325 3515 55345 3535
rect 55345 3515 55350 3535
rect 55320 3510 55350 3515
rect 54955 3450 54985 3480
rect 55065 3450 55095 3480
rect 55175 3450 55205 3480
rect 55285 3450 55315 3480
rect 55395 3450 55425 3480
rect 55505 3450 55535 3480
rect 55615 3450 55645 3480
rect 54610 3370 54640 3400
rect 55010 3355 55040 3385
rect 55120 3355 55150 3385
rect 55010 2715 55040 2745
rect 55230 3355 55260 3385
rect 55120 2715 55150 2745
rect 55340 3355 55370 3385
rect 55230 2715 55260 2745
rect 55450 3355 55480 3385
rect 55340 2715 55370 2745
rect 55560 3355 55590 3385
rect 55450 2715 55480 2745
rect 54955 2670 54985 2700
rect 55065 2670 55095 2700
rect 55175 2670 55205 2700
rect 55285 2670 55315 2700
rect 55395 2670 55425 2700
rect 54610 2610 54640 2640
rect 55315 2635 55345 2640
rect 55315 2615 55320 2635
rect 55320 2615 55340 2635
rect 55340 2615 55345 2635
rect 55315 2610 55345 2615
rect 55560 2715 55590 2745
rect 55505 2670 55535 2700
rect 55615 2670 55645 2700
rect 56010 4110 56040 4140
rect 56130 4110 56160 4140
rect 56250 4110 56280 4140
rect 56370 4110 56400 4140
rect 56490 4110 56520 4140
rect 56610 4110 56640 4140
rect 56730 4110 56760 4140
rect 56070 4045 56100 4075
rect 56010 3655 56040 3685
rect 56190 4045 56220 4075
rect 56130 3655 56160 3685
rect 56310 4045 56340 4075
rect 56250 3655 56280 3685
rect 56430 4045 56460 4075
rect 56370 3655 56400 3685
rect 56550 4045 56580 4075
rect 56490 3655 56520 3685
rect 56670 4045 56700 4075
rect 56610 3655 56640 3685
rect 56730 3655 56760 3685
rect 56070 3610 56100 3640
rect 56190 3610 56220 3640
rect 56310 3610 56340 3640
rect 56430 3610 56460 3640
rect 56550 3610 56580 3640
rect 56670 3610 56700 3640
rect 57150 4730 57180 4760
rect 57210 4755 57240 4760
rect 57210 4735 57215 4755
rect 57215 4735 57235 4755
rect 57235 4735 57240 4755
rect 57210 4730 57240 4735
rect 57500 4755 57530 4760
rect 57500 4735 57505 4755
rect 57505 4735 57525 4755
rect 57525 4735 57530 4755
rect 57500 4730 57530 4735
rect 57560 4730 57590 4760
rect 57680 4755 57710 4760
rect 57680 4735 57685 4755
rect 57685 4735 57705 4755
rect 57705 4735 57710 4755
rect 57680 4730 57710 4735
rect 57090 4325 57120 4355
rect 57560 4325 57590 4355
rect 56940 4225 56970 4255
rect 57576 4295 57606 4300
rect 57576 4275 57581 4295
rect 57581 4275 57601 4295
rect 57601 4275 57606 4295
rect 57576 4270 57606 4275
rect 56885 4170 56915 4200
rect 56400 3580 56430 3585
rect 56400 3560 56405 3580
rect 56405 3560 56425 3580
rect 56425 3560 56430 3580
rect 56400 3555 56430 3560
rect 56840 3555 56870 3585
rect 57140 4215 57170 4245
rect 57620 4215 57650 4245
rect 58010 4170 58040 4200
rect 58125 4170 58155 4200
rect 58245 4170 58275 4200
rect 58365 4170 58395 4200
rect 58485 4170 58515 4200
rect 58605 4170 58635 4200
rect 58725 4170 58755 4200
rect 58845 4170 58875 4200
rect 57040 4110 57070 4140
rect 57160 4110 57190 4140
rect 57280 4110 57310 4140
rect 57400 4110 57430 4140
rect 57520 4110 57550 4140
rect 57640 4110 57670 4140
rect 57760 4110 57790 4140
rect 57100 4045 57130 4075
rect 57040 3655 57070 3685
rect 57220 4045 57250 4075
rect 57160 3655 57190 3685
rect 57340 4045 57370 4075
rect 57280 3655 57310 3685
rect 57460 4045 57490 4075
rect 57400 3655 57430 3685
rect 57580 4045 57610 4075
rect 57520 3655 57550 3685
rect 57700 4045 57730 4075
rect 57640 3655 57670 3685
rect 57760 3655 57790 3685
rect 57100 3610 57130 3640
rect 57220 3610 57250 3640
rect 57340 3610 57370 3640
rect 57460 3610 57490 3640
rect 57580 3610 57610 3640
rect 57700 3610 57730 3640
rect 57370 3580 57400 3585
rect 57370 3560 57375 3580
rect 57375 3560 57395 3580
rect 57395 3560 57400 3580
rect 57370 3555 57400 3560
rect 56930 3510 56960 3540
rect 58185 4045 58215 4075
rect 58305 4045 58335 4075
rect 58185 3655 58215 3685
rect 58425 4045 58455 4075
rect 58305 3655 58335 3685
rect 58545 4045 58575 4075
rect 58425 3655 58455 3685
rect 58665 4045 58695 4075
rect 58545 3655 58575 3685
rect 58785 4045 58815 4075
rect 58665 3655 58695 3685
rect 58785 3655 58815 3685
rect 58055 3610 58085 3640
rect 58125 3610 58155 3640
rect 58245 3610 58275 3640
rect 58365 3610 58395 3640
rect 58485 3610 58515 3640
rect 58605 3610 58635 3640
rect 58725 3610 58755 3640
rect 58845 3610 58875 3640
rect 55760 3450 55790 3480
rect 56280 3450 56310 3480
rect 56390 3450 56420 3480
rect 56500 3450 56530 3480
rect 56610 3450 56640 3480
rect 56720 3450 56750 3480
rect 56830 3450 56860 3480
rect 56940 3450 56970 3480
rect 57050 3450 57080 3480
rect 57160 3450 57190 3480
rect 57270 3450 57300 3480
rect 57380 3450 57410 3480
rect 57490 3450 57520 3480
rect 58010 3450 58040 3480
rect 56335 3405 56365 3435
rect 56445 3360 56475 3390
rect 56335 3270 56365 3300
rect 56145 3225 56175 3255
rect 56035 3090 56065 3120
rect 55940 3040 55970 3070
rect 55990 3065 56020 3070
rect 55990 3045 55995 3065
rect 55995 3045 56015 3065
rect 56015 3045 56020 3065
rect 55990 3040 56020 3045
rect 55760 2765 55790 2795
rect 55715 2610 55745 2640
rect 54300 2565 54330 2595
rect 55450 2565 55480 2595
rect 54250 2470 54280 2500
rect 54955 2515 54985 2545
rect 55615 2515 55645 2545
rect 55010 2470 55040 2500
rect 55120 2470 55150 2500
rect 55230 2470 55260 2500
rect 55340 2470 55370 2500
rect 55450 2470 55480 2500
rect 55560 2470 55590 2500
rect 54765 2170 54795 2200
rect 54300 1880 54330 1910
rect 54450 1540 54485 1545
rect 54450 1515 54455 1540
rect 54455 1515 54480 1540
rect 54480 1515 54485 1540
rect 54450 1510 54485 1515
rect 54510 1540 54545 1545
rect 54510 1515 54515 1540
rect 54515 1515 54540 1540
rect 54540 1515 54545 1540
rect 54510 1510 54545 1515
rect 54570 1540 54605 1545
rect 54570 1515 54575 1540
rect 54575 1515 54600 1540
rect 54600 1515 54605 1540
rect 54570 1510 54605 1515
rect 54630 1540 54665 1545
rect 54630 1515 54635 1540
rect 54635 1515 54660 1540
rect 54660 1515 54665 1540
rect 54630 1510 54665 1515
rect 55065 2425 55095 2455
rect 55175 2425 55205 2455
rect 55065 2195 55095 2200
rect 55065 2175 55070 2195
rect 55070 2175 55090 2195
rect 55090 2175 55095 2195
rect 55065 2170 55095 2175
rect 55285 2425 55315 2455
rect 55175 2195 55205 2200
rect 55175 2175 55180 2195
rect 55180 2175 55200 2195
rect 55200 2175 55205 2195
rect 55175 2170 55205 2175
rect 55395 2425 55425 2455
rect 55285 2195 55315 2200
rect 55285 2175 55290 2195
rect 55290 2175 55310 2195
rect 55310 2175 55315 2195
rect 55285 2170 55315 2175
rect 55505 2425 55535 2455
rect 55395 2195 55425 2200
rect 55395 2175 55400 2195
rect 55400 2175 55420 2195
rect 55420 2175 55425 2195
rect 55395 2170 55425 2175
rect 55505 2195 55535 2200
rect 55505 2175 55510 2195
rect 55510 2175 55530 2195
rect 55530 2175 55535 2195
rect 55505 2170 55535 2175
rect 55010 2125 55040 2155
rect 55120 2125 55150 2155
rect 55230 2125 55260 2155
rect 55340 2125 55370 2155
rect 55450 2125 55480 2155
rect 55560 2125 55590 2155
rect 54955 2080 54985 2110
rect 55615 2080 55645 2110
rect 55760 2515 55790 2545
rect 55315 2045 55345 2050
rect 55315 2025 55320 2045
rect 55320 2025 55340 2045
rect 55340 2025 55345 2045
rect 55315 2020 55345 2025
rect 55715 2020 55745 2050
rect 54955 1955 54985 1985
rect 55615 1955 55645 1985
rect 54810 1865 54840 1895
rect 55010 1910 55040 1940
rect 55120 1910 55150 1940
rect 55230 1910 55260 1940
rect 55340 1910 55370 1940
rect 55450 1910 55480 1940
rect 55560 1910 55590 1940
rect 54810 1510 54840 1540
rect 55065 1865 55095 1895
rect 55175 1865 55205 1895
rect 55065 1525 55095 1555
rect 55285 1865 55315 1895
rect 55175 1525 55205 1555
rect 55395 1865 55425 1895
rect 55285 1525 55315 1555
rect 55505 1865 55535 1895
rect 55395 1525 55425 1555
rect 55505 1525 55535 1555
rect 55850 1905 55880 1935
rect 54575 1455 54605 1485
rect 54765 1455 54795 1485
rect 55010 1480 55040 1510
rect 55120 1480 55150 1510
rect 55230 1480 55260 1510
rect 55340 1480 55370 1510
rect 55450 1480 55480 1510
rect 55560 1480 55590 1510
rect 55760 1480 55790 1510
rect 54955 1435 54985 1465
rect 55615 1435 55645 1465
rect 55850 1435 55880 1465
rect 54455 1390 54485 1420
rect 54735 1295 54765 1325
rect 55340 1295 55370 1325
rect 54300 1175 54330 1205
rect 54990 1220 55020 1250
rect 55190 1220 55220 1250
rect 55390 1220 55420 1250
rect 55590 1220 55620 1250
rect 54800 1175 54830 1205
rect 55090 1175 55120 1205
rect 54735 1145 54770 1150
rect 54735 1120 54740 1145
rect 54740 1120 54765 1145
rect 54765 1120 54770 1145
rect 54735 1115 54770 1120
rect 54795 1145 54830 1150
rect 54795 1120 54800 1145
rect 54800 1120 54825 1145
rect 54825 1120 54830 1145
rect 54795 1115 54830 1120
rect 55290 1175 55320 1205
rect 55090 435 55120 465
rect 55490 1175 55520 1205
rect 55290 435 55320 465
rect 56555 3405 56585 3435
rect 56445 3225 56475 3255
rect 56665 3360 56695 3390
rect 56555 3270 56585 3300
rect 56775 3405 56805 3435
rect 56665 3225 56695 3255
rect 56885 3360 56915 3390
rect 56775 3270 56805 3300
rect 56995 3405 57025 3435
rect 56885 3225 56915 3255
rect 57105 3360 57135 3390
rect 56995 3270 57025 3300
rect 57215 3405 57245 3435
rect 57105 3225 57135 3255
rect 57325 3360 57355 3390
rect 57215 3270 57245 3300
rect 57435 3405 57465 3435
rect 57325 3225 57355 3255
rect 57435 3270 57465 3300
rect 57625 3275 57655 3305
rect 56280 3180 56310 3210
rect 56390 3180 56420 3210
rect 56500 3180 56530 3210
rect 56610 3180 56640 3210
rect 56720 3180 56750 3210
rect 56830 3180 56860 3210
rect 56940 3180 56970 3210
rect 57050 3180 57080 3210
rect 57160 3180 57190 3210
rect 57270 3180 57300 3210
rect 57380 3180 57410 3210
rect 57490 3180 57520 3210
rect 56695 3090 56725 3120
rect 56145 3045 56175 3075
rect 56255 3045 56285 3075
rect 56365 3045 56395 3075
rect 56475 3045 56505 3075
rect 56585 3045 56615 3075
rect 56090 3000 56120 3030
rect 56200 3000 56230 3030
rect 56145 2910 56175 2940
rect 56310 3000 56340 3030
rect 56255 2910 56285 2940
rect 56420 3000 56450 3030
rect 56365 2910 56395 2940
rect 56530 3000 56560 3030
rect 56475 2910 56505 2940
rect 56640 3000 56670 3030
rect 56585 2910 56615 2940
rect 56740 3065 56770 3070
rect 56740 3045 56745 3065
rect 56745 3045 56765 3065
rect 56765 3045 56770 3065
rect 56740 3040 56770 3045
rect 57075 3090 57105 3120
rect 57030 3065 57060 3070
rect 57030 3045 57035 3065
rect 57035 3045 57055 3065
rect 57055 3045 57060 3065
rect 57030 3040 57060 3045
rect 57735 3090 57765 3120
rect 57185 3045 57215 3075
rect 57295 3045 57325 3075
rect 57405 3045 57435 3075
rect 57515 3045 57545 3075
rect 57625 3045 57655 3075
rect 57130 3000 57160 3030
rect 57185 2910 57215 2940
rect 56090 2865 56120 2895
rect 56200 2865 56230 2895
rect 56310 2865 56340 2895
rect 56420 2865 56450 2895
rect 56530 2865 56560 2895
rect 56640 2865 56670 2895
rect 56095 2835 56125 2840
rect 56095 2815 56100 2835
rect 56100 2815 56120 2835
rect 56120 2815 56125 2835
rect 56095 2810 56125 2815
rect 56580 2835 56610 2840
rect 56580 2815 56585 2835
rect 56585 2815 56605 2835
rect 56605 2815 56610 2835
rect 56580 2810 56610 2815
rect 56800 2865 56830 2895
rect 57130 2865 57160 2895
rect 57190 2835 57220 2840
rect 57190 2815 57195 2835
rect 57195 2815 57215 2835
rect 57215 2815 57220 2835
rect 57190 2810 57220 2815
rect 56035 2765 56065 2795
rect 56695 2765 56725 2795
rect 57075 2765 57105 2795
rect 57350 3000 57380 3030
rect 57295 2910 57325 2940
rect 57405 2910 57435 2940
rect 57350 2865 57380 2895
rect 56610 2705 56640 2735
rect 56830 2705 56860 2735
rect 57050 2705 57080 2735
rect 57240 2705 57270 2735
rect 56555 2650 56585 2680
rect 56310 2610 56340 2640
rect 56035 2285 56065 2315
rect 56145 2230 56175 2260
rect 56255 2230 56285 2260
rect 56090 2185 56120 2215
rect 56200 2185 56230 2215
rect 56145 1995 56175 2025
rect 56665 2650 56695 2680
rect 56775 2650 56805 2680
rect 56555 2510 56585 2515
rect 56555 2490 56560 2510
rect 56560 2490 56580 2510
rect 56580 2490 56585 2510
rect 56555 2485 56585 2490
rect 56720 2630 56750 2635
rect 56720 2610 56725 2630
rect 56725 2610 56745 2630
rect 56745 2610 56750 2630
rect 56720 2605 56750 2610
rect 56665 2485 56695 2515
rect 56610 2430 56640 2460
rect 56885 2650 56915 2680
rect 56995 2650 57025 2680
rect 56775 2485 56805 2515
rect 56940 2630 56970 2635
rect 56940 2610 56945 2630
rect 56945 2610 56965 2630
rect 56965 2610 56970 2630
rect 56940 2605 56970 2610
rect 56885 2485 56915 2515
rect 56830 2430 56860 2460
rect 57105 2650 57135 2680
rect 57215 2650 57245 2680
rect 56995 2485 57025 2515
rect 57160 2605 57190 2635
rect 57105 2485 57135 2515
rect 57050 2430 57080 2460
rect 57570 3000 57600 3030
rect 57515 2910 57545 2940
rect 57625 2910 57655 2940
rect 57570 2865 57600 2895
rect 57780 3065 57810 3070
rect 57780 3045 57785 3065
rect 57785 3045 57805 3065
rect 57805 3045 57810 3065
rect 57780 3040 57810 3045
rect 57830 3040 57860 3070
rect 57735 2765 57765 2795
rect 57460 2705 57490 2735
rect 57680 2705 57710 2735
rect 57350 2605 57380 2635
rect 57460 2610 57490 2640
rect 57215 2510 57245 2515
rect 57215 2490 57220 2510
rect 57220 2490 57240 2510
rect 57240 2490 57245 2510
rect 57215 2485 57245 2490
rect 56720 2385 56750 2415
rect 56940 2385 56970 2415
rect 57160 2385 57190 2415
rect 56695 2285 56725 2315
rect 57075 2285 57105 2315
rect 56635 2265 56665 2270
rect 56365 2230 56395 2260
rect 56475 2230 56505 2260
rect 56585 2230 56615 2260
rect 56635 2245 56640 2265
rect 56640 2245 56660 2265
rect 56660 2245 56665 2265
rect 56635 2240 56665 2245
rect 56310 2185 56340 2215
rect 56255 1995 56285 2025
rect 56420 2185 56450 2215
rect 56365 1995 56395 2025
rect 56090 1950 56120 1980
rect 56200 1950 56230 1980
rect 56310 1950 56340 1980
rect 56035 1905 56065 1935
rect 56035 1820 56065 1850
rect 55990 1780 56020 1785
rect 55990 1760 55995 1780
rect 55995 1760 56015 1780
rect 56015 1760 56020 1780
rect 55990 1755 56020 1760
rect 56530 2185 56560 2215
rect 56475 1995 56505 2025
rect 56640 2185 56670 2215
rect 56585 1995 56615 2025
rect 57135 2265 57165 2270
rect 57135 2245 57140 2265
rect 57140 2245 57160 2265
rect 57160 2245 57165 2265
rect 57135 2240 57165 2245
rect 57185 2230 57215 2260
rect 57295 2230 57325 2260
rect 57405 2230 57435 2260
rect 57130 2185 57160 2215
rect 56420 1950 56450 1980
rect 56530 1950 56560 1980
rect 56640 1950 56670 1980
rect 57240 2185 57270 2215
rect 57185 1995 57215 2025
rect 57350 2185 57380 2215
rect 57295 1995 57325 2025
rect 57735 2285 57765 2315
rect 57515 2230 57545 2260
rect 57625 2230 57655 2260
rect 57460 2185 57490 2215
rect 57405 1995 57435 2025
rect 57130 1950 57160 1980
rect 57240 1950 57270 1980
rect 57350 1950 57380 1980
rect 56695 1905 56725 1935
rect 57075 1905 57105 1935
rect 56735 1820 56765 1850
rect 56090 1765 56120 1795
rect 56200 1765 56230 1795
rect 56310 1765 56340 1795
rect 56365 1775 56395 1805
rect 56420 1765 56450 1795
rect 56530 1765 56560 1795
rect 56640 1765 56670 1795
rect 56690 1780 56720 1785
rect 56690 1760 56695 1780
rect 56695 1760 56715 1780
rect 56715 1760 56720 1780
rect 56145 1720 56175 1750
rect 56090 1525 56120 1555
rect 56255 1720 56285 1750
rect 56200 1525 56230 1555
rect 56365 1720 56395 1750
rect 56310 1525 56340 1555
rect 56475 1720 56505 1750
rect 56420 1525 56450 1555
rect 56585 1720 56615 1750
rect 56530 1525 56560 1555
rect 56690 1755 56720 1760
rect 56820 1810 56850 1840
rect 56950 1810 56980 1840
rect 57035 1820 57065 1850
rect 56859 1780 56889 1785
rect 56859 1760 56864 1780
rect 56864 1760 56884 1780
rect 56884 1760 56889 1780
rect 56859 1755 56889 1760
rect 56914 1780 56941 1785
rect 56914 1760 56916 1780
rect 56916 1760 56936 1780
rect 56936 1760 56941 1780
rect 56914 1755 56941 1760
rect 57570 2185 57600 2215
rect 57515 1995 57545 2025
rect 57680 2185 57710 2215
rect 57625 1995 57655 2025
rect 57785 2240 57815 2245
rect 57785 2220 57790 2240
rect 57790 2220 57810 2240
rect 57810 2220 57815 2240
rect 57785 2215 57815 2220
rect 57460 1950 57490 1980
rect 57570 1950 57600 1980
rect 57680 1950 57710 1980
rect 57735 1905 57765 1935
rect 57735 1820 57765 1850
rect 57080 1780 57110 1785
rect 57080 1760 57085 1780
rect 57085 1760 57105 1780
rect 57105 1760 57110 1780
rect 57130 1765 57160 1795
rect 57240 1765 57270 1795
rect 57350 1765 57380 1795
rect 57405 1775 57435 1805
rect 57460 1765 57490 1795
rect 57570 1765 57600 1795
rect 57680 1765 57710 1795
rect 57080 1755 57110 1760
rect 57185 1720 57215 1750
rect 56640 1525 56670 1555
rect 56145 1480 56175 1510
rect 56255 1480 56285 1510
rect 56365 1480 56395 1510
rect 56475 1480 56505 1510
rect 56585 1480 56615 1510
rect 56035 1435 56065 1465
rect 56735 1435 56765 1465
rect 55940 1390 55970 1420
rect 56830 1390 56860 1420
rect 56335 1235 56365 1265
rect 57130 1525 57160 1555
rect 57295 1720 57325 1750
rect 57240 1525 57270 1555
rect 57405 1720 57435 1750
rect 57350 1525 57380 1555
rect 57515 1720 57545 1750
rect 57460 1525 57490 1555
rect 57625 1720 57655 1750
rect 57570 1525 57600 1555
rect 57780 1780 57810 1785
rect 57780 1760 57785 1780
rect 57785 1760 57805 1780
rect 57805 1760 57810 1780
rect 57780 1755 57810 1760
rect 57680 1525 57710 1555
rect 57185 1480 57215 1510
rect 57295 1480 57325 1510
rect 57405 1480 57435 1510
rect 57515 1480 57545 1510
rect 57625 1480 57655 1510
rect 57035 1435 57065 1465
rect 56940 1390 56970 1420
rect 56885 1235 56915 1265
rect 57735 1435 57765 1465
rect 58010 2765 58040 2795
rect 58455 3535 58485 3540
rect 58455 3515 58460 3535
rect 58460 3515 58480 3535
rect 58480 3515 58485 3535
rect 58455 3510 58485 3515
rect 58155 3450 58185 3480
rect 58265 3450 58295 3480
rect 58375 3450 58405 3480
rect 58485 3450 58515 3480
rect 58595 3450 58625 3480
rect 58705 3450 58735 3480
rect 58815 3450 58845 3480
rect 58210 3355 58240 3385
rect 58320 3355 58350 3385
rect 58210 2715 58240 2745
rect 58430 3355 58460 3385
rect 58320 2715 58350 2745
rect 58155 2670 58185 2700
rect 58265 2670 58295 2700
rect 58055 2610 58085 2640
rect 57920 2485 57950 2515
rect 58010 2515 58040 2545
rect 57875 2430 57905 2460
rect 57830 1390 57860 1420
rect 57965 2215 57995 2245
rect 57920 1905 57950 1935
rect 57920 1435 57950 1465
rect 57410 1260 57440 1265
rect 57410 1240 57415 1260
rect 57415 1240 57435 1260
rect 57435 1240 57440 1260
rect 57410 1235 57440 1240
rect 57875 1235 57905 1265
rect 56445 1180 56475 1210
rect 56555 1180 56585 1210
rect 56665 1180 56695 1210
rect 56775 1180 56805 1210
rect 56885 1180 56915 1210
rect 56995 1180 57025 1210
rect 57105 1180 57135 1210
rect 57215 1180 57245 1210
rect 57325 1180 57355 1210
rect 57435 1180 57465 1210
rect 55850 860 55880 890
rect 56225 885 56255 890
rect 56225 865 56230 885
rect 56230 865 56250 885
rect 56250 865 56255 885
rect 56225 860 56255 865
rect 56280 860 56310 890
rect 56390 860 56420 890
rect 55490 435 55520 465
rect 56500 860 56530 890
rect 56610 860 56640 890
rect 56720 860 56750 890
rect 56830 860 56860 890
rect 56940 860 56970 890
rect 57050 860 57080 890
rect 57160 860 57190 890
rect 57270 860 57300 890
rect 57380 860 57410 890
rect 57490 885 57520 890
rect 57490 865 57495 885
rect 57495 865 57515 885
rect 57515 865 57520 885
rect 57490 860 57520 865
rect 57920 850 57950 880
rect 56445 815 56475 845
rect 56555 815 56585 845
rect 56665 815 56695 845
rect 56775 815 56805 845
rect 56885 815 56915 845
rect 56995 815 57025 845
rect 57105 815 57135 845
rect 57215 815 57245 845
rect 57325 815 57355 845
rect 57435 815 57465 845
rect 56545 760 56575 790
rect 56655 760 56685 790
rect 56875 760 56905 790
rect 56490 715 56520 745
rect 56600 740 56630 745
rect 56600 720 56605 740
rect 56605 720 56625 740
rect 56625 720 56630 740
rect 56600 715 56630 720
rect 56545 510 56575 540
rect 56710 715 56740 745
rect 56655 510 56685 540
rect 57045 740 57075 745
rect 57045 720 57050 740
rect 57050 720 57070 740
rect 57070 720 57075 740
rect 57045 715 57075 720
rect 56875 510 56905 540
rect 56490 465 56520 495
rect 56600 465 56630 495
rect 56710 465 56740 495
rect 58540 3355 58570 3385
rect 58430 2715 58460 2745
rect 58650 3355 58680 3385
rect 58540 2715 58570 2745
rect 58760 3355 58790 3385
rect 58650 2715 58680 2745
rect 59160 3370 59190 3400
rect 58760 2715 58790 2745
rect 58375 2670 58405 2700
rect 58485 2670 58515 2700
rect 58595 2670 58625 2700
rect 58705 2670 58735 2700
rect 58815 2670 58845 2700
rect 58455 2635 58485 2640
rect 58455 2615 58460 2635
rect 58460 2615 58480 2635
rect 58480 2615 58485 2635
rect 58455 2610 58485 2615
rect 59160 2610 59190 2640
rect 58320 2565 58350 2595
rect 59470 2565 59500 2595
rect 58155 2515 58185 2545
rect 58815 2515 58845 2545
rect 58210 2470 58240 2500
rect 58320 2470 58350 2500
rect 58430 2470 58460 2500
rect 58540 2470 58570 2500
rect 58650 2470 58680 2500
rect 58760 2470 58790 2500
rect 58265 2425 58295 2455
rect 58375 2425 58405 2455
rect 58265 2195 58295 2200
rect 58265 2175 58270 2195
rect 58270 2175 58290 2195
rect 58290 2175 58295 2195
rect 58265 2170 58295 2175
rect 58485 2425 58515 2455
rect 58375 2195 58405 2200
rect 58375 2175 58380 2195
rect 58380 2175 58400 2195
rect 58400 2175 58405 2195
rect 58375 2170 58405 2175
rect 58595 2425 58625 2455
rect 58485 2195 58515 2200
rect 58485 2175 58490 2195
rect 58490 2175 58510 2195
rect 58510 2175 58515 2195
rect 58485 2170 58515 2175
rect 58705 2425 58735 2455
rect 58595 2195 58625 2200
rect 58595 2175 58600 2195
rect 58600 2175 58620 2195
rect 58620 2175 58625 2195
rect 58595 2170 58625 2175
rect 58705 2195 58735 2200
rect 58705 2175 58710 2195
rect 58710 2175 58730 2195
rect 58730 2175 58735 2195
rect 58705 2170 58735 2175
rect 58210 2125 58240 2155
rect 58320 2125 58350 2155
rect 58430 2125 58460 2155
rect 58540 2125 58570 2155
rect 58650 2125 58680 2155
rect 58760 2125 58790 2155
rect 59005 2170 59035 2200
rect 58155 2080 58185 2110
rect 58815 2080 58845 2110
rect 58055 2020 58085 2050
rect 58455 2045 58485 2050
rect 58455 2025 58460 2045
rect 58460 2025 58480 2045
rect 58480 2025 58485 2045
rect 58455 2020 58485 2025
rect 58155 1955 58185 1985
rect 58815 1955 58845 1985
rect 58210 1910 58240 1940
rect 58320 1910 58350 1940
rect 58430 1910 58460 1940
rect 58540 1910 58570 1940
rect 58650 1910 58680 1940
rect 58760 1910 58790 1940
rect 58265 1865 58295 1895
rect 58375 1865 58405 1895
rect 58265 1525 58295 1555
rect 58485 1865 58515 1895
rect 58375 1525 58405 1555
rect 58595 1865 58625 1895
rect 58485 1525 58515 1555
rect 58705 1865 58735 1895
rect 58595 1525 58625 1555
rect 58705 1525 58735 1555
rect 58960 1865 58990 1895
rect 58010 1480 58040 1510
rect 58210 1480 58240 1510
rect 58320 1480 58350 1510
rect 58430 1480 58460 1510
rect 58540 1480 58570 1510
rect 58650 1480 58680 1510
rect 58760 1480 58790 1510
rect 58960 1510 58990 1540
rect 59520 2470 59550 2500
rect 59470 1880 59500 1910
rect 59135 1540 59170 1545
rect 59135 1515 59140 1540
rect 59140 1515 59165 1540
rect 59165 1515 59170 1540
rect 59135 1510 59170 1515
rect 59195 1540 59230 1545
rect 59195 1515 59200 1540
rect 59200 1515 59225 1540
rect 59225 1515 59230 1540
rect 59195 1510 59230 1515
rect 59255 1540 59290 1545
rect 59255 1515 59260 1540
rect 59260 1515 59285 1540
rect 59285 1515 59290 1540
rect 59255 1510 59290 1515
rect 59315 1540 59350 1545
rect 59315 1515 59320 1540
rect 59320 1515 59345 1540
rect 59345 1515 59350 1540
rect 59315 1510 59350 1515
rect 58155 1435 58185 1465
rect 58815 1435 58845 1465
rect 59005 1455 59035 1485
rect 59195 1455 59225 1485
rect 59315 1390 59345 1420
rect 58435 1295 58465 1325
rect 59040 1295 59070 1325
rect 58185 1220 58215 1250
rect 58385 1220 58415 1250
rect 58585 1220 58615 1250
rect 58785 1220 58815 1250
rect 58285 1175 58315 1205
rect 57965 715 57995 745
rect 58485 1175 58515 1205
rect 58285 435 58315 465
rect 58685 1175 58715 1205
rect 58485 435 58515 465
rect 58975 1175 59005 1205
rect 59470 1175 59500 1205
rect 58975 1145 59010 1150
rect 58975 1120 58980 1145
rect 58980 1120 59005 1145
rect 59005 1120 59010 1145
rect 58975 1115 59010 1120
rect 59035 1145 59070 1150
rect 59035 1120 59040 1145
rect 59040 1120 59065 1145
rect 59065 1120 59070 1145
rect 59035 1115 59070 1120
rect 58685 435 58715 465
rect 54250 365 54280 395
rect 54990 365 55020 395
rect 55190 365 55220 395
rect 55390 365 55420 395
rect 55590 365 55620 395
rect 55850 365 55880 395
rect 56435 365 56465 395
rect 56765 365 56795 395
rect 56885 365 56915 395
rect 57920 365 57950 395
rect 58185 365 58215 395
rect 58385 365 58415 395
rect 58585 365 58615 395
rect 58785 365 58815 395
rect 59520 365 59550 395
rect 56885 -545 56915 -515
<< metal2 >>
rect 56880 6185 56920 6190
rect 56880 6155 56885 6185
rect 56915 6155 56920 6185
rect 56880 6150 56920 6155
rect 56205 4815 56245 4820
rect 56205 4785 56210 4815
rect 56240 4810 56245 4815
rect 56675 4815 56715 4820
rect 56675 4810 56680 4815
rect 56240 4790 56680 4810
rect 56240 4785 56245 4790
rect 56205 4780 56245 4785
rect 56675 4785 56680 4790
rect 56710 4785 56715 4815
rect 56675 4780 56715 4785
rect 57085 4815 57125 4820
rect 57085 4785 57090 4815
rect 57120 4810 57125 4815
rect 57555 4815 57595 4820
rect 57555 4810 57560 4815
rect 57120 4790 57560 4810
rect 57120 4785 57125 4790
rect 57085 4780 57125 4785
rect 57555 4785 57560 4790
rect 57590 4785 57595 4815
rect 57555 4780 57595 4785
rect 56085 4760 56125 4765
rect 56085 4730 56090 4760
rect 56120 4755 56125 4760
rect 56205 4760 56245 4765
rect 56205 4755 56210 4760
rect 56120 4735 56210 4755
rect 56120 4730 56125 4735
rect 56085 4725 56125 4730
rect 56205 4730 56210 4735
rect 56240 4755 56245 4760
rect 56265 4760 56305 4765
rect 56265 4755 56270 4760
rect 56240 4735 56270 4755
rect 56240 4730 56245 4735
rect 56205 4725 56245 4730
rect 56265 4730 56270 4735
rect 56300 4730 56305 4760
rect 56265 4725 56305 4730
rect 56880 4760 56920 4765
rect 56880 4730 56885 4760
rect 56915 4755 56920 4760
rect 57025 4760 57065 4765
rect 57025 4755 57030 4760
rect 56915 4735 57030 4755
rect 56915 4730 56920 4735
rect 56880 4725 56920 4730
rect 57025 4730 57030 4735
rect 57060 4755 57065 4760
rect 57145 4760 57185 4765
rect 57145 4755 57150 4760
rect 57060 4735 57150 4755
rect 57060 4730 57065 4735
rect 57025 4725 57065 4730
rect 57145 4730 57150 4735
rect 57180 4755 57185 4760
rect 57205 4760 57245 4765
rect 57205 4755 57210 4760
rect 57180 4735 57210 4755
rect 57180 4730 57185 4735
rect 57145 4725 57185 4730
rect 57205 4730 57210 4735
rect 57240 4730 57245 4760
rect 57205 4725 57245 4730
rect 57495 4760 57535 4765
rect 57495 4730 57500 4760
rect 57530 4755 57535 4760
rect 57555 4760 57595 4765
rect 57555 4755 57560 4760
rect 57530 4735 57560 4755
rect 57530 4730 57535 4735
rect 57495 4725 57535 4730
rect 57555 4730 57560 4735
rect 57590 4755 57595 4760
rect 57675 4760 57715 4765
rect 57675 4755 57680 4760
rect 57590 4735 57680 4755
rect 57590 4730 57595 4735
rect 57555 4725 57595 4730
rect 57675 4730 57680 4735
rect 57710 4730 57715 4760
rect 57675 4725 57715 4730
rect 56555 4590 56595 4595
rect 56555 4560 56560 4590
rect 56590 4585 56595 4590
rect 56615 4590 56655 4595
rect 56615 4585 56620 4590
rect 56590 4565 56620 4585
rect 56590 4560 56595 4565
rect 56555 4555 56595 4560
rect 56615 4560 56620 4565
rect 56650 4585 56655 4590
rect 56735 4590 56775 4595
rect 56735 4585 56740 4590
rect 56650 4565 56740 4585
rect 56650 4560 56655 4565
rect 56615 4555 56655 4560
rect 56735 4560 56740 4565
rect 56770 4585 56775 4590
rect 56880 4590 56920 4595
rect 56880 4585 56885 4590
rect 56770 4565 56885 4585
rect 56770 4560 56775 4565
rect 56735 4555 56775 4560
rect 56880 4560 56885 4565
rect 56915 4560 56920 4590
rect 56880 4555 56920 4560
rect 56205 4355 56245 4360
rect 56205 4325 56210 4355
rect 56240 4350 56245 4355
rect 56675 4355 56715 4360
rect 56675 4350 56680 4355
rect 56240 4330 56680 4350
rect 56240 4325 56245 4330
rect 56205 4320 56245 4325
rect 56675 4325 56680 4330
rect 56710 4325 56715 4355
rect 56675 4320 56715 4325
rect 57085 4355 57125 4360
rect 57085 4325 57090 4355
rect 57120 4350 57125 4355
rect 57555 4355 57595 4360
rect 57555 4350 57560 4355
rect 57120 4330 57560 4350
rect 57120 4325 57125 4330
rect 57085 4320 57125 4325
rect 57555 4325 57560 4330
rect 57590 4325 57595 4355
rect 57555 4320 57595 4325
rect 56150 4310 56190 4315
rect 56150 4280 56155 4310
rect 56185 4305 56190 4310
rect 56630 4310 56660 4315
rect 56185 4285 56630 4305
rect 56185 4280 56190 4285
rect 56150 4275 56190 4280
rect 56825 4310 56865 4315
rect 56825 4305 56830 4310
rect 56660 4285 56830 4305
rect 56630 4275 56660 4280
rect 56825 4280 56830 4285
rect 56860 4305 56865 4310
rect 56860 4300 57606 4305
rect 56860 4285 57576 4300
rect 56860 4280 56865 4285
rect 56825 4275 56865 4280
rect 57576 4265 57606 4270
rect 56935 4255 56975 4260
rect 56935 4225 56940 4255
rect 56970 4240 56975 4255
rect 57135 4245 57175 4250
rect 57135 4240 57140 4245
rect 56970 4225 57140 4240
rect 56935 4220 57140 4225
rect 57135 4215 57140 4220
rect 57170 4240 57175 4245
rect 57615 4245 57655 4250
rect 57615 4240 57620 4245
rect 57170 4220 57620 4240
rect 57170 4215 57175 4220
rect 57135 4210 57175 4215
rect 57615 4215 57620 4220
rect 57650 4215 57655 4245
rect 57615 4210 57655 4215
rect 54925 4200 54965 4205
rect 54925 4170 54930 4200
rect 54960 4195 54965 4200
rect 55045 4200 55085 4205
rect 55045 4195 55050 4200
rect 54960 4175 55050 4195
rect 54960 4170 54965 4175
rect 54925 4165 54965 4170
rect 55045 4170 55050 4175
rect 55080 4195 55085 4200
rect 55165 4200 55205 4205
rect 55165 4195 55170 4200
rect 55080 4175 55170 4195
rect 55080 4170 55085 4175
rect 55045 4165 55085 4170
rect 55165 4170 55170 4175
rect 55200 4195 55205 4200
rect 55285 4200 55325 4205
rect 55285 4195 55290 4200
rect 55200 4175 55290 4195
rect 55200 4170 55205 4175
rect 55165 4165 55205 4170
rect 55285 4170 55290 4175
rect 55320 4195 55325 4200
rect 55405 4200 55445 4205
rect 55405 4195 55410 4200
rect 55320 4175 55410 4195
rect 55320 4170 55325 4175
rect 55285 4165 55325 4170
rect 55405 4170 55410 4175
rect 55440 4195 55445 4200
rect 55525 4200 55565 4205
rect 55525 4195 55530 4200
rect 55440 4175 55530 4195
rect 55440 4170 55445 4175
rect 55405 4165 55445 4170
rect 55525 4170 55530 4175
rect 55560 4195 55565 4200
rect 55645 4200 55685 4205
rect 55645 4195 55650 4200
rect 55560 4175 55650 4195
rect 55560 4170 55565 4175
rect 55525 4165 55565 4170
rect 55645 4170 55650 4175
rect 55680 4195 55685 4200
rect 55755 4200 55795 4205
rect 55755 4195 55760 4200
rect 55680 4175 55760 4195
rect 55680 4170 55685 4175
rect 55645 4165 55685 4170
rect 55755 4170 55760 4175
rect 55790 4195 55795 4200
rect 56880 4200 56920 4205
rect 56880 4195 56885 4200
rect 55790 4175 56885 4195
rect 55790 4170 55795 4175
rect 55755 4165 55795 4170
rect 56880 4170 56885 4175
rect 56915 4195 56920 4200
rect 58005 4200 58045 4205
rect 58005 4195 58010 4200
rect 56915 4175 58010 4195
rect 56915 4170 56920 4175
rect 56880 4165 56920 4170
rect 58005 4170 58010 4175
rect 58040 4195 58045 4200
rect 58120 4200 58160 4205
rect 58120 4195 58125 4200
rect 58040 4175 58125 4195
rect 58040 4170 58045 4175
rect 58005 4165 58045 4170
rect 58120 4170 58125 4175
rect 58155 4195 58160 4200
rect 58240 4200 58280 4205
rect 58240 4195 58245 4200
rect 58155 4175 58245 4195
rect 58155 4170 58160 4175
rect 58120 4165 58160 4170
rect 58240 4170 58245 4175
rect 58275 4195 58280 4200
rect 58360 4200 58400 4205
rect 58360 4195 58365 4200
rect 58275 4175 58365 4195
rect 58275 4170 58280 4175
rect 58240 4165 58280 4170
rect 58360 4170 58365 4175
rect 58395 4195 58400 4200
rect 58480 4200 58520 4205
rect 58480 4195 58485 4200
rect 58395 4175 58485 4195
rect 58395 4170 58400 4175
rect 58360 4165 58400 4170
rect 58480 4170 58485 4175
rect 58515 4195 58520 4200
rect 58600 4200 58640 4205
rect 58600 4195 58605 4200
rect 58515 4175 58605 4195
rect 58515 4170 58520 4175
rect 58480 4165 58520 4170
rect 58600 4170 58605 4175
rect 58635 4195 58640 4200
rect 58720 4200 58760 4205
rect 58720 4195 58725 4200
rect 58635 4175 58725 4195
rect 58635 4170 58640 4175
rect 58600 4165 58640 4170
rect 58720 4170 58725 4175
rect 58755 4195 58760 4200
rect 58840 4200 58880 4205
rect 58840 4195 58845 4200
rect 58755 4175 58845 4195
rect 58755 4170 58760 4175
rect 58720 4165 58760 4170
rect 58840 4170 58845 4175
rect 58875 4170 58880 4200
rect 58840 4165 58880 4170
rect 56005 4140 56045 4145
rect 56005 4110 56010 4140
rect 56040 4135 56045 4140
rect 56125 4140 56165 4145
rect 56125 4135 56130 4140
rect 56040 4115 56130 4135
rect 56040 4110 56045 4115
rect 56005 4105 56045 4110
rect 56125 4110 56130 4115
rect 56160 4135 56165 4140
rect 56245 4140 56285 4145
rect 56245 4135 56250 4140
rect 56160 4115 56250 4135
rect 56160 4110 56165 4115
rect 56125 4105 56165 4110
rect 56245 4110 56250 4115
rect 56280 4135 56285 4140
rect 56365 4140 56405 4145
rect 56365 4135 56370 4140
rect 56280 4115 56370 4135
rect 56280 4110 56285 4115
rect 56245 4105 56285 4110
rect 56365 4110 56370 4115
rect 56400 4135 56405 4140
rect 56485 4140 56525 4145
rect 56485 4135 56490 4140
rect 56400 4115 56490 4135
rect 56400 4110 56405 4115
rect 56365 4105 56405 4110
rect 56485 4110 56490 4115
rect 56520 4135 56525 4140
rect 56605 4140 56645 4145
rect 56605 4135 56610 4140
rect 56520 4115 56610 4135
rect 56520 4110 56525 4115
rect 56485 4105 56525 4110
rect 56605 4110 56610 4115
rect 56640 4135 56645 4140
rect 56725 4140 56765 4145
rect 56725 4135 56730 4140
rect 56640 4115 56730 4135
rect 56640 4110 56645 4115
rect 56605 4105 56645 4110
rect 56725 4110 56730 4115
rect 56760 4110 56765 4140
rect 56725 4105 56765 4110
rect 57035 4140 57075 4145
rect 57035 4110 57040 4140
rect 57070 4135 57075 4140
rect 57155 4140 57195 4145
rect 57155 4135 57160 4140
rect 57070 4115 57160 4135
rect 57070 4110 57075 4115
rect 57035 4105 57075 4110
rect 57155 4110 57160 4115
rect 57190 4135 57195 4140
rect 57275 4140 57315 4145
rect 57275 4135 57280 4140
rect 57190 4115 57280 4135
rect 57190 4110 57195 4115
rect 57155 4105 57195 4110
rect 57275 4110 57280 4115
rect 57310 4135 57315 4140
rect 57395 4140 57435 4145
rect 57395 4135 57400 4140
rect 57310 4115 57400 4135
rect 57310 4110 57315 4115
rect 57275 4105 57315 4110
rect 57395 4110 57400 4115
rect 57430 4135 57435 4140
rect 57515 4140 57555 4145
rect 57515 4135 57520 4140
rect 57430 4115 57520 4135
rect 57430 4110 57435 4115
rect 57395 4105 57435 4110
rect 57515 4110 57520 4115
rect 57550 4135 57555 4140
rect 57635 4140 57675 4145
rect 57635 4135 57640 4140
rect 57550 4115 57640 4135
rect 57550 4110 57555 4115
rect 57515 4105 57555 4110
rect 57635 4110 57640 4115
rect 57670 4135 57675 4140
rect 57755 4140 57795 4145
rect 57755 4135 57760 4140
rect 57670 4115 57760 4135
rect 57670 4110 57675 4115
rect 57635 4105 57675 4110
rect 57755 4110 57760 4115
rect 57790 4110 57795 4140
rect 57755 4105 57795 4110
rect 54985 4075 55025 4080
rect 54985 4045 54990 4075
rect 55020 4070 55025 4075
rect 55105 4075 55145 4080
rect 55105 4070 55110 4075
rect 55020 4050 55110 4070
rect 55020 4045 55025 4050
rect 54985 4040 55025 4045
rect 55105 4045 55110 4050
rect 55140 4070 55145 4075
rect 55225 4075 55265 4080
rect 55225 4070 55230 4075
rect 55140 4050 55230 4070
rect 55140 4045 55145 4050
rect 55105 4040 55145 4045
rect 55225 4045 55230 4050
rect 55260 4070 55265 4075
rect 55345 4075 55385 4080
rect 55345 4070 55350 4075
rect 55260 4050 55350 4070
rect 55260 4045 55265 4050
rect 55225 4040 55265 4045
rect 55345 4045 55350 4050
rect 55380 4070 55385 4075
rect 55465 4075 55505 4080
rect 55465 4070 55470 4075
rect 55380 4050 55470 4070
rect 55380 4045 55385 4050
rect 55345 4040 55385 4045
rect 55465 4045 55470 4050
rect 55500 4070 55505 4075
rect 55585 4075 55625 4080
rect 55585 4070 55590 4075
rect 55500 4050 55590 4070
rect 55500 4045 55505 4050
rect 55465 4040 55505 4045
rect 55585 4045 55590 4050
rect 55620 4045 55625 4075
rect 55585 4040 55625 4045
rect 56065 4075 56105 4080
rect 56065 4045 56070 4075
rect 56100 4070 56105 4075
rect 56185 4075 56225 4080
rect 56185 4070 56190 4075
rect 56100 4050 56190 4070
rect 56100 4045 56105 4050
rect 56065 4040 56105 4045
rect 56185 4045 56190 4050
rect 56220 4070 56225 4075
rect 56305 4075 56345 4080
rect 56305 4070 56310 4075
rect 56220 4050 56310 4070
rect 56220 4045 56225 4050
rect 56185 4040 56225 4045
rect 56305 4045 56310 4050
rect 56340 4070 56345 4075
rect 56425 4075 56465 4080
rect 56425 4070 56430 4075
rect 56340 4050 56430 4070
rect 56340 4045 56345 4050
rect 56305 4040 56345 4045
rect 56425 4045 56430 4050
rect 56460 4070 56465 4075
rect 56545 4075 56585 4080
rect 56545 4070 56550 4075
rect 56460 4050 56550 4070
rect 56460 4045 56465 4050
rect 56425 4040 56465 4045
rect 56545 4045 56550 4050
rect 56580 4070 56585 4075
rect 56665 4075 56705 4080
rect 56665 4070 56670 4075
rect 56580 4050 56670 4070
rect 56580 4045 56585 4050
rect 56545 4040 56585 4045
rect 56665 4045 56670 4050
rect 56700 4045 56705 4075
rect 56665 4040 56705 4045
rect 57095 4075 57135 4080
rect 57095 4045 57100 4075
rect 57130 4070 57135 4075
rect 57215 4075 57255 4080
rect 57215 4070 57220 4075
rect 57130 4050 57220 4070
rect 57130 4045 57135 4050
rect 57095 4040 57135 4045
rect 57215 4045 57220 4050
rect 57250 4070 57255 4075
rect 57335 4075 57375 4080
rect 57335 4070 57340 4075
rect 57250 4050 57340 4070
rect 57250 4045 57255 4050
rect 57215 4040 57255 4045
rect 57335 4045 57340 4050
rect 57370 4070 57375 4075
rect 57455 4075 57495 4080
rect 57455 4070 57460 4075
rect 57370 4050 57460 4070
rect 57370 4045 57375 4050
rect 57335 4040 57375 4045
rect 57455 4045 57460 4050
rect 57490 4070 57495 4075
rect 57575 4075 57615 4080
rect 57575 4070 57580 4075
rect 57490 4050 57580 4070
rect 57490 4045 57495 4050
rect 57455 4040 57495 4045
rect 57575 4045 57580 4050
rect 57610 4070 57615 4075
rect 57695 4075 57735 4080
rect 57695 4070 57700 4075
rect 57610 4050 57700 4070
rect 57610 4045 57615 4050
rect 57575 4040 57615 4045
rect 57695 4045 57700 4050
rect 57730 4045 57735 4075
rect 57695 4040 57735 4045
rect 58180 4075 58220 4080
rect 58180 4045 58185 4075
rect 58215 4070 58220 4075
rect 58300 4075 58340 4080
rect 58300 4070 58305 4075
rect 58215 4050 58305 4070
rect 58215 4045 58220 4050
rect 58180 4040 58220 4045
rect 58300 4045 58305 4050
rect 58335 4070 58340 4075
rect 58420 4075 58460 4080
rect 58420 4070 58425 4075
rect 58335 4050 58425 4070
rect 58335 4045 58340 4050
rect 58300 4040 58340 4045
rect 58420 4045 58425 4050
rect 58455 4070 58460 4075
rect 58540 4075 58580 4080
rect 58540 4070 58545 4075
rect 58455 4050 58545 4070
rect 58455 4045 58460 4050
rect 58420 4040 58460 4045
rect 58540 4045 58545 4050
rect 58575 4070 58580 4075
rect 58660 4075 58700 4080
rect 58660 4070 58665 4075
rect 58575 4050 58665 4070
rect 58575 4045 58580 4050
rect 58540 4040 58580 4045
rect 58660 4045 58665 4050
rect 58695 4070 58700 4075
rect 58780 4075 58820 4080
rect 58780 4070 58785 4075
rect 58695 4050 58785 4070
rect 58695 4045 58700 4050
rect 58660 4040 58700 4045
rect 58780 4045 58785 4050
rect 58815 4045 58820 4075
rect 58780 4040 58820 4045
rect 54985 3685 55025 3690
rect 54985 3655 54990 3685
rect 55020 3680 55025 3685
rect 55105 3685 55145 3690
rect 55105 3680 55110 3685
rect 55020 3660 55110 3680
rect 55020 3655 55025 3660
rect 54985 3650 55025 3655
rect 55105 3655 55110 3660
rect 55140 3680 55145 3685
rect 55225 3685 55265 3690
rect 55225 3680 55230 3685
rect 55140 3660 55230 3680
rect 55140 3655 55145 3660
rect 55105 3650 55145 3655
rect 55225 3655 55230 3660
rect 55260 3680 55265 3685
rect 55345 3685 55385 3690
rect 55345 3680 55350 3685
rect 55260 3660 55350 3680
rect 55260 3655 55265 3660
rect 55225 3650 55265 3655
rect 55345 3655 55350 3660
rect 55380 3680 55385 3685
rect 55465 3685 55505 3690
rect 55465 3680 55470 3685
rect 55380 3660 55470 3680
rect 55380 3655 55385 3660
rect 55345 3650 55385 3655
rect 55465 3655 55470 3660
rect 55500 3680 55505 3685
rect 55585 3685 55625 3690
rect 55585 3680 55590 3685
rect 55500 3660 55590 3680
rect 55500 3655 55505 3660
rect 55465 3650 55505 3655
rect 55585 3655 55590 3660
rect 55620 3680 55625 3685
rect 56005 3685 56045 3690
rect 56005 3680 56010 3685
rect 55620 3660 56010 3680
rect 55620 3655 55625 3660
rect 55585 3650 55625 3655
rect 56005 3655 56010 3660
rect 56040 3680 56045 3685
rect 56125 3685 56165 3690
rect 56125 3680 56130 3685
rect 56040 3660 56130 3680
rect 56040 3655 56045 3660
rect 56005 3650 56045 3655
rect 56125 3655 56130 3660
rect 56160 3680 56165 3685
rect 56245 3685 56285 3690
rect 56245 3680 56250 3685
rect 56160 3660 56250 3680
rect 56160 3655 56165 3660
rect 56125 3650 56165 3655
rect 56245 3655 56250 3660
rect 56280 3680 56285 3685
rect 56365 3685 56405 3690
rect 56365 3680 56370 3685
rect 56280 3660 56370 3680
rect 56280 3655 56285 3660
rect 56245 3650 56285 3655
rect 56365 3655 56370 3660
rect 56400 3680 56405 3685
rect 56485 3685 56525 3690
rect 56485 3680 56490 3685
rect 56400 3660 56490 3680
rect 56400 3655 56405 3660
rect 56365 3650 56405 3655
rect 56485 3655 56490 3660
rect 56520 3680 56525 3685
rect 56605 3685 56645 3690
rect 56605 3680 56610 3685
rect 56520 3660 56610 3680
rect 56520 3655 56525 3660
rect 56485 3650 56525 3655
rect 56605 3655 56610 3660
rect 56640 3680 56645 3685
rect 56725 3685 56765 3690
rect 56725 3680 56730 3685
rect 56640 3660 56730 3680
rect 56640 3655 56645 3660
rect 56605 3650 56645 3655
rect 56725 3655 56730 3660
rect 56760 3655 56765 3685
rect 56725 3650 56765 3655
rect 57035 3685 57075 3690
rect 57035 3655 57040 3685
rect 57070 3680 57075 3685
rect 57155 3685 57195 3690
rect 57155 3680 57160 3685
rect 57070 3660 57160 3680
rect 57070 3655 57075 3660
rect 57035 3650 57075 3655
rect 57155 3655 57160 3660
rect 57190 3680 57195 3685
rect 57275 3685 57315 3690
rect 57275 3680 57280 3685
rect 57190 3660 57280 3680
rect 57190 3655 57195 3660
rect 57155 3650 57195 3655
rect 57275 3655 57280 3660
rect 57310 3680 57315 3685
rect 57395 3685 57435 3690
rect 57395 3680 57400 3685
rect 57310 3660 57400 3680
rect 57310 3655 57315 3660
rect 57275 3650 57315 3655
rect 57395 3655 57400 3660
rect 57430 3680 57435 3685
rect 57515 3685 57555 3690
rect 57515 3680 57520 3685
rect 57430 3660 57520 3680
rect 57430 3655 57435 3660
rect 57395 3650 57435 3655
rect 57515 3655 57520 3660
rect 57550 3680 57555 3685
rect 57635 3685 57675 3690
rect 57635 3680 57640 3685
rect 57550 3660 57640 3680
rect 57550 3655 57555 3660
rect 57515 3650 57555 3655
rect 57635 3655 57640 3660
rect 57670 3680 57675 3685
rect 57755 3685 57795 3690
rect 57755 3680 57760 3685
rect 57670 3660 57760 3680
rect 57670 3655 57675 3660
rect 57635 3650 57675 3655
rect 57755 3655 57760 3660
rect 57790 3680 57795 3685
rect 58180 3685 58220 3690
rect 58180 3680 58185 3685
rect 57790 3660 58185 3680
rect 57790 3655 57795 3660
rect 57755 3650 57795 3655
rect 58180 3655 58185 3660
rect 58215 3680 58220 3685
rect 58300 3685 58340 3690
rect 58300 3680 58305 3685
rect 58215 3660 58305 3680
rect 58215 3655 58220 3660
rect 58180 3650 58220 3655
rect 58300 3655 58305 3660
rect 58335 3680 58340 3685
rect 58420 3685 58460 3690
rect 58420 3680 58425 3685
rect 58335 3660 58425 3680
rect 58335 3655 58340 3660
rect 58300 3650 58340 3655
rect 58420 3655 58425 3660
rect 58455 3680 58460 3685
rect 58540 3685 58580 3690
rect 58540 3680 58545 3685
rect 58455 3660 58545 3680
rect 58455 3655 58460 3660
rect 58420 3650 58460 3655
rect 58540 3655 58545 3660
rect 58575 3680 58580 3685
rect 58660 3685 58700 3690
rect 58660 3680 58665 3685
rect 58575 3660 58665 3680
rect 58575 3655 58580 3660
rect 58540 3650 58580 3655
rect 58660 3655 58665 3660
rect 58695 3680 58700 3685
rect 58780 3685 58820 3690
rect 58780 3680 58785 3685
rect 58695 3660 58785 3680
rect 58695 3655 58700 3660
rect 58660 3650 58700 3655
rect 58780 3655 58785 3660
rect 58815 3655 58820 3685
rect 58780 3650 58820 3655
rect 54925 3640 54965 3645
rect 54925 3610 54930 3640
rect 54960 3635 54965 3640
rect 55045 3640 55085 3645
rect 55045 3635 55050 3640
rect 54960 3615 55050 3635
rect 54960 3610 54965 3615
rect 54925 3605 54965 3610
rect 55045 3610 55050 3615
rect 55080 3635 55085 3640
rect 55165 3640 55205 3645
rect 55165 3635 55170 3640
rect 55080 3615 55170 3635
rect 55080 3610 55085 3615
rect 55045 3605 55085 3610
rect 55165 3610 55170 3615
rect 55200 3635 55205 3640
rect 55285 3640 55325 3645
rect 55285 3635 55290 3640
rect 55200 3615 55290 3635
rect 55200 3610 55205 3615
rect 55165 3605 55205 3610
rect 55285 3610 55290 3615
rect 55320 3635 55325 3640
rect 55405 3640 55445 3645
rect 55405 3635 55410 3640
rect 55320 3615 55410 3635
rect 55320 3610 55325 3615
rect 55285 3605 55325 3610
rect 55405 3610 55410 3615
rect 55440 3635 55445 3640
rect 55525 3640 55565 3645
rect 55525 3635 55530 3640
rect 55440 3615 55530 3635
rect 55440 3610 55445 3615
rect 55405 3605 55445 3610
rect 55525 3610 55530 3615
rect 55560 3635 55565 3640
rect 55645 3640 55685 3645
rect 55645 3635 55650 3640
rect 55560 3615 55650 3635
rect 55560 3610 55565 3615
rect 55525 3605 55565 3610
rect 55645 3610 55650 3615
rect 55680 3610 55685 3640
rect 55645 3605 55685 3610
rect 55710 3640 55750 3645
rect 55710 3610 55715 3640
rect 55745 3635 55750 3640
rect 56065 3640 56105 3645
rect 56065 3635 56070 3640
rect 55745 3615 56070 3635
rect 55745 3610 55750 3615
rect 55710 3605 55750 3610
rect 56065 3610 56070 3615
rect 56100 3635 56105 3640
rect 56185 3640 56225 3645
rect 56185 3635 56190 3640
rect 56100 3615 56190 3635
rect 56100 3610 56105 3615
rect 56065 3605 56105 3610
rect 56185 3610 56190 3615
rect 56220 3635 56225 3640
rect 56305 3640 56345 3645
rect 56305 3635 56310 3640
rect 56220 3615 56310 3635
rect 56220 3610 56225 3615
rect 56185 3605 56225 3610
rect 56305 3610 56310 3615
rect 56340 3635 56345 3640
rect 56425 3640 56465 3645
rect 56425 3635 56430 3640
rect 56340 3615 56430 3635
rect 56340 3610 56345 3615
rect 56305 3605 56345 3610
rect 56425 3610 56430 3615
rect 56460 3635 56465 3640
rect 56545 3640 56585 3645
rect 56545 3635 56550 3640
rect 56460 3615 56550 3635
rect 56460 3610 56465 3615
rect 56425 3605 56465 3610
rect 56545 3610 56550 3615
rect 56580 3635 56585 3640
rect 56665 3640 56705 3645
rect 56665 3635 56670 3640
rect 56580 3615 56670 3635
rect 56580 3610 56585 3615
rect 56545 3605 56585 3610
rect 56665 3610 56670 3615
rect 56700 3610 56705 3640
rect 56665 3605 56705 3610
rect 57095 3640 57135 3645
rect 57095 3610 57100 3640
rect 57130 3635 57135 3640
rect 57215 3640 57255 3645
rect 57215 3635 57220 3640
rect 57130 3615 57220 3635
rect 57130 3610 57135 3615
rect 57095 3605 57135 3610
rect 57215 3610 57220 3615
rect 57250 3635 57255 3640
rect 57335 3640 57375 3645
rect 57335 3635 57340 3640
rect 57250 3615 57340 3635
rect 57250 3610 57255 3615
rect 57215 3605 57255 3610
rect 57335 3610 57340 3615
rect 57370 3635 57375 3640
rect 57455 3640 57495 3645
rect 57455 3635 57460 3640
rect 57370 3615 57460 3635
rect 57370 3610 57375 3615
rect 57335 3605 57375 3610
rect 57455 3610 57460 3615
rect 57490 3635 57495 3640
rect 57575 3640 57615 3645
rect 57575 3635 57580 3640
rect 57490 3615 57580 3635
rect 57490 3610 57495 3615
rect 57455 3605 57495 3610
rect 57575 3610 57580 3615
rect 57610 3635 57615 3640
rect 57695 3640 57735 3645
rect 57695 3635 57700 3640
rect 57610 3615 57700 3635
rect 57610 3610 57615 3615
rect 57575 3605 57615 3610
rect 57695 3610 57700 3615
rect 57730 3635 57735 3640
rect 58050 3640 58090 3645
rect 58050 3635 58055 3640
rect 57730 3615 58055 3635
rect 57730 3610 57735 3615
rect 57695 3605 57735 3610
rect 58050 3610 58055 3615
rect 58085 3610 58090 3640
rect 58050 3605 58090 3610
rect 58120 3640 58160 3645
rect 58120 3610 58125 3640
rect 58155 3635 58160 3640
rect 58240 3640 58280 3645
rect 58240 3635 58245 3640
rect 58155 3615 58245 3635
rect 58155 3610 58160 3615
rect 58120 3605 58160 3610
rect 58240 3610 58245 3615
rect 58275 3635 58280 3640
rect 58360 3640 58400 3645
rect 58360 3635 58365 3640
rect 58275 3615 58365 3635
rect 58275 3610 58280 3615
rect 58240 3605 58280 3610
rect 58360 3610 58365 3615
rect 58395 3635 58400 3640
rect 58480 3640 58520 3645
rect 58480 3635 58485 3640
rect 58395 3615 58485 3635
rect 58395 3610 58400 3615
rect 58360 3605 58400 3610
rect 58480 3610 58485 3615
rect 58515 3635 58520 3640
rect 58600 3640 58640 3645
rect 58600 3635 58605 3640
rect 58515 3615 58605 3635
rect 58515 3610 58520 3615
rect 58480 3605 58520 3610
rect 58600 3610 58605 3615
rect 58635 3635 58640 3640
rect 58720 3640 58760 3645
rect 58720 3635 58725 3640
rect 58635 3615 58725 3635
rect 58635 3610 58640 3615
rect 58600 3605 58640 3610
rect 58720 3610 58725 3615
rect 58755 3635 58760 3640
rect 58840 3640 58880 3645
rect 58840 3635 58845 3640
rect 58755 3615 58845 3635
rect 58755 3610 58760 3615
rect 58720 3605 58760 3610
rect 58840 3610 58845 3615
rect 58875 3610 58880 3640
rect 58840 3605 58880 3610
rect 56395 3585 56435 3590
rect 56395 3555 56400 3585
rect 56430 3580 56435 3585
rect 56835 3585 56875 3590
rect 56835 3580 56840 3585
rect 56430 3560 56840 3580
rect 56430 3555 56435 3560
rect 56395 3550 56435 3555
rect 56835 3555 56840 3560
rect 56870 3580 56875 3585
rect 57365 3585 57405 3590
rect 57365 3580 57370 3585
rect 56870 3560 57370 3580
rect 56870 3555 56875 3560
rect 56835 3550 56875 3555
rect 57365 3555 57370 3560
rect 57400 3555 57405 3585
rect 57365 3550 57405 3555
rect 55315 3540 55355 3545
rect 55315 3510 55320 3540
rect 55350 3535 55355 3540
rect 56925 3540 56965 3545
rect 56925 3535 56930 3540
rect 55350 3515 56930 3535
rect 55350 3510 55355 3515
rect 55315 3505 55355 3510
rect 56925 3510 56930 3515
rect 56960 3535 56965 3540
rect 58450 3540 58490 3545
rect 58450 3535 58455 3540
rect 56960 3515 58455 3535
rect 56960 3510 56965 3515
rect 56925 3505 56965 3510
rect 58450 3510 58455 3515
rect 58485 3510 58490 3540
rect 58450 3505 58490 3510
rect 54950 3480 54990 3485
rect 54950 3450 54955 3480
rect 54985 3475 54990 3480
rect 55060 3480 55100 3485
rect 55060 3475 55065 3480
rect 54985 3455 55065 3475
rect 54985 3450 54990 3455
rect 54950 3445 54990 3450
rect 55060 3450 55065 3455
rect 55095 3475 55100 3480
rect 55170 3480 55210 3485
rect 55170 3475 55175 3480
rect 55095 3455 55175 3475
rect 55095 3450 55100 3455
rect 55060 3445 55100 3450
rect 55170 3450 55175 3455
rect 55205 3475 55210 3480
rect 55280 3480 55320 3485
rect 55280 3475 55285 3480
rect 55205 3455 55285 3475
rect 55205 3450 55210 3455
rect 55170 3445 55210 3450
rect 55280 3450 55285 3455
rect 55315 3475 55320 3480
rect 55390 3480 55430 3485
rect 55390 3475 55395 3480
rect 55315 3455 55395 3475
rect 55315 3450 55320 3455
rect 55280 3445 55320 3450
rect 55390 3450 55395 3455
rect 55425 3475 55430 3480
rect 55500 3480 55540 3485
rect 55500 3475 55505 3480
rect 55425 3455 55505 3475
rect 55425 3450 55430 3455
rect 55390 3445 55430 3450
rect 55500 3450 55505 3455
rect 55535 3475 55540 3480
rect 55610 3480 55650 3485
rect 55610 3475 55615 3480
rect 55535 3455 55615 3475
rect 55535 3450 55540 3455
rect 55500 3445 55540 3450
rect 55610 3450 55615 3455
rect 55645 3475 55650 3480
rect 55755 3480 55795 3485
rect 55755 3475 55760 3480
rect 55645 3455 55760 3475
rect 55645 3450 55650 3455
rect 55610 3445 55650 3450
rect 55755 3450 55760 3455
rect 55790 3450 55795 3480
rect 55755 3445 55795 3450
rect 56275 3480 56315 3485
rect 56275 3450 56280 3480
rect 56310 3475 56315 3480
rect 56385 3480 56425 3485
rect 56385 3475 56390 3480
rect 56310 3455 56390 3475
rect 56310 3450 56315 3455
rect 56275 3445 56315 3450
rect 56385 3450 56390 3455
rect 56420 3475 56425 3480
rect 56495 3480 56535 3485
rect 56495 3475 56500 3480
rect 56420 3455 56500 3475
rect 56420 3450 56425 3455
rect 56385 3445 56425 3450
rect 56495 3450 56500 3455
rect 56530 3475 56535 3480
rect 56605 3480 56645 3485
rect 56605 3475 56610 3480
rect 56530 3455 56610 3475
rect 56530 3450 56535 3455
rect 56495 3445 56535 3450
rect 56605 3450 56610 3455
rect 56640 3475 56645 3480
rect 56715 3480 56755 3485
rect 56715 3475 56720 3480
rect 56640 3455 56720 3475
rect 56640 3450 56645 3455
rect 56605 3445 56645 3450
rect 56715 3450 56720 3455
rect 56750 3475 56755 3480
rect 56825 3480 56865 3485
rect 56825 3475 56830 3480
rect 56750 3455 56830 3475
rect 56750 3450 56755 3455
rect 56715 3445 56755 3450
rect 56825 3450 56830 3455
rect 56860 3475 56865 3480
rect 56935 3480 56975 3485
rect 56935 3475 56940 3480
rect 56860 3455 56940 3475
rect 56860 3450 56865 3455
rect 56825 3445 56865 3450
rect 56935 3450 56940 3455
rect 56970 3475 56975 3480
rect 57045 3480 57085 3485
rect 57045 3475 57050 3480
rect 56970 3455 57050 3475
rect 56970 3450 56975 3455
rect 56935 3445 56975 3450
rect 57045 3450 57050 3455
rect 57080 3475 57085 3480
rect 57155 3480 57195 3485
rect 57155 3475 57160 3480
rect 57080 3455 57160 3475
rect 57080 3450 57085 3455
rect 57045 3445 57085 3450
rect 57155 3450 57160 3455
rect 57190 3475 57195 3480
rect 57265 3480 57305 3485
rect 57265 3475 57270 3480
rect 57190 3455 57270 3475
rect 57190 3450 57195 3455
rect 57155 3445 57195 3450
rect 57265 3450 57270 3455
rect 57300 3475 57305 3480
rect 57375 3480 57415 3485
rect 57375 3475 57380 3480
rect 57300 3455 57380 3475
rect 57300 3450 57305 3455
rect 57265 3445 57305 3450
rect 57375 3450 57380 3455
rect 57410 3475 57415 3480
rect 57485 3480 57525 3485
rect 57485 3475 57490 3480
rect 57410 3455 57490 3475
rect 57410 3450 57415 3455
rect 57375 3445 57415 3450
rect 57485 3450 57490 3455
rect 57520 3475 57525 3480
rect 58005 3480 58045 3485
rect 58005 3475 58010 3480
rect 57520 3455 58010 3475
rect 57520 3450 57525 3455
rect 57485 3445 57525 3450
rect 58005 3450 58010 3455
rect 58040 3475 58045 3480
rect 58150 3480 58190 3485
rect 58150 3475 58155 3480
rect 58040 3455 58155 3475
rect 58040 3450 58045 3455
rect 58005 3445 58045 3450
rect 58150 3450 58155 3455
rect 58185 3475 58190 3480
rect 58260 3480 58300 3485
rect 58260 3475 58265 3480
rect 58185 3455 58265 3475
rect 58185 3450 58190 3455
rect 58150 3445 58190 3450
rect 58260 3450 58265 3455
rect 58295 3475 58300 3480
rect 58370 3480 58410 3485
rect 58370 3475 58375 3480
rect 58295 3455 58375 3475
rect 58295 3450 58300 3455
rect 58260 3445 58300 3450
rect 58370 3450 58375 3455
rect 58405 3475 58410 3480
rect 58480 3480 58520 3485
rect 58480 3475 58485 3480
rect 58405 3455 58485 3475
rect 58405 3450 58410 3455
rect 58370 3445 58410 3450
rect 58480 3450 58485 3455
rect 58515 3475 58520 3480
rect 58590 3480 58630 3485
rect 58590 3475 58595 3480
rect 58515 3455 58595 3475
rect 58515 3450 58520 3455
rect 58480 3445 58520 3450
rect 58590 3450 58595 3455
rect 58625 3475 58630 3480
rect 58700 3480 58740 3485
rect 58700 3475 58705 3480
rect 58625 3455 58705 3475
rect 58625 3450 58630 3455
rect 58590 3445 58630 3450
rect 58700 3450 58705 3455
rect 58735 3475 58740 3480
rect 58810 3480 58850 3485
rect 58810 3475 58815 3480
rect 58735 3455 58815 3475
rect 58735 3450 58740 3455
rect 58700 3445 58740 3450
rect 58810 3450 58815 3455
rect 58845 3450 58850 3480
rect 58810 3445 58850 3450
rect 56330 3435 56370 3440
rect 56330 3405 56335 3435
rect 56365 3430 56370 3435
rect 56550 3435 56590 3440
rect 56550 3430 56555 3435
rect 56365 3410 56555 3430
rect 56365 3405 56370 3410
rect 54605 3400 54645 3405
rect 56330 3400 56370 3405
rect 56550 3405 56555 3410
rect 56585 3430 56590 3435
rect 56770 3435 56810 3440
rect 56770 3430 56775 3435
rect 56585 3410 56775 3430
rect 56585 3405 56590 3410
rect 56550 3400 56590 3405
rect 56770 3405 56775 3410
rect 56805 3430 56810 3435
rect 56990 3435 57030 3440
rect 56990 3430 56995 3435
rect 56805 3410 56995 3430
rect 56805 3405 56810 3410
rect 56770 3400 56810 3405
rect 56990 3405 56995 3410
rect 57025 3430 57030 3435
rect 57210 3435 57250 3440
rect 57210 3430 57215 3435
rect 57025 3410 57215 3430
rect 57025 3405 57030 3410
rect 56990 3400 57030 3405
rect 57210 3405 57215 3410
rect 57245 3430 57250 3435
rect 57430 3435 57470 3440
rect 57430 3430 57435 3435
rect 57245 3410 57435 3430
rect 57245 3405 57250 3410
rect 57210 3400 57250 3405
rect 57430 3405 57435 3410
rect 57465 3405 57470 3435
rect 57430 3400 57470 3405
rect 59155 3400 59195 3405
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 56440 3390 56480 3395
rect 54605 3365 54645 3370
rect 55005 3385 55045 3390
rect 55005 3355 55010 3385
rect 55040 3380 55045 3385
rect 55115 3385 55155 3390
rect 55115 3380 55120 3385
rect 55040 3360 55120 3380
rect 55040 3355 55045 3360
rect 55005 3350 55045 3355
rect 55115 3355 55120 3360
rect 55150 3380 55155 3385
rect 55225 3385 55265 3390
rect 55225 3380 55230 3385
rect 55150 3360 55230 3380
rect 55150 3355 55155 3360
rect 55115 3350 55155 3355
rect 55225 3355 55230 3360
rect 55260 3380 55265 3385
rect 55335 3385 55375 3390
rect 55335 3380 55340 3385
rect 55260 3360 55340 3380
rect 55260 3355 55265 3360
rect 55225 3350 55265 3355
rect 55335 3355 55340 3360
rect 55370 3380 55375 3385
rect 55445 3385 55485 3390
rect 55445 3380 55450 3385
rect 55370 3360 55450 3380
rect 55370 3355 55375 3360
rect 55335 3350 55375 3355
rect 55445 3355 55450 3360
rect 55480 3380 55485 3385
rect 55555 3385 55595 3390
rect 55555 3380 55560 3385
rect 55480 3360 55560 3380
rect 55480 3355 55485 3360
rect 55445 3350 55485 3355
rect 55555 3355 55560 3360
rect 55590 3355 55595 3385
rect 56440 3360 56445 3390
rect 56475 3385 56480 3390
rect 56660 3390 56700 3395
rect 56660 3385 56665 3390
rect 56475 3365 56665 3385
rect 56475 3360 56480 3365
rect 56440 3355 56480 3360
rect 56660 3360 56665 3365
rect 56695 3385 56700 3390
rect 56880 3390 56920 3395
rect 56880 3385 56885 3390
rect 56695 3365 56885 3385
rect 56695 3360 56700 3365
rect 56660 3355 56700 3360
rect 56880 3360 56885 3365
rect 56915 3385 56920 3390
rect 57100 3390 57140 3395
rect 57100 3385 57105 3390
rect 56915 3365 57105 3385
rect 56915 3360 56920 3365
rect 56880 3355 56920 3360
rect 57100 3360 57105 3365
rect 57135 3385 57140 3390
rect 57320 3390 57360 3395
rect 57320 3385 57325 3390
rect 57135 3365 57325 3385
rect 57135 3360 57140 3365
rect 57100 3355 57140 3360
rect 57320 3360 57325 3365
rect 57355 3360 57360 3390
rect 57320 3355 57360 3360
rect 58205 3385 58245 3390
rect 58205 3355 58210 3385
rect 58240 3380 58245 3385
rect 58315 3385 58355 3390
rect 58315 3380 58320 3385
rect 58240 3360 58320 3380
rect 58240 3355 58245 3360
rect 55555 3350 55595 3355
rect 58205 3350 58245 3355
rect 58315 3355 58320 3360
rect 58350 3380 58355 3385
rect 58425 3385 58465 3390
rect 58425 3380 58430 3385
rect 58350 3360 58430 3380
rect 58350 3355 58355 3360
rect 58315 3350 58355 3355
rect 58425 3355 58430 3360
rect 58460 3380 58465 3385
rect 58535 3385 58575 3390
rect 58535 3380 58540 3385
rect 58460 3360 58540 3380
rect 58460 3355 58465 3360
rect 58425 3350 58465 3355
rect 58535 3355 58540 3360
rect 58570 3380 58575 3385
rect 58645 3385 58685 3390
rect 58645 3380 58650 3385
rect 58570 3360 58650 3380
rect 58570 3355 58575 3360
rect 58535 3350 58575 3355
rect 58645 3355 58650 3360
rect 58680 3380 58685 3385
rect 58755 3385 58795 3390
rect 58755 3380 58760 3385
rect 58680 3360 58760 3380
rect 58680 3355 58685 3360
rect 58645 3350 58685 3355
rect 58755 3355 58760 3360
rect 58790 3355 58795 3385
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 58755 3350 58795 3355
rect 57620 3305 57660 3310
rect 56330 3300 56370 3305
rect 56330 3270 56335 3300
rect 56365 3295 56370 3300
rect 56550 3300 56590 3305
rect 56550 3295 56555 3300
rect 56365 3275 56555 3295
rect 56365 3270 56370 3275
rect 56330 3265 56370 3270
rect 56550 3270 56555 3275
rect 56585 3295 56590 3300
rect 56770 3300 56810 3305
rect 56770 3295 56775 3300
rect 56585 3275 56775 3295
rect 56585 3270 56590 3275
rect 56550 3265 56590 3270
rect 56770 3270 56775 3275
rect 56805 3295 56810 3300
rect 56990 3300 57030 3305
rect 56990 3295 56995 3300
rect 56805 3275 56995 3295
rect 56805 3270 56810 3275
rect 56770 3265 56810 3270
rect 56990 3270 56995 3275
rect 57025 3295 57030 3300
rect 57210 3300 57250 3305
rect 57210 3295 57215 3300
rect 57025 3275 57215 3295
rect 57025 3270 57030 3275
rect 56990 3265 57030 3270
rect 57210 3270 57215 3275
rect 57245 3295 57250 3300
rect 57430 3300 57470 3305
rect 57430 3295 57435 3300
rect 57245 3275 57435 3295
rect 57245 3270 57250 3275
rect 57210 3265 57250 3270
rect 57430 3270 57435 3275
rect 57465 3295 57470 3300
rect 57620 3295 57625 3305
rect 57465 3280 57625 3295
rect 57465 3270 57470 3280
rect 57620 3275 57625 3280
rect 57655 3275 57660 3305
rect 57620 3270 57660 3275
rect 57430 3265 57470 3270
rect 56140 3255 56180 3260
rect 56140 3225 56145 3255
rect 56175 3250 56180 3255
rect 56440 3255 56480 3260
rect 56440 3250 56445 3255
rect 56175 3230 56445 3250
rect 56175 3225 56180 3230
rect 56140 3220 56180 3225
rect 56440 3225 56445 3230
rect 56475 3250 56480 3255
rect 56660 3255 56700 3260
rect 56660 3250 56665 3255
rect 56475 3230 56665 3250
rect 56475 3225 56480 3230
rect 56440 3220 56480 3225
rect 56660 3225 56665 3230
rect 56695 3250 56700 3255
rect 56880 3255 56920 3260
rect 56880 3250 56885 3255
rect 56695 3230 56885 3250
rect 56695 3225 56700 3230
rect 56660 3220 56700 3225
rect 56880 3225 56885 3230
rect 56915 3250 56920 3255
rect 57100 3255 57140 3260
rect 57100 3250 57105 3255
rect 56915 3230 57105 3250
rect 56915 3225 56920 3230
rect 56880 3220 56920 3225
rect 57100 3225 57105 3230
rect 57135 3250 57140 3255
rect 57320 3255 57360 3260
rect 57320 3250 57325 3255
rect 57135 3230 57325 3250
rect 57135 3225 57140 3230
rect 57100 3220 57140 3225
rect 57320 3225 57325 3230
rect 57355 3225 57360 3255
rect 57320 3220 57360 3225
rect 56275 3210 56315 3215
rect 56275 3180 56280 3210
rect 56310 3205 56315 3210
rect 56385 3210 56425 3215
rect 56385 3205 56390 3210
rect 56310 3185 56390 3205
rect 56310 3180 56315 3185
rect 56275 3175 56315 3180
rect 56385 3180 56390 3185
rect 56420 3205 56425 3210
rect 56495 3210 56535 3215
rect 56495 3205 56500 3210
rect 56420 3185 56500 3205
rect 56420 3180 56425 3185
rect 56385 3175 56425 3180
rect 56495 3180 56500 3185
rect 56530 3205 56535 3210
rect 56605 3210 56645 3215
rect 56605 3205 56610 3210
rect 56530 3185 56610 3205
rect 56530 3180 56535 3185
rect 56495 3175 56535 3180
rect 56605 3180 56610 3185
rect 56640 3205 56645 3210
rect 56715 3210 56755 3215
rect 56715 3205 56720 3210
rect 56640 3185 56720 3205
rect 56640 3180 56645 3185
rect 56605 3175 56645 3180
rect 56715 3180 56720 3185
rect 56750 3205 56755 3210
rect 56825 3210 56865 3215
rect 56825 3205 56830 3210
rect 56750 3185 56830 3205
rect 56750 3180 56755 3185
rect 56715 3175 56755 3180
rect 56825 3180 56830 3185
rect 56860 3205 56865 3210
rect 56935 3210 56975 3215
rect 56935 3205 56940 3210
rect 56860 3185 56940 3205
rect 56860 3180 56865 3185
rect 56825 3175 56865 3180
rect 56935 3180 56940 3185
rect 56970 3205 56975 3210
rect 57045 3210 57085 3215
rect 57045 3205 57050 3210
rect 56970 3185 57050 3205
rect 56970 3180 56975 3185
rect 56935 3175 56975 3180
rect 57045 3180 57050 3185
rect 57080 3205 57085 3210
rect 57155 3210 57195 3215
rect 57155 3205 57160 3210
rect 57080 3185 57160 3205
rect 57080 3180 57085 3185
rect 57045 3175 57085 3180
rect 57155 3180 57160 3185
rect 57190 3205 57195 3210
rect 57265 3210 57305 3215
rect 57265 3205 57270 3210
rect 57190 3185 57270 3205
rect 57190 3180 57195 3185
rect 57155 3175 57195 3180
rect 57265 3180 57270 3185
rect 57300 3205 57305 3210
rect 57375 3210 57415 3215
rect 57375 3205 57380 3210
rect 57300 3185 57380 3205
rect 57300 3180 57305 3185
rect 57265 3175 57305 3180
rect 57375 3180 57380 3185
rect 57410 3205 57415 3210
rect 57485 3210 57525 3215
rect 57485 3205 57490 3210
rect 57410 3185 57490 3205
rect 57410 3180 57415 3185
rect 57375 3175 57415 3180
rect 57485 3180 57490 3185
rect 57520 3180 57525 3210
rect 57485 3175 57525 3180
rect 56030 3120 56070 3125
rect 56030 3090 56035 3120
rect 56065 3115 56070 3120
rect 56690 3120 56730 3125
rect 56690 3115 56695 3120
rect 56065 3095 56695 3115
rect 56065 3090 56070 3095
rect 56030 3085 56070 3090
rect 56690 3090 56695 3095
rect 56725 3090 56730 3120
rect 56690 3085 56730 3090
rect 57070 3120 57110 3125
rect 57070 3090 57075 3120
rect 57105 3115 57110 3120
rect 57730 3120 57770 3125
rect 57730 3115 57735 3120
rect 57105 3095 57735 3115
rect 57105 3090 57110 3095
rect 57070 3085 57110 3090
rect 57730 3090 57735 3095
rect 57765 3090 57770 3120
rect 57730 3085 57770 3090
rect 56140 3075 56180 3080
rect 55935 3070 55975 3075
rect 55935 3040 55940 3070
rect 55970 3065 55975 3070
rect 55990 3070 56020 3075
rect 55970 3045 55990 3065
rect 55970 3040 55975 3045
rect 55935 3035 55975 3040
rect 56140 3045 56145 3075
rect 56175 3070 56180 3075
rect 56250 3075 56290 3080
rect 56250 3070 56255 3075
rect 56175 3050 56255 3070
rect 56175 3045 56180 3050
rect 56140 3040 56180 3045
rect 56250 3045 56255 3050
rect 56285 3070 56290 3075
rect 56360 3075 56400 3080
rect 56360 3070 56365 3075
rect 56285 3050 56365 3070
rect 56285 3045 56290 3050
rect 56250 3040 56290 3045
rect 56360 3045 56365 3050
rect 56395 3070 56400 3075
rect 56470 3075 56510 3080
rect 56470 3070 56475 3075
rect 56395 3050 56475 3070
rect 56395 3045 56400 3050
rect 56360 3040 56400 3045
rect 56470 3045 56475 3050
rect 56505 3070 56510 3075
rect 56580 3075 56620 3080
rect 57180 3075 57220 3080
rect 56580 3070 56585 3075
rect 56505 3050 56585 3070
rect 56505 3045 56510 3050
rect 56470 3040 56510 3045
rect 56580 3045 56585 3050
rect 56615 3045 56620 3075
rect 56580 3040 56620 3045
rect 56740 3070 56770 3075
rect 57030 3070 57060 3075
rect 56770 3045 57030 3065
rect 55990 3035 56020 3040
rect 56740 3035 56770 3040
rect 57180 3045 57185 3075
rect 57215 3070 57220 3075
rect 57290 3075 57330 3080
rect 57290 3070 57295 3075
rect 57215 3050 57295 3070
rect 57215 3045 57220 3050
rect 57180 3040 57220 3045
rect 57290 3045 57295 3050
rect 57325 3070 57330 3075
rect 57400 3075 57440 3080
rect 57400 3070 57405 3075
rect 57325 3050 57405 3070
rect 57325 3045 57330 3050
rect 57290 3040 57330 3045
rect 57400 3045 57405 3050
rect 57435 3070 57440 3075
rect 57510 3075 57550 3080
rect 57510 3070 57515 3075
rect 57435 3050 57515 3070
rect 57435 3045 57440 3050
rect 57400 3040 57440 3045
rect 57510 3045 57515 3050
rect 57545 3070 57550 3075
rect 57620 3075 57660 3080
rect 57620 3070 57625 3075
rect 57545 3050 57625 3070
rect 57545 3045 57550 3050
rect 57510 3040 57550 3045
rect 57620 3045 57625 3050
rect 57655 3045 57660 3075
rect 57620 3040 57660 3045
rect 57780 3070 57810 3075
rect 57825 3070 57865 3075
rect 57825 3065 57830 3070
rect 57810 3045 57830 3065
rect 57030 3035 57060 3040
rect 57780 3035 57810 3040
rect 57825 3040 57830 3045
rect 57860 3040 57865 3070
rect 57825 3035 57865 3040
rect 56085 3030 56125 3035
rect 56085 3000 56090 3030
rect 56120 3025 56125 3030
rect 56195 3030 56235 3035
rect 56195 3025 56200 3030
rect 56120 3005 56200 3025
rect 56120 3000 56125 3005
rect 56085 2995 56125 3000
rect 56195 3000 56200 3005
rect 56230 3025 56235 3030
rect 56305 3030 56345 3035
rect 56305 3025 56310 3030
rect 56230 3005 56310 3025
rect 56230 3000 56235 3005
rect 56195 2995 56235 3000
rect 56305 3000 56310 3005
rect 56340 3025 56345 3030
rect 56415 3030 56455 3035
rect 56415 3025 56420 3030
rect 56340 3005 56420 3025
rect 56340 3000 56345 3005
rect 56305 2995 56345 3000
rect 56415 3000 56420 3005
rect 56450 3025 56455 3030
rect 56525 3030 56565 3035
rect 56525 3025 56530 3030
rect 56450 3005 56530 3025
rect 56450 3000 56455 3005
rect 56415 2995 56455 3000
rect 56525 3000 56530 3005
rect 56560 3025 56565 3030
rect 56635 3030 56675 3035
rect 56635 3025 56640 3030
rect 56560 3005 56640 3025
rect 56560 3000 56565 3005
rect 56525 2995 56565 3000
rect 56635 3000 56640 3005
rect 56670 3000 56675 3030
rect 56635 2995 56675 3000
rect 57125 3030 57165 3035
rect 57125 3000 57130 3030
rect 57160 3025 57165 3030
rect 57345 3030 57385 3035
rect 57345 3025 57350 3030
rect 57160 3005 57350 3025
rect 57160 3000 57165 3005
rect 57125 2995 57165 3000
rect 57345 3000 57350 3005
rect 57380 3025 57385 3030
rect 57565 3030 57605 3035
rect 57565 3025 57570 3030
rect 57380 3005 57570 3025
rect 57380 3000 57385 3005
rect 57345 2995 57385 3000
rect 57565 3000 57570 3005
rect 57600 3000 57605 3030
rect 57565 2995 57605 3000
rect 56140 2940 56180 2945
rect 56140 2910 56145 2940
rect 56175 2935 56180 2940
rect 56250 2940 56290 2945
rect 56250 2935 56255 2940
rect 56175 2915 56255 2935
rect 56175 2910 56180 2915
rect 56140 2905 56180 2910
rect 56250 2910 56255 2915
rect 56285 2935 56290 2940
rect 56360 2940 56400 2945
rect 56360 2935 56365 2940
rect 56285 2915 56365 2935
rect 56285 2910 56290 2915
rect 56250 2905 56290 2910
rect 56360 2910 56365 2915
rect 56395 2935 56400 2940
rect 56470 2940 56510 2945
rect 56470 2935 56475 2940
rect 56395 2915 56475 2935
rect 56395 2910 56400 2915
rect 56360 2905 56400 2910
rect 56470 2910 56475 2915
rect 56505 2935 56510 2940
rect 56580 2940 56620 2945
rect 56580 2935 56585 2940
rect 56505 2915 56585 2935
rect 56505 2910 56510 2915
rect 56470 2905 56510 2910
rect 56580 2910 56585 2915
rect 56615 2910 56620 2940
rect 56580 2905 56620 2910
rect 57180 2940 57220 2945
rect 57180 2910 57185 2940
rect 57215 2935 57220 2940
rect 57290 2940 57330 2945
rect 57290 2935 57295 2940
rect 57215 2915 57295 2935
rect 57215 2910 57220 2915
rect 57180 2905 57220 2910
rect 57290 2910 57295 2915
rect 57325 2935 57330 2940
rect 57400 2940 57440 2945
rect 57400 2935 57405 2940
rect 57325 2915 57405 2935
rect 57325 2910 57330 2915
rect 57290 2905 57330 2910
rect 57400 2910 57405 2915
rect 57435 2935 57440 2940
rect 57510 2940 57550 2945
rect 57510 2935 57515 2940
rect 57435 2915 57515 2935
rect 57435 2910 57440 2915
rect 57400 2905 57440 2910
rect 57510 2910 57515 2915
rect 57545 2935 57550 2940
rect 57620 2940 57660 2945
rect 57620 2935 57625 2940
rect 57545 2915 57625 2935
rect 57545 2910 57550 2915
rect 57510 2905 57550 2910
rect 57620 2910 57625 2915
rect 57655 2910 57660 2940
rect 57620 2905 57660 2910
rect 56085 2895 56125 2900
rect 56085 2865 56090 2895
rect 56120 2890 56125 2895
rect 56195 2895 56235 2900
rect 56195 2890 56200 2895
rect 56120 2870 56200 2890
rect 56120 2865 56125 2870
rect 56085 2860 56125 2865
rect 56195 2865 56200 2870
rect 56230 2890 56235 2895
rect 56305 2895 56345 2900
rect 56305 2890 56310 2895
rect 56230 2870 56310 2890
rect 56230 2865 56235 2870
rect 56195 2860 56235 2865
rect 56305 2865 56310 2870
rect 56340 2890 56345 2895
rect 56415 2895 56455 2900
rect 56415 2890 56420 2895
rect 56340 2870 56420 2890
rect 56340 2865 56345 2870
rect 56305 2860 56345 2865
rect 56415 2865 56420 2870
rect 56450 2890 56455 2895
rect 56525 2895 56565 2900
rect 56525 2890 56530 2895
rect 56450 2870 56530 2890
rect 56450 2865 56455 2870
rect 56415 2860 56455 2865
rect 56525 2865 56530 2870
rect 56560 2890 56565 2895
rect 56635 2895 56675 2900
rect 56635 2890 56640 2895
rect 56560 2870 56640 2890
rect 56560 2865 56565 2870
rect 56525 2860 56565 2865
rect 56635 2865 56640 2870
rect 56670 2890 56675 2895
rect 56795 2895 56835 2900
rect 56795 2890 56800 2895
rect 56670 2870 56800 2890
rect 56670 2865 56675 2870
rect 56635 2860 56675 2865
rect 56795 2865 56800 2870
rect 56830 2865 56835 2895
rect 56795 2860 56835 2865
rect 57125 2895 57165 2900
rect 57125 2865 57130 2895
rect 57160 2890 57165 2895
rect 57345 2895 57385 2900
rect 57345 2890 57350 2895
rect 57160 2870 57350 2890
rect 57160 2865 57165 2870
rect 57125 2860 57165 2865
rect 57345 2865 57350 2870
rect 57380 2890 57385 2895
rect 57565 2895 57605 2900
rect 57565 2890 57570 2895
rect 57380 2870 57570 2890
rect 57380 2865 57385 2870
rect 57345 2860 57385 2865
rect 57565 2865 57570 2870
rect 57600 2865 57605 2895
rect 57565 2860 57605 2865
rect 56095 2840 56125 2845
rect 55955 2815 56095 2835
rect 56095 2805 56125 2810
rect 56580 2840 56610 2845
rect 57190 2840 57220 2845
rect 56610 2815 57190 2835
rect 56580 2805 56610 2810
rect 57190 2805 57220 2810
rect 55755 2795 55795 2800
rect 55755 2765 55760 2795
rect 55790 2790 55795 2795
rect 56030 2795 56070 2800
rect 56030 2790 56035 2795
rect 55790 2770 56035 2790
rect 55790 2765 55795 2770
rect 55755 2760 55795 2765
rect 56030 2765 56035 2770
rect 56065 2790 56070 2795
rect 56690 2795 56730 2800
rect 56690 2790 56695 2795
rect 56065 2770 56695 2790
rect 56065 2765 56070 2770
rect 56030 2760 56070 2765
rect 56690 2765 56695 2770
rect 56725 2765 56730 2795
rect 56690 2760 56730 2765
rect 57070 2795 57110 2800
rect 57070 2765 57075 2795
rect 57105 2790 57110 2795
rect 57730 2795 57770 2800
rect 57730 2790 57735 2795
rect 57105 2770 57735 2790
rect 57105 2765 57110 2770
rect 57070 2760 57110 2765
rect 57730 2765 57735 2770
rect 57765 2790 57770 2795
rect 58005 2795 58045 2800
rect 58005 2790 58010 2795
rect 57765 2770 58010 2790
rect 57765 2765 57770 2770
rect 57730 2760 57770 2765
rect 58005 2765 58010 2770
rect 58040 2765 58045 2795
rect 58005 2760 58045 2765
rect 55005 2745 55045 2750
rect 55005 2715 55010 2745
rect 55040 2740 55045 2745
rect 55115 2745 55155 2750
rect 55115 2740 55120 2745
rect 55040 2720 55120 2740
rect 55040 2715 55045 2720
rect 55005 2710 55045 2715
rect 55115 2715 55120 2720
rect 55150 2740 55155 2745
rect 55225 2745 55265 2750
rect 55225 2740 55230 2745
rect 55150 2720 55230 2740
rect 55150 2715 55155 2720
rect 55115 2710 55155 2715
rect 55225 2715 55230 2720
rect 55260 2740 55265 2745
rect 55335 2745 55375 2750
rect 55335 2740 55340 2745
rect 55260 2720 55340 2740
rect 55260 2715 55265 2720
rect 55225 2710 55265 2715
rect 55335 2715 55340 2720
rect 55370 2740 55375 2745
rect 55445 2745 55485 2750
rect 55445 2740 55450 2745
rect 55370 2720 55450 2740
rect 55370 2715 55375 2720
rect 55335 2710 55375 2715
rect 55445 2715 55450 2720
rect 55480 2740 55485 2745
rect 55555 2745 55595 2750
rect 55555 2740 55560 2745
rect 55480 2720 55560 2740
rect 55480 2715 55485 2720
rect 55445 2710 55485 2715
rect 55555 2715 55560 2720
rect 55590 2715 55595 2745
rect 58205 2745 58245 2750
rect 55555 2710 55595 2715
rect 56605 2735 56645 2740
rect 56605 2705 56610 2735
rect 56640 2730 56645 2735
rect 56825 2735 56865 2740
rect 56825 2730 56830 2735
rect 56640 2710 56830 2730
rect 56640 2705 56645 2710
rect 54950 2700 54990 2705
rect 54950 2670 54955 2700
rect 54985 2695 54990 2700
rect 55060 2700 55100 2705
rect 55060 2695 55065 2700
rect 54985 2675 55065 2695
rect 54985 2670 54990 2675
rect 54950 2665 54990 2670
rect 55060 2670 55065 2675
rect 55095 2695 55100 2700
rect 55170 2700 55210 2705
rect 55170 2695 55175 2700
rect 55095 2675 55175 2695
rect 55095 2670 55100 2675
rect 55060 2665 55100 2670
rect 55170 2670 55175 2675
rect 55205 2695 55210 2700
rect 55280 2700 55320 2705
rect 55280 2695 55285 2700
rect 55205 2675 55285 2695
rect 55205 2670 55210 2675
rect 55170 2665 55210 2670
rect 55280 2670 55285 2675
rect 55315 2695 55320 2700
rect 55390 2700 55430 2705
rect 55390 2695 55395 2700
rect 55315 2675 55395 2695
rect 55315 2670 55320 2675
rect 55280 2665 55320 2670
rect 55390 2670 55395 2675
rect 55425 2695 55430 2700
rect 55500 2700 55540 2705
rect 55500 2695 55505 2700
rect 55425 2675 55505 2695
rect 55425 2670 55430 2675
rect 55390 2665 55430 2670
rect 55500 2670 55505 2675
rect 55535 2695 55540 2700
rect 55610 2700 55650 2705
rect 56605 2700 56645 2705
rect 56825 2705 56830 2710
rect 56860 2730 56865 2735
rect 57045 2735 57085 2740
rect 57045 2730 57050 2735
rect 56860 2710 57050 2730
rect 56860 2705 56865 2710
rect 56825 2700 56865 2705
rect 57045 2705 57050 2710
rect 57080 2730 57085 2735
rect 57235 2735 57275 2740
rect 57235 2730 57240 2735
rect 57080 2710 57240 2730
rect 57080 2705 57085 2710
rect 57045 2700 57085 2705
rect 57235 2705 57240 2710
rect 57270 2730 57275 2735
rect 57455 2735 57495 2740
rect 57455 2730 57460 2735
rect 57270 2710 57460 2730
rect 57270 2705 57275 2710
rect 57235 2700 57275 2705
rect 57455 2705 57460 2710
rect 57490 2730 57495 2735
rect 57675 2735 57715 2740
rect 57675 2730 57680 2735
rect 57490 2710 57680 2730
rect 57490 2705 57495 2710
rect 57455 2700 57495 2705
rect 57675 2705 57680 2710
rect 57710 2705 57715 2735
rect 58205 2715 58210 2745
rect 58240 2740 58245 2745
rect 58315 2745 58355 2750
rect 58315 2740 58320 2745
rect 58240 2720 58320 2740
rect 58240 2715 58245 2720
rect 58205 2710 58245 2715
rect 58315 2715 58320 2720
rect 58350 2740 58355 2745
rect 58425 2745 58465 2750
rect 58425 2740 58430 2745
rect 58350 2720 58430 2740
rect 58350 2715 58355 2720
rect 58315 2710 58355 2715
rect 58425 2715 58430 2720
rect 58460 2740 58465 2745
rect 58535 2745 58575 2750
rect 58535 2740 58540 2745
rect 58460 2720 58540 2740
rect 58460 2715 58465 2720
rect 58425 2710 58465 2715
rect 58535 2715 58540 2720
rect 58570 2740 58575 2745
rect 58645 2745 58685 2750
rect 58645 2740 58650 2745
rect 58570 2720 58650 2740
rect 58570 2715 58575 2720
rect 58535 2710 58575 2715
rect 58645 2715 58650 2720
rect 58680 2740 58685 2745
rect 58755 2745 58795 2750
rect 58755 2740 58760 2745
rect 58680 2720 58760 2740
rect 58680 2715 58685 2720
rect 58645 2710 58685 2715
rect 58755 2715 58760 2720
rect 58790 2715 58795 2745
rect 58755 2710 58795 2715
rect 57675 2700 57715 2705
rect 58150 2700 58190 2705
rect 55610 2695 55615 2700
rect 55535 2675 55615 2695
rect 55535 2670 55540 2675
rect 55500 2665 55540 2670
rect 55610 2670 55615 2675
rect 55645 2670 55650 2700
rect 55610 2665 55650 2670
rect 56550 2680 56590 2685
rect 56550 2650 56555 2680
rect 56585 2675 56590 2680
rect 56660 2680 56700 2685
rect 56660 2675 56665 2680
rect 56585 2655 56665 2675
rect 56585 2650 56590 2655
rect 56550 2645 56590 2650
rect 56660 2650 56665 2655
rect 56695 2675 56700 2680
rect 56770 2680 56810 2685
rect 56770 2675 56775 2680
rect 56695 2655 56775 2675
rect 56695 2650 56700 2655
rect 56660 2645 56700 2650
rect 56770 2650 56775 2655
rect 56805 2675 56810 2680
rect 56880 2680 56920 2685
rect 56880 2675 56885 2680
rect 56805 2655 56885 2675
rect 56805 2650 56810 2655
rect 56770 2645 56810 2650
rect 56880 2650 56885 2655
rect 56915 2675 56920 2680
rect 56990 2680 57030 2685
rect 56990 2675 56995 2680
rect 56915 2655 56995 2675
rect 56915 2650 56920 2655
rect 56880 2645 56920 2650
rect 56990 2650 56995 2655
rect 57025 2675 57030 2680
rect 57100 2680 57140 2685
rect 57100 2675 57105 2680
rect 57025 2655 57105 2675
rect 57025 2650 57030 2655
rect 56990 2645 57030 2650
rect 57100 2650 57105 2655
rect 57135 2675 57140 2680
rect 57210 2680 57250 2685
rect 57210 2675 57215 2680
rect 57135 2655 57215 2675
rect 57135 2650 57140 2655
rect 57100 2645 57140 2650
rect 57210 2650 57215 2655
rect 57245 2650 57250 2680
rect 58150 2670 58155 2700
rect 58185 2695 58190 2700
rect 58260 2700 58300 2705
rect 58260 2695 58265 2700
rect 58185 2675 58265 2695
rect 58185 2670 58190 2675
rect 58150 2665 58190 2670
rect 58260 2670 58265 2675
rect 58295 2695 58300 2700
rect 58370 2700 58410 2705
rect 58370 2695 58375 2700
rect 58295 2675 58375 2695
rect 58295 2670 58300 2675
rect 58260 2665 58300 2670
rect 58370 2670 58375 2675
rect 58405 2695 58410 2700
rect 58480 2700 58520 2705
rect 58480 2695 58485 2700
rect 58405 2675 58485 2695
rect 58405 2670 58410 2675
rect 58370 2665 58410 2670
rect 58480 2670 58485 2675
rect 58515 2695 58520 2700
rect 58590 2700 58630 2705
rect 58590 2695 58595 2700
rect 58515 2675 58595 2695
rect 58515 2670 58520 2675
rect 58480 2665 58520 2670
rect 58590 2670 58595 2675
rect 58625 2695 58630 2700
rect 58700 2700 58740 2705
rect 58700 2695 58705 2700
rect 58625 2675 58705 2695
rect 58625 2670 58630 2675
rect 58590 2665 58630 2670
rect 58700 2670 58705 2675
rect 58735 2695 58740 2700
rect 58810 2700 58850 2705
rect 58810 2695 58815 2700
rect 58735 2675 58815 2695
rect 58735 2670 58740 2675
rect 58700 2665 58740 2670
rect 58810 2670 58815 2675
rect 58845 2670 58850 2700
rect 58810 2665 58850 2670
rect 57210 2645 57250 2650
rect 54605 2640 54645 2645
rect 54605 2610 54610 2640
rect 54640 2635 54645 2640
rect 55310 2640 55350 2645
rect 55310 2635 55315 2640
rect 54640 2615 55315 2635
rect 54640 2610 54645 2615
rect 54605 2605 54645 2610
rect 55310 2610 55315 2615
rect 55345 2635 55350 2640
rect 55710 2640 55750 2645
rect 55710 2635 55715 2640
rect 55345 2615 55715 2635
rect 55345 2610 55350 2615
rect 55310 2605 55350 2610
rect 55710 2610 55715 2615
rect 55745 2635 55750 2640
rect 56305 2640 56345 2645
rect 57455 2640 57495 2645
rect 56305 2635 56310 2640
rect 55745 2615 56310 2635
rect 55745 2610 55750 2615
rect 55710 2605 55750 2610
rect 56305 2610 56310 2615
rect 56340 2610 56345 2640
rect 56305 2605 56345 2610
rect 56715 2635 56755 2640
rect 56715 2605 56720 2635
rect 56750 2630 56755 2635
rect 56935 2635 56975 2640
rect 56935 2630 56940 2635
rect 56750 2610 56940 2630
rect 56750 2605 56755 2610
rect 56715 2600 56755 2605
rect 56935 2605 56940 2610
rect 56970 2630 56975 2635
rect 57155 2635 57195 2640
rect 57155 2630 57160 2635
rect 56970 2610 57160 2630
rect 56970 2605 56975 2610
rect 56935 2600 56975 2605
rect 57155 2605 57160 2610
rect 57190 2630 57195 2635
rect 57345 2635 57385 2640
rect 57345 2630 57350 2635
rect 57190 2610 57350 2630
rect 57190 2605 57195 2610
rect 57155 2600 57195 2605
rect 57345 2605 57350 2610
rect 57380 2605 57385 2635
rect 57455 2610 57460 2640
rect 57490 2635 57495 2640
rect 58050 2640 58090 2645
rect 58050 2635 58055 2640
rect 57490 2615 58055 2635
rect 57490 2610 57495 2615
rect 57455 2605 57495 2610
rect 58050 2610 58055 2615
rect 58085 2635 58090 2640
rect 58450 2640 58490 2645
rect 58450 2635 58455 2640
rect 58085 2615 58455 2635
rect 58085 2610 58090 2615
rect 58050 2605 58090 2610
rect 58450 2610 58455 2615
rect 58485 2635 58490 2640
rect 59155 2640 59195 2645
rect 59155 2635 59160 2640
rect 58485 2615 59160 2635
rect 58485 2610 58490 2615
rect 58450 2605 58490 2610
rect 59155 2610 59160 2615
rect 59190 2610 59195 2640
rect 59155 2605 59195 2610
rect 57345 2600 57385 2605
rect 54295 2595 54335 2600
rect 54295 2565 54300 2595
rect 54330 2590 54335 2595
rect 55445 2595 55485 2600
rect 55445 2590 55450 2595
rect 54330 2570 55450 2590
rect 54330 2565 54335 2570
rect 54295 2560 54335 2565
rect 55445 2565 55450 2570
rect 55480 2565 55485 2595
rect 55445 2560 55485 2565
rect 58315 2595 58355 2600
rect 58315 2565 58320 2595
rect 58350 2590 58355 2595
rect 59465 2595 59505 2600
rect 59465 2590 59470 2595
rect 58350 2570 59470 2590
rect 58350 2565 58355 2570
rect 58315 2560 58355 2565
rect 59465 2565 59470 2570
rect 59500 2565 59505 2595
rect 59465 2560 59505 2565
rect 54950 2545 54990 2550
rect 54950 2515 54955 2545
rect 54985 2540 54990 2545
rect 55610 2545 55650 2550
rect 55610 2540 55615 2545
rect 54985 2520 55615 2540
rect 54985 2515 54990 2520
rect 54950 2510 54990 2515
rect 55610 2515 55615 2520
rect 55645 2540 55650 2545
rect 55755 2545 55795 2550
rect 55755 2540 55760 2545
rect 55645 2520 55760 2540
rect 55645 2515 55650 2520
rect 55610 2510 55650 2515
rect 55755 2515 55760 2520
rect 55790 2515 55795 2545
rect 58005 2545 58045 2550
rect 55755 2510 55795 2515
rect 56550 2515 56590 2520
rect 54245 2500 54285 2505
rect 54245 2470 54250 2500
rect 54280 2495 54285 2500
rect 55005 2500 55045 2505
rect 55005 2495 55010 2500
rect 54280 2475 55010 2495
rect 54280 2470 54285 2475
rect 54245 2465 54285 2470
rect 55005 2470 55010 2475
rect 55040 2495 55045 2500
rect 55115 2500 55155 2505
rect 55115 2495 55120 2500
rect 55040 2475 55120 2495
rect 55040 2470 55045 2475
rect 55005 2465 55045 2470
rect 55115 2470 55120 2475
rect 55150 2495 55155 2500
rect 55225 2500 55265 2505
rect 55225 2495 55230 2500
rect 55150 2475 55230 2495
rect 55150 2470 55155 2475
rect 55115 2465 55155 2470
rect 55225 2470 55230 2475
rect 55260 2495 55265 2500
rect 55335 2500 55375 2505
rect 55335 2495 55340 2500
rect 55260 2475 55340 2495
rect 55260 2470 55265 2475
rect 55225 2465 55265 2470
rect 55335 2470 55340 2475
rect 55370 2495 55375 2500
rect 55445 2500 55485 2505
rect 55445 2495 55450 2500
rect 55370 2475 55450 2495
rect 55370 2470 55375 2475
rect 55335 2465 55375 2470
rect 55445 2470 55450 2475
rect 55480 2495 55485 2500
rect 55555 2500 55595 2505
rect 55555 2495 55560 2500
rect 55480 2475 55560 2495
rect 55480 2470 55485 2475
rect 55445 2465 55485 2470
rect 55555 2470 55560 2475
rect 55590 2470 55595 2500
rect 56550 2485 56555 2515
rect 56585 2510 56590 2515
rect 56660 2515 56700 2520
rect 56660 2510 56665 2515
rect 56585 2490 56665 2510
rect 56585 2485 56590 2490
rect 56550 2480 56590 2485
rect 56660 2485 56665 2490
rect 56695 2510 56700 2515
rect 56770 2515 56810 2520
rect 56770 2510 56775 2515
rect 56695 2490 56775 2510
rect 56695 2485 56700 2490
rect 56660 2480 56700 2485
rect 56770 2485 56775 2490
rect 56805 2510 56810 2515
rect 56880 2515 56920 2520
rect 56880 2510 56885 2515
rect 56805 2490 56885 2510
rect 56805 2485 56810 2490
rect 56770 2480 56810 2485
rect 56880 2485 56885 2490
rect 56915 2510 56920 2515
rect 56990 2515 57030 2520
rect 56990 2510 56995 2515
rect 56915 2490 56995 2510
rect 56915 2485 56920 2490
rect 56880 2480 56920 2485
rect 56990 2485 56995 2490
rect 57025 2510 57030 2515
rect 57100 2515 57140 2520
rect 57100 2510 57105 2515
rect 57025 2490 57105 2510
rect 57025 2485 57030 2490
rect 56990 2480 57030 2485
rect 57100 2485 57105 2490
rect 57135 2510 57140 2515
rect 57210 2515 57250 2520
rect 57210 2510 57215 2515
rect 57135 2490 57215 2510
rect 57135 2485 57140 2490
rect 57100 2480 57140 2485
rect 57210 2485 57215 2490
rect 57245 2510 57250 2515
rect 57915 2515 57955 2520
rect 57915 2510 57920 2515
rect 57245 2490 57920 2510
rect 57245 2485 57250 2490
rect 57210 2480 57250 2485
rect 57915 2485 57920 2490
rect 57950 2485 57955 2515
rect 58005 2515 58010 2545
rect 58040 2540 58045 2545
rect 58150 2545 58190 2550
rect 58150 2540 58155 2545
rect 58040 2520 58155 2540
rect 58040 2515 58045 2520
rect 58005 2510 58045 2515
rect 58150 2515 58155 2520
rect 58185 2540 58190 2545
rect 58810 2545 58850 2550
rect 58810 2540 58815 2545
rect 58185 2520 58815 2540
rect 58185 2515 58190 2520
rect 58150 2510 58190 2515
rect 58810 2515 58815 2520
rect 58845 2515 58850 2545
rect 58810 2510 58850 2515
rect 57915 2480 57955 2485
rect 58205 2500 58245 2505
rect 55555 2465 55595 2470
rect 58205 2470 58210 2500
rect 58240 2495 58245 2500
rect 58315 2500 58355 2505
rect 58315 2495 58320 2500
rect 58240 2475 58320 2495
rect 58240 2470 58245 2475
rect 58205 2465 58245 2470
rect 58315 2470 58320 2475
rect 58350 2495 58355 2500
rect 58425 2500 58465 2505
rect 58425 2495 58430 2500
rect 58350 2475 58430 2495
rect 58350 2470 58355 2475
rect 58315 2465 58355 2470
rect 58425 2470 58430 2475
rect 58460 2495 58465 2500
rect 58535 2500 58575 2505
rect 58535 2495 58540 2500
rect 58460 2475 58540 2495
rect 58460 2470 58465 2475
rect 58425 2465 58465 2470
rect 58535 2470 58540 2475
rect 58570 2495 58575 2500
rect 58645 2500 58685 2505
rect 58645 2495 58650 2500
rect 58570 2475 58650 2495
rect 58570 2470 58575 2475
rect 58535 2465 58575 2470
rect 58645 2470 58650 2475
rect 58680 2495 58685 2500
rect 58755 2500 58795 2505
rect 58755 2495 58760 2500
rect 58680 2475 58760 2495
rect 58680 2470 58685 2475
rect 58645 2465 58685 2470
rect 58755 2470 58760 2475
rect 58790 2495 58795 2500
rect 59515 2500 59555 2505
rect 59515 2495 59520 2500
rect 58790 2475 59520 2495
rect 58790 2470 58795 2475
rect 58755 2465 58795 2470
rect 59515 2470 59520 2475
rect 59550 2470 59555 2500
rect 59515 2465 59555 2470
rect 56605 2460 56645 2465
rect 55060 2455 55100 2460
rect 55060 2425 55065 2455
rect 55095 2450 55100 2455
rect 55170 2455 55210 2460
rect 55170 2450 55175 2455
rect 55095 2430 55175 2450
rect 55095 2425 55100 2430
rect 55060 2420 55100 2425
rect 55170 2425 55175 2430
rect 55205 2450 55210 2455
rect 55280 2455 55320 2460
rect 55280 2450 55285 2455
rect 55205 2430 55285 2450
rect 55205 2425 55210 2430
rect 55170 2420 55210 2425
rect 55280 2425 55285 2430
rect 55315 2450 55320 2455
rect 55390 2455 55430 2460
rect 55390 2450 55395 2455
rect 55315 2430 55395 2450
rect 55315 2425 55320 2430
rect 55280 2420 55320 2425
rect 55390 2425 55395 2430
rect 55425 2450 55430 2455
rect 55500 2455 55540 2460
rect 55500 2450 55505 2455
rect 55425 2430 55505 2450
rect 55425 2425 55430 2430
rect 55390 2420 55430 2425
rect 55500 2425 55505 2430
rect 55535 2425 55540 2455
rect 56605 2430 56610 2460
rect 56640 2455 56645 2460
rect 56825 2460 56865 2465
rect 56825 2455 56830 2460
rect 56640 2435 56830 2455
rect 56640 2430 56645 2435
rect 56605 2425 56645 2430
rect 56825 2430 56830 2435
rect 56860 2455 56865 2460
rect 57045 2460 57085 2465
rect 57045 2455 57050 2460
rect 56860 2435 57050 2455
rect 56860 2430 56865 2435
rect 56825 2425 56865 2430
rect 57045 2430 57050 2435
rect 57080 2455 57085 2460
rect 57870 2460 57910 2465
rect 57870 2455 57875 2460
rect 57080 2435 57875 2455
rect 57080 2430 57085 2435
rect 57045 2425 57085 2430
rect 57870 2430 57875 2435
rect 57905 2430 57910 2460
rect 57870 2425 57910 2430
rect 58260 2455 58300 2460
rect 58260 2425 58265 2455
rect 58295 2450 58300 2455
rect 58370 2455 58410 2460
rect 58370 2450 58375 2455
rect 58295 2430 58375 2450
rect 58295 2425 58300 2430
rect 55500 2420 55540 2425
rect 58260 2420 58300 2425
rect 58370 2425 58375 2430
rect 58405 2450 58410 2455
rect 58480 2455 58520 2460
rect 58480 2450 58485 2455
rect 58405 2430 58485 2450
rect 58405 2425 58410 2430
rect 58370 2420 58410 2425
rect 58480 2425 58485 2430
rect 58515 2450 58520 2455
rect 58590 2455 58630 2460
rect 58590 2450 58595 2455
rect 58515 2430 58595 2450
rect 58515 2425 58520 2430
rect 58480 2420 58520 2425
rect 58590 2425 58595 2430
rect 58625 2450 58630 2455
rect 58700 2455 58740 2460
rect 58700 2450 58705 2455
rect 58625 2430 58705 2450
rect 58625 2425 58630 2430
rect 58590 2420 58630 2425
rect 58700 2425 58705 2430
rect 58735 2425 58740 2455
rect 58700 2420 58740 2425
rect 56715 2415 56755 2420
rect 56715 2385 56720 2415
rect 56750 2410 56755 2415
rect 56935 2415 56975 2420
rect 56935 2410 56940 2415
rect 56750 2390 56940 2410
rect 56750 2385 56755 2390
rect 56715 2380 56755 2385
rect 56935 2385 56940 2390
rect 56970 2410 56975 2415
rect 57155 2415 57195 2420
rect 57155 2410 57160 2415
rect 56970 2390 57160 2410
rect 56970 2385 56975 2390
rect 56935 2380 56975 2385
rect 57155 2385 57160 2390
rect 57190 2385 57195 2415
rect 57155 2380 57195 2385
rect 56030 2315 56070 2320
rect 56030 2285 56035 2315
rect 56065 2310 56070 2315
rect 56690 2315 56730 2320
rect 56690 2310 56695 2315
rect 56065 2290 56695 2310
rect 56065 2285 56070 2290
rect 56030 2280 56070 2285
rect 56690 2285 56695 2290
rect 56725 2285 56730 2315
rect 56690 2280 56730 2285
rect 57070 2315 57110 2320
rect 57070 2285 57075 2315
rect 57105 2310 57110 2315
rect 57730 2315 57770 2320
rect 57730 2310 57735 2315
rect 57105 2290 57735 2310
rect 57105 2285 57110 2290
rect 57070 2280 57110 2285
rect 57730 2285 57735 2290
rect 57765 2285 57770 2315
rect 57730 2280 57770 2285
rect 56635 2270 56665 2275
rect 56140 2260 56180 2265
rect 56140 2230 56145 2260
rect 56175 2255 56180 2260
rect 56250 2260 56290 2265
rect 56250 2255 56255 2260
rect 56175 2235 56255 2255
rect 56175 2230 56180 2235
rect 56140 2225 56180 2230
rect 56250 2230 56255 2235
rect 56285 2255 56290 2260
rect 56360 2260 56400 2265
rect 56360 2255 56365 2260
rect 56285 2235 56365 2255
rect 56285 2230 56290 2235
rect 56250 2225 56290 2230
rect 56360 2230 56365 2235
rect 56395 2255 56400 2260
rect 56470 2260 56510 2265
rect 56470 2255 56475 2260
rect 56395 2235 56475 2255
rect 56395 2230 56400 2235
rect 56360 2225 56400 2230
rect 56470 2230 56475 2235
rect 56505 2255 56510 2260
rect 56580 2260 56620 2265
rect 56580 2255 56585 2260
rect 56505 2235 56585 2255
rect 56505 2230 56510 2235
rect 56470 2225 56510 2230
rect 56580 2230 56585 2235
rect 56615 2230 56620 2260
rect 57135 2270 57165 2275
rect 56665 2245 57135 2265
rect 56635 2235 56665 2240
rect 57135 2235 57165 2240
rect 57180 2260 57220 2265
rect 56580 2225 56620 2230
rect 57180 2230 57185 2260
rect 57215 2255 57220 2260
rect 57290 2260 57330 2265
rect 57290 2255 57295 2260
rect 57215 2235 57295 2255
rect 57215 2230 57220 2235
rect 57180 2225 57220 2230
rect 57290 2230 57295 2235
rect 57325 2255 57330 2260
rect 57400 2260 57440 2265
rect 57400 2255 57405 2260
rect 57325 2235 57405 2255
rect 57325 2230 57330 2235
rect 57290 2225 57330 2230
rect 57400 2230 57405 2235
rect 57435 2255 57440 2260
rect 57510 2260 57550 2265
rect 57510 2255 57515 2260
rect 57435 2235 57515 2255
rect 57435 2230 57440 2235
rect 57400 2225 57440 2230
rect 57510 2230 57515 2235
rect 57545 2255 57550 2260
rect 57620 2260 57660 2265
rect 57620 2255 57625 2260
rect 57545 2235 57625 2255
rect 57545 2230 57550 2235
rect 57510 2225 57550 2230
rect 57620 2230 57625 2235
rect 57655 2230 57660 2260
rect 57620 2225 57660 2230
rect 57785 2245 57815 2250
rect 56085 2215 56125 2220
rect 54760 2200 54800 2205
rect 54760 2170 54765 2200
rect 54795 2195 54800 2200
rect 55060 2200 55100 2205
rect 55060 2195 55065 2200
rect 54795 2175 55065 2195
rect 54795 2170 54800 2175
rect 54760 2165 54800 2170
rect 55060 2170 55065 2175
rect 55095 2195 55100 2200
rect 55170 2200 55210 2205
rect 55170 2195 55175 2200
rect 55095 2175 55175 2195
rect 55095 2170 55100 2175
rect 55060 2165 55100 2170
rect 55170 2170 55175 2175
rect 55205 2195 55210 2200
rect 55280 2200 55320 2205
rect 55280 2195 55285 2200
rect 55205 2175 55285 2195
rect 55205 2170 55210 2175
rect 55170 2165 55210 2170
rect 55280 2170 55285 2175
rect 55315 2195 55320 2200
rect 55390 2200 55430 2205
rect 55390 2195 55395 2200
rect 55315 2175 55395 2195
rect 55315 2170 55320 2175
rect 55280 2165 55320 2170
rect 55390 2170 55395 2175
rect 55425 2195 55430 2200
rect 55500 2200 55540 2205
rect 55500 2195 55505 2200
rect 55425 2175 55505 2195
rect 55425 2170 55430 2175
rect 55390 2165 55430 2170
rect 55500 2170 55505 2175
rect 55535 2170 55540 2200
rect 56085 2185 56090 2215
rect 56120 2210 56125 2215
rect 56195 2215 56235 2220
rect 56195 2210 56200 2215
rect 56120 2190 56200 2210
rect 56120 2185 56125 2190
rect 56085 2180 56125 2185
rect 56195 2185 56200 2190
rect 56230 2210 56235 2215
rect 56305 2215 56345 2220
rect 56305 2210 56310 2215
rect 56230 2190 56310 2210
rect 56230 2185 56235 2190
rect 56195 2180 56235 2185
rect 56305 2185 56310 2190
rect 56340 2210 56345 2215
rect 56415 2215 56455 2220
rect 56415 2210 56420 2215
rect 56340 2190 56420 2210
rect 56340 2185 56345 2190
rect 56305 2180 56345 2185
rect 56415 2185 56420 2190
rect 56450 2210 56455 2215
rect 56525 2215 56565 2220
rect 56525 2210 56530 2215
rect 56450 2190 56530 2210
rect 56450 2185 56455 2190
rect 56415 2180 56455 2185
rect 56525 2185 56530 2190
rect 56560 2210 56565 2215
rect 56635 2215 56675 2220
rect 56635 2210 56640 2215
rect 56560 2190 56640 2210
rect 56560 2185 56565 2190
rect 56525 2180 56565 2185
rect 56635 2185 56640 2190
rect 56670 2185 56675 2215
rect 56635 2180 56675 2185
rect 57125 2215 57165 2220
rect 57125 2185 57130 2215
rect 57160 2210 57165 2215
rect 57235 2215 57275 2220
rect 57235 2210 57240 2215
rect 57160 2190 57240 2210
rect 57160 2185 57165 2190
rect 57125 2180 57165 2185
rect 57235 2185 57240 2190
rect 57270 2210 57275 2215
rect 57345 2215 57385 2220
rect 57345 2210 57350 2215
rect 57270 2190 57350 2210
rect 57270 2185 57275 2190
rect 57235 2180 57275 2185
rect 57345 2185 57350 2190
rect 57380 2210 57385 2215
rect 57455 2215 57495 2220
rect 57455 2210 57460 2215
rect 57380 2190 57460 2210
rect 57380 2185 57385 2190
rect 57345 2180 57385 2185
rect 57455 2185 57460 2190
rect 57490 2210 57495 2215
rect 57565 2215 57605 2220
rect 57565 2210 57570 2215
rect 57490 2190 57570 2210
rect 57490 2185 57495 2190
rect 57455 2180 57495 2185
rect 57565 2185 57570 2190
rect 57600 2210 57605 2215
rect 57675 2215 57715 2220
rect 57675 2210 57680 2215
rect 57600 2190 57680 2210
rect 57600 2185 57605 2190
rect 57565 2180 57605 2185
rect 57675 2185 57680 2190
rect 57710 2185 57715 2215
rect 57960 2245 58000 2250
rect 57960 2240 57965 2245
rect 57815 2220 57965 2240
rect 57785 2210 57815 2215
rect 57960 2215 57965 2220
rect 57995 2215 58000 2245
rect 57960 2210 58000 2215
rect 57675 2180 57715 2185
rect 58260 2200 58300 2205
rect 55500 2165 55540 2170
rect 58260 2170 58265 2200
rect 58295 2195 58300 2200
rect 58370 2200 58410 2205
rect 58370 2195 58375 2200
rect 58295 2175 58375 2195
rect 58295 2170 58300 2175
rect 58260 2165 58300 2170
rect 58370 2170 58375 2175
rect 58405 2195 58410 2200
rect 58480 2200 58520 2205
rect 58480 2195 58485 2200
rect 58405 2175 58485 2195
rect 58405 2170 58410 2175
rect 58370 2165 58410 2170
rect 58480 2170 58485 2175
rect 58515 2195 58520 2200
rect 58590 2200 58630 2205
rect 58590 2195 58595 2200
rect 58515 2175 58595 2195
rect 58515 2170 58520 2175
rect 58480 2165 58520 2170
rect 58590 2170 58595 2175
rect 58625 2195 58630 2200
rect 58700 2200 58740 2205
rect 58700 2195 58705 2200
rect 58625 2175 58705 2195
rect 58625 2170 58630 2175
rect 58590 2165 58630 2170
rect 58700 2170 58705 2175
rect 58735 2195 58740 2200
rect 59000 2200 59040 2205
rect 59000 2195 59005 2200
rect 58735 2175 59005 2195
rect 58735 2170 58740 2175
rect 58700 2165 58740 2170
rect 59000 2170 59005 2175
rect 59035 2170 59040 2200
rect 59000 2165 59040 2170
rect 55005 2155 55045 2160
rect 55005 2125 55010 2155
rect 55040 2150 55045 2155
rect 55115 2155 55155 2160
rect 55115 2150 55120 2155
rect 55040 2130 55120 2150
rect 55040 2125 55045 2130
rect 55005 2120 55045 2125
rect 55115 2125 55120 2130
rect 55150 2150 55155 2155
rect 55225 2155 55265 2160
rect 55225 2150 55230 2155
rect 55150 2130 55230 2150
rect 55150 2125 55155 2130
rect 55115 2120 55155 2125
rect 55225 2125 55230 2130
rect 55260 2150 55265 2155
rect 55335 2155 55375 2160
rect 55335 2150 55340 2155
rect 55260 2130 55340 2150
rect 55260 2125 55265 2130
rect 55225 2120 55265 2125
rect 55335 2125 55340 2130
rect 55370 2150 55375 2155
rect 55445 2155 55485 2160
rect 55445 2150 55450 2155
rect 55370 2130 55450 2150
rect 55370 2125 55375 2130
rect 55335 2120 55375 2125
rect 55445 2125 55450 2130
rect 55480 2150 55485 2155
rect 55555 2155 55595 2160
rect 55555 2150 55560 2155
rect 55480 2130 55560 2150
rect 55480 2125 55485 2130
rect 55445 2120 55485 2125
rect 55555 2125 55560 2130
rect 55590 2125 55595 2155
rect 55555 2120 55595 2125
rect 58205 2155 58245 2160
rect 58205 2125 58210 2155
rect 58240 2150 58245 2155
rect 58315 2155 58355 2160
rect 58315 2150 58320 2155
rect 58240 2130 58320 2150
rect 58240 2125 58245 2130
rect 58205 2120 58245 2125
rect 58315 2125 58320 2130
rect 58350 2150 58355 2155
rect 58425 2155 58465 2160
rect 58425 2150 58430 2155
rect 58350 2130 58430 2150
rect 58350 2125 58355 2130
rect 58315 2120 58355 2125
rect 58425 2125 58430 2130
rect 58460 2150 58465 2155
rect 58535 2155 58575 2160
rect 58535 2150 58540 2155
rect 58460 2130 58540 2150
rect 58460 2125 58465 2130
rect 58425 2120 58465 2125
rect 58535 2125 58540 2130
rect 58570 2150 58575 2155
rect 58645 2155 58685 2160
rect 58645 2150 58650 2155
rect 58570 2130 58650 2150
rect 58570 2125 58575 2130
rect 58535 2120 58575 2125
rect 58645 2125 58650 2130
rect 58680 2150 58685 2155
rect 58755 2155 58795 2160
rect 58755 2150 58760 2155
rect 58680 2130 58760 2150
rect 58680 2125 58685 2130
rect 58645 2120 58685 2125
rect 58755 2125 58760 2130
rect 58790 2125 58795 2155
rect 58755 2120 58795 2125
rect 54950 2110 54990 2115
rect 54950 2080 54955 2110
rect 54985 2105 54990 2110
rect 55610 2110 55650 2115
rect 55610 2105 55615 2110
rect 54985 2085 55615 2105
rect 54985 2080 54990 2085
rect 54950 2075 54990 2080
rect 55610 2080 55615 2085
rect 55645 2080 55650 2110
rect 55610 2075 55650 2080
rect 58150 2110 58190 2115
rect 58150 2080 58155 2110
rect 58185 2105 58190 2110
rect 58810 2110 58850 2115
rect 58810 2105 58815 2110
rect 58185 2085 58815 2105
rect 58185 2080 58190 2085
rect 58150 2075 58190 2080
rect 58810 2080 58815 2085
rect 58845 2080 58850 2110
rect 58810 2075 58850 2080
rect 55310 2050 55350 2055
rect 55310 2020 55315 2050
rect 55345 2045 55350 2050
rect 55710 2050 55750 2055
rect 55710 2045 55715 2050
rect 55345 2025 55715 2045
rect 55345 2020 55350 2025
rect 55310 2015 55350 2020
rect 55710 2020 55715 2025
rect 55745 2020 55750 2050
rect 58050 2050 58090 2055
rect 55710 2015 55750 2020
rect 56140 2025 56180 2030
rect 56140 1995 56145 2025
rect 56175 2020 56180 2025
rect 56250 2025 56290 2030
rect 56250 2020 56255 2025
rect 56175 2000 56255 2020
rect 56175 1995 56180 2000
rect 56140 1990 56180 1995
rect 56250 1995 56255 2000
rect 56285 2020 56290 2025
rect 56360 2025 56400 2030
rect 56360 2020 56365 2025
rect 56285 2000 56365 2020
rect 56285 1995 56290 2000
rect 56250 1990 56290 1995
rect 56360 1995 56365 2000
rect 56395 2020 56400 2025
rect 56470 2025 56510 2030
rect 56470 2020 56475 2025
rect 56395 2000 56475 2020
rect 56395 1995 56400 2000
rect 56360 1990 56400 1995
rect 56470 1995 56475 2000
rect 56505 2020 56510 2025
rect 56580 2025 56620 2030
rect 56580 2020 56585 2025
rect 56505 2000 56585 2020
rect 56505 1995 56510 2000
rect 56470 1990 56510 1995
rect 56580 1995 56585 2000
rect 56615 1995 56620 2025
rect 56580 1990 56620 1995
rect 57180 2025 57220 2030
rect 57180 1995 57185 2025
rect 57215 2020 57220 2025
rect 57290 2025 57330 2030
rect 57290 2020 57295 2025
rect 57215 2000 57295 2020
rect 57215 1995 57220 2000
rect 57180 1990 57220 1995
rect 57290 1995 57295 2000
rect 57325 2020 57330 2025
rect 57400 2025 57440 2030
rect 57400 2020 57405 2025
rect 57325 2000 57405 2020
rect 57325 1995 57330 2000
rect 57290 1990 57330 1995
rect 57400 1995 57405 2000
rect 57435 2020 57440 2025
rect 57510 2025 57550 2030
rect 57510 2020 57515 2025
rect 57435 2000 57515 2020
rect 57435 1995 57440 2000
rect 57400 1990 57440 1995
rect 57510 1995 57515 2000
rect 57545 2020 57550 2025
rect 57620 2025 57660 2030
rect 57620 2020 57625 2025
rect 57545 2000 57625 2020
rect 57545 1995 57550 2000
rect 57510 1990 57550 1995
rect 57620 1995 57625 2000
rect 57655 1995 57660 2025
rect 58050 2020 58055 2050
rect 58085 2045 58090 2050
rect 58450 2050 58490 2055
rect 58450 2045 58455 2050
rect 58085 2025 58455 2045
rect 58085 2020 58090 2025
rect 58050 2015 58090 2020
rect 58450 2020 58455 2025
rect 58485 2020 58490 2050
rect 58450 2015 58490 2020
rect 57620 1990 57660 1995
rect 54950 1985 54990 1990
rect 54950 1955 54955 1985
rect 54985 1980 54990 1985
rect 55610 1985 55650 1990
rect 58150 1985 58190 1990
rect 55610 1980 55615 1985
rect 54985 1960 55615 1980
rect 54985 1955 54990 1960
rect 54950 1950 54990 1955
rect 55610 1955 55615 1960
rect 55645 1955 55650 1985
rect 55610 1950 55650 1955
rect 56085 1980 56125 1985
rect 56085 1950 56090 1980
rect 56120 1975 56125 1980
rect 56195 1980 56235 1985
rect 56195 1975 56200 1980
rect 56120 1955 56200 1975
rect 56120 1950 56125 1955
rect 56085 1945 56125 1950
rect 56195 1950 56200 1955
rect 56230 1975 56235 1980
rect 56305 1980 56345 1985
rect 56305 1975 56310 1980
rect 56230 1955 56310 1975
rect 56230 1950 56235 1955
rect 56195 1945 56235 1950
rect 56305 1950 56310 1955
rect 56340 1975 56345 1980
rect 56415 1980 56455 1985
rect 56415 1975 56420 1980
rect 56340 1955 56420 1975
rect 56340 1950 56345 1955
rect 56305 1945 56345 1950
rect 56415 1950 56420 1955
rect 56450 1975 56455 1980
rect 56525 1980 56565 1985
rect 56525 1975 56530 1980
rect 56450 1955 56530 1975
rect 56450 1950 56455 1955
rect 56415 1945 56455 1950
rect 56525 1950 56530 1955
rect 56560 1975 56565 1980
rect 56635 1980 56675 1985
rect 56635 1975 56640 1980
rect 56560 1955 56640 1975
rect 56560 1950 56565 1955
rect 56525 1945 56565 1950
rect 56635 1950 56640 1955
rect 56670 1950 56675 1980
rect 56635 1945 56675 1950
rect 57125 1980 57165 1985
rect 57125 1950 57130 1980
rect 57160 1975 57165 1980
rect 57235 1980 57275 1985
rect 57235 1975 57240 1980
rect 57160 1955 57240 1975
rect 57160 1950 57165 1955
rect 57125 1945 57165 1950
rect 57235 1950 57240 1955
rect 57270 1975 57275 1980
rect 57345 1980 57385 1985
rect 57345 1975 57350 1980
rect 57270 1955 57350 1975
rect 57270 1950 57275 1955
rect 57235 1945 57275 1950
rect 57345 1950 57350 1955
rect 57380 1975 57385 1980
rect 57455 1980 57495 1985
rect 57455 1975 57460 1980
rect 57380 1955 57460 1975
rect 57380 1950 57385 1955
rect 57345 1945 57385 1950
rect 57455 1950 57460 1955
rect 57490 1975 57495 1980
rect 57565 1980 57605 1985
rect 57565 1975 57570 1980
rect 57490 1955 57570 1975
rect 57490 1950 57495 1955
rect 57455 1945 57495 1950
rect 57565 1950 57570 1955
rect 57600 1975 57605 1980
rect 57675 1980 57715 1985
rect 57675 1975 57680 1980
rect 57600 1955 57680 1975
rect 57600 1950 57605 1955
rect 57565 1945 57605 1950
rect 57675 1950 57680 1955
rect 57710 1950 57715 1980
rect 58150 1955 58155 1985
rect 58185 1980 58190 1985
rect 58810 1985 58850 1990
rect 58810 1980 58815 1985
rect 58185 1960 58815 1980
rect 58185 1955 58190 1960
rect 58150 1950 58190 1955
rect 58810 1955 58815 1960
rect 58845 1955 58850 1985
rect 58810 1950 58850 1955
rect 57675 1945 57715 1950
rect 55005 1940 55045 1945
rect 54290 1910 54340 1920
rect 54290 1880 54300 1910
rect 54330 1880 54340 1910
rect 55005 1910 55010 1940
rect 55040 1935 55045 1940
rect 55115 1940 55155 1945
rect 55115 1935 55120 1940
rect 55040 1915 55120 1935
rect 55040 1910 55045 1915
rect 55005 1905 55045 1910
rect 55115 1910 55120 1915
rect 55150 1935 55155 1940
rect 55225 1940 55265 1945
rect 55225 1935 55230 1940
rect 55150 1915 55230 1935
rect 55150 1910 55155 1915
rect 55115 1905 55155 1910
rect 55225 1910 55230 1915
rect 55260 1935 55265 1940
rect 55335 1940 55375 1945
rect 55335 1935 55340 1940
rect 55260 1915 55340 1935
rect 55260 1910 55265 1915
rect 55225 1905 55265 1910
rect 55335 1910 55340 1915
rect 55370 1935 55375 1940
rect 55445 1940 55485 1945
rect 55445 1935 55450 1940
rect 55370 1915 55450 1935
rect 55370 1910 55375 1915
rect 55335 1905 55375 1910
rect 55445 1910 55450 1915
rect 55480 1935 55485 1940
rect 55555 1940 55595 1945
rect 58205 1940 58245 1945
rect 55555 1935 55560 1940
rect 55480 1915 55560 1935
rect 55480 1910 55485 1915
rect 55445 1905 55485 1910
rect 55555 1910 55560 1915
rect 55590 1910 55595 1940
rect 55555 1905 55595 1910
rect 55845 1935 55885 1940
rect 55845 1905 55850 1935
rect 55880 1930 55885 1935
rect 56030 1935 56070 1940
rect 56030 1930 56035 1935
rect 55880 1910 56035 1930
rect 55880 1905 55885 1910
rect 55845 1900 55885 1905
rect 56030 1905 56035 1910
rect 56065 1930 56070 1935
rect 56690 1935 56730 1940
rect 56690 1930 56695 1935
rect 56065 1910 56695 1930
rect 56065 1905 56070 1910
rect 56030 1900 56070 1905
rect 56690 1905 56695 1910
rect 56725 1905 56730 1935
rect 56690 1900 56730 1905
rect 57070 1935 57110 1940
rect 57070 1905 57075 1935
rect 57105 1930 57110 1935
rect 57730 1935 57770 1940
rect 57730 1930 57735 1935
rect 57105 1910 57735 1930
rect 57105 1905 57110 1910
rect 57070 1900 57110 1905
rect 57730 1905 57735 1910
rect 57765 1930 57770 1935
rect 57915 1935 57955 1940
rect 57915 1930 57920 1935
rect 57765 1910 57920 1930
rect 57765 1905 57770 1910
rect 57730 1900 57770 1905
rect 57915 1905 57920 1910
rect 57950 1905 57955 1935
rect 58205 1910 58210 1940
rect 58240 1935 58245 1940
rect 58315 1940 58355 1945
rect 58315 1935 58320 1940
rect 58240 1915 58320 1935
rect 58240 1910 58245 1915
rect 58205 1905 58245 1910
rect 58315 1910 58320 1915
rect 58350 1935 58355 1940
rect 58425 1940 58465 1945
rect 58425 1935 58430 1940
rect 58350 1915 58430 1935
rect 58350 1910 58355 1915
rect 58315 1905 58355 1910
rect 58425 1910 58430 1915
rect 58460 1935 58465 1940
rect 58535 1940 58575 1945
rect 58535 1935 58540 1940
rect 58460 1915 58540 1935
rect 58460 1910 58465 1915
rect 58425 1905 58465 1910
rect 58535 1910 58540 1915
rect 58570 1935 58575 1940
rect 58645 1940 58685 1945
rect 58645 1935 58650 1940
rect 58570 1915 58650 1935
rect 58570 1910 58575 1915
rect 58535 1905 58575 1910
rect 58645 1910 58650 1915
rect 58680 1935 58685 1940
rect 58755 1940 58795 1945
rect 58755 1935 58760 1940
rect 58680 1915 58760 1935
rect 58680 1910 58685 1915
rect 58645 1905 58685 1910
rect 58755 1910 58760 1915
rect 58790 1910 58795 1940
rect 58755 1905 58795 1910
rect 59460 1910 59510 1920
rect 57915 1900 57955 1905
rect 54290 1870 54340 1880
rect 54805 1895 54845 1900
rect 54805 1865 54810 1895
rect 54840 1890 54845 1895
rect 55060 1895 55100 1900
rect 55060 1890 55065 1895
rect 54840 1870 55065 1890
rect 54840 1865 54845 1870
rect 54805 1860 54845 1865
rect 55060 1865 55065 1870
rect 55095 1890 55100 1895
rect 55170 1895 55210 1900
rect 55170 1890 55175 1895
rect 55095 1870 55175 1890
rect 55095 1865 55100 1870
rect 55060 1860 55100 1865
rect 55170 1865 55175 1870
rect 55205 1890 55210 1895
rect 55280 1895 55320 1900
rect 55280 1890 55285 1895
rect 55205 1870 55285 1890
rect 55205 1865 55210 1870
rect 55170 1860 55210 1865
rect 55280 1865 55285 1870
rect 55315 1890 55320 1895
rect 55390 1895 55430 1900
rect 55390 1890 55395 1895
rect 55315 1870 55395 1890
rect 55315 1865 55320 1870
rect 55280 1860 55320 1865
rect 55390 1865 55395 1870
rect 55425 1890 55430 1895
rect 55500 1895 55540 1900
rect 55500 1890 55505 1895
rect 55425 1870 55505 1890
rect 55425 1865 55430 1870
rect 55390 1860 55430 1865
rect 55500 1865 55505 1870
rect 55535 1865 55540 1895
rect 55500 1860 55540 1865
rect 58260 1895 58300 1900
rect 58260 1865 58265 1895
rect 58295 1890 58300 1895
rect 58370 1895 58410 1900
rect 58370 1890 58375 1895
rect 58295 1870 58375 1890
rect 58295 1865 58300 1870
rect 58260 1860 58300 1865
rect 58370 1865 58375 1870
rect 58405 1890 58410 1895
rect 58480 1895 58520 1900
rect 58480 1890 58485 1895
rect 58405 1870 58485 1890
rect 58405 1865 58410 1870
rect 58370 1860 58410 1865
rect 58480 1865 58485 1870
rect 58515 1890 58520 1895
rect 58590 1895 58630 1900
rect 58590 1890 58595 1895
rect 58515 1870 58595 1890
rect 58515 1865 58520 1870
rect 58480 1860 58520 1865
rect 58590 1865 58595 1870
rect 58625 1890 58630 1895
rect 58700 1895 58740 1900
rect 58700 1890 58705 1895
rect 58625 1870 58705 1890
rect 58625 1865 58630 1870
rect 58590 1860 58630 1865
rect 58700 1865 58705 1870
rect 58735 1890 58740 1895
rect 58955 1895 58995 1900
rect 58955 1890 58960 1895
rect 58735 1870 58960 1890
rect 58735 1865 58740 1870
rect 58700 1860 58740 1865
rect 58955 1865 58960 1870
rect 58990 1865 58995 1895
rect 59460 1880 59470 1910
rect 59500 1880 59510 1910
rect 59460 1870 59510 1880
rect 58955 1860 58995 1865
rect 56030 1850 56070 1855
rect 56030 1820 56035 1850
rect 56065 1845 56070 1850
rect 56730 1850 56770 1855
rect 56730 1845 56735 1850
rect 56065 1825 56735 1845
rect 56065 1820 56070 1825
rect 56030 1815 56070 1820
rect 56730 1820 56735 1825
rect 56765 1820 56770 1850
rect 57030 1850 57070 1855
rect 56730 1815 56770 1820
rect 56815 1840 56855 1845
rect 56815 1810 56820 1840
rect 56850 1835 56855 1840
rect 56945 1840 56985 1845
rect 56945 1835 56950 1840
rect 56850 1815 56950 1835
rect 56850 1810 56855 1815
rect 56365 1805 56395 1810
rect 56815 1805 56855 1810
rect 56945 1810 56950 1815
rect 56980 1810 56985 1840
rect 57030 1820 57035 1850
rect 57065 1845 57070 1850
rect 57730 1850 57770 1855
rect 57730 1845 57735 1850
rect 57065 1825 57735 1845
rect 57065 1820 57070 1825
rect 57030 1815 57070 1820
rect 57730 1820 57735 1825
rect 57765 1820 57770 1850
rect 57730 1815 57770 1820
rect 56945 1805 56985 1810
rect 57405 1805 57435 1810
rect 56085 1795 56125 1800
rect 55990 1785 56020 1790
rect 55980 1760 55990 1780
rect 56085 1765 56090 1795
rect 56120 1790 56125 1795
rect 56195 1795 56235 1800
rect 56195 1790 56200 1795
rect 56120 1770 56200 1790
rect 56120 1765 56125 1770
rect 56085 1760 56125 1765
rect 56195 1765 56200 1770
rect 56230 1790 56235 1795
rect 56305 1795 56345 1800
rect 56305 1790 56310 1795
rect 56230 1770 56310 1790
rect 56230 1765 56235 1770
rect 56195 1760 56235 1765
rect 56305 1765 56310 1770
rect 56340 1790 56345 1795
rect 56340 1775 56365 1790
rect 56415 1795 56455 1800
rect 56415 1790 56420 1795
rect 56395 1775 56420 1790
rect 56340 1770 56420 1775
rect 56340 1765 56345 1770
rect 56305 1760 56345 1765
rect 56415 1765 56420 1770
rect 56450 1790 56455 1795
rect 56525 1795 56565 1800
rect 56525 1790 56530 1795
rect 56450 1770 56530 1790
rect 56450 1765 56455 1770
rect 56415 1760 56455 1765
rect 56525 1765 56530 1770
rect 56560 1790 56565 1795
rect 56635 1795 56675 1800
rect 56635 1790 56640 1795
rect 56560 1770 56640 1790
rect 56560 1765 56565 1770
rect 56525 1760 56565 1765
rect 56635 1765 56640 1770
rect 56670 1765 56675 1795
rect 57125 1795 57165 1800
rect 56635 1760 56675 1765
rect 56690 1785 56720 1790
rect 56859 1785 56889 1790
rect 56720 1760 56859 1780
rect 55990 1750 56020 1755
rect 56140 1750 56180 1755
rect 56140 1720 56145 1750
rect 56175 1745 56180 1750
rect 56250 1750 56290 1755
rect 56250 1745 56255 1750
rect 56175 1725 56255 1745
rect 56175 1720 56180 1725
rect 56140 1715 56180 1720
rect 56250 1720 56255 1725
rect 56285 1745 56290 1750
rect 56360 1750 56400 1755
rect 56360 1745 56365 1750
rect 56285 1725 56365 1745
rect 56285 1720 56290 1725
rect 56250 1715 56290 1720
rect 56360 1720 56365 1725
rect 56395 1745 56400 1750
rect 56470 1750 56510 1755
rect 56470 1745 56475 1750
rect 56395 1725 56475 1745
rect 56395 1720 56400 1725
rect 56360 1715 56400 1720
rect 56470 1720 56475 1725
rect 56505 1745 56510 1750
rect 56580 1750 56620 1755
rect 56690 1750 56720 1755
rect 56859 1750 56889 1755
rect 56911 1785 56941 1790
rect 56911 1755 56914 1785
rect 57080 1785 57110 1790
rect 56941 1760 57080 1780
rect 56911 1750 56941 1755
rect 57125 1765 57130 1795
rect 57160 1790 57165 1795
rect 57235 1795 57275 1800
rect 57235 1790 57240 1795
rect 57160 1770 57240 1790
rect 57160 1765 57165 1770
rect 57125 1760 57165 1765
rect 57235 1765 57240 1770
rect 57270 1790 57275 1795
rect 57345 1795 57385 1800
rect 57345 1790 57350 1795
rect 57270 1770 57350 1790
rect 57270 1765 57275 1770
rect 57235 1760 57275 1765
rect 57345 1765 57350 1770
rect 57380 1790 57385 1795
rect 57380 1775 57405 1790
rect 57455 1795 57495 1800
rect 57455 1790 57460 1795
rect 57435 1775 57460 1790
rect 57380 1770 57460 1775
rect 57380 1765 57385 1770
rect 57345 1760 57385 1765
rect 57455 1765 57460 1770
rect 57490 1790 57495 1795
rect 57565 1795 57605 1800
rect 57565 1790 57570 1795
rect 57490 1770 57570 1790
rect 57490 1765 57495 1770
rect 57455 1760 57495 1765
rect 57565 1765 57570 1770
rect 57600 1790 57605 1795
rect 57675 1795 57715 1800
rect 57675 1790 57680 1795
rect 57600 1770 57680 1790
rect 57600 1765 57605 1770
rect 57565 1760 57605 1765
rect 57675 1765 57680 1770
rect 57710 1765 57715 1795
rect 57675 1760 57715 1765
rect 57780 1785 57810 1790
rect 57810 1760 57820 1780
rect 57080 1750 57110 1755
rect 57180 1750 57220 1755
rect 56580 1745 56585 1750
rect 56505 1725 56585 1745
rect 56505 1720 56510 1725
rect 56470 1715 56510 1720
rect 56580 1720 56585 1725
rect 56615 1720 56620 1750
rect 56580 1715 56620 1720
rect 57180 1720 57185 1750
rect 57215 1745 57220 1750
rect 57290 1750 57330 1755
rect 57290 1745 57295 1750
rect 57215 1725 57295 1745
rect 57215 1720 57220 1725
rect 57180 1715 57220 1720
rect 57290 1720 57295 1725
rect 57325 1745 57330 1750
rect 57400 1750 57440 1755
rect 57400 1745 57405 1750
rect 57325 1725 57405 1745
rect 57325 1720 57330 1725
rect 57290 1715 57330 1720
rect 57400 1720 57405 1725
rect 57435 1745 57440 1750
rect 57510 1750 57550 1755
rect 57510 1745 57515 1750
rect 57435 1725 57515 1745
rect 57435 1720 57440 1725
rect 57400 1715 57440 1720
rect 57510 1720 57515 1725
rect 57545 1745 57550 1750
rect 57620 1750 57660 1755
rect 57780 1750 57810 1755
rect 57620 1745 57625 1750
rect 57545 1725 57625 1745
rect 57545 1720 57550 1725
rect 57510 1715 57550 1720
rect 57620 1720 57625 1725
rect 57655 1720 57660 1750
rect 57620 1715 57660 1720
rect 55060 1555 55100 1560
rect 54450 1545 54545 1550
rect 54485 1510 54510 1545
rect 54450 1505 54545 1510
rect 54570 1545 54605 1550
rect 54570 1505 54605 1510
rect 54630 1545 54665 1550
rect 54805 1540 54845 1545
rect 54805 1535 54810 1540
rect 54665 1515 54810 1535
rect 54630 1505 54665 1510
rect 54805 1510 54810 1515
rect 54840 1510 54845 1540
rect 55060 1525 55065 1555
rect 55095 1550 55100 1555
rect 55170 1555 55210 1560
rect 55170 1550 55175 1555
rect 55095 1530 55175 1550
rect 55095 1525 55100 1530
rect 55060 1520 55100 1525
rect 55170 1525 55175 1530
rect 55205 1550 55210 1555
rect 55280 1555 55320 1560
rect 55280 1550 55285 1555
rect 55205 1530 55285 1550
rect 55205 1525 55210 1530
rect 55170 1520 55210 1525
rect 55280 1525 55285 1530
rect 55315 1550 55320 1555
rect 55390 1555 55430 1560
rect 55390 1550 55395 1555
rect 55315 1530 55395 1550
rect 55315 1525 55320 1530
rect 55280 1520 55320 1525
rect 55390 1525 55395 1530
rect 55425 1550 55430 1555
rect 55500 1555 55540 1560
rect 55500 1550 55505 1555
rect 55425 1530 55505 1550
rect 55425 1525 55430 1530
rect 55390 1520 55430 1525
rect 55500 1525 55505 1530
rect 55535 1525 55540 1555
rect 55500 1520 55540 1525
rect 56085 1555 56125 1560
rect 56085 1525 56090 1555
rect 56120 1550 56125 1555
rect 56195 1555 56235 1560
rect 56195 1550 56200 1555
rect 56120 1530 56200 1550
rect 56120 1525 56125 1530
rect 56085 1520 56125 1525
rect 56195 1525 56200 1530
rect 56230 1550 56235 1555
rect 56305 1555 56345 1560
rect 56305 1550 56310 1555
rect 56230 1530 56310 1550
rect 56230 1525 56235 1530
rect 56195 1520 56235 1525
rect 56305 1525 56310 1530
rect 56340 1550 56345 1555
rect 56415 1555 56455 1560
rect 56415 1550 56420 1555
rect 56340 1530 56420 1550
rect 56340 1525 56345 1530
rect 56305 1520 56345 1525
rect 56415 1525 56420 1530
rect 56450 1550 56455 1555
rect 56525 1555 56565 1560
rect 56525 1550 56530 1555
rect 56450 1530 56530 1550
rect 56450 1525 56455 1530
rect 56415 1520 56455 1525
rect 56525 1525 56530 1530
rect 56560 1550 56565 1555
rect 56635 1555 56675 1560
rect 56635 1550 56640 1555
rect 56560 1530 56640 1550
rect 56560 1525 56565 1530
rect 56525 1520 56565 1525
rect 56635 1525 56640 1530
rect 56670 1525 56675 1555
rect 56635 1520 56675 1525
rect 57125 1555 57165 1560
rect 57125 1525 57130 1555
rect 57160 1550 57165 1555
rect 57235 1555 57275 1560
rect 57235 1550 57240 1555
rect 57160 1530 57240 1550
rect 57160 1525 57165 1530
rect 57125 1520 57165 1525
rect 57235 1525 57240 1530
rect 57270 1550 57275 1555
rect 57345 1555 57385 1560
rect 57345 1550 57350 1555
rect 57270 1530 57350 1550
rect 57270 1525 57275 1530
rect 57235 1520 57275 1525
rect 57345 1525 57350 1530
rect 57380 1550 57385 1555
rect 57455 1555 57495 1560
rect 57455 1550 57460 1555
rect 57380 1530 57460 1550
rect 57380 1525 57385 1530
rect 57345 1520 57385 1525
rect 57455 1525 57460 1530
rect 57490 1550 57495 1555
rect 57565 1555 57605 1560
rect 57565 1550 57570 1555
rect 57490 1530 57570 1550
rect 57490 1525 57495 1530
rect 57455 1520 57495 1525
rect 57565 1525 57570 1530
rect 57600 1550 57605 1555
rect 57675 1555 57715 1560
rect 57675 1550 57680 1555
rect 57600 1530 57680 1550
rect 57600 1525 57605 1530
rect 57565 1520 57605 1525
rect 57675 1525 57680 1530
rect 57710 1525 57715 1555
rect 57675 1520 57715 1525
rect 58260 1555 58300 1560
rect 58260 1525 58265 1555
rect 58295 1550 58300 1555
rect 58370 1555 58410 1560
rect 58370 1550 58375 1555
rect 58295 1530 58375 1550
rect 58295 1525 58300 1530
rect 58260 1520 58300 1525
rect 58370 1525 58375 1530
rect 58405 1550 58410 1555
rect 58480 1555 58520 1560
rect 58480 1550 58485 1555
rect 58405 1530 58485 1550
rect 58405 1525 58410 1530
rect 58370 1520 58410 1525
rect 58480 1525 58485 1530
rect 58515 1550 58520 1555
rect 58590 1555 58630 1560
rect 58590 1550 58595 1555
rect 58515 1530 58595 1550
rect 58515 1525 58520 1530
rect 58480 1520 58520 1525
rect 58590 1525 58595 1530
rect 58625 1550 58630 1555
rect 58700 1555 58740 1560
rect 58700 1550 58705 1555
rect 58625 1530 58705 1550
rect 58625 1525 58630 1530
rect 58590 1520 58630 1525
rect 58700 1525 58705 1530
rect 58735 1525 58740 1555
rect 59315 1550 59350 1551
rect 59135 1545 59170 1550
rect 58700 1520 58740 1525
rect 58955 1540 58995 1545
rect 54805 1505 54845 1510
rect 55005 1510 55045 1515
rect 54570 1485 54610 1490
rect 54570 1455 54575 1485
rect 54605 1480 54610 1485
rect 54760 1485 54800 1490
rect 54760 1480 54765 1485
rect 54605 1460 54765 1480
rect 54605 1455 54610 1460
rect 54570 1450 54610 1455
rect 54760 1455 54765 1460
rect 54795 1455 54800 1485
rect 55005 1480 55010 1510
rect 55040 1505 55045 1510
rect 55115 1510 55155 1515
rect 55115 1505 55120 1510
rect 55040 1485 55120 1505
rect 55040 1480 55045 1485
rect 55005 1475 55045 1480
rect 55115 1480 55120 1485
rect 55150 1505 55155 1510
rect 55225 1510 55265 1515
rect 55225 1505 55230 1510
rect 55150 1485 55230 1505
rect 55150 1480 55155 1485
rect 55115 1475 55155 1480
rect 55225 1480 55230 1485
rect 55260 1505 55265 1510
rect 55335 1510 55375 1515
rect 55335 1505 55340 1510
rect 55260 1485 55340 1505
rect 55260 1480 55265 1485
rect 55225 1475 55265 1480
rect 55335 1480 55340 1485
rect 55370 1505 55375 1510
rect 55445 1510 55485 1515
rect 55445 1505 55450 1510
rect 55370 1485 55450 1505
rect 55370 1480 55375 1485
rect 55335 1475 55375 1480
rect 55445 1480 55450 1485
rect 55480 1505 55485 1510
rect 55555 1510 55595 1515
rect 55555 1505 55560 1510
rect 55480 1485 55560 1505
rect 55480 1480 55485 1485
rect 55445 1475 55485 1480
rect 55555 1480 55560 1485
rect 55590 1505 55595 1510
rect 55755 1510 55795 1515
rect 55755 1505 55760 1510
rect 55590 1485 55760 1505
rect 55590 1480 55595 1485
rect 55555 1475 55595 1480
rect 55755 1480 55760 1485
rect 55790 1480 55795 1510
rect 55755 1475 55795 1480
rect 56140 1510 56180 1515
rect 56140 1480 56145 1510
rect 56175 1505 56180 1510
rect 56250 1510 56290 1515
rect 56250 1505 56255 1510
rect 56175 1485 56255 1505
rect 56175 1480 56180 1485
rect 56140 1475 56180 1480
rect 56250 1480 56255 1485
rect 56285 1505 56290 1510
rect 56360 1510 56400 1515
rect 56360 1505 56365 1510
rect 56285 1485 56365 1505
rect 56285 1480 56290 1485
rect 56250 1475 56290 1480
rect 56360 1480 56365 1485
rect 56395 1505 56400 1510
rect 56470 1510 56510 1515
rect 56470 1505 56475 1510
rect 56395 1485 56475 1505
rect 56395 1480 56400 1485
rect 56360 1475 56400 1480
rect 56470 1480 56475 1485
rect 56505 1505 56510 1510
rect 56580 1510 56620 1515
rect 56580 1505 56585 1510
rect 56505 1485 56585 1505
rect 56505 1480 56510 1485
rect 56470 1475 56510 1480
rect 56580 1480 56585 1485
rect 56615 1505 56620 1510
rect 57180 1510 57220 1515
rect 57180 1505 57185 1510
rect 56615 1485 57185 1505
rect 56615 1480 56620 1485
rect 56580 1475 56620 1480
rect 57180 1480 57185 1485
rect 57215 1505 57220 1510
rect 57290 1510 57330 1515
rect 57290 1505 57295 1510
rect 57215 1485 57295 1505
rect 57215 1480 57220 1485
rect 57180 1475 57220 1480
rect 57290 1480 57295 1485
rect 57325 1505 57330 1510
rect 57400 1510 57440 1515
rect 57400 1505 57405 1510
rect 57325 1485 57405 1505
rect 57325 1480 57330 1485
rect 57290 1475 57330 1480
rect 57400 1480 57405 1485
rect 57435 1505 57440 1510
rect 57510 1510 57550 1515
rect 57510 1505 57515 1510
rect 57435 1485 57515 1505
rect 57435 1480 57440 1485
rect 57400 1475 57440 1480
rect 57510 1480 57515 1485
rect 57545 1505 57550 1510
rect 57620 1510 57660 1515
rect 57620 1505 57625 1510
rect 57545 1485 57625 1505
rect 57545 1480 57550 1485
rect 57510 1475 57550 1480
rect 57620 1480 57625 1485
rect 57655 1480 57660 1510
rect 57620 1475 57660 1480
rect 58005 1510 58045 1515
rect 58005 1480 58010 1510
rect 58040 1505 58045 1510
rect 58205 1510 58245 1515
rect 58205 1505 58210 1510
rect 58040 1485 58210 1505
rect 58040 1480 58045 1485
rect 58005 1475 58045 1480
rect 58205 1480 58210 1485
rect 58240 1505 58245 1510
rect 58315 1510 58355 1515
rect 58315 1505 58320 1510
rect 58240 1485 58320 1505
rect 58240 1480 58245 1485
rect 58205 1475 58245 1480
rect 58315 1480 58320 1485
rect 58350 1505 58355 1510
rect 58425 1510 58465 1515
rect 58425 1505 58430 1510
rect 58350 1485 58430 1505
rect 58350 1480 58355 1485
rect 58315 1475 58355 1480
rect 58425 1480 58430 1485
rect 58460 1505 58465 1510
rect 58535 1510 58575 1515
rect 58535 1505 58540 1510
rect 58460 1485 58540 1505
rect 58460 1480 58465 1485
rect 58425 1475 58465 1480
rect 58535 1480 58540 1485
rect 58570 1505 58575 1510
rect 58645 1510 58685 1515
rect 58645 1505 58650 1510
rect 58570 1485 58650 1505
rect 58570 1480 58575 1485
rect 58535 1475 58575 1480
rect 58645 1480 58650 1485
rect 58680 1505 58685 1510
rect 58755 1510 58795 1515
rect 58755 1505 58760 1510
rect 58680 1485 58760 1505
rect 58680 1480 58685 1485
rect 58645 1475 58685 1480
rect 58755 1480 58760 1485
rect 58790 1480 58795 1510
rect 58955 1510 58960 1540
rect 58990 1535 58995 1540
rect 58990 1515 59135 1535
rect 58990 1510 58995 1515
rect 58955 1505 58995 1510
rect 59135 1505 59170 1510
rect 59195 1545 59230 1550
rect 59195 1505 59230 1510
rect 59255 1545 59350 1550
rect 59290 1510 59315 1545
rect 59255 1505 59350 1510
rect 58755 1475 58795 1480
rect 59000 1485 59040 1490
rect 54760 1450 54800 1455
rect 54950 1465 54990 1470
rect 54950 1435 54955 1465
rect 54985 1460 54990 1465
rect 55610 1465 55650 1470
rect 55610 1460 55615 1465
rect 54985 1440 55615 1460
rect 54985 1435 54990 1440
rect 54950 1430 54990 1435
rect 55610 1435 55615 1440
rect 55645 1460 55650 1465
rect 55845 1465 55885 1470
rect 55845 1460 55850 1465
rect 55645 1440 55850 1460
rect 55645 1435 55650 1440
rect 55610 1430 55650 1435
rect 55845 1435 55850 1440
rect 55880 1460 55885 1465
rect 56030 1465 56070 1470
rect 56030 1460 56035 1465
rect 55880 1440 56035 1460
rect 55880 1435 55885 1440
rect 55845 1430 55885 1435
rect 56030 1435 56035 1440
rect 56065 1460 56070 1465
rect 56730 1465 56770 1470
rect 56730 1460 56735 1465
rect 56065 1440 56735 1460
rect 56065 1435 56070 1440
rect 56030 1430 56070 1435
rect 56730 1435 56735 1440
rect 56765 1435 56770 1465
rect 56730 1430 56770 1435
rect 57030 1465 57070 1470
rect 57030 1435 57035 1465
rect 57065 1460 57070 1465
rect 57730 1465 57770 1470
rect 57730 1460 57735 1465
rect 57065 1440 57735 1460
rect 57065 1435 57070 1440
rect 57030 1430 57070 1435
rect 57730 1435 57735 1440
rect 57765 1460 57770 1465
rect 57915 1465 57955 1470
rect 57915 1460 57920 1465
rect 57765 1440 57920 1460
rect 57765 1435 57770 1440
rect 57730 1430 57770 1435
rect 57915 1435 57920 1440
rect 57950 1460 57955 1465
rect 58150 1465 58190 1470
rect 58150 1460 58155 1465
rect 57950 1440 58155 1460
rect 57950 1435 57955 1440
rect 57915 1430 57955 1435
rect 58150 1435 58155 1440
rect 58185 1460 58190 1465
rect 58810 1465 58850 1470
rect 58810 1460 58815 1465
rect 58185 1440 58815 1460
rect 58185 1435 58190 1440
rect 58150 1430 58190 1435
rect 58810 1435 58815 1440
rect 58845 1435 58850 1465
rect 59000 1455 59005 1485
rect 59035 1480 59040 1485
rect 59190 1485 59230 1490
rect 59190 1480 59195 1485
rect 59035 1460 59195 1480
rect 59035 1455 59040 1460
rect 59000 1450 59040 1455
rect 59190 1455 59195 1460
rect 59225 1455 59230 1485
rect 59190 1450 59230 1455
rect 58810 1430 58850 1435
rect 54450 1420 54490 1425
rect 54450 1390 54455 1420
rect 54485 1415 54490 1420
rect 55935 1420 55975 1425
rect 55935 1415 55940 1420
rect 54485 1395 55940 1415
rect 54485 1390 54490 1395
rect 54450 1385 54490 1390
rect 55935 1390 55940 1395
rect 55970 1390 55975 1420
rect 55935 1385 55975 1390
rect 56825 1420 56865 1425
rect 56825 1390 56830 1420
rect 56860 1415 56865 1420
rect 56935 1420 56975 1425
rect 56935 1415 56940 1420
rect 56860 1395 56940 1415
rect 56860 1390 56865 1395
rect 56825 1385 56865 1390
rect 56935 1390 56940 1395
rect 56970 1390 56975 1420
rect 56935 1385 56975 1390
rect 57825 1420 57865 1425
rect 57825 1390 57830 1420
rect 57860 1415 57865 1420
rect 59310 1420 59350 1425
rect 59310 1415 59315 1420
rect 57860 1395 59315 1415
rect 57860 1390 57865 1395
rect 57825 1385 57865 1390
rect 59310 1390 59315 1395
rect 59345 1390 59350 1420
rect 59310 1385 59350 1390
rect 54730 1325 54770 1330
rect 54730 1295 54735 1325
rect 54765 1320 54770 1325
rect 55335 1325 55375 1330
rect 55335 1320 55340 1325
rect 54765 1300 55340 1320
rect 54765 1295 54770 1300
rect 54730 1290 54770 1295
rect 55335 1295 55340 1300
rect 55370 1320 55375 1325
rect 58430 1325 58470 1330
rect 58430 1320 58435 1325
rect 55370 1300 58435 1320
rect 55370 1295 55375 1300
rect 55335 1290 55375 1295
rect 58430 1295 58435 1300
rect 58465 1320 58470 1325
rect 59035 1325 59075 1330
rect 59035 1320 59040 1325
rect 58465 1300 59040 1320
rect 58465 1295 58470 1300
rect 58430 1290 58470 1295
rect 59035 1295 59040 1300
rect 59070 1295 59075 1325
rect 59035 1290 59075 1295
rect 56330 1265 56370 1270
rect 54985 1250 55025 1255
rect 54985 1220 54990 1250
rect 55020 1245 55025 1250
rect 55185 1250 55225 1255
rect 55185 1245 55190 1250
rect 55020 1225 55190 1245
rect 55020 1220 55025 1225
rect 54985 1215 55025 1220
rect 55185 1220 55190 1225
rect 55220 1245 55225 1250
rect 55385 1250 55425 1255
rect 55385 1245 55390 1250
rect 55220 1225 55390 1245
rect 55220 1220 55225 1225
rect 55185 1215 55225 1220
rect 55385 1220 55390 1225
rect 55420 1245 55425 1250
rect 55585 1250 55625 1255
rect 55585 1245 55590 1250
rect 55420 1225 55590 1245
rect 55420 1220 55425 1225
rect 55385 1215 55425 1220
rect 55585 1220 55590 1225
rect 55620 1220 55625 1250
rect 56330 1235 56335 1265
rect 56365 1260 56370 1265
rect 56880 1265 56920 1270
rect 56880 1260 56885 1265
rect 56365 1240 56885 1260
rect 56365 1235 56370 1240
rect 56330 1230 56370 1235
rect 56880 1235 56885 1240
rect 56915 1235 56920 1265
rect 56880 1230 56920 1235
rect 57405 1265 57445 1270
rect 57405 1235 57410 1265
rect 57440 1260 57445 1265
rect 57870 1265 57910 1270
rect 57870 1260 57875 1265
rect 57440 1240 57875 1260
rect 57440 1235 57445 1240
rect 57405 1230 57445 1235
rect 57870 1235 57875 1240
rect 57905 1235 57910 1265
rect 57870 1230 57910 1235
rect 58180 1250 58220 1255
rect 55585 1215 55625 1220
rect 58180 1220 58185 1250
rect 58215 1245 58220 1250
rect 58380 1250 58420 1255
rect 58380 1245 58385 1250
rect 58215 1225 58385 1245
rect 58215 1220 58220 1225
rect 58180 1215 58220 1220
rect 58380 1220 58385 1225
rect 58415 1245 58420 1250
rect 58580 1250 58620 1255
rect 58580 1245 58585 1250
rect 58415 1225 58585 1245
rect 58415 1220 58420 1225
rect 58380 1215 58420 1220
rect 58580 1220 58585 1225
rect 58615 1245 58620 1250
rect 58780 1250 58820 1255
rect 58780 1245 58785 1250
rect 58615 1225 58785 1245
rect 58615 1220 58620 1225
rect 58580 1215 58620 1220
rect 58780 1220 58785 1225
rect 58815 1220 58820 1250
rect 58780 1215 58820 1220
rect 56440 1210 56480 1215
rect 54295 1205 54335 1210
rect 54295 1175 54300 1205
rect 54330 1200 54335 1205
rect 54795 1205 54835 1210
rect 54795 1200 54800 1205
rect 54330 1180 54800 1200
rect 54330 1175 54335 1180
rect 54295 1170 54335 1175
rect 54795 1175 54800 1180
rect 54830 1200 54835 1205
rect 55085 1205 55125 1210
rect 55085 1200 55090 1205
rect 54830 1180 55090 1200
rect 54830 1175 54835 1180
rect 54795 1170 54835 1175
rect 55085 1175 55090 1180
rect 55120 1200 55125 1205
rect 55285 1205 55325 1210
rect 55285 1200 55290 1205
rect 55120 1180 55290 1200
rect 55120 1175 55125 1180
rect 55085 1170 55125 1175
rect 55285 1175 55290 1180
rect 55320 1200 55325 1205
rect 55485 1205 55525 1210
rect 55485 1200 55490 1205
rect 55320 1180 55490 1200
rect 55320 1175 55325 1180
rect 55285 1170 55325 1175
rect 55485 1175 55490 1180
rect 55520 1175 55525 1205
rect 56440 1180 56445 1210
rect 56475 1205 56480 1210
rect 56550 1210 56590 1215
rect 56550 1205 56555 1210
rect 56475 1185 56555 1205
rect 56475 1180 56480 1185
rect 56440 1175 56480 1180
rect 56550 1180 56555 1185
rect 56585 1205 56590 1210
rect 56660 1210 56700 1215
rect 56660 1205 56665 1210
rect 56585 1185 56665 1205
rect 56585 1180 56590 1185
rect 56550 1175 56590 1180
rect 56660 1180 56665 1185
rect 56695 1205 56700 1210
rect 56770 1210 56810 1215
rect 56770 1205 56775 1210
rect 56695 1185 56775 1205
rect 56695 1180 56700 1185
rect 56660 1175 56700 1180
rect 56770 1180 56775 1185
rect 56805 1205 56810 1210
rect 56880 1210 56920 1215
rect 56880 1205 56885 1210
rect 56805 1185 56885 1205
rect 56805 1180 56810 1185
rect 56770 1175 56810 1180
rect 56880 1180 56885 1185
rect 56915 1205 56920 1210
rect 56990 1210 57030 1215
rect 56990 1205 56995 1210
rect 56915 1185 56995 1205
rect 56915 1180 56920 1185
rect 56880 1175 56920 1180
rect 56990 1180 56995 1185
rect 57025 1205 57030 1210
rect 57100 1210 57140 1215
rect 57100 1205 57105 1210
rect 57025 1185 57105 1205
rect 57025 1180 57030 1185
rect 56990 1175 57030 1180
rect 57100 1180 57105 1185
rect 57135 1205 57140 1210
rect 57210 1210 57250 1215
rect 57210 1205 57215 1210
rect 57135 1185 57215 1205
rect 57135 1180 57140 1185
rect 57100 1175 57140 1180
rect 57210 1180 57215 1185
rect 57245 1205 57250 1210
rect 57320 1210 57360 1215
rect 57320 1205 57325 1210
rect 57245 1185 57325 1205
rect 57245 1180 57250 1185
rect 57210 1175 57250 1180
rect 57320 1180 57325 1185
rect 57355 1205 57360 1210
rect 57430 1210 57470 1215
rect 57430 1205 57435 1210
rect 57355 1185 57435 1205
rect 57355 1180 57360 1185
rect 57320 1175 57360 1180
rect 57430 1180 57435 1185
rect 57465 1180 57470 1210
rect 57430 1175 57470 1180
rect 58280 1205 58320 1210
rect 58280 1175 58285 1205
rect 58315 1200 58320 1205
rect 58480 1205 58520 1210
rect 58480 1200 58485 1205
rect 58315 1180 58485 1200
rect 58315 1175 58320 1180
rect 55485 1170 55525 1175
rect 58280 1170 58320 1175
rect 58480 1175 58485 1180
rect 58515 1200 58520 1205
rect 58680 1205 58720 1210
rect 58680 1200 58685 1205
rect 58515 1180 58685 1200
rect 58515 1175 58520 1180
rect 58480 1170 58520 1175
rect 58680 1175 58685 1180
rect 58715 1200 58720 1205
rect 58970 1205 59010 1210
rect 58970 1200 58975 1205
rect 58715 1180 58975 1200
rect 58715 1175 58720 1180
rect 58680 1170 58720 1175
rect 58970 1175 58975 1180
rect 59005 1200 59010 1205
rect 59465 1205 59505 1210
rect 59465 1200 59470 1205
rect 59005 1180 59470 1200
rect 59005 1175 59010 1180
rect 58970 1170 59010 1175
rect 59465 1175 59470 1180
rect 59500 1175 59505 1205
rect 59465 1170 59505 1175
rect 54735 1150 54770 1155
rect 54735 1110 54770 1115
rect 54795 1150 54830 1155
rect 54795 1110 54830 1115
rect 58975 1150 59010 1155
rect 58975 1110 59010 1115
rect 59035 1150 59070 1155
rect 59035 1110 59070 1115
rect 55845 890 55885 895
rect 55845 860 55850 890
rect 55880 885 55885 890
rect 56220 890 56260 895
rect 56220 885 56225 890
rect 55880 865 56225 885
rect 55880 860 55885 865
rect 55845 855 55885 860
rect 56220 860 56225 865
rect 56255 885 56260 890
rect 56275 890 56315 895
rect 56275 885 56280 890
rect 56255 865 56280 885
rect 56255 860 56260 865
rect 56220 855 56260 860
rect 56275 860 56280 865
rect 56310 885 56315 890
rect 56385 890 56425 895
rect 56385 885 56390 890
rect 56310 865 56390 885
rect 56310 860 56315 865
rect 56275 855 56315 860
rect 56385 860 56390 865
rect 56420 885 56425 890
rect 56495 890 56535 895
rect 56495 885 56500 890
rect 56420 865 56500 885
rect 56420 860 56425 865
rect 56385 855 56425 860
rect 56495 860 56500 865
rect 56530 885 56535 890
rect 56605 890 56645 895
rect 56605 885 56610 890
rect 56530 865 56610 885
rect 56530 860 56535 865
rect 56495 855 56535 860
rect 56605 860 56610 865
rect 56640 885 56645 890
rect 56715 890 56755 895
rect 56715 885 56720 890
rect 56640 865 56720 885
rect 56640 860 56645 865
rect 56605 855 56645 860
rect 56715 860 56720 865
rect 56750 885 56755 890
rect 56825 890 56865 895
rect 56825 885 56830 890
rect 56750 865 56830 885
rect 56750 860 56755 865
rect 56715 855 56755 860
rect 56825 860 56830 865
rect 56860 885 56865 890
rect 56935 890 56975 895
rect 56935 885 56940 890
rect 56860 865 56940 885
rect 56860 860 56865 865
rect 56825 855 56865 860
rect 56935 860 56940 865
rect 56970 885 56975 890
rect 57045 890 57085 895
rect 57045 885 57050 890
rect 56970 865 57050 885
rect 56970 860 56975 865
rect 56935 855 56975 860
rect 57045 860 57050 865
rect 57080 885 57085 890
rect 57155 890 57195 895
rect 57155 885 57160 890
rect 57080 865 57160 885
rect 57080 860 57085 865
rect 57045 855 57085 860
rect 57155 860 57160 865
rect 57190 885 57195 890
rect 57265 890 57305 895
rect 57265 885 57270 890
rect 57190 865 57270 885
rect 57190 860 57195 865
rect 57155 855 57195 860
rect 57265 860 57270 865
rect 57300 885 57305 890
rect 57375 890 57415 895
rect 57375 885 57380 890
rect 57300 865 57380 885
rect 57300 860 57305 865
rect 57265 855 57305 860
rect 57375 860 57380 865
rect 57410 885 57415 890
rect 57485 890 57525 895
rect 57485 885 57490 890
rect 57410 865 57490 885
rect 57410 860 57415 865
rect 57375 855 57415 860
rect 57485 860 57490 865
rect 57520 885 57525 890
rect 57520 880 57955 885
rect 57520 865 57920 880
rect 57520 860 57525 865
rect 57485 855 57525 860
rect 57915 850 57920 865
rect 57950 850 57955 880
rect 56440 845 56480 850
rect 56440 815 56445 845
rect 56475 840 56480 845
rect 56550 845 56590 850
rect 56550 840 56555 845
rect 56475 820 56555 840
rect 56475 815 56480 820
rect 56440 810 56480 815
rect 56550 815 56555 820
rect 56585 840 56590 845
rect 56660 845 56700 850
rect 56660 840 56665 845
rect 56585 820 56665 840
rect 56585 815 56590 820
rect 56550 810 56590 815
rect 56660 815 56665 820
rect 56695 840 56700 845
rect 56770 845 56810 850
rect 56770 840 56775 845
rect 56695 820 56775 840
rect 56695 815 56700 820
rect 56660 810 56700 815
rect 56770 815 56775 820
rect 56805 840 56810 845
rect 56880 845 56920 850
rect 56880 840 56885 845
rect 56805 820 56885 840
rect 56805 815 56810 820
rect 56770 810 56810 815
rect 56880 815 56885 820
rect 56915 840 56920 845
rect 56990 845 57030 850
rect 56990 840 56995 845
rect 56915 820 56995 840
rect 56915 815 56920 820
rect 56880 810 56920 815
rect 56990 815 56995 820
rect 57025 840 57030 845
rect 57100 845 57140 850
rect 57100 840 57105 845
rect 57025 820 57105 840
rect 57025 815 57030 820
rect 56990 810 57030 815
rect 57100 815 57105 820
rect 57135 840 57140 845
rect 57210 845 57250 850
rect 57210 840 57215 845
rect 57135 820 57215 840
rect 57135 815 57140 820
rect 57100 810 57140 815
rect 57210 815 57215 820
rect 57245 840 57250 845
rect 57320 845 57360 850
rect 57320 840 57325 845
rect 57245 820 57325 840
rect 57245 815 57250 820
rect 57210 810 57250 815
rect 57320 815 57325 820
rect 57355 840 57360 845
rect 57430 845 57470 850
rect 57915 845 57955 850
rect 57430 840 57435 845
rect 57355 820 57435 840
rect 57355 815 57360 820
rect 57320 810 57360 815
rect 57430 815 57435 820
rect 57465 815 57470 845
rect 57430 810 57470 815
rect 56540 790 56580 795
rect 56540 760 56545 790
rect 56575 785 56580 790
rect 56650 790 56690 795
rect 56650 785 56655 790
rect 56575 765 56655 785
rect 56575 760 56580 765
rect 56540 755 56580 760
rect 56650 760 56655 765
rect 56685 785 56690 790
rect 56870 790 56910 795
rect 56870 785 56875 790
rect 56685 765 56875 785
rect 56685 760 56690 765
rect 56650 755 56690 760
rect 56870 760 56875 765
rect 56905 760 56910 790
rect 56870 755 56910 760
rect 56485 745 56525 750
rect 56485 715 56490 745
rect 56520 740 56525 745
rect 56595 745 56635 750
rect 56595 740 56600 745
rect 56520 720 56600 740
rect 56520 715 56525 720
rect 56485 710 56525 715
rect 56595 715 56600 720
rect 56630 740 56635 745
rect 56705 745 56745 750
rect 56705 740 56710 745
rect 56630 720 56710 740
rect 56630 715 56635 720
rect 56595 710 56635 715
rect 56705 715 56710 720
rect 56740 740 56745 745
rect 57040 745 57080 750
rect 57040 740 57045 745
rect 56740 720 57045 740
rect 56740 715 56745 720
rect 56705 710 56745 715
rect 57040 715 57045 720
rect 57075 740 57080 745
rect 57960 745 58000 750
rect 57960 740 57965 745
rect 57075 720 57965 740
rect 57075 715 57080 720
rect 57040 710 57080 715
rect 57960 715 57965 720
rect 57995 715 58000 745
rect 57960 710 58000 715
rect 56540 540 56580 545
rect 56540 510 56545 540
rect 56575 535 56580 540
rect 56650 540 56690 545
rect 56650 535 56655 540
rect 56575 515 56655 535
rect 56575 510 56580 515
rect 56540 505 56580 510
rect 56650 510 56655 515
rect 56685 535 56690 540
rect 56870 540 56910 545
rect 56870 535 56875 540
rect 56685 515 56875 535
rect 56685 510 56690 515
rect 56650 505 56690 510
rect 56870 510 56875 515
rect 56905 510 56910 540
rect 56870 505 56910 510
rect 56485 495 56525 500
rect 55085 465 55125 470
rect 55085 435 55090 465
rect 55120 460 55125 465
rect 55285 465 55325 470
rect 55285 460 55290 465
rect 55120 440 55290 460
rect 55120 435 55125 440
rect 55085 430 55125 435
rect 55285 435 55290 440
rect 55320 460 55325 465
rect 55485 465 55525 470
rect 55485 460 55490 465
rect 55320 440 55490 460
rect 55320 435 55325 440
rect 55285 430 55325 435
rect 55485 435 55490 440
rect 55520 435 55525 465
rect 56485 465 56490 495
rect 56520 490 56525 495
rect 56595 495 56635 500
rect 56595 490 56600 495
rect 56520 470 56600 490
rect 56520 465 56525 470
rect 56485 460 56525 465
rect 56595 465 56600 470
rect 56630 490 56635 495
rect 56705 495 56745 500
rect 56705 490 56710 495
rect 56630 470 56710 490
rect 56630 465 56635 470
rect 56595 460 56635 465
rect 56705 465 56710 470
rect 56740 465 56745 495
rect 56705 460 56745 465
rect 58280 465 58320 470
rect 55485 430 55525 435
rect 58280 435 58285 465
rect 58315 460 58320 465
rect 58480 465 58520 470
rect 58480 460 58485 465
rect 58315 440 58485 460
rect 58315 435 58320 440
rect 58280 430 58320 435
rect 58480 435 58485 440
rect 58515 460 58520 465
rect 58680 465 58720 470
rect 58680 460 58685 465
rect 58515 440 58685 460
rect 58515 435 58520 440
rect 58480 430 58520 435
rect 58680 435 58685 440
rect 58715 435 58720 465
rect 58680 430 58720 435
rect 54245 395 54285 400
rect 54245 365 54250 395
rect 54280 390 54285 395
rect 54985 395 55025 400
rect 54985 390 54990 395
rect 54280 370 54990 390
rect 54280 365 54285 370
rect 54245 360 54285 365
rect 54985 365 54990 370
rect 55020 390 55025 395
rect 55185 395 55225 400
rect 55185 390 55190 395
rect 55020 370 55190 390
rect 55020 365 55025 370
rect 54985 360 55025 365
rect 55185 365 55190 370
rect 55220 390 55225 395
rect 55385 395 55425 400
rect 55385 390 55390 395
rect 55220 370 55390 390
rect 55220 365 55225 370
rect 55185 360 55225 365
rect 55385 365 55390 370
rect 55420 390 55425 395
rect 55585 395 55625 400
rect 55585 390 55590 395
rect 55420 370 55590 390
rect 55420 365 55425 370
rect 55385 360 55425 365
rect 55585 365 55590 370
rect 55620 390 55625 395
rect 55845 395 55885 400
rect 55845 390 55850 395
rect 55620 370 55850 390
rect 55620 365 55625 370
rect 55585 360 55625 365
rect 55845 365 55850 370
rect 55880 390 55885 395
rect 56430 395 56470 400
rect 56430 390 56435 395
rect 55880 370 56435 390
rect 55880 365 55885 370
rect 55845 360 55885 365
rect 56430 365 56435 370
rect 56465 390 56470 395
rect 56760 395 56800 400
rect 56760 390 56765 395
rect 56465 370 56765 390
rect 56465 365 56470 370
rect 56430 360 56470 365
rect 56760 365 56765 370
rect 56795 390 56800 395
rect 56880 395 56920 400
rect 56880 390 56885 395
rect 56795 370 56885 390
rect 56795 365 56800 370
rect 56760 360 56800 365
rect 56880 365 56885 370
rect 56915 390 56920 395
rect 57915 395 57955 400
rect 57915 390 57920 395
rect 56915 370 57920 390
rect 56915 365 56920 370
rect 56880 360 56920 365
rect 57915 365 57920 370
rect 57950 390 57955 395
rect 58180 395 58220 400
rect 58180 390 58185 395
rect 57950 370 58185 390
rect 57950 365 57955 370
rect 57915 360 57955 365
rect 58180 365 58185 370
rect 58215 390 58220 395
rect 58380 395 58420 400
rect 58380 390 58385 395
rect 58215 370 58385 390
rect 58215 365 58220 370
rect 58180 360 58220 365
rect 58380 365 58385 370
rect 58415 390 58420 395
rect 58580 395 58620 400
rect 58580 390 58585 395
rect 58415 370 58585 390
rect 58415 365 58420 370
rect 58380 360 58420 365
rect 58580 365 58585 370
rect 58615 390 58620 395
rect 58780 395 58820 400
rect 58780 390 58785 395
rect 58615 370 58785 390
rect 58615 365 58620 370
rect 58580 360 58620 365
rect 58780 365 58785 370
rect 58815 390 58820 395
rect 59515 395 59555 400
rect 59515 390 59520 395
rect 58815 370 59520 390
rect 58815 365 58820 370
rect 58780 360 58820 365
rect 59515 365 59520 370
rect 59550 365 59555 395
rect 59515 360 59555 365
rect 56880 -515 56920 -510
rect 56880 -545 56885 -515
rect 56915 -545 56920 -515
rect 56880 -550 56920 -545
<< via2 >>
rect 56885 6155 56915 6185
rect 54610 3370 54640 3400
rect 59160 3370 59190 3400
rect 54300 1880 54330 1910
rect 59470 1880 59500 1910
rect 56885 -545 56915 -515
<< metal3 >>
rect 56875 6190 56925 6195
rect 56875 6150 56880 6190
rect 56920 6150 56925 6190
rect 56875 6145 56925 6150
rect 52410 5770 52640 5855
rect 52760 5770 52990 5855
rect 53110 5770 53340 5855
rect 52410 5720 53340 5770
rect 52410 5625 52640 5720
rect 52760 5625 52990 5720
rect 53110 5625 53340 5720
rect 53460 5625 53690 5855
rect 53810 5625 54040 5855
rect 54160 5625 54390 5855
rect 54510 5625 54740 5855
rect 54860 5625 55090 5855
rect 55210 5625 55440 5855
rect 55560 5625 55790 5855
rect 55910 5625 56140 5855
rect 56260 5625 56490 5855
rect 56610 5625 56840 5855
rect 56960 5625 57190 5855
rect 57310 5625 57540 5855
rect 57660 5625 57890 5855
rect 58010 5625 58240 5855
rect 58360 5625 58590 5855
rect 58710 5625 58940 5855
rect 59060 5625 59290 5855
rect 59410 5625 59640 5855
rect 59760 5625 59990 5855
rect 60110 5625 60340 5855
rect 60460 5770 60690 5855
rect 60810 5770 61040 5855
rect 61160 5770 61390 5855
rect 60460 5720 61390 5770
rect 60460 5625 60690 5720
rect 60810 5625 61040 5720
rect 61160 5625 61390 5720
rect 53200 5505 53250 5625
rect 53550 5505 53600 5625
rect 53900 5505 53950 5625
rect 54250 5505 54300 5625
rect 54600 5505 54650 5625
rect 54950 5505 55000 5625
rect 55300 5505 55350 5625
rect 55650 5505 55700 5625
rect 56000 5505 56050 5625
rect 56350 5505 56400 5625
rect 56700 5505 56750 5625
rect 57050 5505 57100 5625
rect 57400 5505 57450 5625
rect 57750 5505 57800 5625
rect 58100 5505 58150 5625
rect 58450 5505 58500 5625
rect 58800 5505 58850 5625
rect 59150 5505 59200 5625
rect 59500 5505 59550 5625
rect 59850 5505 59900 5625
rect 60200 5505 60250 5625
rect 60550 5505 60600 5625
rect 52410 5420 52640 5505
rect 52760 5420 52990 5505
rect 53110 5420 53340 5505
rect 53460 5420 53690 5505
rect 53810 5420 54040 5505
rect 54160 5420 54390 5505
rect 54510 5420 54740 5505
rect 54860 5420 55090 5505
rect 55210 5420 55440 5505
rect 55560 5420 55790 5505
rect 55910 5420 56140 5505
rect 56260 5420 56490 5505
rect 56610 5420 56840 5505
rect 52410 5370 56840 5420
rect 52410 5275 52640 5370
rect 52760 5275 52990 5370
rect 53110 5275 53340 5370
rect 53460 5275 53690 5370
rect 53810 5275 54040 5370
rect 54160 5275 54390 5370
rect 54510 5275 54740 5370
rect 54860 5275 55090 5370
rect 55210 5275 55440 5370
rect 55560 5275 55790 5370
rect 55910 5275 56140 5370
rect 56260 5275 56490 5370
rect 56610 5275 56840 5370
rect 56960 5420 57190 5505
rect 57310 5420 57540 5505
rect 57660 5420 57890 5505
rect 58010 5420 58240 5505
rect 58360 5420 58590 5505
rect 58710 5420 58940 5505
rect 59060 5420 59290 5505
rect 59410 5420 59640 5505
rect 59760 5420 59990 5505
rect 60110 5420 60340 5505
rect 60460 5420 60690 5505
rect 60810 5420 61040 5505
rect 61160 5420 61390 5505
rect 56960 5370 61390 5420
rect 56960 5275 57190 5370
rect 57310 5275 57540 5370
rect 57660 5275 57890 5370
rect 58010 5275 58240 5370
rect 58360 5275 58590 5370
rect 58710 5275 58940 5370
rect 59060 5275 59290 5370
rect 59410 5275 59640 5370
rect 59760 5275 59990 5370
rect 60110 5275 60340 5370
rect 60460 5275 60690 5370
rect 60810 5275 61040 5370
rect 61160 5275 61390 5370
rect 53200 5155 53250 5275
rect 54250 5155 54300 5275
rect 54600 5155 54650 5275
rect 54950 5155 55000 5275
rect 55300 5155 55350 5275
rect 55650 5155 55700 5275
rect 56000 5155 56050 5275
rect 56350 5155 56400 5275
rect 56700 5155 56750 5275
rect 57050 5155 57100 5275
rect 57400 5155 57450 5275
rect 57750 5155 57800 5275
rect 58100 5155 58150 5275
rect 58450 5155 58500 5275
rect 58800 5155 58850 5275
rect 59150 5155 59200 5275
rect 59500 5155 59550 5275
rect 60550 5155 60600 5275
rect 52410 5070 52640 5155
rect 52760 5070 52990 5155
rect 53110 5070 53340 5155
rect 53460 5070 53690 5155
rect 53810 5070 54040 5155
rect 52410 5020 54040 5070
rect 52410 4925 52640 5020
rect 52760 4925 52990 5020
rect 53110 4925 53340 5020
rect 53460 4925 53690 5020
rect 53810 4925 54040 5020
rect 54160 4925 54390 5155
rect 54510 4925 54740 5155
rect 54860 4925 55090 5155
rect 55210 4925 55440 5155
rect 55560 4925 55790 5155
rect 55910 4925 56140 5155
rect 56260 4925 56490 5155
rect 56610 4925 56840 5155
rect 56960 4925 57190 5155
rect 57310 4925 57540 5155
rect 57660 4925 57890 5155
rect 58010 4925 58240 5155
rect 58360 4925 58590 5155
rect 58710 4925 58940 5155
rect 59060 4925 59290 5155
rect 59410 4925 59640 5155
rect 59760 5070 59990 5155
rect 60110 5070 60340 5155
rect 60460 5070 60690 5155
rect 60810 5070 61040 5155
rect 61160 5070 61390 5155
rect 59760 5020 61390 5070
rect 59760 4925 59990 5020
rect 60110 4925 60340 5020
rect 60460 4925 60690 5020
rect 60810 4925 61040 5020
rect 61160 4925 61390 5020
rect 53200 4805 53250 4925
rect 54250 4805 54300 4925
rect 54600 4805 54650 4925
rect 54950 4805 55000 4925
rect 55300 4805 55350 4925
rect 58450 4805 58500 4925
rect 58800 4805 58850 4925
rect 59150 4805 59200 4925
rect 59500 4805 59550 4925
rect 60550 4805 60600 4925
rect 52410 4720 52640 4805
rect 52760 4720 52990 4805
rect 53110 4720 53340 4805
rect 53460 4720 53690 4805
rect 53810 4720 54040 4805
rect 52410 4670 54040 4720
rect 52410 4575 52640 4670
rect 52760 4575 52990 4670
rect 53110 4575 53340 4670
rect 53460 4575 53690 4670
rect 53810 4575 54040 4670
rect 54160 4575 54390 4805
rect 54510 4575 54740 4805
rect 54860 4575 55090 4805
rect 55210 4575 55440 4805
rect 58360 4575 58590 4805
rect 58710 4575 58940 4805
rect 59060 4575 59290 4805
rect 59410 4575 59640 4805
rect 59760 4720 59990 4805
rect 60110 4720 60340 4805
rect 60460 4720 60690 4805
rect 60810 4720 61040 4805
rect 61160 4720 61390 4805
rect 59760 4670 61390 4720
rect 59760 4575 59990 4670
rect 60110 4575 60340 4670
rect 60460 4575 60690 4670
rect 60810 4575 61040 4670
rect 61160 4575 61390 4670
rect 53200 4455 53250 4575
rect 54250 4455 54300 4575
rect 54600 4455 54650 4575
rect 54950 4455 55000 4575
rect 55300 4455 55350 4575
rect 58450 4455 58500 4575
rect 58800 4455 58850 4575
rect 59150 4455 59200 4575
rect 59500 4455 59550 4575
rect 60550 4455 60600 4575
rect 52410 4370 52640 4455
rect 52760 4370 52990 4455
rect 53110 4370 53340 4455
rect 53460 4370 53690 4455
rect 53810 4370 54040 4455
rect 52410 4320 54040 4370
rect 52410 4225 52640 4320
rect 52760 4225 52990 4320
rect 53110 4225 53340 4320
rect 53460 4225 53690 4320
rect 53810 4225 54040 4320
rect 54160 4225 54390 4455
rect 54510 4225 54740 4455
rect 54860 4225 55090 4455
rect 55210 4225 55440 4455
rect 58360 4225 58590 4455
rect 58710 4225 58940 4455
rect 59060 4225 59290 4455
rect 59410 4225 59640 4455
rect 59760 4370 59990 4455
rect 60110 4370 60340 4455
rect 60460 4370 60690 4455
rect 60810 4370 61040 4455
rect 61160 4370 61390 4455
rect 59760 4320 61390 4370
rect 59760 4225 59990 4320
rect 60110 4225 60340 4320
rect 60460 4225 60690 4320
rect 60810 4225 61040 4320
rect 61160 4225 61390 4320
rect 53200 4105 53250 4225
rect 52410 4020 52640 4105
rect 52760 4020 52990 4105
rect 53110 4020 53340 4105
rect 53460 4020 53690 4105
rect 53810 4020 54040 4105
rect 52410 3970 54040 4020
rect 52410 3875 52640 3970
rect 52760 3875 52990 3970
rect 53110 3875 53340 3970
rect 53460 3875 53690 3970
rect 53810 3875 54040 3970
rect 53200 3755 53250 3875
rect 52410 3670 52640 3755
rect 52760 3670 52990 3755
rect 53110 3670 53340 3755
rect 53460 3670 53690 3755
rect 53810 3670 54040 3755
rect 52410 3620 54040 3670
rect 52410 3525 52640 3620
rect 52760 3525 52990 3620
rect 53110 3525 53340 3620
rect 53460 3525 53690 3620
rect 53810 3525 54040 3620
rect 53200 3405 53250 3525
rect 52410 3320 52640 3405
rect 52760 3320 52990 3405
rect 53110 3320 53340 3405
rect 53460 3320 53690 3405
rect 53810 3320 54040 3405
rect 54605 3400 54645 4225
rect 54605 3370 54610 3400
rect 54640 3370 54645 3400
rect 54605 3365 54645 3370
rect 59155 3400 59195 4225
rect 60550 4105 60600 4225
rect 59760 4020 59990 4105
rect 60110 4020 60340 4105
rect 60460 4020 60690 4105
rect 60810 4020 61040 4105
rect 61160 4020 61390 4105
rect 59760 3970 61390 4020
rect 59760 3875 59990 3970
rect 60110 3875 60340 3970
rect 60460 3875 60690 3970
rect 60810 3875 61040 3970
rect 61160 3875 61390 3970
rect 60550 3755 60600 3875
rect 59760 3670 59990 3755
rect 60110 3670 60340 3755
rect 60460 3670 60690 3755
rect 60810 3670 61040 3755
rect 61160 3670 61390 3755
rect 59760 3620 61390 3670
rect 59760 3525 59990 3620
rect 60110 3525 60340 3620
rect 60460 3525 60690 3620
rect 60810 3525 61040 3620
rect 61160 3525 61390 3620
rect 60550 3405 60600 3525
rect 59155 3370 59160 3400
rect 59190 3370 59195 3400
rect 59155 3365 59195 3370
rect 52410 3270 54040 3320
rect 52410 3175 52640 3270
rect 52760 3175 52990 3270
rect 53110 3175 53340 3270
rect 53460 3175 53690 3270
rect 53810 3175 54040 3270
rect 59760 3320 59990 3405
rect 60110 3320 60340 3405
rect 60460 3320 60690 3405
rect 60810 3320 61040 3405
rect 61160 3320 61390 3405
rect 59760 3270 61390 3320
rect 59760 3175 59990 3270
rect 60110 3175 60340 3270
rect 60460 3175 60690 3270
rect 60810 3175 61040 3270
rect 61160 3175 61390 3270
rect 53200 3055 53250 3175
rect 60550 3055 60600 3175
rect 52410 2970 52640 3055
rect 52760 2970 52990 3055
rect 53110 2970 53340 3055
rect 53460 2970 53690 3055
rect 53810 2970 54040 3055
rect 52410 2920 54040 2970
rect 52410 2825 52640 2920
rect 52760 2825 52990 2920
rect 53110 2825 53340 2920
rect 53460 2825 53690 2920
rect 53810 2825 54040 2920
rect 59760 2970 59990 3055
rect 60110 2970 60340 3055
rect 60460 2970 60690 3055
rect 60810 2970 61040 3055
rect 61160 2970 61390 3055
rect 59760 2920 61390 2970
rect 59760 2825 59990 2920
rect 60110 2825 60340 2920
rect 60460 2825 60690 2920
rect 60810 2825 61040 2920
rect 61160 2825 61390 2920
rect 53200 2705 53250 2825
rect 60550 2705 60600 2825
rect 52410 2620 52640 2705
rect 52760 2620 52990 2705
rect 53110 2620 53340 2705
rect 53460 2620 53690 2705
rect 53810 2620 54040 2705
rect 52410 2570 54040 2620
rect 52410 2475 52640 2570
rect 52760 2475 52990 2570
rect 53110 2475 53340 2570
rect 53460 2475 53690 2570
rect 53810 2475 54040 2570
rect 59760 2620 59990 2705
rect 60110 2620 60340 2705
rect 60460 2620 60690 2705
rect 60810 2620 61040 2705
rect 61160 2620 61390 2705
rect 59760 2570 61390 2620
rect 59760 2475 59990 2570
rect 60110 2475 60340 2570
rect 60460 2475 60690 2570
rect 60810 2475 61040 2570
rect 61160 2475 61390 2570
rect 53200 2355 53250 2475
rect 60550 2355 60600 2475
rect 52410 2270 52640 2355
rect 52760 2270 52990 2355
rect 53110 2270 53340 2355
rect 53460 2270 53690 2355
rect 53810 2270 54040 2355
rect 52410 2220 54040 2270
rect 52410 2125 52640 2220
rect 52760 2125 52990 2220
rect 53110 2125 53340 2220
rect 53460 2125 53690 2220
rect 53810 2125 54040 2220
rect 59760 2270 59990 2355
rect 60110 2270 60340 2355
rect 60460 2270 60690 2355
rect 60810 2270 61040 2355
rect 61160 2270 61390 2355
rect 59760 2220 61390 2270
rect 59760 2125 59990 2220
rect 60110 2125 60340 2220
rect 60460 2125 60690 2220
rect 60810 2125 61040 2220
rect 61160 2125 61390 2220
rect 53200 2005 53250 2125
rect 60550 2005 60600 2125
rect 52410 1920 52640 2005
rect 52760 1920 52990 2005
rect 53110 1920 53340 2005
rect 53460 1920 53690 2005
rect 53810 1920 54040 2005
rect 59760 1920 59990 2005
rect 60110 1920 60340 2005
rect 60460 1920 60690 2005
rect 60810 1920 61040 2005
rect 61160 1920 61390 2005
rect 52410 1870 54040 1920
rect 54290 1915 54340 1920
rect 54290 1875 54295 1915
rect 54335 1875 54340 1915
rect 54290 1870 54340 1875
rect 59460 1915 59510 1920
rect 59460 1875 59465 1915
rect 59505 1875 59510 1915
rect 59460 1870 59510 1875
rect 59760 1870 61390 1920
rect 52410 1775 52640 1870
rect 52760 1775 52990 1870
rect 53110 1775 53340 1870
rect 53460 1775 53690 1870
rect 53810 1775 54040 1870
rect 59760 1775 59990 1870
rect 60110 1775 60340 1870
rect 60460 1775 60690 1870
rect 60810 1775 61040 1870
rect 61160 1775 61390 1870
rect 53200 1655 53250 1775
rect 60550 1655 60600 1775
rect 52410 1570 52640 1655
rect 52760 1570 52990 1655
rect 53110 1570 53340 1655
rect 53460 1570 53690 1655
rect 53810 1570 54040 1655
rect 52410 1520 54040 1570
rect 52410 1425 52640 1520
rect 52760 1425 52990 1520
rect 53110 1425 53340 1520
rect 53460 1425 53690 1520
rect 53810 1425 54040 1520
rect 59760 1570 59990 1655
rect 60110 1570 60340 1655
rect 60460 1570 60690 1655
rect 60810 1570 61040 1655
rect 61160 1570 61390 1655
rect 59760 1520 61390 1570
rect 59760 1425 59990 1520
rect 60110 1425 60340 1520
rect 60460 1425 60690 1520
rect 60810 1425 61040 1520
rect 61160 1425 61390 1520
rect 53200 1305 53250 1425
rect 60550 1305 60600 1425
rect 52410 1220 52640 1305
rect 52760 1220 52990 1305
rect 53110 1220 53340 1305
rect 53460 1220 53690 1305
rect 53810 1220 54040 1305
rect 52410 1170 54040 1220
rect 52410 1075 52640 1170
rect 52760 1075 52990 1170
rect 53110 1075 53340 1170
rect 53460 1075 53690 1170
rect 53810 1075 54040 1170
rect 59760 1220 59990 1305
rect 60110 1220 60340 1305
rect 60460 1220 60690 1305
rect 60810 1220 61040 1305
rect 61160 1220 61390 1305
rect 59760 1170 61390 1220
rect 59760 1075 59990 1170
rect 60110 1075 60340 1170
rect 60460 1075 60690 1170
rect 60810 1075 61040 1170
rect 61160 1075 61390 1170
rect 53200 955 53250 1075
rect 60550 955 60600 1075
rect 52410 870 52640 955
rect 52760 870 52990 955
rect 53110 870 53340 955
rect 53460 870 53690 955
rect 53810 870 54040 955
rect 52410 820 54040 870
rect 52410 725 52640 820
rect 52760 725 52990 820
rect 53110 725 53340 820
rect 53460 725 53690 820
rect 53810 725 54040 820
rect 59760 870 59990 955
rect 60110 870 60340 955
rect 60460 870 60690 955
rect 60810 870 61040 955
rect 61160 870 61390 955
rect 59760 820 61390 870
rect 59760 725 59990 820
rect 60110 725 60340 820
rect 60460 725 60690 820
rect 60810 725 61040 820
rect 61160 725 61390 820
rect 53200 605 53250 725
rect 60550 605 60600 725
rect 52410 520 52640 605
rect 52760 520 52990 605
rect 53110 520 53340 605
rect 53460 520 53690 605
rect 53810 520 54040 605
rect 52410 470 54040 520
rect 52410 375 52640 470
rect 52760 375 52990 470
rect 53110 375 53340 470
rect 53460 375 53690 470
rect 53810 375 54040 470
rect 59760 520 59990 605
rect 60110 520 60340 605
rect 60460 520 60690 605
rect 60810 520 61040 605
rect 61160 520 61390 605
rect 59760 470 61390 520
rect 59760 375 59990 470
rect 60110 375 60340 470
rect 60460 375 60690 470
rect 60810 375 61040 470
rect 61160 375 61390 470
rect 53200 255 53250 375
rect 60550 255 60600 375
rect 52410 170 52640 255
rect 52760 170 52990 255
rect 53110 170 53340 255
rect 53460 170 53690 255
rect 53810 170 54040 255
rect 54160 170 54390 255
rect 54510 170 54740 255
rect 54860 170 55090 255
rect 55210 170 55440 255
rect 55560 170 55790 255
rect 55910 170 56140 255
rect 56260 170 56490 255
rect 56610 170 56840 255
rect 52410 120 56840 170
rect 52410 25 52640 120
rect 52760 25 52990 120
rect 53110 25 53340 120
rect 53460 25 53690 120
rect 53810 25 54040 120
rect 54160 25 54390 120
rect 54510 25 54740 120
rect 54860 25 55090 120
rect 55210 25 55440 120
rect 55560 25 55790 120
rect 55910 25 56140 120
rect 56260 25 56490 120
rect 56610 25 56840 120
rect 56960 170 57190 255
rect 57310 170 57540 255
rect 57660 170 57890 255
rect 58010 170 58240 255
rect 58360 170 58590 255
rect 58710 170 58940 255
rect 59060 170 59290 255
rect 59410 170 59640 255
rect 59760 170 59990 255
rect 60110 170 60340 255
rect 60460 170 60690 255
rect 60810 170 61040 255
rect 61160 170 61390 255
rect 56960 120 61390 170
rect 56960 25 57190 120
rect 57310 25 57540 120
rect 57660 25 57890 120
rect 58010 25 58240 120
rect 58360 25 58590 120
rect 58710 25 58940 120
rect 59060 25 59290 120
rect 59410 25 59640 120
rect 59760 25 59990 120
rect 60110 25 60340 120
rect 60460 25 60690 120
rect 60810 25 61040 120
rect 61160 25 61390 120
rect 53200 -95 53250 25
rect 53550 -95 53600 25
rect 53900 -95 53950 25
rect 54250 -95 54300 25
rect 54600 -95 54650 25
rect 54950 -95 55000 25
rect 55300 -95 55350 25
rect 55650 -95 55700 25
rect 56000 -95 56050 25
rect 56350 -95 56400 25
rect 56700 -95 56750 25
rect 57050 -95 57100 25
rect 57400 -95 57450 25
rect 57750 -95 57800 25
rect 58100 -95 58150 25
rect 58450 -95 58500 25
rect 58800 -95 58850 25
rect 59150 -95 59200 25
rect 59500 -95 59550 25
rect 59850 -95 59900 25
rect 60200 -95 60250 25
rect 60550 -95 60600 25
rect 52410 -180 52640 -95
rect 52760 -180 52990 -95
rect 53110 -180 53340 -95
rect 52410 -230 53340 -180
rect 52410 -325 52640 -230
rect 52760 -325 52990 -230
rect 53110 -325 53340 -230
rect 53460 -325 53690 -95
rect 53810 -325 54040 -95
rect 54160 -325 54390 -95
rect 54510 -325 54740 -95
rect 54860 -325 55090 -95
rect 55210 -325 55440 -95
rect 55560 -325 55790 -95
rect 55910 -325 56140 -95
rect 56260 -325 56490 -95
rect 56610 -325 56840 -95
rect 56960 -325 57190 -95
rect 57310 -325 57540 -95
rect 57660 -325 57890 -95
rect 58010 -325 58240 -95
rect 58360 -325 58590 -95
rect 58710 -325 58940 -95
rect 59060 -325 59290 -95
rect 59410 -325 59640 -95
rect 59760 -325 59990 -95
rect 60110 -325 60340 -95
rect 60460 -180 60690 -95
rect 60810 -180 61040 -95
rect 61160 -180 61390 -95
rect 60460 -230 61390 -180
rect 60460 -325 60690 -230
rect 60810 -325 61040 -230
rect 61160 -325 61390 -230
rect 56875 -510 56925 -505
rect 56875 -550 56880 -510
rect 56920 -550 56925 -510
rect 56875 -555 56925 -550
<< via3 >>
rect 56880 6185 56920 6190
rect 56880 6155 56885 6185
rect 56885 6155 56915 6185
rect 56915 6155 56920 6185
rect 56880 6150 56920 6155
rect 54295 1910 54335 1915
rect 54295 1880 54300 1910
rect 54300 1880 54330 1910
rect 54330 1880 54335 1910
rect 54295 1875 54335 1880
rect 59465 1910 59505 1915
rect 59465 1880 59470 1910
rect 59470 1880 59500 1910
rect 59500 1880 59505 1910
rect 59465 1875 59505 1880
rect 56880 -515 56920 -510
rect 56880 -545 56885 -515
rect 56885 -545 56915 -515
rect 56915 -545 56920 -515
rect 56880 -550 56920 -545
<< mimcap >>
rect 52425 5765 52625 5840
rect 52425 5725 52505 5765
rect 52545 5725 52625 5765
rect 52425 5640 52625 5725
rect 52775 5765 52975 5840
rect 52775 5725 52855 5765
rect 52895 5725 52975 5765
rect 52775 5640 52975 5725
rect 53125 5765 53325 5840
rect 53125 5725 53205 5765
rect 53245 5725 53325 5765
rect 53125 5640 53325 5725
rect 53475 5765 53675 5840
rect 53475 5725 53555 5765
rect 53595 5725 53675 5765
rect 53475 5640 53675 5725
rect 53825 5765 54025 5840
rect 53825 5725 53905 5765
rect 53945 5725 54025 5765
rect 53825 5640 54025 5725
rect 54175 5765 54375 5840
rect 54175 5725 54255 5765
rect 54295 5725 54375 5765
rect 54175 5640 54375 5725
rect 54525 5765 54725 5840
rect 54525 5725 54605 5765
rect 54645 5725 54725 5765
rect 54525 5640 54725 5725
rect 54875 5765 55075 5840
rect 54875 5725 54955 5765
rect 54995 5725 55075 5765
rect 54875 5640 55075 5725
rect 55225 5765 55425 5840
rect 55225 5725 55305 5765
rect 55345 5725 55425 5765
rect 55225 5640 55425 5725
rect 55575 5765 55775 5840
rect 55575 5725 55655 5765
rect 55695 5725 55775 5765
rect 55575 5640 55775 5725
rect 55925 5765 56125 5840
rect 55925 5725 56005 5765
rect 56045 5725 56125 5765
rect 55925 5640 56125 5725
rect 56275 5765 56475 5840
rect 56275 5725 56355 5765
rect 56395 5725 56475 5765
rect 56275 5640 56475 5725
rect 56625 5765 56825 5840
rect 56625 5725 56705 5765
rect 56745 5725 56825 5765
rect 56625 5640 56825 5725
rect 56975 5765 57175 5840
rect 56975 5725 57055 5765
rect 57095 5725 57175 5765
rect 56975 5640 57175 5725
rect 57325 5765 57525 5840
rect 57325 5725 57405 5765
rect 57445 5725 57525 5765
rect 57325 5640 57525 5725
rect 57675 5765 57875 5840
rect 57675 5725 57755 5765
rect 57795 5725 57875 5765
rect 57675 5640 57875 5725
rect 58025 5765 58225 5840
rect 58025 5725 58105 5765
rect 58145 5725 58225 5765
rect 58025 5640 58225 5725
rect 58375 5765 58575 5840
rect 58375 5725 58455 5765
rect 58495 5725 58575 5765
rect 58375 5640 58575 5725
rect 58725 5765 58925 5840
rect 58725 5725 58805 5765
rect 58845 5725 58925 5765
rect 58725 5640 58925 5725
rect 59075 5765 59275 5840
rect 59075 5725 59155 5765
rect 59195 5725 59275 5765
rect 59075 5640 59275 5725
rect 59425 5765 59625 5840
rect 59425 5725 59505 5765
rect 59545 5725 59625 5765
rect 59425 5640 59625 5725
rect 59775 5765 59975 5840
rect 59775 5725 59855 5765
rect 59895 5725 59975 5765
rect 59775 5640 59975 5725
rect 60125 5765 60325 5840
rect 60125 5725 60205 5765
rect 60245 5725 60325 5765
rect 60125 5640 60325 5725
rect 60475 5765 60675 5840
rect 60475 5725 60555 5765
rect 60595 5725 60675 5765
rect 60475 5640 60675 5725
rect 60825 5765 61025 5840
rect 60825 5725 60905 5765
rect 60945 5725 61025 5765
rect 60825 5640 61025 5725
rect 61175 5765 61375 5840
rect 61175 5725 61255 5765
rect 61295 5725 61375 5765
rect 61175 5640 61375 5725
rect 52425 5415 52625 5490
rect 52425 5375 52505 5415
rect 52545 5375 52625 5415
rect 52425 5290 52625 5375
rect 52775 5415 52975 5490
rect 52775 5375 52855 5415
rect 52895 5375 52975 5415
rect 52775 5290 52975 5375
rect 53125 5415 53325 5490
rect 53125 5375 53205 5415
rect 53245 5375 53325 5415
rect 53125 5290 53325 5375
rect 53475 5415 53675 5490
rect 53475 5375 53555 5415
rect 53595 5375 53675 5415
rect 53475 5290 53675 5375
rect 53825 5415 54025 5490
rect 53825 5375 53905 5415
rect 53945 5375 54025 5415
rect 53825 5290 54025 5375
rect 54175 5415 54375 5490
rect 54175 5375 54255 5415
rect 54295 5375 54375 5415
rect 54175 5290 54375 5375
rect 54525 5415 54725 5490
rect 54525 5375 54605 5415
rect 54645 5375 54725 5415
rect 54525 5290 54725 5375
rect 54875 5415 55075 5490
rect 54875 5375 54955 5415
rect 54995 5375 55075 5415
rect 54875 5290 55075 5375
rect 55225 5415 55425 5490
rect 55225 5375 55305 5415
rect 55345 5375 55425 5415
rect 55225 5290 55425 5375
rect 55575 5415 55775 5490
rect 55575 5375 55655 5415
rect 55695 5375 55775 5415
rect 55575 5290 55775 5375
rect 55925 5415 56125 5490
rect 55925 5375 56005 5415
rect 56045 5375 56125 5415
rect 55925 5290 56125 5375
rect 56275 5415 56475 5490
rect 56275 5375 56355 5415
rect 56395 5375 56475 5415
rect 56275 5290 56475 5375
rect 56625 5415 56825 5490
rect 56625 5375 56705 5415
rect 56745 5375 56825 5415
rect 56625 5290 56825 5375
rect 56975 5415 57175 5490
rect 56975 5375 57055 5415
rect 57095 5375 57175 5415
rect 56975 5290 57175 5375
rect 57325 5415 57525 5490
rect 57325 5375 57405 5415
rect 57445 5375 57525 5415
rect 57325 5290 57525 5375
rect 57675 5415 57875 5490
rect 57675 5375 57755 5415
rect 57795 5375 57875 5415
rect 57675 5290 57875 5375
rect 58025 5415 58225 5490
rect 58025 5375 58105 5415
rect 58145 5375 58225 5415
rect 58025 5290 58225 5375
rect 58375 5415 58575 5490
rect 58375 5375 58455 5415
rect 58495 5375 58575 5415
rect 58375 5290 58575 5375
rect 58725 5415 58925 5490
rect 58725 5375 58805 5415
rect 58845 5375 58925 5415
rect 58725 5290 58925 5375
rect 59075 5415 59275 5490
rect 59075 5375 59155 5415
rect 59195 5375 59275 5415
rect 59075 5290 59275 5375
rect 59425 5415 59625 5490
rect 59425 5375 59505 5415
rect 59545 5375 59625 5415
rect 59425 5290 59625 5375
rect 59775 5415 59975 5490
rect 59775 5375 59855 5415
rect 59895 5375 59975 5415
rect 59775 5290 59975 5375
rect 60125 5415 60325 5490
rect 60125 5375 60205 5415
rect 60245 5375 60325 5415
rect 60125 5290 60325 5375
rect 60475 5415 60675 5490
rect 60475 5375 60555 5415
rect 60595 5375 60675 5415
rect 60475 5290 60675 5375
rect 60825 5415 61025 5490
rect 60825 5375 60905 5415
rect 60945 5375 61025 5415
rect 60825 5290 61025 5375
rect 61175 5415 61375 5490
rect 61175 5375 61255 5415
rect 61295 5375 61375 5415
rect 61175 5290 61375 5375
rect 52425 5065 52625 5140
rect 52425 5025 52505 5065
rect 52545 5025 52625 5065
rect 52425 4940 52625 5025
rect 52775 5065 52975 5140
rect 52775 5025 52855 5065
rect 52895 5025 52975 5065
rect 52775 4940 52975 5025
rect 53125 5065 53325 5140
rect 53125 5025 53205 5065
rect 53245 5025 53325 5065
rect 53125 4940 53325 5025
rect 53475 5065 53675 5140
rect 53475 5025 53555 5065
rect 53595 5025 53675 5065
rect 53475 4940 53675 5025
rect 53825 5065 54025 5140
rect 53825 5025 53905 5065
rect 53945 5025 54025 5065
rect 53825 4940 54025 5025
rect 54175 5065 54375 5140
rect 54175 5025 54255 5065
rect 54295 5025 54375 5065
rect 54175 4940 54375 5025
rect 54525 5065 54725 5140
rect 54525 5025 54605 5065
rect 54645 5025 54725 5065
rect 54525 4940 54725 5025
rect 54875 5065 55075 5140
rect 54875 5025 54955 5065
rect 54995 5025 55075 5065
rect 54875 4940 55075 5025
rect 55225 5065 55425 5140
rect 55225 5025 55305 5065
rect 55345 5025 55425 5065
rect 55225 4940 55425 5025
rect 55575 5055 55775 5140
rect 55575 5015 55655 5055
rect 55695 5015 55775 5055
rect 55575 4940 55775 5015
rect 55925 5055 56125 5140
rect 55925 5015 56005 5055
rect 56045 5015 56125 5055
rect 55925 4940 56125 5015
rect 56275 5055 56475 5140
rect 56275 5015 56355 5055
rect 56395 5015 56475 5055
rect 56275 4940 56475 5015
rect 56625 5055 56825 5140
rect 56625 5015 56705 5055
rect 56745 5015 56825 5055
rect 56625 4940 56825 5015
rect 56975 5055 57175 5140
rect 56975 5015 57055 5055
rect 57095 5015 57175 5055
rect 56975 4940 57175 5015
rect 57325 5055 57525 5140
rect 57325 5015 57405 5055
rect 57445 5015 57525 5055
rect 57325 4940 57525 5015
rect 57675 5055 57875 5140
rect 57675 5015 57755 5055
rect 57795 5015 57875 5055
rect 57675 4940 57875 5015
rect 58025 5055 58225 5140
rect 58025 5015 58105 5055
rect 58145 5015 58225 5055
rect 58025 4940 58225 5015
rect 58375 5065 58575 5140
rect 58375 5025 58455 5065
rect 58495 5025 58575 5065
rect 58375 4940 58575 5025
rect 58725 5065 58925 5140
rect 58725 5025 58805 5065
rect 58845 5025 58925 5065
rect 58725 4940 58925 5025
rect 59075 5065 59275 5140
rect 59075 5025 59155 5065
rect 59195 5025 59275 5065
rect 59075 4940 59275 5025
rect 59425 5065 59625 5140
rect 59425 5025 59505 5065
rect 59545 5025 59625 5065
rect 59425 4940 59625 5025
rect 59775 5065 59975 5140
rect 59775 5025 59855 5065
rect 59895 5025 59975 5065
rect 59775 4940 59975 5025
rect 60125 5065 60325 5140
rect 60125 5025 60205 5065
rect 60245 5025 60325 5065
rect 60125 4940 60325 5025
rect 60475 5065 60675 5140
rect 60475 5025 60555 5065
rect 60595 5025 60675 5065
rect 60475 4940 60675 5025
rect 60825 5065 61025 5140
rect 60825 5025 60905 5065
rect 60945 5025 61025 5065
rect 60825 4940 61025 5025
rect 61175 5065 61375 5140
rect 61175 5025 61255 5065
rect 61295 5025 61375 5065
rect 61175 4940 61375 5025
rect 52425 4715 52625 4790
rect 52425 4675 52505 4715
rect 52545 4675 52625 4715
rect 52425 4590 52625 4675
rect 52775 4715 52975 4790
rect 52775 4675 52855 4715
rect 52895 4675 52975 4715
rect 52775 4590 52975 4675
rect 53125 4715 53325 4790
rect 53125 4675 53205 4715
rect 53245 4675 53325 4715
rect 53125 4590 53325 4675
rect 53475 4715 53675 4790
rect 53475 4675 53555 4715
rect 53595 4675 53675 4715
rect 53475 4590 53675 4675
rect 53825 4715 54025 4790
rect 53825 4675 53905 4715
rect 53945 4675 54025 4715
rect 53825 4590 54025 4675
rect 54175 4715 54375 4790
rect 54175 4675 54255 4715
rect 54295 4675 54375 4715
rect 54175 4590 54375 4675
rect 54525 4715 54725 4790
rect 54525 4675 54605 4715
rect 54645 4675 54725 4715
rect 54525 4590 54725 4675
rect 54875 4715 55075 4790
rect 54875 4675 54955 4715
rect 54995 4675 55075 4715
rect 54875 4590 55075 4675
rect 55225 4715 55425 4790
rect 55225 4675 55305 4715
rect 55345 4675 55425 4715
rect 55225 4590 55425 4675
rect 58375 4715 58575 4790
rect 58375 4675 58455 4715
rect 58495 4675 58575 4715
rect 58375 4590 58575 4675
rect 58725 4715 58925 4790
rect 58725 4675 58805 4715
rect 58845 4675 58925 4715
rect 58725 4590 58925 4675
rect 59075 4715 59275 4790
rect 59075 4675 59155 4715
rect 59195 4675 59275 4715
rect 59075 4590 59275 4675
rect 59425 4715 59625 4790
rect 59425 4675 59505 4715
rect 59545 4675 59625 4715
rect 59425 4590 59625 4675
rect 59775 4715 59975 4790
rect 59775 4675 59855 4715
rect 59895 4675 59975 4715
rect 59775 4590 59975 4675
rect 60125 4715 60325 4790
rect 60125 4675 60205 4715
rect 60245 4675 60325 4715
rect 60125 4590 60325 4675
rect 60475 4715 60675 4790
rect 60475 4675 60555 4715
rect 60595 4675 60675 4715
rect 60475 4590 60675 4675
rect 60825 4715 61025 4790
rect 60825 4675 60905 4715
rect 60945 4675 61025 4715
rect 60825 4590 61025 4675
rect 61175 4715 61375 4790
rect 61175 4675 61255 4715
rect 61295 4675 61375 4715
rect 61175 4590 61375 4675
rect 52425 4365 52625 4440
rect 52425 4325 52505 4365
rect 52545 4325 52625 4365
rect 52425 4240 52625 4325
rect 52775 4365 52975 4440
rect 52775 4325 52855 4365
rect 52895 4325 52975 4365
rect 52775 4240 52975 4325
rect 53125 4365 53325 4440
rect 53125 4325 53205 4365
rect 53245 4325 53325 4365
rect 53125 4240 53325 4325
rect 53475 4365 53675 4440
rect 53475 4325 53555 4365
rect 53595 4325 53675 4365
rect 53475 4240 53675 4325
rect 53825 4365 54025 4440
rect 53825 4325 53905 4365
rect 53945 4325 54025 4365
rect 53825 4240 54025 4325
rect 54175 4365 54375 4440
rect 54175 4325 54255 4365
rect 54295 4325 54375 4365
rect 54175 4240 54375 4325
rect 54525 4365 54725 4440
rect 54525 4325 54605 4365
rect 54645 4325 54725 4365
rect 54525 4240 54725 4325
rect 54875 4365 55075 4440
rect 54875 4325 54955 4365
rect 54995 4325 55075 4365
rect 54875 4240 55075 4325
rect 55225 4365 55425 4440
rect 55225 4325 55305 4365
rect 55345 4325 55425 4365
rect 55225 4240 55425 4325
rect 58375 4365 58575 4440
rect 58375 4325 58455 4365
rect 58495 4325 58575 4365
rect 58375 4240 58575 4325
rect 58725 4365 58925 4440
rect 58725 4325 58805 4365
rect 58845 4325 58925 4365
rect 58725 4240 58925 4325
rect 59075 4365 59275 4440
rect 59075 4325 59155 4365
rect 59195 4325 59275 4365
rect 59075 4240 59275 4325
rect 59425 4365 59625 4440
rect 59425 4325 59505 4365
rect 59545 4325 59625 4365
rect 59425 4240 59625 4325
rect 59775 4365 59975 4440
rect 59775 4325 59855 4365
rect 59895 4325 59975 4365
rect 59775 4240 59975 4325
rect 60125 4365 60325 4440
rect 60125 4325 60205 4365
rect 60245 4325 60325 4365
rect 60125 4240 60325 4325
rect 60475 4365 60675 4440
rect 60475 4325 60555 4365
rect 60595 4325 60675 4365
rect 60475 4240 60675 4325
rect 60825 4365 61025 4440
rect 60825 4325 60905 4365
rect 60945 4325 61025 4365
rect 60825 4240 61025 4325
rect 61175 4365 61375 4440
rect 61175 4325 61255 4365
rect 61295 4325 61375 4365
rect 61175 4240 61375 4325
rect 52425 4015 52625 4090
rect 52425 3975 52505 4015
rect 52545 3975 52625 4015
rect 52425 3890 52625 3975
rect 52775 4015 52975 4090
rect 52775 3975 52855 4015
rect 52895 3975 52975 4015
rect 52775 3890 52975 3975
rect 53125 4015 53325 4090
rect 53125 3975 53205 4015
rect 53245 3975 53325 4015
rect 53125 3890 53325 3975
rect 53475 4015 53675 4090
rect 53475 3975 53555 4015
rect 53595 3975 53675 4015
rect 53475 3890 53675 3975
rect 53825 4015 54025 4090
rect 53825 3975 53905 4015
rect 53945 3975 54025 4015
rect 53825 3890 54025 3975
rect 59775 4015 59975 4090
rect 59775 3975 59855 4015
rect 59895 3975 59975 4015
rect 59775 3890 59975 3975
rect 60125 4015 60325 4090
rect 60125 3975 60205 4015
rect 60245 3975 60325 4015
rect 60125 3890 60325 3975
rect 60475 4015 60675 4090
rect 60475 3975 60555 4015
rect 60595 3975 60675 4015
rect 60475 3890 60675 3975
rect 60825 4015 61025 4090
rect 60825 3975 60905 4015
rect 60945 3975 61025 4015
rect 60825 3890 61025 3975
rect 61175 4015 61375 4090
rect 61175 3975 61255 4015
rect 61295 3975 61375 4015
rect 61175 3890 61375 3975
rect 52425 3665 52625 3740
rect 52425 3625 52505 3665
rect 52545 3625 52625 3665
rect 52425 3540 52625 3625
rect 52775 3665 52975 3740
rect 52775 3625 52855 3665
rect 52895 3625 52975 3665
rect 52775 3540 52975 3625
rect 53125 3665 53325 3740
rect 53125 3625 53205 3665
rect 53245 3625 53325 3665
rect 53125 3540 53325 3625
rect 53475 3665 53675 3740
rect 53475 3625 53555 3665
rect 53595 3625 53675 3665
rect 53475 3540 53675 3625
rect 53825 3665 54025 3740
rect 53825 3625 53905 3665
rect 53945 3625 54025 3665
rect 53825 3540 54025 3625
rect 59775 3665 59975 3740
rect 59775 3625 59855 3665
rect 59895 3625 59975 3665
rect 59775 3540 59975 3625
rect 60125 3665 60325 3740
rect 60125 3625 60205 3665
rect 60245 3625 60325 3665
rect 60125 3540 60325 3625
rect 60475 3665 60675 3740
rect 60475 3625 60555 3665
rect 60595 3625 60675 3665
rect 60475 3540 60675 3625
rect 60825 3665 61025 3740
rect 60825 3625 60905 3665
rect 60945 3625 61025 3665
rect 60825 3540 61025 3625
rect 61175 3665 61375 3740
rect 61175 3625 61255 3665
rect 61295 3625 61375 3665
rect 61175 3540 61375 3625
rect 52425 3315 52625 3390
rect 52425 3275 52505 3315
rect 52545 3275 52625 3315
rect 52425 3190 52625 3275
rect 52775 3315 52975 3390
rect 52775 3275 52855 3315
rect 52895 3275 52975 3315
rect 52775 3190 52975 3275
rect 53125 3315 53325 3390
rect 53125 3275 53205 3315
rect 53245 3275 53325 3315
rect 53125 3190 53325 3275
rect 53475 3315 53675 3390
rect 53475 3275 53555 3315
rect 53595 3275 53675 3315
rect 53475 3190 53675 3275
rect 53825 3315 54025 3390
rect 53825 3275 53905 3315
rect 53945 3275 54025 3315
rect 53825 3190 54025 3275
rect 59775 3315 59975 3390
rect 59775 3275 59855 3315
rect 59895 3275 59975 3315
rect 59775 3190 59975 3275
rect 60125 3315 60325 3390
rect 60125 3275 60205 3315
rect 60245 3275 60325 3315
rect 60125 3190 60325 3275
rect 60475 3315 60675 3390
rect 60475 3275 60555 3315
rect 60595 3275 60675 3315
rect 60475 3190 60675 3275
rect 60825 3315 61025 3390
rect 60825 3275 60905 3315
rect 60945 3275 61025 3315
rect 60825 3190 61025 3275
rect 61175 3315 61375 3390
rect 61175 3275 61255 3315
rect 61295 3275 61375 3315
rect 61175 3190 61375 3275
rect 52425 2965 52625 3040
rect 52425 2925 52505 2965
rect 52545 2925 52625 2965
rect 52425 2840 52625 2925
rect 52775 2965 52975 3040
rect 52775 2925 52855 2965
rect 52895 2925 52975 2965
rect 52775 2840 52975 2925
rect 53125 2965 53325 3040
rect 53125 2925 53205 2965
rect 53245 2925 53325 2965
rect 53125 2840 53325 2925
rect 53475 2965 53675 3040
rect 53475 2925 53555 2965
rect 53595 2925 53675 2965
rect 53475 2840 53675 2925
rect 53825 2965 54025 3040
rect 53825 2925 53905 2965
rect 53945 2925 54025 2965
rect 53825 2840 54025 2925
rect 59775 2965 59975 3040
rect 59775 2925 59855 2965
rect 59895 2925 59975 2965
rect 59775 2840 59975 2925
rect 60125 2965 60325 3040
rect 60125 2925 60205 2965
rect 60245 2925 60325 2965
rect 60125 2840 60325 2925
rect 60475 2965 60675 3040
rect 60475 2925 60555 2965
rect 60595 2925 60675 2965
rect 60475 2840 60675 2925
rect 60825 2965 61025 3040
rect 60825 2925 60905 2965
rect 60945 2925 61025 2965
rect 60825 2840 61025 2925
rect 61175 2965 61375 3040
rect 61175 2925 61255 2965
rect 61295 2925 61375 2965
rect 61175 2840 61375 2925
rect 52425 2615 52625 2690
rect 52425 2575 52505 2615
rect 52545 2575 52625 2615
rect 52425 2490 52625 2575
rect 52775 2615 52975 2690
rect 52775 2575 52855 2615
rect 52895 2575 52975 2615
rect 52775 2490 52975 2575
rect 53125 2615 53325 2690
rect 53125 2575 53205 2615
rect 53245 2575 53325 2615
rect 53125 2490 53325 2575
rect 53475 2615 53675 2690
rect 53475 2575 53555 2615
rect 53595 2575 53675 2615
rect 53475 2490 53675 2575
rect 53825 2615 54025 2690
rect 53825 2575 53905 2615
rect 53945 2575 54025 2615
rect 53825 2490 54025 2575
rect 59775 2615 59975 2690
rect 59775 2575 59855 2615
rect 59895 2575 59975 2615
rect 59775 2490 59975 2575
rect 60125 2615 60325 2690
rect 60125 2575 60205 2615
rect 60245 2575 60325 2615
rect 60125 2490 60325 2575
rect 60475 2615 60675 2690
rect 60475 2575 60555 2615
rect 60595 2575 60675 2615
rect 60475 2490 60675 2575
rect 60825 2615 61025 2690
rect 60825 2575 60905 2615
rect 60945 2575 61025 2615
rect 60825 2490 61025 2575
rect 61175 2615 61375 2690
rect 61175 2575 61255 2615
rect 61295 2575 61375 2615
rect 61175 2490 61375 2575
rect 52425 2265 52625 2340
rect 52425 2225 52505 2265
rect 52545 2225 52625 2265
rect 52425 2140 52625 2225
rect 52775 2265 52975 2340
rect 52775 2225 52855 2265
rect 52895 2225 52975 2265
rect 52775 2140 52975 2225
rect 53125 2265 53325 2340
rect 53125 2225 53205 2265
rect 53245 2225 53325 2265
rect 53125 2140 53325 2225
rect 53475 2265 53675 2340
rect 53475 2225 53555 2265
rect 53595 2225 53675 2265
rect 53475 2140 53675 2225
rect 53825 2265 54025 2340
rect 53825 2225 53905 2265
rect 53945 2225 54025 2265
rect 53825 2140 54025 2225
rect 59775 2265 59975 2340
rect 59775 2225 59855 2265
rect 59895 2225 59975 2265
rect 59775 2140 59975 2225
rect 60125 2265 60325 2340
rect 60125 2225 60205 2265
rect 60245 2225 60325 2265
rect 60125 2140 60325 2225
rect 60475 2265 60675 2340
rect 60475 2225 60555 2265
rect 60595 2225 60675 2265
rect 60475 2140 60675 2225
rect 60825 2265 61025 2340
rect 60825 2225 60905 2265
rect 60945 2225 61025 2265
rect 60825 2140 61025 2225
rect 61175 2265 61375 2340
rect 61175 2225 61255 2265
rect 61295 2225 61375 2265
rect 61175 2140 61375 2225
rect 52425 1915 52625 1990
rect 52425 1875 52505 1915
rect 52545 1875 52625 1915
rect 52425 1790 52625 1875
rect 52775 1915 52975 1990
rect 52775 1875 52855 1915
rect 52895 1875 52975 1915
rect 52775 1790 52975 1875
rect 53125 1915 53325 1990
rect 53125 1875 53205 1915
rect 53245 1875 53325 1915
rect 53125 1790 53325 1875
rect 53475 1915 53675 1990
rect 53475 1875 53555 1915
rect 53595 1875 53675 1915
rect 53475 1790 53675 1875
rect 53825 1915 54025 1990
rect 53825 1875 53905 1915
rect 53945 1875 54025 1915
rect 53825 1790 54025 1875
rect 59775 1915 59975 1990
rect 59775 1875 59855 1915
rect 59895 1875 59975 1915
rect 59775 1790 59975 1875
rect 60125 1915 60325 1990
rect 60125 1875 60205 1915
rect 60245 1875 60325 1915
rect 60125 1790 60325 1875
rect 60475 1915 60675 1990
rect 60475 1875 60555 1915
rect 60595 1875 60675 1915
rect 60475 1790 60675 1875
rect 60825 1915 61025 1990
rect 60825 1875 60905 1915
rect 60945 1875 61025 1915
rect 60825 1790 61025 1875
rect 61175 1915 61375 1990
rect 61175 1875 61255 1915
rect 61295 1875 61375 1915
rect 61175 1790 61375 1875
rect 52425 1565 52625 1640
rect 52425 1525 52505 1565
rect 52545 1525 52625 1565
rect 52425 1440 52625 1525
rect 52775 1565 52975 1640
rect 52775 1525 52855 1565
rect 52895 1525 52975 1565
rect 52775 1440 52975 1525
rect 53125 1565 53325 1640
rect 53125 1525 53205 1565
rect 53245 1525 53325 1565
rect 53125 1440 53325 1525
rect 53475 1565 53675 1640
rect 53475 1525 53555 1565
rect 53595 1525 53675 1565
rect 53475 1440 53675 1525
rect 53825 1565 54025 1640
rect 53825 1525 53905 1565
rect 53945 1525 54025 1565
rect 53825 1440 54025 1525
rect 59775 1565 59975 1640
rect 59775 1525 59855 1565
rect 59895 1525 59975 1565
rect 59775 1440 59975 1525
rect 60125 1565 60325 1640
rect 60125 1525 60205 1565
rect 60245 1525 60325 1565
rect 60125 1440 60325 1525
rect 60475 1565 60675 1640
rect 60475 1525 60555 1565
rect 60595 1525 60675 1565
rect 60475 1440 60675 1525
rect 60825 1565 61025 1640
rect 60825 1525 60905 1565
rect 60945 1525 61025 1565
rect 60825 1440 61025 1525
rect 61175 1565 61375 1640
rect 61175 1525 61255 1565
rect 61295 1525 61375 1565
rect 61175 1440 61375 1525
rect 52425 1215 52625 1290
rect 52425 1175 52505 1215
rect 52545 1175 52625 1215
rect 52425 1090 52625 1175
rect 52775 1215 52975 1290
rect 52775 1175 52855 1215
rect 52895 1175 52975 1215
rect 52775 1090 52975 1175
rect 53125 1215 53325 1290
rect 53125 1175 53205 1215
rect 53245 1175 53325 1215
rect 53125 1090 53325 1175
rect 53475 1215 53675 1290
rect 53475 1175 53555 1215
rect 53595 1175 53675 1215
rect 53475 1090 53675 1175
rect 53825 1215 54025 1290
rect 53825 1175 53905 1215
rect 53945 1175 54025 1215
rect 53825 1090 54025 1175
rect 59775 1215 59975 1290
rect 59775 1175 59855 1215
rect 59895 1175 59975 1215
rect 59775 1090 59975 1175
rect 60125 1215 60325 1290
rect 60125 1175 60205 1215
rect 60245 1175 60325 1215
rect 60125 1090 60325 1175
rect 60475 1215 60675 1290
rect 60475 1175 60555 1215
rect 60595 1175 60675 1215
rect 60475 1090 60675 1175
rect 60825 1215 61025 1290
rect 60825 1175 60905 1215
rect 60945 1175 61025 1215
rect 60825 1090 61025 1175
rect 61175 1215 61375 1290
rect 61175 1175 61255 1215
rect 61295 1175 61375 1215
rect 61175 1090 61375 1175
rect 52425 865 52625 940
rect 52425 825 52505 865
rect 52545 825 52625 865
rect 52425 740 52625 825
rect 52775 865 52975 940
rect 52775 825 52855 865
rect 52895 825 52975 865
rect 52775 740 52975 825
rect 53125 865 53325 940
rect 53125 825 53205 865
rect 53245 825 53325 865
rect 53125 740 53325 825
rect 53475 865 53675 940
rect 53475 825 53555 865
rect 53595 825 53675 865
rect 53475 740 53675 825
rect 53825 865 54025 940
rect 53825 825 53905 865
rect 53945 825 54025 865
rect 53825 740 54025 825
rect 59775 865 59975 940
rect 59775 825 59855 865
rect 59895 825 59975 865
rect 59775 740 59975 825
rect 60125 865 60325 940
rect 60125 825 60205 865
rect 60245 825 60325 865
rect 60125 740 60325 825
rect 60475 865 60675 940
rect 60475 825 60555 865
rect 60595 825 60675 865
rect 60475 740 60675 825
rect 60825 865 61025 940
rect 60825 825 60905 865
rect 60945 825 61025 865
rect 60825 740 61025 825
rect 61175 865 61375 940
rect 61175 825 61255 865
rect 61295 825 61375 865
rect 61175 740 61375 825
rect 52425 515 52625 590
rect 52425 475 52505 515
rect 52545 475 52625 515
rect 52425 390 52625 475
rect 52775 515 52975 590
rect 52775 475 52855 515
rect 52895 475 52975 515
rect 52775 390 52975 475
rect 53125 515 53325 590
rect 53125 475 53205 515
rect 53245 475 53325 515
rect 53125 390 53325 475
rect 53475 515 53675 590
rect 53475 475 53555 515
rect 53595 475 53675 515
rect 53475 390 53675 475
rect 53825 515 54025 590
rect 53825 475 53905 515
rect 53945 475 54025 515
rect 53825 390 54025 475
rect 59775 515 59975 590
rect 59775 475 59855 515
rect 59895 475 59975 515
rect 59775 390 59975 475
rect 60125 515 60325 590
rect 60125 475 60205 515
rect 60245 475 60325 515
rect 60125 390 60325 475
rect 60475 515 60675 590
rect 60475 475 60555 515
rect 60595 475 60675 515
rect 60475 390 60675 475
rect 60825 515 61025 590
rect 60825 475 60905 515
rect 60945 475 61025 515
rect 60825 390 61025 475
rect 61175 515 61375 590
rect 61175 475 61255 515
rect 61295 475 61375 515
rect 61175 390 61375 475
rect 52425 165 52625 240
rect 52425 125 52505 165
rect 52545 125 52625 165
rect 52425 40 52625 125
rect 52775 165 52975 240
rect 52775 125 52855 165
rect 52895 125 52975 165
rect 52775 40 52975 125
rect 53125 165 53325 240
rect 53125 125 53205 165
rect 53245 125 53325 165
rect 53125 40 53325 125
rect 53475 165 53675 240
rect 53475 125 53555 165
rect 53595 125 53675 165
rect 53475 40 53675 125
rect 53825 165 54025 240
rect 53825 125 53905 165
rect 53945 125 54025 165
rect 53825 40 54025 125
rect 54175 165 54375 240
rect 54175 125 54255 165
rect 54295 125 54375 165
rect 54175 40 54375 125
rect 54525 165 54725 240
rect 54525 125 54605 165
rect 54645 125 54725 165
rect 54525 40 54725 125
rect 54875 165 55075 240
rect 54875 125 54955 165
rect 54995 125 55075 165
rect 54875 40 55075 125
rect 55225 165 55425 240
rect 55225 125 55305 165
rect 55345 125 55425 165
rect 55225 40 55425 125
rect 55575 165 55775 240
rect 55575 125 55655 165
rect 55695 125 55775 165
rect 55575 40 55775 125
rect 55925 165 56125 240
rect 55925 125 56005 165
rect 56045 125 56125 165
rect 55925 40 56125 125
rect 56275 165 56475 240
rect 56275 125 56355 165
rect 56395 125 56475 165
rect 56275 40 56475 125
rect 56625 165 56825 240
rect 56625 125 56705 165
rect 56745 125 56825 165
rect 56625 40 56825 125
rect 56975 165 57175 240
rect 56975 125 57055 165
rect 57095 125 57175 165
rect 56975 40 57175 125
rect 57325 165 57525 240
rect 57325 125 57405 165
rect 57445 125 57525 165
rect 57325 40 57525 125
rect 57675 165 57875 240
rect 57675 125 57755 165
rect 57795 125 57875 165
rect 57675 40 57875 125
rect 58025 165 58225 240
rect 58025 125 58105 165
rect 58145 125 58225 165
rect 58025 40 58225 125
rect 58375 165 58575 240
rect 58375 125 58455 165
rect 58495 125 58575 165
rect 58375 40 58575 125
rect 58725 165 58925 240
rect 58725 125 58805 165
rect 58845 125 58925 165
rect 58725 40 58925 125
rect 59075 165 59275 240
rect 59075 125 59155 165
rect 59195 125 59275 165
rect 59075 40 59275 125
rect 59425 165 59625 240
rect 59425 125 59505 165
rect 59545 125 59625 165
rect 59425 40 59625 125
rect 59775 165 59975 240
rect 59775 125 59855 165
rect 59895 125 59975 165
rect 59775 40 59975 125
rect 60125 165 60325 240
rect 60125 125 60205 165
rect 60245 125 60325 165
rect 60125 40 60325 125
rect 60475 165 60675 240
rect 60475 125 60555 165
rect 60595 125 60675 165
rect 60475 40 60675 125
rect 60825 165 61025 240
rect 60825 125 60905 165
rect 60945 125 61025 165
rect 60825 40 61025 125
rect 61175 165 61375 240
rect 61175 125 61255 165
rect 61295 125 61375 165
rect 61175 40 61375 125
rect 52425 -185 52625 -110
rect 52425 -225 52505 -185
rect 52545 -225 52625 -185
rect 52425 -310 52625 -225
rect 52775 -185 52975 -110
rect 52775 -225 52855 -185
rect 52895 -225 52975 -185
rect 52775 -310 52975 -225
rect 53125 -185 53325 -110
rect 53125 -225 53205 -185
rect 53245 -225 53325 -185
rect 53125 -310 53325 -225
rect 53475 -185 53675 -110
rect 53475 -225 53555 -185
rect 53595 -225 53675 -185
rect 53475 -310 53675 -225
rect 53825 -185 54025 -110
rect 53825 -225 53905 -185
rect 53945 -225 54025 -185
rect 53825 -310 54025 -225
rect 54175 -185 54375 -110
rect 54175 -225 54255 -185
rect 54295 -225 54375 -185
rect 54175 -310 54375 -225
rect 54525 -185 54725 -110
rect 54525 -225 54605 -185
rect 54645 -225 54725 -185
rect 54525 -310 54725 -225
rect 54875 -185 55075 -110
rect 54875 -225 54955 -185
rect 54995 -225 55075 -185
rect 54875 -310 55075 -225
rect 55225 -185 55425 -110
rect 55225 -225 55305 -185
rect 55345 -225 55425 -185
rect 55225 -310 55425 -225
rect 55575 -185 55775 -110
rect 55575 -225 55655 -185
rect 55695 -225 55775 -185
rect 55575 -310 55775 -225
rect 55925 -185 56125 -110
rect 55925 -225 56005 -185
rect 56045 -225 56125 -185
rect 55925 -310 56125 -225
rect 56275 -185 56475 -110
rect 56275 -225 56355 -185
rect 56395 -225 56475 -185
rect 56275 -310 56475 -225
rect 56625 -185 56825 -110
rect 56625 -225 56705 -185
rect 56745 -225 56825 -185
rect 56625 -310 56825 -225
rect 56975 -185 57175 -110
rect 56975 -225 57055 -185
rect 57095 -225 57175 -185
rect 56975 -310 57175 -225
rect 57325 -185 57525 -110
rect 57325 -225 57405 -185
rect 57445 -225 57525 -185
rect 57325 -310 57525 -225
rect 57675 -185 57875 -110
rect 57675 -225 57755 -185
rect 57795 -225 57875 -185
rect 57675 -310 57875 -225
rect 58025 -185 58225 -110
rect 58025 -225 58105 -185
rect 58145 -225 58225 -185
rect 58025 -310 58225 -225
rect 58375 -185 58575 -110
rect 58375 -225 58455 -185
rect 58495 -225 58575 -185
rect 58375 -310 58575 -225
rect 58725 -185 58925 -110
rect 58725 -225 58805 -185
rect 58845 -225 58925 -185
rect 58725 -310 58925 -225
rect 59075 -185 59275 -110
rect 59075 -225 59155 -185
rect 59195 -225 59275 -185
rect 59075 -310 59275 -225
rect 59425 -185 59625 -110
rect 59425 -225 59505 -185
rect 59545 -225 59625 -185
rect 59425 -310 59625 -225
rect 59775 -185 59975 -110
rect 59775 -225 59855 -185
rect 59895 -225 59975 -185
rect 59775 -310 59975 -225
rect 60125 -185 60325 -110
rect 60125 -225 60205 -185
rect 60245 -225 60325 -185
rect 60125 -310 60325 -225
rect 60475 -185 60675 -110
rect 60475 -225 60555 -185
rect 60595 -225 60675 -185
rect 60475 -310 60675 -225
rect 60825 -185 61025 -110
rect 60825 -225 60905 -185
rect 60945 -225 61025 -185
rect 60825 -310 61025 -225
rect 61175 -185 61375 -110
rect 61175 -225 61255 -185
rect 61295 -225 61375 -185
rect 61175 -310 61375 -225
<< mimcapcontact >>
rect 52505 5725 52545 5765
rect 52855 5725 52895 5765
rect 53205 5725 53245 5765
rect 53555 5725 53595 5765
rect 53905 5725 53945 5765
rect 54255 5725 54295 5765
rect 54605 5725 54645 5765
rect 54955 5725 54995 5765
rect 55305 5725 55345 5765
rect 55655 5725 55695 5765
rect 56005 5725 56045 5765
rect 56355 5725 56395 5765
rect 56705 5725 56745 5765
rect 57055 5725 57095 5765
rect 57405 5725 57445 5765
rect 57755 5725 57795 5765
rect 58105 5725 58145 5765
rect 58455 5725 58495 5765
rect 58805 5725 58845 5765
rect 59155 5725 59195 5765
rect 59505 5725 59545 5765
rect 59855 5725 59895 5765
rect 60205 5725 60245 5765
rect 60555 5725 60595 5765
rect 60905 5725 60945 5765
rect 61255 5725 61295 5765
rect 52505 5375 52545 5415
rect 52855 5375 52895 5415
rect 53205 5375 53245 5415
rect 53555 5375 53595 5415
rect 53905 5375 53945 5415
rect 54255 5375 54295 5415
rect 54605 5375 54645 5415
rect 54955 5375 54995 5415
rect 55305 5375 55345 5415
rect 55655 5375 55695 5415
rect 56005 5375 56045 5415
rect 56355 5375 56395 5415
rect 56705 5375 56745 5415
rect 57055 5375 57095 5415
rect 57405 5375 57445 5415
rect 57755 5375 57795 5415
rect 58105 5375 58145 5415
rect 58455 5375 58495 5415
rect 58805 5375 58845 5415
rect 59155 5375 59195 5415
rect 59505 5375 59545 5415
rect 59855 5375 59895 5415
rect 60205 5375 60245 5415
rect 60555 5375 60595 5415
rect 60905 5375 60945 5415
rect 61255 5375 61295 5415
rect 52505 5025 52545 5065
rect 52855 5025 52895 5065
rect 53205 5025 53245 5065
rect 53555 5025 53595 5065
rect 53905 5025 53945 5065
rect 54255 5025 54295 5065
rect 54605 5025 54645 5065
rect 54955 5025 54995 5065
rect 55305 5025 55345 5065
rect 55655 5015 55695 5055
rect 56005 5015 56045 5055
rect 56355 5015 56395 5055
rect 56705 5015 56745 5055
rect 57055 5015 57095 5055
rect 57405 5015 57445 5055
rect 57755 5015 57795 5055
rect 58105 5015 58145 5055
rect 58455 5025 58495 5065
rect 58805 5025 58845 5065
rect 59155 5025 59195 5065
rect 59505 5025 59545 5065
rect 59855 5025 59895 5065
rect 60205 5025 60245 5065
rect 60555 5025 60595 5065
rect 60905 5025 60945 5065
rect 61255 5025 61295 5065
rect 52505 4675 52545 4715
rect 52855 4675 52895 4715
rect 53205 4675 53245 4715
rect 53555 4675 53595 4715
rect 53905 4675 53945 4715
rect 54255 4675 54295 4715
rect 54605 4675 54645 4715
rect 54955 4675 54995 4715
rect 55305 4675 55345 4715
rect 58455 4675 58495 4715
rect 58805 4675 58845 4715
rect 59155 4675 59195 4715
rect 59505 4675 59545 4715
rect 59855 4675 59895 4715
rect 60205 4675 60245 4715
rect 60555 4675 60595 4715
rect 60905 4675 60945 4715
rect 61255 4675 61295 4715
rect 52505 4325 52545 4365
rect 52855 4325 52895 4365
rect 53205 4325 53245 4365
rect 53555 4325 53595 4365
rect 53905 4325 53945 4365
rect 54255 4325 54295 4365
rect 54605 4325 54645 4365
rect 54955 4325 54995 4365
rect 55305 4325 55345 4365
rect 58455 4325 58495 4365
rect 58805 4325 58845 4365
rect 59155 4325 59195 4365
rect 59505 4325 59545 4365
rect 59855 4325 59895 4365
rect 60205 4325 60245 4365
rect 60555 4325 60595 4365
rect 60905 4325 60945 4365
rect 61255 4325 61295 4365
rect 52505 3975 52545 4015
rect 52855 3975 52895 4015
rect 53205 3975 53245 4015
rect 53555 3975 53595 4015
rect 53905 3975 53945 4015
rect 59855 3975 59895 4015
rect 60205 3975 60245 4015
rect 60555 3975 60595 4015
rect 60905 3975 60945 4015
rect 61255 3975 61295 4015
rect 52505 3625 52545 3665
rect 52855 3625 52895 3665
rect 53205 3625 53245 3665
rect 53555 3625 53595 3665
rect 53905 3625 53945 3665
rect 59855 3625 59895 3665
rect 60205 3625 60245 3665
rect 60555 3625 60595 3665
rect 60905 3625 60945 3665
rect 61255 3625 61295 3665
rect 52505 3275 52545 3315
rect 52855 3275 52895 3315
rect 53205 3275 53245 3315
rect 53555 3275 53595 3315
rect 53905 3275 53945 3315
rect 59855 3275 59895 3315
rect 60205 3275 60245 3315
rect 60555 3275 60595 3315
rect 60905 3275 60945 3315
rect 61255 3275 61295 3315
rect 52505 2925 52545 2965
rect 52855 2925 52895 2965
rect 53205 2925 53245 2965
rect 53555 2925 53595 2965
rect 53905 2925 53945 2965
rect 59855 2925 59895 2965
rect 60205 2925 60245 2965
rect 60555 2925 60595 2965
rect 60905 2925 60945 2965
rect 61255 2925 61295 2965
rect 52505 2575 52545 2615
rect 52855 2575 52895 2615
rect 53205 2575 53245 2615
rect 53555 2575 53595 2615
rect 53905 2575 53945 2615
rect 59855 2575 59895 2615
rect 60205 2575 60245 2615
rect 60555 2575 60595 2615
rect 60905 2575 60945 2615
rect 61255 2575 61295 2615
rect 52505 2225 52545 2265
rect 52855 2225 52895 2265
rect 53205 2225 53245 2265
rect 53555 2225 53595 2265
rect 53905 2225 53945 2265
rect 59855 2225 59895 2265
rect 60205 2225 60245 2265
rect 60555 2225 60595 2265
rect 60905 2225 60945 2265
rect 61255 2225 61295 2265
rect 52505 1875 52545 1915
rect 52855 1875 52895 1915
rect 53205 1875 53245 1915
rect 53555 1875 53595 1915
rect 53905 1875 53945 1915
rect 59855 1875 59895 1915
rect 60205 1875 60245 1915
rect 60555 1875 60595 1915
rect 60905 1875 60945 1915
rect 61255 1875 61295 1915
rect 52505 1525 52545 1565
rect 52855 1525 52895 1565
rect 53205 1525 53245 1565
rect 53555 1525 53595 1565
rect 53905 1525 53945 1565
rect 59855 1525 59895 1565
rect 60205 1525 60245 1565
rect 60555 1525 60595 1565
rect 60905 1525 60945 1565
rect 61255 1525 61295 1565
rect 52505 1175 52545 1215
rect 52855 1175 52895 1215
rect 53205 1175 53245 1215
rect 53555 1175 53595 1215
rect 53905 1175 53945 1215
rect 59855 1175 59895 1215
rect 60205 1175 60245 1215
rect 60555 1175 60595 1215
rect 60905 1175 60945 1215
rect 61255 1175 61295 1215
rect 52505 825 52545 865
rect 52855 825 52895 865
rect 53205 825 53245 865
rect 53555 825 53595 865
rect 53905 825 53945 865
rect 59855 825 59895 865
rect 60205 825 60245 865
rect 60555 825 60595 865
rect 60905 825 60945 865
rect 61255 825 61295 865
rect 52505 475 52545 515
rect 52855 475 52895 515
rect 53205 475 53245 515
rect 53555 475 53595 515
rect 53905 475 53945 515
rect 59855 475 59895 515
rect 60205 475 60245 515
rect 60555 475 60595 515
rect 60905 475 60945 515
rect 61255 475 61295 515
rect 52505 125 52545 165
rect 52855 125 52895 165
rect 53205 125 53245 165
rect 53555 125 53595 165
rect 53905 125 53945 165
rect 54255 125 54295 165
rect 54605 125 54645 165
rect 54955 125 54995 165
rect 55305 125 55345 165
rect 55655 125 55695 165
rect 56005 125 56045 165
rect 56355 125 56395 165
rect 56705 125 56745 165
rect 57055 125 57095 165
rect 57405 125 57445 165
rect 57755 125 57795 165
rect 58105 125 58145 165
rect 58455 125 58495 165
rect 58805 125 58845 165
rect 59155 125 59195 165
rect 59505 125 59545 165
rect 59855 125 59895 165
rect 60205 125 60245 165
rect 60555 125 60595 165
rect 60905 125 60945 165
rect 61255 125 61295 165
rect 52505 -225 52545 -185
rect 52855 -225 52895 -185
rect 53205 -225 53245 -185
rect 53555 -225 53595 -185
rect 53905 -225 53945 -185
rect 54255 -225 54295 -185
rect 54605 -225 54645 -185
rect 54955 -225 54995 -185
rect 55305 -225 55345 -185
rect 55655 -225 55695 -185
rect 56005 -225 56045 -185
rect 56355 -225 56395 -185
rect 56705 -225 56745 -185
rect 57055 -225 57095 -185
rect 57405 -225 57445 -185
rect 57755 -225 57795 -185
rect 58105 -225 58145 -185
rect 58455 -225 58495 -185
rect 58805 -225 58845 -185
rect 59155 -225 59195 -185
rect 59505 -225 59545 -185
rect 59855 -225 59895 -185
rect 60205 -225 60245 -185
rect 60555 -225 60595 -185
rect 60905 -225 60945 -185
rect 61255 -225 61295 -185
<< metal4 >>
rect 51855 6190 61545 6195
rect 51855 6150 56880 6190
rect 56920 6150 61545 6190
rect 51855 6145 61545 6150
rect 52500 5765 53250 5770
rect 52500 5725 52505 5765
rect 52545 5725 52855 5765
rect 52895 5725 53205 5765
rect 53245 5725 53250 5765
rect 52500 5720 53250 5725
rect 53200 5420 53250 5720
rect 53550 5765 53600 5770
rect 53550 5725 53555 5765
rect 53595 5725 53600 5765
rect 53550 5420 53600 5725
rect 53900 5765 53950 5770
rect 53900 5725 53905 5765
rect 53945 5725 53950 5765
rect 53900 5420 53950 5725
rect 54250 5765 54300 5770
rect 54250 5725 54255 5765
rect 54295 5725 54300 5765
rect 54250 5420 54300 5725
rect 54600 5765 54650 5770
rect 54600 5725 54605 5765
rect 54645 5725 54650 5765
rect 54600 5420 54650 5725
rect 54950 5765 55000 5770
rect 54950 5725 54955 5765
rect 54995 5725 55000 5765
rect 54950 5420 55000 5725
rect 55300 5765 55350 5770
rect 55300 5725 55305 5765
rect 55345 5725 55350 5765
rect 55300 5420 55350 5725
rect 55650 5765 55700 5770
rect 55650 5725 55655 5765
rect 55695 5725 55700 5765
rect 55650 5420 55700 5725
rect 56000 5765 56050 5770
rect 56000 5725 56005 5765
rect 56045 5725 56050 5765
rect 56000 5420 56050 5725
rect 56350 5765 56400 5770
rect 56350 5725 56355 5765
rect 56395 5725 56400 5765
rect 56350 5420 56400 5725
rect 56700 5765 56750 5770
rect 56700 5725 56705 5765
rect 56745 5725 56750 5765
rect 56700 5420 56750 5725
rect 52500 5415 56750 5420
rect 52500 5375 52505 5415
rect 52545 5375 52855 5415
rect 52895 5375 53205 5415
rect 53245 5375 53555 5415
rect 53595 5375 53905 5415
rect 53945 5375 54255 5415
rect 54295 5375 54605 5415
rect 54645 5375 54955 5415
rect 54995 5375 55305 5415
rect 55345 5375 55655 5415
rect 55695 5375 56005 5415
rect 56045 5375 56355 5415
rect 56395 5375 56705 5415
rect 56745 5375 56750 5415
rect 52500 5370 56750 5375
rect 53200 5070 53250 5370
rect 52500 5065 53950 5070
rect 52500 5025 52505 5065
rect 52545 5025 52855 5065
rect 52895 5025 53205 5065
rect 53245 5025 53555 5065
rect 53595 5025 53905 5065
rect 53945 5025 53950 5065
rect 52500 5020 53950 5025
rect 54250 5065 54300 5370
rect 54250 5025 54255 5065
rect 54295 5025 54300 5065
rect 53200 4720 53250 5020
rect 52500 4715 53950 4720
rect 52500 4675 52505 4715
rect 52545 4675 52855 4715
rect 52895 4675 53205 4715
rect 53245 4675 53555 4715
rect 53595 4675 53905 4715
rect 53945 4675 53950 4715
rect 52500 4670 53950 4675
rect 54250 4715 54300 5025
rect 54250 4675 54255 4715
rect 54295 4675 54300 4715
rect 53200 4370 53250 4670
rect 52500 4365 53950 4370
rect 52500 4325 52505 4365
rect 52545 4325 52855 4365
rect 52895 4325 53205 4365
rect 53245 4325 53555 4365
rect 53595 4325 53905 4365
rect 53945 4325 53950 4365
rect 52500 4320 53950 4325
rect 54250 4365 54300 4675
rect 54250 4325 54255 4365
rect 54295 4325 54300 4365
rect 54250 4320 54300 4325
rect 54600 5065 54650 5370
rect 54600 5025 54605 5065
rect 54645 5025 54650 5065
rect 54600 4715 54650 5025
rect 54600 4675 54605 4715
rect 54645 4675 54650 4715
rect 54600 4365 54650 4675
rect 54600 4325 54605 4365
rect 54645 4325 54650 4365
rect 54600 4320 54650 4325
rect 54950 5065 55000 5370
rect 54950 5025 54955 5065
rect 54995 5025 55000 5065
rect 54950 4715 55000 5025
rect 54950 4675 54955 4715
rect 54995 4675 55000 4715
rect 54950 4365 55000 4675
rect 54950 4325 54955 4365
rect 54995 4325 55000 4365
rect 54950 4320 55000 4325
rect 55300 5065 55350 5370
rect 55300 5025 55305 5065
rect 55345 5025 55350 5065
rect 55300 4715 55350 5025
rect 55650 5055 55700 5370
rect 55650 5015 55655 5055
rect 55695 5015 55700 5055
rect 55650 5010 55700 5015
rect 56000 5055 56050 5370
rect 56000 5015 56005 5055
rect 56045 5015 56050 5055
rect 56000 5010 56050 5015
rect 56350 5055 56400 5370
rect 56350 5015 56355 5055
rect 56395 5015 56400 5055
rect 56350 5010 56400 5015
rect 56700 5055 56750 5370
rect 56700 5015 56705 5055
rect 56745 5015 56750 5055
rect 56700 5010 56750 5015
rect 57050 5765 57100 5770
rect 57050 5725 57055 5765
rect 57095 5725 57100 5765
rect 57050 5420 57100 5725
rect 57400 5765 57450 5770
rect 57400 5725 57405 5765
rect 57445 5725 57450 5765
rect 57400 5420 57450 5725
rect 57750 5765 57800 5770
rect 57750 5725 57755 5765
rect 57795 5725 57800 5765
rect 57750 5420 57800 5725
rect 58100 5765 58150 5770
rect 58100 5725 58105 5765
rect 58145 5725 58150 5765
rect 58100 5420 58150 5725
rect 58450 5765 58500 5770
rect 58450 5725 58455 5765
rect 58495 5725 58500 5765
rect 58450 5420 58500 5725
rect 58800 5765 58850 5770
rect 58800 5725 58805 5765
rect 58845 5725 58850 5765
rect 58800 5420 58850 5725
rect 59150 5765 59200 5770
rect 59150 5725 59155 5765
rect 59195 5725 59200 5765
rect 59150 5420 59200 5725
rect 59500 5765 59550 5770
rect 59500 5725 59505 5765
rect 59545 5725 59550 5765
rect 59500 5420 59550 5725
rect 59850 5765 59900 5770
rect 59850 5725 59855 5765
rect 59895 5725 59900 5765
rect 59850 5420 59900 5725
rect 60200 5765 60250 5770
rect 60200 5725 60205 5765
rect 60245 5725 60250 5765
rect 60200 5420 60250 5725
rect 60550 5765 61300 5770
rect 60550 5725 60555 5765
rect 60595 5725 60905 5765
rect 60945 5725 61255 5765
rect 61295 5725 61300 5765
rect 60550 5720 61300 5725
rect 60550 5420 60600 5720
rect 57050 5415 61300 5420
rect 57050 5375 57055 5415
rect 57095 5375 57405 5415
rect 57445 5375 57755 5415
rect 57795 5375 58105 5415
rect 58145 5375 58455 5415
rect 58495 5375 58805 5415
rect 58845 5375 59155 5415
rect 59195 5375 59505 5415
rect 59545 5375 59855 5415
rect 59895 5375 60205 5415
rect 60245 5375 60555 5415
rect 60595 5375 60905 5415
rect 60945 5375 61255 5415
rect 61295 5375 61300 5415
rect 57050 5370 61300 5375
rect 57050 5055 57100 5370
rect 57050 5015 57055 5055
rect 57095 5015 57100 5055
rect 57050 5010 57100 5015
rect 57400 5055 57450 5370
rect 57400 5015 57405 5055
rect 57445 5015 57450 5055
rect 57400 5010 57450 5015
rect 57750 5055 57800 5370
rect 57750 5015 57755 5055
rect 57795 5015 57800 5055
rect 57750 5010 57800 5015
rect 58100 5055 58150 5370
rect 58100 5015 58105 5055
rect 58145 5015 58150 5055
rect 58100 5010 58150 5015
rect 58450 5065 58500 5370
rect 58450 5025 58455 5065
rect 58495 5025 58500 5065
rect 55300 4675 55305 4715
rect 55345 4675 55350 4715
rect 55300 4365 55350 4675
rect 55300 4325 55305 4365
rect 55345 4325 55350 4365
rect 55300 4320 55350 4325
rect 58450 4715 58500 5025
rect 58450 4675 58455 4715
rect 58495 4675 58500 4715
rect 58450 4365 58500 4675
rect 58450 4325 58455 4365
rect 58495 4325 58500 4365
rect 58450 4320 58500 4325
rect 58800 5065 58850 5370
rect 58800 5025 58805 5065
rect 58845 5025 58850 5065
rect 58800 4715 58850 5025
rect 58800 4675 58805 4715
rect 58845 4675 58850 4715
rect 58800 4365 58850 4675
rect 58800 4325 58805 4365
rect 58845 4325 58850 4365
rect 58800 4320 58850 4325
rect 59150 5065 59200 5370
rect 59150 5025 59155 5065
rect 59195 5025 59200 5065
rect 59150 4715 59200 5025
rect 59150 4675 59155 4715
rect 59195 4675 59200 4715
rect 59150 4365 59200 4675
rect 59150 4325 59155 4365
rect 59195 4325 59200 4365
rect 59150 4320 59200 4325
rect 59500 5065 59550 5370
rect 60550 5070 60600 5370
rect 59500 5025 59505 5065
rect 59545 5025 59550 5065
rect 59500 4715 59550 5025
rect 59850 5065 61300 5070
rect 59850 5025 59855 5065
rect 59895 5025 60205 5065
rect 60245 5025 60555 5065
rect 60595 5025 60905 5065
rect 60945 5025 61255 5065
rect 61295 5025 61300 5065
rect 59850 5020 61300 5025
rect 60550 4720 60600 5020
rect 59500 4675 59505 4715
rect 59545 4675 59550 4715
rect 59500 4365 59550 4675
rect 59850 4715 61300 4720
rect 59850 4675 59855 4715
rect 59895 4675 60205 4715
rect 60245 4675 60555 4715
rect 60595 4675 60905 4715
rect 60945 4675 61255 4715
rect 61295 4675 61300 4715
rect 59850 4670 61300 4675
rect 60550 4370 60600 4670
rect 59500 4325 59505 4365
rect 59545 4325 59550 4365
rect 59500 4320 59550 4325
rect 59850 4365 61300 4370
rect 59850 4325 59855 4365
rect 59895 4325 60205 4365
rect 60245 4325 60555 4365
rect 60595 4325 60905 4365
rect 60945 4325 61255 4365
rect 61295 4325 61300 4365
rect 59850 4320 61300 4325
rect 53200 4020 53250 4320
rect 60550 4020 60600 4320
rect 52500 4015 53950 4020
rect 52500 3975 52505 4015
rect 52545 3975 52855 4015
rect 52895 3975 53205 4015
rect 53245 3975 53555 4015
rect 53595 3975 53905 4015
rect 53945 3975 53950 4015
rect 52500 3970 53950 3975
rect 59850 4015 61300 4020
rect 59850 3975 59855 4015
rect 59895 3975 60205 4015
rect 60245 3975 60555 4015
rect 60595 3975 60905 4015
rect 60945 3975 61255 4015
rect 61295 3975 61300 4015
rect 59850 3970 61300 3975
rect 53200 3670 53250 3970
rect 60550 3670 60600 3970
rect 52500 3665 53950 3670
rect 52500 3625 52505 3665
rect 52545 3625 52855 3665
rect 52895 3625 53205 3665
rect 53245 3625 53555 3665
rect 53595 3625 53905 3665
rect 53945 3625 53950 3665
rect 52500 3620 53950 3625
rect 59850 3665 61300 3670
rect 59850 3625 59855 3665
rect 59895 3625 60205 3665
rect 60245 3625 60555 3665
rect 60595 3625 60905 3665
rect 60945 3625 61255 3665
rect 61295 3625 61300 3665
rect 59850 3620 61300 3625
rect 53200 3320 53250 3620
rect 60550 3320 60600 3620
rect 52500 3315 53950 3320
rect 52500 3275 52505 3315
rect 52545 3275 52855 3315
rect 52895 3275 53205 3315
rect 53245 3275 53555 3315
rect 53595 3275 53905 3315
rect 53945 3275 53950 3315
rect 52500 3270 53950 3275
rect 59850 3315 61300 3320
rect 59850 3275 59855 3315
rect 59895 3275 60205 3315
rect 60245 3275 60555 3315
rect 60595 3275 60905 3315
rect 60945 3275 61255 3315
rect 61295 3275 61300 3315
rect 59850 3270 61300 3275
rect 53200 2970 53250 3270
rect 60550 2970 60600 3270
rect 52500 2965 53950 2970
rect 52500 2925 52505 2965
rect 52545 2925 52855 2965
rect 52895 2925 53205 2965
rect 53245 2925 53555 2965
rect 53595 2925 53905 2965
rect 53945 2925 53950 2965
rect 52500 2920 53950 2925
rect 59850 2965 61300 2970
rect 59850 2925 59855 2965
rect 59895 2925 60205 2965
rect 60245 2925 60555 2965
rect 60595 2925 60905 2965
rect 60945 2925 61255 2965
rect 61295 2925 61300 2965
rect 59850 2920 61300 2925
rect 53200 2620 53250 2920
rect 60550 2620 60600 2920
rect 52500 2615 53950 2620
rect 52500 2575 52505 2615
rect 52545 2575 52855 2615
rect 52895 2575 53205 2615
rect 53245 2575 53555 2615
rect 53595 2575 53905 2615
rect 53945 2575 53950 2615
rect 52500 2570 53950 2575
rect 59850 2615 61300 2620
rect 59850 2575 59855 2615
rect 59895 2575 60205 2615
rect 60245 2575 60555 2615
rect 60595 2575 60905 2615
rect 60945 2575 61255 2615
rect 61295 2575 61300 2615
rect 59850 2570 61300 2575
rect 53200 2270 53250 2570
rect 60550 2270 60600 2570
rect 52500 2265 53950 2270
rect 52500 2225 52505 2265
rect 52545 2225 52855 2265
rect 52895 2225 53205 2265
rect 53245 2225 53555 2265
rect 53595 2225 53905 2265
rect 53945 2225 53950 2265
rect 52500 2220 53950 2225
rect 59850 2265 61300 2270
rect 59850 2225 59855 2265
rect 59895 2225 60205 2265
rect 60245 2225 60555 2265
rect 60595 2225 60905 2265
rect 60945 2225 61255 2265
rect 61295 2225 61300 2265
rect 59850 2220 61300 2225
rect 53200 1920 53250 2220
rect 60550 1920 60600 2220
rect 52500 1915 54340 1920
rect 52500 1875 52505 1915
rect 52545 1875 52855 1915
rect 52895 1875 53205 1915
rect 53245 1875 53555 1915
rect 53595 1875 53905 1915
rect 53945 1875 54295 1915
rect 54335 1875 54340 1915
rect 52500 1870 54340 1875
rect 59460 1915 61300 1920
rect 59460 1875 59465 1915
rect 59505 1875 59855 1915
rect 59895 1875 60205 1915
rect 60245 1875 60555 1915
rect 60595 1875 60905 1915
rect 60945 1875 61255 1915
rect 61295 1875 61300 1915
rect 59460 1870 61300 1875
rect 53200 1570 53250 1870
rect 60550 1570 60600 1870
rect 52500 1565 53950 1570
rect 52500 1525 52505 1565
rect 52545 1525 52855 1565
rect 52895 1525 53205 1565
rect 53245 1525 53555 1565
rect 53595 1525 53905 1565
rect 53945 1525 53950 1565
rect 52500 1520 53950 1525
rect 59850 1565 61300 1570
rect 59850 1525 59855 1565
rect 59895 1525 60205 1565
rect 60245 1525 60555 1565
rect 60595 1525 60905 1565
rect 60945 1525 61255 1565
rect 61295 1525 61300 1565
rect 59850 1520 61300 1525
rect 53200 1220 53250 1520
rect 60550 1220 60600 1520
rect 52500 1215 53950 1220
rect 52500 1175 52505 1215
rect 52545 1175 52855 1215
rect 52895 1175 53205 1215
rect 53245 1175 53555 1215
rect 53595 1175 53905 1215
rect 53945 1175 53950 1215
rect 52500 1170 53950 1175
rect 59850 1215 61300 1220
rect 59850 1175 59855 1215
rect 59895 1175 60205 1215
rect 60245 1175 60555 1215
rect 60595 1175 60905 1215
rect 60945 1175 61255 1215
rect 61295 1175 61300 1215
rect 59850 1170 61300 1175
rect 53200 870 53250 1170
rect 60550 870 60600 1170
rect 52500 865 53950 870
rect 52500 825 52505 865
rect 52545 825 52855 865
rect 52895 825 53205 865
rect 53245 825 53555 865
rect 53595 825 53905 865
rect 53945 825 53950 865
rect 52500 820 53950 825
rect 59850 865 61300 870
rect 59850 825 59855 865
rect 59895 825 60205 865
rect 60245 825 60555 865
rect 60595 825 60905 865
rect 60945 825 61255 865
rect 61295 825 61300 865
rect 59850 820 61300 825
rect 53200 520 53250 820
rect 60550 520 60600 820
rect 52500 515 53950 520
rect 52500 475 52505 515
rect 52545 475 52855 515
rect 52895 475 53205 515
rect 53245 475 53555 515
rect 53595 475 53905 515
rect 53945 475 53950 515
rect 52500 470 53950 475
rect 59850 515 61300 520
rect 59850 475 59855 515
rect 59895 475 60205 515
rect 60245 475 60555 515
rect 60595 475 60905 515
rect 60945 475 61255 515
rect 61295 475 61300 515
rect 59850 470 61300 475
rect 53200 170 53250 470
rect 60550 170 60600 470
rect 52500 165 56750 170
rect 52500 125 52505 165
rect 52545 125 52855 165
rect 52895 125 53205 165
rect 53245 125 53555 165
rect 53595 125 53905 165
rect 53945 125 54255 165
rect 54295 125 54605 165
rect 54645 125 54955 165
rect 54995 125 55305 165
rect 55345 125 55655 165
rect 55695 125 56005 165
rect 56045 125 56355 165
rect 56395 125 56705 165
rect 56745 125 56750 165
rect 52500 120 56750 125
rect 53200 -180 53250 120
rect 52500 -185 53250 -180
rect 52500 -225 52505 -185
rect 52545 -225 52855 -185
rect 52895 -225 53205 -185
rect 53245 -225 53250 -185
rect 52500 -230 53250 -225
rect 53550 -185 53600 120
rect 53550 -225 53555 -185
rect 53595 -225 53600 -185
rect 53550 -230 53600 -225
rect 53900 -185 53950 120
rect 53900 -225 53905 -185
rect 53945 -225 53950 -185
rect 53900 -230 53950 -225
rect 54250 -185 54300 120
rect 54250 -225 54255 -185
rect 54295 -225 54300 -185
rect 54250 -230 54300 -225
rect 54600 -185 54650 120
rect 54600 -225 54605 -185
rect 54645 -225 54650 -185
rect 54600 -230 54650 -225
rect 54950 -185 55000 120
rect 54950 -225 54955 -185
rect 54995 -225 55000 -185
rect 54950 -230 55000 -225
rect 55300 -185 55350 120
rect 55300 -225 55305 -185
rect 55345 -225 55350 -185
rect 55300 -230 55350 -225
rect 55650 -185 55700 120
rect 55650 -225 55655 -185
rect 55695 -225 55700 -185
rect 55650 -230 55700 -225
rect 56000 -185 56050 120
rect 56000 -225 56005 -185
rect 56045 -225 56050 -185
rect 56000 -230 56050 -225
rect 56350 -185 56400 120
rect 56350 -225 56355 -185
rect 56395 -225 56400 -185
rect 56350 -230 56400 -225
rect 56700 -185 56750 120
rect 56700 -225 56705 -185
rect 56745 -225 56750 -185
rect 56700 -230 56750 -225
rect 57050 165 61300 170
rect 57050 125 57055 165
rect 57095 125 57405 165
rect 57445 125 57755 165
rect 57795 125 58105 165
rect 58145 125 58455 165
rect 58495 125 58805 165
rect 58845 125 59155 165
rect 59195 125 59505 165
rect 59545 125 59855 165
rect 59895 125 60205 165
rect 60245 125 60555 165
rect 60595 125 60905 165
rect 60945 125 61255 165
rect 61295 125 61300 165
rect 57050 120 61300 125
rect 57050 -185 57100 120
rect 57050 -225 57055 -185
rect 57095 -225 57100 -185
rect 57050 -230 57100 -225
rect 57400 -185 57450 120
rect 57400 -225 57405 -185
rect 57445 -225 57450 -185
rect 57400 -230 57450 -225
rect 57750 -185 57800 120
rect 57750 -225 57755 -185
rect 57795 -225 57800 -185
rect 57750 -230 57800 -225
rect 58100 -185 58150 120
rect 58100 -225 58105 -185
rect 58145 -225 58150 -185
rect 58100 -230 58150 -225
rect 58450 -185 58500 120
rect 58450 -225 58455 -185
rect 58495 -225 58500 -185
rect 58450 -230 58500 -225
rect 58800 -185 58850 120
rect 58800 -225 58805 -185
rect 58845 -225 58850 -185
rect 58800 -230 58850 -225
rect 59150 -185 59200 120
rect 59150 -225 59155 -185
rect 59195 -225 59200 -185
rect 59150 -230 59200 -225
rect 59500 -185 59550 120
rect 59500 -225 59505 -185
rect 59545 -225 59550 -185
rect 59500 -230 59550 -225
rect 59850 -185 59900 120
rect 59850 -225 59855 -185
rect 59895 -225 59900 -185
rect 59850 -230 59900 -225
rect 60200 -185 60250 120
rect 60200 -225 60205 -185
rect 60245 -225 60250 -185
rect 60200 -230 60250 -225
rect 60550 -180 60600 120
rect 60550 -185 61300 -180
rect 60550 -225 60555 -185
rect 60595 -225 60905 -185
rect 60945 -225 61255 -185
rect 61295 -225 61300 -185
rect 60550 -230 61300 -225
rect 51855 -510 61545 -505
rect 51855 -550 56880 -510
rect 56920 -550 61545 -510
rect 51855 -555 61545 -550
<< labels >>
flabel metal4 51855 6170 51855 6170 7 FreeSans 800 0 -400 0 VDDA
port 1 w
flabel metal3 59195 3460 59195 3460 3 FreeSans 240 0 80 0 cap_res_X
flabel metal3 54605 3460 54605 3460 7 FreeSans 240 0 -80 0 cap_res_Y
flabel metal4 51855 -530 51855 -530 7 FreeSans 800 0 -400 0 GNDA
port 16 w
flabel metal1 56910 1290 56910 1290 3 FreeSans 200 0 80 0 V_p_mir
flabel metal1 56370 1880 56370 1880 7 FreeSans 240 0 -80 0 VD2
flabel metal1 57430 1875 57430 1875 3 FreeSans 240 0 80 0 VD1
flabel metal2 57720 1300 57720 1300 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal2 57365 4810 57365 4810 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 56455 4810 56455 4810 1 FreeSans 240 0 0 80 Vb2_2
flabel metal1 57220 1285 57220 1285 3 FreeSans 240 0 80 0 V_source
flabel metal1 59485 1170 59485 1170 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 58975 1900 58975 1900 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal2 57000 3515 57000 3515 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56855 3550 56855 3550 5 FreeSans 200 0 0 -80 Vb2
port 5 s
flabel metal2 57865 3660 57865 3660 5 FreeSans 240 0 0 -80 VD3
flabel metal2 55910 3660 55910 3660 5 FreeSans 240 0 0 -80 VD4
flabel metal2 55980 1770 55980 1770 7 FreeSans 240 0 -80 0 VIN+
port 14 w
flabel metal2 57820 1770 57820 1770 3 FreeSans 240 0 80 0 VIN-
port 15 e
flabel metal2 57605 2880 57605 2880 3 FreeSans 200 0 80 0 err_amp_mir
flabel metal2 56900 3065 56900 3065 1 FreeSans 240 0 0 80 V_tot
flabel metal2 57580 2710 57580 2710 5 FreeSans 240 0 0 -80 err_amp_out
flabel metal2 55955 2825 55955 2825 7 FreeSans 200 0 -80 0 V_err_amp_ref
port 12 w
flabel metal1 57455 2625 57455 2625 7 FreeSans 240 0 -80 0 X
flabel metal1 59020 2205 59020 2205 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 54315 1170 54315 1170 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal1 54825 1900 54825 1900 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal1 54780 2205 54780 2205 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 56345 2625 56345 2625 3 FreeSans 240 0 80 0 Y
flabel metal1 57650 3195 57650 3195 3 FreeSans 200 0 80 0 V_err_p
flabel metal1 56140 3240 56140 3240 7 FreeSans 240 0 -80 0 V_er_mir_p
flabel metal1 56795 3145 56795 3145 7 FreeSans 200 0 -80 0 V_err_gate
port 13 w
flabel metal2 56835 515 56835 515 5 FreeSans 240 0 0 -80 Vb1_2
flabel metal1 56955 1810 56955 1810 7 FreeSans 240 0 -80 0 V_tail_gate
port 11 w
flabel metal1 57980 2250 57980 2250 1 FreeSans 200 0 0 80 Vb1
port 6 n
<< end >>
