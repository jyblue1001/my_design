magic
tech sky130A
timestamp 1722810130
<< nwell >>
rect -40 205 170 515
<< nmos >>
rect 30 50 45 150
rect 85 50 100 150
<< pmos >>
rect 30 225 45 425
rect 85 225 100 425
<< ndiff >>
rect -20 130 30 150
rect -20 110 -5 130
rect 15 110 30 130
rect -20 90 30 110
rect -20 70 -5 90
rect 15 70 30 90
rect -20 50 30 70
rect 45 50 85 150
rect 100 130 150 150
rect 100 110 115 130
rect 135 110 150 130
rect 100 90 150 110
rect 100 70 115 90
rect 135 70 150 90
rect 100 50 150 70
<< pdiff >>
rect -20 405 30 425
rect -20 385 -5 405
rect 15 385 30 405
rect -20 360 30 385
rect -20 340 -5 360
rect 15 340 30 360
rect -20 315 30 340
rect -20 295 -5 315
rect 15 295 30 315
rect -20 265 30 295
rect -20 245 -5 265
rect 15 245 30 265
rect -20 225 30 245
rect 45 405 85 425
rect 45 385 55 405
rect 75 385 85 405
rect 45 360 85 385
rect 45 340 55 360
rect 75 340 85 360
rect 45 315 85 340
rect 45 295 55 315
rect 75 295 85 315
rect 45 265 85 295
rect 45 245 55 265
rect 75 245 85 265
rect 45 225 85 245
rect 100 405 150 425
rect 100 385 115 405
rect 135 385 150 405
rect 100 360 150 385
rect 100 340 115 360
rect 135 340 150 360
rect 100 315 150 340
rect 100 295 115 315
rect 135 295 150 315
rect 100 265 150 295
rect 100 245 115 265
rect 135 245 150 265
rect 100 225 150 245
<< ndiffc >>
rect -5 110 15 130
rect -5 70 15 90
rect 115 110 135 130
rect 115 70 135 90
<< pdiffc >>
rect -5 385 15 405
rect -5 340 15 360
rect -5 295 15 315
rect -5 245 15 265
rect 55 385 75 405
rect 55 340 75 360
rect 55 295 75 315
rect 55 245 75 265
rect 115 385 135 405
rect 115 340 135 360
rect 115 295 135 315
rect 115 245 135 265
<< psubdiff >>
rect -20 10 150 20
rect -20 -10 -5 10
rect 15 -10 150 10
rect -20 -20 150 -10
<< nsubdiff >>
rect -20 485 150 495
rect -20 465 -5 485
rect 15 465 55 485
rect 75 465 115 485
rect 135 465 150 485
rect -20 455 150 465
<< psubdiffcont >>
rect -5 -10 15 10
<< nsubdiffcont >>
rect -5 465 15 485
rect 55 465 75 485
rect 115 465 135 485
<< poly >>
rect 30 425 45 440
rect 85 425 100 440
rect 30 200 45 225
rect -10 190 45 200
rect -10 170 0 190
rect 20 170 45 190
rect -10 160 45 170
rect 30 150 45 160
rect 85 200 100 225
rect 85 190 140 200
rect 85 170 110 190
rect 130 170 140 190
rect 85 160 140 170
rect 85 150 100 160
rect 30 35 45 50
rect 85 35 100 50
<< polycont >>
rect 0 170 20 190
rect 110 170 130 190
<< locali >>
rect -10 525 20 530
rect -10 505 -5 525
rect 15 505 20 525
rect -10 485 20 505
rect -10 465 -5 485
rect 15 465 20 485
rect -10 405 20 465
rect -10 385 -5 405
rect 15 385 20 405
rect -10 360 20 385
rect -10 340 -5 360
rect 15 340 20 360
rect -10 315 20 340
rect -10 295 -5 315
rect 15 295 20 315
rect -10 265 20 295
rect -10 245 -5 265
rect 15 245 20 265
rect -10 235 20 245
rect 50 525 80 530
rect 50 505 55 525
rect 75 505 80 525
rect 50 485 80 505
rect 50 465 55 485
rect 75 465 80 485
rect 50 405 80 465
rect 50 385 55 405
rect 75 385 80 405
rect 50 360 80 385
rect 50 340 55 360
rect 75 340 80 360
rect 50 315 80 340
rect 50 295 55 315
rect 75 295 80 315
rect 50 265 80 295
rect 50 245 55 265
rect 75 245 80 265
rect -10 190 30 200
rect -10 170 0 190
rect 20 170 30 190
rect -10 160 30 170
rect 50 140 80 245
rect 110 525 140 530
rect 110 505 115 525
rect 135 505 140 525
rect 110 485 140 505
rect 110 465 115 485
rect 135 465 140 485
rect 110 405 140 465
rect 110 385 115 405
rect 135 385 140 405
rect 110 360 140 385
rect 110 340 115 360
rect 135 340 140 360
rect 110 315 140 340
rect 110 295 115 315
rect 135 295 140 315
rect 110 265 140 295
rect 110 245 115 265
rect 135 245 140 265
rect 110 235 140 245
rect 100 190 140 200
rect 100 170 110 190
rect 130 170 140 190
rect 100 160 140 170
rect -10 130 20 140
rect -10 110 -5 130
rect 15 110 20 130
rect -10 90 20 110
rect -10 70 -5 90
rect 15 70 20 90
rect -10 60 20 70
rect 50 130 140 140
rect 50 110 115 130
rect 135 110 140 130
rect 50 90 140 110
rect 50 70 115 90
rect 135 70 140 90
rect 50 60 140 70
rect -5 10 15 60
rect -10 -25 20 -10
rect -10 -30 140 -25
rect -10 -50 -5 -30
rect 15 -50 55 -30
rect 75 -50 115 -30
rect 135 -50 140 -30
rect -10 -55 140 -50
<< viali >>
rect -5 505 15 525
rect 55 505 75 525
rect 115 505 135 525
rect -5 -50 15 -30
rect 55 -50 75 -30
rect 115 -50 135 -30
<< metal1 >>
rect -20 525 150 535
rect -20 505 -5 525
rect 15 505 55 525
rect 75 505 115 525
rect 135 505 150 525
rect -20 495 150 505
rect -20 -30 150 -20
rect -20 -50 -5 -30
rect 15 -50 55 -30
rect 75 -50 115 -30
rect 135 -50 150 -30
rect -20 -60 150 -50
<< end >>
