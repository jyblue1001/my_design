** sch_path: /foss/designs/my_design/projects/pll/full_pll/magic/tb_pfd_cp_lf_magic.sch
**.subckt tb_pfd_cp_lf_magic
V1 VDD GND 1.8
V2 F_REF GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
V3 F_VCO GND pulse(0 1.8 12ns 1ns 1ns 24ns 50ns)
I1 GND I_IN 100u
x1 V_OUT VDD GND F_REF F_VCO I_IN pfd_cp_lf_magic
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.include /foss/designs/my_design/projects/pll/full_pll/magic/pfd_cp_lf_magic.spice


.option method=gear
.option wnflag=1
.option savecurrents

* V_out initial voltage value for the F_VCO delay of 2ns  (leading)
* .ic v(v_out) = 1.8

* V_out initial voltage value for the F_VCO delay of 12ns (lock condition)
.ic v(v_out) = 0.9

* V_out initial voltage value for the F_VCO delay of 22ns (lagging)
* .ic v(v_out) = 0.0

.control
  save v(f_ref) save v(f_vco) save v(i_in) save v(up_pfd) v(down_pfd) v(up_pfd_b) v(down_pfd_b) v(up) v(up_b) v(down) v(down_b) v(x) v(opamp_out) v(up_input) v(down_input) v(down_gate) v(v_out)
  * save all

  * timestep for exact simulation results
  * tran 5ps 0.5us

  * timestep for faster simulation results
  tran 50ps 0.5us

  remzerovec
  write tb_pfd_cp_lf_magic_8.raw
  set appendwrite

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
