magic
tech sky130A
magscale 1 2
timestamp 1726264562
<< error_p >>
rect 2389 200 2390 201
rect 2390 199 2391 200
rect 2390 -210 2391 -209
rect 2389 -211 2390 -210
rect 250 -2190 251 -2189
rect 649 -2190 650 -2189
rect 249 -2191 250 -2190
rect 650 -2191 651 -2190
rect 1049 -3220 1050 -3219
rect 1450 -3220 1451 -3219
rect 1050 -3221 1051 -3220
rect 1449 -3221 1450 -3220
<< nmos >>
rect 0 200 2790 600
rect 2390 -210 2790 200
rect -10 -610 2790 -210
rect -150 -2190 1050 -1790
rect -150 -3650 250 -2190
rect 650 -3220 1050 -2190
rect 1450 -3220 1850 -1760
rect 650 -3620 1850 -3220
<< ndiff >>
rect -90 580 0 600
rect -90 220 -70 580
rect -30 220 0 580
rect -90 200 0 220
rect -110 -240 -10 -210
rect -110 -580 -80 -240
rect -40 -580 -10 -240
rect -110 -610 -10 -580
rect 1450 -1690 1850 -1660
rect 1450 -1730 1480 -1690
rect 1820 -1730 1850 -1690
rect 1450 -1760 1850 -1730
rect -150 -3680 250 -3650
rect -150 -3720 -130 -3680
rect 230 -3720 250 -3680
rect -150 -3740 250 -3720
<< ndiffc >>
rect -70 220 -30 580
rect -80 -580 -40 -240
rect 1480 -1730 1820 -1690
rect -130 -3720 230 -3680
<< psubdiff >>
rect -180 580 -90 600
rect -180 220 -150 580
rect -110 220 -90 580
rect -180 200 -90 220
rect -150 -3760 250 -3740
rect -150 -3800 -130 -3760
rect 230 -3800 250 -3760
rect -150 -3830 250 -3800
<< psubdiffcont >>
rect -150 220 -110 580
rect -130 -3800 230 -3760
<< poly >>
rect 0 600 2820 630
rect 0 170 2390 200
rect -10 -210 2390 170
rect 2790 -610 2820 600
rect -10 -640 2820 -610
rect -180 -1790 1450 -1760
rect -180 -3650 -150 -1790
rect 250 -3620 650 -2190
rect 1050 -3220 1450 -1790
rect 1850 -3620 1880 -1760
rect 250 -3650 1880 -3620
<< xpolycontact >>
rect 2770 -3034 2908 -2594
rect 2570 -3534 2708 -3094
rect 2570 -4080 2708 -3640
rect 2770 -4080 2908 -3640
<< xpolyres >>
rect 2570 -3640 2708 -3534
rect 2770 -3640 2908 -3034
<< locali >>
rect -170 580 -10 590
rect -170 220 -150 580
rect -110 220 -70 580
rect -30 220 -10 580
rect -170 210 -10 220
rect -100 -240 -20 -220
rect -100 -580 -80 -240
rect -40 -580 -20 -240
rect -100 -600 -20 -580
rect 1460 -1690 1840 -1670
rect 1460 -1730 1480 -1690
rect 1820 -1730 1840 -1690
rect 1460 -1750 1840 -1730
rect -140 -3680 240 -3660
rect -140 -3720 -130 -3680
rect 230 -3720 240 -3680
rect -140 -3760 240 -3720
rect -140 -3800 -130 -3760
rect 230 -3800 240 -3760
rect -140 -3820 240 -3800
<< end >>
