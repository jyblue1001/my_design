** sch_path: /foss/designs/my_design/projects/resistor/xschem_ngspice/resistor20k_xschem.sch
**.subckt resistor20k_xschem
XR2 bot top GND sky130_fd_pr__res_xhigh_po_0p35 L=3.5 mult=1 m=1
**.ends
.GLOBAL GND
.end
